module basic_3000_30000_3500_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_2395,In_1038);
nor U1 (N_1,In_2984,In_713);
or U2 (N_2,In_785,In_414);
nand U3 (N_3,In_483,In_1948);
nor U4 (N_4,In_2246,In_1529);
or U5 (N_5,In_2749,In_988);
and U6 (N_6,In_1440,In_1031);
nand U7 (N_7,In_2489,In_1154);
nand U8 (N_8,In_2173,In_1799);
and U9 (N_9,In_1410,In_2121);
xor U10 (N_10,In_1172,In_1383);
or U11 (N_11,In_2672,In_2095);
xnor U12 (N_12,In_2668,In_1545);
nand U13 (N_13,In_1804,In_2914);
and U14 (N_14,In_2480,In_407);
xor U15 (N_15,In_2429,In_2381);
xnor U16 (N_16,In_2196,In_976);
or U17 (N_17,In_1409,In_2431);
or U18 (N_18,In_2609,In_2306);
nor U19 (N_19,In_2796,In_1144);
nor U20 (N_20,In_1666,In_811);
xnor U21 (N_21,In_2459,In_2159);
nor U22 (N_22,In_646,In_2729);
nor U23 (N_23,In_2709,In_2278);
and U24 (N_24,In_651,In_1023);
nand U25 (N_25,In_2898,In_620);
nor U26 (N_26,In_2469,In_953);
xnor U27 (N_27,In_2276,In_1719);
and U28 (N_28,In_2531,In_2020);
nand U29 (N_29,In_1492,In_2849);
and U30 (N_30,In_2281,In_206);
or U31 (N_31,In_999,In_2228);
xor U32 (N_32,In_2236,In_700);
nand U33 (N_33,In_1504,In_1740);
or U34 (N_34,In_1761,In_1359);
and U35 (N_35,In_1485,In_222);
xor U36 (N_36,In_229,In_2058);
and U37 (N_37,In_2051,In_1380);
or U38 (N_38,In_1446,In_2873);
nand U39 (N_39,In_1803,In_319);
and U40 (N_40,In_1780,In_2837);
nand U41 (N_41,In_358,In_2474);
or U42 (N_42,In_2660,In_2897);
xor U43 (N_43,In_1341,In_317);
nor U44 (N_44,In_2086,In_303);
nand U45 (N_45,In_1551,In_115);
nor U46 (N_46,In_77,In_1113);
and U47 (N_47,In_1795,In_301);
nor U48 (N_48,In_964,In_415);
nand U49 (N_49,In_1094,In_476);
and U50 (N_50,In_2037,In_1473);
and U51 (N_51,In_2560,In_2230);
nand U52 (N_52,In_2985,In_799);
nor U53 (N_53,In_1942,In_2988);
and U54 (N_54,In_1552,In_1371);
nand U55 (N_55,In_2895,In_2846);
or U56 (N_56,In_1775,In_2357);
or U57 (N_57,In_83,In_1064);
and U58 (N_58,In_2225,In_2014);
and U59 (N_59,In_1107,In_1433);
nand U60 (N_60,In_2832,In_252);
xnor U61 (N_61,In_2030,In_2137);
nand U62 (N_62,In_548,In_1497);
and U63 (N_63,In_1053,In_1843);
and U64 (N_64,In_2915,In_1628);
xnor U65 (N_65,In_1702,In_1499);
xor U66 (N_66,In_2118,In_2199);
xor U67 (N_67,In_2272,In_2928);
nor U68 (N_68,In_2958,In_1845);
or U69 (N_69,In_2853,In_47);
nand U70 (N_70,In_436,In_170);
and U71 (N_71,In_1812,In_1862);
xnor U72 (N_72,In_2978,In_1970);
nand U73 (N_73,In_487,In_20);
or U74 (N_74,In_2178,In_2916);
and U75 (N_75,In_162,In_2601);
nand U76 (N_76,In_2691,In_2647);
or U77 (N_77,In_873,In_2102);
nor U78 (N_78,In_2383,In_519);
and U79 (N_79,In_89,In_575);
nor U80 (N_80,In_1721,In_2164);
nand U81 (N_81,In_1275,In_1486);
nand U82 (N_82,In_185,In_395);
nand U83 (N_83,In_372,In_2751);
nor U84 (N_84,In_2857,In_816);
nand U85 (N_85,In_177,In_2645);
or U86 (N_86,In_2420,In_1472);
nand U87 (N_87,In_2448,In_2167);
nor U88 (N_88,In_67,In_1432);
xnor U89 (N_89,In_614,In_709);
nand U90 (N_90,In_2778,In_1387);
nor U91 (N_91,In_585,In_545);
nand U92 (N_92,In_2467,In_1676);
nand U93 (N_93,In_2133,In_2976);
and U94 (N_94,In_2101,In_1561);
nor U95 (N_95,In_2680,In_2097);
or U96 (N_96,In_2863,In_1963);
xnor U97 (N_97,In_1006,In_1832);
xor U98 (N_98,In_2089,In_1568);
nor U99 (N_99,In_2920,In_2106);
xor U100 (N_100,In_1258,In_2659);
xnor U101 (N_101,In_797,In_1151);
or U102 (N_102,In_397,In_2033);
nand U103 (N_103,In_1419,In_2696);
nor U104 (N_104,In_608,In_2867);
xnor U105 (N_105,In_2463,In_335);
and U106 (N_106,In_537,In_2032);
nand U107 (N_107,In_2575,In_408);
xnor U108 (N_108,In_1962,In_69);
and U109 (N_109,In_2762,In_46);
nand U110 (N_110,In_2119,In_2152);
and U111 (N_111,In_778,In_2200);
or U112 (N_112,In_2226,In_648);
or U113 (N_113,In_2370,In_388);
nor U114 (N_114,In_1815,In_1806);
nand U115 (N_115,In_122,In_804);
nor U116 (N_116,In_171,In_2446);
nand U117 (N_117,In_662,In_425);
xnor U118 (N_118,In_793,In_2767);
or U119 (N_119,In_1018,In_2221);
nand U120 (N_120,In_2113,In_12);
nor U121 (N_121,In_239,In_924);
or U122 (N_122,In_1990,In_2845);
nand U123 (N_123,In_231,In_934);
nand U124 (N_124,In_2342,In_1536);
or U125 (N_125,In_1677,In_94);
nor U126 (N_126,In_952,In_1036);
nor U127 (N_127,In_580,In_2638);
nand U128 (N_128,In_1457,In_2124);
or U129 (N_129,In_2507,In_2002);
nor U130 (N_130,In_1496,In_2803);
and U131 (N_131,In_2585,In_589);
xnor U132 (N_132,In_2183,In_2184);
nand U133 (N_133,In_887,In_1967);
nor U134 (N_134,In_2695,In_1562);
and U135 (N_135,In_536,In_2170);
xor U136 (N_136,In_890,In_676);
and U137 (N_137,In_2304,In_2255);
and U138 (N_138,In_2974,In_2242);
xnor U139 (N_139,In_2703,In_769);
and U140 (N_140,In_2850,In_2372);
or U141 (N_141,In_2557,In_2670);
nand U142 (N_142,In_767,In_2082);
and U143 (N_143,In_2043,In_507);
and U144 (N_144,In_2589,In_1878);
nand U145 (N_145,In_325,In_1181);
nor U146 (N_146,In_195,In_2307);
nor U147 (N_147,In_1620,In_1959);
xnor U148 (N_148,In_50,In_1807);
nor U149 (N_149,In_2388,In_484);
xnor U150 (N_150,In_2112,In_1034);
nor U151 (N_151,In_312,In_1695);
and U152 (N_152,In_1136,In_403);
xor U153 (N_153,In_1746,In_2812);
nor U154 (N_154,In_2215,In_2117);
xnor U155 (N_155,In_2540,In_2176);
or U156 (N_156,In_764,In_2339);
nor U157 (N_157,In_1681,In_1789);
or U158 (N_158,In_1917,In_2192);
nand U159 (N_159,In_2235,In_1634);
or U160 (N_160,In_1764,In_1893);
and U161 (N_161,In_1625,In_2499);
xnor U162 (N_162,In_2375,In_967);
nand U163 (N_163,In_508,In_448);
nand U164 (N_164,In_1770,In_2493);
nor U165 (N_165,In_912,In_725);
or U166 (N_166,In_1621,In_2269);
or U167 (N_167,In_526,In_587);
and U168 (N_168,In_219,In_1667);
and U169 (N_169,In_1000,In_404);
nand U170 (N_170,In_1140,In_1032);
and U171 (N_171,In_2579,In_210);
nor U172 (N_172,In_2319,In_865);
xnor U173 (N_173,In_1402,In_1703);
nor U174 (N_174,In_1487,In_1542);
and U175 (N_175,In_204,In_2358);
nor U176 (N_176,In_2338,In_917);
and U177 (N_177,In_503,In_65);
nor U178 (N_178,In_732,In_2071);
nor U179 (N_179,In_169,In_2490);
nor U180 (N_180,In_2013,In_2678);
and U181 (N_181,In_704,In_2788);
nand U182 (N_182,In_1100,In_1960);
and U183 (N_183,In_1350,In_835);
nor U184 (N_184,In_842,In_1065);
xnor U185 (N_185,In_1295,In_1131);
or U186 (N_186,In_1846,In_1170);
or U187 (N_187,In_2041,In_362);
or U188 (N_188,In_2146,In_1459);
or U189 (N_189,In_1294,In_913);
or U190 (N_190,In_783,In_2742);
nand U191 (N_191,In_9,In_2361);
and U192 (N_192,In_1503,In_2053);
xnor U193 (N_193,In_2582,In_13);
and U194 (N_194,In_2295,In_1063);
xor U195 (N_195,In_559,In_2384);
nor U196 (N_196,In_2554,In_187);
and U197 (N_197,In_1632,In_2229);
nand U198 (N_198,In_2072,In_930);
nor U199 (N_199,In_352,In_2959);
nand U200 (N_200,In_45,In_125);
nand U201 (N_201,In_1523,In_1887);
nor U202 (N_202,In_2317,In_2658);
nor U203 (N_203,In_572,In_1161);
and U204 (N_204,In_1156,In_405);
or U205 (N_205,In_440,In_2181);
or U206 (N_206,In_624,In_394);
nand U207 (N_207,In_1995,In_647);
nor U208 (N_208,In_111,In_2539);
and U209 (N_209,In_1830,In_1668);
and U210 (N_210,In_2010,In_1439);
nor U211 (N_211,In_1554,In_1650);
nor U212 (N_212,In_324,In_933);
xnor U213 (N_213,In_1563,In_2801);
nand U214 (N_214,In_859,In_2387);
or U215 (N_215,In_2998,In_2379);
or U216 (N_216,In_546,In_492);
xnor U217 (N_217,In_1757,In_131);
xor U218 (N_218,In_2535,In_381);
and U219 (N_219,In_1927,In_406);
nor U220 (N_220,In_70,In_927);
nand U221 (N_221,In_1362,In_743);
nor U222 (N_222,In_1897,In_318);
or U223 (N_223,In_796,In_2441);
xor U224 (N_224,In_80,In_2016);
and U225 (N_225,In_1796,In_1854);
nand U226 (N_226,In_494,In_2909);
and U227 (N_227,In_1330,In_1193);
or U228 (N_228,In_1430,In_760);
and U229 (N_229,In_1567,In_1988);
or U230 (N_230,In_568,In_1139);
and U231 (N_231,In_2514,In_871);
xor U232 (N_232,In_858,In_1782);
or U233 (N_233,In_262,In_2926);
and U234 (N_234,In_1455,In_741);
nor U235 (N_235,In_260,In_2142);
and U236 (N_236,In_2881,In_322);
nand U237 (N_237,In_1794,In_2689);
and U238 (N_238,In_2508,In_2438);
nor U239 (N_239,In_2889,In_1543);
and U240 (N_240,In_954,In_284);
nor U241 (N_241,In_1838,In_2385);
or U242 (N_242,In_946,In_370);
nor U243 (N_243,In_416,In_1772);
and U244 (N_244,In_2028,In_1072);
xor U245 (N_245,In_2622,In_2313);
nand U246 (N_246,In_1394,In_1324);
and U247 (N_247,In_567,In_2649);
nor U248 (N_248,In_2066,In_1949);
and U249 (N_249,In_2818,In_1802);
or U250 (N_250,In_257,In_2412);
xor U251 (N_251,In_465,In_48);
xnor U252 (N_252,In_191,In_1207);
nand U253 (N_253,In_1048,In_1010);
or U254 (N_254,In_283,In_1743);
nor U255 (N_255,In_2210,In_1723);
and U256 (N_256,In_1541,In_2000);
nand U257 (N_257,In_2746,In_456);
or U258 (N_258,In_867,In_2169);
nand U259 (N_259,In_775,In_1629);
or U260 (N_260,In_1600,In_590);
or U261 (N_261,In_1850,In_2471);
and U262 (N_262,In_1685,In_668);
xor U263 (N_263,In_422,In_1618);
or U264 (N_264,In_1848,In_1644);
nand U265 (N_265,In_14,In_2903);
nor U266 (N_266,In_1379,In_18);
nand U267 (N_267,In_215,In_468);
nor U268 (N_268,In_1343,In_1291);
xor U269 (N_269,In_2791,In_1533);
nand U270 (N_270,In_1786,In_2250);
nand U271 (N_271,In_762,In_1005);
nor U272 (N_272,In_2675,In_2922);
nand U273 (N_273,In_597,In_1711);
and U274 (N_274,In_643,In_2309);
nand U275 (N_275,In_825,In_2847);
nor U276 (N_276,In_2943,In_2894);
and U277 (N_277,In_2820,In_2413);
or U278 (N_278,In_872,In_1649);
xnor U279 (N_279,In_2533,In_473);
nor U280 (N_280,In_2666,In_1531);
and U281 (N_281,In_338,In_2022);
or U282 (N_282,In_457,In_2080);
nand U283 (N_283,In_1706,In_90);
nor U284 (N_284,In_1322,In_1631);
nand U285 (N_285,In_1407,In_76);
xnor U286 (N_286,In_2510,In_1613);
xor U287 (N_287,In_1714,In_1478);
and U288 (N_288,In_1358,In_1236);
xor U289 (N_289,In_1597,In_784);
nor U290 (N_290,In_1248,In_1321);
and U291 (N_291,In_1293,In_176);
and U292 (N_292,In_313,In_2735);
nand U293 (N_293,In_33,In_437);
and U294 (N_294,In_1829,In_1313);
or U295 (N_295,In_1280,In_829);
nand U296 (N_296,In_1548,In_2485);
and U297 (N_297,In_2813,In_1077);
xor U298 (N_298,In_100,In_1469);
xor U299 (N_299,In_2491,In_1654);
or U300 (N_300,In_423,In_103);
xnor U301 (N_301,In_108,In_242);
and U302 (N_302,In_1169,In_2237);
nor U303 (N_303,In_2252,In_2303);
nor U304 (N_304,In_586,In_882);
or U305 (N_305,In_631,In_837);
and U306 (N_306,In_2135,In_10);
and U307 (N_307,In_1194,In_41);
or U308 (N_308,In_1205,In_2581);
nor U309 (N_309,In_1262,In_2563);
nand U310 (N_310,In_2367,In_2064);
and U311 (N_311,In_2565,In_2619);
or U312 (N_312,In_237,In_1817);
nand U313 (N_313,In_2156,In_777);
or U314 (N_314,In_2322,In_2114);
nand U315 (N_315,In_2752,In_1898);
or U316 (N_316,In_211,In_1085);
and U317 (N_317,In_2503,In_1997);
nand U318 (N_318,In_267,In_2267);
or U319 (N_319,In_2782,In_848);
and U320 (N_320,In_1121,In_635);
or U321 (N_321,In_2305,In_1592);
xor U322 (N_322,In_2155,In_61);
or U323 (N_323,In_360,In_155);
xnor U324 (N_324,In_690,In_945);
or U325 (N_325,In_340,In_78);
nand U326 (N_326,In_2817,In_212);
and U327 (N_327,In_2187,In_1749);
xnor U328 (N_328,In_529,In_1678);
or U329 (N_329,In_540,In_1364);
nand U330 (N_330,In_911,In_2404);
xnor U331 (N_331,In_2537,In_399);
and U332 (N_332,In_2781,In_2248);
nand U333 (N_333,In_1471,In_1969);
nor U334 (N_334,In_1283,In_98);
and U335 (N_335,In_2698,In_2435);
or U336 (N_336,In_1996,In_885);
nor U337 (N_337,In_2039,In_2996);
xnor U338 (N_338,In_1813,In_1572);
and U339 (N_339,In_2769,In_1724);
or U340 (N_340,In_1956,In_1411);
nand U341 (N_341,In_1584,In_1093);
or U342 (N_342,In_605,In_616);
or U343 (N_343,In_1431,In_2519);
nand U344 (N_344,In_141,In_670);
nor U345 (N_345,In_1871,In_1828);
or U346 (N_346,In_1544,In_2766);
nand U347 (N_347,In_2650,In_666);
nand U348 (N_348,In_949,In_193);
and U349 (N_349,In_2864,In_1310);
nor U350 (N_350,In_2081,In_2860);
nand U351 (N_351,In_1150,In_236);
nand U352 (N_352,In_1417,In_2925);
xor U353 (N_353,In_909,In_1641);
xnor U354 (N_354,In_1565,In_2344);
or U355 (N_355,In_145,In_2784);
and U356 (N_356,In_2195,In_950);
xor U357 (N_357,In_1404,In_311);
nand U358 (N_358,In_1445,In_2034);
or U359 (N_359,In_2430,In_1537);
and U360 (N_360,In_297,In_2734);
or U361 (N_361,In_2711,In_1664);
nand U362 (N_362,In_2256,In_1346);
and U363 (N_363,In_2015,In_1176);
and U364 (N_364,In_1022,In_2325);
and U365 (N_365,In_1378,In_57);
nor U366 (N_366,In_2440,In_744);
and U367 (N_367,In_596,In_2211);
and U368 (N_368,In_2811,In_474);
nor U369 (N_369,In_1608,In_914);
and U370 (N_370,In_2049,In_2500);
nand U371 (N_371,In_1518,In_16);
nand U372 (N_372,In_2512,In_1722);
nor U373 (N_373,In_652,In_99);
nand U374 (N_374,In_329,In_1429);
and U375 (N_375,In_2201,In_1792);
and U376 (N_376,In_968,In_1449);
xor U377 (N_377,In_2059,In_278);
or U378 (N_378,In_1199,In_936);
nand U379 (N_379,In_2247,In_2263);
and U380 (N_380,In_1259,In_520);
nand U381 (N_381,In_35,In_109);
or U382 (N_382,In_607,In_452);
xor U383 (N_383,In_1734,In_1468);
nor U384 (N_384,In_1221,In_753);
xor U385 (N_385,In_384,In_771);
xor U386 (N_386,In_1708,In_889);
nand U387 (N_387,In_582,In_143);
and U388 (N_388,In_2613,In_818);
nand U389 (N_389,In_813,In_2789);
nand U390 (N_390,In_401,In_1189);
nor U391 (N_391,In_558,In_2296);
nor U392 (N_392,In_1822,In_1556);
and U393 (N_393,In_1135,In_2980);
xnor U394 (N_394,In_893,In_2717);
xnor U395 (N_395,In_140,In_1232);
xor U396 (N_396,In_1538,In_1856);
nor U397 (N_397,In_615,In_997);
or U398 (N_398,In_1869,In_2657);
or U399 (N_399,In_731,In_2783);
nand U400 (N_400,In_1090,In_955);
xnor U401 (N_401,In_2157,In_1267);
and U402 (N_402,In_1576,In_82);
nand U403 (N_403,In_194,In_1247);
or U404 (N_404,In_1937,In_2090);
nand U405 (N_405,In_2175,In_899);
xor U406 (N_406,In_2724,In_525);
nand U407 (N_407,In_2590,In_1281);
nand U408 (N_408,In_2189,In_2913);
or U409 (N_409,In_860,In_530);
and U410 (N_410,In_345,In_2802);
xnor U411 (N_411,In_158,In_634);
nor U412 (N_412,In_2527,In_556);
xnor U413 (N_413,In_981,In_1061);
nand U414 (N_414,In_2606,In_1133);
nor U415 (N_415,In_429,In_2087);
nand U416 (N_416,In_2437,In_2536);
nor U417 (N_417,In_1767,In_1273);
nand U418 (N_418,In_1148,In_2927);
and U419 (N_419,In_2287,In_2807);
xnor U420 (N_420,In_458,In_2405);
nand U421 (N_421,In_5,In_2481);
or U422 (N_422,In_1052,In_1653);
and U423 (N_423,In_1381,In_541);
and U424 (N_424,In_1173,In_1924);
nor U425 (N_425,In_188,In_1765);
xnor U426 (N_426,In_838,In_2671);
or U427 (N_427,In_849,In_1610);
nand U428 (N_428,In_1441,In_1718);
and U429 (N_429,In_189,In_2621);
and U430 (N_430,In_1826,In_1030);
nand U431 (N_431,In_2549,In_2710);
nor U432 (N_432,In_1424,In_1071);
nand U433 (N_433,In_249,In_173);
xnor U434 (N_434,In_1884,In_1532);
nor U435 (N_435,In_593,In_2628);
or U436 (N_436,In_250,In_2244);
xnor U437 (N_437,In_673,In_561);
xnor U438 (N_438,In_30,In_253);
nand U439 (N_439,In_1974,In_1866);
nor U440 (N_440,In_2484,In_1901);
or U441 (N_441,In_789,In_1246);
or U442 (N_442,In_2477,In_2443);
nor U443 (N_443,In_2901,In_233);
or U444 (N_444,In_1980,In_773);
xor U445 (N_445,In_2829,In_1257);
nor U446 (N_446,In_1354,In_2273);
nor U447 (N_447,In_149,In_106);
and U448 (N_448,In_1099,In_1916);
nand U449 (N_449,In_43,In_2940);
or U450 (N_450,In_1195,In_2975);
nand U451 (N_451,In_461,In_2598);
and U452 (N_452,In_2561,In_2054);
xor U453 (N_453,In_2185,In_1149);
xnor U454 (N_454,In_1872,In_432);
nand U455 (N_455,In_601,In_1101);
nand U456 (N_456,In_1278,In_263);
nor U457 (N_457,In_2265,In_1066);
or U458 (N_458,In_2498,In_1372);
nand U459 (N_459,In_579,In_2455);
xnor U460 (N_460,In_1979,In_216);
and U461 (N_461,In_1923,In_2725);
xor U462 (N_462,In_245,In_490);
xnor U463 (N_463,In_1046,In_1211);
nand U464 (N_464,In_1778,In_2445);
and U465 (N_465,In_2130,In_104);
xor U466 (N_466,In_2271,In_1104);
and U467 (N_467,In_296,In_711);
or U468 (N_468,In_2274,In_2518);
and U469 (N_469,In_2346,In_1860);
nand U470 (N_470,In_991,In_308);
xnor U471 (N_471,In_466,In_450);
and U472 (N_472,In_2,In_119);
and U473 (N_473,In_2158,In_1297);
or U474 (N_474,In_1754,In_2422);
xnor U475 (N_475,In_1183,In_2624);
and U476 (N_476,In_2861,In_413);
xnor U477 (N_477,In_1016,In_1344);
nand U478 (N_478,In_214,In_1624);
nor U479 (N_479,In_2006,In_2062);
and U480 (N_480,In_2216,In_888);
xnor U481 (N_481,In_1215,In_2516);
xnor U482 (N_482,In_2029,In_180);
and U483 (N_483,In_1162,In_583);
and U484 (N_484,In_1859,In_516);
or U485 (N_485,In_2017,In_1759);
nand U486 (N_486,In_172,In_1615);
or U487 (N_487,In_241,In_1300);
xnor U488 (N_488,In_1558,In_500);
and U489 (N_489,In_992,In_1540);
or U490 (N_490,In_299,In_290);
xnor U491 (N_491,In_2693,In_273);
xor U492 (N_492,In_2394,In_333);
xor U493 (N_493,In_1527,In_1261);
xor U494 (N_494,In_138,In_1391);
xor U495 (N_495,In_2036,In_113);
xnor U496 (N_496,In_1935,In_2266);
nand U497 (N_497,In_1002,In_431);
nand U498 (N_498,In_1124,In_2068);
nor U499 (N_499,In_2839,In_1386);
xor U500 (N_500,In_854,In_2335);
xor U501 (N_501,In_1302,In_2356);
nor U502 (N_502,In_2883,In_2564);
nor U503 (N_503,In_2100,In_1142);
nor U504 (N_504,In_2629,In_874);
and U505 (N_505,In_2302,In_74);
and U506 (N_506,In_346,In_2763);
nand U507 (N_507,In_2733,In_110);
and U508 (N_508,In_1396,In_2991);
and U509 (N_509,In_1357,In_165);
nand U510 (N_510,In_1037,In_1957);
or U511 (N_511,In_1864,In_1466);
nor U512 (N_512,In_697,In_2760);
nand U513 (N_513,In_576,In_1662);
and U514 (N_514,In_2300,In_511);
or U515 (N_515,In_2482,In_841);
nand U516 (N_516,In_1713,In_2234);
xor U517 (N_517,In_300,In_1886);
xnor U518 (N_518,In_637,In_2591);
nor U519 (N_519,In_2423,In_742);
xnor U520 (N_520,In_1451,In_696);
nor U521 (N_521,In_2902,In_2595);
xor U522 (N_522,In_2132,In_475);
xor U523 (N_523,In_989,In_2292);
xor U524 (N_524,In_428,In_2726);
nor U525 (N_525,In_2562,In_1550);
nand U526 (N_526,In_1530,In_1989);
and U527 (N_527,In_1058,In_39);
nor U528 (N_528,In_36,In_2642);
nor U529 (N_529,In_691,In_780);
xor U530 (N_530,In_1185,In_1382);
xor U531 (N_531,In_2096,In_1867);
and U532 (N_532,In_940,In_674);
nor U533 (N_533,In_1805,In_2223);
xor U534 (N_534,In_1605,In_1647);
nor U535 (N_535,In_1700,In_1798);
or U536 (N_536,In_2611,In_504);
or U537 (N_537,In_1369,In_2125);
nand U538 (N_538,In_1808,In_749);
or U539 (N_539,In_56,In_751);
or U540 (N_540,In_801,In_2824);
nand U541 (N_541,In_980,In_295);
and U542 (N_542,In_1750,In_1516);
or U543 (N_543,In_1814,In_496);
nor U544 (N_544,In_978,In_2063);
or U545 (N_545,In_2804,In_1276);
xnor U546 (N_546,In_75,In_2956);
nand U547 (N_547,In_960,In_482);
nor U548 (N_548,In_1454,In_1405);
and U549 (N_549,In_1506,In_205);
nor U550 (N_550,In_2855,In_1842);
xnor U551 (N_551,In_2227,In_105);
nor U552 (N_552,In_1833,In_121);
or U553 (N_553,In_2060,In_2333);
xnor U554 (N_554,In_1214,In_1907);
and U555 (N_555,In_307,In_2768);
xnor U556 (N_556,In_1129,In_2944);
or U557 (N_557,In_1224,In_2815);
nor U558 (N_558,In_2174,In_19);
and U559 (N_559,In_664,In_351);
xnor U560 (N_560,In_1015,In_2775);
nor U561 (N_561,In_2340,In_2631);
nand U562 (N_562,In_1603,In_2896);
or U563 (N_563,In_2352,In_2955);
xnor U564 (N_564,In_276,In_2912);
or U565 (N_565,In_2947,In_2643);
nor U566 (N_566,In_692,In_2904);
or U567 (N_567,In_2424,In_1951);
xor U568 (N_568,In_549,In_2951);
and U569 (N_569,In_630,In_2744);
or U570 (N_570,In_2261,In_2061);
xor U571 (N_571,In_820,In_380);
nor U572 (N_572,In_1462,In_1643);
and U573 (N_573,In_2900,In_1153);
nand U574 (N_574,In_625,In_2052);
or U575 (N_575,In_2314,In_931);
nor U576 (N_576,In_1694,In_994);
nand U577 (N_577,In_921,In_2398);
nand U578 (N_578,In_315,In_1421);
nand U579 (N_579,In_1375,In_1594);
or U580 (N_580,In_2336,In_1853);
nand U581 (N_581,In_1265,In_2214);
xnor U582 (N_582,In_2663,In_1701);
xor U583 (N_583,In_2929,In_1847);
or U584 (N_584,In_2204,In_1336);
nor U585 (N_585,In_1758,In_832);
nand U586 (N_586,In_1819,In_1645);
xor U587 (N_587,In_1319,In_707);
or U588 (N_588,In_606,In_2910);
nor U589 (N_589,In_354,In_1230);
and U590 (N_590,In_1940,In_2550);
and U591 (N_591,In_971,In_1197);
or U592 (N_592,In_2538,In_560);
nand U593 (N_593,In_2667,In_2993);
and U594 (N_594,In_251,In_95);
xnor U595 (N_595,In_1707,In_1810);
or U596 (N_596,In_2454,In_1385);
nand U597 (N_597,In_641,In_114);
xnor U598 (N_598,In_460,In_948);
nand U599 (N_599,In_175,In_776);
nor U600 (N_600,N_462,N_225);
or U601 (N_601,In_2091,In_2673);
and U602 (N_602,In_1398,In_1717);
or U603 (N_603,In_1687,N_540);
xor U604 (N_604,In_118,In_531);
or U605 (N_605,In_2875,In_2708);
xnor U606 (N_606,In_794,N_356);
or U607 (N_607,In_2136,In_1639);
xor U608 (N_608,N_326,In_1074);
and U609 (N_609,In_1609,In_200);
or U610 (N_610,N_185,In_1515);
or U611 (N_611,N_409,N_29);
and U612 (N_612,In_592,In_2283);
xnor U613 (N_613,N_166,In_1905);
and U614 (N_614,In_2529,N_358);
nand U615 (N_615,In_609,N_299);
nand U616 (N_616,N_191,In_1851);
nand U617 (N_617,In_2131,In_1290);
or U618 (N_618,N_504,In_2021);
xor U619 (N_619,In_2878,In_2786);
xnor U620 (N_620,N_214,In_1976);
or U621 (N_621,N_440,In_1635);
or U622 (N_622,In_721,In_357);
xor U623 (N_623,In_1571,In_1286);
nand U624 (N_624,In_286,N_421);
and U625 (N_625,In_258,N_514);
nor U626 (N_626,N_67,In_2308);
nor U627 (N_627,In_1481,In_1973);
and U628 (N_628,In_1216,N_60);
and U629 (N_629,In_591,In_2198);
or U630 (N_630,N_432,In_718);
nand U631 (N_631,In_2450,N_37);
and U632 (N_632,In_2004,In_1689);
xor U633 (N_633,In_327,In_2679);
nand U634 (N_634,In_1727,In_1768);
nand U635 (N_635,In_2254,In_1092);
nand U636 (N_636,In_1388,In_2723);
and U637 (N_637,N_302,N_518);
or U638 (N_638,In_658,In_671);
nand U639 (N_639,In_1716,In_2241);
or U640 (N_640,In_2664,N_141);
or U641 (N_641,In_748,In_735);
or U642 (N_642,In_152,In_1981);
or U643 (N_643,In_986,In_96);
and U644 (N_644,In_1769,N_571);
or U645 (N_645,N_186,N_99);
nor U646 (N_646,In_1748,In_1159);
nand U647 (N_647,In_190,In_1351);
or U648 (N_648,In_1606,In_1831);
xnor U649 (N_649,In_2683,In_154);
and U650 (N_650,In_349,In_1368);
and U651 (N_651,In_2795,In_855);
or U652 (N_652,In_1491,In_693);
or U653 (N_653,N_447,In_1155);
or U654 (N_654,In_708,N_467);
xnor U655 (N_655,In_2911,N_375);
and U656 (N_656,In_1188,In_1975);
nand U657 (N_657,In_201,In_454);
nor U658 (N_658,In_1498,In_1955);
nand U659 (N_659,In_426,In_2635);
nor U660 (N_660,In_2023,In_1245);
and U661 (N_661,In_565,In_269);
and U662 (N_662,In_1465,In_1611);
or U663 (N_663,In_2686,In_1460);
and U664 (N_664,In_1289,In_1226);
nand U665 (N_665,In_1646,In_1682);
nand U666 (N_666,N_347,In_243);
nand U667 (N_667,N_493,In_259);
xnor U668 (N_668,In_695,In_1243);
and U669 (N_669,In_1470,In_1406);
nand U670 (N_670,In_689,In_92);
nor U671 (N_671,In_969,In_512);
nand U672 (N_672,In_765,N_473);
and U673 (N_673,N_310,In_1834);
or U674 (N_674,In_1880,In_2866);
nand U675 (N_675,N_59,In_1415);
or U676 (N_676,N_291,In_1580);
and U677 (N_677,In_687,N_345);
nor U678 (N_678,In_1448,In_1225);
nand U679 (N_679,In_2277,In_2088);
nand U680 (N_680,N_568,In_132);
nor U681 (N_681,In_411,In_2934);
and U682 (N_682,In_510,In_1587);
nand U683 (N_683,In_2299,In_757);
or U684 (N_684,In_619,N_135);
nand U685 (N_685,N_309,N_523);
nor U686 (N_686,N_258,In_228);
nor U687 (N_687,In_1519,In_2436);
and U688 (N_688,In_595,In_1420);
xnor U689 (N_689,In_2495,In_2094);
xnor U690 (N_690,In_1126,In_2166);
or U691 (N_691,In_186,In_2890);
or U692 (N_692,N_279,In_34);
xnor U693 (N_693,In_2547,N_174);
nor U694 (N_694,In_1968,In_277);
nand U695 (N_695,N_219,In_613);
or U696 (N_696,In_1231,In_1573);
and U697 (N_697,In_2722,In_289);
nand U698 (N_698,In_49,N_15);
nor U699 (N_699,In_2528,In_2148);
nand U700 (N_700,In_806,N_446);
and U701 (N_701,In_2147,In_367);
or U702 (N_702,N_318,N_480);
nand U703 (N_703,In_2777,In_2770);
nand U704 (N_704,In_2773,In_1501);
xnor U705 (N_705,In_1877,In_2186);
nand U706 (N_706,In_2209,N_289);
or U707 (N_707,In_1900,In_908);
and U708 (N_708,In_654,N_579);
or U709 (N_709,In_983,In_1241);
xor U710 (N_710,N_392,In_445);
xnor U711 (N_711,In_1692,N_552);
nand U712 (N_712,In_2754,In_645);
or U713 (N_713,In_2290,In_2470);
and U714 (N_714,In_1946,In_884);
or U715 (N_715,N_300,N_478);
nand U716 (N_716,In_1953,In_1025);
nor U717 (N_717,In_1123,N_50);
or U718 (N_718,In_2594,In_653);
nand U719 (N_719,In_2965,N_58);
nand U720 (N_720,In_1680,In_2736);
xor U721 (N_721,N_574,In_2293);
and U722 (N_722,In_2371,In_1392);
and U723 (N_723,In_570,In_995);
nor U724 (N_724,In_1776,In_1598);
xnor U725 (N_725,In_1876,In_2393);
xnor U726 (N_726,N_249,In_366);
or U727 (N_727,In_2677,In_1081);
xnor U728 (N_728,In_1943,N_445);
nor U729 (N_729,N_260,In_2572);
and U730 (N_730,In_382,In_1999);
xor U731 (N_731,N_100,In_1080);
and U732 (N_732,In_1453,In_527);
or U733 (N_733,In_1068,In_2876);
nand U734 (N_734,In_728,In_1342);
or U735 (N_735,N_283,N_216);
nor U736 (N_736,In_2577,In_1751);
and U737 (N_737,In_1308,In_716);
and U738 (N_738,N_114,In_2665);
nor U739 (N_739,N_17,In_2310);
nand U740 (N_740,In_1906,N_452);
and U741 (N_741,In_959,In_2390);
nor U742 (N_742,In_857,N_117);
nand U743 (N_743,In_1663,N_103);
or U744 (N_744,N_244,In_2559);
and U745 (N_745,In_1235,In_2641);
xnor U746 (N_746,In_752,In_2042);
nor U747 (N_747,In_677,N_450);
xnor U748 (N_748,In_1987,In_305);
nand U749 (N_749,In_1222,In_1233);
or U750 (N_750,In_2835,In_650);
or U751 (N_751,In_341,In_2038);
or U752 (N_752,In_875,In_1141);
nand U753 (N_753,In_1914,In_1903);
and U754 (N_754,N_276,In_2870);
nor U755 (N_755,N_598,In_393);
and U756 (N_756,In_2772,In_2217);
xnor U757 (N_757,In_28,In_2475);
nor U758 (N_758,In_2982,N_266);
nand U759 (N_759,In_1239,In_497);
nor U760 (N_760,In_350,N_465);
xnor U761 (N_761,N_351,In_1298);
nor U762 (N_762,In_1413,N_468);
and U763 (N_763,In_896,In_1986);
xor U764 (N_764,N_284,In_2240);
nand U765 (N_765,N_239,N_542);
and U766 (N_766,N_336,In_2329);
nor U767 (N_767,In_126,In_2140);
or U768 (N_768,In_594,In_2007);
xnor U769 (N_769,In_566,In_32);
nor U770 (N_770,In_2946,In_599);
nor U771 (N_771,In_1024,In_87);
xor U772 (N_772,In_573,In_2257);
xnor U773 (N_773,In_876,In_1895);
nand U774 (N_774,N_88,In_469);
or U775 (N_775,N_394,In_2532);
and U776 (N_776,N_221,In_2171);
or U777 (N_777,N_255,In_462);
nor U778 (N_778,N_362,In_649);
and U779 (N_779,In_681,N_497);
and U780 (N_780,In_1978,N_544);
nor U781 (N_781,N_6,In_961);
xor U782 (N_782,In_1630,In_2779);
or U783 (N_783,In_306,N_261);
xor U784 (N_784,In_528,In_602);
or U785 (N_785,N_23,N_589);
and U786 (N_786,In_2694,In_1652);
xnor U787 (N_787,In_3,N_229);
and U788 (N_788,In_2109,In_962);
nand U789 (N_789,In_1304,In_361);
nor U790 (N_790,In_71,N_321);
or U791 (N_791,In_2354,N_112);
nor U792 (N_792,In_1103,In_182);
or U793 (N_793,N_49,In_990);
nand U794 (N_794,In_2615,In_2347);
nor U795 (N_795,In_2610,N_479);
and U796 (N_796,In_895,In_1400);
nand U797 (N_797,In_2957,N_169);
and U798 (N_798,N_414,In_726);
and U799 (N_799,In_79,In_2522);
xnor U800 (N_800,N_106,In_836);
or U801 (N_801,In_2526,In_1365);
nor U802 (N_802,N_360,In_2620);
and U803 (N_803,N_592,N_28);
xnor U804 (N_804,In_1217,In_359);
or U805 (N_805,In_1585,In_807);
xnor U806 (N_806,In_1559,In_2320);
and U807 (N_807,In_834,In_2750);
nor U808 (N_808,In_199,In_331);
nor U809 (N_809,In_736,In_1797);
or U810 (N_810,In_2432,N_195);
nor U811 (N_811,In_791,In_1152);
nor U812 (N_812,In_839,In_2397);
xor U813 (N_813,In_68,In_1739);
xor U814 (N_814,In_2921,In_944);
nor U815 (N_815,In_433,N_512);
or U816 (N_816,N_156,N_137);
nor U817 (N_817,N_294,In_1693);
nor U818 (N_818,In_495,N_63);
xor U819 (N_819,N_588,N_193);
nor U820 (N_820,In_2962,In_1456);
or U821 (N_821,N_538,N_123);
nand U822 (N_822,In_2476,In_812);
or U823 (N_823,In_639,In_2952);
nand U824 (N_824,In_2588,In_2141);
nor U825 (N_825,N_401,In_2504);
or U826 (N_826,In_373,In_2407);
and U827 (N_827,In_2701,In_1097);
nand U828 (N_828,In_2074,In_1318);
and U829 (N_829,In_642,In_2517);
nor U830 (N_830,In_488,In_2989);
and U831 (N_831,In_803,In_657);
nand U832 (N_832,N_399,In_1809);
and U833 (N_833,In_1240,In_25);
nand U834 (N_834,N_331,In_332);
or U835 (N_835,In_227,In_2759);
nor U836 (N_836,In_1766,In_344);
and U837 (N_837,N_332,In_1069);
xor U838 (N_838,N_378,In_1252);
xnor U839 (N_839,N_209,In_2753);
nand U840 (N_840,In_723,In_843);
and U841 (N_841,In_2755,In_2757);
xor U842 (N_842,In_1134,In_2580);
xor U843 (N_843,N_242,In_2078);
xor U844 (N_844,In_1892,In_1089);
and U845 (N_845,N_419,In_1160);
xnor U846 (N_846,In_2780,N_161);
nand U847 (N_847,In_1434,In_1861);
nand U848 (N_848,In_1335,In_1251);
and U849 (N_849,In_2218,N_7);
xor U850 (N_850,In_247,N_246);
nand U851 (N_851,N_305,In_1993);
nand U852 (N_852,In_2035,In_1132);
or U853 (N_853,N_408,In_1118);
nor U854 (N_854,In_2161,In_2315);
xnor U855 (N_855,In_2655,In_2359);
and U856 (N_856,In_2151,In_2869);
and U857 (N_857,In_1009,In_1930);
nand U858 (N_858,In_1475,In_178);
xor U859 (N_859,In_255,In_1535);
or U860 (N_860,In_996,In_1208);
nand U861 (N_861,N_207,In_453);
and U862 (N_862,In_374,N_140);
and U863 (N_863,In_97,In_756);
xnor U864 (N_864,In_147,In_60);
xnor U865 (N_865,N_434,In_694);
xnor U866 (N_866,In_638,In_1752);
nand U867 (N_867,In_1287,In_321);
xor U868 (N_868,In_1274,N_522);
nor U869 (N_869,In_1477,In_1116);
nand U870 (N_870,N_488,N_439);
nand U871 (N_871,In_790,In_878);
or U872 (N_872,In_1047,N_175);
nor U873 (N_873,In_2380,N_482);
nand U874 (N_874,In_1349,In_2964);
and U875 (N_875,In_786,In_1883);
and U876 (N_876,In_88,In_1686);
nor U877 (N_877,In_2630,N_367);
nor U878 (N_878,N_510,In_1285);
and U879 (N_879,In_2840,In_120);
and U880 (N_880,N_240,In_2122);
xor U881 (N_881,In_481,In_91);
and U882 (N_882,In_1484,N_529);
and U883 (N_883,In_2738,In_1393);
nor U884 (N_884,N_91,In_782);
and U885 (N_885,In_965,N_316);
nand U886 (N_886,In_747,In_136);
and U887 (N_887,N_170,In_163);
nor U888 (N_888,In_2492,In_1824);
nand U889 (N_889,In_1316,In_2525);
xnor U890 (N_890,In_2556,In_2995);
or U891 (N_891,N_183,In_1204);
xor U892 (N_892,In_1827,N_199);
nor U893 (N_893,N_1,In_1043);
or U894 (N_894,In_1888,In_720);
or U895 (N_895,In_1589,In_368);
nand U896 (N_896,In_1332,In_2378);
nand U897 (N_897,In_2906,N_320);
xor U898 (N_898,In_847,In_1539);
nor U899 (N_899,In_1095,N_491);
xnor U900 (N_900,In_442,In_679);
xor U901 (N_901,In_392,In_1377);
or U902 (N_902,In_870,In_2075);
xnor U903 (N_903,In_282,N_585);
nor U904 (N_904,In_202,In_489);
and U905 (N_905,In_1912,In_291);
nor U906 (N_906,In_1709,In_254);
and U907 (N_907,In_1617,In_554);
nor U908 (N_908,N_420,In_1311);
nand U909 (N_909,N_162,N_530);
and U910 (N_910,In_2116,In_2111);
or U911 (N_911,N_304,In_1837);
nand U912 (N_912,In_2165,In_1250);
and U913 (N_913,N_541,In_1705);
or U914 (N_914,N_322,In_1938);
xor U915 (N_915,In_1370,In_957);
or U916 (N_916,N_572,In_2690);
and U917 (N_917,In_2700,In_2249);
nor U918 (N_918,N_487,In_588);
and U919 (N_919,In_1219,In_1690);
or U920 (N_920,N_11,In_1928);
nand U921 (N_921,N_34,In_1008);
or U922 (N_922,N_550,In_1435);
and U923 (N_923,In_1192,N_431);
and U924 (N_924,In_900,N_442);
nand U925 (N_925,In_1062,N_250);
or U926 (N_926,In_746,In_2987);
and U927 (N_927,N_398,In_942);
and U928 (N_928,In_901,In_521);
xor U929 (N_929,In_1356,N_208);
or U930 (N_930,N_329,In_1184);
or U931 (N_931,In_2523,In_2748);
or U932 (N_932,In_563,N_231);
or U933 (N_933,N_376,In_903);
or U934 (N_934,In_471,In_2727);
or U935 (N_935,In_2105,N_9);
or U936 (N_936,In_135,In_2567);
nor U937 (N_937,In_146,In_1929);
nand U938 (N_938,In_265,In_2682);
and U939 (N_939,In_304,In_1726);
and U940 (N_940,In_1163,In_823);
xor U941 (N_941,In_2396,In_2282);
and U942 (N_942,In_2573,N_558);
and U943 (N_943,In_2262,In_2602);
or U944 (N_944,In_701,In_1638);
or U945 (N_945,In_956,N_325);
and U946 (N_946,N_72,In_2050);
nand U947 (N_947,In_209,In_2494);
nand U948 (N_948,N_13,In_2478);
nand U949 (N_949,In_1720,N_554);
and U950 (N_950,In_2134,N_74);
or U951 (N_951,In_2497,In_1526);
and U952 (N_952,In_2364,In_1425);
and U953 (N_953,In_1688,N_136);
xnor U954 (N_954,In_1177,N_150);
nand U955 (N_955,N_527,In_2851);
and U956 (N_956,In_2632,N_27);
nor U957 (N_957,In_2524,In_1110);
nand U958 (N_958,N_350,In_2740);
and U959 (N_959,In_730,In_898);
xnor U960 (N_960,In_678,In_1673);
and U961 (N_961,N_308,In_208);
xor U962 (N_962,In_2076,In_246);
xor U963 (N_963,In_1033,N_181);
or U964 (N_964,In_2521,In_2806);
nor U965 (N_965,In_1070,N_111);
nand U966 (N_966,In_830,In_1187);
xnor U967 (N_967,In_1894,In_150);
and U968 (N_968,In_564,In_2627);
xnor U969 (N_969,In_2858,N_515);
or U970 (N_970,N_425,In_2213);
xor U971 (N_971,N_341,In_347);
nand U972 (N_972,N_430,In_2831);
xnor U973 (N_973,In_2056,N_256);
and U974 (N_974,In_932,N_126);
xnor U975 (N_975,In_439,In_153);
or U976 (N_976,In_1329,In_2541);
or U977 (N_977,In_1306,N_203);
or U978 (N_978,In_925,N_593);
and U979 (N_979,In_1256,N_366);
and U980 (N_980,In_378,In_1931);
nand U981 (N_981,In_2409,In_1309);
or U982 (N_982,In_622,In_542);
or U983 (N_983,In_2923,In_268);
or U984 (N_984,In_2343,In_2421);
and U985 (N_985,In_1614,N_215);
nand U986 (N_986,N_365,In_571);
or U987 (N_987,In_524,N_570);
xnor U988 (N_988,In_2238,N_381);
nand U989 (N_989,In_11,In_1249);
nor U990 (N_990,In_2704,In_562);
nand U991 (N_991,N_86,In_505);
nor U992 (N_992,In_1911,In_2891);
xor U993 (N_993,In_42,In_868);
and U994 (N_994,N_265,In_2070);
nand U995 (N_995,In_2353,In_418);
xnor U996 (N_996,In_1206,In_1744);
or U997 (N_997,In_1190,In_2092);
xor U998 (N_998,N_105,N_164);
nor U999 (N_999,N_139,N_131);
nor U1000 (N_1000,In_1426,In_1333);
nand U1001 (N_1001,N_182,In_491);
nand U1002 (N_1002,N_210,N_357);
nor U1003 (N_1003,N_146,In_21);
nand U1004 (N_1004,In_745,N_511);
nor U1005 (N_1005,In_1553,N_582);
nor U1006 (N_1006,In_846,In_2451);
nand U1007 (N_1007,In_845,In_2258);
xor U1008 (N_1008,In_2408,In_355);
nor U1009 (N_1009,N_92,N_149);
and U1010 (N_1010,N_363,In_667);
nand U1011 (N_1011,In_2596,N_84);
or U1012 (N_1012,In_2019,In_1001);
nand U1013 (N_1013,In_1418,In_517);
xor U1014 (N_1014,In_2530,N_565);
and U1015 (N_1015,In_939,N_24);
xnor U1016 (N_1016,In_226,N_494);
nand U1017 (N_1017,In_181,In_2245);
nor U1018 (N_1018,N_212,In_2716);
or U1019 (N_1019,In_2483,In_1180);
and U1020 (N_1020,In_2488,N_346);
or U1021 (N_1021,In_409,In_2442);
nand U1022 (N_1022,In_2003,N_449);
and U1023 (N_1023,N_546,N_42);
nor U1024 (N_1024,N_18,N_192);
nor U1025 (N_1025,In_656,In_1885);
or U1026 (N_1026,In_1480,N_505);
or U1027 (N_1027,In_1412,In_1282);
xnor U1028 (N_1028,In_2386,N_133);
nand U1029 (N_1029,In_1175,In_438);
nor U1030 (N_1030,In_1972,N_556);
nor U1031 (N_1031,In_1264,In_2950);
or U1032 (N_1032,In_1691,N_448);
nor U1033 (N_1033,N_57,N_5);
and U1034 (N_1034,N_453,In_1966);
xnor U1035 (N_1035,In_2713,N_576);
or U1036 (N_1036,In_1737,In_2224);
and U1037 (N_1037,In_2604,N_40);
or U1038 (N_1038,In_2318,In_750);
and U1039 (N_1039,In_480,In_1422);
nor U1040 (N_1040,N_503,In_1119);
nand U1041 (N_1041,In_1581,In_499);
and U1042 (N_1042,In_2592,In_2025);
nand U1043 (N_1043,In_1041,In_699);
nor U1044 (N_1044,In_2785,In_1619);
and U1045 (N_1045,N_415,N_190);
nand U1046 (N_1046,In_238,N_83);
and U1047 (N_1047,N_38,N_508);
and U1048 (N_1048,In_400,In_58);
and U1049 (N_1049,N_454,In_2805);
xor U1050 (N_1050,In_1604,N_76);
or U1051 (N_1051,In_506,In_2401);
nand U1052 (N_1052,In_644,In_715);
xor U1053 (N_1053,In_817,In_1347);
or U1054 (N_1054,In_1889,N_477);
xor U1055 (N_1055,In_2008,In_1272);
or U1056 (N_1056,In_2905,In_1182);
nor U1057 (N_1057,In_412,N_176);
nand U1058 (N_1058,In_2933,In_2331);
nand U1059 (N_1059,In_684,N_87);
nand U1060 (N_1060,In_2284,In_2578);
nor U1061 (N_1061,N_533,N_80);
nand U1062 (N_1062,In_2419,In_2194);
or U1063 (N_1063,In_632,In_1007);
and U1064 (N_1064,In_1127,In_938);
nand U1065 (N_1065,In_1436,In_1642);
nand U1066 (N_1066,In_2908,N_569);
xor U1067 (N_1067,In_2669,In_1495);
nor U1068 (N_1068,In_2856,In_2264);
or U1069 (N_1069,In_1747,In_1147);
nand U1070 (N_1070,N_56,In_1050);
xnor U1071 (N_1071,In_2464,In_1279);
nor U1072 (N_1072,In_198,In_2544);
and U1073 (N_1073,In_1944,In_2120);
and U1074 (N_1074,In_907,N_402);
xnor U1075 (N_1075,In_1954,In_459);
xnor U1076 (N_1076,In_2219,In_2207);
nand U1077 (N_1077,In_365,In_617);
nand U1078 (N_1078,In_1299,N_8);
xor U1079 (N_1079,N_553,N_561);
nor U1080 (N_1080,In_2834,In_1657);
and U1081 (N_1081,In_2083,In_1253);
or U1082 (N_1082,N_252,In_1186);
and U1083 (N_1083,In_2814,In_2954);
or U1084 (N_1084,In_2055,In_805);
and U1085 (N_1085,In_1616,In_1839);
nor U1086 (N_1086,In_38,N_78);
and U1087 (N_1087,In_116,In_1622);
nor U1088 (N_1088,In_1579,In_1570);
and U1089 (N_1089,In_2981,N_145);
and U1090 (N_1090,In_2797,In_1228);
nor U1091 (N_1091,In_375,In_2279);
and U1092 (N_1092,N_53,In_2208);
or U1093 (N_1093,In_1811,In_1040);
or U1094 (N_1094,In_2968,In_64);
xor U1095 (N_1095,N_22,In_1427);
nand U1096 (N_1096,In_1444,In_1488);
nor U1097 (N_1097,In_424,In_792);
and U1098 (N_1098,In_2542,In_1777);
or U1099 (N_1099,N_204,In_1168);
or U1100 (N_1100,In_2472,In_218);
and U1101 (N_1101,In_2456,N_211);
xor U1102 (N_1102,In_1755,N_97);
nor U1103 (N_1103,N_459,In_669);
and U1104 (N_1104,In_1583,N_275);
nor U1105 (N_1105,In_840,In_1361);
and U1106 (N_1106,In_2960,In_1334);
xnor U1107 (N_1107,In_2833,In_1210);
nand U1108 (N_1108,In_2970,In_2732);
and U1109 (N_1109,In_2886,In_2018);
or U1110 (N_1110,In_1083,In_1710);
nand U1111 (N_1111,In_951,In_53);
or U1112 (N_1112,In_1908,In_443);
xor U1113 (N_1113,N_10,In_207);
nand U1114 (N_1114,In_2360,In_2656);
or U1115 (N_1115,In_2434,In_1882);
nand U1116 (N_1116,In_1626,In_133);
nand U1117 (N_1117,N_509,In_2077);
nand U1118 (N_1118,N_567,In_1841);
xnor U1119 (N_1119,N_313,In_1403);
and U1120 (N_1120,N_257,In_1790);
nor U1121 (N_1121,In_2009,In_1458);
nand U1122 (N_1122,In_754,In_2551);
nor U1123 (N_1123,N_247,N_79);
nand U1124 (N_1124,In_1670,In_430);
nor U1125 (N_1125,In_2505,In_1317);
xor U1126 (N_1126,N_501,In_2979);
nand U1127 (N_1127,In_2699,In_1512);
nand U1128 (N_1128,In_2406,In_2543);
or U1129 (N_1129,In_1476,In_2363);
nand U1130 (N_1130,In_2739,In_156);
and U1131 (N_1131,N_353,In_389);
nor U1132 (N_1132,In_1965,In_1191);
xor U1133 (N_1133,In_1596,In_1363);
nand U1134 (N_1134,In_1896,In_768);
and U1135 (N_1135,In_2681,In_1003);
nor U1136 (N_1136,In_2941,N_423);
xor U1137 (N_1137,N_335,N_274);
nor U1138 (N_1138,In_326,In_470);
xnor U1139 (N_1139,In_2143,In_2345);
and U1140 (N_1140,In_294,In_1117);
nand U1141 (N_1141,In_815,In_2458);
and U1142 (N_1142,N_397,In_993);
and U1143 (N_1143,In_1213,In_1428);
or U1144 (N_1144,In_1315,In_441);
nor U1145 (N_1145,In_1760,N_148);
nor U1146 (N_1146,In_922,N_104);
and U1147 (N_1147,N_463,In_2885);
nor U1148 (N_1148,In_2202,In_2040);
or U1149 (N_1149,In_772,N_259);
nand U1150 (N_1150,N_52,In_2871);
xor U1151 (N_1151,In_1507,In_808);
xnor U1152 (N_1152,In_2103,In_2355);
and U1153 (N_1153,In_2298,In_532);
xor U1154 (N_1154,In_798,In_2280);
nor U1155 (N_1155,N_557,In_1395);
nor U1156 (N_1156,In_717,In_314);
or U1157 (N_1157,N_230,In_1138);
and U1158 (N_1158,In_2994,N_142);
and U1159 (N_1159,In_2110,In_2888);
and U1160 (N_1160,In_281,N_471);
or U1161 (N_1161,In_2644,In_196);
and U1162 (N_1162,In_1012,N_129);
nor U1163 (N_1163,In_866,In_1271);
and U1164 (N_1164,In_2073,In_2737);
and U1165 (N_1165,In_2501,In_1505);
and U1166 (N_1166,In_2179,In_1875);
or U1167 (N_1167,In_2410,N_577);
or U1168 (N_1168,N_206,In_1520);
and U1169 (N_1169,In_427,In_1939);
and U1170 (N_1170,In_2822,In_2586);
nand U1171 (N_1171,N_132,In_1397);
xor U1172 (N_1172,In_627,In_1612);
nand U1173 (N_1173,In_761,In_2351);
xnor U1174 (N_1174,N_348,In_472);
xnor U1175 (N_1175,In_323,N_62);
nand U1176 (N_1176,N_272,In_600);
nand U1177 (N_1177,N_122,In_127);
xnor U1178 (N_1178,N_46,In_2044);
and U1179 (N_1179,In_719,In_1607);
and U1180 (N_1180,In_2816,In_1255);
xnor U1181 (N_1181,In_2460,In_1450);
and U1182 (N_1182,In_982,N_98);
xor U1183 (N_1183,In_1582,In_1665);
or U1184 (N_1184,In_1919,N_171);
or U1185 (N_1185,N_121,N_295);
and U1186 (N_1186,In_2603,N_134);
or U1187 (N_1187,N_19,In_1593);
or U1188 (N_1188,In_660,In_2634);
and U1189 (N_1189,In_680,N_47);
or U1190 (N_1190,In_1816,N_466);
nand U1191 (N_1191,In_2098,N_301);
or U1192 (N_1192,N_520,In_1857);
nor U1193 (N_1193,In_1863,In_1844);
or U1194 (N_1194,In_1868,In_963);
and U1195 (N_1195,In_1374,In_2268);
xnor U1196 (N_1196,In_604,In_2377);
xor U1197 (N_1197,In_2790,In_2399);
nand U1198 (N_1198,N_373,In_550);
xor U1199 (N_1199,In_2324,N_165);
xnor U1200 (N_1200,In_139,N_1028);
nand U1201 (N_1201,In_2633,N_918);
or U1202 (N_1202,N_688,In_734);
and U1203 (N_1203,N_1011,In_1307);
or U1204 (N_1204,N_981,In_1399);
and U1205 (N_1205,In_2144,In_274);
xor U1206 (N_1206,In_1268,N_1155);
nand U1207 (N_1207,In_1575,N_813);
and U1208 (N_1208,In_729,N_167);
xor U1209 (N_1209,N_220,In_1640);
nor U1210 (N_1210,N_948,N_1044);
xor U1211 (N_1211,In_2808,In_330);
xor U1212 (N_1212,N_922,In_1983);
nand U1213 (N_1213,In_467,N_1164);
nor U1214 (N_1214,N_444,In_1467);
or U1215 (N_1215,N_707,N_929);
nand U1216 (N_1216,N_282,N_1085);
and U1217 (N_1217,In_2294,N_108);
nand U1218 (N_1218,N_704,N_804);
and U1219 (N_1219,N_622,N_1032);
and U1220 (N_1220,N_1098,In_2439);
xor U1221 (N_1221,In_455,In_1511);
nor U1222 (N_1222,In_2625,In_2099);
nand U1223 (N_1223,In_2128,N_143);
xnor U1224 (N_1224,In_342,N_14);
or U1225 (N_1225,N_226,In_1783);
and U1226 (N_1226,N_405,In_1292);
and U1227 (N_1227,In_72,In_2349);
and U1228 (N_1228,In_581,In_1345);
nor U1229 (N_1229,In_2452,In_2168);
and U1230 (N_1230,In_557,In_1202);
or U1231 (N_1231,N_768,In_2917);
and U1232 (N_1232,N_406,In_1075);
and U1233 (N_1233,In_86,In_943);
xnor U1234 (N_1234,In_1201,N_389);
and U1235 (N_1235,N_93,In_2479);
and U1236 (N_1236,N_273,In_2794);
or U1237 (N_1237,N_645,N_413);
and U1238 (N_1238,In_1793,In_1513);
nand U1239 (N_1239,In_234,In_2945);
nand U1240 (N_1240,N_548,In_1029);
nor U1241 (N_1241,N_90,N_783);
and U1242 (N_1242,N_535,In_385);
xor U1243 (N_1243,In_2712,N_500);
xnor U1244 (N_1244,N_233,In_1697);
and U1245 (N_1245,N_407,N_532);
xnor U1246 (N_1246,In_2932,N_642);
xor U1247 (N_1247,In_417,N_158);
nor U1248 (N_1248,In_910,N_709);
and U1249 (N_1249,N_950,In_2251);
nand U1250 (N_1250,N_70,N_963);
nand U1251 (N_1251,In_2692,N_575);
or U1252 (N_1252,N_655,In_1223);
nor U1253 (N_1253,N_372,In_2069);
nor U1254 (N_1254,In_1220,In_1698);
nand U1255 (N_1255,In_1742,In_929);
and U1256 (N_1256,In_821,N_1009);
nand U1257 (N_1257,N_1181,N_436);
xor U1258 (N_1258,N_179,In_1636);
xnor U1259 (N_1259,In_1920,In_2706);
nand U1260 (N_1260,N_155,N_780);
or U1261 (N_1261,In_1849,In_1918);
and U1262 (N_1262,N_827,In_2874);
nand U1263 (N_1263,In_1881,N_374);
nand U1264 (N_1264,N_172,N_683);
and U1265 (N_1265,N_382,N_955);
nor U1266 (N_1266,In_2400,In_2027);
and U1267 (N_1267,In_1674,In_1528);
and U1268 (N_1268,N_96,In_1941);
xor U1269 (N_1269,N_587,In_2231);
nor U1270 (N_1270,In_2918,In_2093);
xor U1271 (N_1271,In_610,In_2771);
nor U1272 (N_1272,In_1079,In_1461);
or U1273 (N_1273,N_352,N_153);
xnor U1274 (N_1274,In_2654,N_513);
or U1275 (N_1275,In_2652,In_2260);
nand U1276 (N_1276,In_1637,In_1926);
and U1277 (N_1277,In_1366,N_604);
or U1278 (N_1278,N_649,N_618);
or U1279 (N_1279,N_605,N_782);
nand U1280 (N_1280,In_2253,N_787);
and U1281 (N_1281,In_2127,In_1510);
and U1282 (N_1282,In_603,In_755);
nor U1283 (N_1283,N_441,N_237);
and U1284 (N_1284,In_1627,N_77);
and U1285 (N_1285,In_779,N_403);
nor U1286 (N_1286,In_1745,In_844);
xor U1287 (N_1287,N_410,N_370);
and U1288 (N_1288,In_129,N_241);
or U1289 (N_1289,N_1193,In_814);
nand U1290 (N_1290,In_802,N_770);
and U1291 (N_1291,N_951,N_1185);
nand U1292 (N_1292,N_102,N_721);
and U1293 (N_1293,In_2465,In_672);
nor U1294 (N_1294,N_68,N_699);
nand U1295 (N_1295,In_2558,In_923);
or U1296 (N_1296,In_434,N_615);
and U1297 (N_1297,In_2415,N_1040);
and U1298 (N_1298,In_2365,In_544);
xor U1299 (N_1299,In_2321,N_1022);
nor U1300 (N_1300,N_1114,N_606);
or U1301 (N_1301,In_2877,In_2466);
nor U1302 (N_1302,N_866,N_778);
or U1303 (N_1303,N_160,In_63);
and U1304 (N_1304,In_1874,N_472);
or U1305 (N_1305,In_134,In_640);
and U1306 (N_1306,N_952,N_910);
nand U1307 (N_1307,In_1082,In_2684);
and U1308 (N_1308,N_1119,N_818);
nor U1309 (N_1309,N_641,N_1147);
or U1310 (N_1310,In_2583,N_1162);
nand U1311 (N_1311,N_1152,In_2286);
nand U1312 (N_1312,N_1101,In_2741);
and U1313 (N_1313,In_1902,N_854);
and U1314 (N_1314,In_1932,N_573);
nor U1315 (N_1315,N_700,N_427);
nor U1316 (N_1316,In_2046,In_2674);
and U1317 (N_1317,In_2843,In_1500);
nand U1318 (N_1318,In_1936,In_2545);
and U1319 (N_1319,In_2487,N_380);
xor U1320 (N_1320,In_1339,In_2718);
and U1321 (N_1321,In_1146,In_271);
nor U1322 (N_1322,In_2453,N_187);
xnor U1323 (N_1323,In_535,N_461);
or U1324 (N_1324,N_940,In_213);
xnor U1325 (N_1325,In_2977,N_130);
or U1326 (N_1326,In_2473,In_919);
or U1327 (N_1327,In_2084,N_458);
nand U1328 (N_1328,N_173,N_839);
nor U1329 (N_1329,N_32,N_586);
and U1330 (N_1330,N_760,N_860);
xor U1331 (N_1331,N_1041,N_695);
and U1332 (N_1332,In_17,N_735);
xor U1333 (N_1333,In_800,N_119);
nor U1334 (N_1334,N_673,In_1301);
nor U1335 (N_1335,In_1787,N_819);
or U1336 (N_1336,N_429,N_863);
nor U1337 (N_1337,In_733,N_1123);
xor U1338 (N_1338,In_1137,In_703);
xnor U1339 (N_1339,N_1150,N_844);
or U1340 (N_1340,In_2337,N_644);
xnor U1341 (N_1341,In_1566,N_824);
xor U1342 (N_1342,In_2461,N_621);
xor U1343 (N_1343,In_398,In_2570);
xor U1344 (N_1344,N_722,In_1337);
nor U1345 (N_1345,In_435,N_665);
nor U1346 (N_1346,In_1096,In_1574);
and U1347 (N_1347,N_1087,N_1109);
xor U1348 (N_1348,N_761,In_1961);
xor U1349 (N_1349,In_2715,In_547);
xnor U1350 (N_1350,In_2552,N_781);
or U1351 (N_1351,In_376,N_120);
nand U1352 (N_1352,In_738,In_2449);
nor U1353 (N_1353,In_833,In_66);
nand U1354 (N_1354,N_899,In_1367);
and U1355 (N_1355,In_2301,N_754);
xor U1356 (N_1356,In_1732,In_2948);
xor U1357 (N_1357,N_1143,N_893);
or U1358 (N_1358,In_665,In_2566);
nand U1359 (N_1359,In_59,In_987);
xnor U1360 (N_1360,In_1479,N_698);
or U1361 (N_1361,In_984,In_1013);
xnor U1362 (N_1362,N_163,N_739);
nand U1363 (N_1363,In_1985,In_2182);
or U1364 (N_1364,N_664,In_1971);
and U1365 (N_1365,N_883,N_609);
nor U1366 (N_1366,In_1323,N_1179);
and U1367 (N_1367,N_107,In_1474);
nor U1368 (N_1368,In_2328,In_2362);
and U1369 (N_1369,In_2639,N_1012);
and U1370 (N_1370,In_167,N_1083);
and U1371 (N_1371,N_1003,In_663);
nand U1372 (N_1372,In_2259,N_438);
xor U1373 (N_1373,N_73,N_271);
nor U1374 (N_1374,In_2534,In_309);
or U1375 (N_1375,N_634,N_369);
xor U1376 (N_1376,N_1045,N_563);
nor U1377 (N_1377,In_6,In_1517);
or U1378 (N_1378,In_2688,N_349);
xor U1379 (N_1379,N_985,N_915);
and U1380 (N_1380,N_898,N_1039);
and U1381 (N_1381,N_1105,N_814);
nor U1382 (N_1382,N_109,N_647);
nor U1383 (N_1383,N_980,N_894);
xor U1384 (N_1384,N_178,In_781);
and U1385 (N_1385,N_651,In_2930);
xor U1386 (N_1386,N_595,In_686);
xnor U1387 (N_1387,N_753,N_687);
xor U1388 (N_1388,In_2108,In_225);
nand U1389 (N_1389,In_4,N_603);
or U1390 (N_1390,In_1157,In_23);
nand U1391 (N_1391,In_235,In_1825);
nor U1392 (N_1392,N_612,N_879);
xnor U1393 (N_1393,N_492,N_895);
and U1394 (N_1394,N_507,N_344);
xnor U1395 (N_1395,In_2520,In_2862);
and U1396 (N_1396,N_312,In_1242);
and U1397 (N_1397,N_905,In_386);
or U1398 (N_1398,N_101,In_1004);
nor U1399 (N_1399,N_868,N_1173);
nor U1400 (N_1400,In_2348,N_974);
or U1401 (N_1401,N_433,N_154);
nor U1402 (N_1402,In_1109,N_1030);
nor U1403 (N_1403,In_2496,In_1704);
nand U1404 (N_1404,In_1106,In_2661);
nor U1405 (N_1405,In_879,In_1);
nand U1406 (N_1406,In_975,In_2809);
xor U1407 (N_1407,N_417,In_2756);
xor U1408 (N_1408,N_932,N_1153);
xnor U1409 (N_1409,In_2938,In_2827);
nand U1410 (N_1410,N_831,N_661);
xor U1411 (N_1411,N_267,N_911);
nand U1412 (N_1412,N_1191,In_1730);
nor U1413 (N_1413,N_384,In_244);
and U1414 (N_1414,N_1099,N_285);
xor U1415 (N_1415,In_897,N_800);
or U1416 (N_1416,In_2285,N_243);
or U1417 (N_1417,In_1355,In_1904);
or U1418 (N_1418,In_2001,N_115);
nor U1419 (N_1419,N_338,In_1899);
nand U1420 (N_1420,In_1599,N_490);
nand U1421 (N_1421,N_1175,In_1108);
and U1422 (N_1422,N_941,In_1091);
nand U1423 (N_1423,N_715,In_2220);
xnor U1424 (N_1424,In_2188,In_1659);
xor U1425 (N_1425,In_1353,N_817);
or U1426 (N_1426,In_1591,In_1087);
and U1427 (N_1427,In_339,N_21);
and U1428 (N_1428,N_845,In_501);
nor U1429 (N_1429,In_2787,In_852);
and U1430 (N_1430,N_847,N_639);
xnor U1431 (N_1431,N_931,N_1159);
nor U1432 (N_1432,N_815,In_2731);
or U1433 (N_1433,In_727,In_2893);
nor U1434 (N_1434,In_264,In_850);
or U1435 (N_1435,N_978,N_1142);
nand U1436 (N_1436,In_1122,In_2617);
and U1437 (N_1437,N_772,In_2721);
xor U1438 (N_1438,In_1578,N_1066);
and U1439 (N_1439,N_531,In_2730);
and U1440 (N_1440,N_599,In_2728);
or U1441 (N_1441,N_578,In_1913);
xor U1442 (N_1442,N_1124,In_1076);
nand U1443 (N_1443,In_1774,In_2048);
xor U1444 (N_1444,N_1184,N_51);
nand U1445 (N_1445,N_1075,In_1051);
and U1446 (N_1446,N_303,N_924);
and U1447 (N_1447,In_316,N_218);
xor U1448 (N_1448,In_1128,N_1062);
nor U1449 (N_1449,In_387,N_733);
and U1450 (N_1450,In_1229,N_94);
xnor U1451 (N_1451,N_808,N_1002);
and U1452 (N_1452,N_1174,N_1170);
xor U1453 (N_1453,N_1048,In_1237);
nand U1454 (N_1454,In_1408,In_1756);
and U1455 (N_1455,In_2798,N_470);
xor U1456 (N_1456,N_842,In_1651);
xor U1457 (N_1457,In_880,In_320);
xor U1458 (N_1458,N_1177,In_1166);
and U1459 (N_1459,N_961,In_683);
nand U1460 (N_1460,In_124,N_943);
nand U1461 (N_1461,N_502,N_1140);
or U1462 (N_1462,N_1086,N_516);
nor U1463 (N_1463,N_855,N_549);
xor U1464 (N_1464,N_1063,In_2382);
and U1465 (N_1465,N_993,N_456);
and U1466 (N_1466,N_878,In_1494);
nand U1467 (N_1467,In_1870,In_724);
or U1468 (N_1468,In_1209,N_597);
and U1469 (N_1469,In_128,In_1414);
nand U1470 (N_1470,In_2341,N_517);
nor U1471 (N_1471,N_526,In_2879);
xor U1472 (N_1472,N_871,In_1049);
and U1473 (N_1473,N_773,In_2067);
nand U1474 (N_1474,N_986,N_816);
nand U1475 (N_1475,In_826,N_891);
or U1476 (N_1476,In_1569,In_770);
xnor U1477 (N_1477,N_151,In_851);
nand U1478 (N_1478,N_262,In_1735);
and U1479 (N_1479,In_1958,N_583);
and U1480 (N_1480,N_693,N_913);
and U1481 (N_1481,N_742,In_343);
and U1482 (N_1482,N_789,N_147);
and U1483 (N_1483,In_1588,N_152);
and U1484 (N_1484,In_1277,In_2374);
or U1485 (N_1485,In_2651,In_174);
nand U1486 (N_1486,In_2031,N_1010);
nand U1487 (N_1487,N_264,N_676);
xor U1488 (N_1488,In_2892,In_2509);
nand U1489 (N_1489,N_1115,N_876);
nor U1490 (N_1490,N_315,N_95);
and U1491 (N_1491,In_2825,In_421);
or U1492 (N_1492,In_26,In_288);
nor U1493 (N_1493,N_619,In_31);
xor U1494 (N_1494,In_612,In_1027);
nand U1495 (N_1495,N_1067,N_719);
and U1496 (N_1496,N_959,N_1089);
xnor U1497 (N_1497,In_904,In_1327);
nor U1498 (N_1498,N_853,In_1590);
nand U1499 (N_1499,N_1138,In_1234);
nor U1500 (N_1500,N_904,In_513);
nor U1501 (N_1501,N_180,In_618);
or U1502 (N_1502,In_1699,In_1781);
and U1503 (N_1503,In_1950,In_1086);
nor U1504 (N_1504,N_364,N_1065);
nand U1505 (N_1505,In_810,N_213);
or U1506 (N_1506,In_2139,In_1125);
or U1507 (N_1507,N_600,N_685);
or U1508 (N_1508,In_1060,N_1007);
nand U1509 (N_1509,In_1164,N_886);
nor U1510 (N_1510,In_160,N_238);
and U1511 (N_1511,N_1107,N_455);
xnor U1512 (N_1512,N_631,In_2799);
or U1513 (N_1513,In_623,N_691);
nand U1514 (N_1514,N_1047,In_2571);
nand U1515 (N_1515,N_638,N_16);
xor U1516 (N_1516,In_2852,N_791);
nand U1517 (N_1517,In_795,N_616);
nor U1518 (N_1518,In_478,In_928);
xor U1519 (N_1519,In_514,In_1934);
nor U1520 (N_1520,N_124,In_740);
nor U1521 (N_1521,In_1555,N_607);
nor U1522 (N_1522,In_2593,N_416);
nand U1523 (N_1523,In_1490,N_714);
and U1524 (N_1524,N_437,In_1338);
nor U1525 (N_1525,N_835,In_2416);
and U1526 (N_1526,In_759,In_334);
and U1527 (N_1527,N_795,In_2697);
or U1528 (N_1528,N_900,N_1144);
nor U1529 (N_1529,N_390,In_130);
nand U1530 (N_1530,N_833,In_2793);
and U1531 (N_1531,In_1028,N_1141);
nand U1532 (N_1532,In_328,N_628);
nor U1533 (N_1533,N_613,N_168);
xnor U1534 (N_1534,N_1106,N_988);
nor U1535 (N_1535,N_323,In_1964);
or U1536 (N_1536,N_400,N_297);
or U1537 (N_1537,In_863,N_810);
xnor U1538 (N_1538,In_101,N_877);
nand U1539 (N_1539,N_812,N_1190);
nand U1540 (N_1540,N_1006,In_2828);
xor U1541 (N_1541,N_1056,N_829);
or U1542 (N_1542,N_944,N_1195);
and U1543 (N_1543,In_1102,N_1102);
or U1544 (N_1544,In_2330,In_1489);
or U1545 (N_1545,In_81,N_970);
xnor U1546 (N_1546,N_759,N_547);
xnor U1547 (N_1547,N_1076,N_81);
and U1548 (N_1548,In_2369,N_837);
xnor U1549 (N_1549,N_1192,N_740);
nor U1550 (N_1550,In_2823,N_464);
nor U1551 (N_1551,N_751,N_1059);
xor U1552 (N_1552,In_2884,In_881);
nand U1553 (N_1553,In_485,In_518);
nor U1554 (N_1554,N_971,N_483);
nor U1555 (N_1555,N_966,N_3);
and U1556 (N_1556,In_240,N_765);
nor U1557 (N_1557,In_1549,N_324);
nand U1558 (N_1558,In_293,N_807);
nand U1559 (N_1559,In_266,N_822);
and U1560 (N_1560,N_843,N_627);
and U1561 (N_1561,In_2792,N_1074);
or U1562 (N_1562,In_1733,N_555);
nand U1563 (N_1563,N_1156,In_379);
and U1564 (N_1564,In_533,N_994);
nor U1565 (N_1565,N_387,N_113);
nor U1566 (N_1566,In_2612,N_2);
nor U1567 (N_1567,N_359,In_629);
nor U1568 (N_1568,In_2104,N_474);
nor U1569 (N_1569,In_2800,In_1835);
or U1570 (N_1570,In_1423,In_493);
nor U1571 (N_1571,In_1326,In_809);
or U1572 (N_1572,In_1227,In_1823);
nor U1573 (N_1573,N_689,In_2486);
nand U1574 (N_1574,In_1818,In_232);
nand U1575 (N_1575,N_996,In_920);
xnor U1576 (N_1576,In_1679,N_840);
xor U1577 (N_1577,In_2821,N_906);
or U1578 (N_1578,N_766,In_2024);
xor U1579 (N_1579,N_724,In_2126);
nor U1580 (N_1580,In_979,N_1060);
nand U1581 (N_1581,In_861,N_1132);
nor U1582 (N_1582,In_1437,N_678);
or U1583 (N_1583,N_1199,N_743);
xnor U1584 (N_1584,N_460,In_2275);
xnor U1585 (N_1585,N_902,N_708);
nand U1586 (N_1586,N_790,In_584);
and U1587 (N_1587,In_2899,In_918);
and U1588 (N_1588,N_89,N_793);
nand U1589 (N_1589,In_2997,In_2191);
xnor U1590 (N_1590,In_1171,N_536);
or U1591 (N_1591,In_356,In_2433);
nand U1592 (N_1592,In_287,In_2316);
nand U1593 (N_1593,N_748,In_763);
or U1594 (N_1594,In_633,N_982);
and U1595 (N_1595,In_390,In_1984);
nand U1596 (N_1596,In_2326,In_974);
nand U1597 (N_1597,N_1015,In_1105);
nand U1598 (N_1598,In_2462,N_343);
nand U1599 (N_1599,N_534,In_2160);
nor U1600 (N_1600,N_862,In_611);
nand U1601 (N_1601,N_1103,N_486);
nand U1602 (N_1602,In_2005,N_1188);
or U1603 (N_1603,N_629,N_234);
or U1604 (N_1604,In_2963,In_2587);
nand U1605 (N_1605,N_755,N_608);
or U1606 (N_1606,In_2417,In_1084);
nand U1607 (N_1607,N_1139,N_562);
or U1608 (N_1608,In_2012,In_926);
or U1609 (N_1609,N_989,In_2702);
xnor U1610 (N_1610,N_846,In_1671);
and U1611 (N_1611,N_128,N_1197);
xnor U1612 (N_1612,In_1055,In_224);
or U1613 (N_1613,N_637,N_799);
or U1614 (N_1614,In_2414,In_1389);
and U1615 (N_1615,In_1947,In_1801);
nand U1616 (N_1616,N_908,N_422);
nor U1617 (N_1617,In_248,N_1071);
nor U1618 (N_1618,In_1753,In_2774);
nor U1619 (N_1619,N_236,In_107);
and U1620 (N_1620,In_827,In_1373);
or U1621 (N_1621,In_1325,N_361);
or U1622 (N_1622,N_964,N_385);
or U1623 (N_1623,N_539,In_947);
nor U1624 (N_1624,In_862,In_1039);
xnor U1625 (N_1625,In_2129,N_333);
nand U1626 (N_1626,N_521,N_792);
nor U1627 (N_1627,In_449,N_1033);
nor U1628 (N_1628,N_666,In_2291);
xor U1629 (N_1629,N_1080,In_2937);
or U1630 (N_1630,In_383,N_278);
and U1631 (N_1631,N_54,N_749);
or U1632 (N_1632,In_55,In_410);
nor U1633 (N_1633,In_2747,In_62);
or U1634 (N_1634,N_643,N_729);
and U1635 (N_1635,In_192,In_1288);
or U1636 (N_1636,N_159,In_2844);
nor U1637 (N_1637,N_44,N_889);
or U1638 (N_1638,N_43,In_2138);
or U1639 (N_1639,N_706,N_227);
or U1640 (N_1640,In_1120,In_1675);
nor U1641 (N_1641,In_2764,N_884);
nor U1642 (N_1642,In_998,In_1684);
nand U1643 (N_1643,N_774,In_1855);
or U1644 (N_1644,N_764,In_655);
or U1645 (N_1645,N_1005,N_671);
nand U1646 (N_1646,In_230,In_1376);
and U1647 (N_1647,N_418,N_328);
nand U1648 (N_1648,In_702,N_1158);
or U1649 (N_1649,N_998,N_71);
nor U1650 (N_1650,In_628,In_1595);
nand U1651 (N_1651,N_1126,N_1084);
xnor U1652 (N_1652,N_296,N_85);
xor U1653 (N_1653,In_2239,N_1178);
and U1654 (N_1654,In_523,N_888);
and U1655 (N_1655,In_256,N_48);
xnor U1656 (N_1656,N_611,N_623);
xnor U1657 (N_1657,In_2373,N_716);
xor U1658 (N_1658,N_762,N_1024);
nor U1659 (N_1659,In_2608,In_84);
and U1660 (N_1660,In_2205,In_2605);
and U1661 (N_1661,N_354,N_991);
or U1662 (N_1662,In_2312,In_937);
nand U1663 (N_1663,In_1059,In_2935);
and U1664 (N_1664,In_179,In_2942);
and U1665 (N_1665,In_464,N_857);
nand U1666 (N_1666,N_852,In_1447);
nor U1667 (N_1667,In_166,In_1020);
and U1668 (N_1668,N_694,In_1042);
and U1669 (N_1669,N_235,In_1088);
nor U1670 (N_1670,In_2332,In_1390);
and U1671 (N_1671,In_2653,N_228);
nand U1672 (N_1672,In_758,In_2618);
or U1673 (N_1673,N_1064,N_1148);
and U1674 (N_1674,N_938,N_656);
nor U1675 (N_1675,N_620,N_20);
nor U1676 (N_1676,In_1534,N_596);
or U1677 (N_1677,N_581,N_796);
nand U1678 (N_1678,In_977,In_2154);
and U1679 (N_1679,In_2826,In_2427);
nand U1680 (N_1680,In_1791,N_457);
or U1681 (N_1681,N_670,N_979);
xnor U1682 (N_1682,In_1763,N_712);
and U1683 (N_1683,N_314,In_2637);
and U1684 (N_1684,N_897,N_69);
nor U1685 (N_1685,In_2616,N_1198);
xor U1686 (N_1686,N_1172,In_1998);
nand U1687 (N_1687,N_1051,In_2882);
nor U1688 (N_1688,N_881,In_2546);
nor U1689 (N_1689,N_485,In_1179);
or U1690 (N_1690,N_1013,In_2907);
nor U1691 (N_1691,In_2967,In_1509);
nor U1692 (N_1692,In_1305,In_1546);
and U1693 (N_1693,N_750,In_574);
xnor U1694 (N_1694,N_786,N_803);
or U1695 (N_1695,In_1438,N_355);
or U1696 (N_1696,N_386,N_496);
nor U1697 (N_1697,In_280,N_1031);
nor U1698 (N_1698,N_872,N_1053);
or U1699 (N_1699,N_717,N_1078);
nor U1700 (N_1700,N_973,In_2676);
xor U1701 (N_1701,N_1189,In_302);
nor U1702 (N_1702,In_2418,In_2047);
xnor U1703 (N_1703,N_1129,N_1090);
or U1704 (N_1704,N_675,In_906);
nand U1705 (N_1705,In_1196,N_25);
xnor U1706 (N_1706,In_788,In_551);
or U1707 (N_1707,N_1116,In_2983);
nor U1708 (N_1708,In_1741,In_515);
nor U1709 (N_1709,N_945,In_1696);
nor U1710 (N_1710,In_1669,N_1038);
xnor U1711 (N_1711,In_1800,In_2969);
and U1712 (N_1712,N_82,In_292);
nand U1713 (N_1713,N_340,In_2107);
nand U1714 (N_1714,In_2172,In_1017);
nand U1715 (N_1715,In_685,N_1052);
xnor U1716 (N_1716,In_2707,In_1384);
xnor U1717 (N_1717,N_41,In_1564);
and U1718 (N_1718,N_469,In_1057);
nor U1719 (N_1719,In_2366,N_475);
or U1720 (N_1720,N_640,N_1130);
nor U1721 (N_1721,In_2311,N_726);
or U1722 (N_1722,N_1001,N_590);
xnor U1723 (N_1723,N_626,N_560);
or U1724 (N_1724,In_419,In_1729);
nand U1725 (N_1725,N_377,N_636);
nor U1726 (N_1726,N_1034,In_2924);
nor U1727 (N_1727,In_737,In_279);
nand U1728 (N_1728,In_2868,N_849);
nand U1729 (N_1729,In_1762,In_621);
nor U1730 (N_1730,N_882,N_747);
nor U1731 (N_1731,In_2765,N_697);
xnor U1732 (N_1732,In_2411,N_435);
xor U1733 (N_1733,N_1186,N_887);
nand U1734 (N_1734,In_1648,N_851);
nor U1735 (N_1735,N_0,In_1773);
nor U1736 (N_1736,N_756,In_1601);
nor U1737 (N_1737,In_1263,In_1891);
nor U1738 (N_1738,In_1771,N_391);
and U1739 (N_1739,In_1238,In_1915);
nor U1740 (N_1740,In_2288,N_545);
or U1741 (N_1741,N_702,In_1198);
or U1742 (N_1742,In_2761,N_1122);
or U1743 (N_1743,N_591,In_2232);
nor U1744 (N_1744,N_110,In_2425);
xor U1745 (N_1745,In_902,N_189);
xor U1746 (N_1746,N_936,In_310);
xnor U1747 (N_1747,N_624,In_2569);
nand U1748 (N_1748,In_569,In_2444);
xor U1749 (N_1749,N_919,N_763);
nor U1750 (N_1750,N_404,In_661);
or U1751 (N_1751,N_710,In_1035);
or U1752 (N_1752,N_269,N_489);
or U1753 (N_1753,In_598,In_828);
and U1754 (N_1754,N_1050,N_1118);
and U1755 (N_1755,In_2391,In_1019);
nand U1756 (N_1756,N_371,N_682);
nand U1757 (N_1757,N_412,In_2233);
or U1758 (N_1758,N_669,N_232);
nand U1759 (N_1759,In_7,In_1660);
or U1760 (N_1760,N_825,N_451);
or U1761 (N_1761,N_564,N_738);
and U1762 (N_1762,In_1788,In_2457);
or U1763 (N_1763,N_566,N_1020);
nor U1764 (N_1764,In_1130,In_1200);
and U1765 (N_1765,In_1712,N_1194);
or U1766 (N_1766,N_388,In_2626);
and U1767 (N_1767,In_941,In_2972);
nor U1768 (N_1768,In_1416,In_337);
nand U1769 (N_1769,In_2389,In_1331);
or U1770 (N_1770,N_1137,N_1160);
xnor U1771 (N_1771,N_1077,N_307);
xor U1772 (N_1772,N_1187,In_2949);
or U1773 (N_1773,In_886,N_942);
xnor U1774 (N_1774,N_525,In_148);
nand U1775 (N_1775,In_217,In_1044);
or U1776 (N_1776,N_736,N_12);
and U1777 (N_1777,N_281,N_197);
nor U1778 (N_1778,N_1171,In_2297);
nor U1779 (N_1779,In_157,N_1166);
nor U1780 (N_1780,In_578,In_966);
xor U1781 (N_1781,N_287,N_476);
nor U1782 (N_1782,N_1108,N_946);
and U1783 (N_1783,N_1027,In_1021);
xor U1784 (N_1784,In_2180,In_787);
nand U1785 (N_1785,N_834,In_2819);
xor U1786 (N_1786,In_869,In_2568);
xor U1787 (N_1787,In_463,N_368);
and U1788 (N_1788,N_1133,In_1508);
nand U1789 (N_1789,N_861,N_821);
and U1790 (N_1790,In_1977,In_159);
xnor U1791 (N_1791,In_1779,In_2953);
or U1792 (N_1792,In_774,In_1483);
nand U1793 (N_1793,In_261,N_757);
and U1794 (N_1794,N_1127,In_2836);
nor U1795 (N_1795,N_1035,In_298);
xnor U1796 (N_1796,In_1098,In_2745);
or U1797 (N_1797,N_867,N_869);
nand U1798 (N_1798,In_2392,N_1091);
and U1799 (N_1799,N_424,N_61);
nand U1800 (N_1800,N_1627,N_1332);
and U1801 (N_1801,N_1612,N_1500);
xnor U1802 (N_1802,N_1458,N_1559);
and U1803 (N_1803,N_201,N_1402);
xnor U1804 (N_1804,In_2163,N_1355);
or U1805 (N_1805,N_1630,N_836);
and U1806 (N_1806,In_2162,N_1554);
and U1807 (N_1807,N_1562,N_1294);
xor U1808 (N_1808,N_1359,N_1256);
nand U1809 (N_1809,N_1377,In_1218);
or U1810 (N_1810,In_892,N_506);
and U1811 (N_1811,In_117,N_188);
nor U1812 (N_1812,N_1760,N_1777);
or U1813 (N_1813,N_1254,N_1415);
and U1814 (N_1814,In_1865,In_2838);
xnor U1815 (N_1815,N_1661,N_1633);
and U1816 (N_1816,N_701,In_710);
xor U1817 (N_1817,N_1708,N_1596);
and U1818 (N_1818,N_841,In_1577);
nand U1819 (N_1819,N_1350,N_990);
nor U1820 (N_1820,N_1292,In_2776);
xor U1821 (N_1821,N_1517,N_1602);
nor U1822 (N_1822,In_164,N_1134);
nor U1823 (N_1823,In_1525,N_933);
nor U1824 (N_1824,N_1617,N_1671);
xor U1825 (N_1825,N_1484,In_1026);
and U1826 (N_1826,In_1925,N_1308);
nor U1827 (N_1827,In_2553,N_1358);
and U1828 (N_1828,N_1289,N_1726);
or U1829 (N_1829,In_1514,N_806);
and U1830 (N_1830,N_1681,N_1576);
or U1831 (N_1831,N_1455,In_1879);
and U1832 (N_1832,In_2685,In_819);
or U1833 (N_1833,In_2515,In_336);
xnor U1834 (N_1834,N_1664,N_1326);
nand U1835 (N_1835,N_1683,N_1104);
and U1836 (N_1836,N_1419,N_1548);
and U1837 (N_1837,In_1143,N_196);
nor U1838 (N_1838,N_1678,N_1336);
nand U1839 (N_1839,N_692,N_65);
nor U1840 (N_1840,N_1618,N_1790);
and U1841 (N_1841,N_1776,In_2646);
nand U1842 (N_1842,In_223,N_1516);
and U1843 (N_1843,N_896,N_75);
or U1844 (N_1844,N_1522,N_33);
xnor U1845 (N_1845,N_777,N_1648);
nand U1846 (N_1846,N_1298,N_1004);
or U1847 (N_1847,N_1061,N_66);
and U1848 (N_1848,N_1304,N_809);
nand U1849 (N_1849,N_1729,N_1026);
or U1850 (N_1850,In_705,In_112);
nor U1851 (N_1851,In_1078,N_1333);
or U1852 (N_1852,N_1315,In_2513);
xnor U1853 (N_1853,N_268,N_703);
nor U1854 (N_1854,N_850,N_1736);
and U1855 (N_1855,N_1016,N_1208);
xnor U1856 (N_1856,In_1656,N_1454);
nor U1857 (N_1857,N_1267,N_741);
or U1858 (N_1858,N_1244,N_1501);
nand U1859 (N_1859,N_1518,In_2334);
nand U1860 (N_1860,N_1036,N_1344);
nor U1861 (N_1861,N_1378,N_524);
or U1862 (N_1862,In_552,In_1114);
nand U1863 (N_1863,N_1374,N_617);
nand U1864 (N_1864,N_1204,N_771);
xnor U1865 (N_1865,N_1438,N_1641);
nor U1866 (N_1866,In_2971,N_1673);
xnor U1867 (N_1867,N_1397,N_1669);
or U1868 (N_1868,N_1619,N_1698);
nor U1869 (N_1869,In_538,N_1218);
or U1870 (N_1870,N_1223,N_1423);
xnor U1871 (N_1871,N_1622,In_1014);
nand U1872 (N_1872,N_1589,N_633);
xnor U1873 (N_1873,N_1573,N_1498);
or U1874 (N_1874,N_1734,N_1070);
nand U1875 (N_1875,In_1296,N_1262);
or U1876 (N_1876,N_317,N_1590);
nor U1877 (N_1877,In_1056,N_1381);
xor U1878 (N_1878,N_1329,N_745);
xnor U1879 (N_1879,N_1068,In_1785);
xnor U1880 (N_1880,N_1372,N_248);
and U1881 (N_1881,N_1351,N_293);
or U1882 (N_1882,In_1933,N_976);
xor U1883 (N_1883,N_1369,In_2150);
nor U1884 (N_1884,N_1561,N_858);
xnor U1885 (N_1885,In_1111,N_1079);
xnor U1886 (N_1886,N_1278,N_428);
nor U1887 (N_1887,In_1340,N_1525);
xnor U1888 (N_1888,N_728,In_27);
xor U1889 (N_1889,N_1528,N_1583);
nor U1890 (N_1890,N_1566,N_551);
nor U1891 (N_1891,N_1555,N_1660);
and U1892 (N_1892,N_1183,N_1135);
and U1893 (N_1893,N_1721,In_285);
nand U1894 (N_1894,N_1082,N_1636);
or U1895 (N_1895,In_2919,N_1650);
and U1896 (N_1896,N_1485,N_1462);
xor U1897 (N_1897,N_1788,N_1609);
xor U1898 (N_1898,N_1690,N_997);
or U1899 (N_1899,N_1626,In_853);
or U1900 (N_1900,In_2085,N_1021);
or U1901 (N_1901,N_1774,N_1069);
and U1902 (N_1902,N_650,N_635);
and U1903 (N_1903,In_2502,In_29);
xor U1904 (N_1904,N_1715,N_788);
and U1905 (N_1905,In_2350,N_1496);
xnor U1906 (N_1906,In_1623,N_1713);
and U1907 (N_1907,In_2203,N_686);
nor U1908 (N_1908,In_1352,N_1523);
and U1909 (N_1909,N_776,In_2743);
nand U1910 (N_1910,N_1580,N_31);
and U1911 (N_1911,In_220,N_443);
nor U1912 (N_1912,N_1764,N_1295);
or U1913 (N_1913,N_1686,N_1724);
nor U1914 (N_1914,N_1635,N_1280);
and U1915 (N_1915,In_1314,N_954);
nand U1916 (N_1916,In_44,In_37);
xnor U1917 (N_1917,In_161,N_330);
and U1918 (N_1918,N_730,N_1260);
nand U1919 (N_1919,N_684,N_856);
and U1920 (N_1920,N_1317,N_1117);
xnor U1921 (N_1921,N_1339,N_1533);
or U1922 (N_1922,In_1178,In_1633);
xnor U1923 (N_1923,In_824,In_2447);
xor U1924 (N_1924,N_744,N_1491);
xor U1925 (N_1925,N_1413,N_1416);
and U1926 (N_1926,N_1342,N_205);
nand U1927 (N_1927,N_917,N_1709);
nand U1928 (N_1928,In_197,In_1836);
nand U1929 (N_1929,N_1387,N_1623);
and U1930 (N_1930,N_632,N_1679);
or U1931 (N_1931,N_1530,N_1412);
or U1932 (N_1932,N_1565,N_1795);
and U1933 (N_1933,N_1014,N_157);
xnor U1934 (N_1934,N_1752,N_1328);
and U1935 (N_1935,In_2079,In_1260);
nor U1936 (N_1936,N_1546,In_2986);
nand U1937 (N_1937,In_1683,N_1282);
xnor U1938 (N_1938,N_1780,N_767);
nor U1939 (N_1939,N_1607,N_1442);
nor U1940 (N_1940,N_1285,N_1452);
nand U1941 (N_1941,N_1539,N_1376);
nor U1942 (N_1942,N_1275,In_577);
or U1943 (N_1943,N_972,N_1732);
or U1944 (N_1944,N_1088,In_1602);
nand U1945 (N_1945,N_713,In_1840);
xnor U1946 (N_1946,N_1560,N_1081);
or U1947 (N_1947,N_30,In_856);
nor U1948 (N_1948,In_51,N_253);
xnor U1949 (N_1949,N_559,N_1731);
xor U1950 (N_1950,N_334,In_2966);
and U1951 (N_1951,In_1524,In_1464);
nand U1952 (N_1952,N_1318,In_714);
nand U1953 (N_1953,N_1449,N_1408);
or U1954 (N_1954,N_1476,N_727);
nand U1955 (N_1955,N_797,N_1233);
nand U1956 (N_1956,N_1779,In_1212);
nand U1957 (N_1957,In_1269,N_1386);
and U1958 (N_1958,N_1433,N_1364);
xnor U1959 (N_1959,N_1446,N_1274);
and U1960 (N_1960,N_874,In_2705);
and U1961 (N_1961,N_1743,In_2026);
or U1962 (N_1962,N_668,In_1658);
or U1963 (N_1963,N_1206,N_263);
nand U1964 (N_1964,N_1640,N_1603);
nand U1965 (N_1965,N_1549,N_1401);
or U1966 (N_1966,N_1791,N_1771);
or U1967 (N_1967,N_1424,N_327);
nor U1968 (N_1968,N_1346,N_1582);
or U1969 (N_1969,N_290,In_391);
nand U1970 (N_1970,N_1577,N_1018);
xnor U1971 (N_1971,N_1757,N_1751);
or U1972 (N_1972,In_2403,In_915);
or U1973 (N_1973,N_1793,N_1502);
nor U1974 (N_1974,In_24,N_288);
nor U1975 (N_1975,N_1272,N_1651);
or U1976 (N_1976,N_1579,N_769);
nor U1977 (N_1977,N_1434,N_1427);
and U1978 (N_1978,N_1353,N_1365);
or U1979 (N_1979,N_1472,In_1270);
and U1980 (N_1980,N_1537,In_275);
xor U1981 (N_1981,N_1400,N_1331);
nor U1982 (N_1982,N_280,N_1322);
and U1983 (N_1983,N_859,N_481);
nor U1984 (N_1984,N_1347,In_479);
and U1985 (N_1985,In_2402,N_956);
nand U1986 (N_1986,In_2376,N_1781);
nand U1987 (N_1987,In_144,N_610);
or U1988 (N_1988,N_1456,In_1521);
or U1989 (N_1989,N_1207,In_2190);
xor U1990 (N_1990,N_1391,N_1169);
and U1991 (N_1991,In_221,N_1425);
or U1992 (N_1992,N_1363,N_254);
or U1993 (N_1993,N_1615,N_968);
nand U1994 (N_1994,N_1073,N_828);
or U1995 (N_1995,N_1535,N_1055);
xnor U1996 (N_1996,N_1265,N_1023);
xor U1997 (N_1997,In_502,In_1655);
xnor U1998 (N_1998,N_1538,N_1527);
nand U1999 (N_1999,N_1393,N_1324);
nor U2000 (N_2000,In_2548,N_1741);
and U2001 (N_2001,In_766,N_1513);
nand U2002 (N_2002,N_270,N_1120);
nor U2003 (N_2003,N_1682,In_2848);
xor U2004 (N_2004,N_999,In_688);
and U2005 (N_2005,N_1464,In_102);
and U2006 (N_2006,In_539,N_1493);
and U2007 (N_2007,N_1613,In_2810);
and U2008 (N_2008,N_1421,N_1700);
nor U2009 (N_2009,N_519,In_1115);
nor U2010 (N_2010,In_2600,In_2607);
nor U2011 (N_2011,N_823,N_873);
and U2012 (N_2012,N_1778,N_36);
nand U2013 (N_2013,N_127,N_298);
or U2014 (N_2014,In_1586,In_675);
xnor U2015 (N_2015,N_1587,N_1341);
or U2016 (N_2016,In_1715,N_1634);
xnor U2017 (N_2017,N_928,N_286);
nand U2018 (N_2018,N_1211,In_2153);
and U2019 (N_2019,N_1695,N_1758);
and U2020 (N_2020,N_1490,N_1154);
nor U2021 (N_2021,N_1054,In_396);
nor U2022 (N_2022,In_2859,N_1145);
or U2023 (N_2023,N_1608,N_1281);
nand U2024 (N_2024,N_1478,In_353);
or U2025 (N_2025,N_1799,In_2614);
xor U2026 (N_2026,N_1345,N_55);
nor U2027 (N_2027,N_1146,In_1174);
nand U2028 (N_2028,N_875,In_894);
nand U2029 (N_2029,N_1578,N_1762);
nand U2030 (N_2030,N_1655,N_1745);
and U2031 (N_2031,N_1234,N_1563);
xor U2032 (N_2032,In_1661,N_1246);
nand U2033 (N_2033,N_1136,N_1212);
nand U2034 (N_2034,N_1571,N_1629);
xnor U2035 (N_2035,In_1303,N_1658);
and U2036 (N_2036,N_916,N_1058);
nor U2037 (N_2037,N_1646,N_711);
nor U2038 (N_2038,N_1654,In_543);
nor U2039 (N_2039,N_1665,In_1725);
or U2040 (N_2040,N_1049,N_1335);
and U2041 (N_2041,In_864,N_677);
nor U2042 (N_2042,N_1180,N_1453);
nor U2043 (N_2043,In_555,N_1092);
xor U2044 (N_2044,N_1691,N_319);
and U2045 (N_2045,N_1642,In_1728);
nand U2046 (N_2046,N_125,N_1540);
or U2047 (N_2047,N_947,In_2468);
xnor U2048 (N_2048,In_1073,In_1502);
or U2049 (N_2049,N_1477,In_2842);
nand U2050 (N_2050,N_484,N_1570);
nand U2051 (N_2051,In_1165,N_200);
and U2052 (N_2052,N_920,In_1992);
nand U2053 (N_2053,In_905,N_1475);
nor U2054 (N_2054,In_522,N_45);
nand U2055 (N_2055,N_1529,N_1725);
nor U2056 (N_2056,In_739,N_1542);
nor U2057 (N_2057,In_371,N_1699);
and U2058 (N_2058,N_342,N_848);
xnor U2059 (N_2059,N_601,N_1763);
or U2060 (N_2060,N_1149,N_1459);
nand U2061 (N_2061,N_737,N_1247);
xor U2062 (N_2062,N_625,N_1266);
nand U2063 (N_2063,N_1486,N_1524);
nor U2064 (N_2064,N_1371,N_1270);
and U2065 (N_2065,N_543,In_272);
or U2066 (N_2066,In_2323,N_1722);
nor U2067 (N_2067,In_477,In_52);
nand U2068 (N_2068,N_1514,In_1821);
and U2069 (N_2069,N_1675,N_1783);
nor U2070 (N_2070,N_987,N_1046);
and U2071 (N_2071,N_1659,N_865);
and U2072 (N_2072,N_1653,N_1742);
and U2073 (N_2073,In_1254,N_1775);
xor U2074 (N_2074,N_396,N_1604);
nand U2075 (N_2075,N_960,N_1382);
xnor U2076 (N_2076,N_965,In_831);
and U2077 (N_2077,N_1313,In_534);
xor U2078 (N_2078,N_1689,N_731);
xor U2079 (N_2079,In_2197,N_725);
or U2080 (N_2080,In_2057,N_1754);
nand U2081 (N_2081,N_984,In_402);
xor U2082 (N_2082,N_1447,In_1463);
xor U2083 (N_2083,N_1744,N_1787);
nand U2084 (N_2084,N_1553,In_1560);
xor U2085 (N_2085,N_177,N_1319);
nand U2086 (N_2086,N_39,N_1644);
xor U2087 (N_2087,In_1054,N_775);
nor U2088 (N_2088,N_1383,N_1672);
and U2089 (N_2089,N_1767,N_1309);
or U2090 (N_2090,In_2149,In_698);
and U2091 (N_2091,N_892,N_949);
xor U2092 (N_2092,N_1738,N_926);
xnor U2093 (N_2093,N_1759,N_925);
and U2094 (N_2094,N_1259,N_1296);
nand U2095 (N_2095,N_1588,N_657);
or U2096 (N_2096,N_696,N_1239);
xnor U2097 (N_2097,N_679,N_1503);
xor U2098 (N_2098,N_1547,N_1214);
nor U2099 (N_2099,In_498,N_1394);
nand U2100 (N_2100,N_1568,N_222);
and U2101 (N_2101,In_1284,In_377);
and U2102 (N_2102,N_1461,In_822);
nor U2103 (N_2103,N_723,In_2636);
and U2104 (N_2104,In_2887,N_1789);
and U2105 (N_2105,N_983,N_1151);
nand U2106 (N_2106,N_907,N_537);
or U2107 (N_2107,N_1794,N_1210);
xor U2108 (N_2108,In_626,N_1228);
and U2109 (N_2109,N_1473,N_277);
xnor U2110 (N_2110,In_935,N_1242);
or U2111 (N_2111,N_1704,N_958);
and U2112 (N_2112,In_970,In_1244);
xor U2113 (N_2113,N_1017,N_1610);
or U2114 (N_2114,N_1111,N_1747);
nand U2115 (N_2115,N_1599,N_1506);
xnor U2116 (N_2116,N_1688,N_779);
or U2117 (N_2117,N_1483,N_1288);
nor U2118 (N_2118,In_1145,In_2990);
and U2119 (N_2119,N_1385,N_1652);
nor U2120 (N_2120,N_1448,In_8);
or U2121 (N_2121,N_1311,N_1600);
and U2122 (N_2122,N_1720,In_2426);
xor U2123 (N_2123,N_1222,In_1873);
nand U2124 (N_2124,N_1354,N_1357);
or U2125 (N_2125,In_1328,In_1910);
or U2126 (N_2126,N_1666,N_1645);
nand U2127 (N_2127,N_1249,N_1263);
or U2128 (N_2128,In_420,N_1586);
nand U2129 (N_2129,N_499,N_1569);
nor U2130 (N_2130,In_2243,In_0);
nand U2131 (N_2131,In_2584,N_1723);
nand U2132 (N_2132,N_1361,N_1238);
or U2133 (N_2133,N_1676,In_2854);
nand U2134 (N_2134,N_1255,N_1268);
nand U2135 (N_2135,N_995,N_1420);
or U2136 (N_2136,N_1403,N_1598);
nor U2137 (N_2137,In_15,N_1209);
or U2138 (N_2138,N_1432,N_1306);
and U2139 (N_2139,N_1511,In_2872);
xnor U2140 (N_2140,In_1852,In_85);
nand U2141 (N_2141,N_1417,In_1442);
or U2142 (N_2142,N_1521,N_1414);
or U2143 (N_2143,N_1436,N_194);
nor U2144 (N_2144,N_1657,N_1440);
and U2145 (N_2145,N_1782,In_2973);
or U2146 (N_2146,N_1597,In_2640);
or U2147 (N_2147,N_1662,N_1410);
nand U2148 (N_2148,N_1301,N_1094);
and U2149 (N_2149,N_1110,N_64);
xnor U2150 (N_2150,N_801,In_2865);
xor U2151 (N_2151,N_957,N_864);
and U2152 (N_2152,N_1656,N_1325);
nor U2153 (N_2153,N_930,N_1277);
nor U2154 (N_2154,N_1470,In_183);
nand U2155 (N_2155,N_1167,N_1739);
xnor U2156 (N_2156,N_1241,In_2123);
xnor U2157 (N_2157,N_1221,N_1668);
or U2158 (N_2158,N_1445,N_1457);
nor U2159 (N_2159,N_939,N_1718);
or U2160 (N_2160,In_636,N_1591);
or U2161 (N_2161,In_2623,N_395);
nor U2162 (N_2162,In_985,N_1380);
nand U2163 (N_2163,N_1029,In_1452);
and U2164 (N_2164,N_1340,In_916);
and U2165 (N_2165,N_1235,N_1287);
nor U2166 (N_2166,N_1231,N_967);
xor U2167 (N_2167,In_877,N_1443);
nor U2168 (N_2168,N_1431,N_1240);
or U2169 (N_2169,In_2011,N_1220);
nor U2170 (N_2170,N_1405,N_1245);
nor U2171 (N_2171,In_1266,In_364);
nand U2172 (N_2172,N_885,N_630);
xnor U2173 (N_2173,In_2270,In_1672);
nor U2174 (N_2174,N_1362,N_245);
nand U2175 (N_2175,N_1307,N_1687);
nor U2176 (N_2176,In_1158,N_1439);
nand U2177 (N_2177,N_1711,In_151);
nor U2178 (N_2178,N_1515,N_1677);
or U2179 (N_2179,N_1388,N_1392);
nand U2180 (N_2180,N_1705,N_224);
nand U2181 (N_2181,N_1426,N_1494);
nand U2182 (N_2182,In_444,N_498);
or U2183 (N_2183,N_1567,N_1585);
and U2184 (N_2184,N_811,In_2576);
nor U2185 (N_2185,N_1463,N_1581);
xor U2186 (N_2186,N_1112,N_802);
xor U2187 (N_2187,N_118,In_1991);
or U2188 (N_2188,N_658,N_1601);
and U2189 (N_2189,N_1343,In_2939);
nand U2190 (N_2190,N_663,N_1482);
nand U2191 (N_2191,N_1200,N_975);
nand U2192 (N_2192,N_1230,N_26);
nor U2193 (N_2193,In_2936,N_935);
xnor U2194 (N_2194,N_977,In_1443);
nor U2195 (N_2195,In_973,N_1526);
nor U2196 (N_2196,N_1356,N_1786);
or U2197 (N_2197,In_1203,N_393);
or U2198 (N_2198,N_1283,N_1250);
nand U2199 (N_2199,N_1334,In_706);
or U2200 (N_2200,N_1628,N_758);
nor U2201 (N_2201,N_1113,N_662);
nor U2202 (N_2202,In_2714,N_969);
or U2203 (N_2203,In_1736,N_1670);
nand U2204 (N_2204,N_1248,N_1552);
or U2205 (N_2205,N_1253,In_2687);
nand U2206 (N_2206,In_93,N_1302);
nand U2207 (N_2207,In_1557,N_1727);
nor U2208 (N_2208,In_2045,N_1753);
and U2209 (N_2209,N_1418,N_1625);
nand U2210 (N_2210,In_2999,N_1205);
nor U2211 (N_2211,N_1466,N_306);
xnor U2212 (N_2212,N_1766,In_142);
nor U2213 (N_2213,In_722,N_1019);
nor U2214 (N_2214,N_1251,N_1606);
and U2215 (N_2215,N_1703,N_1202);
nor U2216 (N_2216,In_1320,N_1303);
nor U2217 (N_2217,N_580,N_1243);
and U2218 (N_2218,In_1360,In_1909);
nand U2219 (N_2219,N_339,N_426);
nand U2220 (N_2220,In_1890,N_1798);
and U2221 (N_2221,In_2065,N_1685);
nand U2222 (N_2222,N_1232,N_1226);
or U2223 (N_2223,In_2193,N_1163);
and U2224 (N_2224,N_681,N_1271);
nor U2225 (N_2225,N_832,N_830);
or U2226 (N_2226,N_667,N_1437);
nand U2227 (N_2227,N_826,N_1225);
and U2228 (N_2228,In_1738,N_1203);
or U2229 (N_2229,N_1749,In_972);
and U2230 (N_2230,N_680,N_1697);
and U2231 (N_2231,In_1493,In_1112);
or U2232 (N_2232,In_1011,In_363);
or U2233 (N_2233,N_1495,N_184);
nor U2234 (N_2234,N_1637,N_705);
and U2235 (N_2235,N_1785,N_870);
or U2236 (N_2236,N_1499,N_1614);
nand U2237 (N_2237,N_1093,N_912);
or U2238 (N_2238,N_1095,In_22);
nor U2239 (N_2239,In_2648,In_73);
and U2240 (N_2240,N_805,N_1509);
nor U2241 (N_2241,N_1730,N_653);
and U2242 (N_2242,N_1131,N_1488);
or U2243 (N_2243,N_1217,N_1100);
or U2244 (N_2244,In_2961,In_1312);
nor U2245 (N_2245,N_1373,N_660);
xor U2246 (N_2246,N_1284,N_1168);
or U2247 (N_2247,N_1536,N_1750);
xor U2248 (N_2248,N_1543,N_1216);
xor U2249 (N_2249,N_1680,In_54);
or U2250 (N_2250,N_1594,N_934);
xnor U2251 (N_2251,N_1575,N_217);
or U2252 (N_2252,N_1097,N_1701);
xor U2253 (N_2253,N_1411,In_1731);
or U2254 (N_2254,N_1398,N_614);
or U2255 (N_2255,N_1712,N_1692);
or U2256 (N_2256,N_937,N_1352);
xor U2257 (N_2257,N_379,N_1631);
nor U2258 (N_2258,N_1375,In_40);
nor U2259 (N_2259,N_1765,N_1684);
xor U2260 (N_2260,In_2830,N_1649);
nor U2261 (N_2261,N_1314,N_1505);
xor U2262 (N_2262,N_223,N_1707);
nand U2263 (N_2263,N_1770,In_2177);
xor U2264 (N_2264,N_914,N_1746);
or U2265 (N_2265,N_1395,N_1674);
or U2266 (N_2266,N_1384,In_712);
or U2267 (N_2267,N_654,N_1406);
and U2268 (N_2268,N_1286,N_1532);
or U2269 (N_2269,N_1176,N_1497);
and U2270 (N_2270,N_1293,N_798);
or U2271 (N_2271,N_1632,N_1072);
nor U2272 (N_2272,In_2880,N_1428);
and U2273 (N_2273,N_1468,N_674);
xor U2274 (N_2274,N_1702,N_1330);
xor U2275 (N_2275,N_1769,N_921);
or U2276 (N_2276,N_1215,N_1574);
and U2277 (N_2277,N_1276,N_1430);
xnor U2278 (N_2278,N_1279,In_168);
nand U2279 (N_2279,N_1327,N_1441);
nor U2280 (N_2280,N_1551,N_1663);
or U2281 (N_2281,N_1716,N_1469);
nor U2282 (N_2282,N_648,N_1310);
xor U2283 (N_2283,N_672,N_528);
and U2284 (N_2284,N_1465,N_1258);
xor U2285 (N_2285,N_1756,N_1492);
or U2286 (N_2286,In_1858,N_1227);
and U2287 (N_2287,In_447,N_1337);
and U2288 (N_2288,In_1401,N_1611);
and U2289 (N_2289,In_2662,N_1057);
and U2290 (N_2290,N_1504,In_486);
nor U2291 (N_2291,N_890,N_1300);
xor U2292 (N_2292,In_682,N_1556);
or U2293 (N_2293,In_1820,N_1768);
nand U2294 (N_2294,In_184,N_311);
and U2295 (N_2295,In_1522,In_2115);
nand U2296 (N_2296,N_1201,N_1450);
and U2297 (N_2297,N_251,N_718);
or U2298 (N_2298,N_1037,N_1321);
or U2299 (N_2299,N_411,N_909);
xnor U2300 (N_2300,N_1639,In_2841);
nor U2301 (N_2301,N_1121,N_690);
or U2302 (N_2302,N_1784,N_1291);
nand U2303 (N_2303,N_1545,N_1564);
nand U2304 (N_2304,N_1297,N_953);
nor U2305 (N_2305,N_1000,In_1167);
nor U2306 (N_2306,N_1508,N_720);
xnor U2307 (N_2307,In_2992,N_1368);
or U2308 (N_2308,N_659,N_1261);
and U2309 (N_2309,In_509,In_1952);
nor U2310 (N_2310,N_901,N_1595);
xor U2311 (N_2311,In_1922,N_1257);
nor U2312 (N_2312,In_2758,N_1165);
or U2313 (N_2313,N_1696,N_1796);
xnor U2314 (N_2314,N_1429,N_820);
nand U2315 (N_2315,In_2368,In_137);
and U2316 (N_2316,N_1422,In_2428);
nor U2317 (N_2317,N_1710,In_1348);
nand U2318 (N_2318,N_1593,N_1761);
nand U2319 (N_2319,N_1323,N_1507);
nand U2320 (N_2320,N_1320,N_1480);
nand U2321 (N_2321,N_1299,N_1219);
nor U2322 (N_2322,N_1755,In_2719);
nand U2323 (N_2323,N_1735,N_1620);
nand U2324 (N_2324,N_1512,N_1592);
nor U2325 (N_2325,N_1396,N_903);
and U2326 (N_2326,N_1213,N_1728);
nand U2327 (N_2327,In_1067,N_292);
or U2328 (N_2328,N_927,N_1316);
xnor U2329 (N_2329,In_1547,N_1125);
nand U2330 (N_2330,In_659,N_383);
nor U2331 (N_2331,N_1435,In_2212);
nor U2332 (N_2332,N_202,N_1534);
nand U2333 (N_2333,N_1733,In_1921);
and U2334 (N_2334,N_1460,In_553);
or U2335 (N_2335,N_1008,N_1667);
nand U2336 (N_2336,N_746,In_203);
and U2337 (N_2337,In_958,N_1474);
nand U2338 (N_2338,N_594,In_270);
xor U2339 (N_2339,N_1531,N_962);
and U2340 (N_2340,N_1717,N_1584);
xnor U2341 (N_2341,In_1945,N_1043);
nor U2342 (N_2342,In_891,In_2511);
nand U2343 (N_2343,N_1312,N_1273);
and U2344 (N_2344,N_1647,N_1616);
and U2345 (N_2345,N_1196,N_337);
nor U2346 (N_2346,N_144,N_1467);
and U2347 (N_2347,N_1541,N_992);
and U2348 (N_2348,N_1748,In_2599);
or U2349 (N_2349,N_784,N_1161);
nor U2350 (N_2350,N_1370,N_1719);
or U2351 (N_2351,N_116,In_2574);
nand U2352 (N_2352,N_1305,N_1714);
nand U2353 (N_2353,N_1182,In_2206);
xnor U2354 (N_2354,N_1290,In_451);
nand U2355 (N_2355,N_1269,In_1784);
or U2356 (N_2356,N_1404,N_1740);
and U2357 (N_2357,N_1621,N_1237);
nand U2358 (N_2358,N_1510,N_752);
nor U2359 (N_2359,In_883,In_2555);
nor U2360 (N_2360,In_446,N_652);
xnor U2361 (N_2361,N_1264,N_646);
and U2362 (N_2362,N_1557,N_1643);
or U2363 (N_2363,N_1550,N_1605);
and U2364 (N_2364,In_1994,In_2597);
xnor U2365 (N_2365,N_1797,N_495);
xnor U2366 (N_2366,N_1338,N_1451);
and U2367 (N_2367,N_1792,N_1624);
nor U2368 (N_2368,N_35,N_1042);
xor U2369 (N_2369,N_1519,N_1379);
nor U2370 (N_2370,In_369,N_1096);
nand U2371 (N_2371,In_2327,In_1045);
and U2372 (N_2372,N_1348,N_4);
nor U2373 (N_2373,N_838,N_1224);
nor U2374 (N_2374,N_1229,N_584);
and U2375 (N_2375,N_1349,In_2222);
or U2376 (N_2376,N_794,N_1399);
nand U2377 (N_2377,N_1409,N_1389);
xor U2378 (N_2378,N_1360,In_2506);
nor U2379 (N_2379,N_880,N_1638);
and U2380 (N_2380,N_1252,N_1366);
nor U2381 (N_2381,N_923,N_1737);
and U2382 (N_2382,N_1128,N_1694);
or U2383 (N_2383,N_602,N_198);
and U2384 (N_2384,In_1982,N_1773);
nand U2385 (N_2385,N_1025,N_138);
xnor U2386 (N_2386,N_1487,N_1471);
xor U2387 (N_2387,N_1706,N_1520);
and U2388 (N_2388,N_1444,In_2145);
or U2389 (N_2389,N_1407,N_1390);
xor U2390 (N_2390,In_2289,N_1772);
nand U2391 (N_2391,In_2720,N_1157);
or U2392 (N_2392,N_1544,N_1489);
xor U2393 (N_2393,In_2931,In_348);
xor U2394 (N_2394,N_1479,N_1558);
or U2395 (N_2395,N_734,N_1693);
or U2396 (N_2396,N_785,N_1481);
nor U2397 (N_2397,N_1367,N_1236);
and U2398 (N_2398,N_732,N_1572);
nor U2399 (N_2399,In_123,In_1482);
nand U2400 (N_2400,N_2032,N_1899);
nand U2401 (N_2401,N_2162,N_2232);
and U2402 (N_2402,N_2240,N_2226);
xnor U2403 (N_2403,N_2230,N_2269);
or U2404 (N_2404,N_2391,N_2354);
nor U2405 (N_2405,N_2197,N_1861);
or U2406 (N_2406,N_2255,N_2348);
or U2407 (N_2407,N_2059,N_1869);
xnor U2408 (N_2408,N_2022,N_2143);
or U2409 (N_2409,N_1975,N_2082);
nand U2410 (N_2410,N_2178,N_2218);
and U2411 (N_2411,N_2183,N_2243);
or U2412 (N_2412,N_1888,N_2170);
xor U2413 (N_2413,N_2261,N_2225);
nand U2414 (N_2414,N_1843,N_2185);
nand U2415 (N_2415,N_1953,N_2333);
nor U2416 (N_2416,N_2236,N_2139);
or U2417 (N_2417,N_2064,N_2308);
xnor U2418 (N_2418,N_2161,N_2380);
nand U2419 (N_2419,N_2128,N_2033);
or U2420 (N_2420,N_1946,N_2325);
or U2421 (N_2421,N_2223,N_2062);
or U2422 (N_2422,N_2012,N_2219);
nor U2423 (N_2423,N_2123,N_2028);
nand U2424 (N_2424,N_2165,N_2211);
xnor U2425 (N_2425,N_1878,N_2205);
nand U2426 (N_2426,N_2051,N_2208);
and U2427 (N_2427,N_2277,N_1894);
xnor U2428 (N_2428,N_2374,N_1974);
xor U2429 (N_2429,N_2387,N_2210);
nand U2430 (N_2430,N_2155,N_2041);
xor U2431 (N_2431,N_2036,N_2390);
or U2432 (N_2432,N_1933,N_1945);
nor U2433 (N_2433,N_2166,N_1854);
nand U2434 (N_2434,N_2086,N_2147);
nand U2435 (N_2435,N_2074,N_2238);
or U2436 (N_2436,N_2010,N_1885);
nand U2437 (N_2437,N_1973,N_2376);
and U2438 (N_2438,N_1817,N_2253);
nand U2439 (N_2439,N_2151,N_2350);
or U2440 (N_2440,N_2202,N_1971);
or U2441 (N_2441,N_1827,N_2259);
and U2442 (N_2442,N_1836,N_2357);
nor U2443 (N_2443,N_1962,N_2173);
nand U2444 (N_2444,N_2326,N_2043);
xor U2445 (N_2445,N_2105,N_2196);
nand U2446 (N_2446,N_2181,N_2224);
nand U2447 (N_2447,N_1872,N_2201);
nand U2448 (N_2448,N_2368,N_1956);
and U2449 (N_2449,N_2172,N_2245);
nor U2450 (N_2450,N_1852,N_2246);
and U2451 (N_2451,N_1858,N_2373);
nor U2452 (N_2452,N_1951,N_1830);
xnor U2453 (N_2453,N_2334,N_2177);
xnor U2454 (N_2454,N_2382,N_2054);
and U2455 (N_2455,N_2003,N_2169);
nor U2456 (N_2456,N_2399,N_1984);
xnor U2457 (N_2457,N_2108,N_2369);
and U2458 (N_2458,N_1926,N_1844);
and U2459 (N_2459,N_2055,N_1823);
xnor U2460 (N_2460,N_1874,N_1967);
nand U2461 (N_2461,N_1922,N_2008);
nand U2462 (N_2462,N_1941,N_1821);
or U2463 (N_2463,N_2204,N_1845);
nand U2464 (N_2464,N_2264,N_2132);
nor U2465 (N_2465,N_2356,N_1949);
nor U2466 (N_2466,N_2363,N_1914);
nor U2467 (N_2467,N_2100,N_2145);
and U2468 (N_2468,N_2347,N_2384);
xor U2469 (N_2469,N_2285,N_2228);
nor U2470 (N_2470,N_2362,N_2154);
or U2471 (N_2471,N_1842,N_2341);
and U2472 (N_2472,N_2372,N_2278);
nand U2473 (N_2473,N_1996,N_1921);
or U2474 (N_2474,N_1832,N_2013);
xor U2475 (N_2475,N_2053,N_2254);
xor U2476 (N_2476,N_2340,N_2011);
and U2477 (N_2477,N_1859,N_2052);
or U2478 (N_2478,N_2093,N_1970);
nand U2479 (N_2479,N_1896,N_2297);
nor U2480 (N_2480,N_2018,N_2294);
xnor U2481 (N_2481,N_2088,N_2396);
or U2482 (N_2482,N_2316,N_2256);
nor U2483 (N_2483,N_2258,N_2042);
and U2484 (N_2484,N_2009,N_1847);
nor U2485 (N_2485,N_1960,N_2150);
or U2486 (N_2486,N_1800,N_2090);
nand U2487 (N_2487,N_2379,N_2038);
and U2488 (N_2488,N_2275,N_1811);
xnor U2489 (N_2489,N_2079,N_2107);
nand U2490 (N_2490,N_1983,N_2284);
or U2491 (N_2491,N_1875,N_2026);
nand U2492 (N_2492,N_2195,N_2135);
nor U2493 (N_2493,N_2104,N_2199);
nor U2494 (N_2494,N_2077,N_2194);
and U2495 (N_2495,N_1828,N_2098);
or U2496 (N_2496,N_2184,N_1904);
xnor U2497 (N_2497,N_1988,N_2206);
and U2498 (N_2498,N_1955,N_2187);
or U2499 (N_2499,N_2260,N_1989);
or U2500 (N_2500,N_1994,N_1911);
nor U2501 (N_2501,N_1870,N_1952);
nand U2502 (N_2502,N_1839,N_2298);
nand U2503 (N_2503,N_2229,N_2320);
and U2504 (N_2504,N_2231,N_2114);
xnor U2505 (N_2505,N_2319,N_2159);
nor U2506 (N_2506,N_1871,N_2014);
nor U2507 (N_2507,N_1934,N_2176);
or U2508 (N_2508,N_2152,N_2276);
nand U2509 (N_2509,N_2371,N_2078);
or U2510 (N_2510,N_1912,N_2241);
or U2511 (N_2511,N_1818,N_1909);
and U2512 (N_2512,N_1923,N_2004);
and U2513 (N_2513,N_2214,N_2359);
nand U2514 (N_2514,N_1978,N_1924);
or U2515 (N_2515,N_2081,N_2191);
and U2516 (N_2516,N_1895,N_1893);
and U2517 (N_2517,N_1980,N_1822);
and U2518 (N_2518,N_2314,N_2303);
nand U2519 (N_2519,N_1925,N_2366);
and U2520 (N_2520,N_2156,N_2186);
xnor U2521 (N_2521,N_1939,N_2133);
and U2522 (N_2522,N_2392,N_1824);
or U2523 (N_2523,N_1860,N_2227);
xor U2524 (N_2524,N_2283,N_2058);
and U2525 (N_2525,N_2335,N_2250);
xor U2526 (N_2526,N_2083,N_2029);
and U2527 (N_2527,N_1927,N_2293);
or U2528 (N_2528,N_1940,N_2321);
nand U2529 (N_2529,N_2160,N_2279);
xor U2530 (N_2530,N_1881,N_2274);
or U2531 (N_2531,N_2257,N_1856);
or U2532 (N_2532,N_2127,N_2346);
xnor U2533 (N_2533,N_2304,N_1918);
nand U2534 (N_2534,N_1812,N_2300);
nand U2535 (N_2535,N_1834,N_1809);
nand U2536 (N_2536,N_2383,N_2237);
nor U2537 (N_2537,N_2398,N_2328);
nor U2538 (N_2538,N_1903,N_2153);
or U2539 (N_2539,N_1950,N_2061);
nand U2540 (N_2540,N_2272,N_2149);
nand U2541 (N_2541,N_2096,N_1961);
or U2542 (N_2542,N_2365,N_2031);
and U2543 (N_2543,N_2358,N_2394);
or U2544 (N_2544,N_2244,N_1906);
nand U2545 (N_2545,N_1917,N_1807);
and U2546 (N_2546,N_2137,N_2289);
nand U2547 (N_2547,N_1966,N_1882);
nand U2548 (N_2548,N_2377,N_2024);
and U2549 (N_2549,N_2097,N_1846);
and U2550 (N_2550,N_2116,N_1877);
nand U2551 (N_2551,N_1819,N_1902);
nand U2552 (N_2552,N_2103,N_2212);
nand U2553 (N_2553,N_2112,N_2126);
nor U2554 (N_2554,N_1937,N_2315);
and U2555 (N_2555,N_2040,N_2305);
nand U2556 (N_2556,N_1943,N_1813);
or U2557 (N_2557,N_1976,N_1897);
or U2558 (N_2558,N_1837,N_2189);
nor U2559 (N_2559,N_2361,N_1814);
or U2560 (N_2560,N_1947,N_2235);
xor U2561 (N_2561,N_1816,N_1972);
and U2562 (N_2562,N_1993,N_1958);
and U2563 (N_2563,N_1954,N_2066);
and U2564 (N_2564,N_2327,N_2020);
or U2565 (N_2565,N_2179,N_1831);
nand U2566 (N_2566,N_1915,N_1805);
nand U2567 (N_2567,N_2175,N_2273);
xnor U2568 (N_2568,N_1803,N_2252);
nor U2569 (N_2569,N_1806,N_2134);
nor U2570 (N_2570,N_2337,N_2095);
and U2571 (N_2571,N_2288,N_2084);
nand U2572 (N_2572,N_2266,N_2209);
nand U2573 (N_2573,N_2332,N_2131);
xor U2574 (N_2574,N_1883,N_2101);
nor U2575 (N_2575,N_2047,N_2158);
xor U2576 (N_2576,N_1930,N_1889);
or U2577 (N_2577,N_2251,N_2023);
nand U2578 (N_2578,N_2296,N_1908);
xnor U2579 (N_2579,N_2270,N_2046);
nand U2580 (N_2580,N_2087,N_2389);
and U2581 (N_2581,N_2342,N_2085);
nor U2582 (N_2582,N_1810,N_2217);
and U2583 (N_2583,N_2234,N_2027);
xor U2584 (N_2584,N_2069,N_2353);
nand U2585 (N_2585,N_2089,N_2068);
xnor U2586 (N_2586,N_2073,N_2375);
and U2587 (N_2587,N_2386,N_1898);
xnor U2588 (N_2588,N_1985,N_2044);
nor U2589 (N_2589,N_2242,N_2249);
nand U2590 (N_2590,N_1957,N_1853);
or U2591 (N_2591,N_1979,N_2050);
or U2592 (N_2592,N_2048,N_2072);
xor U2593 (N_2593,N_1995,N_2306);
and U2594 (N_2594,N_2109,N_1876);
xnor U2595 (N_2595,N_1965,N_1892);
nand U2596 (N_2596,N_1820,N_2351);
nand U2597 (N_2597,N_2203,N_2092);
or U2598 (N_2598,N_1849,N_1944);
xnor U2599 (N_2599,N_2343,N_2002);
or U2600 (N_2600,N_2193,N_1884);
and U2601 (N_2601,N_2349,N_2280);
or U2602 (N_2602,N_2322,N_2338);
xor U2603 (N_2603,N_2129,N_1802);
xnor U2604 (N_2604,N_2324,N_1910);
nor U2605 (N_2605,N_2281,N_2080);
nor U2606 (N_2606,N_2309,N_1920);
or U2607 (N_2607,N_1907,N_2397);
or U2608 (N_2608,N_2265,N_1913);
and U2609 (N_2609,N_2282,N_1931);
nor U2610 (N_2610,N_2213,N_2142);
nor U2611 (N_2611,N_2295,N_2140);
nand U2612 (N_2612,N_2071,N_2037);
and U2613 (N_2613,N_2345,N_2113);
nor U2614 (N_2614,N_2312,N_1887);
and U2615 (N_2615,N_2121,N_2395);
xor U2616 (N_2616,N_2000,N_2001);
and U2617 (N_2617,N_2174,N_2025);
or U2618 (N_2618,N_1835,N_1850);
and U2619 (N_2619,N_2130,N_1929);
and U2620 (N_2620,N_2367,N_2122);
and U2621 (N_2621,N_1900,N_2336);
and U2622 (N_2622,N_2070,N_2118);
and U2623 (N_2623,N_1886,N_2364);
nor U2624 (N_2624,N_2302,N_1891);
nor U2625 (N_2625,N_1905,N_2125);
nand U2626 (N_2626,N_2019,N_2291);
or U2627 (N_2627,N_2076,N_1841);
xnor U2628 (N_2628,N_1948,N_1997);
or U2629 (N_2629,N_2124,N_2290);
nand U2630 (N_2630,N_2163,N_2310);
or U2631 (N_2631,N_2286,N_2007);
nor U2632 (N_2632,N_2063,N_2360);
xnor U2633 (N_2633,N_2091,N_2057);
xnor U2634 (N_2634,N_1977,N_1928);
and U2635 (N_2635,N_1829,N_2094);
nor U2636 (N_2636,N_2015,N_1938);
and U2637 (N_2637,N_1936,N_2311);
nand U2638 (N_2638,N_1840,N_2331);
or U2639 (N_2639,N_2263,N_2207);
nand U2640 (N_2640,N_1857,N_2006);
nor U2641 (N_2641,N_1868,N_2198);
or U2642 (N_2642,N_1826,N_2344);
nor U2643 (N_2643,N_1968,N_2188);
and U2644 (N_2644,N_2388,N_1986);
xor U2645 (N_2645,N_2039,N_2110);
and U2646 (N_2646,N_2292,N_1851);
nand U2647 (N_2647,N_2370,N_1999);
or U2648 (N_2648,N_2182,N_1942);
nor U2649 (N_2649,N_2164,N_1866);
or U2650 (N_2650,N_1815,N_2067);
and U2651 (N_2651,N_1969,N_1865);
nor U2652 (N_2652,N_1867,N_2355);
nand U2653 (N_2653,N_2141,N_2099);
or U2654 (N_2654,N_1838,N_2299);
and U2655 (N_2655,N_1804,N_2301);
and U2656 (N_2656,N_2157,N_1992);
nand U2657 (N_2657,N_2215,N_1890);
nand U2658 (N_2658,N_2111,N_1932);
and U2659 (N_2659,N_2385,N_2115);
nor U2660 (N_2660,N_1864,N_2247);
or U2661 (N_2661,N_1991,N_2065);
nand U2662 (N_2662,N_2248,N_2200);
and U2663 (N_2663,N_2268,N_2287);
nand U2664 (N_2664,N_2262,N_2216);
xor U2665 (N_2665,N_2222,N_2221);
xnor U2666 (N_2666,N_2146,N_1873);
xnor U2667 (N_2667,N_2138,N_2381);
nor U2668 (N_2668,N_2117,N_2075);
nor U2669 (N_2669,N_1801,N_1916);
nand U2670 (N_2670,N_2318,N_2317);
and U2671 (N_2671,N_1919,N_2016);
and U2672 (N_2672,N_2267,N_2329);
xnor U2673 (N_2673,N_2021,N_1963);
nor U2674 (N_2674,N_2393,N_2106);
xor U2675 (N_2675,N_2323,N_1825);
and U2676 (N_2676,N_1855,N_2119);
nor U2677 (N_2677,N_2233,N_2220);
nor U2678 (N_2678,N_2190,N_1901);
and U2679 (N_2679,N_2352,N_2378);
or U2680 (N_2680,N_2136,N_2060);
nor U2681 (N_2681,N_2120,N_1987);
nor U2682 (N_2682,N_2167,N_2313);
or U2683 (N_2683,N_2035,N_2034);
and U2684 (N_2684,N_2144,N_1981);
and U2685 (N_2685,N_2330,N_2271);
nor U2686 (N_2686,N_2049,N_2005);
and U2687 (N_2687,N_1990,N_1808);
nor U2688 (N_2688,N_2307,N_2339);
nand U2689 (N_2689,N_2056,N_2171);
xor U2690 (N_2690,N_2168,N_2045);
and U2691 (N_2691,N_2192,N_1862);
and U2692 (N_2692,N_1982,N_1964);
and U2693 (N_2693,N_1863,N_2102);
nand U2694 (N_2694,N_1959,N_2239);
nor U2695 (N_2695,N_1833,N_2148);
or U2696 (N_2696,N_1880,N_1848);
and U2697 (N_2697,N_2030,N_2017);
and U2698 (N_2698,N_1879,N_2180);
nor U2699 (N_2699,N_1935,N_1998);
xnor U2700 (N_2700,N_2275,N_2133);
xnor U2701 (N_2701,N_2324,N_2020);
nor U2702 (N_2702,N_2054,N_2207);
xnor U2703 (N_2703,N_2319,N_1815);
or U2704 (N_2704,N_1854,N_1863);
nand U2705 (N_2705,N_2331,N_1856);
and U2706 (N_2706,N_1891,N_2090);
xnor U2707 (N_2707,N_2126,N_2087);
nand U2708 (N_2708,N_2287,N_2011);
nor U2709 (N_2709,N_1928,N_1979);
nor U2710 (N_2710,N_2248,N_2194);
or U2711 (N_2711,N_2341,N_2133);
nand U2712 (N_2712,N_2294,N_1998);
or U2713 (N_2713,N_2362,N_2088);
nor U2714 (N_2714,N_1937,N_1843);
nand U2715 (N_2715,N_2296,N_1909);
nand U2716 (N_2716,N_2099,N_2278);
xnor U2717 (N_2717,N_1883,N_2335);
and U2718 (N_2718,N_2080,N_1804);
or U2719 (N_2719,N_2257,N_1836);
and U2720 (N_2720,N_2012,N_2204);
and U2721 (N_2721,N_2145,N_1886);
nor U2722 (N_2722,N_2049,N_2073);
xnor U2723 (N_2723,N_2174,N_1942);
and U2724 (N_2724,N_2266,N_2231);
or U2725 (N_2725,N_2130,N_2384);
nor U2726 (N_2726,N_2360,N_2284);
nor U2727 (N_2727,N_1825,N_1984);
nor U2728 (N_2728,N_2117,N_2103);
or U2729 (N_2729,N_1973,N_1929);
and U2730 (N_2730,N_2072,N_2039);
or U2731 (N_2731,N_2005,N_1936);
xor U2732 (N_2732,N_2295,N_2044);
and U2733 (N_2733,N_2326,N_1922);
xor U2734 (N_2734,N_2348,N_2201);
nor U2735 (N_2735,N_1868,N_1860);
nand U2736 (N_2736,N_2096,N_1952);
or U2737 (N_2737,N_2169,N_1826);
nand U2738 (N_2738,N_2186,N_2180);
nand U2739 (N_2739,N_1808,N_2009);
xor U2740 (N_2740,N_1805,N_2288);
nor U2741 (N_2741,N_2264,N_2108);
nor U2742 (N_2742,N_2184,N_2017);
and U2743 (N_2743,N_2095,N_2117);
or U2744 (N_2744,N_2062,N_2357);
and U2745 (N_2745,N_2324,N_1940);
or U2746 (N_2746,N_2080,N_2116);
or U2747 (N_2747,N_1852,N_1994);
nor U2748 (N_2748,N_1940,N_2029);
nor U2749 (N_2749,N_2332,N_2366);
and U2750 (N_2750,N_1986,N_2090);
nand U2751 (N_2751,N_2324,N_1880);
nor U2752 (N_2752,N_2375,N_1835);
nor U2753 (N_2753,N_1861,N_2277);
xnor U2754 (N_2754,N_2323,N_1943);
or U2755 (N_2755,N_1944,N_2254);
or U2756 (N_2756,N_2194,N_2040);
or U2757 (N_2757,N_1899,N_1829);
nor U2758 (N_2758,N_2373,N_1828);
or U2759 (N_2759,N_1911,N_2253);
nor U2760 (N_2760,N_2022,N_1843);
xor U2761 (N_2761,N_1969,N_2058);
nand U2762 (N_2762,N_1813,N_2232);
or U2763 (N_2763,N_1896,N_2291);
nor U2764 (N_2764,N_2381,N_2112);
and U2765 (N_2765,N_2351,N_1817);
nor U2766 (N_2766,N_1867,N_2313);
nor U2767 (N_2767,N_1944,N_2288);
or U2768 (N_2768,N_2227,N_2165);
xor U2769 (N_2769,N_2194,N_1832);
nor U2770 (N_2770,N_2117,N_2233);
xor U2771 (N_2771,N_2330,N_1850);
or U2772 (N_2772,N_2189,N_2111);
xnor U2773 (N_2773,N_2184,N_2140);
nor U2774 (N_2774,N_1917,N_1808);
nor U2775 (N_2775,N_1977,N_1893);
or U2776 (N_2776,N_2178,N_2308);
nand U2777 (N_2777,N_1841,N_2127);
and U2778 (N_2778,N_1855,N_1997);
and U2779 (N_2779,N_2168,N_2111);
nor U2780 (N_2780,N_1841,N_1933);
or U2781 (N_2781,N_2228,N_2185);
nand U2782 (N_2782,N_2106,N_2182);
xnor U2783 (N_2783,N_2179,N_2396);
or U2784 (N_2784,N_2362,N_1805);
or U2785 (N_2785,N_1960,N_2385);
and U2786 (N_2786,N_2106,N_2056);
nor U2787 (N_2787,N_2070,N_2030);
or U2788 (N_2788,N_2213,N_2043);
and U2789 (N_2789,N_2140,N_2045);
or U2790 (N_2790,N_1944,N_2299);
and U2791 (N_2791,N_2139,N_2331);
nand U2792 (N_2792,N_2203,N_2053);
and U2793 (N_2793,N_2245,N_2185);
xnor U2794 (N_2794,N_2108,N_2136);
or U2795 (N_2795,N_2267,N_2025);
xnor U2796 (N_2796,N_2252,N_2141);
nor U2797 (N_2797,N_1959,N_2133);
xor U2798 (N_2798,N_2353,N_1929);
xnor U2799 (N_2799,N_2119,N_2248);
or U2800 (N_2800,N_2046,N_1916);
xnor U2801 (N_2801,N_1937,N_2276);
xor U2802 (N_2802,N_2302,N_1927);
nand U2803 (N_2803,N_2186,N_1912);
nor U2804 (N_2804,N_2335,N_1937);
nor U2805 (N_2805,N_2271,N_2301);
nor U2806 (N_2806,N_2309,N_1982);
nor U2807 (N_2807,N_2213,N_2288);
nand U2808 (N_2808,N_2184,N_1800);
nand U2809 (N_2809,N_2222,N_2297);
and U2810 (N_2810,N_1808,N_2032);
and U2811 (N_2811,N_2270,N_2160);
or U2812 (N_2812,N_1967,N_2125);
and U2813 (N_2813,N_2184,N_1848);
xor U2814 (N_2814,N_1990,N_1927);
nor U2815 (N_2815,N_2134,N_1970);
nor U2816 (N_2816,N_2012,N_2300);
and U2817 (N_2817,N_1947,N_2325);
nand U2818 (N_2818,N_2278,N_2228);
nand U2819 (N_2819,N_2033,N_2084);
and U2820 (N_2820,N_1913,N_2077);
nor U2821 (N_2821,N_2182,N_2153);
xnor U2822 (N_2822,N_2127,N_2123);
or U2823 (N_2823,N_1879,N_1963);
and U2824 (N_2824,N_1896,N_2220);
nor U2825 (N_2825,N_1931,N_1911);
nand U2826 (N_2826,N_2372,N_1824);
nor U2827 (N_2827,N_1913,N_1933);
and U2828 (N_2828,N_1919,N_2119);
nor U2829 (N_2829,N_2096,N_1927);
nand U2830 (N_2830,N_2243,N_2039);
and U2831 (N_2831,N_1889,N_1853);
nor U2832 (N_2832,N_2286,N_2262);
nor U2833 (N_2833,N_2322,N_2381);
nor U2834 (N_2834,N_1917,N_1913);
or U2835 (N_2835,N_1875,N_2007);
nor U2836 (N_2836,N_2040,N_1973);
and U2837 (N_2837,N_1952,N_2123);
xnor U2838 (N_2838,N_2329,N_2061);
nand U2839 (N_2839,N_2319,N_1921);
xnor U2840 (N_2840,N_2225,N_1988);
xor U2841 (N_2841,N_2175,N_2185);
xnor U2842 (N_2842,N_1894,N_2319);
nand U2843 (N_2843,N_2308,N_1816);
nor U2844 (N_2844,N_2389,N_1988);
and U2845 (N_2845,N_2147,N_2196);
nand U2846 (N_2846,N_2207,N_2142);
xnor U2847 (N_2847,N_1907,N_2125);
nand U2848 (N_2848,N_2036,N_2072);
and U2849 (N_2849,N_2053,N_2047);
or U2850 (N_2850,N_2195,N_1869);
or U2851 (N_2851,N_2240,N_2213);
or U2852 (N_2852,N_1867,N_2230);
and U2853 (N_2853,N_2035,N_2003);
or U2854 (N_2854,N_2153,N_2340);
nand U2855 (N_2855,N_1891,N_1903);
nor U2856 (N_2856,N_2184,N_2059);
or U2857 (N_2857,N_2392,N_1865);
or U2858 (N_2858,N_2203,N_2145);
xor U2859 (N_2859,N_2091,N_2196);
or U2860 (N_2860,N_1824,N_2386);
or U2861 (N_2861,N_2231,N_2138);
or U2862 (N_2862,N_2306,N_2033);
nand U2863 (N_2863,N_2297,N_2148);
nor U2864 (N_2864,N_2185,N_1928);
and U2865 (N_2865,N_1818,N_1837);
xnor U2866 (N_2866,N_1952,N_1886);
nand U2867 (N_2867,N_2311,N_1939);
nand U2868 (N_2868,N_2053,N_1907);
nand U2869 (N_2869,N_2146,N_2303);
xor U2870 (N_2870,N_1817,N_2051);
xor U2871 (N_2871,N_2378,N_1904);
or U2872 (N_2872,N_1915,N_2320);
nand U2873 (N_2873,N_1945,N_2146);
nor U2874 (N_2874,N_2027,N_2102);
nor U2875 (N_2875,N_2274,N_2367);
nor U2876 (N_2876,N_1992,N_2237);
nand U2877 (N_2877,N_2101,N_1800);
and U2878 (N_2878,N_1949,N_2359);
or U2879 (N_2879,N_2087,N_2203);
or U2880 (N_2880,N_1861,N_2073);
or U2881 (N_2881,N_2114,N_2096);
nand U2882 (N_2882,N_2247,N_2281);
or U2883 (N_2883,N_2056,N_2100);
nand U2884 (N_2884,N_2097,N_2146);
or U2885 (N_2885,N_2361,N_2268);
or U2886 (N_2886,N_1868,N_1803);
or U2887 (N_2887,N_1935,N_1822);
xor U2888 (N_2888,N_2118,N_2105);
nand U2889 (N_2889,N_2088,N_2036);
and U2890 (N_2890,N_2012,N_2120);
xnor U2891 (N_2891,N_2204,N_2179);
and U2892 (N_2892,N_2225,N_1876);
and U2893 (N_2893,N_2087,N_2383);
nor U2894 (N_2894,N_2339,N_2164);
nand U2895 (N_2895,N_2253,N_2318);
or U2896 (N_2896,N_2294,N_2168);
nor U2897 (N_2897,N_2213,N_1909);
nand U2898 (N_2898,N_2080,N_2347);
and U2899 (N_2899,N_2362,N_2093);
nand U2900 (N_2900,N_1966,N_2129);
nand U2901 (N_2901,N_2249,N_1928);
xor U2902 (N_2902,N_2091,N_1991);
nand U2903 (N_2903,N_2154,N_2344);
or U2904 (N_2904,N_1872,N_1970);
and U2905 (N_2905,N_2325,N_2218);
nor U2906 (N_2906,N_2213,N_1992);
and U2907 (N_2907,N_2259,N_1893);
xnor U2908 (N_2908,N_1920,N_2293);
nand U2909 (N_2909,N_2009,N_2126);
nand U2910 (N_2910,N_2355,N_2080);
nand U2911 (N_2911,N_2230,N_2366);
nand U2912 (N_2912,N_1953,N_2087);
or U2913 (N_2913,N_2023,N_1968);
nor U2914 (N_2914,N_2120,N_2124);
xor U2915 (N_2915,N_1985,N_2133);
nand U2916 (N_2916,N_2234,N_1938);
xor U2917 (N_2917,N_2353,N_2213);
xnor U2918 (N_2918,N_2171,N_2146);
nand U2919 (N_2919,N_1984,N_1884);
xnor U2920 (N_2920,N_1839,N_1810);
or U2921 (N_2921,N_1856,N_2294);
xnor U2922 (N_2922,N_2033,N_2335);
xnor U2923 (N_2923,N_2325,N_2353);
or U2924 (N_2924,N_2064,N_1968);
or U2925 (N_2925,N_2281,N_2290);
or U2926 (N_2926,N_1998,N_1801);
nand U2927 (N_2927,N_2368,N_1994);
and U2928 (N_2928,N_2209,N_2156);
or U2929 (N_2929,N_1861,N_2247);
nand U2930 (N_2930,N_2231,N_2179);
and U2931 (N_2931,N_2096,N_1843);
xor U2932 (N_2932,N_2329,N_2360);
or U2933 (N_2933,N_1921,N_2363);
xor U2934 (N_2934,N_2245,N_2101);
nand U2935 (N_2935,N_2189,N_2168);
and U2936 (N_2936,N_2181,N_2032);
nor U2937 (N_2937,N_1930,N_1960);
nor U2938 (N_2938,N_2368,N_2268);
and U2939 (N_2939,N_1920,N_2270);
xnor U2940 (N_2940,N_2350,N_2076);
nor U2941 (N_2941,N_2388,N_1978);
and U2942 (N_2942,N_2050,N_1884);
nor U2943 (N_2943,N_2164,N_2344);
xor U2944 (N_2944,N_1941,N_2225);
and U2945 (N_2945,N_1858,N_2303);
xnor U2946 (N_2946,N_2303,N_2277);
nor U2947 (N_2947,N_1978,N_2073);
or U2948 (N_2948,N_2090,N_1879);
and U2949 (N_2949,N_1865,N_2385);
nand U2950 (N_2950,N_1840,N_2108);
nor U2951 (N_2951,N_1868,N_2162);
xnor U2952 (N_2952,N_1959,N_2372);
nand U2953 (N_2953,N_2154,N_2071);
or U2954 (N_2954,N_2093,N_2261);
or U2955 (N_2955,N_1848,N_1924);
nor U2956 (N_2956,N_2062,N_1955);
xor U2957 (N_2957,N_2275,N_1800);
or U2958 (N_2958,N_2018,N_2308);
nand U2959 (N_2959,N_2396,N_2287);
and U2960 (N_2960,N_1915,N_1961);
nand U2961 (N_2961,N_1864,N_1936);
or U2962 (N_2962,N_2165,N_2007);
nor U2963 (N_2963,N_2272,N_1876);
and U2964 (N_2964,N_1911,N_2044);
and U2965 (N_2965,N_1902,N_2241);
nor U2966 (N_2966,N_1988,N_1880);
nor U2967 (N_2967,N_1965,N_2370);
nor U2968 (N_2968,N_2363,N_1976);
xnor U2969 (N_2969,N_1963,N_2048);
nand U2970 (N_2970,N_2352,N_2290);
nor U2971 (N_2971,N_2171,N_1998);
or U2972 (N_2972,N_2153,N_2033);
nor U2973 (N_2973,N_2080,N_2177);
or U2974 (N_2974,N_2036,N_1971);
or U2975 (N_2975,N_2188,N_2323);
and U2976 (N_2976,N_2137,N_1841);
nor U2977 (N_2977,N_1800,N_2140);
or U2978 (N_2978,N_2013,N_2108);
nand U2979 (N_2979,N_2201,N_2114);
and U2980 (N_2980,N_1958,N_2103);
nand U2981 (N_2981,N_2070,N_2344);
nand U2982 (N_2982,N_2066,N_1976);
or U2983 (N_2983,N_2042,N_2398);
nand U2984 (N_2984,N_2183,N_1851);
and U2985 (N_2985,N_1920,N_2130);
nand U2986 (N_2986,N_1979,N_1873);
nor U2987 (N_2987,N_2373,N_2344);
xor U2988 (N_2988,N_1957,N_2057);
or U2989 (N_2989,N_2314,N_2304);
or U2990 (N_2990,N_1942,N_1810);
and U2991 (N_2991,N_1881,N_2221);
nand U2992 (N_2992,N_2174,N_2367);
or U2993 (N_2993,N_2077,N_2086);
or U2994 (N_2994,N_1961,N_2056);
xnor U2995 (N_2995,N_2276,N_2194);
or U2996 (N_2996,N_1928,N_1832);
xnor U2997 (N_2997,N_2320,N_1918);
nor U2998 (N_2998,N_2190,N_2208);
and U2999 (N_2999,N_2216,N_2286);
or U3000 (N_3000,N_2654,N_2524);
xnor U3001 (N_3001,N_2769,N_2479);
nand U3002 (N_3002,N_2408,N_2993);
nor U3003 (N_3003,N_2675,N_2625);
and U3004 (N_3004,N_2568,N_2768);
or U3005 (N_3005,N_2532,N_2452);
and U3006 (N_3006,N_2771,N_2717);
or U3007 (N_3007,N_2629,N_2642);
xnor U3008 (N_3008,N_2487,N_2605);
nor U3009 (N_3009,N_2517,N_2521);
nor U3010 (N_3010,N_2480,N_2696);
and U3011 (N_3011,N_2502,N_2732);
nand U3012 (N_3012,N_2709,N_2857);
or U3013 (N_3013,N_2514,N_2926);
xnor U3014 (N_3014,N_2948,N_2982);
nand U3015 (N_3015,N_2655,N_2825);
xor U3016 (N_3016,N_2423,N_2535);
and U3017 (N_3017,N_2402,N_2976);
or U3018 (N_3018,N_2927,N_2753);
nand U3019 (N_3019,N_2551,N_2988);
and U3020 (N_3020,N_2538,N_2458);
xor U3021 (N_3021,N_2766,N_2958);
and U3022 (N_3022,N_2876,N_2519);
nand U3023 (N_3023,N_2561,N_2497);
and U3024 (N_3024,N_2481,N_2965);
nor U3025 (N_3025,N_2541,N_2752);
nand U3026 (N_3026,N_2566,N_2811);
or U3027 (N_3027,N_2909,N_2758);
and U3028 (N_3028,N_2503,N_2903);
xnor U3029 (N_3029,N_2516,N_2567);
or U3030 (N_3030,N_2898,N_2492);
xnor U3031 (N_3031,N_2688,N_2546);
nor U3032 (N_3032,N_2936,N_2735);
or U3033 (N_3033,N_2460,N_2456);
and U3034 (N_3034,N_2728,N_2729);
nand U3035 (N_3035,N_2457,N_2777);
xnor U3036 (N_3036,N_2809,N_2829);
nor U3037 (N_3037,N_2540,N_2499);
nand U3038 (N_3038,N_2704,N_2400);
nand U3039 (N_3039,N_2639,N_2646);
or U3040 (N_3040,N_2987,N_2484);
xnor U3041 (N_3041,N_2755,N_2881);
nand U3042 (N_3042,N_2421,N_2464);
nor U3043 (N_3043,N_2974,N_2872);
nor U3044 (N_3044,N_2870,N_2565);
nor U3045 (N_3045,N_2527,N_2469);
nor U3046 (N_3046,N_2840,N_2944);
xor U3047 (N_3047,N_2865,N_2961);
nand U3048 (N_3048,N_2427,N_2859);
or U3049 (N_3049,N_2520,N_2947);
xnor U3050 (N_3050,N_2433,N_2883);
xnor U3051 (N_3051,N_2939,N_2558);
xnor U3052 (N_3052,N_2589,N_2784);
or U3053 (N_3053,N_2813,N_2573);
nand U3054 (N_3054,N_2760,N_2489);
xnor U3055 (N_3055,N_2679,N_2610);
nand U3056 (N_3056,N_2957,N_2648);
nand U3057 (N_3057,N_2761,N_2619);
or U3058 (N_3058,N_2448,N_2543);
and U3059 (N_3059,N_2860,N_2962);
xnor U3060 (N_3060,N_2575,N_2673);
and U3061 (N_3061,N_2842,N_2801);
xnor U3062 (N_3062,N_2830,N_2416);
xnor U3063 (N_3063,N_2434,N_2645);
nand U3064 (N_3064,N_2737,N_2530);
nand U3065 (N_3065,N_2618,N_2733);
or U3066 (N_3066,N_2963,N_2496);
nand U3067 (N_3067,N_2879,N_2498);
xor U3068 (N_3068,N_2432,N_2415);
and U3069 (N_3069,N_2592,N_2967);
and U3070 (N_3070,N_2966,N_2627);
xor U3071 (N_3071,N_2506,N_2716);
nor U3072 (N_3072,N_2607,N_2756);
xnor U3073 (N_3073,N_2807,N_2689);
nor U3074 (N_3074,N_2485,N_2582);
xnor U3075 (N_3075,N_2938,N_2658);
and U3076 (N_3076,N_2933,N_2803);
nor U3077 (N_3077,N_2711,N_2653);
nand U3078 (N_3078,N_2604,N_2461);
xor U3079 (N_3079,N_2742,N_2429);
nand U3080 (N_3080,N_2741,N_2690);
or U3081 (N_3081,N_2624,N_2955);
xnor U3082 (N_3082,N_2925,N_2996);
nor U3083 (N_3083,N_2907,N_2725);
nor U3084 (N_3084,N_2921,N_2792);
xnor U3085 (N_3085,N_2867,N_2826);
nand U3086 (N_3086,N_2483,N_2700);
xor U3087 (N_3087,N_2477,N_2796);
xor U3088 (N_3088,N_2832,N_2536);
and U3089 (N_3089,N_2425,N_2914);
and U3090 (N_3090,N_2413,N_2467);
and U3091 (N_3091,N_2978,N_2552);
xor U3092 (N_3092,N_2578,N_2971);
and U3093 (N_3093,N_2763,N_2950);
or U3094 (N_3094,N_2633,N_2476);
and U3095 (N_3095,N_2710,N_2775);
and U3096 (N_3096,N_2686,N_2613);
nand U3097 (N_3097,N_2439,N_2699);
nand U3098 (N_3098,N_2637,N_2869);
xor U3099 (N_3099,N_2892,N_2919);
or U3100 (N_3100,N_2684,N_2804);
nor U3101 (N_3101,N_2972,N_2577);
and U3102 (N_3102,N_2923,N_2856);
xnor U3103 (N_3103,N_2652,N_2937);
nor U3104 (N_3104,N_2705,N_2436);
nor U3105 (N_3105,N_2672,N_2749);
and U3106 (N_3106,N_2922,N_2435);
or U3107 (N_3107,N_2443,N_2897);
nand U3108 (N_3108,N_2726,N_2960);
or U3109 (N_3109,N_2471,N_2409);
nor U3110 (N_3110,N_2977,N_2776);
nor U3111 (N_3111,N_2975,N_2598);
xor U3112 (N_3112,N_2647,N_2664);
or U3113 (N_3113,N_2419,N_2587);
xor U3114 (N_3114,N_2547,N_2523);
nor U3115 (N_3115,N_2422,N_2992);
xnor U3116 (N_3116,N_2871,N_2841);
nand U3117 (N_3117,N_2848,N_2537);
xor U3118 (N_3118,N_2703,N_2828);
xor U3119 (N_3119,N_2849,N_2852);
or U3120 (N_3120,N_2437,N_2990);
nor U3121 (N_3121,N_2544,N_2600);
or U3122 (N_3122,N_2449,N_2632);
or U3123 (N_3123,N_2671,N_2494);
xor U3124 (N_3124,N_2823,N_2681);
xnor U3125 (N_3125,N_2946,N_2884);
and U3126 (N_3126,N_2863,N_2640);
nor U3127 (N_3127,N_2727,N_2724);
and U3128 (N_3128,N_2949,N_2586);
and U3129 (N_3129,N_2738,N_2593);
xnor U3130 (N_3130,N_2656,N_2781);
or U3131 (N_3131,N_2953,N_2790);
nor U3132 (N_3132,N_2821,N_2942);
nand U3133 (N_3133,N_2431,N_2877);
nor U3134 (N_3134,N_2626,N_2956);
and U3135 (N_3135,N_2968,N_2782);
xnor U3136 (N_3136,N_2820,N_2526);
or U3137 (N_3137,N_2579,N_2845);
nand U3138 (N_3138,N_2912,N_2562);
or U3139 (N_3139,N_2698,N_2542);
nor U3140 (N_3140,N_2878,N_2574);
and U3141 (N_3141,N_2644,N_2445);
xor U3142 (N_3142,N_2602,N_2899);
nand U3143 (N_3143,N_2814,N_2585);
or U3144 (N_3144,N_2864,N_2844);
xnor U3145 (N_3145,N_2571,N_2563);
and U3146 (N_3146,N_2723,N_2455);
xor U3147 (N_3147,N_2930,N_2470);
and U3148 (N_3148,N_2695,N_2910);
and U3149 (N_3149,N_2734,N_2858);
nor U3150 (N_3150,N_2887,N_2838);
or U3151 (N_3151,N_2720,N_2918);
nor U3152 (N_3152,N_2472,N_2465);
or U3153 (N_3153,N_2611,N_2559);
or U3154 (N_3154,N_2708,N_2615);
and U3155 (N_3155,N_2410,N_2691);
nand U3156 (N_3156,N_2687,N_2442);
or U3157 (N_3157,N_2683,N_2808);
nand U3158 (N_3158,N_2905,N_2951);
nand U3159 (N_3159,N_2660,N_2855);
nand U3160 (N_3160,N_2407,N_2555);
xnor U3161 (N_3161,N_2793,N_2983);
xnor U3162 (N_3162,N_2474,N_2504);
xnor U3163 (N_3163,N_2875,N_2995);
xnor U3164 (N_3164,N_2508,N_2650);
nand U3165 (N_3165,N_2453,N_2534);
nor U3166 (N_3166,N_2981,N_2603);
nand U3167 (N_3167,N_2843,N_2818);
and U3168 (N_3168,N_2420,N_2482);
nand U3169 (N_3169,N_2446,N_2634);
or U3170 (N_3170,N_2989,N_2780);
nor U3171 (N_3171,N_2641,N_2659);
xnor U3172 (N_3172,N_2682,N_2512);
xor U3173 (N_3173,N_2430,N_2952);
and U3174 (N_3174,N_2454,N_2412);
and U3175 (N_3175,N_2731,N_2623);
nand U3176 (N_3176,N_2511,N_2835);
nand U3177 (N_3177,N_2815,N_2557);
nand U3178 (N_3178,N_2583,N_2740);
xnor U3179 (N_3179,N_2513,N_2928);
nor U3180 (N_3180,N_2817,N_2490);
and U3181 (N_3181,N_2450,N_2553);
nand U3182 (N_3182,N_2822,N_2697);
and U3183 (N_3183,N_2556,N_2772);
xnor U3184 (N_3184,N_2588,N_2486);
or U3185 (N_3185,N_2406,N_2500);
or U3186 (N_3186,N_2570,N_2764);
nand U3187 (N_3187,N_2836,N_2522);
xor U3188 (N_3188,N_2676,N_2888);
xnor U3189 (N_3189,N_2649,N_2596);
or U3190 (N_3190,N_2934,N_2806);
nor U3191 (N_3191,N_2874,N_2904);
xor U3192 (N_3192,N_2440,N_2787);
or U3193 (N_3193,N_2631,N_2783);
and U3194 (N_3194,N_2564,N_2959);
and U3195 (N_3195,N_2518,N_2560);
or U3196 (N_3196,N_2451,N_2964);
nor U3197 (N_3197,N_2591,N_2721);
and U3198 (N_3198,N_2621,N_2663);
nand U3199 (N_3199,N_2831,N_2861);
xor U3200 (N_3200,N_2706,N_2507);
and U3201 (N_3201,N_2417,N_2873);
xor U3202 (N_3202,N_2794,N_2473);
nor U3203 (N_3203,N_2447,N_2707);
nor U3204 (N_3204,N_2911,N_2750);
nor U3205 (N_3205,N_2539,N_2935);
and U3206 (N_3206,N_2765,N_2924);
nand U3207 (N_3207,N_2594,N_2515);
nand U3208 (N_3208,N_2712,N_2463);
or U3209 (N_3209,N_2620,N_2833);
xnor U3210 (N_3210,N_2894,N_2901);
nor U3211 (N_3211,N_2751,N_2674);
nand U3212 (N_3212,N_2979,N_2661);
or U3213 (N_3213,N_2779,N_2880);
xor U3214 (N_3214,N_2920,N_2590);
nand U3215 (N_3215,N_2932,N_2773);
xnor U3216 (N_3216,N_2501,N_2789);
xor U3217 (N_3217,N_2612,N_2510);
nand U3218 (N_3218,N_2748,N_2630);
nand U3219 (N_3219,N_2668,N_2509);
nand U3220 (N_3220,N_2529,N_2985);
nand U3221 (N_3221,N_2597,N_2713);
xor U3222 (N_3222,N_2908,N_2576);
or U3223 (N_3223,N_2569,N_2931);
xnor U3224 (N_3224,N_2945,N_2418);
nor U3225 (N_3225,N_2669,N_2719);
nor U3226 (N_3226,N_2846,N_2785);
xor U3227 (N_3227,N_2882,N_2614);
nand U3228 (N_3228,N_2984,N_2616);
and U3229 (N_3229,N_2827,N_2493);
nor U3230 (N_3230,N_2778,N_2617);
nand U3231 (N_3231,N_2940,N_2545);
xnor U3232 (N_3232,N_2913,N_2678);
nor U3233 (N_3233,N_2886,N_2628);
xor U3234 (N_3234,N_2608,N_2837);
nand U3235 (N_3235,N_2662,N_2969);
and U3236 (N_3236,N_2403,N_2770);
and U3237 (N_3237,N_2730,N_2638);
and U3238 (N_3238,N_2525,N_2572);
nor U3239 (N_3239,N_2736,N_2424);
nor U3240 (N_3240,N_2428,N_2609);
nor U3241 (N_3241,N_2991,N_2666);
or U3242 (N_3242,N_2797,N_2595);
nand U3243 (N_3243,N_2606,N_2999);
nor U3244 (N_3244,N_2757,N_2798);
nand U3245 (N_3245,N_2715,N_2805);
or U3246 (N_3246,N_2890,N_2810);
or U3247 (N_3247,N_2441,N_2722);
nand U3248 (N_3248,N_2462,N_2906);
nor U3249 (N_3249,N_2466,N_2692);
and U3250 (N_3250,N_2970,N_2657);
or U3251 (N_3251,N_2444,N_2895);
or U3252 (N_3252,N_2550,N_2788);
nand U3253 (N_3253,N_2739,N_2665);
xnor U3254 (N_3254,N_2973,N_2531);
and U3255 (N_3255,N_2854,N_2404);
or U3256 (N_3256,N_2548,N_2701);
or U3257 (N_3257,N_2554,N_2819);
nand U3258 (N_3258,N_2405,N_2980);
and U3259 (N_3259,N_2411,N_2853);
or U3260 (N_3260,N_2685,N_2702);
nor U3261 (N_3261,N_2601,N_2714);
or U3262 (N_3262,N_2847,N_2816);
nor U3263 (N_3263,N_2986,N_2426);
xnor U3264 (N_3264,N_2488,N_2834);
xnor U3265 (N_3265,N_2917,N_2468);
xnor U3266 (N_3266,N_2533,N_2718);
and U3267 (N_3267,N_2998,N_2693);
nand U3268 (N_3268,N_2599,N_2580);
xnor U3269 (N_3269,N_2850,N_2795);
and U3270 (N_3270,N_2954,N_2900);
or U3271 (N_3271,N_2800,N_2851);
xnor U3272 (N_3272,N_2581,N_2812);
nand U3273 (N_3273,N_2745,N_2994);
nor U3274 (N_3274,N_2746,N_2896);
nand U3275 (N_3275,N_2743,N_2862);
or U3276 (N_3276,N_2893,N_2791);
nor U3277 (N_3277,N_2786,N_2902);
or U3278 (N_3278,N_2495,N_2929);
nand U3279 (N_3279,N_2802,N_2401);
and U3280 (N_3280,N_2478,N_2635);
nand U3281 (N_3281,N_2889,N_2414);
nand U3282 (N_3282,N_2584,N_2680);
or U3283 (N_3283,N_2677,N_2866);
xor U3284 (N_3284,N_2438,N_2505);
nand U3285 (N_3285,N_2549,N_2767);
xnor U3286 (N_3286,N_2868,N_2636);
and U3287 (N_3287,N_2799,N_2747);
or U3288 (N_3288,N_2651,N_2622);
or U3289 (N_3289,N_2824,N_2916);
and U3290 (N_3290,N_2744,N_2459);
and U3291 (N_3291,N_2754,N_2839);
nor U3292 (N_3292,N_2891,N_2774);
nand U3293 (N_3293,N_2528,N_2762);
xnor U3294 (N_3294,N_2667,N_2694);
nand U3295 (N_3295,N_2941,N_2885);
nand U3296 (N_3296,N_2475,N_2491);
nand U3297 (N_3297,N_2997,N_2670);
nand U3298 (N_3298,N_2943,N_2643);
nor U3299 (N_3299,N_2759,N_2915);
nand U3300 (N_3300,N_2454,N_2890);
and U3301 (N_3301,N_2631,N_2960);
and U3302 (N_3302,N_2498,N_2842);
xnor U3303 (N_3303,N_2586,N_2424);
nor U3304 (N_3304,N_2523,N_2918);
and U3305 (N_3305,N_2744,N_2449);
nand U3306 (N_3306,N_2434,N_2906);
and U3307 (N_3307,N_2809,N_2777);
nor U3308 (N_3308,N_2568,N_2994);
nor U3309 (N_3309,N_2596,N_2668);
nand U3310 (N_3310,N_2744,N_2650);
nor U3311 (N_3311,N_2990,N_2544);
nand U3312 (N_3312,N_2581,N_2629);
or U3313 (N_3313,N_2813,N_2606);
or U3314 (N_3314,N_2548,N_2629);
xor U3315 (N_3315,N_2623,N_2467);
and U3316 (N_3316,N_2968,N_2520);
xor U3317 (N_3317,N_2843,N_2530);
xnor U3318 (N_3318,N_2770,N_2462);
nor U3319 (N_3319,N_2431,N_2503);
or U3320 (N_3320,N_2491,N_2734);
or U3321 (N_3321,N_2644,N_2559);
xnor U3322 (N_3322,N_2624,N_2753);
nor U3323 (N_3323,N_2527,N_2473);
nand U3324 (N_3324,N_2851,N_2909);
xnor U3325 (N_3325,N_2606,N_2409);
nor U3326 (N_3326,N_2960,N_2775);
and U3327 (N_3327,N_2594,N_2401);
nand U3328 (N_3328,N_2998,N_2498);
xor U3329 (N_3329,N_2866,N_2892);
or U3330 (N_3330,N_2756,N_2817);
nor U3331 (N_3331,N_2620,N_2434);
or U3332 (N_3332,N_2624,N_2705);
nand U3333 (N_3333,N_2877,N_2798);
or U3334 (N_3334,N_2852,N_2716);
or U3335 (N_3335,N_2435,N_2586);
and U3336 (N_3336,N_2752,N_2474);
or U3337 (N_3337,N_2697,N_2702);
xor U3338 (N_3338,N_2893,N_2990);
nor U3339 (N_3339,N_2514,N_2638);
xnor U3340 (N_3340,N_2913,N_2907);
nor U3341 (N_3341,N_2604,N_2944);
and U3342 (N_3342,N_2785,N_2402);
or U3343 (N_3343,N_2470,N_2727);
or U3344 (N_3344,N_2635,N_2547);
xor U3345 (N_3345,N_2416,N_2806);
xnor U3346 (N_3346,N_2881,N_2891);
and U3347 (N_3347,N_2687,N_2709);
or U3348 (N_3348,N_2492,N_2435);
xor U3349 (N_3349,N_2631,N_2995);
nor U3350 (N_3350,N_2647,N_2815);
or U3351 (N_3351,N_2973,N_2415);
or U3352 (N_3352,N_2816,N_2683);
xnor U3353 (N_3353,N_2569,N_2879);
and U3354 (N_3354,N_2811,N_2479);
xnor U3355 (N_3355,N_2735,N_2712);
nor U3356 (N_3356,N_2461,N_2557);
nor U3357 (N_3357,N_2951,N_2568);
nand U3358 (N_3358,N_2668,N_2569);
nor U3359 (N_3359,N_2494,N_2749);
nor U3360 (N_3360,N_2744,N_2746);
xnor U3361 (N_3361,N_2612,N_2820);
xnor U3362 (N_3362,N_2919,N_2723);
xnor U3363 (N_3363,N_2579,N_2610);
and U3364 (N_3364,N_2929,N_2783);
or U3365 (N_3365,N_2533,N_2548);
nor U3366 (N_3366,N_2708,N_2934);
or U3367 (N_3367,N_2818,N_2450);
nand U3368 (N_3368,N_2502,N_2761);
and U3369 (N_3369,N_2540,N_2472);
nand U3370 (N_3370,N_2459,N_2444);
nand U3371 (N_3371,N_2890,N_2487);
nand U3372 (N_3372,N_2617,N_2937);
and U3373 (N_3373,N_2480,N_2981);
xor U3374 (N_3374,N_2569,N_2741);
and U3375 (N_3375,N_2535,N_2511);
or U3376 (N_3376,N_2611,N_2574);
and U3377 (N_3377,N_2992,N_2695);
and U3378 (N_3378,N_2766,N_2691);
or U3379 (N_3379,N_2436,N_2960);
xnor U3380 (N_3380,N_2657,N_2887);
and U3381 (N_3381,N_2945,N_2613);
nand U3382 (N_3382,N_2405,N_2534);
xnor U3383 (N_3383,N_2824,N_2606);
nand U3384 (N_3384,N_2883,N_2577);
and U3385 (N_3385,N_2981,N_2846);
and U3386 (N_3386,N_2499,N_2819);
nor U3387 (N_3387,N_2676,N_2419);
and U3388 (N_3388,N_2739,N_2794);
xnor U3389 (N_3389,N_2996,N_2510);
nand U3390 (N_3390,N_2421,N_2472);
nor U3391 (N_3391,N_2676,N_2677);
xnor U3392 (N_3392,N_2489,N_2980);
nor U3393 (N_3393,N_2684,N_2762);
and U3394 (N_3394,N_2655,N_2923);
nor U3395 (N_3395,N_2980,N_2565);
nand U3396 (N_3396,N_2687,N_2498);
nand U3397 (N_3397,N_2463,N_2466);
nor U3398 (N_3398,N_2603,N_2581);
nand U3399 (N_3399,N_2439,N_2417);
xnor U3400 (N_3400,N_2743,N_2896);
and U3401 (N_3401,N_2496,N_2537);
xnor U3402 (N_3402,N_2607,N_2609);
or U3403 (N_3403,N_2592,N_2568);
xnor U3404 (N_3404,N_2935,N_2410);
nand U3405 (N_3405,N_2475,N_2999);
xnor U3406 (N_3406,N_2839,N_2472);
nor U3407 (N_3407,N_2776,N_2878);
and U3408 (N_3408,N_2841,N_2891);
or U3409 (N_3409,N_2946,N_2488);
xor U3410 (N_3410,N_2838,N_2755);
or U3411 (N_3411,N_2953,N_2618);
or U3412 (N_3412,N_2518,N_2851);
xor U3413 (N_3413,N_2869,N_2500);
nor U3414 (N_3414,N_2454,N_2599);
and U3415 (N_3415,N_2443,N_2946);
and U3416 (N_3416,N_2961,N_2937);
or U3417 (N_3417,N_2521,N_2887);
or U3418 (N_3418,N_2472,N_2635);
nand U3419 (N_3419,N_2497,N_2721);
and U3420 (N_3420,N_2934,N_2518);
nand U3421 (N_3421,N_2520,N_2633);
nor U3422 (N_3422,N_2462,N_2862);
xnor U3423 (N_3423,N_2866,N_2864);
or U3424 (N_3424,N_2842,N_2798);
xnor U3425 (N_3425,N_2593,N_2456);
xnor U3426 (N_3426,N_2880,N_2860);
nor U3427 (N_3427,N_2501,N_2590);
nand U3428 (N_3428,N_2504,N_2981);
nor U3429 (N_3429,N_2802,N_2844);
nand U3430 (N_3430,N_2633,N_2649);
nand U3431 (N_3431,N_2410,N_2753);
xnor U3432 (N_3432,N_2672,N_2746);
nand U3433 (N_3433,N_2868,N_2504);
nor U3434 (N_3434,N_2763,N_2957);
nor U3435 (N_3435,N_2760,N_2784);
nand U3436 (N_3436,N_2503,N_2523);
xnor U3437 (N_3437,N_2953,N_2599);
xor U3438 (N_3438,N_2842,N_2508);
nand U3439 (N_3439,N_2852,N_2899);
xor U3440 (N_3440,N_2917,N_2782);
or U3441 (N_3441,N_2930,N_2473);
or U3442 (N_3442,N_2776,N_2546);
nand U3443 (N_3443,N_2789,N_2712);
nand U3444 (N_3444,N_2516,N_2524);
nor U3445 (N_3445,N_2520,N_2488);
and U3446 (N_3446,N_2533,N_2569);
xnor U3447 (N_3447,N_2685,N_2634);
or U3448 (N_3448,N_2844,N_2728);
nand U3449 (N_3449,N_2456,N_2779);
xor U3450 (N_3450,N_2919,N_2800);
nor U3451 (N_3451,N_2629,N_2734);
and U3452 (N_3452,N_2929,N_2907);
xnor U3453 (N_3453,N_2999,N_2518);
and U3454 (N_3454,N_2728,N_2826);
nor U3455 (N_3455,N_2841,N_2621);
xor U3456 (N_3456,N_2622,N_2932);
or U3457 (N_3457,N_2680,N_2473);
nand U3458 (N_3458,N_2479,N_2450);
xor U3459 (N_3459,N_2525,N_2541);
nor U3460 (N_3460,N_2841,N_2984);
or U3461 (N_3461,N_2722,N_2616);
xor U3462 (N_3462,N_2406,N_2849);
and U3463 (N_3463,N_2675,N_2615);
nand U3464 (N_3464,N_2645,N_2534);
xor U3465 (N_3465,N_2511,N_2503);
and U3466 (N_3466,N_2496,N_2834);
and U3467 (N_3467,N_2735,N_2854);
xnor U3468 (N_3468,N_2409,N_2896);
nor U3469 (N_3469,N_2921,N_2911);
xnor U3470 (N_3470,N_2594,N_2835);
nand U3471 (N_3471,N_2968,N_2700);
or U3472 (N_3472,N_2935,N_2605);
nor U3473 (N_3473,N_2942,N_2501);
xor U3474 (N_3474,N_2609,N_2470);
or U3475 (N_3475,N_2561,N_2772);
nor U3476 (N_3476,N_2665,N_2717);
nor U3477 (N_3477,N_2587,N_2939);
xor U3478 (N_3478,N_2943,N_2760);
or U3479 (N_3479,N_2659,N_2625);
or U3480 (N_3480,N_2742,N_2801);
nand U3481 (N_3481,N_2922,N_2912);
and U3482 (N_3482,N_2883,N_2668);
xor U3483 (N_3483,N_2636,N_2813);
nand U3484 (N_3484,N_2741,N_2724);
and U3485 (N_3485,N_2790,N_2915);
xnor U3486 (N_3486,N_2554,N_2970);
nor U3487 (N_3487,N_2774,N_2474);
xnor U3488 (N_3488,N_2634,N_2556);
xnor U3489 (N_3489,N_2866,N_2973);
or U3490 (N_3490,N_2680,N_2750);
or U3491 (N_3491,N_2619,N_2639);
and U3492 (N_3492,N_2508,N_2930);
or U3493 (N_3493,N_2955,N_2421);
or U3494 (N_3494,N_2474,N_2788);
nand U3495 (N_3495,N_2876,N_2730);
nand U3496 (N_3496,N_2903,N_2909);
and U3497 (N_3497,N_2512,N_2607);
or U3498 (N_3498,N_2481,N_2401);
or U3499 (N_3499,N_2861,N_2864);
nand U3500 (N_3500,N_2716,N_2812);
xor U3501 (N_3501,N_2897,N_2714);
nor U3502 (N_3502,N_2894,N_2524);
nand U3503 (N_3503,N_2868,N_2872);
and U3504 (N_3504,N_2941,N_2593);
and U3505 (N_3505,N_2411,N_2581);
xnor U3506 (N_3506,N_2819,N_2951);
nor U3507 (N_3507,N_2861,N_2986);
and U3508 (N_3508,N_2821,N_2752);
or U3509 (N_3509,N_2422,N_2921);
nand U3510 (N_3510,N_2726,N_2991);
nor U3511 (N_3511,N_2415,N_2843);
and U3512 (N_3512,N_2728,N_2481);
nor U3513 (N_3513,N_2781,N_2999);
xnor U3514 (N_3514,N_2420,N_2577);
or U3515 (N_3515,N_2874,N_2952);
xor U3516 (N_3516,N_2818,N_2496);
and U3517 (N_3517,N_2910,N_2602);
xor U3518 (N_3518,N_2444,N_2702);
xor U3519 (N_3519,N_2513,N_2719);
and U3520 (N_3520,N_2952,N_2695);
or U3521 (N_3521,N_2900,N_2894);
nand U3522 (N_3522,N_2930,N_2896);
xnor U3523 (N_3523,N_2678,N_2804);
xnor U3524 (N_3524,N_2772,N_2608);
or U3525 (N_3525,N_2798,N_2745);
and U3526 (N_3526,N_2624,N_2559);
and U3527 (N_3527,N_2934,N_2622);
or U3528 (N_3528,N_2585,N_2916);
and U3529 (N_3529,N_2677,N_2651);
and U3530 (N_3530,N_2742,N_2909);
nor U3531 (N_3531,N_2758,N_2604);
xnor U3532 (N_3532,N_2680,N_2774);
nand U3533 (N_3533,N_2865,N_2422);
nor U3534 (N_3534,N_2875,N_2733);
xor U3535 (N_3535,N_2524,N_2688);
and U3536 (N_3536,N_2967,N_2541);
nand U3537 (N_3537,N_2611,N_2707);
xnor U3538 (N_3538,N_2557,N_2472);
and U3539 (N_3539,N_2694,N_2425);
nand U3540 (N_3540,N_2649,N_2487);
and U3541 (N_3541,N_2700,N_2789);
nor U3542 (N_3542,N_2975,N_2416);
xor U3543 (N_3543,N_2796,N_2704);
or U3544 (N_3544,N_2517,N_2456);
or U3545 (N_3545,N_2944,N_2593);
nor U3546 (N_3546,N_2880,N_2987);
xnor U3547 (N_3547,N_2463,N_2723);
nor U3548 (N_3548,N_2822,N_2840);
xnor U3549 (N_3549,N_2424,N_2898);
and U3550 (N_3550,N_2590,N_2897);
nor U3551 (N_3551,N_2430,N_2712);
and U3552 (N_3552,N_2541,N_2599);
nor U3553 (N_3553,N_2743,N_2645);
nor U3554 (N_3554,N_2722,N_2897);
nor U3555 (N_3555,N_2813,N_2963);
nand U3556 (N_3556,N_2840,N_2428);
xor U3557 (N_3557,N_2854,N_2857);
or U3558 (N_3558,N_2925,N_2993);
or U3559 (N_3559,N_2926,N_2742);
and U3560 (N_3560,N_2509,N_2730);
nand U3561 (N_3561,N_2827,N_2928);
nor U3562 (N_3562,N_2446,N_2713);
nand U3563 (N_3563,N_2854,N_2951);
and U3564 (N_3564,N_2405,N_2605);
and U3565 (N_3565,N_2677,N_2632);
nand U3566 (N_3566,N_2939,N_2985);
or U3567 (N_3567,N_2891,N_2524);
xnor U3568 (N_3568,N_2495,N_2914);
nand U3569 (N_3569,N_2615,N_2841);
nor U3570 (N_3570,N_2628,N_2983);
nand U3571 (N_3571,N_2849,N_2708);
and U3572 (N_3572,N_2823,N_2616);
or U3573 (N_3573,N_2819,N_2927);
and U3574 (N_3574,N_2739,N_2997);
nor U3575 (N_3575,N_2613,N_2734);
nor U3576 (N_3576,N_2540,N_2411);
xor U3577 (N_3577,N_2613,N_2527);
nand U3578 (N_3578,N_2757,N_2928);
and U3579 (N_3579,N_2597,N_2525);
xnor U3580 (N_3580,N_2589,N_2743);
nor U3581 (N_3581,N_2789,N_2865);
nor U3582 (N_3582,N_2973,N_2751);
xor U3583 (N_3583,N_2789,N_2891);
nor U3584 (N_3584,N_2615,N_2444);
nor U3585 (N_3585,N_2437,N_2750);
xor U3586 (N_3586,N_2748,N_2876);
nand U3587 (N_3587,N_2767,N_2920);
nand U3588 (N_3588,N_2443,N_2605);
xnor U3589 (N_3589,N_2994,N_2905);
xor U3590 (N_3590,N_2439,N_2940);
nand U3591 (N_3591,N_2458,N_2894);
and U3592 (N_3592,N_2859,N_2473);
and U3593 (N_3593,N_2736,N_2899);
and U3594 (N_3594,N_2854,N_2732);
or U3595 (N_3595,N_2907,N_2627);
nand U3596 (N_3596,N_2743,N_2882);
and U3597 (N_3597,N_2517,N_2423);
nand U3598 (N_3598,N_2691,N_2476);
and U3599 (N_3599,N_2796,N_2998);
or U3600 (N_3600,N_3016,N_3557);
nor U3601 (N_3601,N_3410,N_3247);
or U3602 (N_3602,N_3260,N_3297);
xnor U3603 (N_3603,N_3519,N_3525);
nand U3604 (N_3604,N_3457,N_3267);
nor U3605 (N_3605,N_3492,N_3469);
nor U3606 (N_3606,N_3331,N_3039);
or U3607 (N_3607,N_3282,N_3143);
nor U3608 (N_3608,N_3361,N_3046);
xor U3609 (N_3609,N_3293,N_3007);
xnor U3610 (N_3610,N_3438,N_3202);
nand U3611 (N_3611,N_3356,N_3238);
nor U3612 (N_3612,N_3230,N_3350);
and U3613 (N_3613,N_3522,N_3237);
and U3614 (N_3614,N_3246,N_3548);
nand U3615 (N_3615,N_3572,N_3164);
and U3616 (N_3616,N_3565,N_3471);
or U3617 (N_3617,N_3132,N_3552);
and U3618 (N_3618,N_3179,N_3461);
nor U3619 (N_3619,N_3270,N_3015);
xnor U3620 (N_3620,N_3449,N_3428);
nand U3621 (N_3621,N_3562,N_3261);
xor U3622 (N_3622,N_3500,N_3392);
xor U3623 (N_3623,N_3545,N_3540);
xnor U3624 (N_3624,N_3386,N_3288);
nand U3625 (N_3625,N_3248,N_3152);
or U3626 (N_3626,N_3187,N_3294);
and U3627 (N_3627,N_3117,N_3052);
and U3628 (N_3628,N_3254,N_3125);
or U3629 (N_3629,N_3466,N_3221);
and U3630 (N_3630,N_3532,N_3534);
nand U3631 (N_3631,N_3343,N_3319);
xor U3632 (N_3632,N_3505,N_3272);
nor U3633 (N_3633,N_3579,N_3121);
xnor U3634 (N_3634,N_3581,N_3175);
and U3635 (N_3635,N_3127,N_3307);
and U3636 (N_3636,N_3425,N_3145);
xnor U3637 (N_3637,N_3169,N_3369);
and U3638 (N_3638,N_3385,N_3456);
or U3639 (N_3639,N_3064,N_3227);
xnor U3640 (N_3640,N_3442,N_3334);
xnor U3641 (N_3641,N_3516,N_3543);
or U3642 (N_3642,N_3234,N_3104);
xnor U3643 (N_3643,N_3223,N_3089);
or U3644 (N_3644,N_3274,N_3322);
and U3645 (N_3645,N_3339,N_3542);
nand U3646 (N_3646,N_3596,N_3417);
nor U3647 (N_3647,N_3368,N_3012);
nor U3648 (N_3648,N_3549,N_3035);
nor U3649 (N_3649,N_3496,N_3241);
and U3650 (N_3650,N_3154,N_3521);
or U3651 (N_3651,N_3219,N_3036);
nor U3652 (N_3652,N_3062,N_3515);
or U3653 (N_3653,N_3533,N_3108);
xor U3654 (N_3654,N_3439,N_3196);
nor U3655 (N_3655,N_3362,N_3432);
or U3656 (N_3656,N_3054,N_3537);
xor U3657 (N_3657,N_3389,N_3049);
and U3658 (N_3658,N_3100,N_3002);
or U3659 (N_3659,N_3069,N_3199);
nor U3660 (N_3660,N_3470,N_3013);
nand U3661 (N_3661,N_3275,N_3024);
xnor U3662 (N_3662,N_3393,N_3245);
xnor U3663 (N_3663,N_3437,N_3277);
nand U3664 (N_3664,N_3053,N_3530);
xor U3665 (N_3665,N_3130,N_3001);
and U3666 (N_3666,N_3255,N_3376);
nor U3667 (N_3667,N_3563,N_3303);
and U3668 (N_3668,N_3229,N_3379);
nor U3669 (N_3669,N_3093,N_3355);
nor U3670 (N_3670,N_3050,N_3008);
or U3671 (N_3671,N_3463,N_3299);
or U3672 (N_3672,N_3281,N_3589);
xor U3673 (N_3673,N_3416,N_3110);
nand U3674 (N_3674,N_3406,N_3091);
and U3675 (N_3675,N_3066,N_3535);
xor U3676 (N_3676,N_3258,N_3482);
or U3677 (N_3677,N_3239,N_3210);
xor U3678 (N_3678,N_3155,N_3375);
and U3679 (N_3679,N_3484,N_3259);
or U3680 (N_3680,N_3403,N_3330);
nand U3681 (N_3681,N_3569,N_3390);
or U3682 (N_3682,N_3311,N_3118);
and U3683 (N_3683,N_3030,N_3273);
nand U3684 (N_3684,N_3211,N_3149);
nor U3685 (N_3685,N_3341,N_3233);
and U3686 (N_3686,N_3265,N_3398);
nor U3687 (N_3687,N_3538,N_3289);
nor U3688 (N_3688,N_3226,N_3171);
xnor U3689 (N_3689,N_3306,N_3436);
nand U3690 (N_3690,N_3166,N_3119);
xor U3691 (N_3691,N_3163,N_3168);
nor U3692 (N_3692,N_3364,N_3550);
and U3693 (N_3693,N_3023,N_3590);
or U3694 (N_3694,N_3314,N_3480);
or U3695 (N_3695,N_3494,N_3367);
nand U3696 (N_3696,N_3508,N_3347);
nand U3697 (N_3697,N_3031,N_3101);
nor U3698 (N_3698,N_3252,N_3283);
xnor U3699 (N_3699,N_3178,N_3065);
nand U3700 (N_3700,N_3597,N_3291);
nor U3701 (N_3701,N_3358,N_3559);
nand U3702 (N_3702,N_3387,N_3526);
and U3703 (N_3703,N_3266,N_3317);
and U3704 (N_3704,N_3029,N_3147);
nand U3705 (N_3705,N_3251,N_3194);
nor U3706 (N_3706,N_3305,N_3408);
or U3707 (N_3707,N_3595,N_3577);
and U3708 (N_3708,N_3099,N_3140);
nand U3709 (N_3709,N_3420,N_3158);
and U3710 (N_3710,N_3103,N_3366);
nor U3711 (N_3711,N_3045,N_3431);
nand U3712 (N_3712,N_3014,N_3396);
nor U3713 (N_3713,N_3573,N_3536);
xnor U3714 (N_3714,N_3399,N_3215);
xor U3715 (N_3715,N_3043,N_3176);
nor U3716 (N_3716,N_3422,N_3198);
nand U3717 (N_3717,N_3181,N_3413);
nor U3718 (N_3718,N_3427,N_3560);
xnor U3719 (N_3719,N_3075,N_3446);
or U3720 (N_3720,N_3025,N_3197);
nand U3721 (N_3721,N_3539,N_3354);
and U3722 (N_3722,N_3070,N_3424);
or U3723 (N_3723,N_3019,N_3076);
or U3724 (N_3724,N_3074,N_3123);
or U3725 (N_3725,N_3495,N_3512);
and U3726 (N_3726,N_3468,N_3598);
xor U3727 (N_3727,N_3524,N_3224);
or U3728 (N_3728,N_3115,N_3477);
nor U3729 (N_3729,N_3060,N_3360);
or U3730 (N_3730,N_3326,N_3095);
and U3731 (N_3731,N_3243,N_3337);
or U3732 (N_3732,N_3483,N_3503);
nor U3733 (N_3733,N_3055,N_3200);
nor U3734 (N_3734,N_3308,N_3284);
or U3735 (N_3735,N_3381,N_3280);
xnor U3736 (N_3736,N_3129,N_3593);
nor U3737 (N_3737,N_3113,N_3434);
xnor U3738 (N_3738,N_3310,N_3068);
and U3739 (N_3739,N_3490,N_3185);
and U3740 (N_3740,N_3498,N_3137);
nand U3741 (N_3741,N_3286,N_3271);
and U3742 (N_3742,N_3038,N_3418);
or U3743 (N_3743,N_3373,N_3067);
or U3744 (N_3744,N_3374,N_3397);
nor U3745 (N_3745,N_3489,N_3454);
xor U3746 (N_3746,N_3208,N_3455);
xor U3747 (N_3747,N_3131,N_3586);
xor U3748 (N_3748,N_3574,N_3499);
or U3749 (N_3749,N_3440,N_3378);
or U3750 (N_3750,N_3201,N_3502);
nand U3751 (N_3751,N_3122,N_3527);
or U3752 (N_3752,N_3567,N_3443);
and U3753 (N_3753,N_3333,N_3472);
nor U3754 (N_3754,N_3059,N_3186);
xnor U3755 (N_3755,N_3004,N_3300);
nand U3756 (N_3756,N_3491,N_3313);
or U3757 (N_3757,N_3507,N_3106);
nor U3758 (N_3758,N_3182,N_3017);
nor U3759 (N_3759,N_3298,N_3405);
or U3760 (N_3760,N_3409,N_3193);
nor U3761 (N_3761,N_3180,N_3142);
or U3762 (N_3762,N_3384,N_3531);
nor U3763 (N_3763,N_3566,N_3128);
or U3764 (N_3764,N_3162,N_3336);
or U3765 (N_3765,N_3287,N_3380);
or U3766 (N_3766,N_3365,N_3412);
nor U3767 (N_3767,N_3433,N_3599);
nand U3768 (N_3768,N_3514,N_3027);
and U3769 (N_3769,N_3085,N_3558);
xor U3770 (N_3770,N_3098,N_3033);
or U3771 (N_3771,N_3585,N_3444);
nor U3772 (N_3772,N_3555,N_3086);
nand U3773 (N_3773,N_3421,N_3005);
nand U3774 (N_3774,N_3203,N_3034);
or U3775 (N_3775,N_3415,N_3309);
xor U3776 (N_3776,N_3269,N_3081);
nand U3777 (N_3777,N_3506,N_3316);
and U3778 (N_3778,N_3077,N_3020);
xnor U3779 (N_3779,N_3195,N_3032);
nand U3780 (N_3780,N_3414,N_3304);
xor U3781 (N_3781,N_3071,N_3096);
nor U3782 (N_3782,N_3395,N_3458);
nor U3783 (N_3783,N_3473,N_3445);
nand U3784 (N_3784,N_3006,N_3167);
nor U3785 (N_3785,N_3231,N_3325);
nand U3786 (N_3786,N_3570,N_3429);
nand U3787 (N_3787,N_3173,N_3497);
and U3788 (N_3788,N_3301,N_3544);
nand U3789 (N_3789,N_3450,N_3553);
and U3790 (N_3790,N_3134,N_3587);
nand U3791 (N_3791,N_3292,N_3547);
and U3792 (N_3792,N_3107,N_3467);
nor U3793 (N_3793,N_3150,N_3112);
and U3794 (N_3794,N_3357,N_3353);
nor U3795 (N_3795,N_3047,N_3584);
nand U3796 (N_3796,N_3236,N_3235);
or U3797 (N_3797,N_3401,N_3160);
and U3798 (N_3798,N_3009,N_3441);
xnor U3799 (N_3799,N_3411,N_3486);
xor U3800 (N_3800,N_3504,N_3592);
xor U3801 (N_3801,N_3509,N_3188);
xor U3802 (N_3802,N_3591,N_3352);
xnor U3803 (N_3803,N_3323,N_3189);
nor U3804 (N_3804,N_3138,N_3102);
nor U3805 (N_3805,N_3370,N_3161);
xor U3806 (N_3806,N_3568,N_3092);
nand U3807 (N_3807,N_3133,N_3459);
xor U3808 (N_3808,N_3109,N_3232);
nor U3809 (N_3809,N_3476,N_3391);
xnor U3810 (N_3810,N_3529,N_3351);
or U3811 (N_3811,N_3513,N_3148);
or U3812 (N_3812,N_3213,N_3453);
nand U3813 (N_3813,N_3580,N_3146);
and U3814 (N_3814,N_3359,N_3426);
or U3815 (N_3815,N_3262,N_3296);
or U3816 (N_3816,N_3153,N_3090);
xor U3817 (N_3817,N_3157,N_3372);
xnor U3818 (N_3818,N_3192,N_3225);
xor U3819 (N_3819,N_3315,N_3402);
or U3820 (N_3820,N_3217,N_3430);
nand U3821 (N_3821,N_3487,N_3183);
and U3822 (N_3822,N_3464,N_3087);
or U3823 (N_3823,N_3207,N_3051);
nor U3824 (N_3824,N_3022,N_3377);
or U3825 (N_3825,N_3478,N_3320);
or U3826 (N_3826,N_3041,N_3465);
or U3827 (N_3827,N_3249,N_3321);
and U3828 (N_3828,N_3312,N_3072);
and U3829 (N_3829,N_3242,N_3061);
xor U3830 (N_3830,N_3204,N_3554);
nor U3831 (N_3831,N_3080,N_3268);
xor U3832 (N_3832,N_3481,N_3493);
xnor U3833 (N_3833,N_3010,N_3250);
nor U3834 (N_3834,N_3578,N_3407);
nor U3835 (N_3835,N_3165,N_3510);
and U3836 (N_3836,N_3105,N_3528);
or U3837 (N_3837,N_3342,N_3551);
xor U3838 (N_3838,N_3063,N_3139);
nand U3839 (N_3839,N_3058,N_3363);
xnor U3840 (N_3840,N_3214,N_3400);
xnor U3841 (N_3841,N_3575,N_3170);
nor U3842 (N_3842,N_3114,N_3571);
nor U3843 (N_3843,N_3044,N_3003);
or U3844 (N_3844,N_3518,N_3040);
and U3845 (N_3845,N_3244,N_3345);
and U3846 (N_3846,N_3037,N_3371);
nand U3847 (N_3847,N_3073,N_3257);
or U3848 (N_3848,N_3448,N_3561);
nor U3849 (N_3849,N_3388,N_3256);
nor U3850 (N_3850,N_3088,N_3462);
or U3851 (N_3851,N_3348,N_3346);
nor U3852 (N_3852,N_3159,N_3057);
nand U3853 (N_3853,N_3460,N_3151);
nor U3854 (N_3854,N_3338,N_3276);
and U3855 (N_3855,N_3135,N_3588);
nand U3856 (N_3856,N_3290,N_3517);
nor U3857 (N_3857,N_3141,N_3501);
and U3858 (N_3858,N_3028,N_3156);
xor U3859 (N_3859,N_3329,N_3488);
or U3860 (N_3860,N_3048,N_3000);
or U3861 (N_3861,N_3324,N_3011);
or U3862 (N_3862,N_3253,N_3279);
nand U3863 (N_3863,N_3382,N_3452);
nand U3864 (N_3864,N_3594,N_3228);
xnor U3865 (N_3865,N_3190,N_3332);
and U3866 (N_3866,N_3564,N_3479);
or U3867 (N_3867,N_3511,N_3344);
nand U3868 (N_3868,N_3318,N_3419);
nor U3869 (N_3869,N_3126,N_3383);
or U3870 (N_3870,N_3447,N_3328);
and U3871 (N_3871,N_3079,N_3205);
nand U3872 (N_3872,N_3084,N_3177);
xnor U3873 (N_3873,N_3451,N_3124);
xor U3874 (N_3874,N_3523,N_3172);
or U3875 (N_3875,N_3191,N_3435);
nand U3876 (N_3876,N_3018,N_3335);
xnor U3877 (N_3877,N_3404,N_3546);
nand U3878 (N_3878,N_3520,N_3206);
nor U3879 (N_3879,N_3097,N_3263);
or U3880 (N_3880,N_3026,N_3184);
and U3881 (N_3881,N_3485,N_3082);
and U3882 (N_3882,N_3264,N_3136);
xor U3883 (N_3883,N_3216,N_3218);
xnor U3884 (N_3884,N_3285,N_3349);
or U3885 (N_3885,N_3042,N_3094);
xnor U3886 (N_3886,N_3116,N_3056);
nor U3887 (N_3887,N_3222,N_3475);
or U3888 (N_3888,N_3174,N_3278);
or U3889 (N_3889,N_3302,N_3220);
or U3890 (N_3890,N_3582,N_3078);
nand U3891 (N_3891,N_3144,N_3240);
nand U3892 (N_3892,N_3576,N_3340);
and U3893 (N_3893,N_3209,N_3111);
xor U3894 (N_3894,N_3541,N_3083);
and U3895 (N_3895,N_3021,N_3583);
and U3896 (N_3896,N_3295,N_3327);
and U3897 (N_3897,N_3556,N_3120);
nand U3898 (N_3898,N_3423,N_3394);
or U3899 (N_3899,N_3474,N_3212);
nand U3900 (N_3900,N_3521,N_3409);
xor U3901 (N_3901,N_3080,N_3044);
or U3902 (N_3902,N_3288,N_3118);
or U3903 (N_3903,N_3522,N_3423);
or U3904 (N_3904,N_3207,N_3490);
xor U3905 (N_3905,N_3378,N_3522);
nand U3906 (N_3906,N_3507,N_3086);
or U3907 (N_3907,N_3317,N_3472);
nor U3908 (N_3908,N_3303,N_3177);
nor U3909 (N_3909,N_3209,N_3489);
xor U3910 (N_3910,N_3207,N_3026);
and U3911 (N_3911,N_3061,N_3554);
xor U3912 (N_3912,N_3329,N_3126);
nand U3913 (N_3913,N_3362,N_3211);
nor U3914 (N_3914,N_3477,N_3122);
and U3915 (N_3915,N_3364,N_3378);
and U3916 (N_3916,N_3529,N_3506);
nand U3917 (N_3917,N_3198,N_3277);
nor U3918 (N_3918,N_3018,N_3567);
and U3919 (N_3919,N_3121,N_3506);
xnor U3920 (N_3920,N_3052,N_3275);
xnor U3921 (N_3921,N_3373,N_3483);
or U3922 (N_3922,N_3529,N_3451);
nand U3923 (N_3923,N_3442,N_3213);
xnor U3924 (N_3924,N_3069,N_3216);
nand U3925 (N_3925,N_3248,N_3463);
nor U3926 (N_3926,N_3104,N_3176);
nor U3927 (N_3927,N_3185,N_3592);
or U3928 (N_3928,N_3117,N_3297);
and U3929 (N_3929,N_3246,N_3586);
or U3930 (N_3930,N_3265,N_3374);
nor U3931 (N_3931,N_3528,N_3152);
or U3932 (N_3932,N_3523,N_3317);
xor U3933 (N_3933,N_3359,N_3536);
nand U3934 (N_3934,N_3047,N_3297);
or U3935 (N_3935,N_3518,N_3086);
nor U3936 (N_3936,N_3145,N_3106);
nor U3937 (N_3937,N_3239,N_3472);
xor U3938 (N_3938,N_3067,N_3199);
or U3939 (N_3939,N_3203,N_3217);
nor U3940 (N_3940,N_3276,N_3155);
or U3941 (N_3941,N_3031,N_3395);
xor U3942 (N_3942,N_3452,N_3102);
xor U3943 (N_3943,N_3489,N_3457);
or U3944 (N_3944,N_3514,N_3128);
nand U3945 (N_3945,N_3351,N_3272);
nand U3946 (N_3946,N_3586,N_3334);
nor U3947 (N_3947,N_3111,N_3497);
nor U3948 (N_3948,N_3000,N_3512);
and U3949 (N_3949,N_3281,N_3285);
nand U3950 (N_3950,N_3233,N_3391);
and U3951 (N_3951,N_3357,N_3334);
and U3952 (N_3952,N_3145,N_3068);
and U3953 (N_3953,N_3403,N_3472);
and U3954 (N_3954,N_3542,N_3408);
and U3955 (N_3955,N_3260,N_3145);
xor U3956 (N_3956,N_3009,N_3584);
and U3957 (N_3957,N_3364,N_3243);
xor U3958 (N_3958,N_3073,N_3239);
nand U3959 (N_3959,N_3044,N_3491);
and U3960 (N_3960,N_3063,N_3330);
or U3961 (N_3961,N_3581,N_3447);
or U3962 (N_3962,N_3526,N_3277);
nor U3963 (N_3963,N_3537,N_3073);
or U3964 (N_3964,N_3333,N_3033);
nand U3965 (N_3965,N_3098,N_3535);
or U3966 (N_3966,N_3521,N_3086);
nand U3967 (N_3967,N_3081,N_3360);
xnor U3968 (N_3968,N_3154,N_3393);
and U3969 (N_3969,N_3373,N_3271);
xor U3970 (N_3970,N_3372,N_3143);
nor U3971 (N_3971,N_3500,N_3574);
nor U3972 (N_3972,N_3070,N_3193);
or U3973 (N_3973,N_3376,N_3012);
nand U3974 (N_3974,N_3029,N_3079);
nor U3975 (N_3975,N_3112,N_3566);
xnor U3976 (N_3976,N_3044,N_3216);
or U3977 (N_3977,N_3093,N_3526);
nor U3978 (N_3978,N_3397,N_3084);
and U3979 (N_3979,N_3422,N_3121);
or U3980 (N_3980,N_3427,N_3122);
nand U3981 (N_3981,N_3478,N_3216);
nor U3982 (N_3982,N_3391,N_3330);
or U3983 (N_3983,N_3427,N_3406);
nor U3984 (N_3984,N_3298,N_3524);
nand U3985 (N_3985,N_3167,N_3410);
or U3986 (N_3986,N_3098,N_3077);
xnor U3987 (N_3987,N_3463,N_3447);
nor U3988 (N_3988,N_3110,N_3515);
or U3989 (N_3989,N_3309,N_3180);
or U3990 (N_3990,N_3332,N_3527);
nand U3991 (N_3991,N_3504,N_3432);
and U3992 (N_3992,N_3089,N_3203);
xnor U3993 (N_3993,N_3558,N_3329);
nor U3994 (N_3994,N_3573,N_3447);
xnor U3995 (N_3995,N_3057,N_3299);
and U3996 (N_3996,N_3282,N_3460);
xnor U3997 (N_3997,N_3468,N_3234);
or U3998 (N_3998,N_3529,N_3114);
or U3999 (N_3999,N_3373,N_3100);
and U4000 (N_4000,N_3354,N_3058);
xor U4001 (N_4001,N_3589,N_3465);
nor U4002 (N_4002,N_3010,N_3457);
nand U4003 (N_4003,N_3556,N_3097);
nor U4004 (N_4004,N_3002,N_3017);
and U4005 (N_4005,N_3238,N_3186);
xnor U4006 (N_4006,N_3456,N_3318);
nand U4007 (N_4007,N_3513,N_3594);
or U4008 (N_4008,N_3408,N_3219);
xor U4009 (N_4009,N_3117,N_3266);
nor U4010 (N_4010,N_3576,N_3582);
xor U4011 (N_4011,N_3226,N_3168);
nor U4012 (N_4012,N_3496,N_3139);
xor U4013 (N_4013,N_3449,N_3239);
or U4014 (N_4014,N_3070,N_3272);
xnor U4015 (N_4015,N_3437,N_3154);
xor U4016 (N_4016,N_3457,N_3312);
xnor U4017 (N_4017,N_3231,N_3240);
and U4018 (N_4018,N_3289,N_3429);
or U4019 (N_4019,N_3383,N_3567);
nand U4020 (N_4020,N_3464,N_3250);
nand U4021 (N_4021,N_3458,N_3318);
nand U4022 (N_4022,N_3130,N_3303);
and U4023 (N_4023,N_3516,N_3175);
nand U4024 (N_4024,N_3112,N_3442);
nor U4025 (N_4025,N_3549,N_3438);
nor U4026 (N_4026,N_3276,N_3523);
nand U4027 (N_4027,N_3015,N_3115);
nand U4028 (N_4028,N_3202,N_3471);
nand U4029 (N_4029,N_3124,N_3549);
xor U4030 (N_4030,N_3349,N_3594);
nand U4031 (N_4031,N_3027,N_3429);
nor U4032 (N_4032,N_3380,N_3099);
nand U4033 (N_4033,N_3077,N_3396);
nand U4034 (N_4034,N_3127,N_3228);
xnor U4035 (N_4035,N_3284,N_3262);
and U4036 (N_4036,N_3385,N_3531);
and U4037 (N_4037,N_3063,N_3151);
xnor U4038 (N_4038,N_3055,N_3462);
nand U4039 (N_4039,N_3153,N_3193);
nand U4040 (N_4040,N_3587,N_3011);
nand U4041 (N_4041,N_3181,N_3480);
or U4042 (N_4042,N_3053,N_3072);
or U4043 (N_4043,N_3076,N_3330);
or U4044 (N_4044,N_3131,N_3064);
and U4045 (N_4045,N_3255,N_3197);
nand U4046 (N_4046,N_3465,N_3279);
or U4047 (N_4047,N_3278,N_3048);
xnor U4048 (N_4048,N_3216,N_3389);
xnor U4049 (N_4049,N_3238,N_3477);
and U4050 (N_4050,N_3452,N_3034);
and U4051 (N_4051,N_3270,N_3063);
and U4052 (N_4052,N_3200,N_3344);
xor U4053 (N_4053,N_3582,N_3472);
nor U4054 (N_4054,N_3150,N_3057);
or U4055 (N_4055,N_3507,N_3470);
nor U4056 (N_4056,N_3146,N_3188);
nand U4057 (N_4057,N_3468,N_3193);
or U4058 (N_4058,N_3149,N_3462);
nand U4059 (N_4059,N_3077,N_3232);
nand U4060 (N_4060,N_3388,N_3595);
nand U4061 (N_4061,N_3530,N_3066);
nand U4062 (N_4062,N_3289,N_3299);
and U4063 (N_4063,N_3398,N_3552);
nand U4064 (N_4064,N_3274,N_3225);
or U4065 (N_4065,N_3158,N_3595);
and U4066 (N_4066,N_3102,N_3281);
and U4067 (N_4067,N_3365,N_3199);
nand U4068 (N_4068,N_3332,N_3562);
or U4069 (N_4069,N_3398,N_3203);
and U4070 (N_4070,N_3032,N_3158);
nor U4071 (N_4071,N_3554,N_3574);
nand U4072 (N_4072,N_3501,N_3418);
or U4073 (N_4073,N_3082,N_3515);
or U4074 (N_4074,N_3313,N_3146);
nand U4075 (N_4075,N_3490,N_3136);
xnor U4076 (N_4076,N_3458,N_3335);
xor U4077 (N_4077,N_3575,N_3169);
nor U4078 (N_4078,N_3516,N_3384);
or U4079 (N_4079,N_3003,N_3546);
and U4080 (N_4080,N_3227,N_3151);
xor U4081 (N_4081,N_3439,N_3477);
nor U4082 (N_4082,N_3404,N_3020);
and U4083 (N_4083,N_3177,N_3130);
nor U4084 (N_4084,N_3500,N_3220);
nor U4085 (N_4085,N_3035,N_3427);
nand U4086 (N_4086,N_3026,N_3192);
nand U4087 (N_4087,N_3104,N_3036);
nand U4088 (N_4088,N_3007,N_3271);
nor U4089 (N_4089,N_3098,N_3534);
xor U4090 (N_4090,N_3090,N_3517);
and U4091 (N_4091,N_3066,N_3155);
and U4092 (N_4092,N_3353,N_3173);
nand U4093 (N_4093,N_3191,N_3576);
and U4094 (N_4094,N_3107,N_3119);
and U4095 (N_4095,N_3159,N_3133);
and U4096 (N_4096,N_3126,N_3314);
and U4097 (N_4097,N_3437,N_3460);
or U4098 (N_4098,N_3139,N_3358);
and U4099 (N_4099,N_3204,N_3113);
nand U4100 (N_4100,N_3320,N_3567);
or U4101 (N_4101,N_3025,N_3307);
nor U4102 (N_4102,N_3324,N_3145);
nor U4103 (N_4103,N_3058,N_3105);
nor U4104 (N_4104,N_3475,N_3339);
and U4105 (N_4105,N_3469,N_3544);
xnor U4106 (N_4106,N_3122,N_3258);
xor U4107 (N_4107,N_3587,N_3043);
and U4108 (N_4108,N_3091,N_3465);
and U4109 (N_4109,N_3533,N_3561);
nor U4110 (N_4110,N_3012,N_3299);
or U4111 (N_4111,N_3391,N_3505);
and U4112 (N_4112,N_3209,N_3220);
nand U4113 (N_4113,N_3463,N_3162);
and U4114 (N_4114,N_3118,N_3407);
nand U4115 (N_4115,N_3480,N_3148);
and U4116 (N_4116,N_3149,N_3189);
nor U4117 (N_4117,N_3247,N_3549);
or U4118 (N_4118,N_3583,N_3194);
xnor U4119 (N_4119,N_3525,N_3570);
xnor U4120 (N_4120,N_3588,N_3496);
nand U4121 (N_4121,N_3295,N_3336);
xor U4122 (N_4122,N_3255,N_3015);
xnor U4123 (N_4123,N_3195,N_3141);
and U4124 (N_4124,N_3002,N_3444);
or U4125 (N_4125,N_3597,N_3556);
and U4126 (N_4126,N_3365,N_3023);
and U4127 (N_4127,N_3461,N_3558);
nand U4128 (N_4128,N_3249,N_3136);
xnor U4129 (N_4129,N_3238,N_3468);
or U4130 (N_4130,N_3134,N_3556);
and U4131 (N_4131,N_3140,N_3105);
nand U4132 (N_4132,N_3090,N_3580);
or U4133 (N_4133,N_3422,N_3204);
nor U4134 (N_4134,N_3012,N_3358);
nand U4135 (N_4135,N_3364,N_3466);
xor U4136 (N_4136,N_3267,N_3098);
and U4137 (N_4137,N_3003,N_3359);
xor U4138 (N_4138,N_3225,N_3277);
nor U4139 (N_4139,N_3597,N_3494);
or U4140 (N_4140,N_3534,N_3297);
nor U4141 (N_4141,N_3215,N_3401);
nor U4142 (N_4142,N_3070,N_3107);
or U4143 (N_4143,N_3262,N_3033);
and U4144 (N_4144,N_3367,N_3551);
or U4145 (N_4145,N_3290,N_3453);
nor U4146 (N_4146,N_3214,N_3285);
and U4147 (N_4147,N_3351,N_3490);
or U4148 (N_4148,N_3507,N_3592);
nand U4149 (N_4149,N_3379,N_3517);
and U4150 (N_4150,N_3125,N_3548);
nor U4151 (N_4151,N_3517,N_3415);
and U4152 (N_4152,N_3289,N_3567);
and U4153 (N_4153,N_3436,N_3472);
or U4154 (N_4154,N_3447,N_3100);
xor U4155 (N_4155,N_3503,N_3021);
nand U4156 (N_4156,N_3124,N_3233);
nor U4157 (N_4157,N_3021,N_3211);
and U4158 (N_4158,N_3014,N_3495);
or U4159 (N_4159,N_3297,N_3111);
xnor U4160 (N_4160,N_3025,N_3498);
nand U4161 (N_4161,N_3011,N_3137);
or U4162 (N_4162,N_3328,N_3178);
or U4163 (N_4163,N_3373,N_3201);
nor U4164 (N_4164,N_3372,N_3165);
or U4165 (N_4165,N_3361,N_3490);
nor U4166 (N_4166,N_3387,N_3543);
or U4167 (N_4167,N_3206,N_3537);
nor U4168 (N_4168,N_3322,N_3091);
or U4169 (N_4169,N_3420,N_3513);
xor U4170 (N_4170,N_3400,N_3471);
and U4171 (N_4171,N_3251,N_3094);
and U4172 (N_4172,N_3356,N_3114);
nand U4173 (N_4173,N_3076,N_3589);
nand U4174 (N_4174,N_3343,N_3261);
xor U4175 (N_4175,N_3099,N_3223);
nand U4176 (N_4176,N_3378,N_3033);
and U4177 (N_4177,N_3171,N_3127);
and U4178 (N_4178,N_3483,N_3480);
and U4179 (N_4179,N_3471,N_3234);
nand U4180 (N_4180,N_3279,N_3343);
or U4181 (N_4181,N_3210,N_3533);
or U4182 (N_4182,N_3304,N_3310);
and U4183 (N_4183,N_3052,N_3516);
xor U4184 (N_4184,N_3109,N_3216);
nor U4185 (N_4185,N_3561,N_3443);
xnor U4186 (N_4186,N_3507,N_3384);
nor U4187 (N_4187,N_3426,N_3030);
and U4188 (N_4188,N_3087,N_3284);
or U4189 (N_4189,N_3341,N_3207);
xor U4190 (N_4190,N_3141,N_3576);
or U4191 (N_4191,N_3314,N_3330);
or U4192 (N_4192,N_3069,N_3533);
and U4193 (N_4193,N_3588,N_3444);
nand U4194 (N_4194,N_3552,N_3298);
nor U4195 (N_4195,N_3272,N_3392);
xor U4196 (N_4196,N_3592,N_3243);
nor U4197 (N_4197,N_3264,N_3212);
or U4198 (N_4198,N_3084,N_3081);
nor U4199 (N_4199,N_3440,N_3381);
nor U4200 (N_4200,N_3638,N_3990);
nand U4201 (N_4201,N_4196,N_3628);
or U4202 (N_4202,N_3823,N_3946);
or U4203 (N_4203,N_3917,N_3716);
xnor U4204 (N_4204,N_3674,N_3878);
xor U4205 (N_4205,N_3707,N_4161);
xor U4206 (N_4206,N_3774,N_3689);
and U4207 (N_4207,N_3789,N_4007);
xnor U4208 (N_4208,N_3755,N_4146);
xor U4209 (N_4209,N_3943,N_4117);
nor U4210 (N_4210,N_4049,N_4110);
xnor U4211 (N_4211,N_3736,N_3907);
xnor U4212 (N_4212,N_3659,N_3658);
nand U4213 (N_4213,N_3935,N_3937);
or U4214 (N_4214,N_3934,N_3957);
and U4215 (N_4215,N_3792,N_3999);
or U4216 (N_4216,N_4043,N_4154);
xor U4217 (N_4217,N_3810,N_4119);
or U4218 (N_4218,N_3657,N_3858);
xnor U4219 (N_4219,N_3874,N_3720);
xnor U4220 (N_4220,N_4030,N_3992);
or U4221 (N_4221,N_3710,N_3717);
xnor U4222 (N_4222,N_4099,N_4014);
and U4223 (N_4223,N_4063,N_3954);
nor U4224 (N_4224,N_3600,N_4003);
and U4225 (N_4225,N_4139,N_4097);
xnor U4226 (N_4226,N_3651,N_3904);
nor U4227 (N_4227,N_3682,N_3699);
or U4228 (N_4228,N_3884,N_4194);
and U4229 (N_4229,N_4101,N_4142);
and U4230 (N_4230,N_3741,N_3773);
nor U4231 (N_4231,N_3841,N_3980);
xor U4232 (N_4232,N_4090,N_3967);
nand U4233 (N_4233,N_4048,N_4164);
nor U4234 (N_4234,N_3860,N_3897);
xor U4235 (N_4235,N_3760,N_3681);
or U4236 (N_4236,N_3742,N_4165);
xor U4237 (N_4237,N_3795,N_4172);
and U4238 (N_4238,N_3777,N_3608);
or U4239 (N_4239,N_3619,N_4198);
xnor U4240 (N_4240,N_3863,N_3632);
xor U4241 (N_4241,N_3613,N_3728);
or U4242 (N_4242,N_3840,N_3708);
nand U4243 (N_4243,N_4183,N_3704);
xor U4244 (N_4244,N_3988,N_3656);
nor U4245 (N_4245,N_3743,N_3969);
or U4246 (N_4246,N_4078,N_3664);
nor U4247 (N_4247,N_3861,N_3997);
nor U4248 (N_4248,N_3756,N_3703);
nand U4249 (N_4249,N_4122,N_4088);
or U4250 (N_4250,N_3695,N_3796);
nand U4251 (N_4251,N_4096,N_4190);
or U4252 (N_4252,N_4103,N_3791);
nor U4253 (N_4253,N_3763,N_3782);
nand U4254 (N_4254,N_4051,N_4153);
nor U4255 (N_4255,N_4020,N_4121);
and U4256 (N_4256,N_3733,N_3601);
or U4257 (N_4257,N_3855,N_3962);
and U4258 (N_4258,N_3652,N_3690);
xnor U4259 (N_4259,N_4176,N_3891);
xor U4260 (N_4260,N_4187,N_4150);
nor U4261 (N_4261,N_3642,N_3993);
nor U4262 (N_4262,N_3625,N_4108);
nand U4263 (N_4263,N_4126,N_3781);
xor U4264 (N_4264,N_3916,N_4156);
nand U4265 (N_4265,N_3768,N_3872);
nor U4266 (N_4266,N_3772,N_4174);
nor U4267 (N_4267,N_4180,N_3623);
and U4268 (N_4268,N_3800,N_3824);
and U4269 (N_4269,N_4076,N_3888);
xnor U4270 (N_4270,N_3744,N_3815);
nor U4271 (N_4271,N_3764,N_3746);
nand U4272 (N_4272,N_4045,N_3955);
nand U4273 (N_4273,N_3953,N_3844);
nor U4274 (N_4274,N_4042,N_4177);
nor U4275 (N_4275,N_3668,N_3856);
nor U4276 (N_4276,N_4107,N_3867);
and U4277 (N_4277,N_4105,N_4009);
nor U4278 (N_4278,N_3759,N_3762);
or U4279 (N_4279,N_4114,N_3678);
nor U4280 (N_4280,N_3942,N_3665);
or U4281 (N_4281,N_3940,N_3846);
and U4282 (N_4282,N_3958,N_3731);
xor U4283 (N_4283,N_3926,N_3821);
nand U4284 (N_4284,N_4140,N_3732);
nor U4285 (N_4285,N_3948,N_3718);
or U4286 (N_4286,N_4016,N_4124);
nand U4287 (N_4287,N_3661,N_4116);
or U4288 (N_4288,N_3735,N_4129);
nand U4289 (N_4289,N_4072,N_4035);
nand U4290 (N_4290,N_3713,N_3910);
or U4291 (N_4291,N_3802,N_3603);
or U4292 (N_4292,N_3620,N_4132);
nand U4293 (N_4293,N_3711,N_4143);
xnor U4294 (N_4294,N_4037,N_3751);
nand U4295 (N_4295,N_3672,N_3694);
nand U4296 (N_4296,N_4133,N_3783);
or U4297 (N_4297,N_3837,N_3780);
or U4298 (N_4298,N_4015,N_4098);
xor U4299 (N_4299,N_3941,N_3696);
nor U4300 (N_4300,N_3831,N_3998);
xnor U4301 (N_4301,N_3947,N_3982);
and U4302 (N_4302,N_4024,N_3684);
or U4303 (N_4303,N_4111,N_4064);
and U4304 (N_4304,N_3881,N_4120);
nor U4305 (N_4305,N_3790,N_3828);
nor U4306 (N_4306,N_3983,N_3912);
xnor U4307 (N_4307,N_3859,N_3750);
and U4308 (N_4308,N_3626,N_3706);
or U4309 (N_4309,N_3775,N_4080);
xor U4310 (N_4310,N_3921,N_3933);
or U4311 (N_4311,N_3676,N_3911);
nor U4312 (N_4312,N_3972,N_3893);
or U4313 (N_4313,N_4004,N_3932);
nor U4314 (N_4314,N_3938,N_4027);
nor U4315 (N_4315,N_3637,N_3956);
or U4316 (N_4316,N_3719,N_4085);
nor U4317 (N_4317,N_3857,N_4145);
xnor U4318 (N_4318,N_3922,N_3639);
xor U4319 (N_4319,N_3989,N_3776);
and U4320 (N_4320,N_4001,N_4199);
nor U4321 (N_4321,N_3739,N_4025);
nor U4322 (N_4322,N_4029,N_3974);
or U4323 (N_4323,N_3987,N_3865);
and U4324 (N_4324,N_4141,N_3927);
nand U4325 (N_4325,N_3849,N_3692);
nor U4326 (N_4326,N_3675,N_3757);
nor U4327 (N_4327,N_3968,N_3687);
nand U4328 (N_4328,N_4059,N_3712);
or U4329 (N_4329,N_4022,N_3648);
nor U4330 (N_4330,N_3877,N_3970);
xnor U4331 (N_4331,N_3753,N_3666);
nor U4332 (N_4332,N_3747,N_3622);
or U4333 (N_4333,N_4012,N_3729);
and U4334 (N_4334,N_3929,N_3787);
or U4335 (N_4335,N_3965,N_3793);
nor U4336 (N_4336,N_3645,N_3723);
nor U4337 (N_4337,N_4131,N_4047);
nor U4338 (N_4338,N_3767,N_3701);
and U4339 (N_4339,N_3890,N_3848);
or U4340 (N_4340,N_4005,N_3818);
or U4341 (N_4341,N_4056,N_3680);
nor U4342 (N_4342,N_4152,N_3944);
or U4343 (N_4343,N_3852,N_3770);
nand U4344 (N_4344,N_3646,N_3727);
nor U4345 (N_4345,N_3838,N_3901);
nand U4346 (N_4346,N_3709,N_3918);
xor U4347 (N_4347,N_4044,N_3900);
or U4348 (N_4348,N_3612,N_3914);
xor U4349 (N_4349,N_3794,N_3685);
nand U4350 (N_4350,N_4192,N_3930);
and U4351 (N_4351,N_3977,N_4109);
xnor U4352 (N_4352,N_4128,N_3730);
nor U4353 (N_4353,N_3995,N_4070);
nand U4354 (N_4354,N_3928,N_3906);
nor U4355 (N_4355,N_3816,N_3850);
xnor U4356 (N_4356,N_4036,N_3640);
xnor U4357 (N_4357,N_3715,N_3931);
xor U4358 (N_4358,N_4054,N_4082);
nand U4359 (N_4359,N_4055,N_4134);
nand U4360 (N_4360,N_4157,N_4106);
and U4361 (N_4361,N_3905,N_3845);
xor U4362 (N_4362,N_3961,N_4125);
and U4363 (N_4363,N_3984,N_4130);
nand U4364 (N_4364,N_3978,N_3761);
and U4365 (N_4365,N_3631,N_3740);
xor U4366 (N_4366,N_4017,N_3679);
or U4367 (N_4367,N_3805,N_3667);
nand U4368 (N_4368,N_3809,N_3827);
and U4369 (N_4369,N_4040,N_3976);
xnor U4370 (N_4370,N_4195,N_3839);
xnor U4371 (N_4371,N_3876,N_3871);
nor U4372 (N_4372,N_4135,N_4178);
xnor U4373 (N_4373,N_4094,N_3721);
or U4374 (N_4374,N_4053,N_4188);
or U4375 (N_4375,N_3745,N_3804);
xor U4376 (N_4376,N_3722,N_3610);
or U4377 (N_4377,N_4158,N_4093);
nor U4378 (N_4378,N_4175,N_3811);
xnor U4379 (N_4379,N_4184,N_4091);
and U4380 (N_4380,N_3886,N_4127);
nand U4381 (N_4381,N_3605,N_3996);
nor U4382 (N_4382,N_4112,N_3683);
nand U4383 (N_4383,N_3749,N_4067);
and U4384 (N_4384,N_3862,N_3950);
nand U4385 (N_4385,N_3644,N_4060);
nor U4386 (N_4386,N_3985,N_3691);
or U4387 (N_4387,N_4046,N_4197);
xnor U4388 (N_4388,N_4113,N_3766);
and U4389 (N_4389,N_4170,N_3892);
xor U4390 (N_4390,N_3662,N_4100);
nand U4391 (N_4391,N_3959,N_3836);
xnor U4392 (N_4392,N_3633,N_3653);
nand U4393 (N_4393,N_4031,N_4034);
xnor U4394 (N_4394,N_3788,N_4050);
or U4395 (N_4395,N_3909,N_4074);
nor U4396 (N_4396,N_3686,N_3971);
xor U4397 (N_4397,N_4166,N_4137);
and U4398 (N_4398,N_3634,N_3797);
and U4399 (N_4399,N_4081,N_3864);
or U4400 (N_4400,N_4002,N_4104);
nand U4401 (N_4401,N_3785,N_3835);
xor U4402 (N_4402,N_3737,N_4039);
and U4403 (N_4403,N_3896,N_4167);
xnor U4404 (N_4404,N_4052,N_4061);
and U4405 (N_4405,N_3808,N_3758);
nand U4406 (N_4406,N_4102,N_3847);
nor U4407 (N_4407,N_3812,N_3677);
xor U4408 (N_4408,N_3611,N_3643);
nand U4409 (N_4409,N_3842,N_3923);
xor U4410 (N_4410,N_3834,N_4148);
xor U4411 (N_4411,N_3616,N_3964);
nor U4412 (N_4412,N_4041,N_3829);
xnor U4413 (N_4413,N_3925,N_3883);
nor U4414 (N_4414,N_3615,N_3991);
nand U4415 (N_4415,N_4087,N_4149);
xor U4416 (N_4416,N_4182,N_3986);
nand U4417 (N_4417,N_3630,N_4138);
nand U4418 (N_4418,N_4011,N_4069);
or U4419 (N_4419,N_3660,N_4066);
or U4420 (N_4420,N_3994,N_3882);
nand U4421 (N_4421,N_4075,N_3673);
or U4422 (N_4422,N_3949,N_3803);
nor U4423 (N_4423,N_4033,N_3843);
nand U4424 (N_4424,N_4169,N_3973);
nor U4425 (N_4425,N_3908,N_3830);
or U4426 (N_4426,N_3779,N_3945);
nor U4427 (N_4427,N_4083,N_3960);
or U4428 (N_4428,N_3963,N_3650);
nor U4429 (N_4429,N_4057,N_3817);
and U4430 (N_4430,N_3754,N_4006);
nand U4431 (N_4431,N_3726,N_3966);
nor U4432 (N_4432,N_3913,N_3688);
xnor U4433 (N_4433,N_3799,N_3641);
nand U4434 (N_4434,N_4115,N_4136);
nand U4435 (N_4435,N_3702,N_3895);
nor U4436 (N_4436,N_3655,N_3705);
and U4437 (N_4437,N_3866,N_4163);
nor U4438 (N_4438,N_4018,N_4155);
nand U4439 (N_4439,N_3814,N_3979);
xor U4440 (N_4440,N_3629,N_4010);
xor U4441 (N_4441,N_3853,N_4023);
xnor U4442 (N_4442,N_3894,N_4181);
xnor U4443 (N_4443,N_4092,N_4144);
and U4444 (N_4444,N_3697,N_3898);
nand U4445 (N_4445,N_4193,N_3820);
and U4446 (N_4446,N_3765,N_4065);
xor U4447 (N_4447,N_3698,N_4147);
or U4448 (N_4448,N_3602,N_3924);
xnor U4449 (N_4449,N_3663,N_3952);
or U4450 (N_4450,N_4151,N_3870);
nor U4451 (N_4451,N_3784,N_3769);
xor U4452 (N_4452,N_4089,N_3738);
nor U4453 (N_4453,N_3649,N_4189);
and U4454 (N_4454,N_3854,N_4123);
nand U4455 (N_4455,N_3609,N_3734);
nand U4456 (N_4456,N_3636,N_3825);
and U4457 (N_4457,N_3899,N_4168);
and U4458 (N_4458,N_3975,N_3606);
nor U4459 (N_4459,N_3868,N_3902);
nor U4460 (N_4460,N_4077,N_3714);
nor U4461 (N_4461,N_4028,N_3725);
or U4462 (N_4462,N_4160,N_3951);
or U4463 (N_4463,N_3873,N_3617);
and U4464 (N_4464,N_4095,N_3822);
nor U4465 (N_4465,N_3670,N_3981);
or U4466 (N_4466,N_4008,N_4032);
nand U4467 (N_4467,N_3627,N_4191);
nor U4468 (N_4468,N_4073,N_3903);
xor U4469 (N_4469,N_3875,N_4185);
or U4470 (N_4470,N_3801,N_4118);
nand U4471 (N_4471,N_3671,N_3819);
nand U4472 (N_4472,N_4084,N_4173);
nor U4473 (N_4473,N_4086,N_3604);
nor U4474 (N_4474,N_4186,N_3771);
or U4475 (N_4475,N_3832,N_4068);
and U4476 (N_4476,N_3826,N_3869);
and U4477 (N_4477,N_3806,N_4021);
xor U4478 (N_4478,N_3833,N_3798);
nand U4479 (N_4479,N_4019,N_4162);
xor U4480 (N_4480,N_3889,N_3936);
nand U4481 (N_4481,N_3778,N_3693);
nor U4482 (N_4482,N_4026,N_3786);
and U4483 (N_4483,N_3880,N_3939);
and U4484 (N_4484,N_3700,N_3813);
nand U4485 (N_4485,N_4062,N_3851);
nand U4486 (N_4486,N_4058,N_3614);
nand U4487 (N_4487,N_4038,N_3654);
nor U4488 (N_4488,N_3885,N_3618);
and U4489 (N_4489,N_3915,N_3621);
and U4490 (N_4490,N_3887,N_3647);
or U4491 (N_4491,N_4000,N_4171);
xnor U4492 (N_4492,N_3669,N_3919);
nor U4493 (N_4493,N_3607,N_4159);
or U4494 (N_4494,N_3752,N_3635);
and U4495 (N_4495,N_3748,N_4071);
and U4496 (N_4496,N_4013,N_4179);
or U4497 (N_4497,N_3807,N_3879);
or U4498 (N_4498,N_3920,N_3624);
nor U4499 (N_4499,N_3724,N_4079);
nor U4500 (N_4500,N_3998,N_4188);
nand U4501 (N_4501,N_3645,N_3924);
and U4502 (N_4502,N_3715,N_4064);
nor U4503 (N_4503,N_3924,N_3839);
and U4504 (N_4504,N_3816,N_3944);
nor U4505 (N_4505,N_3602,N_3793);
nor U4506 (N_4506,N_4058,N_3784);
nor U4507 (N_4507,N_3860,N_3752);
nor U4508 (N_4508,N_3853,N_3914);
xor U4509 (N_4509,N_3957,N_3712);
nand U4510 (N_4510,N_3806,N_3776);
nor U4511 (N_4511,N_4018,N_4154);
nand U4512 (N_4512,N_3889,N_3855);
xor U4513 (N_4513,N_4045,N_3945);
xnor U4514 (N_4514,N_3694,N_4107);
xor U4515 (N_4515,N_3971,N_3688);
nand U4516 (N_4516,N_3950,N_3883);
xor U4517 (N_4517,N_3962,N_3718);
or U4518 (N_4518,N_3766,N_3763);
and U4519 (N_4519,N_4058,N_4080);
nand U4520 (N_4520,N_3861,N_3941);
or U4521 (N_4521,N_3968,N_3724);
or U4522 (N_4522,N_3896,N_3761);
xor U4523 (N_4523,N_3829,N_3640);
nor U4524 (N_4524,N_3606,N_3786);
nand U4525 (N_4525,N_3708,N_4081);
xnor U4526 (N_4526,N_4159,N_3735);
or U4527 (N_4527,N_3668,N_3633);
xor U4528 (N_4528,N_3842,N_4042);
or U4529 (N_4529,N_3605,N_4103);
nand U4530 (N_4530,N_3763,N_3907);
nor U4531 (N_4531,N_4077,N_4059);
nor U4532 (N_4532,N_4071,N_4182);
nand U4533 (N_4533,N_4010,N_3950);
nand U4534 (N_4534,N_4172,N_3967);
xnor U4535 (N_4535,N_3718,N_3887);
and U4536 (N_4536,N_3959,N_4014);
nand U4537 (N_4537,N_3825,N_3720);
and U4538 (N_4538,N_4066,N_4164);
xnor U4539 (N_4539,N_3625,N_3792);
xor U4540 (N_4540,N_4011,N_3770);
or U4541 (N_4541,N_3611,N_3789);
nor U4542 (N_4542,N_3807,N_4136);
or U4543 (N_4543,N_3980,N_3746);
xor U4544 (N_4544,N_3871,N_3919);
nand U4545 (N_4545,N_3959,N_4107);
nor U4546 (N_4546,N_3845,N_4112);
xor U4547 (N_4547,N_3956,N_4011);
nor U4548 (N_4548,N_3723,N_3987);
xnor U4549 (N_4549,N_4019,N_3989);
or U4550 (N_4550,N_3616,N_3613);
and U4551 (N_4551,N_4008,N_3882);
xor U4552 (N_4552,N_4190,N_3858);
or U4553 (N_4553,N_3725,N_4102);
xnor U4554 (N_4554,N_3994,N_4043);
and U4555 (N_4555,N_3791,N_3663);
nor U4556 (N_4556,N_3852,N_4193);
nor U4557 (N_4557,N_3766,N_3730);
and U4558 (N_4558,N_4097,N_3698);
or U4559 (N_4559,N_4028,N_3651);
nand U4560 (N_4560,N_3795,N_3784);
and U4561 (N_4561,N_3826,N_3853);
or U4562 (N_4562,N_3826,N_4112);
nand U4563 (N_4563,N_4126,N_3646);
and U4564 (N_4564,N_4149,N_3989);
nand U4565 (N_4565,N_3647,N_3728);
nor U4566 (N_4566,N_3765,N_4005);
or U4567 (N_4567,N_3853,N_3877);
nand U4568 (N_4568,N_3631,N_3965);
xor U4569 (N_4569,N_3799,N_3947);
nor U4570 (N_4570,N_4080,N_4032);
nor U4571 (N_4571,N_4153,N_3986);
or U4572 (N_4572,N_3634,N_4092);
nand U4573 (N_4573,N_4149,N_4113);
xor U4574 (N_4574,N_3859,N_4141);
and U4575 (N_4575,N_3926,N_3657);
nand U4576 (N_4576,N_3792,N_3619);
or U4577 (N_4577,N_3842,N_3986);
or U4578 (N_4578,N_3756,N_3628);
nor U4579 (N_4579,N_3897,N_3635);
and U4580 (N_4580,N_3834,N_3970);
and U4581 (N_4581,N_4184,N_4198);
and U4582 (N_4582,N_3700,N_3856);
xor U4583 (N_4583,N_4061,N_3755);
or U4584 (N_4584,N_3856,N_3637);
and U4585 (N_4585,N_4026,N_3728);
nor U4586 (N_4586,N_3985,N_3870);
nor U4587 (N_4587,N_4021,N_3685);
nand U4588 (N_4588,N_3603,N_3700);
nand U4589 (N_4589,N_4030,N_3632);
or U4590 (N_4590,N_3895,N_3973);
or U4591 (N_4591,N_4013,N_3723);
nor U4592 (N_4592,N_3917,N_4164);
nor U4593 (N_4593,N_3809,N_4087);
xor U4594 (N_4594,N_3948,N_3671);
and U4595 (N_4595,N_4188,N_3746);
or U4596 (N_4596,N_3971,N_4087);
xor U4597 (N_4597,N_4107,N_3829);
or U4598 (N_4598,N_4037,N_3984);
or U4599 (N_4599,N_4131,N_4178);
and U4600 (N_4600,N_4040,N_3855);
nor U4601 (N_4601,N_4119,N_3889);
nand U4602 (N_4602,N_4176,N_3656);
xnor U4603 (N_4603,N_3839,N_3901);
or U4604 (N_4604,N_4045,N_3768);
nand U4605 (N_4605,N_4157,N_3630);
nor U4606 (N_4606,N_3731,N_4124);
nor U4607 (N_4607,N_4042,N_3811);
or U4608 (N_4608,N_4196,N_3777);
nand U4609 (N_4609,N_3736,N_4097);
xor U4610 (N_4610,N_3704,N_3868);
nor U4611 (N_4611,N_3783,N_3640);
nand U4612 (N_4612,N_3809,N_3910);
or U4613 (N_4613,N_3851,N_4157);
xor U4614 (N_4614,N_3792,N_3637);
nor U4615 (N_4615,N_3756,N_4060);
nor U4616 (N_4616,N_3725,N_4059);
or U4617 (N_4617,N_3825,N_4006);
xnor U4618 (N_4618,N_4162,N_3983);
nor U4619 (N_4619,N_3726,N_4049);
xor U4620 (N_4620,N_3615,N_3933);
and U4621 (N_4621,N_4074,N_3734);
xnor U4622 (N_4622,N_4180,N_4008);
and U4623 (N_4623,N_4193,N_3935);
or U4624 (N_4624,N_3767,N_3973);
xnor U4625 (N_4625,N_4186,N_4162);
nand U4626 (N_4626,N_4161,N_3976);
xnor U4627 (N_4627,N_4083,N_3959);
and U4628 (N_4628,N_3621,N_3946);
or U4629 (N_4629,N_3742,N_4062);
nand U4630 (N_4630,N_4144,N_3872);
nor U4631 (N_4631,N_3863,N_3620);
nand U4632 (N_4632,N_3752,N_3977);
nand U4633 (N_4633,N_4046,N_3690);
nor U4634 (N_4634,N_4000,N_3906);
and U4635 (N_4635,N_3750,N_3681);
or U4636 (N_4636,N_4002,N_4128);
xor U4637 (N_4637,N_3999,N_3655);
nand U4638 (N_4638,N_3847,N_4038);
nand U4639 (N_4639,N_3614,N_4148);
nor U4640 (N_4640,N_4117,N_3917);
and U4641 (N_4641,N_3623,N_3694);
nand U4642 (N_4642,N_4101,N_4090);
nand U4643 (N_4643,N_3824,N_3941);
or U4644 (N_4644,N_3605,N_3800);
xnor U4645 (N_4645,N_4023,N_4095);
and U4646 (N_4646,N_3959,N_3894);
nand U4647 (N_4647,N_3886,N_3818);
or U4648 (N_4648,N_3706,N_4111);
nand U4649 (N_4649,N_3967,N_4106);
or U4650 (N_4650,N_4068,N_4044);
and U4651 (N_4651,N_4014,N_4174);
and U4652 (N_4652,N_3662,N_4077);
and U4653 (N_4653,N_4161,N_4147);
nor U4654 (N_4654,N_4156,N_3854);
nor U4655 (N_4655,N_3703,N_4053);
xor U4656 (N_4656,N_4153,N_3806);
or U4657 (N_4657,N_4191,N_3684);
or U4658 (N_4658,N_3872,N_3830);
nor U4659 (N_4659,N_3989,N_3938);
or U4660 (N_4660,N_4167,N_3887);
nor U4661 (N_4661,N_3672,N_3704);
xor U4662 (N_4662,N_3896,N_4151);
nand U4663 (N_4663,N_3927,N_4047);
nor U4664 (N_4664,N_4107,N_4181);
nor U4665 (N_4665,N_3785,N_4097);
and U4666 (N_4666,N_3805,N_3982);
or U4667 (N_4667,N_3645,N_3904);
xnor U4668 (N_4668,N_3683,N_3785);
or U4669 (N_4669,N_3602,N_3791);
nor U4670 (N_4670,N_4162,N_3779);
nand U4671 (N_4671,N_4111,N_4042);
nor U4672 (N_4672,N_3999,N_3689);
and U4673 (N_4673,N_3962,N_3866);
xnor U4674 (N_4674,N_3904,N_4016);
xor U4675 (N_4675,N_3755,N_3629);
and U4676 (N_4676,N_3638,N_3908);
and U4677 (N_4677,N_3979,N_3699);
xnor U4678 (N_4678,N_3817,N_3847);
nor U4679 (N_4679,N_3771,N_3710);
xnor U4680 (N_4680,N_4104,N_3616);
or U4681 (N_4681,N_4198,N_3873);
xor U4682 (N_4682,N_4010,N_3680);
nand U4683 (N_4683,N_3824,N_4133);
nor U4684 (N_4684,N_3782,N_3892);
and U4685 (N_4685,N_3673,N_3627);
xor U4686 (N_4686,N_4162,N_4166);
and U4687 (N_4687,N_3960,N_4157);
nor U4688 (N_4688,N_3844,N_3939);
and U4689 (N_4689,N_3654,N_3687);
nor U4690 (N_4690,N_3614,N_3752);
nand U4691 (N_4691,N_4131,N_3615);
nor U4692 (N_4692,N_3875,N_3602);
and U4693 (N_4693,N_4107,N_3673);
or U4694 (N_4694,N_4182,N_3847);
or U4695 (N_4695,N_4118,N_3604);
nor U4696 (N_4696,N_4053,N_3904);
nor U4697 (N_4697,N_3939,N_3617);
and U4698 (N_4698,N_3853,N_3712);
nor U4699 (N_4699,N_3974,N_3765);
nor U4700 (N_4700,N_4143,N_3970);
and U4701 (N_4701,N_3740,N_3705);
and U4702 (N_4702,N_3812,N_4132);
and U4703 (N_4703,N_4082,N_3948);
nand U4704 (N_4704,N_3970,N_4041);
or U4705 (N_4705,N_3858,N_3928);
nor U4706 (N_4706,N_3615,N_3856);
nor U4707 (N_4707,N_3733,N_3947);
nor U4708 (N_4708,N_3929,N_3635);
or U4709 (N_4709,N_3794,N_3625);
xor U4710 (N_4710,N_3663,N_3762);
and U4711 (N_4711,N_3646,N_4042);
and U4712 (N_4712,N_3714,N_3661);
and U4713 (N_4713,N_4127,N_4135);
or U4714 (N_4714,N_3619,N_4062);
or U4715 (N_4715,N_3626,N_3864);
xor U4716 (N_4716,N_4170,N_4126);
nand U4717 (N_4717,N_3831,N_3992);
and U4718 (N_4718,N_3753,N_4055);
xnor U4719 (N_4719,N_3647,N_3964);
nand U4720 (N_4720,N_4145,N_3643);
nand U4721 (N_4721,N_4115,N_4085);
or U4722 (N_4722,N_4114,N_3891);
and U4723 (N_4723,N_4183,N_3778);
xor U4724 (N_4724,N_4143,N_4080);
nand U4725 (N_4725,N_4159,N_4074);
and U4726 (N_4726,N_3725,N_3638);
and U4727 (N_4727,N_3949,N_3942);
or U4728 (N_4728,N_3752,N_3692);
and U4729 (N_4729,N_4144,N_3804);
nand U4730 (N_4730,N_3947,N_3705);
or U4731 (N_4731,N_3694,N_3933);
and U4732 (N_4732,N_3699,N_3871);
or U4733 (N_4733,N_4060,N_3896);
and U4734 (N_4734,N_3611,N_3705);
and U4735 (N_4735,N_4028,N_3911);
nand U4736 (N_4736,N_3620,N_3655);
nor U4737 (N_4737,N_4131,N_3626);
nor U4738 (N_4738,N_3866,N_3773);
nor U4739 (N_4739,N_3655,N_3755);
nor U4740 (N_4740,N_3702,N_3869);
xor U4741 (N_4741,N_4140,N_4166);
and U4742 (N_4742,N_3620,N_3646);
nor U4743 (N_4743,N_4183,N_4142);
nand U4744 (N_4744,N_3982,N_3811);
xor U4745 (N_4745,N_3837,N_3758);
nor U4746 (N_4746,N_3850,N_3863);
nand U4747 (N_4747,N_4084,N_3749);
nor U4748 (N_4748,N_4169,N_3872);
nand U4749 (N_4749,N_3921,N_3752);
and U4750 (N_4750,N_3953,N_3910);
and U4751 (N_4751,N_4095,N_4064);
xor U4752 (N_4752,N_3836,N_3691);
and U4753 (N_4753,N_3807,N_4139);
xnor U4754 (N_4754,N_4144,N_3849);
or U4755 (N_4755,N_3791,N_3960);
xor U4756 (N_4756,N_3981,N_3692);
xnor U4757 (N_4757,N_3838,N_4067);
or U4758 (N_4758,N_3668,N_3979);
or U4759 (N_4759,N_3654,N_3993);
nor U4760 (N_4760,N_3809,N_3691);
xnor U4761 (N_4761,N_3932,N_4146);
nand U4762 (N_4762,N_3994,N_3975);
or U4763 (N_4763,N_3659,N_3955);
nand U4764 (N_4764,N_3720,N_3832);
and U4765 (N_4765,N_3789,N_3927);
xnor U4766 (N_4766,N_3922,N_4150);
and U4767 (N_4767,N_4090,N_3796);
or U4768 (N_4768,N_3615,N_4142);
xor U4769 (N_4769,N_3777,N_4126);
or U4770 (N_4770,N_3932,N_4047);
or U4771 (N_4771,N_3770,N_4080);
or U4772 (N_4772,N_4182,N_3837);
and U4773 (N_4773,N_3946,N_3913);
xor U4774 (N_4774,N_3700,N_4050);
nor U4775 (N_4775,N_3930,N_4096);
xnor U4776 (N_4776,N_4047,N_3936);
or U4777 (N_4777,N_4134,N_3769);
xor U4778 (N_4778,N_4111,N_4134);
or U4779 (N_4779,N_4138,N_3647);
nor U4780 (N_4780,N_4123,N_3956);
nor U4781 (N_4781,N_3697,N_3872);
xnor U4782 (N_4782,N_3702,N_4067);
xnor U4783 (N_4783,N_3805,N_4106);
and U4784 (N_4784,N_3782,N_3714);
xor U4785 (N_4785,N_4184,N_3732);
and U4786 (N_4786,N_3954,N_4005);
and U4787 (N_4787,N_4102,N_3839);
nor U4788 (N_4788,N_3804,N_4162);
nand U4789 (N_4789,N_3730,N_3885);
nor U4790 (N_4790,N_3778,N_3773);
xnor U4791 (N_4791,N_4111,N_3645);
xnor U4792 (N_4792,N_4143,N_3636);
and U4793 (N_4793,N_4053,N_4199);
nor U4794 (N_4794,N_4152,N_3793);
xor U4795 (N_4795,N_3720,N_4140);
and U4796 (N_4796,N_3640,N_3995);
and U4797 (N_4797,N_4139,N_3808);
or U4798 (N_4798,N_4011,N_4186);
or U4799 (N_4799,N_3978,N_3818);
xor U4800 (N_4800,N_4734,N_4375);
xor U4801 (N_4801,N_4264,N_4775);
nand U4802 (N_4802,N_4787,N_4533);
nand U4803 (N_4803,N_4571,N_4242);
nand U4804 (N_4804,N_4629,N_4667);
nor U4805 (N_4805,N_4245,N_4272);
nor U4806 (N_4806,N_4500,N_4753);
xor U4807 (N_4807,N_4411,N_4399);
nor U4808 (N_4808,N_4423,N_4436);
or U4809 (N_4809,N_4593,N_4567);
nand U4810 (N_4810,N_4613,N_4581);
and U4811 (N_4811,N_4679,N_4605);
nor U4812 (N_4812,N_4281,N_4678);
xnor U4813 (N_4813,N_4204,N_4381);
xor U4814 (N_4814,N_4441,N_4530);
nor U4815 (N_4815,N_4582,N_4284);
nor U4816 (N_4816,N_4563,N_4603);
or U4817 (N_4817,N_4365,N_4614);
nor U4818 (N_4818,N_4637,N_4633);
xnor U4819 (N_4819,N_4665,N_4287);
and U4820 (N_4820,N_4539,N_4340);
nor U4821 (N_4821,N_4774,N_4231);
xor U4822 (N_4822,N_4451,N_4797);
or U4823 (N_4823,N_4414,N_4564);
nor U4824 (N_4824,N_4244,N_4410);
nand U4825 (N_4825,N_4290,N_4486);
nand U4826 (N_4826,N_4298,N_4367);
or U4827 (N_4827,N_4764,N_4599);
and U4828 (N_4828,N_4219,N_4396);
nand U4829 (N_4829,N_4417,N_4624);
and U4830 (N_4830,N_4589,N_4235);
nor U4831 (N_4831,N_4346,N_4283);
and U4832 (N_4832,N_4526,N_4454);
nand U4833 (N_4833,N_4241,N_4523);
or U4834 (N_4834,N_4368,N_4370);
xnor U4835 (N_4835,N_4401,N_4543);
xor U4836 (N_4836,N_4202,N_4675);
and U4837 (N_4837,N_4345,N_4583);
and U4838 (N_4838,N_4259,N_4700);
nor U4839 (N_4839,N_4542,N_4519);
or U4840 (N_4840,N_4507,N_4262);
nor U4841 (N_4841,N_4630,N_4650);
nor U4842 (N_4842,N_4501,N_4251);
xor U4843 (N_4843,N_4254,N_4329);
and U4844 (N_4844,N_4600,N_4347);
and U4845 (N_4845,N_4587,N_4333);
xor U4846 (N_4846,N_4331,N_4225);
nor U4847 (N_4847,N_4766,N_4521);
nor U4848 (N_4848,N_4409,N_4322);
nand U4849 (N_4849,N_4491,N_4769);
and U4850 (N_4850,N_4692,N_4348);
or U4851 (N_4851,N_4361,N_4209);
and U4852 (N_4852,N_4779,N_4560);
nor U4853 (N_4853,N_4460,N_4795);
nor U4854 (N_4854,N_4724,N_4555);
and U4855 (N_4855,N_4529,N_4458);
nor U4856 (N_4856,N_4383,N_4655);
and U4857 (N_4857,N_4404,N_4638);
or U4858 (N_4858,N_4738,N_4471);
and U4859 (N_4859,N_4301,N_4658);
and U4860 (N_4860,N_4377,N_4628);
xnor U4861 (N_4861,N_4720,N_4391);
xor U4862 (N_4862,N_4336,N_4573);
and U4863 (N_4863,N_4598,N_4360);
nand U4864 (N_4864,N_4757,N_4308);
nand U4865 (N_4865,N_4550,N_4577);
nand U4866 (N_4866,N_4709,N_4228);
nand U4867 (N_4867,N_4611,N_4395);
xor U4868 (N_4868,N_4747,N_4479);
nor U4869 (N_4869,N_4648,N_4594);
and U4870 (N_4870,N_4495,N_4371);
nand U4871 (N_4871,N_4698,N_4349);
nand U4872 (N_4872,N_4616,N_4615);
xor U4873 (N_4873,N_4783,N_4554);
nor U4874 (N_4874,N_4776,N_4540);
xor U4875 (N_4875,N_4403,N_4740);
nand U4876 (N_4876,N_4496,N_4296);
nand U4877 (N_4877,N_4325,N_4257);
xnor U4878 (N_4878,N_4444,N_4269);
nor U4879 (N_4879,N_4355,N_4492);
or U4880 (N_4880,N_4392,N_4278);
or U4881 (N_4881,N_4666,N_4626);
nor U4882 (N_4882,N_4211,N_4768);
nand U4883 (N_4883,N_4545,N_4697);
or U4884 (N_4884,N_4440,N_4236);
nand U4885 (N_4885,N_4645,N_4223);
and U4886 (N_4886,N_4758,N_4681);
nand U4887 (N_4887,N_4782,N_4721);
or U4888 (N_4888,N_4565,N_4247);
xor U4889 (N_4889,N_4473,N_4708);
nand U4890 (N_4890,N_4536,N_4310);
xor U4891 (N_4891,N_4464,N_4690);
nor U4892 (N_4892,N_4636,N_4323);
or U4893 (N_4893,N_4732,N_4684);
or U4894 (N_4894,N_4785,N_4644);
nor U4895 (N_4895,N_4482,N_4651);
xor U4896 (N_4896,N_4380,N_4514);
or U4897 (N_4897,N_4618,N_4229);
nand U4898 (N_4898,N_4386,N_4256);
nand U4899 (N_4899,N_4435,N_4452);
nor U4900 (N_4900,N_4745,N_4227);
and U4901 (N_4901,N_4232,N_4270);
and U4902 (N_4902,N_4639,N_4237);
and U4903 (N_4903,N_4670,N_4457);
nand U4904 (N_4904,N_4448,N_4341);
xor U4905 (N_4905,N_4233,N_4557);
nand U4906 (N_4906,N_4796,N_4799);
or U4907 (N_4907,N_4522,N_4316);
nand U4908 (N_4908,N_4297,N_4574);
xor U4909 (N_4909,N_4499,N_4206);
and U4910 (N_4910,N_4324,N_4652);
nand U4911 (N_4911,N_4389,N_4788);
and U4912 (N_4912,N_4714,N_4427);
and U4913 (N_4913,N_4311,N_4596);
nor U4914 (N_4914,N_4777,N_4425);
or U4915 (N_4915,N_4754,N_4713);
xnor U4916 (N_4916,N_4718,N_4489);
nand U4917 (N_4917,N_4749,N_4561);
nor U4918 (N_4918,N_4252,N_4673);
nand U4919 (N_4919,N_4504,N_4619);
and U4920 (N_4920,N_4717,N_4685);
nor U4921 (N_4921,N_4216,N_4218);
or U4922 (N_4922,N_4657,N_4729);
nor U4923 (N_4923,N_4369,N_4248);
nor U4924 (N_4924,N_4664,N_4663);
nor U4925 (N_4925,N_4275,N_4748);
xor U4926 (N_4926,N_4602,N_4344);
nand U4927 (N_4927,N_4765,N_4627);
nor U4928 (N_4928,N_4695,N_4510);
and U4929 (N_4929,N_4334,N_4511);
nand U4930 (N_4930,N_4789,N_4699);
nand U4931 (N_4931,N_4798,N_4632);
or U4932 (N_4932,N_4366,N_4794);
nor U4933 (N_4933,N_4453,N_4541);
nor U4934 (N_4934,N_4544,N_4622);
nor U4935 (N_4935,N_4570,N_4635);
nor U4936 (N_4936,N_4439,N_4601);
xor U4937 (N_4937,N_4537,N_4730);
nand U4938 (N_4938,N_4586,N_4413);
xnor U4939 (N_4939,N_4480,N_4475);
and U4940 (N_4940,N_4559,N_4295);
nand U4941 (N_4941,N_4286,N_4226);
and U4942 (N_4942,N_4741,N_4552);
xnor U4943 (N_4943,N_4442,N_4406);
and U4944 (N_4944,N_4688,N_4761);
and U4945 (N_4945,N_4304,N_4481);
xor U4946 (N_4946,N_4736,N_4320);
xor U4947 (N_4947,N_4597,N_4327);
nor U4948 (N_4948,N_4398,N_4750);
nor U4949 (N_4949,N_4277,N_4470);
nor U4950 (N_4950,N_4659,N_4502);
or U4951 (N_4951,N_4512,N_4609);
nor U4952 (N_4952,N_4646,N_4474);
nor U4953 (N_4953,N_4640,N_4434);
xnor U4954 (N_4954,N_4465,N_4484);
xnor U4955 (N_4955,N_4727,N_4677);
xor U4956 (N_4956,N_4584,N_4483);
nor U4957 (N_4957,N_4781,N_4300);
nand U4958 (N_4958,N_4548,N_4494);
nand U4959 (N_4959,N_4531,N_4437);
nand U4960 (N_4960,N_4590,N_4315);
nand U4961 (N_4961,N_4362,N_4686);
and U4962 (N_4962,N_4210,N_4641);
xor U4963 (N_4963,N_4691,N_4469);
nand U4964 (N_4964,N_4430,N_4382);
nand U4965 (N_4965,N_4706,N_4566);
nor U4966 (N_4966,N_4505,N_4710);
and U4967 (N_4967,N_4438,N_4466);
nand U4968 (N_4968,N_4488,N_4289);
xor U4969 (N_4969,N_4595,N_4656);
nand U4970 (N_4970,N_4468,N_4607);
or U4971 (N_4971,N_4513,N_4220);
xnor U4972 (N_4972,N_4379,N_4671);
nor U4973 (N_4973,N_4532,N_4402);
or U4974 (N_4974,N_4342,N_4535);
and U4975 (N_4975,N_4472,N_4255);
nand U4976 (N_4976,N_4376,N_4591);
nand U4977 (N_4977,N_4756,N_4549);
nor U4978 (N_4978,N_4224,N_4763);
nand U4979 (N_4979,N_4378,N_4508);
xnor U4980 (N_4980,N_4767,N_4354);
nand U4981 (N_4981,N_4580,N_4445);
or U4982 (N_4982,N_4373,N_4343);
or U4983 (N_4983,N_4770,N_4653);
and U4984 (N_4984,N_4213,N_4265);
xnor U4985 (N_4985,N_4604,N_4267);
xnor U4986 (N_4986,N_4722,N_4551);
or U4987 (N_4987,N_4707,N_4762);
nand U4988 (N_4988,N_4556,N_4705);
and U4989 (N_4989,N_4791,N_4205);
and U4990 (N_4990,N_4493,N_4447);
nor U4991 (N_4991,N_4517,N_4680);
nor U4992 (N_4992,N_4528,N_4385);
nand U4993 (N_4993,N_4222,N_4352);
nor U4994 (N_4994,N_4631,N_4271);
nand U4995 (N_4995,N_4412,N_4498);
nor U4996 (N_4996,N_4372,N_4234);
xnor U4997 (N_4997,N_4728,N_4478);
nand U4998 (N_4998,N_4203,N_4759);
nand U4999 (N_4999,N_4357,N_4485);
nor U5000 (N_5000,N_4506,N_4520);
or U5001 (N_5001,N_4703,N_4608);
or U5002 (N_5002,N_4291,N_4249);
xor U5003 (N_5003,N_4433,N_4418);
xnor U5004 (N_5004,N_4456,N_4790);
nor U5005 (N_5005,N_4294,N_4682);
or U5006 (N_5006,N_4746,N_4778);
xor U5007 (N_5007,N_4702,N_4687);
and U5008 (N_5008,N_4588,N_4674);
nand U5009 (N_5009,N_4649,N_4742);
nand U5010 (N_5010,N_4612,N_4450);
or U5011 (N_5011,N_4459,N_4303);
nor U5012 (N_5012,N_4317,N_4527);
xnor U5013 (N_5013,N_4731,N_4585);
nand U5014 (N_5014,N_4306,N_4704);
xor U5015 (N_5015,N_4246,N_4328);
and U5016 (N_5016,N_4643,N_4363);
nand U5017 (N_5017,N_4693,N_4351);
nand U5018 (N_5018,N_4307,N_4250);
or U5019 (N_5019,N_4752,N_4288);
nor U5020 (N_5020,N_4339,N_4208);
nor U5021 (N_5021,N_4200,N_4230);
nand U5022 (N_5022,N_4515,N_4476);
nor U5023 (N_5023,N_4621,N_4715);
or U5024 (N_5024,N_4592,N_4518);
and U5025 (N_5025,N_4302,N_4672);
nand U5026 (N_5026,N_4268,N_4719);
nand U5027 (N_5027,N_4792,N_4266);
or U5028 (N_5028,N_4394,N_4579);
nor U5029 (N_5029,N_4538,N_4274);
or U5030 (N_5030,N_4516,N_4712);
xnor U5031 (N_5031,N_4524,N_4725);
nor U5032 (N_5032,N_4420,N_4422);
or U5033 (N_5033,N_4280,N_4553);
or U5034 (N_5034,N_4562,N_4558);
or U5035 (N_5035,N_4276,N_4771);
nand U5036 (N_5036,N_4497,N_4625);
xor U5037 (N_5037,N_4617,N_4487);
and U5038 (N_5038,N_4669,N_4760);
nand U5039 (N_5039,N_4773,N_4668);
nor U5040 (N_5040,N_4575,N_4258);
nor U5041 (N_5041,N_4694,N_4353);
xor U5042 (N_5042,N_4477,N_4240);
and U5043 (N_5043,N_4337,N_4314);
xnor U5044 (N_5044,N_4578,N_4490);
nand U5045 (N_5045,N_4534,N_4739);
and U5046 (N_5046,N_4647,N_4689);
or U5047 (N_5047,N_4282,N_4569);
or U5048 (N_5048,N_4426,N_4330);
xnor U5049 (N_5049,N_4285,N_4390);
nand U5050 (N_5050,N_4784,N_4321);
and U5051 (N_5051,N_4356,N_4733);
xnor U5052 (N_5052,N_4239,N_4620);
nor U5053 (N_5053,N_4431,N_4547);
xnor U5054 (N_5054,N_4429,N_4201);
nand U5055 (N_5055,N_4509,N_4318);
and U5056 (N_5056,N_4503,N_4623);
nand U5057 (N_5057,N_4326,N_4743);
nor U5058 (N_5058,N_4467,N_4716);
or U5059 (N_5059,N_4207,N_4662);
or U5060 (N_5060,N_4393,N_4546);
nor U5061 (N_5061,N_4217,N_4463);
nand U5062 (N_5062,N_4292,N_4374);
nand U5063 (N_5063,N_4455,N_4735);
xnor U5064 (N_5064,N_4263,N_4572);
xnor U5065 (N_5065,N_4408,N_4260);
and U5066 (N_5066,N_4568,N_4221);
and U5067 (N_5067,N_4273,N_4384);
xor U5068 (N_5068,N_4421,N_4786);
xnor U5069 (N_5069,N_4751,N_4335);
nor U5070 (N_5070,N_4446,N_4683);
nand U5071 (N_5071,N_4388,N_4364);
and U5072 (N_5072,N_4755,N_4212);
and U5073 (N_5073,N_4701,N_4238);
nor U5074 (N_5074,N_4793,N_4696);
or U5075 (N_5075,N_4305,N_4660);
nand U5076 (N_5076,N_4654,N_4424);
xor U5077 (N_5077,N_4215,N_4279);
or U5078 (N_5078,N_4780,N_4243);
nand U5079 (N_5079,N_4634,N_4711);
or U5080 (N_5080,N_4359,N_4350);
or U5081 (N_5081,N_4610,N_4419);
nand U5082 (N_5082,N_4415,N_4214);
nor U5083 (N_5083,N_4407,N_4358);
nor U5084 (N_5084,N_4606,N_4443);
or U5085 (N_5085,N_4676,N_4400);
nand U5086 (N_5086,N_4309,N_4293);
xor U5087 (N_5087,N_4299,N_4461);
and U5088 (N_5088,N_4405,N_4416);
nor U5089 (N_5089,N_4723,N_4462);
or U5090 (N_5090,N_4428,N_4661);
nor U5091 (N_5091,N_4726,N_4319);
xnor U5092 (N_5092,N_4432,N_4772);
or U5093 (N_5093,N_4744,N_4332);
nor U5094 (N_5094,N_4397,N_4338);
nor U5095 (N_5095,N_4525,N_4642);
nand U5096 (N_5096,N_4261,N_4576);
xnor U5097 (N_5097,N_4387,N_4737);
xnor U5098 (N_5098,N_4449,N_4312);
nor U5099 (N_5099,N_4313,N_4253);
xor U5100 (N_5100,N_4519,N_4426);
nand U5101 (N_5101,N_4489,N_4394);
and U5102 (N_5102,N_4527,N_4227);
nand U5103 (N_5103,N_4636,N_4392);
nand U5104 (N_5104,N_4629,N_4263);
xor U5105 (N_5105,N_4272,N_4641);
nor U5106 (N_5106,N_4474,N_4542);
xnor U5107 (N_5107,N_4282,N_4217);
nor U5108 (N_5108,N_4724,N_4275);
and U5109 (N_5109,N_4399,N_4381);
or U5110 (N_5110,N_4228,N_4501);
and U5111 (N_5111,N_4373,N_4307);
nor U5112 (N_5112,N_4380,N_4617);
xnor U5113 (N_5113,N_4612,N_4202);
or U5114 (N_5114,N_4401,N_4459);
or U5115 (N_5115,N_4628,N_4584);
xnor U5116 (N_5116,N_4362,N_4215);
nor U5117 (N_5117,N_4508,N_4617);
nand U5118 (N_5118,N_4778,N_4306);
nand U5119 (N_5119,N_4293,N_4725);
nor U5120 (N_5120,N_4678,N_4788);
or U5121 (N_5121,N_4690,N_4631);
nand U5122 (N_5122,N_4481,N_4490);
and U5123 (N_5123,N_4493,N_4617);
or U5124 (N_5124,N_4513,N_4542);
xor U5125 (N_5125,N_4623,N_4681);
xor U5126 (N_5126,N_4572,N_4482);
xnor U5127 (N_5127,N_4244,N_4694);
nor U5128 (N_5128,N_4204,N_4425);
and U5129 (N_5129,N_4490,N_4581);
xor U5130 (N_5130,N_4677,N_4365);
nand U5131 (N_5131,N_4267,N_4254);
nand U5132 (N_5132,N_4788,N_4533);
xor U5133 (N_5133,N_4620,N_4397);
or U5134 (N_5134,N_4713,N_4702);
xnor U5135 (N_5135,N_4515,N_4523);
or U5136 (N_5136,N_4390,N_4467);
and U5137 (N_5137,N_4491,N_4571);
nor U5138 (N_5138,N_4282,N_4664);
xor U5139 (N_5139,N_4222,N_4216);
xor U5140 (N_5140,N_4662,N_4231);
nand U5141 (N_5141,N_4625,N_4558);
nand U5142 (N_5142,N_4374,N_4620);
nor U5143 (N_5143,N_4462,N_4642);
or U5144 (N_5144,N_4281,N_4716);
and U5145 (N_5145,N_4797,N_4754);
nand U5146 (N_5146,N_4370,N_4594);
and U5147 (N_5147,N_4425,N_4592);
xor U5148 (N_5148,N_4565,N_4725);
or U5149 (N_5149,N_4669,N_4218);
xnor U5150 (N_5150,N_4580,N_4794);
or U5151 (N_5151,N_4782,N_4538);
and U5152 (N_5152,N_4799,N_4709);
or U5153 (N_5153,N_4600,N_4648);
nand U5154 (N_5154,N_4598,N_4541);
nand U5155 (N_5155,N_4675,N_4557);
or U5156 (N_5156,N_4201,N_4254);
or U5157 (N_5157,N_4561,N_4299);
nand U5158 (N_5158,N_4202,N_4574);
nand U5159 (N_5159,N_4766,N_4604);
nor U5160 (N_5160,N_4331,N_4597);
nor U5161 (N_5161,N_4278,N_4433);
nand U5162 (N_5162,N_4302,N_4594);
and U5163 (N_5163,N_4508,N_4779);
and U5164 (N_5164,N_4698,N_4567);
and U5165 (N_5165,N_4329,N_4262);
xnor U5166 (N_5166,N_4465,N_4651);
nand U5167 (N_5167,N_4729,N_4668);
or U5168 (N_5168,N_4484,N_4435);
nor U5169 (N_5169,N_4664,N_4285);
and U5170 (N_5170,N_4299,N_4316);
nor U5171 (N_5171,N_4426,N_4447);
or U5172 (N_5172,N_4268,N_4273);
xor U5173 (N_5173,N_4706,N_4279);
and U5174 (N_5174,N_4637,N_4747);
or U5175 (N_5175,N_4430,N_4317);
nand U5176 (N_5176,N_4300,N_4758);
nor U5177 (N_5177,N_4224,N_4558);
nand U5178 (N_5178,N_4358,N_4775);
nor U5179 (N_5179,N_4437,N_4351);
or U5180 (N_5180,N_4339,N_4292);
nand U5181 (N_5181,N_4773,N_4562);
or U5182 (N_5182,N_4238,N_4778);
xor U5183 (N_5183,N_4241,N_4749);
nor U5184 (N_5184,N_4683,N_4298);
nand U5185 (N_5185,N_4365,N_4227);
and U5186 (N_5186,N_4226,N_4369);
and U5187 (N_5187,N_4260,N_4474);
or U5188 (N_5188,N_4552,N_4267);
nor U5189 (N_5189,N_4203,N_4760);
or U5190 (N_5190,N_4500,N_4443);
and U5191 (N_5191,N_4773,N_4786);
and U5192 (N_5192,N_4203,N_4618);
and U5193 (N_5193,N_4572,N_4664);
or U5194 (N_5194,N_4701,N_4713);
or U5195 (N_5195,N_4767,N_4713);
or U5196 (N_5196,N_4745,N_4463);
nor U5197 (N_5197,N_4746,N_4490);
or U5198 (N_5198,N_4584,N_4462);
or U5199 (N_5199,N_4305,N_4206);
and U5200 (N_5200,N_4223,N_4370);
or U5201 (N_5201,N_4360,N_4325);
nand U5202 (N_5202,N_4278,N_4320);
nand U5203 (N_5203,N_4255,N_4520);
nand U5204 (N_5204,N_4571,N_4655);
nand U5205 (N_5205,N_4275,N_4624);
or U5206 (N_5206,N_4424,N_4412);
nor U5207 (N_5207,N_4430,N_4692);
nand U5208 (N_5208,N_4646,N_4352);
or U5209 (N_5209,N_4663,N_4572);
and U5210 (N_5210,N_4462,N_4570);
nor U5211 (N_5211,N_4699,N_4726);
xnor U5212 (N_5212,N_4282,N_4426);
or U5213 (N_5213,N_4264,N_4787);
and U5214 (N_5214,N_4653,N_4643);
nand U5215 (N_5215,N_4762,N_4770);
nor U5216 (N_5216,N_4393,N_4504);
xor U5217 (N_5217,N_4350,N_4523);
nor U5218 (N_5218,N_4690,N_4405);
xnor U5219 (N_5219,N_4630,N_4573);
xor U5220 (N_5220,N_4433,N_4214);
xor U5221 (N_5221,N_4320,N_4494);
xnor U5222 (N_5222,N_4708,N_4678);
nor U5223 (N_5223,N_4762,N_4712);
nand U5224 (N_5224,N_4242,N_4440);
or U5225 (N_5225,N_4509,N_4240);
or U5226 (N_5226,N_4266,N_4525);
xor U5227 (N_5227,N_4325,N_4713);
nand U5228 (N_5228,N_4235,N_4397);
and U5229 (N_5229,N_4265,N_4379);
xor U5230 (N_5230,N_4526,N_4790);
and U5231 (N_5231,N_4385,N_4354);
nor U5232 (N_5232,N_4770,N_4776);
nand U5233 (N_5233,N_4375,N_4223);
nand U5234 (N_5234,N_4741,N_4229);
xnor U5235 (N_5235,N_4692,N_4771);
nor U5236 (N_5236,N_4648,N_4392);
xor U5237 (N_5237,N_4678,N_4316);
xor U5238 (N_5238,N_4259,N_4441);
nor U5239 (N_5239,N_4719,N_4678);
nand U5240 (N_5240,N_4664,N_4547);
nor U5241 (N_5241,N_4550,N_4480);
and U5242 (N_5242,N_4261,N_4302);
nor U5243 (N_5243,N_4789,N_4650);
nand U5244 (N_5244,N_4294,N_4775);
nor U5245 (N_5245,N_4506,N_4491);
and U5246 (N_5246,N_4448,N_4467);
or U5247 (N_5247,N_4279,N_4694);
xor U5248 (N_5248,N_4734,N_4755);
or U5249 (N_5249,N_4662,N_4376);
and U5250 (N_5250,N_4493,N_4646);
nand U5251 (N_5251,N_4543,N_4379);
nor U5252 (N_5252,N_4796,N_4533);
or U5253 (N_5253,N_4493,N_4254);
xnor U5254 (N_5254,N_4640,N_4611);
nand U5255 (N_5255,N_4552,N_4516);
or U5256 (N_5256,N_4580,N_4265);
nand U5257 (N_5257,N_4450,N_4513);
nor U5258 (N_5258,N_4448,N_4599);
nor U5259 (N_5259,N_4593,N_4210);
and U5260 (N_5260,N_4314,N_4523);
nand U5261 (N_5261,N_4718,N_4221);
xor U5262 (N_5262,N_4314,N_4386);
xnor U5263 (N_5263,N_4773,N_4493);
xnor U5264 (N_5264,N_4389,N_4507);
nor U5265 (N_5265,N_4376,N_4442);
or U5266 (N_5266,N_4547,N_4673);
or U5267 (N_5267,N_4669,N_4509);
nand U5268 (N_5268,N_4292,N_4512);
nor U5269 (N_5269,N_4727,N_4382);
xor U5270 (N_5270,N_4399,N_4748);
xor U5271 (N_5271,N_4702,N_4769);
nor U5272 (N_5272,N_4267,N_4583);
nor U5273 (N_5273,N_4731,N_4215);
nand U5274 (N_5274,N_4463,N_4698);
nor U5275 (N_5275,N_4254,N_4453);
or U5276 (N_5276,N_4741,N_4369);
xor U5277 (N_5277,N_4459,N_4426);
nand U5278 (N_5278,N_4318,N_4567);
xor U5279 (N_5279,N_4320,N_4479);
or U5280 (N_5280,N_4484,N_4326);
nand U5281 (N_5281,N_4749,N_4671);
and U5282 (N_5282,N_4514,N_4759);
nand U5283 (N_5283,N_4200,N_4343);
nand U5284 (N_5284,N_4677,N_4752);
nand U5285 (N_5285,N_4707,N_4678);
nand U5286 (N_5286,N_4418,N_4613);
nand U5287 (N_5287,N_4446,N_4212);
nand U5288 (N_5288,N_4607,N_4661);
and U5289 (N_5289,N_4749,N_4357);
or U5290 (N_5290,N_4734,N_4221);
or U5291 (N_5291,N_4342,N_4781);
nand U5292 (N_5292,N_4259,N_4616);
and U5293 (N_5293,N_4712,N_4778);
or U5294 (N_5294,N_4216,N_4485);
nor U5295 (N_5295,N_4744,N_4363);
nand U5296 (N_5296,N_4481,N_4517);
or U5297 (N_5297,N_4367,N_4215);
or U5298 (N_5298,N_4491,N_4702);
nor U5299 (N_5299,N_4657,N_4771);
xnor U5300 (N_5300,N_4776,N_4238);
nand U5301 (N_5301,N_4344,N_4354);
nand U5302 (N_5302,N_4768,N_4760);
or U5303 (N_5303,N_4314,N_4357);
nand U5304 (N_5304,N_4342,N_4557);
xnor U5305 (N_5305,N_4354,N_4498);
nor U5306 (N_5306,N_4236,N_4435);
nand U5307 (N_5307,N_4370,N_4744);
nand U5308 (N_5308,N_4713,N_4661);
and U5309 (N_5309,N_4422,N_4716);
or U5310 (N_5310,N_4636,N_4629);
nand U5311 (N_5311,N_4757,N_4272);
nor U5312 (N_5312,N_4466,N_4511);
and U5313 (N_5313,N_4723,N_4394);
xor U5314 (N_5314,N_4639,N_4556);
nand U5315 (N_5315,N_4360,N_4792);
and U5316 (N_5316,N_4547,N_4638);
xnor U5317 (N_5317,N_4617,N_4751);
or U5318 (N_5318,N_4626,N_4205);
xnor U5319 (N_5319,N_4501,N_4700);
nand U5320 (N_5320,N_4793,N_4227);
nand U5321 (N_5321,N_4308,N_4384);
and U5322 (N_5322,N_4309,N_4499);
nand U5323 (N_5323,N_4576,N_4792);
nor U5324 (N_5324,N_4497,N_4752);
or U5325 (N_5325,N_4672,N_4682);
or U5326 (N_5326,N_4229,N_4300);
xor U5327 (N_5327,N_4309,N_4506);
nor U5328 (N_5328,N_4405,N_4371);
nor U5329 (N_5329,N_4257,N_4387);
or U5330 (N_5330,N_4765,N_4331);
xor U5331 (N_5331,N_4539,N_4232);
nor U5332 (N_5332,N_4776,N_4404);
and U5333 (N_5333,N_4403,N_4330);
and U5334 (N_5334,N_4382,N_4664);
nand U5335 (N_5335,N_4746,N_4749);
nor U5336 (N_5336,N_4672,N_4745);
nand U5337 (N_5337,N_4499,N_4742);
nor U5338 (N_5338,N_4676,N_4458);
nor U5339 (N_5339,N_4383,N_4612);
nor U5340 (N_5340,N_4412,N_4530);
xor U5341 (N_5341,N_4747,N_4629);
xor U5342 (N_5342,N_4611,N_4465);
or U5343 (N_5343,N_4259,N_4591);
or U5344 (N_5344,N_4274,N_4672);
nand U5345 (N_5345,N_4765,N_4494);
or U5346 (N_5346,N_4504,N_4362);
nand U5347 (N_5347,N_4465,N_4299);
or U5348 (N_5348,N_4213,N_4471);
or U5349 (N_5349,N_4669,N_4610);
nor U5350 (N_5350,N_4730,N_4626);
and U5351 (N_5351,N_4340,N_4484);
nand U5352 (N_5352,N_4235,N_4776);
xor U5353 (N_5353,N_4319,N_4476);
xor U5354 (N_5354,N_4278,N_4331);
or U5355 (N_5355,N_4209,N_4649);
nand U5356 (N_5356,N_4468,N_4566);
or U5357 (N_5357,N_4451,N_4642);
and U5358 (N_5358,N_4356,N_4551);
or U5359 (N_5359,N_4634,N_4758);
nor U5360 (N_5360,N_4602,N_4407);
nor U5361 (N_5361,N_4319,N_4388);
xor U5362 (N_5362,N_4612,N_4617);
nor U5363 (N_5363,N_4638,N_4598);
nor U5364 (N_5364,N_4437,N_4282);
and U5365 (N_5365,N_4358,N_4726);
and U5366 (N_5366,N_4613,N_4500);
nor U5367 (N_5367,N_4229,N_4349);
and U5368 (N_5368,N_4207,N_4336);
and U5369 (N_5369,N_4226,N_4385);
nor U5370 (N_5370,N_4368,N_4453);
or U5371 (N_5371,N_4508,N_4618);
nor U5372 (N_5372,N_4646,N_4425);
xor U5373 (N_5373,N_4334,N_4606);
and U5374 (N_5374,N_4711,N_4482);
nand U5375 (N_5375,N_4552,N_4762);
nand U5376 (N_5376,N_4716,N_4261);
xnor U5377 (N_5377,N_4288,N_4544);
and U5378 (N_5378,N_4414,N_4459);
and U5379 (N_5379,N_4634,N_4335);
nand U5380 (N_5380,N_4557,N_4630);
nand U5381 (N_5381,N_4758,N_4437);
nand U5382 (N_5382,N_4619,N_4552);
or U5383 (N_5383,N_4714,N_4429);
and U5384 (N_5384,N_4740,N_4481);
and U5385 (N_5385,N_4239,N_4716);
nor U5386 (N_5386,N_4714,N_4306);
nand U5387 (N_5387,N_4662,N_4692);
xor U5388 (N_5388,N_4601,N_4674);
nor U5389 (N_5389,N_4584,N_4550);
and U5390 (N_5390,N_4660,N_4626);
nand U5391 (N_5391,N_4405,N_4606);
nand U5392 (N_5392,N_4528,N_4427);
xor U5393 (N_5393,N_4539,N_4451);
or U5394 (N_5394,N_4788,N_4423);
and U5395 (N_5395,N_4213,N_4566);
nor U5396 (N_5396,N_4554,N_4547);
and U5397 (N_5397,N_4471,N_4418);
and U5398 (N_5398,N_4694,N_4280);
or U5399 (N_5399,N_4416,N_4714);
nor U5400 (N_5400,N_4919,N_4921);
and U5401 (N_5401,N_5137,N_5190);
nand U5402 (N_5402,N_5395,N_5320);
nand U5403 (N_5403,N_5000,N_4900);
nand U5404 (N_5404,N_5111,N_5005);
nand U5405 (N_5405,N_5260,N_5308);
or U5406 (N_5406,N_5200,N_5258);
xor U5407 (N_5407,N_5007,N_4975);
nand U5408 (N_5408,N_5339,N_4869);
nand U5409 (N_5409,N_5052,N_5332);
and U5410 (N_5410,N_4882,N_5094);
and U5411 (N_5411,N_4951,N_4842);
and U5412 (N_5412,N_5098,N_4848);
nand U5413 (N_5413,N_4952,N_5170);
xnor U5414 (N_5414,N_5152,N_5041);
nand U5415 (N_5415,N_5364,N_5374);
nor U5416 (N_5416,N_5344,N_5149);
and U5417 (N_5417,N_4844,N_5133);
or U5418 (N_5418,N_5159,N_4861);
and U5419 (N_5419,N_5286,N_4903);
xor U5420 (N_5420,N_4956,N_5150);
or U5421 (N_5421,N_4945,N_4831);
nand U5422 (N_5422,N_5178,N_4814);
nor U5423 (N_5423,N_5036,N_5165);
nor U5424 (N_5424,N_4899,N_5168);
nor U5425 (N_5425,N_5251,N_4853);
or U5426 (N_5426,N_5132,N_4867);
and U5427 (N_5427,N_5342,N_5011);
and U5428 (N_5428,N_5363,N_5303);
nand U5429 (N_5429,N_4858,N_4875);
nor U5430 (N_5430,N_5086,N_4823);
xor U5431 (N_5431,N_4863,N_5390);
or U5432 (N_5432,N_5093,N_4877);
xnor U5433 (N_5433,N_5256,N_5375);
or U5434 (N_5434,N_5201,N_5311);
xor U5435 (N_5435,N_5001,N_5026);
xnor U5436 (N_5436,N_5250,N_4826);
xnor U5437 (N_5437,N_5044,N_4990);
nand U5438 (N_5438,N_5046,N_4930);
nor U5439 (N_5439,N_5230,N_4908);
nand U5440 (N_5440,N_5072,N_4907);
xnor U5441 (N_5441,N_4935,N_4818);
or U5442 (N_5442,N_5232,N_5184);
and U5443 (N_5443,N_5009,N_5373);
xnor U5444 (N_5444,N_5182,N_5157);
xor U5445 (N_5445,N_5143,N_5199);
xor U5446 (N_5446,N_5075,N_5291);
nor U5447 (N_5447,N_4983,N_5108);
and U5448 (N_5448,N_4839,N_5349);
nor U5449 (N_5449,N_4854,N_5281);
nor U5450 (N_5450,N_4896,N_4891);
and U5451 (N_5451,N_4970,N_5037);
nand U5452 (N_5452,N_5119,N_5128);
and U5453 (N_5453,N_5099,N_5144);
and U5454 (N_5454,N_5361,N_5326);
and U5455 (N_5455,N_4878,N_5126);
nor U5456 (N_5456,N_4906,N_5279);
xor U5457 (N_5457,N_4874,N_5204);
xor U5458 (N_5458,N_5097,N_5155);
xor U5459 (N_5459,N_4810,N_5218);
nor U5460 (N_5460,N_5255,N_5302);
xor U5461 (N_5461,N_4885,N_4909);
nor U5462 (N_5462,N_4841,N_4954);
and U5463 (N_5463,N_4929,N_5181);
nand U5464 (N_5464,N_4847,N_5307);
or U5465 (N_5465,N_5027,N_5338);
nand U5466 (N_5466,N_5248,N_5234);
or U5467 (N_5467,N_5317,N_4991);
and U5468 (N_5468,N_5039,N_4911);
and U5469 (N_5469,N_5171,N_4941);
nor U5470 (N_5470,N_4996,N_5348);
or U5471 (N_5471,N_5070,N_4856);
xor U5472 (N_5472,N_4862,N_5154);
or U5473 (N_5473,N_4984,N_5221);
and U5474 (N_5474,N_5240,N_5387);
nor U5475 (N_5475,N_5136,N_5147);
and U5476 (N_5476,N_5369,N_4802);
xor U5477 (N_5477,N_5219,N_5063);
nor U5478 (N_5478,N_5354,N_5213);
nand U5479 (N_5479,N_5372,N_5092);
and U5480 (N_5480,N_4803,N_5224);
xor U5481 (N_5481,N_5129,N_4840);
nand U5482 (N_5482,N_5145,N_5319);
and U5483 (N_5483,N_5306,N_4923);
xor U5484 (N_5484,N_5151,N_4827);
nor U5485 (N_5485,N_4946,N_5254);
nand U5486 (N_5486,N_5022,N_5162);
nand U5487 (N_5487,N_5069,N_4998);
nand U5488 (N_5488,N_5140,N_5288);
and U5489 (N_5489,N_4947,N_5167);
nand U5490 (N_5490,N_4905,N_4922);
or U5491 (N_5491,N_5225,N_4817);
and U5492 (N_5492,N_5280,N_4944);
nand U5493 (N_5493,N_4948,N_5025);
xor U5494 (N_5494,N_5135,N_5187);
or U5495 (N_5495,N_5183,N_5077);
nand U5496 (N_5496,N_5214,N_5379);
nor U5497 (N_5497,N_5276,N_5310);
nand U5498 (N_5498,N_4825,N_4913);
and U5499 (N_5499,N_5090,N_5067);
and U5500 (N_5500,N_5125,N_5314);
nand U5501 (N_5501,N_4808,N_5004);
nand U5502 (N_5502,N_5360,N_4821);
nand U5503 (N_5503,N_4979,N_5362);
and U5504 (N_5504,N_5083,N_5223);
nand U5505 (N_5505,N_4912,N_4883);
and U5506 (N_5506,N_5180,N_5381);
or U5507 (N_5507,N_5220,N_4809);
nand U5508 (N_5508,N_5212,N_5292);
and U5509 (N_5509,N_5050,N_5085);
nor U5510 (N_5510,N_5122,N_5239);
nand U5511 (N_5511,N_5206,N_4961);
and U5512 (N_5512,N_5355,N_5247);
and U5513 (N_5513,N_5068,N_4849);
or U5514 (N_5514,N_5327,N_4881);
and U5515 (N_5515,N_5029,N_5043);
and U5516 (N_5516,N_5089,N_5301);
and U5517 (N_5517,N_4925,N_5104);
or U5518 (N_5518,N_5203,N_5146);
xnor U5519 (N_5519,N_5179,N_5282);
or U5520 (N_5520,N_5261,N_4931);
nand U5521 (N_5521,N_4981,N_4894);
and U5522 (N_5522,N_5296,N_5350);
and U5523 (N_5523,N_5321,N_4835);
nor U5524 (N_5524,N_5065,N_5138);
or U5525 (N_5525,N_5298,N_5018);
and U5526 (N_5526,N_5262,N_4936);
nand U5527 (N_5527,N_5335,N_4997);
nand U5528 (N_5528,N_5116,N_4959);
or U5529 (N_5529,N_4958,N_5346);
or U5530 (N_5530,N_4924,N_5019);
nand U5531 (N_5531,N_5396,N_5345);
or U5532 (N_5532,N_4904,N_5356);
and U5533 (N_5533,N_4887,N_5377);
xnor U5534 (N_5534,N_5048,N_5117);
nor U5535 (N_5535,N_5285,N_5031);
or U5536 (N_5536,N_5392,N_4864);
nor U5537 (N_5537,N_4829,N_5141);
or U5538 (N_5538,N_5283,N_5134);
nand U5539 (N_5539,N_5318,N_5290);
nor U5540 (N_5540,N_5388,N_4940);
or U5541 (N_5541,N_5289,N_5188);
xnor U5542 (N_5542,N_5278,N_5002);
nor U5543 (N_5543,N_5231,N_5228);
nor U5544 (N_5544,N_5185,N_4898);
nor U5545 (N_5545,N_5079,N_5120);
xnor U5546 (N_5546,N_4837,N_5323);
and U5547 (N_5547,N_5193,N_5160);
nor U5548 (N_5548,N_5299,N_5367);
nand U5549 (N_5549,N_5123,N_5233);
xnor U5550 (N_5550,N_5268,N_5366);
or U5551 (N_5551,N_5365,N_5166);
xnor U5552 (N_5552,N_5236,N_5164);
and U5553 (N_5553,N_4830,N_4889);
nor U5554 (N_5554,N_5257,N_5352);
or U5555 (N_5555,N_5066,N_5294);
or U5556 (N_5556,N_4880,N_5161);
nand U5557 (N_5557,N_4805,N_4914);
nand U5558 (N_5558,N_4972,N_5192);
or U5559 (N_5559,N_4942,N_5186);
nand U5560 (N_5560,N_5358,N_5091);
or U5561 (N_5561,N_4801,N_5386);
or U5562 (N_5562,N_5101,N_5341);
and U5563 (N_5563,N_5191,N_4992);
and U5564 (N_5564,N_5370,N_4813);
xor U5565 (N_5565,N_4845,N_5107);
nand U5566 (N_5566,N_5347,N_5081);
xnor U5567 (N_5567,N_5024,N_4901);
nand U5568 (N_5568,N_5383,N_5391);
or U5569 (N_5569,N_5252,N_5131);
nand U5570 (N_5570,N_4812,N_4870);
nand U5571 (N_5571,N_5163,N_4815);
and U5572 (N_5572,N_5304,N_4932);
nand U5573 (N_5573,N_5028,N_5270);
nand U5574 (N_5574,N_4957,N_5238);
and U5575 (N_5575,N_4977,N_5003);
or U5576 (N_5576,N_5053,N_4832);
nor U5577 (N_5577,N_4859,N_5194);
or U5578 (N_5578,N_5118,N_4860);
and U5579 (N_5579,N_4938,N_5353);
nor U5580 (N_5580,N_4824,N_5343);
and U5581 (N_5581,N_4963,N_5045);
xor U5582 (N_5582,N_5095,N_5158);
xor U5583 (N_5583,N_5080,N_4852);
or U5584 (N_5584,N_5084,N_4804);
and U5585 (N_5585,N_4933,N_5226);
and U5586 (N_5586,N_5062,N_4822);
nor U5587 (N_5587,N_5035,N_5249);
xor U5588 (N_5588,N_4879,N_5176);
nand U5589 (N_5589,N_5013,N_5385);
or U5590 (N_5590,N_5210,N_5102);
or U5591 (N_5591,N_4836,N_5114);
nor U5592 (N_5592,N_5017,N_4916);
or U5593 (N_5593,N_4974,N_5380);
and U5594 (N_5594,N_4971,N_5061);
nor U5595 (N_5595,N_5284,N_5078);
or U5596 (N_5596,N_4868,N_5351);
xor U5597 (N_5597,N_5269,N_5293);
or U5598 (N_5598,N_5047,N_4866);
xnor U5599 (N_5599,N_4987,N_5274);
and U5600 (N_5600,N_4865,N_5038);
and U5601 (N_5601,N_4937,N_4886);
and U5602 (N_5602,N_5087,N_4902);
and U5603 (N_5603,N_5242,N_4846);
nand U5604 (N_5604,N_5227,N_5244);
nand U5605 (N_5605,N_5336,N_5216);
and U5606 (N_5606,N_5267,N_5305);
or U5607 (N_5607,N_5175,N_5331);
nor U5608 (N_5608,N_5325,N_4816);
xor U5609 (N_5609,N_5273,N_5246);
nor U5610 (N_5610,N_4871,N_4806);
nand U5611 (N_5611,N_5329,N_5121);
xor U5612 (N_5612,N_4915,N_5371);
and U5613 (N_5613,N_5020,N_5202);
nor U5614 (N_5614,N_4966,N_4872);
xnor U5615 (N_5615,N_5115,N_5015);
nand U5616 (N_5616,N_4876,N_5198);
and U5617 (N_5617,N_4943,N_5127);
and U5618 (N_5618,N_5197,N_4934);
nor U5619 (N_5619,N_5169,N_5110);
xor U5620 (N_5620,N_4995,N_5368);
or U5621 (N_5621,N_5008,N_5034);
xnor U5622 (N_5622,N_4895,N_4850);
or U5623 (N_5623,N_5109,N_4910);
xor U5624 (N_5624,N_5312,N_4811);
xnor U5625 (N_5625,N_5139,N_5174);
nor U5626 (N_5626,N_4988,N_5315);
xnor U5627 (N_5627,N_5056,N_4918);
xnor U5628 (N_5628,N_4807,N_4851);
xnor U5629 (N_5629,N_4989,N_5058);
or U5630 (N_5630,N_4980,N_5215);
or U5631 (N_5631,N_4838,N_4967);
or U5632 (N_5632,N_5074,N_4927);
and U5633 (N_5633,N_4968,N_5054);
or U5634 (N_5634,N_4955,N_4843);
nand U5635 (N_5635,N_5012,N_4917);
or U5636 (N_5636,N_5113,N_5195);
nand U5637 (N_5637,N_4994,N_4978);
xnor U5638 (N_5638,N_5010,N_5266);
and U5639 (N_5639,N_5376,N_5082);
xor U5640 (N_5640,N_5397,N_5106);
xnor U5641 (N_5641,N_5271,N_4890);
nor U5642 (N_5642,N_4893,N_5259);
nand U5643 (N_5643,N_5211,N_5275);
nor U5644 (N_5644,N_5040,N_5148);
or U5645 (N_5645,N_5156,N_5064);
and U5646 (N_5646,N_5059,N_5399);
xnor U5647 (N_5647,N_5235,N_5324);
nor U5648 (N_5648,N_5105,N_5300);
or U5649 (N_5649,N_5322,N_5253);
nand U5650 (N_5650,N_4888,N_5049);
nand U5651 (N_5651,N_5297,N_5209);
or U5652 (N_5652,N_4857,N_5100);
and U5653 (N_5653,N_4884,N_4962);
or U5654 (N_5654,N_5088,N_5173);
xnor U5655 (N_5655,N_5055,N_4960);
xor U5656 (N_5656,N_4926,N_5205);
and U5657 (N_5657,N_5124,N_5328);
nand U5658 (N_5658,N_5023,N_4833);
or U5659 (N_5659,N_4969,N_4985);
xor U5660 (N_5660,N_5394,N_5222);
and U5661 (N_5661,N_5032,N_5217);
nor U5662 (N_5662,N_5189,N_5389);
nand U5663 (N_5663,N_5316,N_4892);
or U5664 (N_5664,N_4834,N_5309);
nor U5665 (N_5665,N_4920,N_4964);
and U5666 (N_5666,N_5277,N_5243);
nor U5667 (N_5667,N_5103,N_4953);
nand U5668 (N_5668,N_5153,N_5357);
nor U5669 (N_5669,N_5060,N_5096);
and U5670 (N_5670,N_4873,N_5021);
and U5671 (N_5671,N_5130,N_5393);
or U5672 (N_5672,N_4855,N_4828);
and U5673 (N_5673,N_5265,N_4820);
and U5674 (N_5674,N_5340,N_5073);
nand U5675 (N_5675,N_5245,N_5207);
or U5676 (N_5676,N_4973,N_5177);
and U5677 (N_5677,N_5051,N_4982);
or U5678 (N_5678,N_4993,N_5142);
and U5679 (N_5679,N_5030,N_5334);
or U5680 (N_5680,N_5071,N_5333);
or U5681 (N_5681,N_4965,N_5172);
or U5682 (N_5682,N_4999,N_5295);
nor U5683 (N_5683,N_5016,N_5313);
nand U5684 (N_5684,N_5196,N_5014);
or U5685 (N_5685,N_5229,N_5112);
and U5686 (N_5686,N_4976,N_5264);
or U5687 (N_5687,N_5076,N_5398);
and U5688 (N_5688,N_5287,N_5382);
and U5689 (N_5689,N_5378,N_5337);
or U5690 (N_5690,N_5057,N_5330);
or U5691 (N_5691,N_4950,N_5384);
nor U5692 (N_5692,N_4819,N_5272);
xor U5693 (N_5693,N_4897,N_4949);
xor U5694 (N_5694,N_5033,N_4986);
or U5695 (N_5695,N_5006,N_5241);
and U5696 (N_5696,N_5237,N_4800);
or U5697 (N_5697,N_4928,N_5359);
and U5698 (N_5698,N_4939,N_5263);
nor U5699 (N_5699,N_5208,N_5042);
or U5700 (N_5700,N_5014,N_4884);
nand U5701 (N_5701,N_4896,N_5167);
or U5702 (N_5702,N_4981,N_5118);
nor U5703 (N_5703,N_5013,N_5377);
nor U5704 (N_5704,N_4918,N_5297);
or U5705 (N_5705,N_5279,N_5150);
nand U5706 (N_5706,N_5193,N_5231);
or U5707 (N_5707,N_5392,N_5078);
and U5708 (N_5708,N_5017,N_4878);
xor U5709 (N_5709,N_4966,N_5035);
nand U5710 (N_5710,N_5139,N_5221);
xnor U5711 (N_5711,N_4892,N_4984);
or U5712 (N_5712,N_5179,N_5262);
nand U5713 (N_5713,N_5150,N_5325);
nor U5714 (N_5714,N_5288,N_5194);
and U5715 (N_5715,N_5078,N_5232);
nand U5716 (N_5716,N_5203,N_5193);
xnor U5717 (N_5717,N_5218,N_5188);
xnor U5718 (N_5718,N_4861,N_4939);
nand U5719 (N_5719,N_5231,N_5128);
nor U5720 (N_5720,N_5251,N_5176);
nand U5721 (N_5721,N_4866,N_4974);
xnor U5722 (N_5722,N_5000,N_5069);
or U5723 (N_5723,N_5079,N_5226);
nor U5724 (N_5724,N_5352,N_5346);
nand U5725 (N_5725,N_5138,N_5047);
and U5726 (N_5726,N_4935,N_5058);
or U5727 (N_5727,N_4934,N_5133);
nor U5728 (N_5728,N_5254,N_4906);
nor U5729 (N_5729,N_5019,N_5316);
or U5730 (N_5730,N_5395,N_4880);
and U5731 (N_5731,N_5075,N_5213);
or U5732 (N_5732,N_5320,N_4841);
and U5733 (N_5733,N_4906,N_5276);
or U5734 (N_5734,N_5119,N_5276);
nand U5735 (N_5735,N_5177,N_4964);
xor U5736 (N_5736,N_5326,N_4898);
nor U5737 (N_5737,N_5291,N_4859);
nand U5738 (N_5738,N_4897,N_4816);
nand U5739 (N_5739,N_5132,N_5095);
or U5740 (N_5740,N_4983,N_5020);
or U5741 (N_5741,N_5327,N_5155);
nand U5742 (N_5742,N_4845,N_5204);
and U5743 (N_5743,N_5087,N_4830);
xnor U5744 (N_5744,N_5169,N_5359);
or U5745 (N_5745,N_4887,N_4918);
and U5746 (N_5746,N_5389,N_5179);
nor U5747 (N_5747,N_5001,N_5115);
nand U5748 (N_5748,N_5382,N_5043);
or U5749 (N_5749,N_5171,N_5284);
and U5750 (N_5750,N_5200,N_5127);
and U5751 (N_5751,N_4952,N_5155);
and U5752 (N_5752,N_4887,N_5321);
nor U5753 (N_5753,N_5277,N_5042);
or U5754 (N_5754,N_5099,N_5201);
nand U5755 (N_5755,N_5244,N_5181);
xnor U5756 (N_5756,N_4830,N_4850);
nor U5757 (N_5757,N_5190,N_4803);
xor U5758 (N_5758,N_4942,N_4961);
xor U5759 (N_5759,N_5398,N_5361);
xor U5760 (N_5760,N_5232,N_4853);
nand U5761 (N_5761,N_5170,N_5268);
or U5762 (N_5762,N_4909,N_4877);
or U5763 (N_5763,N_4944,N_4926);
nand U5764 (N_5764,N_5291,N_4826);
or U5765 (N_5765,N_5053,N_5071);
xor U5766 (N_5766,N_4885,N_5131);
nor U5767 (N_5767,N_5263,N_5279);
nor U5768 (N_5768,N_5000,N_5378);
or U5769 (N_5769,N_5194,N_5051);
and U5770 (N_5770,N_5285,N_4956);
and U5771 (N_5771,N_4810,N_5305);
nand U5772 (N_5772,N_5229,N_5009);
xor U5773 (N_5773,N_4988,N_5322);
nand U5774 (N_5774,N_5164,N_5221);
nand U5775 (N_5775,N_5140,N_5095);
and U5776 (N_5776,N_5025,N_5156);
and U5777 (N_5777,N_5100,N_5057);
nor U5778 (N_5778,N_5154,N_5230);
nor U5779 (N_5779,N_5334,N_5002);
and U5780 (N_5780,N_5175,N_5131);
nand U5781 (N_5781,N_5139,N_4926);
nand U5782 (N_5782,N_5011,N_5323);
and U5783 (N_5783,N_5359,N_5144);
nand U5784 (N_5784,N_5001,N_4990);
and U5785 (N_5785,N_5373,N_5104);
and U5786 (N_5786,N_5191,N_4809);
xnor U5787 (N_5787,N_5250,N_5151);
and U5788 (N_5788,N_5339,N_5365);
nand U5789 (N_5789,N_5067,N_5387);
or U5790 (N_5790,N_4814,N_5258);
nand U5791 (N_5791,N_5027,N_5260);
nor U5792 (N_5792,N_5226,N_5193);
and U5793 (N_5793,N_5073,N_4994);
xor U5794 (N_5794,N_4817,N_5201);
nand U5795 (N_5795,N_4848,N_5021);
or U5796 (N_5796,N_5298,N_5287);
nand U5797 (N_5797,N_5072,N_5267);
nand U5798 (N_5798,N_5326,N_5042);
and U5799 (N_5799,N_5202,N_5219);
or U5800 (N_5800,N_5046,N_4868);
nand U5801 (N_5801,N_5079,N_4956);
and U5802 (N_5802,N_5112,N_5263);
nand U5803 (N_5803,N_5059,N_5375);
or U5804 (N_5804,N_5022,N_5186);
and U5805 (N_5805,N_4809,N_4842);
xor U5806 (N_5806,N_5388,N_4852);
xor U5807 (N_5807,N_5145,N_5026);
or U5808 (N_5808,N_4914,N_5250);
and U5809 (N_5809,N_4974,N_4918);
nor U5810 (N_5810,N_5319,N_4915);
and U5811 (N_5811,N_5196,N_4992);
nor U5812 (N_5812,N_5298,N_5253);
or U5813 (N_5813,N_5024,N_5165);
and U5814 (N_5814,N_4881,N_4869);
xor U5815 (N_5815,N_5285,N_5356);
xnor U5816 (N_5816,N_5105,N_5072);
and U5817 (N_5817,N_4906,N_4892);
or U5818 (N_5818,N_4825,N_4934);
xor U5819 (N_5819,N_4959,N_5319);
and U5820 (N_5820,N_5078,N_4824);
nand U5821 (N_5821,N_4813,N_4863);
and U5822 (N_5822,N_4953,N_5004);
or U5823 (N_5823,N_5373,N_5198);
and U5824 (N_5824,N_4958,N_5318);
xor U5825 (N_5825,N_4991,N_5358);
nand U5826 (N_5826,N_4869,N_5229);
nor U5827 (N_5827,N_5269,N_5386);
xor U5828 (N_5828,N_4947,N_5034);
or U5829 (N_5829,N_5359,N_5287);
nor U5830 (N_5830,N_4927,N_5397);
or U5831 (N_5831,N_5160,N_4977);
or U5832 (N_5832,N_4928,N_5054);
or U5833 (N_5833,N_5068,N_4880);
and U5834 (N_5834,N_4858,N_5365);
or U5835 (N_5835,N_5268,N_5311);
nor U5836 (N_5836,N_5374,N_5113);
or U5837 (N_5837,N_4813,N_4935);
or U5838 (N_5838,N_5111,N_5347);
xor U5839 (N_5839,N_4999,N_5080);
or U5840 (N_5840,N_5235,N_5229);
xnor U5841 (N_5841,N_5109,N_4905);
nor U5842 (N_5842,N_5060,N_5250);
or U5843 (N_5843,N_4876,N_4812);
nor U5844 (N_5844,N_5374,N_4859);
nand U5845 (N_5845,N_5253,N_5096);
nand U5846 (N_5846,N_5314,N_5216);
nand U5847 (N_5847,N_4941,N_5102);
nor U5848 (N_5848,N_4826,N_5103);
nor U5849 (N_5849,N_4928,N_4931);
nand U5850 (N_5850,N_5087,N_5363);
xnor U5851 (N_5851,N_4800,N_5155);
and U5852 (N_5852,N_5070,N_4968);
nand U5853 (N_5853,N_4840,N_4953);
and U5854 (N_5854,N_4832,N_5111);
nand U5855 (N_5855,N_5064,N_5216);
nor U5856 (N_5856,N_4806,N_4860);
and U5857 (N_5857,N_5399,N_5130);
or U5858 (N_5858,N_5248,N_5081);
nor U5859 (N_5859,N_4943,N_5082);
nor U5860 (N_5860,N_5082,N_5157);
nor U5861 (N_5861,N_4807,N_5395);
xnor U5862 (N_5862,N_5373,N_5081);
or U5863 (N_5863,N_5270,N_5015);
and U5864 (N_5864,N_5395,N_5348);
or U5865 (N_5865,N_4914,N_5137);
xor U5866 (N_5866,N_4840,N_4800);
or U5867 (N_5867,N_4977,N_4930);
nor U5868 (N_5868,N_5120,N_5074);
and U5869 (N_5869,N_5005,N_5239);
and U5870 (N_5870,N_5177,N_5313);
or U5871 (N_5871,N_4959,N_4938);
or U5872 (N_5872,N_4910,N_5019);
and U5873 (N_5873,N_4821,N_4809);
nor U5874 (N_5874,N_5101,N_5365);
nand U5875 (N_5875,N_5172,N_5320);
xnor U5876 (N_5876,N_5124,N_4932);
and U5877 (N_5877,N_4801,N_5249);
xnor U5878 (N_5878,N_5130,N_4902);
nand U5879 (N_5879,N_4979,N_4872);
or U5880 (N_5880,N_4934,N_5144);
nor U5881 (N_5881,N_5229,N_4832);
and U5882 (N_5882,N_5247,N_5291);
nand U5883 (N_5883,N_5223,N_4944);
or U5884 (N_5884,N_5081,N_5101);
nor U5885 (N_5885,N_5183,N_4863);
xor U5886 (N_5886,N_4899,N_5366);
nand U5887 (N_5887,N_5285,N_5075);
nand U5888 (N_5888,N_5242,N_5273);
and U5889 (N_5889,N_4837,N_5008);
xor U5890 (N_5890,N_4935,N_4955);
xnor U5891 (N_5891,N_5095,N_5188);
or U5892 (N_5892,N_5239,N_5199);
or U5893 (N_5893,N_5210,N_4913);
or U5894 (N_5894,N_4812,N_4838);
xnor U5895 (N_5895,N_5010,N_5089);
or U5896 (N_5896,N_5364,N_5082);
xnor U5897 (N_5897,N_4996,N_4858);
nand U5898 (N_5898,N_4881,N_5036);
xnor U5899 (N_5899,N_5397,N_4982);
or U5900 (N_5900,N_5249,N_5241);
or U5901 (N_5901,N_5353,N_5351);
and U5902 (N_5902,N_4802,N_5209);
and U5903 (N_5903,N_5394,N_5201);
nor U5904 (N_5904,N_5076,N_5168);
or U5905 (N_5905,N_5118,N_4862);
or U5906 (N_5906,N_5364,N_4959);
or U5907 (N_5907,N_5019,N_5180);
or U5908 (N_5908,N_5017,N_5081);
nand U5909 (N_5909,N_4952,N_5348);
xor U5910 (N_5910,N_4878,N_5358);
or U5911 (N_5911,N_4831,N_5249);
or U5912 (N_5912,N_4942,N_5203);
xnor U5913 (N_5913,N_5246,N_5313);
nand U5914 (N_5914,N_5345,N_4808);
nand U5915 (N_5915,N_5373,N_4895);
or U5916 (N_5916,N_5128,N_5347);
or U5917 (N_5917,N_5024,N_5150);
xor U5918 (N_5918,N_5040,N_4826);
xnor U5919 (N_5919,N_5151,N_5155);
xor U5920 (N_5920,N_5318,N_4935);
xor U5921 (N_5921,N_5299,N_5353);
and U5922 (N_5922,N_5164,N_5321);
or U5923 (N_5923,N_5096,N_5395);
xor U5924 (N_5924,N_4892,N_5259);
xnor U5925 (N_5925,N_5343,N_4917);
nor U5926 (N_5926,N_5323,N_4950);
xnor U5927 (N_5927,N_5178,N_5398);
xnor U5928 (N_5928,N_5373,N_5036);
xor U5929 (N_5929,N_5023,N_5120);
nor U5930 (N_5930,N_4932,N_4866);
nor U5931 (N_5931,N_5343,N_5215);
xnor U5932 (N_5932,N_5264,N_4985);
and U5933 (N_5933,N_5374,N_4913);
nand U5934 (N_5934,N_5165,N_4954);
or U5935 (N_5935,N_4960,N_5206);
xnor U5936 (N_5936,N_5381,N_4992);
and U5937 (N_5937,N_4882,N_5025);
and U5938 (N_5938,N_5303,N_4843);
nand U5939 (N_5939,N_4874,N_5056);
nand U5940 (N_5940,N_5104,N_4808);
xnor U5941 (N_5941,N_5021,N_5395);
nand U5942 (N_5942,N_5259,N_5323);
nor U5943 (N_5943,N_5312,N_5184);
nand U5944 (N_5944,N_4994,N_5074);
and U5945 (N_5945,N_5116,N_5064);
nor U5946 (N_5946,N_5324,N_5044);
and U5947 (N_5947,N_5297,N_4829);
xor U5948 (N_5948,N_4919,N_4877);
nand U5949 (N_5949,N_5206,N_4839);
nand U5950 (N_5950,N_5176,N_5078);
nand U5951 (N_5951,N_5076,N_5346);
xor U5952 (N_5952,N_4936,N_5153);
xnor U5953 (N_5953,N_4872,N_5193);
xor U5954 (N_5954,N_5098,N_5173);
or U5955 (N_5955,N_4901,N_5195);
or U5956 (N_5956,N_5334,N_5380);
or U5957 (N_5957,N_5289,N_5082);
nor U5958 (N_5958,N_5281,N_5272);
nand U5959 (N_5959,N_4843,N_5386);
nand U5960 (N_5960,N_5141,N_5101);
nor U5961 (N_5961,N_5061,N_5366);
nand U5962 (N_5962,N_5159,N_5394);
xnor U5963 (N_5963,N_4941,N_5018);
and U5964 (N_5964,N_5255,N_4898);
and U5965 (N_5965,N_5234,N_4806);
or U5966 (N_5966,N_5060,N_4866);
nand U5967 (N_5967,N_4904,N_4891);
xor U5968 (N_5968,N_5069,N_5062);
or U5969 (N_5969,N_4859,N_4825);
xnor U5970 (N_5970,N_4893,N_4858);
nor U5971 (N_5971,N_5390,N_5226);
xnor U5972 (N_5972,N_5261,N_5057);
nor U5973 (N_5973,N_4806,N_4814);
xnor U5974 (N_5974,N_5066,N_5010);
nand U5975 (N_5975,N_5388,N_5317);
nor U5976 (N_5976,N_4986,N_5338);
nand U5977 (N_5977,N_5305,N_5069);
and U5978 (N_5978,N_4991,N_4906);
and U5979 (N_5979,N_5077,N_4939);
nand U5980 (N_5980,N_5250,N_4833);
nand U5981 (N_5981,N_5134,N_4809);
nand U5982 (N_5982,N_4967,N_4931);
xnor U5983 (N_5983,N_5044,N_5184);
nor U5984 (N_5984,N_5367,N_4948);
nor U5985 (N_5985,N_5307,N_4992);
or U5986 (N_5986,N_4842,N_5319);
or U5987 (N_5987,N_5306,N_4944);
nor U5988 (N_5988,N_5020,N_4916);
nand U5989 (N_5989,N_5125,N_5152);
nand U5990 (N_5990,N_5158,N_5363);
nor U5991 (N_5991,N_5235,N_4865);
xor U5992 (N_5992,N_4988,N_5122);
xnor U5993 (N_5993,N_4865,N_5041);
nor U5994 (N_5994,N_5353,N_4982);
nand U5995 (N_5995,N_5086,N_4887);
and U5996 (N_5996,N_5382,N_5310);
and U5997 (N_5997,N_5107,N_5045);
nand U5998 (N_5998,N_5211,N_4866);
and U5999 (N_5999,N_5335,N_5169);
or U6000 (N_6000,N_5831,N_5714);
and U6001 (N_6001,N_5424,N_5922);
and U6002 (N_6002,N_5745,N_5582);
xnor U6003 (N_6003,N_5559,N_5854);
nor U6004 (N_6004,N_5778,N_5614);
nand U6005 (N_6005,N_5526,N_5796);
and U6006 (N_6006,N_5679,N_5902);
nor U6007 (N_6007,N_5690,N_5988);
xnor U6008 (N_6008,N_5979,N_5755);
or U6009 (N_6009,N_5704,N_5877);
nor U6010 (N_6010,N_5449,N_5956);
xor U6011 (N_6011,N_5895,N_5828);
or U6012 (N_6012,N_5867,N_5475);
or U6013 (N_6013,N_5550,N_5490);
xor U6014 (N_6014,N_5918,N_5729);
nand U6015 (N_6015,N_5676,N_5842);
nand U6016 (N_6016,N_5980,N_5777);
nand U6017 (N_6017,N_5914,N_5827);
xor U6018 (N_6018,N_5650,N_5900);
and U6019 (N_6019,N_5546,N_5554);
and U6020 (N_6020,N_5955,N_5558);
nand U6021 (N_6021,N_5579,N_5586);
xnor U6022 (N_6022,N_5939,N_5557);
and U6023 (N_6023,N_5468,N_5438);
or U6024 (N_6024,N_5499,N_5625);
or U6025 (N_6025,N_5869,N_5887);
nand U6026 (N_6026,N_5835,N_5686);
nor U6027 (N_6027,N_5441,N_5991);
or U6028 (N_6028,N_5949,N_5801);
xor U6029 (N_6029,N_5508,N_5551);
or U6030 (N_6030,N_5618,N_5505);
nand U6031 (N_6031,N_5765,N_5595);
xor U6032 (N_6032,N_5717,N_5760);
and U6033 (N_6033,N_5797,N_5965);
nor U6034 (N_6034,N_5450,N_5758);
and U6035 (N_6035,N_5472,N_5699);
and U6036 (N_6036,N_5581,N_5705);
or U6037 (N_6037,N_5541,N_5658);
and U6038 (N_6038,N_5478,N_5616);
or U6039 (N_6039,N_5888,N_5532);
xnor U6040 (N_6040,N_5992,N_5969);
nand U6041 (N_6041,N_5569,N_5556);
and U6042 (N_6042,N_5773,N_5401);
nor U6043 (N_6043,N_5839,N_5931);
and U6044 (N_6044,N_5696,N_5908);
nand U6045 (N_6045,N_5665,N_5452);
nor U6046 (N_6046,N_5728,N_5862);
and U6047 (N_6047,N_5471,N_5549);
nor U6048 (N_6048,N_5523,N_5788);
and U6049 (N_6049,N_5738,N_5935);
nor U6050 (N_6050,N_5975,N_5772);
or U6051 (N_6051,N_5510,N_5488);
or U6052 (N_6052,N_5832,N_5400);
and U6053 (N_6053,N_5824,N_5632);
or U6054 (N_6054,N_5740,N_5837);
nand U6055 (N_6055,N_5821,N_5563);
nand U6056 (N_6056,N_5756,N_5775);
nand U6057 (N_6057,N_5409,N_5495);
or U6058 (N_6058,N_5764,N_5851);
xnor U6059 (N_6059,N_5890,N_5711);
and U6060 (N_6060,N_5783,N_5455);
and U6061 (N_6061,N_5722,N_5730);
nor U6062 (N_6062,N_5480,N_5570);
xnor U6063 (N_6063,N_5873,N_5746);
xor U6064 (N_6064,N_5689,N_5572);
and U6065 (N_6065,N_5652,N_5709);
and U6066 (N_6066,N_5713,N_5973);
xor U6067 (N_6067,N_5637,N_5612);
or U6068 (N_6068,N_5989,N_5601);
or U6069 (N_6069,N_5448,N_5840);
nor U6070 (N_6070,N_5420,N_5896);
xnor U6071 (N_6071,N_5798,N_5810);
and U6072 (N_6072,N_5583,N_5522);
nand U6073 (N_6073,N_5863,N_5410);
xor U6074 (N_6074,N_5677,N_5574);
xor U6075 (N_6075,N_5429,N_5985);
xnor U6076 (N_6076,N_5911,N_5566);
or U6077 (N_6077,N_5720,N_5836);
xnor U6078 (N_6078,N_5520,N_5608);
or U6079 (N_6079,N_5474,N_5805);
xor U6080 (N_6080,N_5970,N_5750);
nor U6081 (N_6081,N_5633,N_5402);
nor U6082 (N_6082,N_5669,N_5536);
xor U6083 (N_6083,N_5803,N_5754);
and U6084 (N_6084,N_5963,N_5707);
xor U6085 (N_6085,N_5678,N_5509);
nor U6086 (N_6086,N_5500,N_5997);
nor U6087 (N_6087,N_5501,N_5850);
and U6088 (N_6088,N_5539,N_5567);
and U6089 (N_6089,N_5893,N_5990);
nand U6090 (N_6090,N_5858,N_5855);
and U6091 (N_6091,N_5953,N_5693);
or U6092 (N_6092,N_5675,N_5958);
and U6093 (N_6093,N_5811,N_5562);
and U6094 (N_6094,N_5636,N_5710);
and U6095 (N_6095,N_5957,N_5721);
nand U6096 (N_6096,N_5876,N_5642);
or U6097 (N_6097,N_5629,N_5643);
and U6098 (N_6098,N_5919,N_5687);
xor U6099 (N_6099,N_5882,N_5597);
nand U6100 (N_6100,N_5437,N_5433);
xnor U6101 (N_6101,N_5647,N_5761);
nand U6102 (N_6102,N_5626,N_5683);
nand U6103 (N_6103,N_5602,N_5681);
or U6104 (N_6104,N_5848,N_5528);
nor U6105 (N_6105,N_5912,N_5735);
xnor U6106 (N_6106,N_5431,N_5596);
and U6107 (N_6107,N_5723,N_5763);
nand U6108 (N_6108,N_5819,N_5892);
and U6109 (N_6109,N_5732,N_5903);
nor U6110 (N_6110,N_5483,N_5627);
or U6111 (N_6111,N_5826,N_5793);
and U6112 (N_6112,N_5898,N_5981);
nand U6113 (N_6113,N_5415,N_5942);
nand U6114 (N_6114,N_5418,N_5782);
and U6115 (N_6115,N_5927,N_5640);
nand U6116 (N_6116,N_5639,N_5535);
nor U6117 (N_6117,N_5630,N_5680);
nor U6118 (N_6118,N_5591,N_5886);
and U6119 (N_6119,N_5544,N_5947);
or U6120 (N_6120,N_5878,N_5414);
xor U6121 (N_6121,N_5611,N_5664);
or U6122 (N_6122,N_5940,N_5571);
nand U6123 (N_6123,N_5790,N_5460);
xor U6124 (N_6124,N_5982,N_5830);
nor U6125 (N_6125,N_5847,N_5426);
nand U6126 (N_6126,N_5458,N_5496);
and U6127 (N_6127,N_5482,N_5820);
nand U6128 (N_6128,N_5874,N_5945);
nand U6129 (N_6129,N_5430,N_5565);
nor U6130 (N_6130,N_5883,N_5530);
xnor U6131 (N_6131,N_5785,N_5511);
or U6132 (N_6132,N_5432,N_5906);
nand U6133 (N_6133,N_5994,N_5527);
and U6134 (N_6134,N_5879,N_5870);
or U6135 (N_6135,N_5814,N_5917);
xnor U6136 (N_6136,N_5673,N_5628);
nand U6137 (N_6137,N_5845,N_5897);
and U6138 (N_6138,N_5904,N_5833);
or U6139 (N_6139,N_5457,N_5787);
and U6140 (N_6140,N_5708,N_5408);
or U6141 (N_6141,N_5959,N_5660);
and U6142 (N_6142,N_5610,N_5473);
nor U6143 (N_6143,N_5434,N_5808);
nand U6144 (N_6144,N_5884,N_5484);
or U6145 (N_6145,N_5964,N_5674);
xnor U6146 (N_6146,N_5852,N_5446);
or U6147 (N_6147,N_5987,N_5998);
nand U6148 (N_6148,N_5776,N_5789);
nand U6149 (N_6149,N_5491,N_5442);
or U6150 (N_6150,N_5712,N_5593);
or U6151 (N_6151,N_5419,N_5654);
xor U6152 (N_6152,N_5620,N_5469);
nor U6153 (N_6153,N_5802,N_5477);
nor U6154 (N_6154,N_5463,N_5967);
xnor U6155 (N_6155,N_5771,N_5866);
or U6156 (N_6156,N_5668,N_5759);
nand U6157 (N_6157,N_5493,N_5751);
xor U6158 (N_6158,N_5823,N_5966);
nand U6159 (N_6159,N_5466,N_5464);
nor U6160 (N_6160,N_5584,N_5641);
xor U6161 (N_6161,N_5568,N_5531);
and U6162 (N_6162,N_5860,N_5781);
nand U6163 (N_6163,N_5894,N_5791);
xnor U6164 (N_6164,N_5443,N_5701);
or U6165 (N_6165,N_5984,N_5706);
xnor U6166 (N_6166,N_5916,N_5671);
xor U6167 (N_6167,N_5816,N_5698);
xnor U6168 (N_6168,N_5844,N_5983);
nand U6169 (N_6169,N_5932,N_5933);
and U6170 (N_6170,N_5909,N_5435);
xor U6171 (N_6171,N_5752,N_5749);
xor U6172 (N_6172,N_5649,N_5733);
and U6173 (N_6173,N_5993,N_5615);
xnor U6174 (N_6174,N_5807,N_5515);
xor U6175 (N_6175,N_5972,N_5951);
nand U6176 (N_6176,N_5407,N_5604);
and U6177 (N_6177,N_5659,N_5503);
and U6178 (N_6178,N_5498,N_5857);
nor U6179 (N_6179,N_5774,N_5417);
nand U6180 (N_6180,N_5403,N_5747);
nor U6181 (N_6181,N_5489,N_5743);
xnor U6182 (N_6182,N_5928,N_5538);
xor U6183 (N_6183,N_5779,N_5470);
or U6184 (N_6184,N_5999,N_5757);
or U6185 (N_6185,N_5739,N_5507);
nor U6186 (N_6186,N_5971,N_5621);
nor U6187 (N_6187,N_5891,N_5946);
or U6188 (N_6188,N_5421,N_5548);
or U6189 (N_6189,N_5924,N_5413);
nand U6190 (N_6190,N_5519,N_5542);
or U6191 (N_6191,N_5692,N_5920);
nand U6192 (N_6192,N_5838,N_5962);
and U6193 (N_6193,N_5880,N_5651);
xnor U6194 (N_6194,N_5986,N_5841);
or U6195 (N_6195,N_5913,N_5881);
nor U6196 (N_6196,N_5829,N_5447);
nand U6197 (N_6197,N_5697,N_5599);
xor U6198 (N_6198,N_5588,N_5516);
xor U6199 (N_6199,N_5813,N_5436);
nor U6200 (N_6200,N_5818,N_5533);
xnor U6201 (N_6201,N_5948,N_5792);
xor U6202 (N_6202,N_5767,N_5938);
nor U6203 (N_6203,N_5631,N_5724);
or U6204 (N_6204,N_5768,N_5657);
xnor U6205 (N_6205,N_5502,N_5667);
xor U6206 (N_6206,N_5545,N_5968);
nor U6207 (N_6207,N_5428,N_5405);
xnor U6208 (N_6208,N_5547,N_5555);
and U6209 (N_6209,N_5512,N_5825);
nand U6210 (N_6210,N_5638,N_5537);
and U6211 (N_6211,N_5451,N_5634);
xnor U6212 (N_6212,N_5961,N_5577);
or U6213 (N_6213,N_5794,N_5622);
nor U6214 (N_6214,N_5974,N_5952);
nand U6215 (N_6215,N_5529,N_5748);
xor U6216 (N_6216,N_5623,N_5694);
nand U6217 (N_6217,N_5494,N_5609);
nor U6218 (N_6218,N_5427,N_5589);
and U6219 (N_6219,N_5655,N_5521);
or U6220 (N_6220,N_5861,N_5573);
or U6221 (N_6221,N_5753,N_5461);
or U6222 (N_6222,N_5929,N_5590);
or U6223 (N_6223,N_5444,N_5404);
and U6224 (N_6224,N_5865,N_5726);
xor U6225 (N_6225,N_5624,N_5486);
or U6226 (N_6226,N_5587,N_5718);
nand U6227 (N_6227,N_5425,N_5804);
nor U6228 (N_6228,N_5762,N_5619);
xnor U6229 (N_6229,N_5485,N_5815);
nor U6230 (N_6230,N_5411,N_5766);
or U6231 (N_6231,N_5943,N_5666);
or U6232 (N_6232,N_5481,N_5926);
nor U6233 (N_6233,N_5492,N_5534);
and U6234 (N_6234,N_5644,N_5737);
and U6235 (N_6235,N_5580,N_5716);
and U6236 (N_6236,N_5476,N_5497);
nand U6237 (N_6237,N_5684,N_5670);
nor U6238 (N_6238,N_5700,N_5944);
nand U6239 (N_6239,N_5688,N_5937);
xnor U6240 (N_6240,N_5784,N_5635);
xnor U6241 (N_6241,N_5853,N_5817);
nand U6242 (N_6242,N_5682,N_5923);
xnor U6243 (N_6243,N_5504,N_5525);
and U6244 (N_6244,N_5954,N_5795);
or U6245 (N_6245,N_5822,N_5809);
or U6246 (N_6246,N_5786,N_5653);
or U6247 (N_6247,N_5479,N_5849);
and U6248 (N_6248,N_5662,N_5741);
or U6249 (N_6249,N_5467,N_5769);
and U6250 (N_6250,N_5440,N_5770);
nor U6251 (N_6251,N_5416,N_5517);
or U6252 (N_6252,N_5744,N_5846);
and U6253 (N_6253,N_5976,N_5552);
nor U6254 (N_6254,N_5871,N_5663);
or U6255 (N_6255,N_5422,N_5950);
and U6256 (N_6256,N_5702,N_5864);
or U6257 (N_6257,N_5843,N_5607);
nand U6258 (N_6258,N_5695,N_5524);
and U6259 (N_6259,N_5648,N_5872);
nand U6260 (N_6260,N_5606,N_5603);
or U6261 (N_6261,N_5930,N_5453);
xnor U6262 (N_6262,N_5941,N_5899);
or U6263 (N_6263,N_5934,N_5685);
or U6264 (N_6264,N_5465,N_5834);
nor U6265 (N_6265,N_5978,N_5423);
and U6266 (N_6266,N_5715,N_5412);
and U6267 (N_6267,N_5605,N_5905);
nor U6268 (N_6268,N_5598,N_5734);
nor U6269 (N_6269,N_5672,N_5799);
nand U6270 (N_6270,N_5439,N_5727);
nor U6271 (N_6271,N_5506,N_5600);
or U6272 (N_6272,N_5736,N_5885);
or U6273 (N_6273,N_5553,N_5543);
or U6274 (N_6274,N_5915,N_5703);
nand U6275 (N_6275,N_5936,N_5645);
nor U6276 (N_6276,N_5725,N_5456);
or U6277 (N_6277,N_5613,N_5910);
or U6278 (N_6278,N_5576,N_5925);
nand U6279 (N_6279,N_5487,N_5514);
xnor U6280 (N_6280,N_5875,N_5661);
or U6281 (N_6281,N_5921,N_5901);
and U6282 (N_6282,N_5462,N_5646);
or U6283 (N_6283,N_5856,N_5513);
or U6284 (N_6284,N_5977,N_5889);
xnor U6285 (N_6285,N_5868,N_5742);
nor U6286 (N_6286,N_5459,N_5454);
nand U6287 (N_6287,N_5806,N_5564);
nor U6288 (N_6288,N_5731,N_5561);
xnor U6289 (N_6289,N_5445,N_5578);
xnor U6290 (N_6290,N_5540,N_5656);
and U6291 (N_6291,N_5575,N_5780);
and U6292 (N_6292,N_5859,N_5907);
nor U6293 (N_6293,N_5719,N_5594);
xnor U6294 (N_6294,N_5960,N_5691);
nor U6295 (N_6295,N_5560,N_5812);
or U6296 (N_6296,N_5406,N_5585);
or U6297 (N_6297,N_5800,N_5995);
nand U6298 (N_6298,N_5518,N_5996);
xor U6299 (N_6299,N_5617,N_5592);
and U6300 (N_6300,N_5552,N_5691);
nand U6301 (N_6301,N_5431,N_5841);
xnor U6302 (N_6302,N_5461,N_5573);
xnor U6303 (N_6303,N_5653,N_5706);
nand U6304 (N_6304,N_5755,N_5947);
or U6305 (N_6305,N_5434,N_5561);
nor U6306 (N_6306,N_5894,N_5955);
nand U6307 (N_6307,N_5440,N_5810);
xnor U6308 (N_6308,N_5866,N_5897);
nand U6309 (N_6309,N_5421,N_5517);
nor U6310 (N_6310,N_5564,N_5807);
nand U6311 (N_6311,N_5569,N_5774);
xor U6312 (N_6312,N_5604,N_5987);
nand U6313 (N_6313,N_5699,N_5707);
and U6314 (N_6314,N_5495,N_5725);
xnor U6315 (N_6315,N_5497,N_5824);
xnor U6316 (N_6316,N_5535,N_5439);
nand U6317 (N_6317,N_5507,N_5729);
nor U6318 (N_6318,N_5895,N_5585);
nor U6319 (N_6319,N_5819,N_5687);
or U6320 (N_6320,N_5620,N_5530);
nand U6321 (N_6321,N_5569,N_5778);
or U6322 (N_6322,N_5856,N_5553);
and U6323 (N_6323,N_5531,N_5553);
nand U6324 (N_6324,N_5601,N_5534);
and U6325 (N_6325,N_5598,N_5559);
and U6326 (N_6326,N_5918,N_5731);
and U6327 (N_6327,N_5717,N_5805);
and U6328 (N_6328,N_5851,N_5451);
and U6329 (N_6329,N_5629,N_5481);
nand U6330 (N_6330,N_5608,N_5646);
nand U6331 (N_6331,N_5806,N_5761);
nand U6332 (N_6332,N_5957,N_5596);
nor U6333 (N_6333,N_5723,N_5740);
nand U6334 (N_6334,N_5638,N_5802);
xnor U6335 (N_6335,N_5429,N_5496);
and U6336 (N_6336,N_5634,N_5473);
and U6337 (N_6337,N_5738,N_5607);
or U6338 (N_6338,N_5662,N_5919);
nor U6339 (N_6339,N_5647,N_5997);
nor U6340 (N_6340,N_5477,N_5770);
and U6341 (N_6341,N_5473,N_5772);
nor U6342 (N_6342,N_5487,N_5652);
xor U6343 (N_6343,N_5509,N_5596);
nand U6344 (N_6344,N_5755,N_5865);
nand U6345 (N_6345,N_5464,N_5561);
nand U6346 (N_6346,N_5592,N_5977);
nor U6347 (N_6347,N_5871,N_5722);
or U6348 (N_6348,N_5875,N_5704);
xnor U6349 (N_6349,N_5803,N_5557);
xnor U6350 (N_6350,N_5729,N_5726);
nand U6351 (N_6351,N_5993,N_5445);
and U6352 (N_6352,N_5904,N_5566);
or U6353 (N_6353,N_5956,N_5818);
xnor U6354 (N_6354,N_5684,N_5469);
or U6355 (N_6355,N_5568,N_5444);
xor U6356 (N_6356,N_5469,N_5846);
nand U6357 (N_6357,N_5533,N_5448);
nand U6358 (N_6358,N_5501,N_5547);
or U6359 (N_6359,N_5834,N_5773);
nand U6360 (N_6360,N_5559,N_5539);
xor U6361 (N_6361,N_5911,N_5650);
nor U6362 (N_6362,N_5789,N_5660);
xor U6363 (N_6363,N_5716,N_5959);
or U6364 (N_6364,N_5921,N_5631);
or U6365 (N_6365,N_5877,N_5527);
nand U6366 (N_6366,N_5660,N_5729);
nand U6367 (N_6367,N_5768,N_5770);
xnor U6368 (N_6368,N_5657,N_5805);
xnor U6369 (N_6369,N_5517,N_5953);
or U6370 (N_6370,N_5734,N_5691);
or U6371 (N_6371,N_5752,N_5961);
nand U6372 (N_6372,N_5881,N_5656);
or U6373 (N_6373,N_5941,N_5734);
xor U6374 (N_6374,N_5452,N_5501);
xor U6375 (N_6375,N_5643,N_5505);
xor U6376 (N_6376,N_5681,N_5497);
nand U6377 (N_6377,N_5452,N_5785);
and U6378 (N_6378,N_5945,N_5460);
nor U6379 (N_6379,N_5821,N_5850);
or U6380 (N_6380,N_5749,N_5598);
xor U6381 (N_6381,N_5576,N_5951);
nor U6382 (N_6382,N_5857,N_5431);
xnor U6383 (N_6383,N_5978,N_5550);
xor U6384 (N_6384,N_5974,N_5823);
and U6385 (N_6385,N_5587,N_5486);
nand U6386 (N_6386,N_5496,N_5614);
or U6387 (N_6387,N_5739,N_5434);
nor U6388 (N_6388,N_5935,N_5889);
and U6389 (N_6389,N_5675,N_5505);
xor U6390 (N_6390,N_5524,N_5917);
and U6391 (N_6391,N_5519,N_5539);
nand U6392 (N_6392,N_5833,N_5691);
or U6393 (N_6393,N_5421,N_5499);
xnor U6394 (N_6394,N_5840,N_5793);
and U6395 (N_6395,N_5973,N_5504);
nor U6396 (N_6396,N_5997,N_5802);
nor U6397 (N_6397,N_5710,N_5739);
xor U6398 (N_6398,N_5604,N_5451);
and U6399 (N_6399,N_5414,N_5859);
xnor U6400 (N_6400,N_5831,N_5481);
and U6401 (N_6401,N_5873,N_5435);
and U6402 (N_6402,N_5672,N_5496);
or U6403 (N_6403,N_5430,N_5522);
and U6404 (N_6404,N_5915,N_5580);
xnor U6405 (N_6405,N_5546,N_5812);
xnor U6406 (N_6406,N_5739,N_5889);
and U6407 (N_6407,N_5680,N_5597);
or U6408 (N_6408,N_5852,N_5470);
or U6409 (N_6409,N_5808,N_5930);
or U6410 (N_6410,N_5649,N_5831);
nor U6411 (N_6411,N_5715,N_5782);
nand U6412 (N_6412,N_5745,N_5426);
and U6413 (N_6413,N_5831,N_5405);
nand U6414 (N_6414,N_5802,N_5980);
or U6415 (N_6415,N_5863,N_5534);
nor U6416 (N_6416,N_5770,N_5450);
or U6417 (N_6417,N_5905,N_5778);
nor U6418 (N_6418,N_5500,N_5783);
or U6419 (N_6419,N_5994,N_5885);
or U6420 (N_6420,N_5751,N_5691);
xor U6421 (N_6421,N_5895,N_5790);
nor U6422 (N_6422,N_5487,N_5427);
nand U6423 (N_6423,N_5764,N_5669);
or U6424 (N_6424,N_5830,N_5581);
nor U6425 (N_6425,N_5645,N_5684);
or U6426 (N_6426,N_5892,N_5863);
or U6427 (N_6427,N_5532,N_5470);
xnor U6428 (N_6428,N_5410,N_5702);
or U6429 (N_6429,N_5641,N_5917);
xnor U6430 (N_6430,N_5799,N_5655);
or U6431 (N_6431,N_5802,N_5985);
xnor U6432 (N_6432,N_5673,N_5859);
nand U6433 (N_6433,N_5923,N_5426);
or U6434 (N_6434,N_5992,N_5717);
xnor U6435 (N_6435,N_5520,N_5518);
nor U6436 (N_6436,N_5475,N_5443);
nand U6437 (N_6437,N_5666,N_5973);
or U6438 (N_6438,N_5675,N_5900);
nand U6439 (N_6439,N_5604,N_5654);
nor U6440 (N_6440,N_5853,N_5537);
xnor U6441 (N_6441,N_5438,N_5702);
or U6442 (N_6442,N_5902,N_5466);
and U6443 (N_6443,N_5402,N_5890);
nor U6444 (N_6444,N_5724,N_5457);
nand U6445 (N_6445,N_5459,N_5499);
xnor U6446 (N_6446,N_5546,N_5464);
nor U6447 (N_6447,N_5531,N_5801);
or U6448 (N_6448,N_5578,N_5552);
nand U6449 (N_6449,N_5773,N_5976);
or U6450 (N_6450,N_5698,N_5687);
or U6451 (N_6451,N_5788,N_5643);
or U6452 (N_6452,N_5837,N_5733);
nor U6453 (N_6453,N_5895,N_5709);
and U6454 (N_6454,N_5563,N_5688);
nor U6455 (N_6455,N_5800,N_5575);
or U6456 (N_6456,N_5663,N_5603);
xor U6457 (N_6457,N_5543,N_5796);
nand U6458 (N_6458,N_5810,N_5641);
nor U6459 (N_6459,N_5830,N_5693);
nor U6460 (N_6460,N_5861,N_5648);
xnor U6461 (N_6461,N_5751,N_5864);
nand U6462 (N_6462,N_5938,N_5678);
and U6463 (N_6463,N_5514,N_5980);
and U6464 (N_6464,N_5871,N_5423);
xnor U6465 (N_6465,N_5595,N_5954);
or U6466 (N_6466,N_5969,N_5830);
nor U6467 (N_6467,N_5747,N_5713);
and U6468 (N_6468,N_5524,N_5753);
xnor U6469 (N_6469,N_5836,N_5985);
xnor U6470 (N_6470,N_5861,N_5412);
nor U6471 (N_6471,N_5823,N_5416);
or U6472 (N_6472,N_5890,N_5658);
or U6473 (N_6473,N_5577,N_5769);
nand U6474 (N_6474,N_5422,N_5898);
xnor U6475 (N_6475,N_5646,N_5846);
xor U6476 (N_6476,N_5557,N_5438);
nand U6477 (N_6477,N_5609,N_5962);
nor U6478 (N_6478,N_5667,N_5521);
nand U6479 (N_6479,N_5503,N_5529);
nand U6480 (N_6480,N_5424,N_5852);
and U6481 (N_6481,N_5644,N_5886);
nand U6482 (N_6482,N_5821,N_5963);
nor U6483 (N_6483,N_5568,N_5622);
nor U6484 (N_6484,N_5594,N_5712);
or U6485 (N_6485,N_5548,N_5418);
xnor U6486 (N_6486,N_5448,N_5450);
nand U6487 (N_6487,N_5805,N_5708);
or U6488 (N_6488,N_5854,N_5570);
nand U6489 (N_6489,N_5580,N_5652);
nand U6490 (N_6490,N_5815,N_5905);
and U6491 (N_6491,N_5736,N_5741);
and U6492 (N_6492,N_5611,N_5840);
xor U6493 (N_6493,N_5968,N_5690);
and U6494 (N_6494,N_5403,N_5672);
nor U6495 (N_6495,N_5946,N_5957);
xor U6496 (N_6496,N_5625,N_5986);
xnor U6497 (N_6497,N_5926,N_5685);
xor U6498 (N_6498,N_5787,N_5575);
or U6499 (N_6499,N_5593,N_5925);
xor U6500 (N_6500,N_5616,N_5810);
xor U6501 (N_6501,N_5942,N_5792);
and U6502 (N_6502,N_5502,N_5574);
nor U6503 (N_6503,N_5597,N_5761);
and U6504 (N_6504,N_5723,N_5730);
nor U6505 (N_6505,N_5924,N_5755);
and U6506 (N_6506,N_5736,N_5505);
nand U6507 (N_6507,N_5739,N_5621);
or U6508 (N_6508,N_5463,N_5772);
xor U6509 (N_6509,N_5745,N_5434);
and U6510 (N_6510,N_5427,N_5949);
nor U6511 (N_6511,N_5435,N_5850);
nand U6512 (N_6512,N_5425,N_5731);
nor U6513 (N_6513,N_5413,N_5954);
and U6514 (N_6514,N_5608,N_5585);
and U6515 (N_6515,N_5452,N_5688);
nor U6516 (N_6516,N_5817,N_5880);
nand U6517 (N_6517,N_5640,N_5689);
and U6518 (N_6518,N_5662,N_5614);
nand U6519 (N_6519,N_5645,N_5415);
nor U6520 (N_6520,N_5640,N_5860);
xnor U6521 (N_6521,N_5685,N_5845);
or U6522 (N_6522,N_5931,N_5952);
or U6523 (N_6523,N_5839,N_5405);
nor U6524 (N_6524,N_5964,N_5735);
xor U6525 (N_6525,N_5568,N_5433);
nand U6526 (N_6526,N_5925,N_5439);
or U6527 (N_6527,N_5494,N_5782);
nor U6528 (N_6528,N_5518,N_5465);
xnor U6529 (N_6529,N_5818,N_5834);
nor U6530 (N_6530,N_5549,N_5496);
nand U6531 (N_6531,N_5810,N_5719);
nand U6532 (N_6532,N_5514,N_5879);
nand U6533 (N_6533,N_5956,N_5409);
nand U6534 (N_6534,N_5456,N_5748);
nand U6535 (N_6535,N_5901,N_5504);
nand U6536 (N_6536,N_5956,N_5404);
nand U6537 (N_6537,N_5770,N_5901);
nand U6538 (N_6538,N_5464,N_5631);
or U6539 (N_6539,N_5447,N_5483);
and U6540 (N_6540,N_5816,N_5614);
nand U6541 (N_6541,N_5913,N_5719);
or U6542 (N_6542,N_5401,N_5433);
and U6543 (N_6543,N_5540,N_5835);
or U6544 (N_6544,N_5858,N_5642);
nand U6545 (N_6545,N_5836,N_5782);
xnor U6546 (N_6546,N_5656,N_5867);
and U6547 (N_6547,N_5866,N_5696);
nor U6548 (N_6548,N_5615,N_5990);
nor U6549 (N_6549,N_5686,N_5579);
or U6550 (N_6550,N_5781,N_5520);
or U6551 (N_6551,N_5683,N_5780);
nand U6552 (N_6552,N_5972,N_5692);
xor U6553 (N_6553,N_5947,N_5942);
or U6554 (N_6554,N_5725,N_5655);
and U6555 (N_6555,N_5707,N_5906);
and U6556 (N_6556,N_5763,N_5503);
and U6557 (N_6557,N_5899,N_5871);
xnor U6558 (N_6558,N_5854,N_5610);
xor U6559 (N_6559,N_5424,N_5719);
nor U6560 (N_6560,N_5651,N_5691);
nand U6561 (N_6561,N_5598,N_5916);
nor U6562 (N_6562,N_5991,N_5552);
xnor U6563 (N_6563,N_5909,N_5840);
nor U6564 (N_6564,N_5814,N_5801);
nand U6565 (N_6565,N_5432,N_5635);
and U6566 (N_6566,N_5836,N_5523);
xor U6567 (N_6567,N_5645,N_5874);
nor U6568 (N_6568,N_5757,N_5547);
nand U6569 (N_6569,N_5971,N_5535);
and U6570 (N_6570,N_5642,N_5935);
xor U6571 (N_6571,N_5784,N_5453);
xor U6572 (N_6572,N_5985,N_5853);
xnor U6573 (N_6573,N_5917,N_5673);
and U6574 (N_6574,N_5494,N_5698);
xnor U6575 (N_6575,N_5714,N_5991);
xnor U6576 (N_6576,N_5616,N_5473);
or U6577 (N_6577,N_5909,N_5983);
and U6578 (N_6578,N_5889,N_5717);
or U6579 (N_6579,N_5880,N_5579);
or U6580 (N_6580,N_5881,N_5828);
or U6581 (N_6581,N_5766,N_5886);
and U6582 (N_6582,N_5702,N_5978);
xor U6583 (N_6583,N_5437,N_5622);
or U6584 (N_6584,N_5454,N_5810);
nand U6585 (N_6585,N_5695,N_5692);
nor U6586 (N_6586,N_5912,N_5496);
and U6587 (N_6587,N_5927,N_5408);
xor U6588 (N_6588,N_5897,N_5694);
or U6589 (N_6589,N_5676,N_5915);
nand U6590 (N_6590,N_5676,N_5562);
xnor U6591 (N_6591,N_5904,N_5706);
nor U6592 (N_6592,N_5580,N_5632);
nor U6593 (N_6593,N_5910,N_5944);
nor U6594 (N_6594,N_5680,N_5642);
or U6595 (N_6595,N_5411,N_5881);
nand U6596 (N_6596,N_5553,N_5420);
and U6597 (N_6597,N_5799,N_5504);
xnor U6598 (N_6598,N_5697,N_5506);
nor U6599 (N_6599,N_5880,N_5528);
or U6600 (N_6600,N_6269,N_6292);
nand U6601 (N_6601,N_6094,N_6090);
nor U6602 (N_6602,N_6405,N_6215);
xor U6603 (N_6603,N_6080,N_6125);
or U6604 (N_6604,N_6183,N_6501);
xnor U6605 (N_6605,N_6087,N_6120);
nand U6606 (N_6606,N_6345,N_6192);
xnor U6607 (N_6607,N_6248,N_6377);
nor U6608 (N_6608,N_6329,N_6239);
xnor U6609 (N_6609,N_6364,N_6028);
or U6610 (N_6610,N_6427,N_6394);
nor U6611 (N_6611,N_6121,N_6399);
xnor U6612 (N_6612,N_6548,N_6092);
or U6613 (N_6613,N_6016,N_6164);
or U6614 (N_6614,N_6050,N_6168);
or U6615 (N_6615,N_6521,N_6596);
xor U6616 (N_6616,N_6440,N_6065);
or U6617 (N_6617,N_6519,N_6115);
xnor U6618 (N_6618,N_6277,N_6064);
xnor U6619 (N_6619,N_6063,N_6367);
xor U6620 (N_6620,N_6328,N_6268);
xor U6621 (N_6621,N_6251,N_6363);
and U6622 (N_6622,N_6294,N_6143);
nand U6623 (N_6623,N_6321,N_6347);
nand U6624 (N_6624,N_6078,N_6332);
or U6625 (N_6625,N_6290,N_6571);
nand U6626 (N_6626,N_6299,N_6151);
nor U6627 (N_6627,N_6003,N_6441);
xnor U6628 (N_6628,N_6395,N_6306);
or U6629 (N_6629,N_6376,N_6576);
or U6630 (N_6630,N_6033,N_6132);
xor U6631 (N_6631,N_6404,N_6100);
and U6632 (N_6632,N_6538,N_6022);
nand U6633 (N_6633,N_6463,N_6040);
xnor U6634 (N_6634,N_6017,N_6498);
nand U6635 (N_6635,N_6263,N_6072);
or U6636 (N_6636,N_6439,N_6049);
or U6637 (N_6637,N_6230,N_6195);
and U6638 (N_6638,N_6134,N_6560);
xor U6639 (N_6639,N_6265,N_6129);
and U6640 (N_6640,N_6423,N_6071);
nor U6641 (N_6641,N_6341,N_6213);
and U6642 (N_6642,N_6414,N_6553);
nand U6643 (N_6643,N_6160,N_6169);
or U6644 (N_6644,N_6261,N_6459);
and U6645 (N_6645,N_6371,N_6079);
or U6646 (N_6646,N_6336,N_6275);
nor U6647 (N_6647,N_6450,N_6549);
xnor U6648 (N_6648,N_6199,N_6447);
or U6649 (N_6649,N_6211,N_6180);
xor U6650 (N_6650,N_6550,N_6235);
nor U6651 (N_6651,N_6485,N_6006);
nand U6652 (N_6652,N_6547,N_6042);
xor U6653 (N_6653,N_6297,N_6249);
nor U6654 (N_6654,N_6231,N_6518);
or U6655 (N_6655,N_6597,N_6257);
xnor U6656 (N_6656,N_6303,N_6153);
and U6657 (N_6657,N_6055,N_6526);
xor U6658 (N_6658,N_6021,N_6014);
xor U6659 (N_6659,N_6047,N_6599);
and U6660 (N_6660,N_6334,N_6059);
nand U6661 (N_6661,N_6166,N_6044);
nor U6662 (N_6662,N_6242,N_6529);
or U6663 (N_6663,N_6130,N_6256);
and U6664 (N_6664,N_6206,N_6552);
nor U6665 (N_6665,N_6219,N_6058);
and U6666 (N_6666,N_6496,N_6315);
nand U6667 (N_6667,N_6267,N_6031);
nor U6668 (N_6668,N_6537,N_6456);
xor U6669 (N_6669,N_6171,N_6532);
and U6670 (N_6670,N_6146,N_6595);
xnor U6671 (N_6671,N_6449,N_6343);
nand U6672 (N_6672,N_6259,N_6075);
nand U6673 (N_6673,N_6309,N_6389);
and U6674 (N_6674,N_6188,N_6305);
and U6675 (N_6675,N_6051,N_6073);
nand U6676 (N_6676,N_6531,N_6454);
and U6677 (N_6677,N_6477,N_6539);
or U6678 (N_6678,N_6159,N_6530);
nor U6679 (N_6679,N_6380,N_6438);
nand U6680 (N_6680,N_6346,N_6127);
xor U6681 (N_6681,N_6264,N_6397);
or U6682 (N_6682,N_6535,N_6013);
or U6683 (N_6683,N_6434,N_6417);
and U6684 (N_6684,N_6430,N_6509);
and U6685 (N_6685,N_6296,N_6157);
nand U6686 (N_6686,N_6546,N_6262);
nor U6687 (N_6687,N_6588,N_6109);
nor U6688 (N_6688,N_6032,N_6384);
xnor U6689 (N_6689,N_6174,N_6322);
or U6690 (N_6690,N_6173,N_6407);
or U6691 (N_6691,N_6133,N_6279);
nand U6692 (N_6692,N_6103,N_6005);
or U6693 (N_6693,N_6077,N_6435);
xor U6694 (N_6694,N_6422,N_6339);
xor U6695 (N_6695,N_6551,N_6524);
nor U6696 (N_6696,N_6432,N_6409);
nand U6697 (N_6697,N_6489,N_6245);
or U6698 (N_6698,N_6375,N_6408);
nor U6699 (N_6699,N_6291,N_6392);
xnor U6700 (N_6700,N_6184,N_6254);
nand U6701 (N_6701,N_6220,N_6563);
xor U6702 (N_6702,N_6431,N_6577);
or U6703 (N_6703,N_6383,N_6554);
xnor U6704 (N_6704,N_6098,N_6562);
or U6705 (N_6705,N_6210,N_6196);
nand U6706 (N_6706,N_6070,N_6411);
or U6707 (N_6707,N_6214,N_6243);
and U6708 (N_6708,N_6372,N_6379);
and U6709 (N_6709,N_6591,N_6015);
nor U6710 (N_6710,N_6574,N_6410);
nor U6711 (N_6711,N_6301,N_6507);
and U6712 (N_6712,N_6302,N_6488);
and U6713 (N_6713,N_6359,N_6057);
nor U6714 (N_6714,N_6444,N_6106);
nor U6715 (N_6715,N_6118,N_6038);
nor U6716 (N_6716,N_6490,N_6253);
nand U6717 (N_6717,N_6217,N_6114);
and U6718 (N_6718,N_6326,N_6340);
or U6719 (N_6719,N_6009,N_6515);
nor U6720 (N_6720,N_6240,N_6478);
nand U6721 (N_6721,N_6579,N_6473);
or U6722 (N_6722,N_6419,N_6216);
nor U6723 (N_6723,N_6209,N_6433);
and U6724 (N_6724,N_6357,N_6027);
nand U6725 (N_6725,N_6402,N_6154);
nand U6726 (N_6726,N_6493,N_6398);
xor U6727 (N_6727,N_6482,N_6293);
or U6728 (N_6728,N_6274,N_6429);
and U6729 (N_6729,N_6483,N_6298);
nand U6730 (N_6730,N_6580,N_6572);
or U6731 (N_6731,N_6481,N_6480);
nor U6732 (N_6732,N_6084,N_6234);
xor U6733 (N_6733,N_6415,N_6469);
or U6734 (N_6734,N_6101,N_6320);
and U6735 (N_6735,N_6095,N_6052);
and U6736 (N_6736,N_6587,N_6226);
nand U6737 (N_6737,N_6452,N_6557);
nor U6738 (N_6738,N_6285,N_6112);
nand U6739 (N_6739,N_6185,N_6246);
or U6740 (N_6740,N_6286,N_6083);
and U6741 (N_6741,N_6228,N_6337);
or U6742 (N_6742,N_6138,N_6499);
nand U6743 (N_6743,N_6324,N_6108);
xor U6744 (N_6744,N_6559,N_6594);
nand U6745 (N_6745,N_6018,N_6494);
nand U6746 (N_6746,N_6360,N_6351);
xnor U6747 (N_6747,N_6037,N_6026);
and U6748 (N_6748,N_6443,N_6569);
xor U6749 (N_6749,N_6053,N_6179);
nand U6750 (N_6750,N_6190,N_6500);
xor U6751 (N_6751,N_6505,N_6012);
xor U6752 (N_6752,N_6102,N_6474);
nor U6753 (N_6753,N_6270,N_6046);
and U6754 (N_6754,N_6391,N_6224);
or U6755 (N_6755,N_6119,N_6203);
nor U6756 (N_6756,N_6445,N_6522);
nand U6757 (N_6757,N_6155,N_6247);
and U6758 (N_6758,N_6034,N_6178);
nand U6759 (N_6759,N_6545,N_6283);
and U6760 (N_6760,N_6568,N_6487);
nor U6761 (N_6761,N_6222,N_6428);
xor U6762 (N_6762,N_6388,N_6314);
nand U6763 (N_6763,N_6089,N_6139);
nand U6764 (N_6764,N_6140,N_6163);
nor U6765 (N_6765,N_6227,N_6378);
xor U6766 (N_6766,N_6122,N_6289);
nor U6767 (N_6767,N_6317,N_6088);
xnor U6768 (N_6768,N_6370,N_6528);
nand U6769 (N_6769,N_6510,N_6204);
or U6770 (N_6770,N_6066,N_6497);
xor U6771 (N_6771,N_6479,N_6177);
xnor U6772 (N_6772,N_6491,N_6096);
xor U6773 (N_6773,N_6202,N_6421);
xnor U6774 (N_6774,N_6319,N_6255);
nor U6775 (N_6775,N_6312,N_6374);
and U6776 (N_6776,N_6205,N_6288);
xnor U6777 (N_6777,N_6416,N_6131);
xnor U6778 (N_6778,N_6401,N_6544);
nand U6779 (N_6779,N_6221,N_6011);
xor U6780 (N_6780,N_6123,N_6460);
nand U6781 (N_6781,N_6502,N_6271);
or U6782 (N_6782,N_6516,N_6187);
xor U6783 (N_6783,N_6197,N_6091);
nand U6784 (N_6784,N_6250,N_6193);
or U6785 (N_6785,N_6582,N_6476);
nor U6786 (N_6786,N_6584,N_6467);
or U6787 (N_6787,N_6097,N_6307);
or U6788 (N_6788,N_6369,N_6523);
nor U6789 (N_6789,N_6280,N_6461);
xor U6790 (N_6790,N_6426,N_6311);
or U6791 (N_6791,N_6495,N_6135);
nor U6792 (N_6792,N_6471,N_6331);
or U6793 (N_6793,N_6074,N_6000);
or U6794 (N_6794,N_6152,N_6273);
and U6795 (N_6795,N_6508,N_6472);
nand U6796 (N_6796,N_6099,N_6503);
nor U6797 (N_6797,N_6442,N_6313);
or U6798 (N_6798,N_6350,N_6578);
nand U6799 (N_6799,N_6464,N_6468);
and U6800 (N_6800,N_6327,N_6069);
nand U6801 (N_6801,N_6586,N_6534);
and U6802 (N_6802,N_6284,N_6212);
xor U6803 (N_6803,N_6393,N_6276);
and U6804 (N_6804,N_6382,N_6540);
or U6805 (N_6805,N_6282,N_6258);
nand U6806 (N_6806,N_6186,N_6024);
xnor U6807 (N_6807,N_6525,N_6082);
nor U6808 (N_6808,N_6161,N_6054);
or U6809 (N_6809,N_6086,N_6353);
or U6810 (N_6810,N_6381,N_6036);
nand U6811 (N_6811,N_6573,N_6061);
or U6812 (N_6812,N_6373,N_6300);
nand U6813 (N_6813,N_6541,N_6107);
xnor U6814 (N_6814,N_6451,N_6175);
xor U6815 (N_6815,N_6278,N_6223);
and U6816 (N_6816,N_6342,N_6325);
nor U6817 (N_6817,N_6062,N_6366);
nor U6818 (N_6818,N_6150,N_6542);
xor U6819 (N_6819,N_6076,N_6352);
xor U6820 (N_6820,N_6330,N_6144);
and U6821 (N_6821,N_6182,N_6260);
xor U6822 (N_6822,N_6295,N_6425);
or U6823 (N_6823,N_6565,N_6002);
and U6824 (N_6824,N_6176,N_6007);
and U6825 (N_6825,N_6349,N_6218);
nand U6826 (N_6826,N_6465,N_6068);
and U6827 (N_6827,N_6145,N_6111);
nand U6828 (N_6828,N_6592,N_6358);
or U6829 (N_6829,N_6043,N_6010);
nand U6830 (N_6830,N_6385,N_6492);
xor U6831 (N_6831,N_6041,N_6067);
nand U6832 (N_6832,N_6520,N_6462);
nor U6833 (N_6833,N_6170,N_6232);
and U6834 (N_6834,N_6335,N_6148);
xnor U6835 (N_6835,N_6593,N_6566);
xor U6836 (N_6836,N_6413,N_6241);
xor U6837 (N_6837,N_6004,N_6589);
nor U6838 (N_6838,N_6172,N_6244);
xor U6839 (N_6839,N_6048,N_6019);
or U6840 (N_6840,N_6035,N_6412);
or U6841 (N_6841,N_6287,N_6181);
nor U6842 (N_6842,N_6475,N_6400);
nor U6843 (N_6843,N_6142,N_6453);
nor U6844 (N_6844,N_6020,N_6201);
nor U6845 (N_6845,N_6128,N_6355);
nand U6846 (N_6846,N_6470,N_6598);
or U6847 (N_6847,N_6198,N_6167);
xnor U6848 (N_6848,N_6455,N_6238);
or U6849 (N_6849,N_6390,N_6001);
nor U6850 (N_6850,N_6564,N_6030);
and U6851 (N_6851,N_6126,N_6446);
nand U6852 (N_6852,N_6008,N_6533);
nand U6853 (N_6853,N_6506,N_6581);
or U6854 (N_6854,N_6418,N_6513);
xnor U6855 (N_6855,N_6361,N_6396);
nor U6856 (N_6856,N_6527,N_6457);
and U6857 (N_6857,N_6029,N_6200);
or U6858 (N_6858,N_6272,N_6344);
nand U6859 (N_6859,N_6104,N_6466);
nand U6860 (N_6860,N_6354,N_6437);
or U6861 (N_6861,N_6060,N_6333);
nor U6862 (N_6862,N_6512,N_6039);
or U6863 (N_6863,N_6081,N_6458);
or U6864 (N_6864,N_6484,N_6165);
nor U6865 (N_6865,N_6567,N_6025);
xnor U6866 (N_6866,N_6093,N_6556);
nor U6867 (N_6867,N_6045,N_6448);
or U6868 (N_6868,N_6348,N_6308);
nand U6869 (N_6869,N_6194,N_6229);
or U6870 (N_6870,N_6517,N_6561);
or U6871 (N_6871,N_6141,N_6124);
and U6872 (N_6872,N_6158,N_6252);
xnor U6873 (N_6873,N_6225,N_6555);
xnor U6874 (N_6874,N_6310,N_6583);
and U6875 (N_6875,N_6585,N_6117);
nor U6876 (N_6876,N_6420,N_6436);
nand U6877 (N_6877,N_6162,N_6136);
and U6878 (N_6878,N_6323,N_6110);
xnor U6879 (N_6879,N_6116,N_6316);
nor U6880 (N_6880,N_6207,N_6362);
or U6881 (N_6881,N_6156,N_6266);
nand U6882 (N_6882,N_6365,N_6543);
or U6883 (N_6883,N_6368,N_6318);
and U6884 (N_6884,N_6424,N_6304);
nor U6885 (N_6885,N_6189,N_6237);
nand U6886 (N_6886,N_6281,N_6147);
nor U6887 (N_6887,N_6105,N_6233);
nor U6888 (N_6888,N_6590,N_6504);
or U6889 (N_6889,N_6387,N_6149);
or U6890 (N_6890,N_6403,N_6558);
xor U6891 (N_6891,N_6486,N_6113);
nand U6892 (N_6892,N_6511,N_6236);
nand U6893 (N_6893,N_6536,N_6208);
nor U6894 (N_6894,N_6023,N_6137);
or U6895 (N_6895,N_6085,N_6575);
xor U6896 (N_6896,N_6514,N_6386);
xnor U6897 (N_6897,N_6191,N_6338);
nand U6898 (N_6898,N_6570,N_6406);
nand U6899 (N_6899,N_6356,N_6056);
and U6900 (N_6900,N_6599,N_6375);
xor U6901 (N_6901,N_6097,N_6271);
or U6902 (N_6902,N_6369,N_6349);
nor U6903 (N_6903,N_6221,N_6068);
and U6904 (N_6904,N_6411,N_6500);
nand U6905 (N_6905,N_6070,N_6233);
xnor U6906 (N_6906,N_6582,N_6434);
xnor U6907 (N_6907,N_6599,N_6344);
xnor U6908 (N_6908,N_6129,N_6488);
and U6909 (N_6909,N_6072,N_6325);
and U6910 (N_6910,N_6262,N_6573);
or U6911 (N_6911,N_6386,N_6453);
and U6912 (N_6912,N_6448,N_6247);
and U6913 (N_6913,N_6566,N_6351);
and U6914 (N_6914,N_6475,N_6007);
or U6915 (N_6915,N_6350,N_6042);
nor U6916 (N_6916,N_6070,N_6244);
or U6917 (N_6917,N_6493,N_6033);
nand U6918 (N_6918,N_6209,N_6121);
nand U6919 (N_6919,N_6095,N_6504);
nand U6920 (N_6920,N_6478,N_6156);
and U6921 (N_6921,N_6143,N_6225);
nand U6922 (N_6922,N_6286,N_6329);
xnor U6923 (N_6923,N_6445,N_6341);
or U6924 (N_6924,N_6538,N_6029);
xnor U6925 (N_6925,N_6424,N_6008);
xor U6926 (N_6926,N_6174,N_6222);
xnor U6927 (N_6927,N_6046,N_6174);
xnor U6928 (N_6928,N_6194,N_6071);
or U6929 (N_6929,N_6493,N_6512);
nor U6930 (N_6930,N_6001,N_6341);
xor U6931 (N_6931,N_6596,N_6173);
nor U6932 (N_6932,N_6316,N_6534);
and U6933 (N_6933,N_6308,N_6179);
nor U6934 (N_6934,N_6574,N_6466);
or U6935 (N_6935,N_6428,N_6079);
and U6936 (N_6936,N_6048,N_6265);
nand U6937 (N_6937,N_6530,N_6031);
and U6938 (N_6938,N_6416,N_6553);
or U6939 (N_6939,N_6182,N_6084);
and U6940 (N_6940,N_6474,N_6124);
nor U6941 (N_6941,N_6088,N_6476);
xnor U6942 (N_6942,N_6165,N_6391);
nand U6943 (N_6943,N_6370,N_6188);
nand U6944 (N_6944,N_6098,N_6277);
xor U6945 (N_6945,N_6167,N_6140);
nand U6946 (N_6946,N_6006,N_6120);
and U6947 (N_6947,N_6165,N_6140);
nand U6948 (N_6948,N_6486,N_6215);
or U6949 (N_6949,N_6019,N_6025);
nor U6950 (N_6950,N_6130,N_6028);
xor U6951 (N_6951,N_6293,N_6216);
xnor U6952 (N_6952,N_6076,N_6348);
nor U6953 (N_6953,N_6413,N_6438);
and U6954 (N_6954,N_6151,N_6285);
or U6955 (N_6955,N_6222,N_6245);
nor U6956 (N_6956,N_6297,N_6131);
nor U6957 (N_6957,N_6024,N_6234);
nand U6958 (N_6958,N_6510,N_6577);
or U6959 (N_6959,N_6195,N_6280);
nor U6960 (N_6960,N_6491,N_6372);
xor U6961 (N_6961,N_6278,N_6109);
xnor U6962 (N_6962,N_6091,N_6229);
nor U6963 (N_6963,N_6257,N_6076);
or U6964 (N_6964,N_6222,N_6322);
xnor U6965 (N_6965,N_6354,N_6564);
and U6966 (N_6966,N_6272,N_6030);
and U6967 (N_6967,N_6329,N_6291);
nand U6968 (N_6968,N_6403,N_6179);
or U6969 (N_6969,N_6556,N_6124);
xor U6970 (N_6970,N_6106,N_6429);
nand U6971 (N_6971,N_6553,N_6316);
or U6972 (N_6972,N_6554,N_6242);
nand U6973 (N_6973,N_6203,N_6581);
nand U6974 (N_6974,N_6099,N_6394);
nor U6975 (N_6975,N_6278,N_6188);
nand U6976 (N_6976,N_6532,N_6584);
and U6977 (N_6977,N_6069,N_6575);
and U6978 (N_6978,N_6251,N_6460);
nand U6979 (N_6979,N_6055,N_6436);
xor U6980 (N_6980,N_6381,N_6551);
nor U6981 (N_6981,N_6520,N_6432);
or U6982 (N_6982,N_6169,N_6224);
and U6983 (N_6983,N_6224,N_6485);
xor U6984 (N_6984,N_6381,N_6429);
nand U6985 (N_6985,N_6449,N_6318);
or U6986 (N_6986,N_6352,N_6110);
and U6987 (N_6987,N_6035,N_6426);
nor U6988 (N_6988,N_6522,N_6018);
nor U6989 (N_6989,N_6359,N_6064);
xor U6990 (N_6990,N_6168,N_6015);
nand U6991 (N_6991,N_6248,N_6598);
or U6992 (N_6992,N_6103,N_6379);
xor U6993 (N_6993,N_6201,N_6532);
and U6994 (N_6994,N_6484,N_6302);
nand U6995 (N_6995,N_6406,N_6599);
nor U6996 (N_6996,N_6492,N_6250);
nand U6997 (N_6997,N_6297,N_6364);
and U6998 (N_6998,N_6082,N_6232);
xnor U6999 (N_6999,N_6264,N_6411);
nor U7000 (N_7000,N_6343,N_6242);
xnor U7001 (N_7001,N_6440,N_6130);
xor U7002 (N_7002,N_6432,N_6593);
nand U7003 (N_7003,N_6454,N_6383);
and U7004 (N_7004,N_6277,N_6063);
and U7005 (N_7005,N_6510,N_6480);
nand U7006 (N_7006,N_6239,N_6348);
xnor U7007 (N_7007,N_6114,N_6091);
and U7008 (N_7008,N_6209,N_6102);
nand U7009 (N_7009,N_6086,N_6408);
nand U7010 (N_7010,N_6466,N_6100);
or U7011 (N_7011,N_6482,N_6337);
and U7012 (N_7012,N_6408,N_6576);
nor U7013 (N_7013,N_6368,N_6567);
or U7014 (N_7014,N_6235,N_6218);
xor U7015 (N_7015,N_6103,N_6186);
or U7016 (N_7016,N_6437,N_6179);
nor U7017 (N_7017,N_6454,N_6542);
nand U7018 (N_7018,N_6244,N_6087);
xnor U7019 (N_7019,N_6561,N_6210);
nand U7020 (N_7020,N_6025,N_6117);
nand U7021 (N_7021,N_6072,N_6314);
xor U7022 (N_7022,N_6284,N_6592);
nor U7023 (N_7023,N_6001,N_6025);
nand U7024 (N_7024,N_6385,N_6235);
or U7025 (N_7025,N_6129,N_6492);
or U7026 (N_7026,N_6268,N_6410);
nand U7027 (N_7027,N_6333,N_6436);
xor U7028 (N_7028,N_6045,N_6536);
and U7029 (N_7029,N_6124,N_6397);
nor U7030 (N_7030,N_6511,N_6071);
nand U7031 (N_7031,N_6053,N_6335);
nand U7032 (N_7032,N_6050,N_6550);
and U7033 (N_7033,N_6267,N_6114);
and U7034 (N_7034,N_6208,N_6044);
xnor U7035 (N_7035,N_6049,N_6205);
nand U7036 (N_7036,N_6404,N_6024);
nor U7037 (N_7037,N_6248,N_6164);
or U7038 (N_7038,N_6434,N_6196);
or U7039 (N_7039,N_6584,N_6361);
xnor U7040 (N_7040,N_6219,N_6231);
or U7041 (N_7041,N_6085,N_6000);
nor U7042 (N_7042,N_6151,N_6074);
nand U7043 (N_7043,N_6285,N_6356);
nor U7044 (N_7044,N_6173,N_6336);
or U7045 (N_7045,N_6571,N_6319);
and U7046 (N_7046,N_6050,N_6443);
nor U7047 (N_7047,N_6569,N_6429);
nand U7048 (N_7048,N_6037,N_6134);
or U7049 (N_7049,N_6051,N_6180);
nor U7050 (N_7050,N_6379,N_6071);
nand U7051 (N_7051,N_6261,N_6387);
or U7052 (N_7052,N_6522,N_6521);
nor U7053 (N_7053,N_6426,N_6531);
xnor U7054 (N_7054,N_6103,N_6117);
and U7055 (N_7055,N_6102,N_6499);
xor U7056 (N_7056,N_6458,N_6485);
nor U7057 (N_7057,N_6275,N_6215);
and U7058 (N_7058,N_6596,N_6555);
xor U7059 (N_7059,N_6012,N_6467);
nand U7060 (N_7060,N_6312,N_6013);
or U7061 (N_7061,N_6299,N_6515);
nand U7062 (N_7062,N_6052,N_6030);
nand U7063 (N_7063,N_6249,N_6171);
nand U7064 (N_7064,N_6491,N_6172);
or U7065 (N_7065,N_6038,N_6095);
nor U7066 (N_7066,N_6474,N_6339);
nand U7067 (N_7067,N_6103,N_6279);
and U7068 (N_7068,N_6025,N_6129);
nand U7069 (N_7069,N_6441,N_6310);
nor U7070 (N_7070,N_6333,N_6057);
nand U7071 (N_7071,N_6169,N_6431);
nor U7072 (N_7072,N_6282,N_6444);
nand U7073 (N_7073,N_6444,N_6220);
or U7074 (N_7074,N_6375,N_6217);
nand U7075 (N_7075,N_6124,N_6574);
nor U7076 (N_7076,N_6156,N_6436);
and U7077 (N_7077,N_6120,N_6113);
nor U7078 (N_7078,N_6553,N_6110);
nor U7079 (N_7079,N_6025,N_6409);
or U7080 (N_7080,N_6341,N_6386);
nor U7081 (N_7081,N_6234,N_6517);
xor U7082 (N_7082,N_6244,N_6429);
and U7083 (N_7083,N_6219,N_6509);
nand U7084 (N_7084,N_6595,N_6325);
nor U7085 (N_7085,N_6247,N_6489);
and U7086 (N_7086,N_6334,N_6187);
and U7087 (N_7087,N_6507,N_6070);
nor U7088 (N_7088,N_6164,N_6367);
nor U7089 (N_7089,N_6007,N_6067);
nor U7090 (N_7090,N_6504,N_6094);
xor U7091 (N_7091,N_6371,N_6045);
nor U7092 (N_7092,N_6177,N_6151);
or U7093 (N_7093,N_6146,N_6581);
nand U7094 (N_7094,N_6093,N_6557);
nor U7095 (N_7095,N_6302,N_6584);
nand U7096 (N_7096,N_6440,N_6136);
and U7097 (N_7097,N_6333,N_6446);
nor U7098 (N_7098,N_6488,N_6025);
xnor U7099 (N_7099,N_6008,N_6119);
and U7100 (N_7100,N_6176,N_6361);
or U7101 (N_7101,N_6145,N_6213);
nor U7102 (N_7102,N_6298,N_6017);
and U7103 (N_7103,N_6253,N_6208);
nor U7104 (N_7104,N_6253,N_6197);
or U7105 (N_7105,N_6151,N_6222);
and U7106 (N_7106,N_6395,N_6147);
and U7107 (N_7107,N_6146,N_6379);
xor U7108 (N_7108,N_6301,N_6175);
xor U7109 (N_7109,N_6459,N_6552);
xor U7110 (N_7110,N_6200,N_6298);
or U7111 (N_7111,N_6000,N_6135);
and U7112 (N_7112,N_6091,N_6563);
and U7113 (N_7113,N_6002,N_6490);
nor U7114 (N_7114,N_6226,N_6341);
xnor U7115 (N_7115,N_6423,N_6512);
xor U7116 (N_7116,N_6067,N_6586);
nand U7117 (N_7117,N_6237,N_6380);
xor U7118 (N_7118,N_6180,N_6542);
nor U7119 (N_7119,N_6549,N_6322);
xor U7120 (N_7120,N_6580,N_6313);
and U7121 (N_7121,N_6033,N_6276);
or U7122 (N_7122,N_6286,N_6362);
nand U7123 (N_7123,N_6484,N_6399);
xor U7124 (N_7124,N_6065,N_6533);
or U7125 (N_7125,N_6187,N_6587);
or U7126 (N_7126,N_6033,N_6570);
nor U7127 (N_7127,N_6252,N_6268);
and U7128 (N_7128,N_6536,N_6274);
or U7129 (N_7129,N_6588,N_6366);
and U7130 (N_7130,N_6527,N_6238);
or U7131 (N_7131,N_6019,N_6309);
nand U7132 (N_7132,N_6410,N_6540);
or U7133 (N_7133,N_6083,N_6529);
and U7134 (N_7134,N_6390,N_6460);
or U7135 (N_7135,N_6050,N_6394);
nand U7136 (N_7136,N_6390,N_6498);
or U7137 (N_7137,N_6135,N_6181);
or U7138 (N_7138,N_6484,N_6518);
xnor U7139 (N_7139,N_6113,N_6524);
xnor U7140 (N_7140,N_6321,N_6410);
xnor U7141 (N_7141,N_6122,N_6380);
xnor U7142 (N_7142,N_6472,N_6521);
or U7143 (N_7143,N_6267,N_6593);
nand U7144 (N_7144,N_6550,N_6080);
nor U7145 (N_7145,N_6489,N_6273);
xnor U7146 (N_7146,N_6123,N_6219);
nor U7147 (N_7147,N_6541,N_6536);
xor U7148 (N_7148,N_6278,N_6429);
nand U7149 (N_7149,N_6262,N_6496);
and U7150 (N_7150,N_6138,N_6011);
nor U7151 (N_7151,N_6342,N_6418);
or U7152 (N_7152,N_6160,N_6222);
and U7153 (N_7153,N_6288,N_6101);
and U7154 (N_7154,N_6036,N_6500);
nand U7155 (N_7155,N_6364,N_6003);
or U7156 (N_7156,N_6521,N_6152);
nand U7157 (N_7157,N_6464,N_6558);
or U7158 (N_7158,N_6482,N_6265);
nand U7159 (N_7159,N_6287,N_6379);
xnor U7160 (N_7160,N_6360,N_6264);
nor U7161 (N_7161,N_6105,N_6544);
nand U7162 (N_7162,N_6079,N_6520);
xor U7163 (N_7163,N_6265,N_6327);
xor U7164 (N_7164,N_6208,N_6362);
xor U7165 (N_7165,N_6027,N_6391);
nand U7166 (N_7166,N_6275,N_6309);
xnor U7167 (N_7167,N_6211,N_6437);
or U7168 (N_7168,N_6505,N_6134);
or U7169 (N_7169,N_6514,N_6261);
xnor U7170 (N_7170,N_6099,N_6498);
xor U7171 (N_7171,N_6476,N_6422);
or U7172 (N_7172,N_6134,N_6296);
nor U7173 (N_7173,N_6428,N_6395);
or U7174 (N_7174,N_6159,N_6427);
or U7175 (N_7175,N_6386,N_6056);
nor U7176 (N_7176,N_6368,N_6080);
xnor U7177 (N_7177,N_6476,N_6543);
or U7178 (N_7178,N_6138,N_6437);
nor U7179 (N_7179,N_6352,N_6401);
xor U7180 (N_7180,N_6102,N_6350);
nand U7181 (N_7181,N_6591,N_6257);
or U7182 (N_7182,N_6138,N_6116);
nand U7183 (N_7183,N_6135,N_6354);
xor U7184 (N_7184,N_6136,N_6255);
nor U7185 (N_7185,N_6279,N_6557);
or U7186 (N_7186,N_6263,N_6462);
or U7187 (N_7187,N_6374,N_6175);
nor U7188 (N_7188,N_6395,N_6242);
xor U7189 (N_7189,N_6154,N_6321);
xor U7190 (N_7190,N_6536,N_6393);
nand U7191 (N_7191,N_6142,N_6187);
or U7192 (N_7192,N_6095,N_6533);
nor U7193 (N_7193,N_6376,N_6284);
and U7194 (N_7194,N_6548,N_6495);
xnor U7195 (N_7195,N_6183,N_6554);
or U7196 (N_7196,N_6329,N_6004);
or U7197 (N_7197,N_6156,N_6087);
or U7198 (N_7198,N_6020,N_6268);
and U7199 (N_7199,N_6502,N_6483);
and U7200 (N_7200,N_6907,N_6629);
and U7201 (N_7201,N_6936,N_6722);
xor U7202 (N_7202,N_7192,N_6710);
nor U7203 (N_7203,N_6805,N_6918);
or U7204 (N_7204,N_7170,N_6843);
or U7205 (N_7205,N_7136,N_6715);
or U7206 (N_7206,N_6638,N_6712);
nor U7207 (N_7207,N_6892,N_6991);
nor U7208 (N_7208,N_7072,N_6724);
nand U7209 (N_7209,N_6913,N_6741);
nor U7210 (N_7210,N_6791,N_6995);
nor U7211 (N_7211,N_6611,N_7066);
xor U7212 (N_7212,N_7199,N_7169);
nor U7213 (N_7213,N_7133,N_6940);
or U7214 (N_7214,N_6957,N_7116);
nand U7215 (N_7215,N_7099,N_6975);
and U7216 (N_7216,N_7112,N_6880);
or U7217 (N_7217,N_6736,N_7076);
nand U7218 (N_7218,N_6842,N_6732);
nor U7219 (N_7219,N_6824,N_6883);
and U7220 (N_7220,N_6766,N_6993);
xnor U7221 (N_7221,N_6790,N_6604);
xnor U7222 (N_7222,N_6651,N_6989);
nor U7223 (N_7223,N_6770,N_6920);
nor U7224 (N_7224,N_6970,N_7057);
and U7225 (N_7225,N_6828,N_6941);
and U7226 (N_7226,N_6779,N_6894);
or U7227 (N_7227,N_6683,N_6745);
xnor U7228 (N_7228,N_6927,N_6674);
or U7229 (N_7229,N_6740,N_6847);
and U7230 (N_7230,N_6632,N_6665);
and U7231 (N_7231,N_6742,N_6716);
nand U7232 (N_7232,N_6752,N_6846);
xor U7233 (N_7233,N_6753,N_7115);
nand U7234 (N_7234,N_6788,N_6681);
or U7235 (N_7235,N_6614,N_7138);
nor U7236 (N_7236,N_6688,N_6747);
xor U7237 (N_7237,N_6622,N_7106);
and U7238 (N_7238,N_7001,N_6902);
nor U7239 (N_7239,N_6896,N_7068);
and U7240 (N_7240,N_7080,N_6666);
or U7241 (N_7241,N_6776,N_6690);
nor U7242 (N_7242,N_7025,N_7065);
nor U7243 (N_7243,N_6871,N_6663);
or U7244 (N_7244,N_6773,N_7155);
nor U7245 (N_7245,N_6985,N_7096);
nor U7246 (N_7246,N_6755,N_7172);
nand U7247 (N_7247,N_6679,N_6911);
xnor U7248 (N_7248,N_7189,N_7056);
xnor U7249 (N_7249,N_6998,N_6877);
or U7250 (N_7250,N_6930,N_6875);
and U7251 (N_7251,N_7043,N_6699);
nor U7252 (N_7252,N_6659,N_6744);
or U7253 (N_7253,N_6691,N_7139);
nor U7254 (N_7254,N_7154,N_6761);
and U7255 (N_7255,N_6804,N_7044);
or U7256 (N_7256,N_6785,N_6719);
or U7257 (N_7257,N_7107,N_6729);
nand U7258 (N_7258,N_7059,N_6973);
and U7259 (N_7259,N_6831,N_6780);
nor U7260 (N_7260,N_6728,N_6654);
xnor U7261 (N_7261,N_7165,N_6763);
nor U7262 (N_7262,N_6648,N_7181);
or U7263 (N_7263,N_7120,N_7013);
nand U7264 (N_7264,N_7187,N_6643);
nor U7265 (N_7265,N_6646,N_6981);
nand U7266 (N_7266,N_7020,N_6727);
nor U7267 (N_7267,N_6762,N_6713);
or U7268 (N_7268,N_6702,N_7078);
and U7269 (N_7269,N_7041,N_6774);
nand U7270 (N_7270,N_6647,N_6943);
xor U7271 (N_7271,N_6881,N_7122);
nor U7272 (N_7272,N_6898,N_7088);
nand U7273 (N_7273,N_6910,N_6900);
or U7274 (N_7274,N_6721,N_6932);
or U7275 (N_7275,N_6867,N_6882);
nor U7276 (N_7276,N_6677,N_6811);
xor U7277 (N_7277,N_6855,N_6983);
nor U7278 (N_7278,N_6864,N_6820);
and U7279 (N_7279,N_6609,N_6796);
xnor U7280 (N_7280,N_7017,N_6873);
nand U7281 (N_7281,N_7042,N_6992);
xnor U7282 (N_7282,N_6612,N_6600);
and U7283 (N_7283,N_7027,N_6678);
nand U7284 (N_7284,N_6714,N_6759);
nor U7285 (N_7285,N_7144,N_6619);
and U7286 (N_7286,N_6966,N_6778);
or U7287 (N_7287,N_7033,N_6809);
or U7288 (N_7288,N_6644,N_6825);
and U7289 (N_7289,N_6784,N_6959);
xor U7290 (N_7290,N_6947,N_6925);
and U7291 (N_7291,N_7161,N_7153);
nor U7292 (N_7292,N_7186,N_7117);
nor U7293 (N_7293,N_6968,N_7123);
nor U7294 (N_7294,N_6962,N_6834);
nor U7295 (N_7295,N_7007,N_6792);
xor U7296 (N_7296,N_7082,N_6720);
nand U7297 (N_7297,N_7190,N_7119);
nor U7298 (N_7298,N_6706,N_6851);
nor U7299 (N_7299,N_6765,N_7127);
nor U7300 (N_7300,N_6997,N_6772);
nand U7301 (N_7301,N_7178,N_7171);
and U7302 (N_7302,N_6689,N_6810);
nand U7303 (N_7303,N_7128,N_6664);
and U7304 (N_7304,N_7022,N_7104);
nand U7305 (N_7305,N_6929,N_7159);
nand U7306 (N_7306,N_7142,N_6750);
xor U7307 (N_7307,N_7074,N_6613);
nor U7308 (N_7308,N_6781,N_6803);
xnor U7309 (N_7309,N_6703,N_7048);
xor U7310 (N_7310,N_7094,N_6708);
nor U7311 (N_7311,N_7029,N_6908);
nor U7312 (N_7312,N_6960,N_6661);
and U7313 (N_7313,N_6617,N_6833);
or U7314 (N_7314,N_7150,N_7188);
or U7315 (N_7315,N_7129,N_6857);
xnor U7316 (N_7316,N_6686,N_6839);
or U7317 (N_7317,N_7184,N_7091);
and U7318 (N_7318,N_6764,N_6705);
or U7319 (N_7319,N_6606,N_7162);
nand U7320 (N_7320,N_6837,N_6829);
nor U7321 (N_7321,N_6923,N_6808);
nand U7322 (N_7322,N_7028,N_7002);
nor U7323 (N_7323,N_6931,N_7167);
and U7324 (N_7324,N_6642,N_7149);
or U7325 (N_7325,N_6967,N_6958);
and U7326 (N_7326,N_6977,N_7132);
nor U7327 (N_7327,N_6948,N_7182);
nand U7328 (N_7328,N_7004,N_7180);
or U7329 (N_7329,N_7198,N_6601);
or U7330 (N_7330,N_6668,N_6965);
and U7331 (N_7331,N_7095,N_7111);
and U7332 (N_7332,N_6826,N_6639);
nand U7333 (N_7333,N_6903,N_6869);
xnor U7334 (N_7334,N_6701,N_7008);
nand U7335 (N_7335,N_7049,N_6746);
nor U7336 (N_7336,N_6897,N_6658);
nor U7337 (N_7337,N_6982,N_6726);
or U7338 (N_7338,N_7124,N_6696);
or U7339 (N_7339,N_6856,N_7024);
nand U7340 (N_7340,N_6836,N_6933);
nor U7341 (N_7341,N_6944,N_7174);
and U7342 (N_7342,N_6636,N_7075);
xor U7343 (N_7343,N_6640,N_6733);
xnor U7344 (N_7344,N_7166,N_6969);
xor U7345 (N_7345,N_7193,N_6942);
nor U7346 (N_7346,N_6974,N_6799);
xor U7347 (N_7347,N_6602,N_7064);
and U7348 (N_7348,N_7173,N_6950);
nor U7349 (N_7349,N_6771,N_6734);
and U7350 (N_7350,N_7101,N_6980);
or U7351 (N_7351,N_7023,N_6626);
xnor U7352 (N_7352,N_6886,N_6704);
xor U7353 (N_7353,N_6783,N_6621);
or U7354 (N_7354,N_7040,N_6961);
or U7355 (N_7355,N_7121,N_6874);
nor U7356 (N_7356,N_6756,N_6650);
xnor U7357 (N_7357,N_7126,N_7021);
and U7358 (N_7358,N_6945,N_6868);
nor U7359 (N_7359,N_6812,N_7016);
or U7360 (N_7360,N_7090,N_6634);
xnor U7361 (N_7361,N_6937,N_7137);
nor U7362 (N_7362,N_6798,N_6813);
xor U7363 (N_7363,N_7191,N_6687);
nor U7364 (N_7364,N_6832,N_7110);
nor U7365 (N_7365,N_6922,N_6916);
xor U7366 (N_7366,N_6955,N_6655);
nand U7367 (N_7367,N_6939,N_6861);
nor U7368 (N_7368,N_7010,N_6858);
nand U7369 (N_7369,N_6972,N_6737);
nor U7370 (N_7370,N_7054,N_6879);
and U7371 (N_7371,N_7168,N_6624);
or U7372 (N_7372,N_6860,N_7026);
nor U7373 (N_7373,N_7047,N_7073);
xnor U7374 (N_7374,N_6794,N_7197);
xor U7375 (N_7375,N_6899,N_6641);
and U7376 (N_7376,N_6802,N_7185);
or U7377 (N_7377,N_6835,N_7005);
and U7378 (N_7378,N_6814,N_7070);
xor U7379 (N_7379,N_6738,N_7046);
xor U7380 (N_7380,N_6840,N_6618);
nor U7381 (N_7381,N_7103,N_6637);
or U7382 (N_7382,N_7079,N_6673);
nor U7383 (N_7383,N_7050,N_7194);
nand U7384 (N_7384,N_6623,N_6775);
xor U7385 (N_7385,N_7034,N_6935);
xor U7386 (N_7386,N_6928,N_7061);
nor U7387 (N_7387,N_6964,N_7031);
nor U7388 (N_7388,N_6986,N_6730);
xnor U7389 (N_7389,N_6692,N_7086);
nand U7390 (N_7390,N_7014,N_6627);
and U7391 (N_7391,N_7196,N_6633);
nor U7392 (N_7392,N_6603,N_6718);
nor U7393 (N_7393,N_6806,N_6693);
or U7394 (N_7394,N_6978,N_6996);
or U7395 (N_7395,N_6707,N_7163);
and U7396 (N_7396,N_6789,N_6676);
nand U7397 (N_7397,N_6854,N_6723);
and U7398 (N_7398,N_7164,N_7151);
nand U7399 (N_7399,N_6859,N_7018);
nand U7400 (N_7400,N_7053,N_7100);
xnor U7401 (N_7401,N_6797,N_7081);
nand U7402 (N_7402,N_6987,N_7060);
xnor U7403 (N_7403,N_7098,N_6767);
or U7404 (N_7404,N_7009,N_7030);
and U7405 (N_7405,N_6801,N_7152);
xor U7406 (N_7406,N_6953,N_7105);
and U7407 (N_7407,N_7179,N_7052);
nand U7408 (N_7408,N_6917,N_6795);
nand U7409 (N_7409,N_6615,N_6845);
xor U7410 (N_7410,N_7158,N_6865);
and U7411 (N_7411,N_6984,N_6608);
or U7412 (N_7412,N_6751,N_6862);
nand U7413 (N_7413,N_7000,N_7134);
and U7414 (N_7414,N_6616,N_6895);
or U7415 (N_7415,N_6963,N_7032);
nor U7416 (N_7416,N_6994,N_6905);
xnor U7417 (N_7417,N_6697,N_7125);
nand U7418 (N_7418,N_6946,N_6853);
or U7419 (N_7419,N_7077,N_6680);
nor U7420 (N_7420,N_6660,N_7148);
xnor U7421 (N_7421,N_7118,N_6850);
or U7422 (N_7422,N_6652,N_6669);
nand U7423 (N_7423,N_6891,N_6887);
or U7424 (N_7424,N_6876,N_7006);
and U7425 (N_7425,N_6631,N_6830);
xor U7426 (N_7426,N_6635,N_7102);
and U7427 (N_7427,N_6971,N_7195);
or U7428 (N_7428,N_6757,N_6954);
nand U7429 (N_7429,N_6934,N_7083);
and U7430 (N_7430,N_7012,N_6682);
xnor U7431 (N_7431,N_6926,N_6717);
and U7432 (N_7432,N_6988,N_6787);
or U7433 (N_7433,N_6976,N_7156);
or U7434 (N_7434,N_6844,N_6656);
or U7435 (N_7435,N_6711,N_7085);
nor U7436 (N_7436,N_6725,N_7063);
nor U7437 (N_7437,N_7051,N_6700);
nor U7438 (N_7438,N_6884,N_6786);
xor U7439 (N_7439,N_6672,N_7037);
or U7440 (N_7440,N_6657,N_7160);
nand U7441 (N_7441,N_7087,N_6956);
nor U7442 (N_7442,N_7135,N_6885);
nand U7443 (N_7443,N_6671,N_6739);
xor U7444 (N_7444,N_6754,N_6915);
and U7445 (N_7445,N_7141,N_6769);
and U7446 (N_7446,N_6760,N_6870);
xor U7447 (N_7447,N_6684,N_7093);
xnor U7448 (N_7448,N_6823,N_6695);
or U7449 (N_7449,N_6819,N_6849);
nor U7450 (N_7450,N_6889,N_6610);
or U7451 (N_7451,N_7015,N_6893);
xor U7452 (N_7452,N_7113,N_6649);
nand U7453 (N_7453,N_6605,N_6777);
nor U7454 (N_7454,N_7039,N_7084);
or U7455 (N_7455,N_6748,N_6866);
nor U7456 (N_7456,N_6951,N_7011);
nand U7457 (N_7457,N_7183,N_6888);
nor U7458 (N_7458,N_7058,N_6667);
or U7459 (N_7459,N_7036,N_7097);
and U7460 (N_7460,N_6906,N_6912);
xnor U7461 (N_7461,N_6620,N_6919);
nand U7462 (N_7462,N_6949,N_6793);
nor U7463 (N_7463,N_6743,N_6904);
or U7464 (N_7464,N_7108,N_6800);
nand U7465 (N_7465,N_6841,N_7019);
nand U7466 (N_7466,N_7114,N_6863);
nor U7467 (N_7467,N_6818,N_6782);
xnor U7468 (N_7468,N_6731,N_6924);
or U7469 (N_7469,N_6979,N_7089);
xnor U7470 (N_7470,N_7177,N_7146);
nand U7471 (N_7471,N_6952,N_6698);
or U7472 (N_7472,N_6625,N_7003);
or U7473 (N_7473,N_6838,N_7175);
or U7474 (N_7474,N_6645,N_6848);
and U7475 (N_7475,N_6914,N_6815);
nor U7476 (N_7476,N_6735,N_6901);
and U7477 (N_7477,N_7067,N_7176);
or U7478 (N_7478,N_7071,N_7130);
nand U7479 (N_7479,N_6817,N_6872);
nor U7480 (N_7480,N_7045,N_6758);
nand U7481 (N_7481,N_7062,N_6685);
nor U7482 (N_7482,N_6768,N_6827);
xnor U7483 (N_7483,N_7145,N_7140);
and U7484 (N_7484,N_6694,N_7143);
or U7485 (N_7485,N_6999,N_6749);
xnor U7486 (N_7486,N_6653,N_6852);
and U7487 (N_7487,N_6890,N_6630);
nand U7488 (N_7488,N_6709,N_7035);
xnor U7489 (N_7489,N_7038,N_6938);
and U7490 (N_7490,N_6816,N_6821);
nor U7491 (N_7491,N_7109,N_6909);
nand U7492 (N_7492,N_7131,N_7069);
nor U7493 (N_7493,N_6662,N_7147);
and U7494 (N_7494,N_6822,N_6628);
and U7495 (N_7495,N_6607,N_6807);
or U7496 (N_7496,N_6990,N_6921);
nand U7497 (N_7497,N_7157,N_6670);
and U7498 (N_7498,N_7092,N_6878);
or U7499 (N_7499,N_7055,N_6675);
or U7500 (N_7500,N_6925,N_7041);
and U7501 (N_7501,N_6721,N_7056);
or U7502 (N_7502,N_6771,N_7045);
xor U7503 (N_7503,N_6933,N_6994);
nor U7504 (N_7504,N_6997,N_7182);
xnor U7505 (N_7505,N_6720,N_7050);
xnor U7506 (N_7506,N_6879,N_6792);
nor U7507 (N_7507,N_6745,N_7117);
or U7508 (N_7508,N_6744,N_7114);
nand U7509 (N_7509,N_6856,N_7126);
nor U7510 (N_7510,N_6817,N_6675);
xor U7511 (N_7511,N_7005,N_6757);
or U7512 (N_7512,N_6935,N_7028);
nand U7513 (N_7513,N_7171,N_7118);
nor U7514 (N_7514,N_6685,N_6896);
xor U7515 (N_7515,N_6881,N_7113);
and U7516 (N_7516,N_6756,N_6620);
and U7517 (N_7517,N_6603,N_6704);
and U7518 (N_7518,N_7101,N_6738);
and U7519 (N_7519,N_6618,N_7043);
nor U7520 (N_7520,N_6702,N_7197);
xnor U7521 (N_7521,N_7058,N_6749);
or U7522 (N_7522,N_6733,N_7131);
xor U7523 (N_7523,N_6710,N_7052);
and U7524 (N_7524,N_6989,N_7080);
nand U7525 (N_7525,N_7111,N_6965);
nor U7526 (N_7526,N_6830,N_6904);
or U7527 (N_7527,N_6624,N_6660);
xnor U7528 (N_7528,N_6757,N_6621);
xor U7529 (N_7529,N_7082,N_6627);
nor U7530 (N_7530,N_6764,N_6661);
nor U7531 (N_7531,N_6707,N_6753);
and U7532 (N_7532,N_6819,N_6881);
nor U7533 (N_7533,N_6682,N_6715);
xor U7534 (N_7534,N_6862,N_6962);
nor U7535 (N_7535,N_7104,N_6726);
and U7536 (N_7536,N_7074,N_6743);
and U7537 (N_7537,N_7045,N_7194);
or U7538 (N_7538,N_6836,N_7195);
nor U7539 (N_7539,N_7174,N_7009);
nand U7540 (N_7540,N_6919,N_7092);
or U7541 (N_7541,N_6812,N_6638);
xor U7542 (N_7542,N_6756,N_6702);
or U7543 (N_7543,N_6682,N_7017);
nor U7544 (N_7544,N_6874,N_6614);
nor U7545 (N_7545,N_7021,N_7153);
xor U7546 (N_7546,N_7037,N_6792);
xnor U7547 (N_7547,N_7125,N_6648);
nand U7548 (N_7548,N_6746,N_7164);
or U7549 (N_7549,N_7034,N_6801);
xor U7550 (N_7550,N_7102,N_7004);
or U7551 (N_7551,N_6962,N_7167);
and U7552 (N_7552,N_7121,N_6967);
and U7553 (N_7553,N_7103,N_7183);
nor U7554 (N_7554,N_6808,N_7019);
nand U7555 (N_7555,N_7190,N_6995);
and U7556 (N_7556,N_6652,N_7158);
nand U7557 (N_7557,N_6792,N_7126);
xnor U7558 (N_7558,N_6752,N_7112);
nor U7559 (N_7559,N_7159,N_7174);
nor U7560 (N_7560,N_7126,N_6853);
nand U7561 (N_7561,N_7115,N_6829);
nand U7562 (N_7562,N_6874,N_7009);
nand U7563 (N_7563,N_6695,N_6984);
or U7564 (N_7564,N_7129,N_7084);
or U7565 (N_7565,N_6884,N_7105);
nand U7566 (N_7566,N_7014,N_6898);
xor U7567 (N_7567,N_6997,N_6777);
or U7568 (N_7568,N_7004,N_6817);
xnor U7569 (N_7569,N_6875,N_6988);
and U7570 (N_7570,N_6908,N_6784);
nand U7571 (N_7571,N_6779,N_7149);
or U7572 (N_7572,N_7132,N_6856);
and U7573 (N_7573,N_7105,N_6655);
and U7574 (N_7574,N_7054,N_6914);
and U7575 (N_7575,N_7017,N_7098);
or U7576 (N_7576,N_7008,N_6651);
or U7577 (N_7577,N_6789,N_6787);
nand U7578 (N_7578,N_6609,N_6648);
xnor U7579 (N_7579,N_6841,N_6834);
or U7580 (N_7580,N_6675,N_6999);
or U7581 (N_7581,N_7117,N_6983);
nor U7582 (N_7582,N_6671,N_6969);
and U7583 (N_7583,N_7179,N_7140);
xnor U7584 (N_7584,N_6950,N_7115);
and U7585 (N_7585,N_7037,N_6880);
xnor U7586 (N_7586,N_6884,N_7194);
nand U7587 (N_7587,N_7163,N_7191);
nand U7588 (N_7588,N_7111,N_7040);
nor U7589 (N_7589,N_7146,N_6615);
nor U7590 (N_7590,N_6865,N_6945);
nand U7591 (N_7591,N_7052,N_6751);
nand U7592 (N_7592,N_6686,N_6828);
nor U7593 (N_7593,N_6958,N_6740);
xor U7594 (N_7594,N_6986,N_6902);
nand U7595 (N_7595,N_6827,N_6868);
nand U7596 (N_7596,N_7185,N_6715);
or U7597 (N_7597,N_7103,N_7023);
or U7598 (N_7598,N_7075,N_6859);
and U7599 (N_7599,N_6610,N_6783);
xnor U7600 (N_7600,N_6866,N_6822);
and U7601 (N_7601,N_6746,N_6783);
xor U7602 (N_7602,N_6639,N_6981);
xnor U7603 (N_7603,N_6971,N_7157);
or U7604 (N_7604,N_6712,N_6914);
nor U7605 (N_7605,N_6860,N_7059);
xor U7606 (N_7606,N_6957,N_6781);
and U7607 (N_7607,N_6743,N_7146);
nand U7608 (N_7608,N_7072,N_6706);
or U7609 (N_7609,N_6674,N_6745);
and U7610 (N_7610,N_6946,N_7155);
and U7611 (N_7611,N_6924,N_7089);
nand U7612 (N_7612,N_6869,N_7070);
nor U7613 (N_7613,N_6927,N_6610);
nor U7614 (N_7614,N_6651,N_7165);
nor U7615 (N_7615,N_6962,N_7081);
xnor U7616 (N_7616,N_7055,N_6738);
or U7617 (N_7617,N_6907,N_7095);
and U7618 (N_7618,N_6787,N_6898);
or U7619 (N_7619,N_7019,N_7165);
xor U7620 (N_7620,N_7181,N_6858);
nand U7621 (N_7621,N_6679,N_6885);
nor U7622 (N_7622,N_6873,N_6832);
nand U7623 (N_7623,N_6637,N_7052);
xnor U7624 (N_7624,N_6657,N_7011);
and U7625 (N_7625,N_7089,N_7057);
nor U7626 (N_7626,N_6748,N_6741);
or U7627 (N_7627,N_7143,N_6771);
or U7628 (N_7628,N_6744,N_7106);
xnor U7629 (N_7629,N_6838,N_7128);
xnor U7630 (N_7630,N_6993,N_6847);
xnor U7631 (N_7631,N_6961,N_6956);
xor U7632 (N_7632,N_6731,N_6908);
or U7633 (N_7633,N_6615,N_6757);
and U7634 (N_7634,N_6643,N_7047);
xnor U7635 (N_7635,N_7067,N_7022);
nand U7636 (N_7636,N_6747,N_6888);
nand U7637 (N_7637,N_6891,N_6712);
and U7638 (N_7638,N_7190,N_6925);
or U7639 (N_7639,N_7035,N_7134);
and U7640 (N_7640,N_6753,N_7037);
and U7641 (N_7641,N_6980,N_6755);
or U7642 (N_7642,N_6808,N_7155);
nand U7643 (N_7643,N_6816,N_7133);
nor U7644 (N_7644,N_6875,N_6824);
nand U7645 (N_7645,N_7094,N_7088);
or U7646 (N_7646,N_6658,N_7143);
and U7647 (N_7647,N_6888,N_7151);
xor U7648 (N_7648,N_7177,N_7020);
nand U7649 (N_7649,N_7024,N_7048);
xor U7650 (N_7650,N_6821,N_7197);
or U7651 (N_7651,N_6719,N_6806);
xor U7652 (N_7652,N_7133,N_7175);
or U7653 (N_7653,N_6717,N_7045);
xnor U7654 (N_7654,N_6707,N_6742);
nand U7655 (N_7655,N_6610,N_6848);
nor U7656 (N_7656,N_6770,N_6677);
nand U7657 (N_7657,N_6864,N_6721);
xnor U7658 (N_7658,N_6795,N_6721);
nor U7659 (N_7659,N_6987,N_6638);
xor U7660 (N_7660,N_6637,N_6805);
or U7661 (N_7661,N_6898,N_6667);
or U7662 (N_7662,N_7181,N_6605);
nor U7663 (N_7663,N_6964,N_6607);
nand U7664 (N_7664,N_6642,N_6830);
nand U7665 (N_7665,N_7017,N_6998);
xnor U7666 (N_7666,N_7153,N_7191);
nor U7667 (N_7667,N_7143,N_7027);
and U7668 (N_7668,N_7028,N_6803);
xnor U7669 (N_7669,N_7128,N_7086);
or U7670 (N_7670,N_6905,N_6809);
or U7671 (N_7671,N_6673,N_7151);
nand U7672 (N_7672,N_7054,N_7110);
nor U7673 (N_7673,N_6677,N_7017);
nor U7674 (N_7674,N_6699,N_6811);
xnor U7675 (N_7675,N_7148,N_7005);
nand U7676 (N_7676,N_6990,N_6633);
or U7677 (N_7677,N_7068,N_7013);
and U7678 (N_7678,N_6721,N_6771);
nand U7679 (N_7679,N_7106,N_6729);
or U7680 (N_7680,N_6931,N_6969);
nor U7681 (N_7681,N_6710,N_6930);
xor U7682 (N_7682,N_6965,N_6947);
xor U7683 (N_7683,N_6957,N_6915);
xor U7684 (N_7684,N_6765,N_6916);
and U7685 (N_7685,N_6940,N_6760);
or U7686 (N_7686,N_7050,N_6834);
xnor U7687 (N_7687,N_7178,N_6641);
nand U7688 (N_7688,N_6887,N_6617);
xor U7689 (N_7689,N_6993,N_7069);
xor U7690 (N_7690,N_7125,N_7027);
xor U7691 (N_7691,N_6922,N_7099);
xor U7692 (N_7692,N_6742,N_7086);
nand U7693 (N_7693,N_6737,N_6924);
nand U7694 (N_7694,N_7168,N_7162);
or U7695 (N_7695,N_6705,N_6991);
or U7696 (N_7696,N_6948,N_7191);
nand U7697 (N_7697,N_7166,N_6604);
and U7698 (N_7698,N_7044,N_6876);
or U7699 (N_7699,N_6798,N_6745);
or U7700 (N_7700,N_7050,N_6821);
nand U7701 (N_7701,N_6733,N_6642);
and U7702 (N_7702,N_7020,N_6723);
or U7703 (N_7703,N_7177,N_6623);
nand U7704 (N_7704,N_7075,N_7026);
nor U7705 (N_7705,N_6743,N_6788);
or U7706 (N_7706,N_6904,N_6861);
and U7707 (N_7707,N_7106,N_6968);
xnor U7708 (N_7708,N_6860,N_6922);
nor U7709 (N_7709,N_6649,N_6784);
or U7710 (N_7710,N_6717,N_6807);
and U7711 (N_7711,N_7118,N_7078);
or U7712 (N_7712,N_7106,N_7006);
nand U7713 (N_7713,N_7198,N_7049);
nand U7714 (N_7714,N_6966,N_7079);
nor U7715 (N_7715,N_6844,N_6996);
xor U7716 (N_7716,N_7012,N_6701);
xnor U7717 (N_7717,N_6954,N_6858);
nand U7718 (N_7718,N_6909,N_7194);
xor U7719 (N_7719,N_7059,N_7157);
xnor U7720 (N_7720,N_6915,N_6620);
or U7721 (N_7721,N_6980,N_6851);
nor U7722 (N_7722,N_6737,N_6986);
nand U7723 (N_7723,N_7007,N_6636);
nand U7724 (N_7724,N_7103,N_6780);
or U7725 (N_7725,N_6880,N_7074);
xor U7726 (N_7726,N_6894,N_7185);
xnor U7727 (N_7727,N_7163,N_6924);
nand U7728 (N_7728,N_7120,N_6951);
or U7729 (N_7729,N_7037,N_6627);
and U7730 (N_7730,N_6919,N_6951);
or U7731 (N_7731,N_6708,N_6744);
nor U7732 (N_7732,N_6849,N_7098);
or U7733 (N_7733,N_6901,N_6787);
or U7734 (N_7734,N_6719,N_6850);
nand U7735 (N_7735,N_7040,N_6928);
nor U7736 (N_7736,N_6942,N_6914);
or U7737 (N_7737,N_7101,N_7173);
xnor U7738 (N_7738,N_6977,N_6711);
or U7739 (N_7739,N_7106,N_6753);
xor U7740 (N_7740,N_6659,N_6809);
nand U7741 (N_7741,N_6758,N_7194);
and U7742 (N_7742,N_7007,N_7021);
nand U7743 (N_7743,N_6956,N_6698);
nand U7744 (N_7744,N_6748,N_6807);
or U7745 (N_7745,N_7063,N_6634);
nand U7746 (N_7746,N_6617,N_7123);
and U7747 (N_7747,N_6821,N_6958);
nand U7748 (N_7748,N_7183,N_6622);
nand U7749 (N_7749,N_6652,N_7047);
xnor U7750 (N_7750,N_6714,N_6755);
xor U7751 (N_7751,N_7102,N_6800);
nand U7752 (N_7752,N_6846,N_7138);
xnor U7753 (N_7753,N_6914,N_6775);
nor U7754 (N_7754,N_6815,N_6685);
xnor U7755 (N_7755,N_6786,N_7148);
nor U7756 (N_7756,N_6843,N_7021);
xnor U7757 (N_7757,N_7108,N_7101);
or U7758 (N_7758,N_6981,N_6676);
xor U7759 (N_7759,N_7126,N_6801);
nand U7760 (N_7760,N_6903,N_6736);
nand U7761 (N_7761,N_6676,N_7033);
nand U7762 (N_7762,N_6638,N_7100);
nand U7763 (N_7763,N_6630,N_7051);
nand U7764 (N_7764,N_6692,N_6696);
or U7765 (N_7765,N_6714,N_6908);
and U7766 (N_7766,N_7067,N_7065);
and U7767 (N_7767,N_6717,N_7181);
and U7768 (N_7768,N_6844,N_6622);
nand U7769 (N_7769,N_7098,N_7076);
and U7770 (N_7770,N_7126,N_7053);
or U7771 (N_7771,N_7038,N_6803);
nor U7772 (N_7772,N_7044,N_6917);
nand U7773 (N_7773,N_6927,N_6735);
xor U7774 (N_7774,N_7148,N_7113);
or U7775 (N_7775,N_7130,N_6931);
nand U7776 (N_7776,N_7174,N_6610);
or U7777 (N_7777,N_6890,N_6725);
nor U7778 (N_7778,N_7139,N_7175);
and U7779 (N_7779,N_7189,N_6905);
or U7780 (N_7780,N_7150,N_6854);
or U7781 (N_7781,N_7193,N_6957);
nand U7782 (N_7782,N_7168,N_6626);
or U7783 (N_7783,N_6663,N_6605);
nor U7784 (N_7784,N_6992,N_7197);
nand U7785 (N_7785,N_6922,N_7107);
nand U7786 (N_7786,N_7070,N_6910);
or U7787 (N_7787,N_7144,N_6699);
xnor U7788 (N_7788,N_6701,N_7173);
or U7789 (N_7789,N_7176,N_6999);
nor U7790 (N_7790,N_7087,N_6828);
xor U7791 (N_7791,N_6750,N_7111);
nor U7792 (N_7792,N_7158,N_6632);
nor U7793 (N_7793,N_7070,N_6688);
nor U7794 (N_7794,N_6927,N_6837);
and U7795 (N_7795,N_6615,N_6894);
and U7796 (N_7796,N_6994,N_7133);
or U7797 (N_7797,N_7146,N_6636);
and U7798 (N_7798,N_6715,N_6894);
nand U7799 (N_7799,N_6917,N_6652);
and U7800 (N_7800,N_7786,N_7266);
xnor U7801 (N_7801,N_7619,N_7315);
nand U7802 (N_7802,N_7685,N_7797);
and U7803 (N_7803,N_7639,N_7226);
nor U7804 (N_7804,N_7218,N_7389);
nand U7805 (N_7805,N_7366,N_7348);
nand U7806 (N_7806,N_7485,N_7722);
and U7807 (N_7807,N_7547,N_7728);
and U7808 (N_7808,N_7751,N_7654);
nor U7809 (N_7809,N_7692,N_7531);
and U7810 (N_7810,N_7541,N_7573);
nand U7811 (N_7811,N_7408,N_7232);
nor U7812 (N_7812,N_7688,N_7788);
nor U7813 (N_7813,N_7529,N_7571);
xnor U7814 (N_7814,N_7718,N_7337);
nand U7815 (N_7815,N_7755,N_7445);
nor U7816 (N_7816,N_7488,N_7320);
or U7817 (N_7817,N_7523,N_7332);
nor U7818 (N_7818,N_7505,N_7411);
nor U7819 (N_7819,N_7511,N_7578);
nand U7820 (N_7820,N_7597,N_7607);
and U7821 (N_7821,N_7720,N_7508);
nor U7822 (N_7822,N_7768,N_7438);
nand U7823 (N_7823,N_7741,N_7596);
xnor U7824 (N_7824,N_7633,N_7361);
xor U7825 (N_7825,N_7455,N_7624);
and U7826 (N_7826,N_7663,N_7785);
nand U7827 (N_7827,N_7612,N_7657);
nor U7828 (N_7828,N_7668,N_7672);
nand U7829 (N_7829,N_7598,N_7662);
or U7830 (N_7830,N_7482,N_7664);
xnor U7831 (N_7831,N_7223,N_7393);
or U7832 (N_7832,N_7609,N_7414);
xnor U7833 (N_7833,N_7453,N_7757);
or U7834 (N_7834,N_7795,N_7739);
or U7835 (N_7835,N_7431,N_7250);
or U7836 (N_7836,N_7477,N_7373);
nand U7837 (N_7837,N_7342,N_7263);
and U7838 (N_7838,N_7655,N_7420);
or U7839 (N_7839,N_7271,N_7409);
nor U7840 (N_7840,N_7355,N_7748);
nor U7841 (N_7841,N_7790,N_7333);
and U7842 (N_7842,N_7632,N_7673);
nor U7843 (N_7843,N_7585,N_7303);
xnor U7844 (N_7844,N_7225,N_7273);
xnor U7845 (N_7845,N_7686,N_7599);
nor U7846 (N_7846,N_7392,N_7636);
nand U7847 (N_7847,N_7564,N_7527);
nor U7848 (N_7848,N_7298,N_7563);
and U7849 (N_7849,N_7721,N_7209);
nand U7850 (N_7850,N_7487,N_7614);
and U7851 (N_7851,N_7550,N_7693);
and U7852 (N_7852,N_7454,N_7635);
and U7853 (N_7853,N_7725,N_7424);
xnor U7854 (N_7854,N_7500,N_7778);
nor U7855 (N_7855,N_7690,N_7615);
or U7856 (N_7856,N_7317,N_7717);
nand U7857 (N_7857,N_7306,N_7435);
xor U7858 (N_7858,N_7709,N_7534);
and U7859 (N_7859,N_7467,N_7308);
or U7860 (N_7860,N_7386,N_7416);
or U7861 (N_7861,N_7759,N_7283);
and U7862 (N_7862,N_7257,N_7479);
xnor U7863 (N_7863,N_7764,N_7203);
xor U7864 (N_7864,N_7377,N_7566);
xor U7865 (N_7865,N_7284,N_7666);
nand U7866 (N_7866,N_7753,N_7542);
nand U7867 (N_7867,N_7740,N_7448);
nand U7868 (N_7868,N_7781,N_7407);
or U7869 (N_7869,N_7429,N_7208);
nor U7870 (N_7870,N_7572,N_7265);
or U7871 (N_7871,N_7696,N_7490);
nor U7872 (N_7872,N_7282,N_7552);
and U7873 (N_7873,N_7754,N_7618);
xnor U7874 (N_7874,N_7553,N_7695);
xor U7875 (N_7875,N_7352,N_7227);
or U7876 (N_7876,N_7346,N_7702);
nand U7877 (N_7877,N_7697,N_7770);
xor U7878 (N_7878,N_7796,N_7684);
or U7879 (N_7879,N_7360,N_7787);
or U7880 (N_7880,N_7592,N_7267);
xor U7881 (N_7881,N_7470,N_7396);
xnor U7882 (N_7882,N_7460,N_7325);
or U7883 (N_7883,N_7545,N_7322);
and U7884 (N_7884,N_7533,N_7275);
nand U7885 (N_7885,N_7581,N_7792);
nand U7886 (N_7886,N_7365,N_7749);
nand U7887 (N_7887,N_7210,N_7574);
nand U7888 (N_7888,N_7558,N_7628);
and U7889 (N_7889,N_7756,N_7241);
or U7890 (N_7890,N_7319,N_7510);
or U7891 (N_7891,N_7653,N_7595);
nor U7892 (N_7892,N_7665,N_7425);
or U7893 (N_7893,N_7437,N_7736);
xor U7894 (N_7894,N_7670,N_7214);
nor U7895 (N_7895,N_7499,N_7334);
nor U7896 (N_7896,N_7743,N_7606);
and U7897 (N_7897,N_7674,N_7551);
nand U7898 (N_7898,N_7486,N_7459);
nand U7899 (N_7899,N_7538,N_7703);
xor U7900 (N_7900,N_7339,N_7400);
nor U7901 (N_7901,N_7652,N_7602);
nand U7902 (N_7902,N_7212,N_7388);
and U7903 (N_7903,N_7643,N_7710);
nand U7904 (N_7904,N_7216,N_7731);
xor U7905 (N_7905,N_7671,N_7474);
nor U7906 (N_7906,N_7447,N_7752);
and U7907 (N_7907,N_7421,N_7561);
xor U7908 (N_7908,N_7577,N_7313);
nor U7909 (N_7909,N_7760,N_7517);
xor U7910 (N_7910,N_7481,N_7548);
nand U7911 (N_7911,N_7773,N_7291);
nor U7912 (N_7912,N_7648,N_7469);
nand U7913 (N_7913,N_7343,N_7237);
nand U7914 (N_7914,N_7353,N_7213);
xnor U7915 (N_7915,N_7289,N_7516);
nand U7916 (N_7916,N_7262,N_7428);
nor U7917 (N_7917,N_7627,N_7323);
xnor U7918 (N_7918,N_7415,N_7476);
and U7919 (N_7919,N_7626,N_7277);
xnor U7920 (N_7920,N_7766,N_7590);
or U7921 (N_7921,N_7395,N_7309);
nor U7922 (N_7922,N_7496,N_7582);
nand U7923 (N_7923,N_7798,N_7642);
nand U7924 (N_7924,N_7629,N_7625);
nand U7925 (N_7925,N_7616,N_7507);
nor U7926 (N_7926,N_7682,N_7364);
xnor U7927 (N_7927,N_7274,N_7234);
or U7928 (N_7928,N_7557,N_7704);
and U7929 (N_7929,N_7245,N_7789);
and U7930 (N_7930,N_7535,N_7280);
nand U7931 (N_7931,N_7699,N_7726);
xor U7932 (N_7932,N_7600,N_7379);
nor U7933 (N_7933,N_7347,N_7371);
and U7934 (N_7934,N_7771,N_7502);
nand U7935 (N_7935,N_7401,N_7363);
nand U7936 (N_7936,N_7276,N_7270);
and U7937 (N_7937,N_7418,N_7784);
nand U7938 (N_7938,N_7587,N_7576);
xnor U7939 (N_7939,N_7368,N_7242);
and U7940 (N_7940,N_7465,N_7583);
nor U7941 (N_7941,N_7777,N_7405);
and U7942 (N_7942,N_7555,N_7520);
xnor U7943 (N_7943,N_7473,N_7656);
and U7944 (N_7944,N_7433,N_7249);
nand U7945 (N_7945,N_7412,N_7525);
nand U7946 (N_7946,N_7559,N_7205);
xnor U7947 (N_7947,N_7794,N_7514);
or U7948 (N_7948,N_7630,N_7314);
nand U7949 (N_7949,N_7734,N_7281);
and U7950 (N_7950,N_7236,N_7349);
or U7951 (N_7951,N_7480,N_7229);
and U7952 (N_7952,N_7640,N_7336);
nor U7953 (N_7953,N_7747,N_7436);
nor U7954 (N_7954,N_7732,N_7567);
xnor U7955 (N_7955,N_7712,N_7378);
nand U7956 (N_7956,N_7610,N_7296);
and U7957 (N_7957,N_7530,N_7316);
xor U7958 (N_7958,N_7675,N_7307);
xnor U7959 (N_7959,N_7367,N_7617);
nor U7960 (N_7960,N_7374,N_7345);
nor U7961 (N_7961,N_7518,N_7432);
and U7962 (N_7962,N_7466,N_7501);
xnor U7963 (N_7963,N_7341,N_7427);
xnor U7964 (N_7964,N_7680,N_7338);
and U7965 (N_7965,N_7586,N_7492);
xor U7966 (N_7966,N_7536,N_7260);
or U7967 (N_7967,N_7761,N_7750);
and U7968 (N_7968,N_7515,N_7406);
nand U7969 (N_7969,N_7248,N_7272);
nor U7970 (N_7970,N_7522,N_7247);
or U7971 (N_7971,N_7758,N_7713);
and U7972 (N_7972,N_7397,N_7532);
xnor U7973 (N_7973,N_7637,N_7575);
or U7974 (N_7974,N_7509,N_7782);
or U7975 (N_7975,N_7239,N_7278);
or U7976 (N_7976,N_7677,N_7321);
and U7977 (N_7977,N_7204,N_7442);
xnor U7978 (N_7978,N_7285,N_7200);
or U7979 (N_7979,N_7495,N_7791);
nand U7980 (N_7980,N_7410,N_7201);
nor U7981 (N_7981,N_7434,N_7261);
xnor U7982 (N_7982,N_7661,N_7290);
or U7983 (N_7983,N_7799,N_7694);
and U7984 (N_7984,N_7570,N_7252);
or U7985 (N_7985,N_7310,N_7591);
nor U7986 (N_7986,N_7745,N_7330);
or U7987 (N_7987,N_7294,N_7601);
and U7988 (N_7988,N_7464,N_7344);
or U7989 (N_7989,N_7255,N_7312);
nor U7990 (N_7990,N_7651,N_7351);
nor U7991 (N_7991,N_7390,N_7472);
and U7992 (N_7992,N_7611,N_7372);
and U7993 (N_7993,N_7579,N_7484);
and U7994 (N_7994,N_7475,N_7235);
or U7995 (N_7995,N_7659,N_7658);
or U7996 (N_7996,N_7258,N_7644);
nand U7997 (N_7997,N_7569,N_7256);
nand U7998 (N_7998,N_7705,N_7449);
nand U7999 (N_7999,N_7506,N_7776);
xor U8000 (N_8000,N_7299,N_7620);
or U8001 (N_8001,N_7384,N_7783);
and U8002 (N_8002,N_7793,N_7546);
xor U8003 (N_8003,N_7621,N_7254);
xnor U8004 (N_8004,N_7382,N_7593);
or U8005 (N_8005,N_7549,N_7327);
nand U8006 (N_8006,N_7498,N_7707);
and U8007 (N_8007,N_7780,N_7269);
nor U8008 (N_8008,N_7737,N_7305);
xnor U8009 (N_8009,N_7471,N_7251);
or U8010 (N_8010,N_7422,N_7253);
or U8011 (N_8011,N_7383,N_7376);
xor U8012 (N_8012,N_7413,N_7613);
nand U8013 (N_8013,N_7729,N_7526);
or U8014 (N_8014,N_7451,N_7311);
or U8015 (N_8015,N_7207,N_7300);
nand U8016 (N_8016,N_7774,N_7715);
and U8017 (N_8017,N_7391,N_7733);
nor U8018 (N_8018,N_7556,N_7206);
or U8019 (N_8019,N_7678,N_7419);
xor U8020 (N_8020,N_7667,N_7562);
nor U8021 (N_8021,N_7369,N_7439);
nor U8022 (N_8022,N_7727,N_7603);
nand U8023 (N_8023,N_7238,N_7608);
nor U8024 (N_8024,N_7669,N_7244);
nor U8025 (N_8025,N_7356,N_7497);
nor U8026 (N_8026,N_7647,N_7701);
nor U8027 (N_8027,N_7634,N_7403);
nand U8028 (N_8028,N_7228,N_7426);
and U8029 (N_8029,N_7302,N_7240);
nand U8030 (N_8030,N_7660,N_7354);
nor U8031 (N_8031,N_7394,N_7358);
xor U8032 (N_8032,N_7708,N_7691);
nor U8033 (N_8033,N_7493,N_7404);
xnor U8034 (N_8034,N_7463,N_7537);
nand U8035 (N_8035,N_7211,N_7233);
and U8036 (N_8036,N_7243,N_7452);
or U8037 (N_8037,N_7259,N_7221);
or U8038 (N_8038,N_7350,N_7217);
and U8039 (N_8039,N_7646,N_7494);
xnor U8040 (N_8040,N_7735,N_7623);
nand U8041 (N_8041,N_7645,N_7524);
xor U8042 (N_8042,N_7588,N_7594);
and U8043 (N_8043,N_7723,N_7744);
nor U8044 (N_8044,N_7304,N_7335);
nand U8045 (N_8045,N_7554,N_7268);
xnor U8046 (N_8046,N_7700,N_7443);
or U8047 (N_8047,N_7698,N_7219);
nor U8048 (N_8048,N_7292,N_7444);
and U8049 (N_8049,N_7220,N_7402);
nand U8050 (N_8050,N_7456,N_7746);
and U8051 (N_8051,N_7279,N_7458);
xnor U8052 (N_8052,N_7417,N_7687);
nand U8053 (N_8053,N_7503,N_7326);
or U8054 (N_8054,N_7539,N_7544);
nor U8055 (N_8055,N_7775,N_7769);
and U8056 (N_8056,N_7457,N_7478);
and U8057 (N_8057,N_7224,N_7540);
xor U8058 (N_8058,N_7560,N_7286);
and U8059 (N_8059,N_7340,N_7398);
nand U8060 (N_8060,N_7331,N_7711);
nor U8061 (N_8061,N_7297,N_7767);
nor U8062 (N_8062,N_7638,N_7706);
xor U8063 (N_8063,N_7568,N_7264);
nand U8064 (N_8064,N_7580,N_7719);
xnor U8065 (N_8065,N_7762,N_7779);
or U8066 (N_8066,N_7649,N_7521);
and U8067 (N_8067,N_7604,N_7375);
nand U8068 (N_8068,N_7589,N_7222);
nand U8069 (N_8069,N_7716,N_7446);
and U8070 (N_8070,N_7288,N_7230);
or U8071 (N_8071,N_7430,N_7519);
nor U8072 (N_8072,N_7742,N_7468);
and U8073 (N_8073,N_7440,N_7381);
nand U8074 (N_8074,N_7483,N_7287);
and U8075 (N_8075,N_7681,N_7513);
nor U8076 (N_8076,N_7324,N_7528);
nor U8077 (N_8077,N_7683,N_7679);
and U8078 (N_8078,N_7462,N_7301);
xnor U8079 (N_8079,N_7202,N_7724);
nand U8080 (N_8080,N_7441,N_7461);
nor U8081 (N_8081,N_7423,N_7357);
nand U8082 (N_8082,N_7380,N_7370);
or U8083 (N_8083,N_7450,N_7385);
nor U8084 (N_8084,N_7738,N_7512);
nand U8085 (N_8085,N_7714,N_7676);
and U8086 (N_8086,N_7359,N_7399);
nand U8087 (N_8087,N_7293,N_7772);
and U8088 (N_8088,N_7491,N_7763);
xor U8089 (N_8089,N_7504,N_7622);
nand U8090 (N_8090,N_7246,N_7689);
and U8091 (N_8091,N_7631,N_7295);
and U8092 (N_8092,N_7650,N_7489);
xnor U8093 (N_8093,N_7328,N_7730);
or U8094 (N_8094,N_7641,N_7231);
and U8095 (N_8095,N_7543,N_7387);
nand U8096 (N_8096,N_7215,N_7318);
and U8097 (N_8097,N_7362,N_7329);
and U8098 (N_8098,N_7565,N_7765);
nand U8099 (N_8099,N_7584,N_7605);
xnor U8100 (N_8100,N_7444,N_7630);
nand U8101 (N_8101,N_7445,N_7578);
nor U8102 (N_8102,N_7792,N_7794);
nor U8103 (N_8103,N_7661,N_7299);
and U8104 (N_8104,N_7343,N_7746);
xnor U8105 (N_8105,N_7282,N_7255);
and U8106 (N_8106,N_7492,N_7781);
nand U8107 (N_8107,N_7799,N_7268);
xnor U8108 (N_8108,N_7696,N_7726);
or U8109 (N_8109,N_7286,N_7509);
xor U8110 (N_8110,N_7589,N_7392);
or U8111 (N_8111,N_7451,N_7726);
nor U8112 (N_8112,N_7243,N_7713);
and U8113 (N_8113,N_7668,N_7396);
or U8114 (N_8114,N_7320,N_7393);
or U8115 (N_8115,N_7644,N_7702);
nand U8116 (N_8116,N_7326,N_7782);
nand U8117 (N_8117,N_7569,N_7755);
or U8118 (N_8118,N_7262,N_7684);
and U8119 (N_8119,N_7730,N_7204);
nand U8120 (N_8120,N_7337,N_7284);
and U8121 (N_8121,N_7774,N_7506);
and U8122 (N_8122,N_7521,N_7714);
xor U8123 (N_8123,N_7233,N_7569);
or U8124 (N_8124,N_7290,N_7319);
xnor U8125 (N_8125,N_7512,N_7550);
or U8126 (N_8126,N_7264,N_7660);
nor U8127 (N_8127,N_7335,N_7618);
and U8128 (N_8128,N_7231,N_7431);
nor U8129 (N_8129,N_7666,N_7489);
or U8130 (N_8130,N_7752,N_7522);
nor U8131 (N_8131,N_7282,N_7259);
nand U8132 (N_8132,N_7701,N_7686);
nand U8133 (N_8133,N_7743,N_7337);
or U8134 (N_8134,N_7273,N_7415);
or U8135 (N_8135,N_7519,N_7457);
or U8136 (N_8136,N_7254,N_7670);
or U8137 (N_8137,N_7605,N_7449);
and U8138 (N_8138,N_7713,N_7638);
nor U8139 (N_8139,N_7307,N_7238);
or U8140 (N_8140,N_7792,N_7258);
xor U8141 (N_8141,N_7685,N_7225);
nand U8142 (N_8142,N_7553,N_7599);
xor U8143 (N_8143,N_7546,N_7739);
and U8144 (N_8144,N_7467,N_7477);
nand U8145 (N_8145,N_7346,N_7784);
and U8146 (N_8146,N_7519,N_7576);
nor U8147 (N_8147,N_7490,N_7287);
nand U8148 (N_8148,N_7455,N_7552);
nor U8149 (N_8149,N_7555,N_7474);
nand U8150 (N_8150,N_7713,N_7368);
and U8151 (N_8151,N_7353,N_7370);
nand U8152 (N_8152,N_7468,N_7547);
xor U8153 (N_8153,N_7725,N_7668);
nand U8154 (N_8154,N_7687,N_7655);
nand U8155 (N_8155,N_7605,N_7395);
nand U8156 (N_8156,N_7569,N_7292);
xor U8157 (N_8157,N_7202,N_7786);
xor U8158 (N_8158,N_7447,N_7685);
nand U8159 (N_8159,N_7732,N_7479);
nand U8160 (N_8160,N_7709,N_7402);
xor U8161 (N_8161,N_7442,N_7295);
or U8162 (N_8162,N_7256,N_7610);
nand U8163 (N_8163,N_7479,N_7597);
or U8164 (N_8164,N_7451,N_7730);
nand U8165 (N_8165,N_7390,N_7209);
xor U8166 (N_8166,N_7430,N_7385);
and U8167 (N_8167,N_7332,N_7327);
or U8168 (N_8168,N_7461,N_7559);
nand U8169 (N_8169,N_7350,N_7731);
or U8170 (N_8170,N_7239,N_7531);
xor U8171 (N_8171,N_7698,N_7239);
nor U8172 (N_8172,N_7550,N_7325);
nor U8173 (N_8173,N_7523,N_7376);
nand U8174 (N_8174,N_7707,N_7592);
nor U8175 (N_8175,N_7290,N_7468);
xnor U8176 (N_8176,N_7300,N_7619);
and U8177 (N_8177,N_7441,N_7466);
xnor U8178 (N_8178,N_7283,N_7637);
nor U8179 (N_8179,N_7627,N_7538);
nor U8180 (N_8180,N_7695,N_7735);
nor U8181 (N_8181,N_7795,N_7286);
nor U8182 (N_8182,N_7683,N_7601);
xor U8183 (N_8183,N_7597,N_7583);
nand U8184 (N_8184,N_7685,N_7342);
nor U8185 (N_8185,N_7732,N_7717);
nand U8186 (N_8186,N_7230,N_7784);
xor U8187 (N_8187,N_7277,N_7433);
nor U8188 (N_8188,N_7657,N_7429);
xor U8189 (N_8189,N_7393,N_7457);
or U8190 (N_8190,N_7265,N_7588);
nand U8191 (N_8191,N_7236,N_7699);
xnor U8192 (N_8192,N_7623,N_7772);
or U8193 (N_8193,N_7491,N_7617);
and U8194 (N_8194,N_7355,N_7545);
or U8195 (N_8195,N_7338,N_7667);
or U8196 (N_8196,N_7770,N_7457);
or U8197 (N_8197,N_7698,N_7517);
xnor U8198 (N_8198,N_7728,N_7208);
and U8199 (N_8199,N_7692,N_7272);
nand U8200 (N_8200,N_7720,N_7717);
xor U8201 (N_8201,N_7290,N_7768);
and U8202 (N_8202,N_7530,N_7760);
xor U8203 (N_8203,N_7376,N_7425);
nand U8204 (N_8204,N_7294,N_7464);
nor U8205 (N_8205,N_7497,N_7636);
nand U8206 (N_8206,N_7425,N_7213);
nor U8207 (N_8207,N_7311,N_7490);
or U8208 (N_8208,N_7398,N_7685);
nor U8209 (N_8209,N_7663,N_7732);
or U8210 (N_8210,N_7710,N_7479);
and U8211 (N_8211,N_7299,N_7354);
nand U8212 (N_8212,N_7272,N_7579);
and U8213 (N_8213,N_7441,N_7742);
or U8214 (N_8214,N_7677,N_7505);
nor U8215 (N_8215,N_7489,N_7392);
or U8216 (N_8216,N_7537,N_7765);
and U8217 (N_8217,N_7799,N_7292);
xnor U8218 (N_8218,N_7533,N_7448);
nor U8219 (N_8219,N_7611,N_7417);
or U8220 (N_8220,N_7304,N_7798);
nand U8221 (N_8221,N_7289,N_7298);
xnor U8222 (N_8222,N_7664,N_7396);
nor U8223 (N_8223,N_7307,N_7544);
nand U8224 (N_8224,N_7774,N_7653);
or U8225 (N_8225,N_7476,N_7593);
or U8226 (N_8226,N_7730,N_7301);
nor U8227 (N_8227,N_7300,N_7426);
nor U8228 (N_8228,N_7309,N_7656);
xnor U8229 (N_8229,N_7484,N_7687);
nor U8230 (N_8230,N_7482,N_7636);
nor U8231 (N_8231,N_7512,N_7786);
nand U8232 (N_8232,N_7367,N_7548);
xnor U8233 (N_8233,N_7458,N_7726);
xor U8234 (N_8234,N_7393,N_7701);
or U8235 (N_8235,N_7761,N_7379);
xnor U8236 (N_8236,N_7205,N_7767);
nand U8237 (N_8237,N_7659,N_7350);
nand U8238 (N_8238,N_7692,N_7611);
xnor U8239 (N_8239,N_7494,N_7303);
nand U8240 (N_8240,N_7642,N_7275);
and U8241 (N_8241,N_7509,N_7263);
xor U8242 (N_8242,N_7393,N_7492);
or U8243 (N_8243,N_7334,N_7263);
xnor U8244 (N_8244,N_7691,N_7244);
nor U8245 (N_8245,N_7736,N_7610);
nor U8246 (N_8246,N_7618,N_7504);
nor U8247 (N_8247,N_7232,N_7420);
nand U8248 (N_8248,N_7549,N_7624);
and U8249 (N_8249,N_7617,N_7335);
nor U8250 (N_8250,N_7507,N_7677);
nand U8251 (N_8251,N_7474,N_7424);
and U8252 (N_8252,N_7256,N_7659);
nor U8253 (N_8253,N_7480,N_7734);
xnor U8254 (N_8254,N_7389,N_7449);
or U8255 (N_8255,N_7726,N_7590);
xnor U8256 (N_8256,N_7378,N_7681);
nand U8257 (N_8257,N_7543,N_7623);
and U8258 (N_8258,N_7748,N_7741);
or U8259 (N_8259,N_7584,N_7782);
nand U8260 (N_8260,N_7424,N_7247);
and U8261 (N_8261,N_7513,N_7342);
nor U8262 (N_8262,N_7398,N_7566);
or U8263 (N_8263,N_7743,N_7233);
nor U8264 (N_8264,N_7762,N_7636);
or U8265 (N_8265,N_7473,N_7438);
nor U8266 (N_8266,N_7644,N_7506);
xor U8267 (N_8267,N_7483,N_7795);
xor U8268 (N_8268,N_7642,N_7512);
nor U8269 (N_8269,N_7446,N_7674);
nand U8270 (N_8270,N_7354,N_7251);
nand U8271 (N_8271,N_7312,N_7348);
or U8272 (N_8272,N_7287,N_7424);
or U8273 (N_8273,N_7386,N_7341);
xor U8274 (N_8274,N_7303,N_7423);
nor U8275 (N_8275,N_7755,N_7303);
xnor U8276 (N_8276,N_7508,N_7348);
xnor U8277 (N_8277,N_7559,N_7789);
xnor U8278 (N_8278,N_7469,N_7454);
xor U8279 (N_8279,N_7420,N_7477);
xnor U8280 (N_8280,N_7547,N_7524);
nor U8281 (N_8281,N_7200,N_7617);
or U8282 (N_8282,N_7402,N_7602);
and U8283 (N_8283,N_7500,N_7678);
or U8284 (N_8284,N_7500,N_7630);
nor U8285 (N_8285,N_7554,N_7422);
xnor U8286 (N_8286,N_7695,N_7207);
and U8287 (N_8287,N_7740,N_7328);
or U8288 (N_8288,N_7709,N_7620);
or U8289 (N_8289,N_7514,N_7636);
nand U8290 (N_8290,N_7619,N_7736);
nor U8291 (N_8291,N_7425,N_7419);
or U8292 (N_8292,N_7585,N_7460);
and U8293 (N_8293,N_7295,N_7768);
xnor U8294 (N_8294,N_7335,N_7279);
or U8295 (N_8295,N_7384,N_7795);
nor U8296 (N_8296,N_7396,N_7748);
or U8297 (N_8297,N_7273,N_7481);
xnor U8298 (N_8298,N_7353,N_7560);
nor U8299 (N_8299,N_7515,N_7402);
and U8300 (N_8300,N_7630,N_7665);
and U8301 (N_8301,N_7316,N_7370);
nand U8302 (N_8302,N_7539,N_7557);
xnor U8303 (N_8303,N_7693,N_7706);
or U8304 (N_8304,N_7608,N_7369);
or U8305 (N_8305,N_7497,N_7319);
and U8306 (N_8306,N_7520,N_7386);
or U8307 (N_8307,N_7302,N_7791);
nand U8308 (N_8308,N_7427,N_7668);
nand U8309 (N_8309,N_7228,N_7677);
xnor U8310 (N_8310,N_7529,N_7539);
and U8311 (N_8311,N_7212,N_7694);
xnor U8312 (N_8312,N_7636,N_7294);
nor U8313 (N_8313,N_7658,N_7378);
nand U8314 (N_8314,N_7731,N_7453);
nor U8315 (N_8315,N_7636,N_7435);
nand U8316 (N_8316,N_7430,N_7603);
xnor U8317 (N_8317,N_7484,N_7533);
nor U8318 (N_8318,N_7221,N_7673);
nor U8319 (N_8319,N_7695,N_7598);
xnor U8320 (N_8320,N_7330,N_7401);
nand U8321 (N_8321,N_7319,N_7546);
nor U8322 (N_8322,N_7714,N_7760);
and U8323 (N_8323,N_7695,N_7541);
and U8324 (N_8324,N_7266,N_7540);
and U8325 (N_8325,N_7431,N_7255);
and U8326 (N_8326,N_7389,N_7785);
xor U8327 (N_8327,N_7478,N_7542);
or U8328 (N_8328,N_7385,N_7271);
nor U8329 (N_8329,N_7640,N_7276);
or U8330 (N_8330,N_7468,N_7253);
xor U8331 (N_8331,N_7470,N_7286);
xor U8332 (N_8332,N_7743,N_7568);
nand U8333 (N_8333,N_7745,N_7346);
nand U8334 (N_8334,N_7432,N_7392);
and U8335 (N_8335,N_7594,N_7751);
xnor U8336 (N_8336,N_7591,N_7571);
xor U8337 (N_8337,N_7415,N_7233);
nand U8338 (N_8338,N_7597,N_7548);
and U8339 (N_8339,N_7357,N_7538);
nor U8340 (N_8340,N_7522,N_7328);
and U8341 (N_8341,N_7612,N_7420);
or U8342 (N_8342,N_7207,N_7626);
or U8343 (N_8343,N_7711,N_7315);
or U8344 (N_8344,N_7327,N_7708);
nor U8345 (N_8345,N_7515,N_7506);
nor U8346 (N_8346,N_7757,N_7695);
and U8347 (N_8347,N_7748,N_7416);
nand U8348 (N_8348,N_7782,N_7348);
or U8349 (N_8349,N_7262,N_7352);
or U8350 (N_8350,N_7623,N_7224);
nor U8351 (N_8351,N_7632,N_7571);
nand U8352 (N_8352,N_7397,N_7279);
nor U8353 (N_8353,N_7221,N_7322);
and U8354 (N_8354,N_7627,N_7392);
or U8355 (N_8355,N_7562,N_7260);
nor U8356 (N_8356,N_7323,N_7349);
xor U8357 (N_8357,N_7357,N_7385);
and U8358 (N_8358,N_7541,N_7374);
and U8359 (N_8359,N_7468,N_7549);
nand U8360 (N_8360,N_7754,N_7224);
nor U8361 (N_8361,N_7505,N_7664);
or U8362 (N_8362,N_7625,N_7219);
and U8363 (N_8363,N_7727,N_7764);
xnor U8364 (N_8364,N_7459,N_7569);
and U8365 (N_8365,N_7564,N_7250);
nand U8366 (N_8366,N_7362,N_7571);
nor U8367 (N_8367,N_7351,N_7611);
and U8368 (N_8368,N_7523,N_7300);
and U8369 (N_8369,N_7662,N_7565);
or U8370 (N_8370,N_7229,N_7386);
nor U8371 (N_8371,N_7601,N_7726);
xor U8372 (N_8372,N_7675,N_7498);
or U8373 (N_8373,N_7213,N_7479);
or U8374 (N_8374,N_7560,N_7536);
nand U8375 (N_8375,N_7406,N_7391);
and U8376 (N_8376,N_7733,N_7354);
nor U8377 (N_8377,N_7773,N_7535);
xor U8378 (N_8378,N_7212,N_7403);
or U8379 (N_8379,N_7493,N_7594);
nand U8380 (N_8380,N_7489,N_7262);
nand U8381 (N_8381,N_7612,N_7705);
or U8382 (N_8382,N_7709,N_7329);
xnor U8383 (N_8383,N_7720,N_7514);
and U8384 (N_8384,N_7778,N_7775);
or U8385 (N_8385,N_7390,N_7659);
or U8386 (N_8386,N_7445,N_7698);
xor U8387 (N_8387,N_7463,N_7727);
and U8388 (N_8388,N_7210,N_7206);
nand U8389 (N_8389,N_7621,N_7220);
nor U8390 (N_8390,N_7684,N_7717);
and U8391 (N_8391,N_7285,N_7775);
nand U8392 (N_8392,N_7489,N_7492);
or U8393 (N_8393,N_7795,N_7606);
and U8394 (N_8394,N_7321,N_7615);
nand U8395 (N_8395,N_7668,N_7209);
nand U8396 (N_8396,N_7204,N_7676);
nor U8397 (N_8397,N_7321,N_7517);
nand U8398 (N_8398,N_7310,N_7459);
nand U8399 (N_8399,N_7291,N_7429);
or U8400 (N_8400,N_8326,N_8273);
nand U8401 (N_8401,N_8118,N_7871);
xnor U8402 (N_8402,N_8318,N_7833);
and U8403 (N_8403,N_8036,N_8054);
nand U8404 (N_8404,N_7874,N_7901);
nor U8405 (N_8405,N_8007,N_8065);
or U8406 (N_8406,N_7851,N_8089);
and U8407 (N_8407,N_8372,N_8158);
nand U8408 (N_8408,N_8191,N_8321);
and U8409 (N_8409,N_8019,N_8307);
and U8410 (N_8410,N_7900,N_8251);
xnor U8411 (N_8411,N_7811,N_8346);
xor U8412 (N_8412,N_8051,N_7890);
nand U8413 (N_8413,N_8300,N_8109);
and U8414 (N_8414,N_7841,N_8210);
nor U8415 (N_8415,N_8357,N_7870);
nor U8416 (N_8416,N_8004,N_7946);
nand U8417 (N_8417,N_8341,N_8181);
nand U8418 (N_8418,N_8121,N_8388);
nand U8419 (N_8419,N_8042,N_8186);
xor U8420 (N_8420,N_8205,N_8258);
xnor U8421 (N_8421,N_7828,N_8085);
nor U8422 (N_8422,N_8136,N_8267);
xnor U8423 (N_8423,N_7985,N_8241);
and U8424 (N_8424,N_7827,N_7896);
or U8425 (N_8425,N_8268,N_8200);
nand U8426 (N_8426,N_7826,N_8132);
and U8427 (N_8427,N_7978,N_8365);
or U8428 (N_8428,N_8142,N_8285);
nor U8429 (N_8429,N_8069,N_8304);
or U8430 (N_8430,N_7962,N_7865);
or U8431 (N_8431,N_7913,N_8030);
nand U8432 (N_8432,N_7824,N_8246);
or U8433 (N_8433,N_8367,N_8391);
or U8434 (N_8434,N_8112,N_8339);
or U8435 (N_8435,N_8049,N_8182);
or U8436 (N_8436,N_8274,N_8392);
and U8437 (N_8437,N_8249,N_7937);
xnor U8438 (N_8438,N_7810,N_7869);
nand U8439 (N_8439,N_8068,N_8298);
or U8440 (N_8440,N_8359,N_7873);
nand U8441 (N_8441,N_8232,N_8043);
nand U8442 (N_8442,N_8102,N_8034);
nor U8443 (N_8443,N_7989,N_8343);
nor U8444 (N_8444,N_8187,N_8399);
nand U8445 (N_8445,N_8235,N_8344);
xor U8446 (N_8446,N_8302,N_7808);
or U8447 (N_8447,N_7941,N_8101);
and U8448 (N_8448,N_7894,N_7880);
xor U8449 (N_8449,N_8259,N_8203);
nand U8450 (N_8450,N_7816,N_8296);
nand U8451 (N_8451,N_7991,N_7943);
and U8452 (N_8452,N_7909,N_8292);
and U8453 (N_8453,N_8199,N_8384);
nand U8454 (N_8454,N_8070,N_8322);
or U8455 (N_8455,N_8312,N_7858);
and U8456 (N_8456,N_8192,N_8381);
nand U8457 (N_8457,N_7812,N_7912);
nand U8458 (N_8458,N_7961,N_8373);
xnor U8459 (N_8459,N_8166,N_8234);
xnor U8460 (N_8460,N_8299,N_7883);
and U8461 (N_8461,N_8082,N_8333);
or U8462 (N_8462,N_8347,N_7936);
xnor U8463 (N_8463,N_8035,N_8281);
or U8464 (N_8464,N_8330,N_8100);
nor U8465 (N_8465,N_8371,N_7945);
or U8466 (N_8466,N_8272,N_7916);
and U8467 (N_8467,N_8092,N_7971);
xnor U8468 (N_8468,N_7881,N_8348);
and U8469 (N_8469,N_7846,N_8024);
nor U8470 (N_8470,N_8047,N_8215);
and U8471 (N_8471,N_8309,N_8176);
xor U8472 (N_8472,N_7845,N_8099);
and U8473 (N_8473,N_8290,N_7859);
xnor U8474 (N_8474,N_8012,N_8243);
and U8475 (N_8475,N_7829,N_8002);
nand U8476 (N_8476,N_8340,N_7932);
xor U8477 (N_8477,N_8147,N_7879);
nand U8478 (N_8478,N_8233,N_7903);
xor U8479 (N_8479,N_7821,N_8150);
or U8480 (N_8480,N_8264,N_8319);
or U8481 (N_8481,N_7839,N_8239);
or U8482 (N_8482,N_8140,N_8098);
or U8483 (N_8483,N_7997,N_8366);
and U8484 (N_8484,N_7818,N_8238);
xor U8485 (N_8485,N_8308,N_8013);
or U8486 (N_8486,N_7999,N_7897);
and U8487 (N_8487,N_8072,N_8214);
or U8488 (N_8488,N_7995,N_8360);
xnor U8489 (N_8489,N_8156,N_7847);
xor U8490 (N_8490,N_8288,N_8354);
nand U8491 (N_8491,N_7944,N_8248);
nand U8492 (N_8492,N_7918,N_8114);
or U8493 (N_8493,N_8057,N_8219);
nand U8494 (N_8494,N_8025,N_8189);
xor U8495 (N_8495,N_8066,N_8113);
xnor U8496 (N_8496,N_8120,N_8311);
and U8497 (N_8497,N_7996,N_8084);
xor U8498 (N_8498,N_8055,N_8332);
or U8499 (N_8499,N_8379,N_8198);
and U8500 (N_8500,N_8064,N_7804);
and U8501 (N_8501,N_8208,N_8095);
nand U8502 (N_8502,N_8301,N_7959);
nor U8503 (N_8503,N_8244,N_7877);
and U8504 (N_8504,N_7927,N_8173);
xor U8505 (N_8505,N_8270,N_8393);
nand U8506 (N_8506,N_7835,N_8096);
or U8507 (N_8507,N_8094,N_7921);
nand U8508 (N_8508,N_8293,N_7954);
nor U8509 (N_8509,N_7875,N_7853);
or U8510 (N_8510,N_7957,N_7963);
nor U8511 (N_8511,N_8141,N_8387);
nor U8512 (N_8512,N_8106,N_8152);
nor U8513 (N_8513,N_7805,N_8190);
or U8514 (N_8514,N_7919,N_7914);
nand U8515 (N_8515,N_8044,N_8011);
nor U8516 (N_8516,N_7942,N_8265);
xnor U8517 (N_8517,N_7972,N_8317);
nor U8518 (N_8518,N_8336,N_8133);
and U8519 (N_8519,N_8017,N_8088);
xnor U8520 (N_8520,N_7861,N_7930);
xor U8521 (N_8521,N_7905,N_8240);
xnor U8522 (N_8522,N_8124,N_8380);
nor U8523 (N_8523,N_8079,N_8236);
nand U8524 (N_8524,N_8223,N_7822);
nand U8525 (N_8525,N_8029,N_7837);
and U8526 (N_8526,N_8131,N_8335);
xnor U8527 (N_8527,N_7888,N_8342);
and U8528 (N_8528,N_7935,N_8389);
and U8529 (N_8529,N_7809,N_8144);
or U8530 (N_8530,N_8217,N_7948);
nand U8531 (N_8531,N_8289,N_7975);
or U8532 (N_8532,N_7966,N_8374);
and U8533 (N_8533,N_7863,N_7817);
and U8534 (N_8534,N_8209,N_8039);
and U8535 (N_8535,N_8040,N_7979);
nor U8536 (N_8536,N_8279,N_8327);
xor U8537 (N_8537,N_8104,N_8129);
nor U8538 (N_8538,N_8168,N_7848);
xor U8539 (N_8539,N_7928,N_8139);
xnor U8540 (N_8540,N_8382,N_8180);
nand U8541 (N_8541,N_8155,N_7907);
nor U8542 (N_8542,N_7815,N_8256);
nor U8543 (N_8543,N_8378,N_7860);
nand U8544 (N_8544,N_8395,N_7974);
and U8545 (N_8545,N_8398,N_7862);
nand U8546 (N_8546,N_8277,N_7986);
xnor U8547 (N_8547,N_7915,N_8328);
and U8548 (N_8548,N_7849,N_7938);
nor U8549 (N_8549,N_8071,N_7855);
or U8550 (N_8550,N_8253,N_8172);
nand U8551 (N_8551,N_7977,N_8216);
nand U8552 (N_8552,N_8127,N_8169);
and U8553 (N_8553,N_8247,N_8148);
and U8554 (N_8554,N_7953,N_8355);
and U8555 (N_8555,N_8027,N_8314);
nor U8556 (N_8556,N_8159,N_8083);
nor U8557 (N_8557,N_7856,N_8278);
or U8558 (N_8558,N_8003,N_7806);
xor U8559 (N_8559,N_8245,N_8196);
nor U8560 (N_8560,N_8154,N_8294);
and U8561 (N_8561,N_7884,N_8226);
xnor U8562 (N_8562,N_8162,N_8038);
xor U8563 (N_8563,N_8165,N_8093);
nor U8564 (N_8564,N_7960,N_8060);
or U8565 (N_8565,N_8397,N_8107);
nand U8566 (N_8566,N_8345,N_8016);
xnor U8567 (N_8567,N_8194,N_8211);
nand U8568 (N_8568,N_8356,N_8151);
and U8569 (N_8569,N_8364,N_8174);
xor U8570 (N_8570,N_7814,N_8237);
nor U8571 (N_8571,N_8390,N_8143);
xnor U8572 (N_8572,N_8052,N_8287);
and U8573 (N_8573,N_8282,N_8263);
nand U8574 (N_8574,N_8207,N_7940);
and U8575 (N_8575,N_7850,N_8179);
nand U8576 (N_8576,N_8185,N_8188);
or U8577 (N_8577,N_7825,N_8023);
and U8578 (N_8578,N_8212,N_8091);
and U8579 (N_8579,N_8349,N_8275);
or U8580 (N_8580,N_8284,N_8010);
and U8581 (N_8581,N_7801,N_8087);
and U8582 (N_8582,N_7949,N_7952);
xnor U8583 (N_8583,N_8032,N_8213);
nor U8584 (N_8584,N_8313,N_7802);
xnor U8585 (N_8585,N_7934,N_7813);
nor U8586 (N_8586,N_8291,N_7898);
nor U8587 (N_8587,N_7889,N_8103);
or U8588 (N_8588,N_8197,N_7939);
or U8589 (N_8589,N_7904,N_7982);
nand U8590 (N_8590,N_8170,N_8204);
nor U8591 (N_8591,N_8164,N_8048);
or U8592 (N_8592,N_7902,N_8184);
xor U8593 (N_8593,N_7840,N_8334);
nand U8594 (N_8594,N_8167,N_7908);
nand U8595 (N_8595,N_8115,N_8316);
and U8596 (N_8596,N_8376,N_8145);
nand U8597 (N_8597,N_8061,N_8105);
xor U8598 (N_8598,N_7842,N_8160);
or U8599 (N_8599,N_8086,N_8271);
and U8600 (N_8600,N_8260,N_8053);
xnor U8601 (N_8601,N_7976,N_8134);
nand U8602 (N_8602,N_7998,N_8254);
nor U8603 (N_8603,N_8269,N_8178);
xor U8604 (N_8604,N_8078,N_8261);
or U8605 (N_8605,N_8266,N_8050);
or U8606 (N_8606,N_7906,N_8058);
nand U8607 (N_8607,N_8077,N_8255);
nor U8608 (N_8608,N_8362,N_8161);
nor U8609 (N_8609,N_8126,N_8351);
xnor U8610 (N_8610,N_8081,N_8171);
nor U8611 (N_8611,N_8000,N_8280);
or U8612 (N_8612,N_8138,N_8006);
nand U8613 (N_8613,N_7967,N_7800);
and U8614 (N_8614,N_8020,N_8369);
nor U8615 (N_8615,N_8076,N_8225);
xnor U8616 (N_8616,N_7973,N_8163);
or U8617 (N_8617,N_8009,N_7882);
nor U8618 (N_8618,N_8022,N_7852);
nor U8619 (N_8619,N_7964,N_8276);
xnor U8620 (N_8620,N_8324,N_7920);
nand U8621 (N_8621,N_7892,N_8018);
and U8622 (N_8622,N_7838,N_7831);
xnor U8623 (N_8623,N_8153,N_8074);
and U8624 (N_8624,N_8128,N_8242);
or U8625 (N_8625,N_8117,N_7981);
nor U8626 (N_8626,N_8297,N_8059);
and U8627 (N_8627,N_8286,N_8283);
xnor U8628 (N_8628,N_8046,N_8368);
and U8629 (N_8629,N_8337,N_7984);
or U8630 (N_8630,N_8386,N_7878);
xnor U8631 (N_8631,N_8177,N_8125);
nor U8632 (N_8632,N_8224,N_7969);
or U8633 (N_8633,N_8252,N_7947);
and U8634 (N_8634,N_8329,N_8222);
xnor U8635 (N_8635,N_8228,N_8157);
xnor U8636 (N_8636,N_8310,N_7857);
or U8637 (N_8637,N_7866,N_7836);
or U8638 (N_8638,N_8111,N_8119);
and U8639 (N_8639,N_8005,N_7992);
nand U8640 (N_8640,N_7876,N_7925);
nor U8641 (N_8641,N_8067,N_8193);
xor U8642 (N_8642,N_8375,N_7950);
or U8643 (N_8643,N_7990,N_7854);
nor U8644 (N_8644,N_8227,N_8097);
nor U8645 (N_8645,N_8394,N_7830);
or U8646 (N_8646,N_8146,N_8033);
xnor U8647 (N_8647,N_8075,N_8202);
or U8648 (N_8648,N_7823,N_8221);
nor U8649 (N_8649,N_8220,N_7868);
nand U8650 (N_8650,N_7910,N_7899);
xor U8651 (N_8651,N_7931,N_8195);
xnor U8652 (N_8652,N_8108,N_7872);
or U8653 (N_8653,N_7924,N_7933);
and U8654 (N_8654,N_8363,N_8130);
or U8655 (N_8655,N_8358,N_8303);
xnor U8656 (N_8656,N_8352,N_7983);
xor U8657 (N_8657,N_8350,N_8385);
nor U8658 (N_8658,N_8028,N_7893);
nand U8659 (N_8659,N_7929,N_7843);
and U8660 (N_8660,N_8037,N_7803);
nor U8661 (N_8661,N_8031,N_7844);
or U8662 (N_8662,N_8295,N_8361);
or U8663 (N_8663,N_8123,N_7926);
nand U8664 (N_8664,N_7951,N_8183);
or U8665 (N_8665,N_8250,N_8175);
xor U8666 (N_8666,N_8001,N_8257);
xnor U8667 (N_8667,N_7987,N_8325);
nor U8668 (N_8668,N_7885,N_8315);
and U8669 (N_8669,N_8063,N_7895);
nor U8670 (N_8670,N_7864,N_8383);
or U8671 (N_8671,N_7911,N_8218);
nand U8672 (N_8672,N_8045,N_7820);
or U8673 (N_8673,N_7867,N_7965);
xnor U8674 (N_8674,N_8331,N_8073);
and U8675 (N_8675,N_7819,N_8137);
xor U8676 (N_8676,N_8206,N_8116);
nand U8677 (N_8677,N_8306,N_7970);
nand U8678 (N_8678,N_8201,N_7887);
xnor U8679 (N_8679,N_8377,N_8014);
or U8680 (N_8680,N_8229,N_8008);
xor U8681 (N_8681,N_8135,N_7891);
nor U8682 (N_8682,N_7923,N_7956);
and U8683 (N_8683,N_8305,N_8110);
nand U8684 (N_8684,N_7922,N_8396);
and U8685 (N_8685,N_8353,N_8021);
xnor U8686 (N_8686,N_7988,N_7886);
and U8687 (N_8687,N_8056,N_8062);
xor U8688 (N_8688,N_8090,N_8320);
or U8689 (N_8689,N_8262,N_7834);
xnor U8690 (N_8690,N_7968,N_8122);
nand U8691 (N_8691,N_8015,N_8041);
or U8692 (N_8692,N_7980,N_7917);
and U8693 (N_8693,N_8323,N_7955);
and U8694 (N_8694,N_8230,N_8149);
xor U8695 (N_8695,N_7993,N_8231);
nand U8696 (N_8696,N_8026,N_7994);
nand U8697 (N_8697,N_8338,N_7958);
nand U8698 (N_8698,N_8370,N_7807);
and U8699 (N_8699,N_8080,N_7832);
xor U8700 (N_8700,N_7957,N_8064);
xnor U8701 (N_8701,N_7899,N_7862);
nor U8702 (N_8702,N_7917,N_7972);
or U8703 (N_8703,N_8212,N_7899);
xor U8704 (N_8704,N_7856,N_7831);
or U8705 (N_8705,N_7987,N_8236);
or U8706 (N_8706,N_7915,N_8213);
or U8707 (N_8707,N_8251,N_8311);
nand U8708 (N_8708,N_8280,N_7977);
or U8709 (N_8709,N_8174,N_8204);
or U8710 (N_8710,N_8354,N_7828);
nand U8711 (N_8711,N_8240,N_8333);
nor U8712 (N_8712,N_7854,N_7816);
nand U8713 (N_8713,N_7818,N_7946);
nor U8714 (N_8714,N_8075,N_8167);
and U8715 (N_8715,N_8126,N_8036);
and U8716 (N_8716,N_8237,N_8012);
nor U8717 (N_8717,N_8369,N_8135);
or U8718 (N_8718,N_8231,N_8306);
nor U8719 (N_8719,N_8141,N_8383);
nand U8720 (N_8720,N_8172,N_7819);
and U8721 (N_8721,N_8040,N_8146);
or U8722 (N_8722,N_7804,N_8354);
xnor U8723 (N_8723,N_8294,N_8038);
or U8724 (N_8724,N_7905,N_8229);
nand U8725 (N_8725,N_8064,N_8163);
or U8726 (N_8726,N_8022,N_8166);
nand U8727 (N_8727,N_8193,N_8045);
nor U8728 (N_8728,N_8272,N_8230);
xor U8729 (N_8729,N_8124,N_8240);
and U8730 (N_8730,N_8276,N_7986);
and U8731 (N_8731,N_8394,N_7982);
nand U8732 (N_8732,N_7997,N_7872);
nor U8733 (N_8733,N_8315,N_8198);
nor U8734 (N_8734,N_7832,N_7913);
and U8735 (N_8735,N_8000,N_8130);
and U8736 (N_8736,N_7924,N_8216);
nor U8737 (N_8737,N_7978,N_8010);
and U8738 (N_8738,N_8228,N_8122);
and U8739 (N_8739,N_8172,N_7996);
xnor U8740 (N_8740,N_7999,N_8188);
xnor U8741 (N_8741,N_8397,N_8338);
nand U8742 (N_8742,N_8094,N_8151);
xor U8743 (N_8743,N_8290,N_8170);
nand U8744 (N_8744,N_8304,N_8224);
nor U8745 (N_8745,N_8127,N_8397);
or U8746 (N_8746,N_8070,N_8259);
nand U8747 (N_8747,N_8248,N_8193);
nand U8748 (N_8748,N_8373,N_8253);
or U8749 (N_8749,N_8180,N_8286);
nand U8750 (N_8750,N_8001,N_7884);
nand U8751 (N_8751,N_8311,N_8248);
and U8752 (N_8752,N_7892,N_8329);
nor U8753 (N_8753,N_8299,N_8366);
nand U8754 (N_8754,N_7986,N_8347);
nand U8755 (N_8755,N_8135,N_7933);
nor U8756 (N_8756,N_8281,N_8384);
or U8757 (N_8757,N_8277,N_8084);
or U8758 (N_8758,N_8366,N_7860);
nor U8759 (N_8759,N_7850,N_8197);
and U8760 (N_8760,N_7858,N_7985);
or U8761 (N_8761,N_7829,N_8232);
nor U8762 (N_8762,N_7931,N_8121);
xor U8763 (N_8763,N_7974,N_8223);
nand U8764 (N_8764,N_7938,N_8126);
xnor U8765 (N_8765,N_7890,N_8344);
nand U8766 (N_8766,N_8248,N_8266);
or U8767 (N_8767,N_8328,N_8280);
and U8768 (N_8768,N_7935,N_7978);
and U8769 (N_8769,N_7918,N_8181);
xor U8770 (N_8770,N_8044,N_7954);
nor U8771 (N_8771,N_7878,N_8299);
nor U8772 (N_8772,N_8141,N_7911);
and U8773 (N_8773,N_8339,N_8226);
nand U8774 (N_8774,N_8115,N_8178);
or U8775 (N_8775,N_8235,N_7909);
nor U8776 (N_8776,N_8292,N_8369);
and U8777 (N_8777,N_7845,N_7954);
and U8778 (N_8778,N_8252,N_8143);
or U8779 (N_8779,N_8298,N_7984);
nor U8780 (N_8780,N_8311,N_8094);
nand U8781 (N_8781,N_8213,N_8171);
nand U8782 (N_8782,N_7912,N_8194);
nor U8783 (N_8783,N_8020,N_7912);
or U8784 (N_8784,N_7829,N_8229);
or U8785 (N_8785,N_8123,N_8245);
xor U8786 (N_8786,N_8136,N_7986);
xnor U8787 (N_8787,N_8072,N_8211);
xor U8788 (N_8788,N_8189,N_8181);
nor U8789 (N_8789,N_8312,N_8105);
nand U8790 (N_8790,N_8251,N_7971);
nor U8791 (N_8791,N_7918,N_7991);
and U8792 (N_8792,N_8089,N_8248);
and U8793 (N_8793,N_8311,N_8330);
and U8794 (N_8794,N_7849,N_7980);
and U8795 (N_8795,N_8362,N_8220);
or U8796 (N_8796,N_8305,N_8202);
and U8797 (N_8797,N_8190,N_8165);
and U8798 (N_8798,N_8309,N_7910);
nand U8799 (N_8799,N_8103,N_8206);
and U8800 (N_8800,N_8346,N_8377);
xnor U8801 (N_8801,N_8020,N_8388);
or U8802 (N_8802,N_8091,N_7932);
xor U8803 (N_8803,N_8246,N_7804);
xnor U8804 (N_8804,N_8219,N_8277);
or U8805 (N_8805,N_8195,N_7976);
nor U8806 (N_8806,N_7892,N_8251);
nand U8807 (N_8807,N_7894,N_8165);
nor U8808 (N_8808,N_7930,N_8228);
nor U8809 (N_8809,N_8239,N_8350);
and U8810 (N_8810,N_8377,N_8340);
nand U8811 (N_8811,N_8008,N_7995);
and U8812 (N_8812,N_8072,N_8015);
or U8813 (N_8813,N_7803,N_8148);
nand U8814 (N_8814,N_7827,N_7954);
or U8815 (N_8815,N_8228,N_7937);
nor U8816 (N_8816,N_8083,N_8122);
nand U8817 (N_8817,N_7909,N_8022);
xor U8818 (N_8818,N_8161,N_7831);
and U8819 (N_8819,N_8109,N_8087);
and U8820 (N_8820,N_8015,N_8334);
or U8821 (N_8821,N_8140,N_8391);
or U8822 (N_8822,N_8084,N_7836);
and U8823 (N_8823,N_8071,N_8373);
nand U8824 (N_8824,N_7960,N_7810);
or U8825 (N_8825,N_8115,N_8392);
xnor U8826 (N_8826,N_8165,N_8255);
nor U8827 (N_8827,N_8323,N_7936);
nor U8828 (N_8828,N_7958,N_8116);
nor U8829 (N_8829,N_8188,N_7806);
xnor U8830 (N_8830,N_7906,N_8230);
nor U8831 (N_8831,N_8347,N_8187);
and U8832 (N_8832,N_8231,N_8378);
or U8833 (N_8833,N_7962,N_8062);
nand U8834 (N_8834,N_7841,N_8355);
nor U8835 (N_8835,N_8021,N_8083);
and U8836 (N_8836,N_7939,N_7934);
and U8837 (N_8837,N_8372,N_8043);
and U8838 (N_8838,N_8117,N_8073);
or U8839 (N_8839,N_8010,N_8341);
or U8840 (N_8840,N_8058,N_7931);
and U8841 (N_8841,N_8227,N_8269);
or U8842 (N_8842,N_7986,N_7951);
and U8843 (N_8843,N_7907,N_8376);
or U8844 (N_8844,N_7816,N_7813);
or U8845 (N_8845,N_7974,N_8128);
and U8846 (N_8846,N_8389,N_7843);
or U8847 (N_8847,N_7908,N_8098);
and U8848 (N_8848,N_7837,N_8079);
nand U8849 (N_8849,N_8094,N_7993);
or U8850 (N_8850,N_7869,N_7988);
nand U8851 (N_8851,N_8175,N_8024);
or U8852 (N_8852,N_7806,N_7909);
nor U8853 (N_8853,N_8005,N_8034);
and U8854 (N_8854,N_8358,N_7850);
or U8855 (N_8855,N_7869,N_8358);
xnor U8856 (N_8856,N_8191,N_8125);
nand U8857 (N_8857,N_8284,N_8327);
nor U8858 (N_8858,N_8088,N_8035);
nor U8859 (N_8859,N_8318,N_8348);
and U8860 (N_8860,N_8399,N_8103);
or U8861 (N_8861,N_8088,N_8078);
nand U8862 (N_8862,N_8372,N_8008);
and U8863 (N_8863,N_8102,N_7980);
nand U8864 (N_8864,N_8089,N_8066);
xor U8865 (N_8865,N_8024,N_7838);
or U8866 (N_8866,N_8374,N_8366);
xor U8867 (N_8867,N_8207,N_8396);
nand U8868 (N_8868,N_8288,N_8231);
nor U8869 (N_8869,N_7847,N_8254);
nand U8870 (N_8870,N_8384,N_7980);
nand U8871 (N_8871,N_8044,N_7801);
and U8872 (N_8872,N_8188,N_7874);
or U8873 (N_8873,N_7882,N_8299);
xor U8874 (N_8874,N_8268,N_8223);
nand U8875 (N_8875,N_8367,N_8080);
xnor U8876 (N_8876,N_8179,N_8012);
nor U8877 (N_8877,N_8231,N_8048);
xnor U8878 (N_8878,N_8258,N_8241);
nor U8879 (N_8879,N_8399,N_8363);
and U8880 (N_8880,N_8023,N_8307);
xor U8881 (N_8881,N_8023,N_7876);
or U8882 (N_8882,N_8204,N_7802);
xnor U8883 (N_8883,N_8337,N_8022);
xor U8884 (N_8884,N_8006,N_8218);
or U8885 (N_8885,N_8009,N_8375);
nand U8886 (N_8886,N_7962,N_7976);
or U8887 (N_8887,N_8088,N_8326);
xnor U8888 (N_8888,N_8298,N_7961);
xnor U8889 (N_8889,N_8251,N_8079);
and U8890 (N_8890,N_8276,N_8300);
xnor U8891 (N_8891,N_8258,N_8319);
or U8892 (N_8892,N_8326,N_7967);
xor U8893 (N_8893,N_8264,N_8103);
nor U8894 (N_8894,N_8140,N_7885);
nand U8895 (N_8895,N_8307,N_8300);
xor U8896 (N_8896,N_8047,N_7849);
nor U8897 (N_8897,N_7860,N_8148);
nand U8898 (N_8898,N_8049,N_8246);
nor U8899 (N_8899,N_8302,N_8213);
nand U8900 (N_8900,N_8260,N_8013);
nand U8901 (N_8901,N_8180,N_8173);
nand U8902 (N_8902,N_8197,N_7852);
nor U8903 (N_8903,N_7862,N_8041);
or U8904 (N_8904,N_8227,N_8180);
nor U8905 (N_8905,N_8121,N_8086);
or U8906 (N_8906,N_7819,N_7914);
nor U8907 (N_8907,N_8228,N_7922);
and U8908 (N_8908,N_8370,N_7912);
xor U8909 (N_8909,N_8106,N_7890);
or U8910 (N_8910,N_8025,N_7815);
or U8911 (N_8911,N_8364,N_8370);
nand U8912 (N_8912,N_7999,N_7991);
xor U8913 (N_8913,N_8035,N_7910);
nand U8914 (N_8914,N_7854,N_8199);
nor U8915 (N_8915,N_8063,N_8206);
nand U8916 (N_8916,N_7843,N_8272);
and U8917 (N_8917,N_8378,N_8205);
nor U8918 (N_8918,N_7894,N_8055);
nor U8919 (N_8919,N_8165,N_8262);
nand U8920 (N_8920,N_8056,N_8318);
nand U8921 (N_8921,N_8232,N_8364);
or U8922 (N_8922,N_7815,N_8328);
and U8923 (N_8923,N_7832,N_7997);
and U8924 (N_8924,N_8395,N_7802);
or U8925 (N_8925,N_8325,N_8365);
nor U8926 (N_8926,N_8226,N_8172);
xor U8927 (N_8927,N_8225,N_8397);
nor U8928 (N_8928,N_8376,N_7884);
nand U8929 (N_8929,N_8387,N_8277);
nor U8930 (N_8930,N_8177,N_7805);
xor U8931 (N_8931,N_8354,N_8367);
nor U8932 (N_8932,N_8152,N_8301);
nor U8933 (N_8933,N_8288,N_8091);
and U8934 (N_8934,N_8239,N_8053);
xnor U8935 (N_8935,N_7914,N_8242);
nor U8936 (N_8936,N_8049,N_8228);
and U8937 (N_8937,N_7823,N_8385);
nand U8938 (N_8938,N_8159,N_7934);
and U8939 (N_8939,N_8018,N_7908);
nand U8940 (N_8940,N_8247,N_8090);
nand U8941 (N_8941,N_7916,N_8091);
or U8942 (N_8942,N_7804,N_8341);
and U8943 (N_8943,N_7933,N_8027);
nand U8944 (N_8944,N_7833,N_8227);
xnor U8945 (N_8945,N_8273,N_7842);
nand U8946 (N_8946,N_8147,N_8326);
and U8947 (N_8947,N_8377,N_7903);
or U8948 (N_8948,N_7962,N_8077);
or U8949 (N_8949,N_8141,N_8202);
xor U8950 (N_8950,N_7875,N_7940);
or U8951 (N_8951,N_7912,N_8384);
xnor U8952 (N_8952,N_8082,N_7883);
and U8953 (N_8953,N_7969,N_7912);
nor U8954 (N_8954,N_8288,N_8083);
nor U8955 (N_8955,N_7942,N_8040);
and U8956 (N_8956,N_8069,N_8155);
nand U8957 (N_8957,N_7821,N_8193);
nor U8958 (N_8958,N_8295,N_7897);
nor U8959 (N_8959,N_8182,N_8307);
or U8960 (N_8960,N_8023,N_8044);
and U8961 (N_8961,N_8342,N_7962);
or U8962 (N_8962,N_8357,N_7926);
nand U8963 (N_8963,N_8349,N_8391);
xnor U8964 (N_8964,N_7816,N_7819);
or U8965 (N_8965,N_8199,N_8171);
nand U8966 (N_8966,N_8290,N_7948);
nor U8967 (N_8967,N_8269,N_8368);
nor U8968 (N_8968,N_8319,N_8326);
xnor U8969 (N_8969,N_8365,N_8245);
and U8970 (N_8970,N_8072,N_8330);
nand U8971 (N_8971,N_8185,N_7837);
xor U8972 (N_8972,N_7990,N_8208);
nand U8973 (N_8973,N_8366,N_8315);
nand U8974 (N_8974,N_8086,N_8065);
nand U8975 (N_8975,N_7994,N_8042);
or U8976 (N_8976,N_8338,N_8050);
nand U8977 (N_8977,N_8203,N_8134);
xor U8978 (N_8978,N_7816,N_7974);
or U8979 (N_8979,N_7858,N_7993);
and U8980 (N_8980,N_8009,N_8115);
xnor U8981 (N_8981,N_8248,N_8287);
xor U8982 (N_8982,N_7992,N_7892);
or U8983 (N_8983,N_7927,N_8080);
xnor U8984 (N_8984,N_7926,N_8399);
nor U8985 (N_8985,N_7848,N_7857);
and U8986 (N_8986,N_8188,N_8083);
or U8987 (N_8987,N_8353,N_8102);
xnor U8988 (N_8988,N_8180,N_8261);
nor U8989 (N_8989,N_8304,N_8026);
and U8990 (N_8990,N_8000,N_7832);
xnor U8991 (N_8991,N_7865,N_8082);
nor U8992 (N_8992,N_7880,N_8265);
and U8993 (N_8993,N_8128,N_8058);
nor U8994 (N_8994,N_8061,N_8068);
or U8995 (N_8995,N_8062,N_8055);
xor U8996 (N_8996,N_8052,N_8069);
nor U8997 (N_8997,N_7883,N_8331);
or U8998 (N_8998,N_8365,N_8243);
nor U8999 (N_8999,N_8257,N_7966);
nand U9000 (N_9000,N_8615,N_8450);
and U9001 (N_9001,N_8406,N_8432);
nand U9002 (N_9002,N_8880,N_8889);
and U9003 (N_9003,N_8991,N_8545);
nor U9004 (N_9004,N_8617,N_8518);
and U9005 (N_9005,N_8431,N_8820);
nand U9006 (N_9006,N_8415,N_8500);
or U9007 (N_9007,N_8683,N_8954);
nand U9008 (N_9008,N_8596,N_8412);
and U9009 (N_9009,N_8514,N_8665);
nand U9010 (N_9010,N_8928,N_8802);
xor U9011 (N_9011,N_8911,N_8945);
xor U9012 (N_9012,N_8987,N_8635);
nor U9013 (N_9013,N_8875,N_8738);
and U9014 (N_9014,N_8976,N_8739);
or U9015 (N_9015,N_8582,N_8870);
xnor U9016 (N_9016,N_8805,N_8819);
or U9017 (N_9017,N_8498,N_8686);
nor U9018 (N_9018,N_8897,N_8599);
or U9019 (N_9019,N_8790,N_8536);
nor U9020 (N_9020,N_8562,N_8751);
xor U9021 (N_9021,N_8939,N_8730);
nor U9022 (N_9022,N_8898,N_8999);
or U9023 (N_9023,N_8851,N_8970);
xor U9024 (N_9024,N_8586,N_8769);
xor U9025 (N_9025,N_8778,N_8620);
xor U9026 (N_9026,N_8784,N_8994);
or U9027 (N_9027,N_8828,N_8534);
and U9028 (N_9028,N_8591,N_8749);
xnor U9029 (N_9029,N_8499,N_8728);
xor U9030 (N_9030,N_8697,N_8678);
or U9031 (N_9031,N_8888,N_8566);
nor U9032 (N_9032,N_8800,N_8465);
nor U9033 (N_9033,N_8578,N_8853);
nand U9034 (N_9034,N_8677,N_8867);
and U9035 (N_9035,N_8878,N_8899);
or U9036 (N_9036,N_8680,N_8983);
xnor U9037 (N_9037,N_8786,N_8447);
or U9038 (N_9038,N_8919,N_8785);
and U9039 (N_9039,N_8882,N_8905);
or U9040 (N_9040,N_8794,N_8977);
or U9041 (N_9041,N_8759,N_8768);
xnor U9042 (N_9042,N_8410,N_8585);
xor U9043 (N_9043,N_8468,N_8424);
and U9044 (N_9044,N_8703,N_8411);
or U9045 (N_9045,N_8868,N_8670);
nand U9046 (N_9046,N_8496,N_8404);
and U9047 (N_9047,N_8764,N_8509);
and U9048 (N_9048,N_8783,N_8681);
nand U9049 (N_9049,N_8832,N_8548);
nand U9050 (N_9050,N_8829,N_8957);
nor U9051 (N_9051,N_8843,N_8955);
and U9052 (N_9052,N_8540,N_8815);
xnor U9053 (N_9053,N_8484,N_8572);
nand U9054 (N_9054,N_8873,N_8717);
and U9055 (N_9055,N_8732,N_8634);
or U9056 (N_9056,N_8542,N_8936);
or U9057 (N_9057,N_8975,N_8906);
nor U9058 (N_9058,N_8440,N_8709);
nand U9059 (N_9059,N_8520,N_8750);
nor U9060 (N_9060,N_8611,N_8511);
nor U9061 (N_9061,N_8948,N_8527);
xnor U9062 (N_9062,N_8667,N_8877);
and U9063 (N_9063,N_8429,N_8672);
and U9064 (N_9064,N_8477,N_8487);
nor U9065 (N_9065,N_8806,N_8831);
or U9066 (N_9066,N_8973,N_8796);
and U9067 (N_9067,N_8760,N_8910);
nor U9068 (N_9068,N_8598,N_8425);
nand U9069 (N_9069,N_8864,N_8510);
xor U9070 (N_9070,N_8782,N_8671);
nand U9071 (N_9071,N_8731,N_8743);
xnor U9072 (N_9072,N_8658,N_8524);
and U9073 (N_9073,N_8933,N_8619);
xnor U9074 (N_9074,N_8988,N_8687);
nor U9075 (N_9075,N_8744,N_8736);
xor U9076 (N_9076,N_8834,N_8632);
nand U9077 (N_9077,N_8644,N_8814);
and U9078 (N_9078,N_8418,N_8961);
or U9079 (N_9079,N_8812,N_8921);
or U9080 (N_9080,N_8584,N_8435);
nand U9081 (N_9081,N_8696,N_8701);
or U9082 (N_9082,N_8923,N_8568);
xnor U9083 (N_9083,N_8869,N_8444);
and U9084 (N_9084,N_8449,N_8443);
xor U9085 (N_9085,N_8689,N_8439);
or U9086 (N_9086,N_8559,N_8849);
xor U9087 (N_9087,N_8879,N_8756);
nor U9088 (N_9088,N_8525,N_8846);
nor U9089 (N_9089,N_8475,N_8663);
nor U9090 (N_9090,N_8699,N_8716);
or U9091 (N_9091,N_8854,N_8929);
or U9092 (N_9092,N_8734,N_8633);
or U9093 (N_9093,N_8592,N_8902);
and U9094 (N_9094,N_8638,N_8629);
nor U9095 (N_9095,N_8795,N_8940);
nand U9096 (N_9096,N_8807,N_8771);
nor U9097 (N_9097,N_8555,N_8816);
or U9098 (N_9098,N_8522,N_8420);
xor U9099 (N_9099,N_8452,N_8554);
xnor U9100 (N_9100,N_8881,N_8925);
or U9101 (N_9101,N_8523,N_8883);
and U9102 (N_9102,N_8579,N_8922);
nor U9103 (N_9103,N_8757,N_8456);
or U9104 (N_9104,N_8413,N_8727);
and U9105 (N_9105,N_8789,N_8946);
and U9106 (N_9106,N_8996,N_8886);
and U9107 (N_9107,N_8947,N_8564);
or U9108 (N_9108,N_8859,N_8551);
and U9109 (N_9109,N_8469,N_8981);
and U9110 (N_9110,N_8588,N_8984);
or U9111 (N_9111,N_8850,N_8521);
nand U9112 (N_9112,N_8648,N_8623);
or U9113 (N_9113,N_8824,N_8942);
nand U9114 (N_9114,N_8676,N_8647);
nor U9115 (N_9115,N_8405,N_8715);
nor U9116 (N_9116,N_8752,N_8773);
or U9117 (N_9117,N_8914,N_8417);
nand U9118 (N_9118,N_8855,N_8426);
or U9119 (N_9119,N_8614,N_8753);
and U9120 (N_9120,N_8577,N_8645);
xnor U9121 (N_9121,N_8995,N_8594);
nor U9122 (N_9122,N_8613,N_8721);
xor U9123 (N_9123,N_8442,N_8941);
nor U9124 (N_9124,N_8493,N_8628);
and U9125 (N_9125,N_8966,N_8664);
xnor U9126 (N_9126,N_8747,N_8655);
nor U9127 (N_9127,N_8675,N_8978);
and U9128 (N_9128,N_8561,N_8626);
or U9129 (N_9129,N_8400,N_8421);
nor U9130 (N_9130,N_8479,N_8958);
nor U9131 (N_9131,N_8949,N_8746);
and U9132 (N_9132,N_8822,N_8865);
or U9133 (N_9133,N_8506,N_8950);
nor U9134 (N_9134,N_8871,N_8702);
nor U9135 (N_9135,N_8766,N_8863);
or U9136 (N_9136,N_8791,N_8809);
xnor U9137 (N_9137,N_8470,N_8932);
or U9138 (N_9138,N_8430,N_8765);
and U9139 (N_9139,N_8774,N_8489);
and U9140 (N_9140,N_8720,N_8856);
nor U9141 (N_9141,N_8595,N_8685);
nand U9142 (N_9142,N_8546,N_8916);
and U9143 (N_9143,N_8445,N_8616);
nand U9144 (N_9144,N_8740,N_8971);
xor U9145 (N_9145,N_8913,N_8488);
nand U9146 (N_9146,N_8963,N_8688);
and U9147 (N_9147,N_8446,N_8642);
nand U9148 (N_9148,N_8893,N_8472);
xor U9149 (N_9149,N_8714,N_8494);
xnor U9150 (N_9150,N_8847,N_8967);
nor U9151 (N_9151,N_8894,N_8486);
or U9152 (N_9152,N_8901,N_8840);
nand U9153 (N_9153,N_8907,N_8758);
or U9154 (N_9154,N_8462,N_8982);
or U9155 (N_9155,N_8917,N_8892);
nor U9156 (N_9156,N_8567,N_8985);
and U9157 (N_9157,N_8508,N_8735);
and U9158 (N_9158,N_8640,N_8575);
nor U9159 (N_9159,N_8428,N_8772);
nand U9160 (N_9160,N_8679,N_8654);
nor U9161 (N_9161,N_8622,N_8833);
or U9162 (N_9162,N_8643,N_8700);
or U9163 (N_9163,N_8825,N_8550);
and U9164 (N_9164,N_8581,N_8974);
nand U9165 (N_9165,N_8777,N_8968);
and U9166 (N_9166,N_8733,N_8725);
nand U9167 (N_9167,N_8476,N_8872);
and U9168 (N_9168,N_8636,N_8501);
nor U9169 (N_9169,N_8433,N_8682);
nand U9170 (N_9170,N_8775,N_8673);
or U9171 (N_9171,N_8798,N_8920);
xor U9172 (N_9172,N_8660,N_8637);
xnor U9173 (N_9173,N_8528,N_8454);
or U9174 (N_9174,N_8571,N_8729);
xor U9175 (N_9175,N_8674,N_8537);
or U9176 (N_9176,N_8801,N_8693);
and U9177 (N_9177,N_8770,N_8866);
and U9178 (N_9178,N_8530,N_8504);
and U9179 (N_9179,N_8817,N_8531);
nor U9180 (N_9180,N_8538,N_8533);
nor U9181 (N_9181,N_8659,N_8558);
or U9182 (N_9182,N_8606,N_8603);
or U9183 (N_9183,N_8818,N_8839);
xnor U9184 (N_9184,N_8964,N_8482);
nor U9185 (N_9185,N_8560,N_8926);
nand U9186 (N_9186,N_8896,N_8780);
nor U9187 (N_9187,N_8838,N_8997);
xnor U9188 (N_9188,N_8990,N_8669);
or U9189 (N_9189,N_8705,N_8960);
and U9190 (N_9190,N_8952,N_8480);
nand U9191 (N_9191,N_8793,N_8419);
or U9192 (N_9192,N_8587,N_8767);
or U9193 (N_9193,N_8503,N_8556);
and U9194 (N_9194,N_8438,N_8737);
and U9195 (N_9195,N_8485,N_8827);
nand U9196 (N_9196,N_8535,N_8653);
and U9197 (N_9197,N_8631,N_8726);
nor U9198 (N_9198,N_8808,N_8691);
xnor U9199 (N_9199,N_8908,N_8719);
nor U9200 (N_9200,N_8836,N_8745);
or U9201 (N_9201,N_8570,N_8403);
and U9202 (N_9202,N_8876,N_8507);
or U9203 (N_9203,N_8861,N_8437);
or U9204 (N_9204,N_8458,N_8972);
xnor U9205 (N_9205,N_8912,N_8505);
xor U9206 (N_9206,N_8857,N_8666);
xor U9207 (N_9207,N_8762,N_8483);
nor U9208 (N_9208,N_8407,N_8993);
nand U9209 (N_9209,N_8969,N_8512);
xor U9210 (N_9210,N_8965,N_8414);
xnor U9211 (N_9211,N_8884,N_8448);
nor U9212 (N_9212,N_8776,N_8455);
or U9213 (N_9213,N_8552,N_8694);
xnor U9214 (N_9214,N_8549,N_8698);
or U9215 (N_9215,N_8401,N_8529);
nand U9216 (N_9216,N_8710,N_8610);
nand U9217 (N_9217,N_8516,N_8837);
xor U9218 (N_9218,N_8605,N_8662);
and U9219 (N_9219,N_8779,N_8848);
nand U9220 (N_9220,N_8541,N_8463);
nor U9221 (N_9221,N_8422,N_8711);
or U9222 (N_9222,N_8813,N_8722);
xnor U9223 (N_9223,N_8656,N_8630);
nor U9224 (N_9224,N_8600,N_8885);
or U9225 (N_9225,N_8434,N_8574);
nor U9226 (N_9226,N_8755,N_8989);
nor U9227 (N_9227,N_8427,N_8589);
xor U9228 (N_9228,N_8491,N_8909);
xnor U9229 (N_9229,N_8895,N_8951);
nand U9230 (N_9230,N_8441,N_8986);
nor U9231 (N_9231,N_8704,N_8607);
xor U9232 (N_9232,N_8841,N_8690);
and U9233 (N_9233,N_8748,N_8810);
or U9234 (N_9234,N_8497,N_8826);
or U9235 (N_9235,N_8953,N_8597);
xor U9236 (N_9236,N_8845,N_8891);
or U9237 (N_9237,N_8513,N_8517);
nor U9238 (N_9238,N_8924,N_8918);
xor U9239 (N_9239,N_8763,N_8708);
and U9240 (N_9240,N_8706,N_8811);
nor U9241 (N_9241,N_8641,N_8937);
nor U9242 (N_9242,N_8646,N_8569);
nand U9243 (N_9243,N_8539,N_8478);
nor U9244 (N_9244,N_8639,N_8565);
and U9245 (N_9245,N_8423,N_8580);
nand U9246 (N_9246,N_8787,N_8821);
xor U9247 (N_9247,N_8612,N_8842);
and U9248 (N_9248,N_8803,N_8461);
xor U9249 (N_9249,N_8621,N_8980);
nor U9250 (N_9250,N_8601,N_8695);
and U9251 (N_9251,N_8915,N_8904);
xnor U9252 (N_9252,N_8609,N_8627);
nand U9253 (N_9253,N_8979,N_8451);
nor U9254 (N_9254,N_8887,N_8502);
nor U9255 (N_9255,N_8652,N_8944);
nor U9256 (N_9256,N_8657,N_8473);
nand U9257 (N_9257,N_8495,N_8835);
nand U9258 (N_9258,N_8618,N_8799);
nand U9259 (N_9259,N_8724,N_8625);
nor U9260 (N_9260,N_8935,N_8466);
xor U9261 (N_9261,N_8474,N_8862);
nand U9262 (N_9262,N_8467,N_8934);
nand U9263 (N_9263,N_8741,N_8436);
nor U9264 (N_9264,N_8707,N_8651);
xnor U9265 (N_9265,N_8547,N_8649);
nor U9266 (N_9266,N_8858,N_8797);
or U9267 (N_9267,N_8792,N_8563);
or U9268 (N_9268,N_8713,N_8692);
nand U9269 (N_9269,N_8712,N_8471);
or U9270 (N_9270,N_8874,N_8416);
xnor U9271 (N_9271,N_8938,N_8742);
or U9272 (N_9272,N_8804,N_8823);
nor U9273 (N_9273,N_8464,N_8481);
xor U9274 (N_9274,N_8408,N_8723);
xor U9275 (N_9275,N_8624,N_8962);
nand U9276 (N_9276,N_8998,N_8602);
xnor U9277 (N_9277,N_8532,N_8890);
xnor U9278 (N_9278,N_8402,N_8576);
and U9279 (N_9279,N_8830,N_8459);
nor U9280 (N_9280,N_8515,N_8604);
nor U9281 (N_9281,N_8526,N_8788);
and U9282 (N_9282,N_8927,N_8959);
and U9283 (N_9283,N_8409,N_8718);
nand U9284 (N_9284,N_8544,N_8956);
and U9285 (N_9285,N_8492,N_8453);
nor U9286 (N_9286,N_8593,N_8852);
or U9287 (N_9287,N_8860,N_8761);
nand U9288 (N_9288,N_8930,N_8931);
and U9289 (N_9289,N_8943,N_8781);
nand U9290 (N_9290,N_8844,N_8519);
or U9291 (N_9291,N_8590,N_8543);
xor U9292 (N_9292,N_8903,N_8573);
xnor U9293 (N_9293,N_8557,N_8650);
nor U9294 (N_9294,N_8668,N_8583);
nand U9295 (N_9295,N_8490,N_8553);
nand U9296 (N_9296,N_8457,N_8460);
and U9297 (N_9297,N_8661,N_8608);
nor U9298 (N_9298,N_8684,N_8754);
nor U9299 (N_9299,N_8992,N_8900);
nor U9300 (N_9300,N_8417,N_8488);
xnor U9301 (N_9301,N_8821,N_8956);
nor U9302 (N_9302,N_8872,N_8890);
xor U9303 (N_9303,N_8949,N_8668);
nor U9304 (N_9304,N_8747,N_8549);
and U9305 (N_9305,N_8840,N_8528);
nand U9306 (N_9306,N_8549,N_8817);
or U9307 (N_9307,N_8818,N_8718);
nand U9308 (N_9308,N_8619,N_8517);
and U9309 (N_9309,N_8467,N_8739);
xnor U9310 (N_9310,N_8784,N_8415);
and U9311 (N_9311,N_8529,N_8431);
nor U9312 (N_9312,N_8410,N_8658);
nand U9313 (N_9313,N_8516,N_8822);
xnor U9314 (N_9314,N_8960,N_8569);
and U9315 (N_9315,N_8705,N_8947);
nor U9316 (N_9316,N_8753,N_8788);
xor U9317 (N_9317,N_8701,N_8434);
nor U9318 (N_9318,N_8921,N_8950);
xor U9319 (N_9319,N_8755,N_8902);
or U9320 (N_9320,N_8823,N_8655);
or U9321 (N_9321,N_8546,N_8774);
nor U9322 (N_9322,N_8698,N_8944);
and U9323 (N_9323,N_8626,N_8728);
nor U9324 (N_9324,N_8429,N_8400);
nor U9325 (N_9325,N_8584,N_8454);
xnor U9326 (N_9326,N_8916,N_8892);
nand U9327 (N_9327,N_8942,N_8491);
nor U9328 (N_9328,N_8968,N_8674);
xnor U9329 (N_9329,N_8948,N_8573);
or U9330 (N_9330,N_8795,N_8956);
nand U9331 (N_9331,N_8555,N_8818);
xor U9332 (N_9332,N_8677,N_8545);
nand U9333 (N_9333,N_8823,N_8571);
nor U9334 (N_9334,N_8669,N_8963);
nand U9335 (N_9335,N_8538,N_8703);
xnor U9336 (N_9336,N_8811,N_8561);
xnor U9337 (N_9337,N_8748,N_8752);
xor U9338 (N_9338,N_8960,N_8805);
xor U9339 (N_9339,N_8731,N_8604);
nand U9340 (N_9340,N_8776,N_8427);
or U9341 (N_9341,N_8970,N_8531);
nand U9342 (N_9342,N_8589,N_8727);
or U9343 (N_9343,N_8714,N_8627);
and U9344 (N_9344,N_8954,N_8590);
or U9345 (N_9345,N_8648,N_8553);
nor U9346 (N_9346,N_8712,N_8657);
and U9347 (N_9347,N_8895,N_8713);
or U9348 (N_9348,N_8628,N_8946);
or U9349 (N_9349,N_8613,N_8697);
and U9350 (N_9350,N_8956,N_8453);
and U9351 (N_9351,N_8702,N_8786);
nor U9352 (N_9352,N_8744,N_8908);
nor U9353 (N_9353,N_8762,N_8884);
nand U9354 (N_9354,N_8563,N_8980);
or U9355 (N_9355,N_8696,N_8831);
xor U9356 (N_9356,N_8707,N_8781);
or U9357 (N_9357,N_8510,N_8862);
nand U9358 (N_9358,N_8708,N_8688);
nand U9359 (N_9359,N_8920,N_8800);
and U9360 (N_9360,N_8552,N_8548);
nor U9361 (N_9361,N_8441,N_8508);
and U9362 (N_9362,N_8405,N_8476);
or U9363 (N_9363,N_8698,N_8757);
and U9364 (N_9364,N_8844,N_8907);
nor U9365 (N_9365,N_8494,N_8656);
nand U9366 (N_9366,N_8614,N_8721);
xor U9367 (N_9367,N_8610,N_8446);
xor U9368 (N_9368,N_8651,N_8916);
nor U9369 (N_9369,N_8457,N_8848);
xnor U9370 (N_9370,N_8510,N_8903);
or U9371 (N_9371,N_8703,N_8822);
nand U9372 (N_9372,N_8746,N_8614);
nand U9373 (N_9373,N_8565,N_8981);
xnor U9374 (N_9374,N_8959,N_8416);
xor U9375 (N_9375,N_8939,N_8648);
or U9376 (N_9376,N_8989,N_8437);
and U9377 (N_9377,N_8940,N_8881);
xor U9378 (N_9378,N_8780,N_8447);
nand U9379 (N_9379,N_8958,N_8626);
and U9380 (N_9380,N_8948,N_8985);
xnor U9381 (N_9381,N_8424,N_8987);
nor U9382 (N_9382,N_8419,N_8469);
and U9383 (N_9383,N_8778,N_8625);
and U9384 (N_9384,N_8809,N_8698);
xor U9385 (N_9385,N_8650,N_8540);
or U9386 (N_9386,N_8954,N_8657);
xnor U9387 (N_9387,N_8696,N_8690);
xor U9388 (N_9388,N_8840,N_8937);
nor U9389 (N_9389,N_8476,N_8404);
nor U9390 (N_9390,N_8610,N_8575);
or U9391 (N_9391,N_8727,N_8982);
or U9392 (N_9392,N_8402,N_8415);
xor U9393 (N_9393,N_8642,N_8841);
or U9394 (N_9394,N_8898,N_8438);
nand U9395 (N_9395,N_8864,N_8584);
or U9396 (N_9396,N_8853,N_8953);
or U9397 (N_9397,N_8755,N_8616);
or U9398 (N_9398,N_8532,N_8940);
xor U9399 (N_9399,N_8957,N_8575);
and U9400 (N_9400,N_8925,N_8719);
nor U9401 (N_9401,N_8754,N_8487);
and U9402 (N_9402,N_8900,N_8908);
nor U9403 (N_9403,N_8470,N_8747);
nor U9404 (N_9404,N_8963,N_8496);
and U9405 (N_9405,N_8787,N_8702);
and U9406 (N_9406,N_8689,N_8772);
or U9407 (N_9407,N_8801,N_8623);
nand U9408 (N_9408,N_8869,N_8503);
nor U9409 (N_9409,N_8782,N_8970);
nor U9410 (N_9410,N_8424,N_8899);
xnor U9411 (N_9411,N_8953,N_8945);
xnor U9412 (N_9412,N_8918,N_8519);
or U9413 (N_9413,N_8412,N_8819);
and U9414 (N_9414,N_8594,N_8768);
or U9415 (N_9415,N_8704,N_8491);
and U9416 (N_9416,N_8658,N_8461);
or U9417 (N_9417,N_8654,N_8461);
nand U9418 (N_9418,N_8614,N_8404);
nand U9419 (N_9419,N_8714,N_8988);
nor U9420 (N_9420,N_8688,N_8410);
nand U9421 (N_9421,N_8573,N_8866);
or U9422 (N_9422,N_8855,N_8481);
nand U9423 (N_9423,N_8740,N_8616);
and U9424 (N_9424,N_8882,N_8626);
nor U9425 (N_9425,N_8620,N_8413);
xor U9426 (N_9426,N_8511,N_8423);
nor U9427 (N_9427,N_8560,N_8907);
and U9428 (N_9428,N_8833,N_8632);
or U9429 (N_9429,N_8701,N_8757);
nor U9430 (N_9430,N_8675,N_8600);
nand U9431 (N_9431,N_8709,N_8759);
and U9432 (N_9432,N_8563,N_8871);
xnor U9433 (N_9433,N_8620,N_8964);
nor U9434 (N_9434,N_8773,N_8601);
nand U9435 (N_9435,N_8423,N_8581);
nor U9436 (N_9436,N_8557,N_8606);
and U9437 (N_9437,N_8539,N_8522);
or U9438 (N_9438,N_8980,N_8788);
nor U9439 (N_9439,N_8501,N_8764);
nand U9440 (N_9440,N_8493,N_8601);
xnor U9441 (N_9441,N_8556,N_8636);
or U9442 (N_9442,N_8551,N_8650);
nor U9443 (N_9443,N_8400,N_8966);
nor U9444 (N_9444,N_8564,N_8926);
nor U9445 (N_9445,N_8523,N_8470);
xnor U9446 (N_9446,N_8772,N_8635);
and U9447 (N_9447,N_8494,N_8658);
nand U9448 (N_9448,N_8894,N_8773);
or U9449 (N_9449,N_8966,N_8893);
and U9450 (N_9450,N_8913,N_8774);
nor U9451 (N_9451,N_8896,N_8664);
nor U9452 (N_9452,N_8526,N_8897);
and U9453 (N_9453,N_8675,N_8661);
nand U9454 (N_9454,N_8858,N_8413);
xnor U9455 (N_9455,N_8673,N_8402);
xnor U9456 (N_9456,N_8432,N_8777);
or U9457 (N_9457,N_8518,N_8623);
or U9458 (N_9458,N_8449,N_8837);
and U9459 (N_9459,N_8900,N_8522);
nand U9460 (N_9460,N_8539,N_8826);
or U9461 (N_9461,N_8845,N_8810);
or U9462 (N_9462,N_8584,N_8983);
nor U9463 (N_9463,N_8768,N_8531);
and U9464 (N_9464,N_8758,N_8883);
nand U9465 (N_9465,N_8961,N_8654);
nand U9466 (N_9466,N_8519,N_8942);
and U9467 (N_9467,N_8780,N_8908);
and U9468 (N_9468,N_8733,N_8453);
nor U9469 (N_9469,N_8561,N_8906);
or U9470 (N_9470,N_8832,N_8837);
nor U9471 (N_9471,N_8953,N_8589);
nor U9472 (N_9472,N_8943,N_8436);
or U9473 (N_9473,N_8704,N_8413);
and U9474 (N_9474,N_8978,N_8585);
xor U9475 (N_9475,N_8758,N_8689);
and U9476 (N_9476,N_8661,N_8882);
xnor U9477 (N_9477,N_8748,N_8450);
or U9478 (N_9478,N_8565,N_8796);
nor U9479 (N_9479,N_8686,N_8479);
or U9480 (N_9480,N_8728,N_8850);
nand U9481 (N_9481,N_8422,N_8579);
nand U9482 (N_9482,N_8574,N_8553);
nand U9483 (N_9483,N_8632,N_8758);
nor U9484 (N_9484,N_8972,N_8916);
nand U9485 (N_9485,N_8798,N_8506);
and U9486 (N_9486,N_8695,N_8611);
or U9487 (N_9487,N_8575,N_8554);
xnor U9488 (N_9488,N_8744,N_8403);
xnor U9489 (N_9489,N_8492,N_8655);
xnor U9490 (N_9490,N_8935,N_8447);
or U9491 (N_9491,N_8471,N_8926);
nor U9492 (N_9492,N_8723,N_8697);
nand U9493 (N_9493,N_8824,N_8985);
xnor U9494 (N_9494,N_8972,N_8928);
nand U9495 (N_9495,N_8798,N_8556);
nand U9496 (N_9496,N_8920,N_8456);
nor U9497 (N_9497,N_8901,N_8929);
and U9498 (N_9498,N_8649,N_8858);
xnor U9499 (N_9499,N_8632,N_8418);
nand U9500 (N_9500,N_8506,N_8567);
xor U9501 (N_9501,N_8794,N_8407);
nand U9502 (N_9502,N_8687,N_8854);
xnor U9503 (N_9503,N_8862,N_8554);
nor U9504 (N_9504,N_8725,N_8993);
nor U9505 (N_9505,N_8612,N_8436);
nand U9506 (N_9506,N_8714,N_8412);
and U9507 (N_9507,N_8899,N_8466);
nor U9508 (N_9508,N_8943,N_8869);
nand U9509 (N_9509,N_8630,N_8948);
and U9510 (N_9510,N_8661,N_8724);
xnor U9511 (N_9511,N_8903,N_8437);
nand U9512 (N_9512,N_8619,N_8629);
xnor U9513 (N_9513,N_8794,N_8674);
xor U9514 (N_9514,N_8779,N_8405);
or U9515 (N_9515,N_8823,N_8677);
or U9516 (N_9516,N_8650,N_8581);
xnor U9517 (N_9517,N_8696,N_8705);
nor U9518 (N_9518,N_8947,N_8688);
and U9519 (N_9519,N_8444,N_8509);
nor U9520 (N_9520,N_8548,N_8496);
xor U9521 (N_9521,N_8851,N_8917);
and U9522 (N_9522,N_8982,N_8675);
and U9523 (N_9523,N_8860,N_8728);
nor U9524 (N_9524,N_8832,N_8834);
xor U9525 (N_9525,N_8558,N_8601);
nor U9526 (N_9526,N_8616,N_8548);
or U9527 (N_9527,N_8816,N_8757);
nand U9528 (N_9528,N_8463,N_8755);
nand U9529 (N_9529,N_8820,N_8578);
nor U9530 (N_9530,N_8462,N_8699);
or U9531 (N_9531,N_8729,N_8720);
nand U9532 (N_9532,N_8626,N_8571);
nand U9533 (N_9533,N_8896,N_8560);
or U9534 (N_9534,N_8973,N_8660);
xnor U9535 (N_9535,N_8596,N_8875);
xnor U9536 (N_9536,N_8757,N_8869);
or U9537 (N_9537,N_8548,N_8938);
nand U9538 (N_9538,N_8990,N_8931);
nor U9539 (N_9539,N_8736,N_8879);
xnor U9540 (N_9540,N_8909,N_8462);
and U9541 (N_9541,N_8619,N_8470);
xnor U9542 (N_9542,N_8486,N_8991);
nand U9543 (N_9543,N_8671,N_8576);
or U9544 (N_9544,N_8659,N_8965);
nor U9545 (N_9545,N_8631,N_8441);
nor U9546 (N_9546,N_8607,N_8635);
nor U9547 (N_9547,N_8908,N_8553);
xnor U9548 (N_9548,N_8439,N_8660);
nand U9549 (N_9549,N_8415,N_8592);
or U9550 (N_9550,N_8792,N_8920);
nand U9551 (N_9551,N_8863,N_8444);
or U9552 (N_9552,N_8503,N_8976);
and U9553 (N_9553,N_8405,N_8470);
nor U9554 (N_9554,N_8790,N_8943);
or U9555 (N_9555,N_8657,N_8424);
or U9556 (N_9556,N_8687,N_8819);
xor U9557 (N_9557,N_8745,N_8756);
nor U9558 (N_9558,N_8818,N_8893);
and U9559 (N_9559,N_8670,N_8958);
or U9560 (N_9560,N_8592,N_8787);
nand U9561 (N_9561,N_8429,N_8987);
xnor U9562 (N_9562,N_8561,N_8711);
nor U9563 (N_9563,N_8807,N_8820);
and U9564 (N_9564,N_8662,N_8836);
xor U9565 (N_9565,N_8805,N_8560);
nor U9566 (N_9566,N_8506,N_8645);
or U9567 (N_9567,N_8710,N_8861);
and U9568 (N_9568,N_8799,N_8905);
nand U9569 (N_9569,N_8461,N_8928);
and U9570 (N_9570,N_8620,N_8452);
and U9571 (N_9571,N_8951,N_8885);
and U9572 (N_9572,N_8520,N_8725);
nor U9573 (N_9573,N_8859,N_8989);
or U9574 (N_9574,N_8607,N_8974);
and U9575 (N_9575,N_8944,N_8713);
or U9576 (N_9576,N_8919,N_8552);
nor U9577 (N_9577,N_8780,N_8717);
or U9578 (N_9578,N_8840,N_8549);
nand U9579 (N_9579,N_8550,N_8910);
nand U9580 (N_9580,N_8507,N_8466);
xnor U9581 (N_9581,N_8659,N_8499);
nor U9582 (N_9582,N_8522,N_8547);
nor U9583 (N_9583,N_8860,N_8409);
nor U9584 (N_9584,N_8772,N_8836);
and U9585 (N_9585,N_8422,N_8835);
nor U9586 (N_9586,N_8914,N_8760);
nand U9587 (N_9587,N_8544,N_8624);
nor U9588 (N_9588,N_8493,N_8645);
or U9589 (N_9589,N_8489,N_8448);
xnor U9590 (N_9590,N_8777,N_8871);
and U9591 (N_9591,N_8849,N_8674);
nand U9592 (N_9592,N_8738,N_8712);
or U9593 (N_9593,N_8890,N_8801);
nor U9594 (N_9594,N_8991,N_8519);
and U9595 (N_9595,N_8726,N_8452);
or U9596 (N_9596,N_8761,N_8760);
xor U9597 (N_9597,N_8873,N_8943);
nand U9598 (N_9598,N_8951,N_8465);
or U9599 (N_9599,N_8923,N_8691);
xor U9600 (N_9600,N_9550,N_9409);
or U9601 (N_9601,N_9197,N_9446);
xor U9602 (N_9602,N_9144,N_9212);
nand U9603 (N_9603,N_9054,N_9165);
nor U9604 (N_9604,N_9045,N_9385);
nor U9605 (N_9605,N_9585,N_9583);
nand U9606 (N_9606,N_9528,N_9463);
xor U9607 (N_9607,N_9376,N_9452);
or U9608 (N_9608,N_9386,N_9420);
nand U9609 (N_9609,N_9450,N_9106);
nand U9610 (N_9610,N_9082,N_9189);
or U9611 (N_9611,N_9220,N_9505);
xor U9612 (N_9612,N_9545,N_9160);
and U9613 (N_9613,N_9531,N_9187);
and U9614 (N_9614,N_9564,N_9401);
xnor U9615 (N_9615,N_9374,N_9179);
nor U9616 (N_9616,N_9461,N_9108);
or U9617 (N_9617,N_9534,N_9544);
and U9618 (N_9618,N_9001,N_9367);
nor U9619 (N_9619,N_9053,N_9091);
nand U9620 (N_9620,N_9042,N_9566);
xnor U9621 (N_9621,N_9181,N_9047);
xor U9622 (N_9622,N_9083,N_9225);
nor U9623 (N_9623,N_9097,N_9396);
or U9624 (N_9624,N_9590,N_9475);
or U9625 (N_9625,N_9280,N_9019);
nand U9626 (N_9626,N_9041,N_9195);
nand U9627 (N_9627,N_9056,N_9427);
nand U9628 (N_9628,N_9482,N_9365);
nor U9629 (N_9629,N_9278,N_9388);
nand U9630 (N_9630,N_9138,N_9369);
xnor U9631 (N_9631,N_9006,N_9209);
and U9632 (N_9632,N_9524,N_9312);
nand U9633 (N_9633,N_9215,N_9440);
xnor U9634 (N_9634,N_9556,N_9236);
xnor U9635 (N_9635,N_9422,N_9473);
xnor U9636 (N_9636,N_9497,N_9368);
nor U9637 (N_9637,N_9502,N_9314);
nand U9638 (N_9638,N_9148,N_9582);
and U9639 (N_9639,N_9355,N_9559);
nand U9640 (N_9640,N_9008,N_9346);
nor U9641 (N_9641,N_9009,N_9309);
and U9642 (N_9642,N_9222,N_9481);
xnor U9643 (N_9643,N_9168,N_9134);
nand U9644 (N_9644,N_9494,N_9486);
nand U9645 (N_9645,N_9443,N_9162);
nand U9646 (N_9646,N_9244,N_9541);
nand U9647 (N_9647,N_9205,N_9594);
and U9648 (N_9648,N_9400,N_9533);
xnor U9649 (N_9649,N_9230,N_9086);
nor U9650 (N_9650,N_9542,N_9261);
and U9651 (N_9651,N_9335,N_9132);
nor U9652 (N_9652,N_9393,N_9003);
or U9653 (N_9653,N_9057,N_9119);
and U9654 (N_9654,N_9202,N_9254);
nor U9655 (N_9655,N_9589,N_9288);
nand U9656 (N_9656,N_9078,N_9276);
nand U9657 (N_9657,N_9338,N_9188);
xor U9658 (N_9658,N_9291,N_9477);
nand U9659 (N_9659,N_9273,N_9437);
and U9660 (N_9660,N_9044,N_9251);
nor U9661 (N_9661,N_9158,N_9429);
xor U9662 (N_9662,N_9077,N_9128);
or U9663 (N_9663,N_9577,N_9570);
or U9664 (N_9664,N_9432,N_9336);
and U9665 (N_9665,N_9064,N_9139);
nor U9666 (N_9666,N_9479,N_9522);
xor U9667 (N_9667,N_9467,N_9483);
nand U9668 (N_9668,N_9269,N_9571);
or U9669 (N_9669,N_9063,N_9038);
xor U9670 (N_9670,N_9048,N_9485);
and U9671 (N_9671,N_9184,N_9107);
xor U9672 (N_9672,N_9404,N_9306);
nand U9673 (N_9673,N_9166,N_9032);
nand U9674 (N_9674,N_9348,N_9296);
xor U9675 (N_9675,N_9352,N_9286);
nor U9676 (N_9676,N_9394,N_9024);
and U9677 (N_9677,N_9444,N_9208);
nand U9678 (N_9678,N_9358,N_9152);
nand U9679 (N_9679,N_9458,N_9334);
nand U9680 (N_9680,N_9087,N_9118);
or U9681 (N_9681,N_9238,N_9298);
or U9682 (N_9682,N_9176,N_9243);
or U9683 (N_9683,N_9249,N_9421);
nand U9684 (N_9684,N_9098,N_9115);
xnor U9685 (N_9685,N_9370,N_9340);
xnor U9686 (N_9686,N_9381,N_9584);
nor U9687 (N_9687,N_9242,N_9506);
nand U9688 (N_9688,N_9532,N_9092);
nor U9689 (N_9689,N_9468,N_9080);
xnor U9690 (N_9690,N_9426,N_9117);
nand U9691 (N_9691,N_9123,N_9052);
or U9692 (N_9692,N_9035,N_9178);
nand U9693 (N_9693,N_9297,N_9228);
and U9694 (N_9694,N_9445,N_9265);
and U9695 (N_9695,N_9096,N_9214);
and U9696 (N_9696,N_9331,N_9007);
or U9697 (N_9697,N_9313,N_9126);
nand U9698 (N_9698,N_9026,N_9263);
xor U9699 (N_9699,N_9449,N_9538);
nand U9700 (N_9700,N_9022,N_9407);
nand U9701 (N_9701,N_9345,N_9224);
or U9702 (N_9702,N_9329,N_9198);
and U9703 (N_9703,N_9402,N_9471);
and U9704 (N_9704,N_9282,N_9151);
nor U9705 (N_9705,N_9289,N_9216);
nor U9706 (N_9706,N_9241,N_9558);
nand U9707 (N_9707,N_9435,N_9543);
nand U9708 (N_9708,N_9448,N_9130);
nor U9709 (N_9709,N_9015,N_9527);
and U9710 (N_9710,N_9120,N_9223);
xor U9711 (N_9711,N_9303,N_9516);
xor U9712 (N_9712,N_9513,N_9030);
xor U9713 (N_9713,N_9510,N_9040);
or U9714 (N_9714,N_9462,N_9167);
nor U9715 (N_9715,N_9507,N_9598);
xor U9716 (N_9716,N_9354,N_9549);
xor U9717 (N_9717,N_9147,N_9302);
nand U9718 (N_9718,N_9438,N_9266);
nand U9719 (N_9719,N_9563,N_9163);
nor U9720 (N_9720,N_9501,N_9530);
xor U9721 (N_9721,N_9295,N_9509);
nand U9722 (N_9722,N_9460,N_9455);
or U9723 (N_9723,N_9259,N_9267);
xor U9724 (N_9724,N_9546,N_9536);
and U9725 (N_9725,N_9020,N_9182);
xnor U9726 (N_9726,N_9379,N_9177);
xor U9727 (N_9727,N_9363,N_9327);
or U9728 (N_9728,N_9256,N_9114);
or U9729 (N_9729,N_9308,N_9454);
nor U9730 (N_9730,N_9010,N_9116);
or U9731 (N_9731,N_9157,N_9560);
and U9732 (N_9732,N_9232,N_9525);
nand U9733 (N_9733,N_9068,N_9043);
and U9734 (N_9734,N_9090,N_9153);
xnor U9735 (N_9735,N_9362,N_9466);
nand U9736 (N_9736,N_9592,N_9557);
xnor U9737 (N_9737,N_9397,N_9074);
xnor U9738 (N_9738,N_9033,N_9279);
nor U9739 (N_9739,N_9561,N_9492);
xor U9740 (N_9740,N_9478,N_9299);
xnor U9741 (N_9741,N_9457,N_9172);
xnor U9742 (N_9742,N_9547,N_9217);
xor U9743 (N_9743,N_9226,N_9219);
or U9744 (N_9744,N_9360,N_9499);
xor U9745 (N_9745,N_9060,N_9412);
nand U9746 (N_9746,N_9073,N_9218);
nor U9747 (N_9747,N_9465,N_9099);
xor U9748 (N_9748,N_9002,N_9332);
nor U9749 (N_9749,N_9136,N_9121);
nor U9750 (N_9750,N_9490,N_9075);
nand U9751 (N_9751,N_9565,N_9428);
xnor U9752 (N_9752,N_9587,N_9529);
or U9753 (N_9753,N_9011,N_9129);
or U9754 (N_9754,N_9239,N_9287);
and U9755 (N_9755,N_9375,N_9210);
and U9756 (N_9756,N_9262,N_9055);
nand U9757 (N_9757,N_9413,N_9277);
or U9758 (N_9758,N_9089,N_9496);
nand U9759 (N_9759,N_9018,N_9599);
or U9760 (N_9760,N_9447,N_9310);
or U9761 (N_9761,N_9206,N_9240);
nor U9762 (N_9762,N_9004,N_9112);
nor U9763 (N_9763,N_9095,N_9211);
xor U9764 (N_9764,N_9135,N_9192);
xnor U9765 (N_9765,N_9343,N_9380);
nor U9766 (N_9766,N_9029,N_9233);
or U9767 (N_9767,N_9000,N_9349);
nand U9768 (N_9768,N_9316,N_9065);
or U9769 (N_9769,N_9037,N_9495);
nor U9770 (N_9770,N_9569,N_9359);
nor U9771 (N_9771,N_9100,N_9307);
nand U9772 (N_9772,N_9127,N_9164);
xor U9773 (N_9773,N_9392,N_9150);
xor U9774 (N_9774,N_9328,N_9416);
or U9775 (N_9775,N_9555,N_9377);
nand U9776 (N_9776,N_9341,N_9039);
and U9777 (N_9777,N_9325,N_9597);
nor U9778 (N_9778,N_9079,N_9229);
xnor U9779 (N_9779,N_9398,N_9200);
nor U9780 (N_9780,N_9133,N_9156);
nand U9781 (N_9781,N_9292,N_9433);
and U9782 (N_9782,N_9204,N_9567);
xnor U9783 (N_9783,N_9474,N_9050);
and U9784 (N_9784,N_9387,N_9517);
nand U9785 (N_9785,N_9441,N_9025);
xor U9786 (N_9786,N_9146,N_9105);
or U9787 (N_9787,N_9161,N_9183);
nor U9788 (N_9788,N_9285,N_9453);
xor U9789 (N_9789,N_9484,N_9072);
or U9790 (N_9790,N_9470,N_9154);
or U9791 (N_9791,N_9500,N_9175);
nor U9792 (N_9792,N_9250,N_9104);
or U9793 (N_9793,N_9382,N_9084);
nand U9794 (N_9794,N_9351,N_9201);
and U9795 (N_9795,N_9491,N_9081);
or U9796 (N_9796,N_9061,N_9318);
nor U9797 (N_9797,N_9058,N_9572);
xnor U9798 (N_9798,N_9012,N_9270);
nand U9799 (N_9799,N_9361,N_9399);
xor U9800 (N_9800,N_9034,N_9535);
xor U9801 (N_9801,N_9149,N_9070);
nand U9802 (N_9802,N_9311,N_9539);
xnor U9803 (N_9803,N_9319,N_9431);
xor U9804 (N_9804,N_9562,N_9304);
nor U9805 (N_9805,N_9456,N_9554);
and U9806 (N_9806,N_9272,N_9028);
or U9807 (N_9807,N_9122,N_9264);
and U9808 (N_9808,N_9321,N_9498);
nand U9809 (N_9809,N_9260,N_9476);
or U9810 (N_9810,N_9442,N_9066);
and U9811 (N_9811,N_9364,N_9537);
or U9812 (N_9812,N_9575,N_9185);
nand U9813 (N_9813,N_9186,N_9221);
xor U9814 (N_9814,N_9094,N_9005);
xnor U9815 (N_9815,N_9579,N_9451);
nor U9816 (N_9816,N_9586,N_9523);
nand U9817 (N_9817,N_9252,N_9323);
nand U9818 (N_9818,N_9111,N_9551);
xnor U9819 (N_9819,N_9417,N_9140);
xor U9820 (N_9820,N_9596,N_9353);
xnor U9821 (N_9821,N_9194,N_9142);
nor U9822 (N_9822,N_9419,N_9268);
xnor U9823 (N_9823,N_9344,N_9464);
nor U9824 (N_9824,N_9085,N_9322);
or U9825 (N_9825,N_9580,N_9076);
nor U9826 (N_9826,N_9493,N_9518);
nand U9827 (N_9827,N_9548,N_9014);
nand U9828 (N_9828,N_9190,N_9013);
or U9829 (N_9829,N_9257,N_9487);
xor U9830 (N_9830,N_9235,N_9406);
nor U9831 (N_9831,N_9021,N_9390);
nor U9832 (N_9832,N_9342,N_9300);
or U9833 (N_9833,N_9071,N_9339);
and U9834 (N_9834,N_9283,N_9036);
or U9835 (N_9835,N_9436,N_9103);
and U9836 (N_9836,N_9027,N_9519);
nand U9837 (N_9837,N_9389,N_9581);
or U9838 (N_9838,N_9290,N_9424);
nand U9839 (N_9839,N_9237,N_9301);
and U9840 (N_9840,N_9520,N_9434);
nand U9841 (N_9841,N_9016,N_9294);
or U9842 (N_9842,N_9143,N_9411);
nor U9843 (N_9843,N_9405,N_9526);
nor U9844 (N_9844,N_9227,N_9383);
xor U9845 (N_9845,N_9330,N_9488);
and U9846 (N_9846,N_9511,N_9350);
nand U9847 (N_9847,N_9508,N_9333);
xor U9848 (N_9848,N_9423,N_9540);
or U9849 (N_9849,N_9046,N_9356);
or U9850 (N_9850,N_9504,N_9088);
nor U9851 (N_9851,N_9109,N_9125);
nor U9852 (N_9852,N_9203,N_9315);
nor U9853 (N_9853,N_9503,N_9588);
or U9854 (N_9854,N_9595,N_9410);
xor U9855 (N_9855,N_9403,N_9320);
nand U9856 (N_9856,N_9378,N_9366);
xor U9857 (N_9857,N_9337,N_9049);
nor U9858 (N_9858,N_9408,N_9576);
or U9859 (N_9859,N_9199,N_9425);
and U9860 (N_9860,N_9207,N_9141);
xor U9861 (N_9861,N_9101,N_9512);
or U9862 (N_9862,N_9031,N_9110);
xnor U9863 (N_9863,N_9489,N_9271);
nand U9864 (N_9864,N_9062,N_9067);
and U9865 (N_9865,N_9255,N_9514);
xor U9866 (N_9866,N_9193,N_9069);
nand U9867 (N_9867,N_9317,N_9414);
or U9868 (N_9868,N_9059,N_9155);
nor U9869 (N_9869,N_9196,N_9124);
and U9870 (N_9870,N_9247,N_9113);
nor U9871 (N_9871,N_9591,N_9430);
xor U9872 (N_9872,N_9293,N_9371);
nor U9873 (N_9873,N_9180,N_9472);
or U9874 (N_9874,N_9159,N_9174);
or U9875 (N_9875,N_9418,N_9552);
or U9876 (N_9876,N_9170,N_9415);
nand U9877 (N_9877,N_9305,N_9573);
xnor U9878 (N_9878,N_9553,N_9017);
nand U9879 (N_9879,N_9372,N_9213);
nor U9880 (N_9880,N_9234,N_9137);
and U9881 (N_9881,N_9275,N_9023);
nor U9882 (N_9882,N_9191,N_9373);
xnor U9883 (N_9883,N_9568,N_9274);
nor U9884 (N_9884,N_9324,N_9347);
or U9885 (N_9885,N_9357,N_9593);
or U9886 (N_9886,N_9231,N_9326);
or U9887 (N_9887,N_9395,N_9102);
or U9888 (N_9888,N_9051,N_9169);
nor U9889 (N_9889,N_9131,N_9469);
or U9890 (N_9890,N_9384,N_9459);
or U9891 (N_9891,N_9574,N_9246);
or U9892 (N_9892,N_9284,N_9093);
xnor U9893 (N_9893,N_9391,N_9258);
nor U9894 (N_9894,N_9439,N_9515);
or U9895 (N_9895,N_9578,N_9145);
nand U9896 (N_9896,N_9245,N_9480);
xor U9897 (N_9897,N_9253,N_9521);
or U9898 (N_9898,N_9248,N_9171);
or U9899 (N_9899,N_9173,N_9281);
or U9900 (N_9900,N_9211,N_9110);
nand U9901 (N_9901,N_9264,N_9427);
nand U9902 (N_9902,N_9230,N_9554);
or U9903 (N_9903,N_9127,N_9093);
xor U9904 (N_9904,N_9544,N_9395);
or U9905 (N_9905,N_9549,N_9552);
xor U9906 (N_9906,N_9213,N_9006);
or U9907 (N_9907,N_9112,N_9314);
nand U9908 (N_9908,N_9229,N_9077);
xor U9909 (N_9909,N_9233,N_9243);
xor U9910 (N_9910,N_9488,N_9015);
xor U9911 (N_9911,N_9518,N_9206);
xor U9912 (N_9912,N_9086,N_9522);
xnor U9913 (N_9913,N_9554,N_9259);
nand U9914 (N_9914,N_9035,N_9491);
and U9915 (N_9915,N_9395,N_9068);
xor U9916 (N_9916,N_9095,N_9028);
or U9917 (N_9917,N_9050,N_9107);
or U9918 (N_9918,N_9096,N_9422);
and U9919 (N_9919,N_9273,N_9349);
nor U9920 (N_9920,N_9576,N_9445);
and U9921 (N_9921,N_9501,N_9455);
nor U9922 (N_9922,N_9580,N_9586);
and U9923 (N_9923,N_9309,N_9399);
xor U9924 (N_9924,N_9297,N_9498);
and U9925 (N_9925,N_9068,N_9430);
xor U9926 (N_9926,N_9325,N_9259);
xnor U9927 (N_9927,N_9273,N_9204);
nor U9928 (N_9928,N_9516,N_9383);
nor U9929 (N_9929,N_9328,N_9009);
or U9930 (N_9930,N_9489,N_9341);
nand U9931 (N_9931,N_9244,N_9530);
xor U9932 (N_9932,N_9012,N_9598);
nor U9933 (N_9933,N_9523,N_9441);
nor U9934 (N_9934,N_9539,N_9448);
nand U9935 (N_9935,N_9471,N_9317);
nor U9936 (N_9936,N_9327,N_9104);
xor U9937 (N_9937,N_9356,N_9283);
nand U9938 (N_9938,N_9566,N_9528);
nand U9939 (N_9939,N_9219,N_9040);
nor U9940 (N_9940,N_9472,N_9247);
or U9941 (N_9941,N_9355,N_9360);
nor U9942 (N_9942,N_9447,N_9507);
or U9943 (N_9943,N_9172,N_9482);
or U9944 (N_9944,N_9568,N_9558);
or U9945 (N_9945,N_9450,N_9351);
or U9946 (N_9946,N_9563,N_9382);
xnor U9947 (N_9947,N_9013,N_9054);
nor U9948 (N_9948,N_9249,N_9517);
xor U9949 (N_9949,N_9029,N_9427);
nor U9950 (N_9950,N_9191,N_9124);
and U9951 (N_9951,N_9366,N_9480);
and U9952 (N_9952,N_9067,N_9232);
nand U9953 (N_9953,N_9574,N_9298);
xor U9954 (N_9954,N_9302,N_9110);
xnor U9955 (N_9955,N_9326,N_9138);
nand U9956 (N_9956,N_9404,N_9279);
xnor U9957 (N_9957,N_9511,N_9056);
nor U9958 (N_9958,N_9270,N_9208);
xor U9959 (N_9959,N_9228,N_9416);
and U9960 (N_9960,N_9377,N_9236);
or U9961 (N_9961,N_9369,N_9354);
or U9962 (N_9962,N_9185,N_9399);
xor U9963 (N_9963,N_9463,N_9273);
xnor U9964 (N_9964,N_9428,N_9133);
or U9965 (N_9965,N_9282,N_9391);
nor U9966 (N_9966,N_9180,N_9450);
nor U9967 (N_9967,N_9081,N_9170);
and U9968 (N_9968,N_9366,N_9344);
and U9969 (N_9969,N_9091,N_9111);
nand U9970 (N_9970,N_9003,N_9574);
and U9971 (N_9971,N_9527,N_9165);
nand U9972 (N_9972,N_9594,N_9097);
nor U9973 (N_9973,N_9436,N_9592);
nand U9974 (N_9974,N_9356,N_9357);
and U9975 (N_9975,N_9314,N_9219);
and U9976 (N_9976,N_9378,N_9504);
xor U9977 (N_9977,N_9274,N_9358);
nand U9978 (N_9978,N_9276,N_9327);
and U9979 (N_9979,N_9202,N_9096);
nand U9980 (N_9980,N_9098,N_9336);
and U9981 (N_9981,N_9026,N_9553);
or U9982 (N_9982,N_9319,N_9099);
nand U9983 (N_9983,N_9417,N_9035);
or U9984 (N_9984,N_9047,N_9249);
xnor U9985 (N_9985,N_9294,N_9571);
nand U9986 (N_9986,N_9152,N_9544);
or U9987 (N_9987,N_9064,N_9387);
nand U9988 (N_9988,N_9380,N_9116);
or U9989 (N_9989,N_9482,N_9501);
nor U9990 (N_9990,N_9385,N_9186);
nand U9991 (N_9991,N_9067,N_9273);
or U9992 (N_9992,N_9436,N_9039);
nand U9993 (N_9993,N_9051,N_9221);
nand U9994 (N_9994,N_9009,N_9395);
nor U9995 (N_9995,N_9518,N_9029);
or U9996 (N_9996,N_9544,N_9417);
and U9997 (N_9997,N_9092,N_9510);
xnor U9998 (N_9998,N_9501,N_9100);
or U9999 (N_9999,N_9448,N_9200);
and U10000 (N_10000,N_9171,N_9139);
xor U10001 (N_10001,N_9125,N_9063);
xor U10002 (N_10002,N_9577,N_9554);
nand U10003 (N_10003,N_9002,N_9371);
or U10004 (N_10004,N_9197,N_9531);
and U10005 (N_10005,N_9502,N_9187);
nor U10006 (N_10006,N_9461,N_9135);
nand U10007 (N_10007,N_9449,N_9120);
and U10008 (N_10008,N_9552,N_9414);
nor U10009 (N_10009,N_9412,N_9094);
or U10010 (N_10010,N_9463,N_9154);
nand U10011 (N_10011,N_9190,N_9311);
and U10012 (N_10012,N_9473,N_9305);
and U10013 (N_10013,N_9420,N_9321);
nand U10014 (N_10014,N_9387,N_9288);
and U10015 (N_10015,N_9089,N_9202);
or U10016 (N_10016,N_9004,N_9288);
and U10017 (N_10017,N_9296,N_9065);
xnor U10018 (N_10018,N_9020,N_9562);
nor U10019 (N_10019,N_9042,N_9092);
nor U10020 (N_10020,N_9055,N_9426);
nor U10021 (N_10021,N_9512,N_9295);
or U10022 (N_10022,N_9330,N_9328);
and U10023 (N_10023,N_9131,N_9551);
or U10024 (N_10024,N_9497,N_9063);
and U10025 (N_10025,N_9162,N_9523);
and U10026 (N_10026,N_9087,N_9318);
or U10027 (N_10027,N_9052,N_9452);
and U10028 (N_10028,N_9556,N_9290);
or U10029 (N_10029,N_9228,N_9474);
nand U10030 (N_10030,N_9281,N_9204);
nand U10031 (N_10031,N_9308,N_9316);
or U10032 (N_10032,N_9317,N_9240);
nand U10033 (N_10033,N_9354,N_9143);
and U10034 (N_10034,N_9544,N_9170);
nand U10035 (N_10035,N_9089,N_9596);
and U10036 (N_10036,N_9588,N_9271);
nand U10037 (N_10037,N_9188,N_9089);
xor U10038 (N_10038,N_9003,N_9168);
nand U10039 (N_10039,N_9237,N_9315);
and U10040 (N_10040,N_9347,N_9559);
and U10041 (N_10041,N_9597,N_9315);
nor U10042 (N_10042,N_9394,N_9022);
nand U10043 (N_10043,N_9446,N_9058);
nand U10044 (N_10044,N_9337,N_9016);
xnor U10045 (N_10045,N_9373,N_9321);
nor U10046 (N_10046,N_9072,N_9273);
nor U10047 (N_10047,N_9479,N_9219);
and U10048 (N_10048,N_9594,N_9331);
nand U10049 (N_10049,N_9582,N_9264);
and U10050 (N_10050,N_9112,N_9072);
xnor U10051 (N_10051,N_9050,N_9156);
or U10052 (N_10052,N_9177,N_9323);
or U10053 (N_10053,N_9241,N_9335);
nor U10054 (N_10054,N_9526,N_9386);
and U10055 (N_10055,N_9568,N_9161);
nor U10056 (N_10056,N_9303,N_9100);
nor U10057 (N_10057,N_9219,N_9527);
nor U10058 (N_10058,N_9491,N_9435);
nor U10059 (N_10059,N_9185,N_9204);
and U10060 (N_10060,N_9557,N_9506);
or U10061 (N_10061,N_9435,N_9038);
or U10062 (N_10062,N_9401,N_9039);
and U10063 (N_10063,N_9458,N_9200);
or U10064 (N_10064,N_9105,N_9145);
nor U10065 (N_10065,N_9356,N_9471);
and U10066 (N_10066,N_9068,N_9108);
or U10067 (N_10067,N_9475,N_9464);
nor U10068 (N_10068,N_9367,N_9306);
or U10069 (N_10069,N_9236,N_9296);
nor U10070 (N_10070,N_9212,N_9477);
and U10071 (N_10071,N_9110,N_9332);
nor U10072 (N_10072,N_9256,N_9343);
nor U10073 (N_10073,N_9180,N_9379);
and U10074 (N_10074,N_9577,N_9247);
nor U10075 (N_10075,N_9078,N_9384);
nand U10076 (N_10076,N_9428,N_9373);
and U10077 (N_10077,N_9468,N_9052);
nand U10078 (N_10078,N_9052,N_9286);
nand U10079 (N_10079,N_9540,N_9495);
and U10080 (N_10080,N_9360,N_9309);
xnor U10081 (N_10081,N_9030,N_9194);
or U10082 (N_10082,N_9583,N_9216);
nand U10083 (N_10083,N_9005,N_9586);
xor U10084 (N_10084,N_9182,N_9174);
xor U10085 (N_10085,N_9484,N_9064);
and U10086 (N_10086,N_9014,N_9595);
and U10087 (N_10087,N_9349,N_9004);
nor U10088 (N_10088,N_9338,N_9077);
nand U10089 (N_10089,N_9306,N_9016);
nand U10090 (N_10090,N_9053,N_9378);
nand U10091 (N_10091,N_9522,N_9045);
or U10092 (N_10092,N_9108,N_9093);
xor U10093 (N_10093,N_9146,N_9019);
or U10094 (N_10094,N_9314,N_9225);
nand U10095 (N_10095,N_9571,N_9305);
or U10096 (N_10096,N_9304,N_9359);
or U10097 (N_10097,N_9387,N_9484);
nor U10098 (N_10098,N_9278,N_9503);
nand U10099 (N_10099,N_9230,N_9454);
nor U10100 (N_10100,N_9062,N_9113);
or U10101 (N_10101,N_9206,N_9461);
and U10102 (N_10102,N_9219,N_9595);
nand U10103 (N_10103,N_9402,N_9341);
xnor U10104 (N_10104,N_9444,N_9119);
nand U10105 (N_10105,N_9406,N_9018);
xor U10106 (N_10106,N_9066,N_9186);
nand U10107 (N_10107,N_9306,N_9112);
and U10108 (N_10108,N_9424,N_9354);
or U10109 (N_10109,N_9328,N_9570);
and U10110 (N_10110,N_9350,N_9473);
nand U10111 (N_10111,N_9342,N_9572);
or U10112 (N_10112,N_9473,N_9321);
xnor U10113 (N_10113,N_9489,N_9386);
or U10114 (N_10114,N_9350,N_9048);
nor U10115 (N_10115,N_9181,N_9462);
xor U10116 (N_10116,N_9113,N_9573);
or U10117 (N_10117,N_9585,N_9325);
nand U10118 (N_10118,N_9503,N_9053);
nor U10119 (N_10119,N_9495,N_9062);
nand U10120 (N_10120,N_9096,N_9054);
nand U10121 (N_10121,N_9595,N_9593);
nand U10122 (N_10122,N_9107,N_9450);
xnor U10123 (N_10123,N_9071,N_9243);
xnor U10124 (N_10124,N_9031,N_9255);
nor U10125 (N_10125,N_9519,N_9174);
nand U10126 (N_10126,N_9049,N_9479);
and U10127 (N_10127,N_9117,N_9302);
nor U10128 (N_10128,N_9081,N_9370);
or U10129 (N_10129,N_9123,N_9489);
or U10130 (N_10130,N_9015,N_9391);
or U10131 (N_10131,N_9399,N_9096);
nand U10132 (N_10132,N_9144,N_9376);
or U10133 (N_10133,N_9059,N_9015);
xnor U10134 (N_10134,N_9437,N_9400);
or U10135 (N_10135,N_9215,N_9091);
or U10136 (N_10136,N_9273,N_9597);
xnor U10137 (N_10137,N_9446,N_9077);
nor U10138 (N_10138,N_9406,N_9258);
or U10139 (N_10139,N_9165,N_9461);
nor U10140 (N_10140,N_9428,N_9349);
or U10141 (N_10141,N_9378,N_9282);
and U10142 (N_10142,N_9553,N_9572);
nor U10143 (N_10143,N_9370,N_9102);
and U10144 (N_10144,N_9562,N_9130);
xnor U10145 (N_10145,N_9489,N_9593);
xnor U10146 (N_10146,N_9500,N_9040);
nand U10147 (N_10147,N_9530,N_9151);
nor U10148 (N_10148,N_9342,N_9044);
and U10149 (N_10149,N_9035,N_9140);
nor U10150 (N_10150,N_9231,N_9297);
nand U10151 (N_10151,N_9293,N_9467);
and U10152 (N_10152,N_9359,N_9374);
and U10153 (N_10153,N_9067,N_9229);
or U10154 (N_10154,N_9148,N_9499);
nand U10155 (N_10155,N_9265,N_9492);
nand U10156 (N_10156,N_9082,N_9005);
nand U10157 (N_10157,N_9249,N_9219);
nand U10158 (N_10158,N_9106,N_9300);
xor U10159 (N_10159,N_9383,N_9316);
xor U10160 (N_10160,N_9036,N_9012);
nor U10161 (N_10161,N_9521,N_9535);
xnor U10162 (N_10162,N_9436,N_9244);
xor U10163 (N_10163,N_9098,N_9589);
and U10164 (N_10164,N_9222,N_9438);
or U10165 (N_10165,N_9538,N_9048);
nor U10166 (N_10166,N_9548,N_9357);
nor U10167 (N_10167,N_9571,N_9463);
and U10168 (N_10168,N_9197,N_9352);
xnor U10169 (N_10169,N_9514,N_9257);
xnor U10170 (N_10170,N_9242,N_9065);
nand U10171 (N_10171,N_9362,N_9581);
or U10172 (N_10172,N_9321,N_9148);
nand U10173 (N_10173,N_9183,N_9019);
xnor U10174 (N_10174,N_9557,N_9031);
and U10175 (N_10175,N_9413,N_9337);
xnor U10176 (N_10176,N_9069,N_9575);
or U10177 (N_10177,N_9155,N_9276);
nand U10178 (N_10178,N_9040,N_9515);
nor U10179 (N_10179,N_9209,N_9559);
xnor U10180 (N_10180,N_9103,N_9597);
nor U10181 (N_10181,N_9145,N_9480);
and U10182 (N_10182,N_9020,N_9232);
or U10183 (N_10183,N_9357,N_9318);
nor U10184 (N_10184,N_9416,N_9476);
nand U10185 (N_10185,N_9368,N_9538);
nor U10186 (N_10186,N_9053,N_9308);
or U10187 (N_10187,N_9575,N_9105);
or U10188 (N_10188,N_9117,N_9424);
and U10189 (N_10189,N_9261,N_9018);
and U10190 (N_10190,N_9454,N_9513);
and U10191 (N_10191,N_9272,N_9390);
xor U10192 (N_10192,N_9219,N_9351);
or U10193 (N_10193,N_9139,N_9571);
xor U10194 (N_10194,N_9022,N_9540);
nor U10195 (N_10195,N_9351,N_9076);
or U10196 (N_10196,N_9350,N_9297);
and U10197 (N_10197,N_9598,N_9085);
or U10198 (N_10198,N_9380,N_9595);
nand U10199 (N_10199,N_9205,N_9169);
nor U10200 (N_10200,N_10073,N_9817);
or U10201 (N_10201,N_10058,N_10151);
xor U10202 (N_10202,N_9748,N_10064);
and U10203 (N_10203,N_10159,N_9901);
or U10204 (N_10204,N_9984,N_10066);
nand U10205 (N_10205,N_9736,N_10124);
and U10206 (N_10206,N_10027,N_9742);
xnor U10207 (N_10207,N_9853,N_9770);
or U10208 (N_10208,N_10034,N_9902);
and U10209 (N_10209,N_9882,N_9785);
nand U10210 (N_10210,N_10088,N_10148);
or U10211 (N_10211,N_9603,N_9836);
nand U10212 (N_10212,N_9932,N_10031);
and U10213 (N_10213,N_10111,N_10154);
nor U10214 (N_10214,N_9686,N_9943);
xnor U10215 (N_10215,N_9680,N_10099);
xor U10216 (N_10216,N_9655,N_9828);
or U10217 (N_10217,N_9967,N_9780);
nand U10218 (N_10218,N_9638,N_9757);
or U10219 (N_10219,N_10108,N_10186);
nand U10220 (N_10220,N_10050,N_10030);
nor U10221 (N_10221,N_10060,N_9701);
and U10222 (N_10222,N_10097,N_9672);
nor U10223 (N_10223,N_9904,N_9760);
or U10224 (N_10224,N_10117,N_9809);
or U10225 (N_10225,N_9740,N_9936);
and U10226 (N_10226,N_10150,N_9894);
nor U10227 (N_10227,N_9703,N_9776);
nand U10228 (N_10228,N_10129,N_9887);
nor U10229 (N_10229,N_9648,N_10133);
nor U10230 (N_10230,N_10198,N_9766);
xor U10231 (N_10231,N_9966,N_10072);
nor U10232 (N_10232,N_9940,N_9965);
xnor U10233 (N_10233,N_9697,N_9633);
or U10234 (N_10234,N_9634,N_9691);
nand U10235 (N_10235,N_10195,N_10176);
nand U10236 (N_10236,N_9824,N_9820);
and U10237 (N_10237,N_9924,N_9617);
nand U10238 (N_10238,N_10011,N_10162);
nand U10239 (N_10239,N_10112,N_9641);
nor U10240 (N_10240,N_9751,N_10074);
xor U10241 (N_10241,N_9865,N_9654);
xnor U10242 (N_10242,N_10080,N_10093);
nor U10243 (N_10243,N_9790,N_9895);
nand U10244 (N_10244,N_9732,N_9679);
and U10245 (N_10245,N_9918,N_9771);
or U10246 (N_10246,N_9601,N_9645);
nand U10247 (N_10247,N_9713,N_9955);
nor U10248 (N_10248,N_9976,N_9723);
and U10249 (N_10249,N_9781,N_9805);
xnor U10250 (N_10250,N_9752,N_9621);
nand U10251 (N_10251,N_9840,N_9835);
nor U10252 (N_10252,N_10192,N_10067);
nand U10253 (N_10253,N_10103,N_9899);
and U10254 (N_10254,N_9667,N_9610);
nand U10255 (N_10255,N_9682,N_9992);
xnor U10256 (N_10256,N_10098,N_10063);
or U10257 (N_10257,N_9643,N_9636);
nand U10258 (N_10258,N_10052,N_9661);
nor U10259 (N_10259,N_9879,N_9741);
or U10260 (N_10260,N_10106,N_9812);
and U10261 (N_10261,N_9606,N_9874);
nor U10262 (N_10262,N_9928,N_9864);
nand U10263 (N_10263,N_9993,N_9685);
nand U10264 (N_10264,N_9816,N_9807);
nand U10265 (N_10265,N_9717,N_9880);
nand U10266 (N_10266,N_10191,N_9744);
xnor U10267 (N_10267,N_9861,N_9969);
nor U10268 (N_10268,N_9750,N_9960);
nand U10269 (N_10269,N_10168,N_9782);
nand U10270 (N_10270,N_9854,N_9825);
and U10271 (N_10271,N_9930,N_10130);
nand U10272 (N_10272,N_9962,N_9803);
xor U10273 (N_10273,N_9669,N_10042);
and U10274 (N_10274,N_9905,N_10116);
or U10275 (N_10275,N_9908,N_10002);
and U10276 (N_10276,N_9843,N_9659);
or U10277 (N_10277,N_9954,N_9614);
nand U10278 (N_10278,N_9725,N_10024);
nor U10279 (N_10279,N_10156,N_9794);
nor U10280 (N_10280,N_10166,N_9791);
or U10281 (N_10281,N_10086,N_9897);
and U10282 (N_10282,N_9871,N_10037);
xor U10283 (N_10283,N_9793,N_9778);
nor U10284 (N_10284,N_9755,N_9665);
and U10285 (N_10285,N_10183,N_10178);
nand U10286 (N_10286,N_10015,N_9656);
nor U10287 (N_10287,N_10045,N_10180);
or U10288 (N_10288,N_9640,N_9935);
nand U10289 (N_10289,N_9831,N_10101);
and U10290 (N_10290,N_9886,N_10081);
xor U10291 (N_10291,N_9762,N_9796);
nand U10292 (N_10292,N_10170,N_9964);
nor U10293 (N_10293,N_9818,N_10100);
and U10294 (N_10294,N_9844,N_10122);
or U10295 (N_10295,N_10118,N_9728);
nand U10296 (N_10296,N_9647,N_10033);
nand U10297 (N_10297,N_9709,N_10181);
nand U10298 (N_10298,N_9759,N_9738);
nor U10299 (N_10299,N_9852,N_9758);
nand U10300 (N_10300,N_9799,N_9891);
xnor U10301 (N_10301,N_9699,N_9716);
and U10302 (N_10302,N_9737,N_9810);
or U10303 (N_10303,N_9666,N_9658);
nand U10304 (N_10304,N_10075,N_9600);
xor U10305 (N_10305,N_10018,N_10059);
nand U10306 (N_10306,N_9869,N_10000);
nor U10307 (N_10307,N_10012,N_9784);
xor U10308 (N_10308,N_9849,N_9909);
nor U10309 (N_10309,N_10127,N_10190);
and U10310 (N_10310,N_9921,N_10092);
and U10311 (N_10311,N_10115,N_9959);
nand U10312 (N_10312,N_9772,N_9972);
xor U10313 (N_10313,N_10004,N_10175);
or U10314 (N_10314,N_9911,N_9689);
xnor U10315 (N_10315,N_9994,N_9963);
xnor U10316 (N_10316,N_10105,N_10141);
nand U10317 (N_10317,N_9779,N_10120);
or U10318 (N_10318,N_10007,N_10062);
xnor U10319 (N_10319,N_9729,N_9848);
nor U10320 (N_10320,N_9811,N_9743);
xor U10321 (N_10321,N_10149,N_10025);
or U10322 (N_10322,N_10121,N_9756);
and U10323 (N_10323,N_9980,N_9607);
or U10324 (N_10324,N_10140,N_10163);
nand U10325 (N_10325,N_9734,N_9800);
nand U10326 (N_10326,N_10006,N_9813);
and U10327 (N_10327,N_9674,N_9868);
nand U10328 (N_10328,N_10090,N_9917);
and U10329 (N_10329,N_10169,N_9925);
nor U10330 (N_10330,N_9653,N_10102);
and U10331 (N_10331,N_9683,N_9764);
and U10332 (N_10332,N_9730,N_9884);
and U10333 (N_10333,N_9620,N_9920);
and U10334 (N_10334,N_10039,N_10003);
nor U10335 (N_10335,N_9765,N_9704);
or U10336 (N_10336,N_9767,N_9892);
nand U10337 (N_10337,N_9945,N_10053);
nor U10338 (N_10338,N_9979,N_9989);
and U10339 (N_10339,N_9602,N_9727);
nand U10340 (N_10340,N_10114,N_10173);
nor U10341 (N_10341,N_10022,N_9931);
or U10342 (N_10342,N_9907,N_10085);
or U10343 (N_10343,N_10158,N_9624);
xor U10344 (N_10344,N_10132,N_9870);
xor U10345 (N_10345,N_9958,N_9613);
or U10346 (N_10346,N_9628,N_9690);
nand U10347 (N_10347,N_9650,N_9681);
or U10348 (N_10348,N_9783,N_10135);
or U10349 (N_10349,N_9754,N_9974);
or U10350 (N_10350,N_9625,N_9919);
nor U10351 (N_10351,N_10054,N_10019);
or U10352 (N_10352,N_9660,N_9923);
nor U10353 (N_10353,N_9986,N_9939);
xnor U10354 (N_10354,N_9858,N_9627);
xor U10355 (N_10355,N_10137,N_10083);
nand U10356 (N_10356,N_9823,N_9644);
xnor U10357 (N_10357,N_10185,N_9673);
nor U10358 (N_10358,N_10094,N_9684);
and U10359 (N_10359,N_9846,N_9941);
xor U10360 (N_10360,N_9998,N_10167);
or U10361 (N_10361,N_9705,N_9878);
nand U10362 (N_10362,N_9995,N_9949);
nand U10363 (N_10363,N_9970,N_9857);
and U10364 (N_10364,N_9706,N_9956);
and U10365 (N_10365,N_9707,N_9637);
nor U10366 (N_10366,N_10177,N_10189);
nand U10367 (N_10367,N_10143,N_9837);
nand U10368 (N_10368,N_10020,N_9719);
nor U10369 (N_10369,N_9692,N_9611);
nor U10370 (N_10370,N_10155,N_9626);
nor U10371 (N_10371,N_9842,N_9652);
nor U10372 (N_10372,N_9670,N_9657);
nand U10373 (N_10373,N_9838,N_9988);
nand U10374 (N_10374,N_9718,N_9881);
and U10375 (N_10375,N_10028,N_9639);
nand U10376 (N_10376,N_9850,N_9677);
xor U10377 (N_10377,N_10144,N_9826);
xor U10378 (N_10378,N_10036,N_9847);
nand U10379 (N_10379,N_9944,N_10160);
xnor U10380 (N_10380,N_9876,N_9642);
or U10381 (N_10381,N_10047,N_9971);
nand U10382 (N_10382,N_9663,N_10021);
nand U10383 (N_10383,N_9951,N_10146);
nor U10384 (N_10384,N_9795,N_9630);
nand U10385 (N_10385,N_9786,N_9604);
xor U10386 (N_10386,N_9910,N_10070);
nor U10387 (N_10387,N_10187,N_9866);
xor U10388 (N_10388,N_9753,N_9834);
nand U10389 (N_10389,N_9877,N_10139);
nand U10390 (N_10390,N_9773,N_9906);
nand U10391 (N_10391,N_10119,N_9792);
nand U10392 (N_10392,N_10076,N_9619);
nor U10393 (N_10393,N_9635,N_9933);
xor U10394 (N_10394,N_9618,N_9987);
or U10395 (N_10395,N_9903,N_9623);
nor U10396 (N_10396,N_9711,N_10145);
or U10397 (N_10397,N_9832,N_10082);
nand U10398 (N_10398,N_10048,N_9726);
nor U10399 (N_10399,N_10153,N_9739);
nand U10400 (N_10400,N_10184,N_9950);
xnor U10401 (N_10401,N_9676,N_9675);
nand U10402 (N_10402,N_9720,N_10147);
nand U10403 (N_10403,N_9859,N_9804);
and U10404 (N_10404,N_9815,N_10065);
and U10405 (N_10405,N_10126,N_9646);
and U10406 (N_10406,N_10091,N_9608);
xor U10407 (N_10407,N_9763,N_9863);
and U10408 (N_10408,N_10164,N_9622);
xor U10409 (N_10409,N_9733,N_9937);
or U10410 (N_10410,N_9615,N_9822);
and U10411 (N_10411,N_9916,N_9698);
and U10412 (N_10412,N_10049,N_9662);
nor U10413 (N_10413,N_9808,N_10079);
xor U10414 (N_10414,N_9983,N_9712);
nor U10415 (N_10415,N_9806,N_9774);
or U10416 (N_10416,N_10056,N_10078);
xor U10417 (N_10417,N_9724,N_9851);
or U10418 (N_10418,N_10138,N_10013);
or U10419 (N_10419,N_10016,N_9668);
nand U10420 (N_10420,N_10008,N_10068);
nor U10421 (N_10421,N_9845,N_10040);
xor U10422 (N_10422,N_9890,N_10161);
and U10423 (N_10423,N_10010,N_10032);
nand U10424 (N_10424,N_10179,N_9629);
xor U10425 (N_10425,N_9695,N_9860);
and U10426 (N_10426,N_9900,N_9814);
and U10427 (N_10427,N_10174,N_9888);
nand U10428 (N_10428,N_10199,N_9769);
nand U10429 (N_10429,N_10005,N_9873);
xor U10430 (N_10430,N_9746,N_10125);
and U10431 (N_10431,N_10171,N_9829);
nand U10432 (N_10432,N_9801,N_9787);
nand U10433 (N_10433,N_9721,N_9632);
nor U10434 (N_10434,N_9981,N_9889);
nand U10435 (N_10435,N_9839,N_9749);
or U10436 (N_10436,N_9953,N_9605);
xnor U10437 (N_10437,N_9671,N_9929);
xnor U10438 (N_10438,N_9922,N_9651);
xnor U10439 (N_10439,N_10128,N_10188);
nand U10440 (N_10440,N_10057,N_10104);
nand U10441 (N_10441,N_10142,N_9898);
nor U10442 (N_10442,N_10087,N_9687);
nor U10443 (N_10443,N_9990,N_9693);
and U10444 (N_10444,N_9997,N_9612);
xnor U10445 (N_10445,N_9688,N_10182);
and U10446 (N_10446,N_9999,N_9649);
nand U10447 (N_10447,N_9761,N_9631);
nand U10448 (N_10448,N_9872,N_10055);
or U10449 (N_10449,N_10051,N_10157);
nand U10450 (N_10450,N_9946,N_10113);
nor U10451 (N_10451,N_9927,N_10001);
xnor U10452 (N_10452,N_10009,N_9973);
nand U10453 (N_10453,N_10095,N_9788);
or U10454 (N_10454,N_9616,N_9883);
xor U10455 (N_10455,N_10014,N_9914);
xnor U10456 (N_10456,N_9714,N_9968);
or U10457 (N_10457,N_9802,N_9819);
nor U10458 (N_10458,N_9942,N_10026);
and U10459 (N_10459,N_9827,N_9694);
nor U10460 (N_10460,N_10165,N_9912);
xnor U10461 (N_10461,N_10044,N_10136);
or U10462 (N_10462,N_10077,N_10029);
or U10463 (N_10463,N_9867,N_9862);
nor U10464 (N_10464,N_9982,N_9841);
nand U10465 (N_10465,N_10134,N_9715);
xnor U10466 (N_10466,N_9833,N_9985);
xor U10467 (N_10467,N_10038,N_9856);
xnor U10468 (N_10468,N_9696,N_9977);
nor U10469 (N_10469,N_10152,N_10193);
nor U10470 (N_10470,N_9710,N_9747);
nor U10471 (N_10471,N_10017,N_10123);
xnor U10472 (N_10472,N_9789,N_9777);
nand U10473 (N_10473,N_9609,N_9797);
nor U10474 (N_10474,N_10131,N_10069);
xor U10475 (N_10475,N_10194,N_9975);
and U10476 (N_10476,N_9798,N_9893);
xor U10477 (N_10477,N_9938,N_10023);
nand U10478 (N_10478,N_10196,N_9821);
nand U10479 (N_10479,N_9952,N_9913);
xnor U10480 (N_10480,N_9957,N_10089);
xor U10481 (N_10481,N_9664,N_9947);
xor U10482 (N_10482,N_9896,N_10172);
and U10483 (N_10483,N_10084,N_9885);
xor U10484 (N_10484,N_10035,N_10107);
xnor U10485 (N_10485,N_10041,N_9830);
nor U10486 (N_10486,N_9722,N_9700);
nor U10487 (N_10487,N_9745,N_10197);
or U10488 (N_10488,N_10071,N_10061);
nor U10489 (N_10489,N_10109,N_9768);
xor U10490 (N_10490,N_9678,N_9735);
and U10491 (N_10491,N_9926,N_9991);
and U10492 (N_10492,N_10110,N_9915);
and U10493 (N_10493,N_9875,N_9948);
and U10494 (N_10494,N_9731,N_9775);
nand U10495 (N_10495,N_9708,N_9978);
nor U10496 (N_10496,N_10096,N_9996);
or U10497 (N_10497,N_10043,N_9855);
nand U10498 (N_10498,N_9961,N_10046);
nand U10499 (N_10499,N_9934,N_9702);
nor U10500 (N_10500,N_9932,N_9926);
nand U10501 (N_10501,N_9903,N_9899);
xnor U10502 (N_10502,N_9660,N_9630);
nand U10503 (N_10503,N_9659,N_9906);
xor U10504 (N_10504,N_9829,N_10004);
nor U10505 (N_10505,N_9744,N_9900);
nor U10506 (N_10506,N_9829,N_9621);
and U10507 (N_10507,N_9702,N_9973);
and U10508 (N_10508,N_9737,N_10015);
or U10509 (N_10509,N_10157,N_9911);
xor U10510 (N_10510,N_9911,N_10121);
nand U10511 (N_10511,N_9653,N_9983);
nor U10512 (N_10512,N_10110,N_10131);
xor U10513 (N_10513,N_9868,N_9821);
and U10514 (N_10514,N_10135,N_9718);
nand U10515 (N_10515,N_10008,N_10152);
or U10516 (N_10516,N_10104,N_10112);
and U10517 (N_10517,N_9743,N_9764);
nand U10518 (N_10518,N_9968,N_9604);
and U10519 (N_10519,N_9769,N_9931);
nor U10520 (N_10520,N_9995,N_9638);
or U10521 (N_10521,N_9765,N_10150);
xnor U10522 (N_10522,N_9898,N_10058);
and U10523 (N_10523,N_10143,N_10077);
and U10524 (N_10524,N_9836,N_9699);
and U10525 (N_10525,N_9783,N_10127);
nor U10526 (N_10526,N_9809,N_9816);
nor U10527 (N_10527,N_9707,N_10150);
or U10528 (N_10528,N_9770,N_10053);
and U10529 (N_10529,N_9932,N_9791);
nand U10530 (N_10530,N_10052,N_9965);
xor U10531 (N_10531,N_9805,N_10061);
xor U10532 (N_10532,N_9722,N_10021);
nand U10533 (N_10533,N_10195,N_10088);
nor U10534 (N_10534,N_10177,N_9936);
nor U10535 (N_10535,N_9852,N_9630);
nor U10536 (N_10536,N_9728,N_10113);
nand U10537 (N_10537,N_9696,N_10013);
or U10538 (N_10538,N_9799,N_10113);
or U10539 (N_10539,N_9751,N_9857);
and U10540 (N_10540,N_9620,N_9949);
nand U10541 (N_10541,N_9683,N_9755);
nor U10542 (N_10542,N_9994,N_10089);
nor U10543 (N_10543,N_10135,N_9922);
or U10544 (N_10544,N_10103,N_9605);
nor U10545 (N_10545,N_10067,N_9831);
or U10546 (N_10546,N_9896,N_10054);
and U10547 (N_10547,N_9813,N_9773);
xor U10548 (N_10548,N_9824,N_10033);
xor U10549 (N_10549,N_10193,N_9644);
nor U10550 (N_10550,N_9749,N_9931);
nand U10551 (N_10551,N_9764,N_9845);
nand U10552 (N_10552,N_10154,N_10030);
xor U10553 (N_10553,N_9663,N_9886);
and U10554 (N_10554,N_10156,N_9803);
and U10555 (N_10555,N_9765,N_10177);
or U10556 (N_10556,N_9985,N_10102);
nor U10557 (N_10557,N_10182,N_9809);
nand U10558 (N_10558,N_9920,N_9918);
nand U10559 (N_10559,N_10188,N_10103);
xor U10560 (N_10560,N_10031,N_9987);
and U10561 (N_10561,N_9840,N_9656);
or U10562 (N_10562,N_10154,N_10078);
or U10563 (N_10563,N_9614,N_10147);
nor U10564 (N_10564,N_9672,N_9949);
or U10565 (N_10565,N_10193,N_9640);
or U10566 (N_10566,N_10010,N_10177);
nand U10567 (N_10567,N_10069,N_10163);
xor U10568 (N_10568,N_10093,N_9784);
nand U10569 (N_10569,N_9807,N_10060);
nor U10570 (N_10570,N_9889,N_10091);
nor U10571 (N_10571,N_9935,N_10013);
xor U10572 (N_10572,N_9658,N_9637);
xor U10573 (N_10573,N_10123,N_10099);
or U10574 (N_10574,N_9920,N_9962);
xor U10575 (N_10575,N_10169,N_9929);
or U10576 (N_10576,N_10023,N_10175);
xor U10577 (N_10577,N_9754,N_9610);
nor U10578 (N_10578,N_10086,N_9880);
and U10579 (N_10579,N_10002,N_10071);
nand U10580 (N_10580,N_9991,N_9625);
nor U10581 (N_10581,N_9864,N_9810);
xor U10582 (N_10582,N_9876,N_10160);
nand U10583 (N_10583,N_9826,N_9814);
xor U10584 (N_10584,N_9801,N_9777);
or U10585 (N_10585,N_9791,N_9826);
xor U10586 (N_10586,N_9693,N_9944);
and U10587 (N_10587,N_10164,N_9821);
nand U10588 (N_10588,N_9992,N_9829);
nand U10589 (N_10589,N_9982,N_9754);
nor U10590 (N_10590,N_9723,N_9985);
nand U10591 (N_10591,N_9749,N_9760);
nor U10592 (N_10592,N_9666,N_9925);
nand U10593 (N_10593,N_9622,N_10188);
nor U10594 (N_10594,N_10133,N_10120);
xnor U10595 (N_10595,N_10193,N_9866);
nor U10596 (N_10596,N_10060,N_9973);
nor U10597 (N_10597,N_10196,N_10130);
xor U10598 (N_10598,N_9633,N_9682);
nand U10599 (N_10599,N_9964,N_9711);
and U10600 (N_10600,N_9735,N_10142);
and U10601 (N_10601,N_9975,N_9920);
or U10602 (N_10602,N_10153,N_10013);
nand U10603 (N_10603,N_9836,N_9814);
or U10604 (N_10604,N_9881,N_9703);
nand U10605 (N_10605,N_9807,N_10096);
or U10606 (N_10606,N_10023,N_10047);
and U10607 (N_10607,N_9600,N_10069);
and U10608 (N_10608,N_9894,N_9994);
or U10609 (N_10609,N_9912,N_10170);
or U10610 (N_10610,N_9733,N_9608);
nor U10611 (N_10611,N_9868,N_9632);
xnor U10612 (N_10612,N_10088,N_9729);
xor U10613 (N_10613,N_9882,N_9766);
nand U10614 (N_10614,N_9785,N_9754);
and U10615 (N_10615,N_10104,N_10156);
and U10616 (N_10616,N_9757,N_9707);
xnor U10617 (N_10617,N_9932,N_10109);
nand U10618 (N_10618,N_10126,N_9740);
and U10619 (N_10619,N_9757,N_10055);
and U10620 (N_10620,N_9733,N_9838);
nor U10621 (N_10621,N_9793,N_9742);
nor U10622 (N_10622,N_9804,N_9828);
and U10623 (N_10623,N_10081,N_9971);
nor U10624 (N_10624,N_9639,N_9601);
xor U10625 (N_10625,N_10066,N_9827);
nand U10626 (N_10626,N_9818,N_9677);
and U10627 (N_10627,N_9684,N_9708);
nand U10628 (N_10628,N_10153,N_9958);
or U10629 (N_10629,N_9767,N_9722);
or U10630 (N_10630,N_10085,N_10176);
xnor U10631 (N_10631,N_10060,N_10165);
nor U10632 (N_10632,N_9635,N_10139);
xor U10633 (N_10633,N_9974,N_10087);
nor U10634 (N_10634,N_9842,N_9882);
nor U10635 (N_10635,N_9749,N_10004);
xor U10636 (N_10636,N_9880,N_10168);
and U10637 (N_10637,N_9970,N_9816);
nor U10638 (N_10638,N_9618,N_9936);
nand U10639 (N_10639,N_9659,N_10143);
and U10640 (N_10640,N_9698,N_9684);
or U10641 (N_10641,N_9664,N_9658);
and U10642 (N_10642,N_10010,N_10041);
or U10643 (N_10643,N_9810,N_9923);
or U10644 (N_10644,N_9733,N_9602);
nor U10645 (N_10645,N_10156,N_9772);
nor U10646 (N_10646,N_9844,N_9854);
or U10647 (N_10647,N_9944,N_9870);
and U10648 (N_10648,N_10113,N_9761);
nor U10649 (N_10649,N_9872,N_9937);
xnor U10650 (N_10650,N_9759,N_9812);
xnor U10651 (N_10651,N_9805,N_9961);
nor U10652 (N_10652,N_9849,N_9605);
or U10653 (N_10653,N_9823,N_10174);
nand U10654 (N_10654,N_9792,N_9801);
or U10655 (N_10655,N_9778,N_9676);
nor U10656 (N_10656,N_10036,N_10063);
and U10657 (N_10657,N_9916,N_9963);
or U10658 (N_10658,N_9701,N_9680);
or U10659 (N_10659,N_10148,N_9669);
nor U10660 (N_10660,N_10020,N_9670);
and U10661 (N_10661,N_9634,N_9885);
nor U10662 (N_10662,N_9776,N_9745);
nand U10663 (N_10663,N_9826,N_9625);
nand U10664 (N_10664,N_9741,N_10030);
nand U10665 (N_10665,N_10172,N_9847);
nand U10666 (N_10666,N_9754,N_9987);
nand U10667 (N_10667,N_10156,N_9784);
and U10668 (N_10668,N_9661,N_9985);
nand U10669 (N_10669,N_9673,N_9868);
nand U10670 (N_10670,N_10118,N_9664);
nand U10671 (N_10671,N_9727,N_10005);
and U10672 (N_10672,N_9920,N_9949);
and U10673 (N_10673,N_10174,N_10126);
nor U10674 (N_10674,N_9949,N_9638);
nand U10675 (N_10675,N_10121,N_9766);
and U10676 (N_10676,N_10072,N_9630);
xnor U10677 (N_10677,N_9681,N_10142);
nand U10678 (N_10678,N_9664,N_9857);
and U10679 (N_10679,N_10104,N_10005);
xnor U10680 (N_10680,N_10028,N_9996);
and U10681 (N_10681,N_9644,N_9647);
and U10682 (N_10682,N_9846,N_10182);
and U10683 (N_10683,N_9688,N_9967);
nor U10684 (N_10684,N_9637,N_10076);
nand U10685 (N_10685,N_10050,N_10039);
xor U10686 (N_10686,N_9978,N_9806);
nor U10687 (N_10687,N_10140,N_9625);
or U10688 (N_10688,N_10032,N_9704);
or U10689 (N_10689,N_9674,N_9799);
or U10690 (N_10690,N_9883,N_9943);
or U10691 (N_10691,N_10031,N_9967);
nand U10692 (N_10692,N_9828,N_10127);
nor U10693 (N_10693,N_10068,N_10154);
nand U10694 (N_10694,N_9878,N_9994);
nand U10695 (N_10695,N_10168,N_10105);
nor U10696 (N_10696,N_9648,N_9616);
xor U10697 (N_10697,N_9734,N_10127);
nand U10698 (N_10698,N_10172,N_9977);
nor U10699 (N_10699,N_10049,N_10190);
or U10700 (N_10700,N_10168,N_9792);
nor U10701 (N_10701,N_9612,N_9956);
nor U10702 (N_10702,N_10178,N_9946);
nand U10703 (N_10703,N_9698,N_10034);
nand U10704 (N_10704,N_9683,N_9837);
and U10705 (N_10705,N_9894,N_10075);
nand U10706 (N_10706,N_9773,N_9775);
xnor U10707 (N_10707,N_10122,N_10027);
nor U10708 (N_10708,N_9718,N_9798);
or U10709 (N_10709,N_9959,N_9611);
xnor U10710 (N_10710,N_10191,N_10140);
and U10711 (N_10711,N_10154,N_9729);
nand U10712 (N_10712,N_10013,N_9843);
or U10713 (N_10713,N_9713,N_10144);
xnor U10714 (N_10714,N_9824,N_9807);
nor U10715 (N_10715,N_9858,N_9689);
and U10716 (N_10716,N_9865,N_10124);
or U10717 (N_10717,N_9698,N_9910);
and U10718 (N_10718,N_9831,N_9790);
nor U10719 (N_10719,N_10103,N_9613);
and U10720 (N_10720,N_9970,N_10017);
xnor U10721 (N_10721,N_9848,N_9605);
or U10722 (N_10722,N_10044,N_10079);
nand U10723 (N_10723,N_9910,N_9660);
xnor U10724 (N_10724,N_9909,N_10034);
or U10725 (N_10725,N_10082,N_10041);
and U10726 (N_10726,N_9639,N_9612);
and U10727 (N_10727,N_9704,N_9947);
nand U10728 (N_10728,N_10015,N_9918);
and U10729 (N_10729,N_9917,N_9786);
or U10730 (N_10730,N_9755,N_9886);
xor U10731 (N_10731,N_10011,N_9773);
nor U10732 (N_10732,N_9659,N_10021);
nor U10733 (N_10733,N_9949,N_9725);
xor U10734 (N_10734,N_9902,N_10132);
xor U10735 (N_10735,N_10102,N_9954);
or U10736 (N_10736,N_10030,N_9709);
or U10737 (N_10737,N_10033,N_9792);
and U10738 (N_10738,N_9969,N_9888);
nor U10739 (N_10739,N_9850,N_9882);
nor U10740 (N_10740,N_9839,N_9668);
nand U10741 (N_10741,N_10129,N_9718);
and U10742 (N_10742,N_9691,N_10086);
or U10743 (N_10743,N_10039,N_9880);
nor U10744 (N_10744,N_9848,N_9938);
or U10745 (N_10745,N_10080,N_9856);
or U10746 (N_10746,N_10033,N_9727);
or U10747 (N_10747,N_10085,N_9937);
or U10748 (N_10748,N_9843,N_10017);
nand U10749 (N_10749,N_9744,N_9876);
nand U10750 (N_10750,N_9941,N_10094);
or U10751 (N_10751,N_10168,N_9707);
nand U10752 (N_10752,N_9771,N_10035);
nor U10753 (N_10753,N_9665,N_9629);
and U10754 (N_10754,N_10175,N_10015);
or U10755 (N_10755,N_9686,N_9620);
and U10756 (N_10756,N_9640,N_9602);
xnor U10757 (N_10757,N_9813,N_9744);
xor U10758 (N_10758,N_9879,N_9697);
or U10759 (N_10759,N_9986,N_9705);
xnor U10760 (N_10760,N_9690,N_9890);
nor U10761 (N_10761,N_10151,N_10040);
and U10762 (N_10762,N_10179,N_9897);
xor U10763 (N_10763,N_9638,N_9809);
xnor U10764 (N_10764,N_9866,N_9757);
nor U10765 (N_10765,N_9903,N_9883);
nand U10766 (N_10766,N_9773,N_10022);
nor U10767 (N_10767,N_9980,N_10105);
xor U10768 (N_10768,N_10144,N_9954);
nor U10769 (N_10769,N_9690,N_9855);
xor U10770 (N_10770,N_9755,N_9815);
and U10771 (N_10771,N_9944,N_9804);
xor U10772 (N_10772,N_9716,N_9998);
xor U10773 (N_10773,N_10126,N_10127);
nand U10774 (N_10774,N_10169,N_10096);
nor U10775 (N_10775,N_10089,N_10113);
and U10776 (N_10776,N_9867,N_10051);
and U10777 (N_10777,N_10150,N_10112);
or U10778 (N_10778,N_9647,N_9798);
or U10779 (N_10779,N_9973,N_9780);
nand U10780 (N_10780,N_9898,N_9706);
nand U10781 (N_10781,N_9992,N_10115);
or U10782 (N_10782,N_9859,N_9631);
nor U10783 (N_10783,N_9886,N_9827);
and U10784 (N_10784,N_9845,N_9783);
or U10785 (N_10785,N_9851,N_9998);
nor U10786 (N_10786,N_10196,N_9676);
and U10787 (N_10787,N_10143,N_9963);
or U10788 (N_10788,N_10132,N_9605);
and U10789 (N_10789,N_9772,N_9712);
and U10790 (N_10790,N_9769,N_9921);
and U10791 (N_10791,N_10146,N_9861);
or U10792 (N_10792,N_10091,N_10140);
or U10793 (N_10793,N_9784,N_10150);
and U10794 (N_10794,N_10043,N_9888);
nand U10795 (N_10795,N_9821,N_9861);
nor U10796 (N_10796,N_9609,N_9675);
and U10797 (N_10797,N_10087,N_9880);
or U10798 (N_10798,N_9986,N_9742);
or U10799 (N_10799,N_9888,N_9652);
or U10800 (N_10800,N_10299,N_10415);
or U10801 (N_10801,N_10755,N_10399);
nand U10802 (N_10802,N_10343,N_10651);
or U10803 (N_10803,N_10376,N_10291);
nand U10804 (N_10804,N_10735,N_10567);
or U10805 (N_10805,N_10360,N_10468);
nor U10806 (N_10806,N_10236,N_10362);
nand U10807 (N_10807,N_10201,N_10326);
nand U10808 (N_10808,N_10336,N_10564);
or U10809 (N_10809,N_10633,N_10698);
nand U10810 (N_10810,N_10589,N_10391);
xor U10811 (N_10811,N_10680,N_10750);
nor U10812 (N_10812,N_10620,N_10444);
nand U10813 (N_10813,N_10699,N_10456);
nand U10814 (N_10814,N_10737,N_10548);
or U10815 (N_10815,N_10597,N_10264);
nand U10816 (N_10816,N_10792,N_10216);
xnor U10817 (N_10817,N_10208,N_10785);
or U10818 (N_10818,N_10358,N_10563);
or U10819 (N_10819,N_10733,N_10443);
nor U10820 (N_10820,N_10372,N_10587);
xor U10821 (N_10821,N_10780,N_10333);
nor U10822 (N_10822,N_10635,N_10740);
nor U10823 (N_10823,N_10572,N_10774);
nor U10824 (N_10824,N_10252,N_10647);
and U10825 (N_10825,N_10777,N_10380);
nor U10826 (N_10826,N_10576,N_10571);
or U10827 (N_10827,N_10294,N_10498);
nor U10828 (N_10828,N_10307,N_10310);
nand U10829 (N_10829,N_10256,N_10794);
and U10830 (N_10830,N_10344,N_10531);
nor U10831 (N_10831,N_10775,N_10405);
nand U10832 (N_10832,N_10428,N_10617);
nor U10833 (N_10833,N_10561,N_10400);
nand U10834 (N_10834,N_10345,N_10664);
nand U10835 (N_10835,N_10267,N_10791);
xnor U10836 (N_10836,N_10583,N_10782);
nor U10837 (N_10837,N_10215,N_10254);
nand U10838 (N_10838,N_10233,N_10555);
or U10839 (N_10839,N_10793,N_10662);
and U10840 (N_10840,N_10608,N_10560);
and U10841 (N_10841,N_10387,N_10761);
or U10842 (N_10842,N_10705,N_10243);
nand U10843 (N_10843,N_10667,N_10276);
nor U10844 (N_10844,N_10437,N_10363);
and U10845 (N_10845,N_10370,N_10205);
nor U10846 (N_10846,N_10258,N_10547);
nand U10847 (N_10847,N_10454,N_10776);
and U10848 (N_10848,N_10656,N_10230);
xnor U10849 (N_10849,N_10600,N_10432);
or U10850 (N_10850,N_10237,N_10287);
nor U10851 (N_10851,N_10674,N_10787);
nand U10852 (N_10852,N_10574,N_10210);
xor U10853 (N_10853,N_10732,N_10537);
nor U10854 (N_10854,N_10628,N_10729);
nor U10855 (N_10855,N_10371,N_10588);
nor U10856 (N_10856,N_10632,N_10591);
or U10857 (N_10857,N_10293,N_10753);
nand U10858 (N_10858,N_10337,N_10211);
nand U10859 (N_10859,N_10402,N_10631);
and U10860 (N_10860,N_10749,N_10408);
or U10861 (N_10861,N_10390,N_10356);
xor U10862 (N_10862,N_10594,N_10275);
nor U10863 (N_10863,N_10511,N_10320);
and U10864 (N_10864,N_10206,N_10709);
nand U10865 (N_10865,N_10687,N_10623);
nor U10866 (N_10866,N_10655,N_10477);
xnor U10867 (N_10867,N_10259,N_10523);
or U10868 (N_10868,N_10661,N_10673);
nor U10869 (N_10869,N_10719,N_10306);
nand U10870 (N_10870,N_10678,N_10551);
or U10871 (N_10871,N_10378,N_10644);
xnor U10872 (N_10872,N_10481,N_10229);
nor U10873 (N_10873,N_10706,N_10604);
xnor U10874 (N_10874,N_10424,N_10420);
nor U10875 (N_10875,N_10442,N_10247);
nand U10876 (N_10876,N_10579,N_10253);
or U10877 (N_10877,N_10557,N_10431);
or U10878 (N_10878,N_10495,N_10743);
xnor U10879 (N_10879,N_10240,N_10228);
nand U10880 (N_10880,N_10319,N_10701);
nor U10881 (N_10881,N_10332,N_10317);
nand U10882 (N_10882,N_10772,N_10781);
or U10883 (N_10883,N_10262,N_10734);
nand U10884 (N_10884,N_10438,N_10550);
nand U10885 (N_10885,N_10412,N_10500);
xor U10886 (N_10886,N_10342,N_10666);
nor U10887 (N_10887,N_10465,N_10538);
and U10888 (N_10888,N_10463,N_10469);
xnor U10889 (N_10889,N_10368,N_10377);
nor U10890 (N_10890,N_10725,N_10611);
nor U10891 (N_10891,N_10760,N_10383);
and U10892 (N_10892,N_10273,N_10249);
or U10893 (N_10893,N_10417,N_10328);
or U10894 (N_10894,N_10747,N_10475);
xnor U10895 (N_10895,N_10271,N_10354);
or U10896 (N_10896,N_10445,N_10744);
and U10897 (N_10897,N_10578,N_10621);
xnor U10898 (N_10898,N_10489,N_10395);
nand U10899 (N_10899,N_10278,N_10492);
xor U10900 (N_10900,N_10334,N_10462);
or U10901 (N_10901,N_10688,N_10488);
and U10902 (N_10902,N_10795,N_10321);
or U10903 (N_10903,N_10440,N_10450);
and U10904 (N_10904,N_10426,N_10448);
nor U10905 (N_10905,N_10464,N_10212);
or U10906 (N_10906,N_10718,N_10527);
xnor U10907 (N_10907,N_10250,N_10409);
nor U10908 (N_10908,N_10672,N_10392);
xnor U10909 (N_10909,N_10593,N_10452);
xnor U10910 (N_10910,N_10241,N_10364);
xnor U10911 (N_10911,N_10541,N_10502);
and U10912 (N_10912,N_10351,N_10446);
or U10913 (N_10913,N_10542,N_10601);
or U10914 (N_10914,N_10798,N_10365);
nand U10915 (N_10915,N_10742,N_10657);
nand U10916 (N_10916,N_10312,N_10219);
xor U10917 (N_10917,N_10757,N_10738);
nand U10918 (N_10918,N_10289,N_10285);
nor U10919 (N_10919,N_10353,N_10668);
or U10920 (N_10920,N_10418,N_10416);
or U10921 (N_10921,N_10730,N_10491);
nand U10922 (N_10922,N_10501,N_10677);
nor U10923 (N_10923,N_10634,N_10374);
and U10924 (N_10924,N_10435,N_10643);
nor U10925 (N_10925,N_10717,N_10348);
xnor U10926 (N_10926,N_10690,N_10494);
xor U10927 (N_10927,N_10231,N_10352);
nor U10928 (N_10928,N_10441,N_10302);
and U10929 (N_10929,N_10539,N_10327);
or U10930 (N_10930,N_10754,N_10727);
nand U10931 (N_10931,N_10707,N_10487);
nor U10932 (N_10932,N_10375,N_10367);
or U10933 (N_10933,N_10286,N_10692);
or U10934 (N_10934,N_10545,N_10640);
xnor U10935 (N_10935,N_10283,N_10427);
xor U10936 (N_10936,N_10313,N_10316);
and U10937 (N_10937,N_10473,N_10203);
xnor U10938 (N_10938,N_10603,N_10654);
nand U10939 (N_10939,N_10478,N_10663);
nor U10940 (N_10940,N_10304,N_10235);
and U10941 (N_10941,N_10771,N_10533);
or U10942 (N_10942,N_10386,N_10756);
and U10943 (N_10943,N_10619,N_10482);
nor U10944 (N_10944,N_10214,N_10516);
nor U10945 (N_10945,N_10669,N_10708);
or U10946 (N_10946,N_10769,N_10762);
xor U10947 (N_10947,N_10568,N_10300);
and U10948 (N_10948,N_10496,N_10357);
nand U10949 (N_10949,N_10484,N_10512);
xor U10950 (N_10950,N_10503,N_10288);
xnor U10951 (N_10951,N_10268,N_10222);
xor U10952 (N_10952,N_10765,N_10297);
xnor U10953 (N_10953,N_10586,N_10685);
xnor U10954 (N_10954,N_10245,N_10242);
nand U10955 (N_10955,N_10549,N_10410);
nor U10956 (N_10956,N_10540,N_10339);
xor U10957 (N_10957,N_10712,N_10460);
or U10958 (N_10958,N_10459,N_10279);
nand U10959 (N_10959,N_10748,N_10269);
or U10960 (N_10960,N_10789,N_10627);
nor U10961 (N_10961,N_10394,N_10493);
nand U10962 (N_10962,N_10556,N_10329);
nand U10963 (N_10963,N_10679,N_10255);
or U10964 (N_10964,N_10758,N_10778);
xor U10965 (N_10965,N_10315,N_10499);
nand U10966 (N_10966,N_10260,N_10366);
nand U10967 (N_10967,N_10615,N_10303);
or U10968 (N_10968,N_10385,N_10414);
xnor U10969 (N_10969,N_10263,N_10728);
nor U10970 (N_10970,N_10421,N_10277);
nand U10971 (N_10971,N_10266,N_10466);
nand U10972 (N_10972,N_10209,N_10703);
and U10973 (N_10973,N_10696,N_10483);
and U10974 (N_10974,N_10246,N_10507);
xnor U10975 (N_10975,N_10244,N_10553);
or U10976 (N_10976,N_10517,N_10425);
nor U10977 (N_10977,N_10722,N_10388);
and U10978 (N_10978,N_10340,N_10711);
or U10979 (N_10979,N_10751,N_10347);
nor U10980 (N_10980,N_10455,N_10311);
xnor U10981 (N_10981,N_10726,N_10514);
nand U10982 (N_10982,N_10763,N_10381);
or U10983 (N_10983,N_10474,N_10535);
and U10984 (N_10984,N_10693,N_10786);
nand U10985 (N_10985,N_10715,N_10683);
and U10986 (N_10986,N_10767,N_10797);
or U10987 (N_10987,N_10788,N_10565);
nor U10988 (N_10988,N_10575,N_10301);
xor U10989 (N_10989,N_10532,N_10359);
nand U10990 (N_10990,N_10626,N_10773);
nor U10991 (N_10991,N_10389,N_10265);
nand U10992 (N_10992,N_10704,N_10613);
or U10993 (N_10993,N_10436,N_10423);
or U10994 (N_10994,N_10239,N_10534);
nor U10995 (N_10995,N_10783,N_10659);
nand U10996 (N_10996,N_10447,N_10650);
and U10997 (N_10997,N_10606,N_10232);
or U10998 (N_10998,N_10544,N_10251);
nor U10999 (N_10999,N_10665,N_10379);
xor U11000 (N_11000,N_10518,N_10261);
and U11001 (N_11001,N_10689,N_10472);
xnor U11002 (N_11002,N_10309,N_10295);
and U11003 (N_11003,N_10433,N_10434);
or U11004 (N_11004,N_10612,N_10716);
xnor U11005 (N_11005,N_10403,N_10552);
nor U11006 (N_11006,N_10224,N_10622);
xor U11007 (N_11007,N_10768,N_10585);
xor U11008 (N_11008,N_10731,N_10697);
nor U11009 (N_11009,N_10530,N_10595);
and U11010 (N_11010,N_10373,N_10720);
xnor U11011 (N_11011,N_10207,N_10471);
or U11012 (N_11012,N_10524,N_10515);
and U11013 (N_11013,N_10526,N_10681);
nand U11014 (N_11014,N_10330,N_10598);
xor U11015 (N_11015,N_10398,N_10457);
and U11016 (N_11016,N_10658,N_10520);
and U11017 (N_11017,N_10636,N_10453);
nor U11018 (N_11018,N_10280,N_10325);
xnor U11019 (N_11019,N_10225,N_10355);
nor U11020 (N_11020,N_10582,N_10554);
or U11021 (N_11021,N_10397,N_10723);
nor U11022 (N_11022,N_10660,N_10648);
xor U11023 (N_11023,N_10779,N_10234);
and U11024 (N_11024,N_10314,N_10509);
xor U11025 (N_11025,N_10618,N_10404);
or U11026 (N_11026,N_10584,N_10684);
and U11027 (N_11027,N_10308,N_10671);
nand U11028 (N_11028,N_10270,N_10741);
and U11029 (N_11029,N_10573,N_10519);
nand U11030 (N_11030,N_10525,N_10486);
or U11031 (N_11031,N_10322,N_10318);
and U11032 (N_11032,N_10558,N_10653);
or U11033 (N_11033,N_10419,N_10467);
or U11034 (N_11034,N_10479,N_10625);
nand U11035 (N_11035,N_10570,N_10637);
nor U11036 (N_11036,N_10724,N_10770);
nand U11037 (N_11037,N_10562,N_10449);
or U11038 (N_11038,N_10305,N_10226);
or U11039 (N_11039,N_10642,N_10508);
or U11040 (N_11040,N_10700,N_10610);
nor U11041 (N_11041,N_10646,N_10335);
or U11042 (N_11042,N_10675,N_10248);
xor U11043 (N_11043,N_10670,N_10736);
nor U11044 (N_11044,N_10413,N_10590);
xnor U11045 (N_11045,N_10323,N_10213);
or U11046 (N_11046,N_10745,N_10349);
or U11047 (N_11047,N_10350,N_10504);
and U11048 (N_11048,N_10691,N_10202);
and U11049 (N_11049,N_10296,N_10506);
xnor U11050 (N_11050,N_10361,N_10580);
or U11051 (N_11051,N_10513,N_10624);
and U11052 (N_11052,N_10292,N_10505);
xor U11053 (N_11053,N_10766,N_10694);
or U11054 (N_11054,N_10566,N_10543);
nand U11055 (N_11055,N_10639,N_10714);
or U11056 (N_11056,N_10490,N_10223);
and U11057 (N_11057,N_10204,N_10238);
nor U11058 (N_11058,N_10217,N_10739);
nor U11059 (N_11059,N_10227,N_10616);
and U11060 (N_11060,N_10605,N_10759);
nand U11061 (N_11061,N_10396,N_10599);
nand U11062 (N_11062,N_10609,N_10695);
or U11063 (N_11063,N_10281,N_10422);
and U11064 (N_11064,N_10581,N_10470);
and U11065 (N_11065,N_10220,N_10369);
or U11066 (N_11066,N_10406,N_10393);
and U11067 (N_11067,N_10569,N_10401);
and U11068 (N_11068,N_10686,N_10614);
nor U11069 (N_11069,N_10461,N_10274);
nor U11070 (N_11070,N_10284,N_10592);
xnor U11071 (N_11071,N_10218,N_10607);
nor U11072 (N_11072,N_10682,N_10799);
xor U11073 (N_11073,N_10324,N_10577);
xor U11074 (N_11074,N_10338,N_10752);
xor U11075 (N_11075,N_10559,N_10796);
and U11076 (N_11076,N_10257,N_10764);
xnor U11077 (N_11077,N_10298,N_10536);
or U11078 (N_11078,N_10407,N_10630);
nand U11079 (N_11079,N_10522,N_10451);
or U11080 (N_11080,N_10430,N_10546);
nand U11081 (N_11081,N_10713,N_10341);
or U11082 (N_11082,N_10676,N_10746);
nor U11083 (N_11083,N_10476,N_10382);
nor U11084 (N_11084,N_10439,N_10497);
xor U11085 (N_11085,N_10645,N_10510);
and U11086 (N_11086,N_10629,N_10272);
and U11087 (N_11087,N_10528,N_10710);
xor U11088 (N_11088,N_10485,N_10596);
nand U11089 (N_11089,N_10641,N_10429);
or U11090 (N_11090,N_10529,N_10221);
xor U11091 (N_11091,N_10638,N_10784);
nor U11092 (N_11092,N_10649,N_10458);
and U11093 (N_11093,N_10282,N_10521);
or U11094 (N_11094,N_10480,N_10200);
or U11095 (N_11095,N_10652,N_10331);
nand U11096 (N_11096,N_10290,N_10411);
or U11097 (N_11097,N_10346,N_10602);
nor U11098 (N_11098,N_10790,N_10721);
and U11099 (N_11099,N_10702,N_10384);
or U11100 (N_11100,N_10676,N_10519);
nor U11101 (N_11101,N_10209,N_10264);
or U11102 (N_11102,N_10422,N_10261);
or U11103 (N_11103,N_10711,N_10759);
nand U11104 (N_11104,N_10761,N_10519);
nor U11105 (N_11105,N_10658,N_10717);
xor U11106 (N_11106,N_10750,N_10639);
nand U11107 (N_11107,N_10547,N_10659);
nand U11108 (N_11108,N_10281,N_10715);
nor U11109 (N_11109,N_10719,N_10520);
xnor U11110 (N_11110,N_10308,N_10608);
and U11111 (N_11111,N_10771,N_10404);
xnor U11112 (N_11112,N_10390,N_10549);
and U11113 (N_11113,N_10593,N_10446);
xnor U11114 (N_11114,N_10737,N_10726);
nor U11115 (N_11115,N_10395,N_10636);
and U11116 (N_11116,N_10457,N_10633);
and U11117 (N_11117,N_10291,N_10605);
nand U11118 (N_11118,N_10525,N_10626);
and U11119 (N_11119,N_10384,N_10265);
or U11120 (N_11120,N_10372,N_10428);
nor U11121 (N_11121,N_10310,N_10787);
or U11122 (N_11122,N_10313,N_10362);
nand U11123 (N_11123,N_10721,N_10307);
or U11124 (N_11124,N_10630,N_10293);
nor U11125 (N_11125,N_10785,N_10459);
xor U11126 (N_11126,N_10217,N_10484);
nor U11127 (N_11127,N_10388,N_10551);
or U11128 (N_11128,N_10728,N_10379);
nand U11129 (N_11129,N_10389,N_10762);
nand U11130 (N_11130,N_10232,N_10473);
nand U11131 (N_11131,N_10574,N_10347);
nand U11132 (N_11132,N_10714,N_10740);
nor U11133 (N_11133,N_10658,N_10316);
nor U11134 (N_11134,N_10289,N_10342);
nor U11135 (N_11135,N_10773,N_10425);
nand U11136 (N_11136,N_10426,N_10394);
nor U11137 (N_11137,N_10309,N_10651);
nand U11138 (N_11138,N_10525,N_10289);
or U11139 (N_11139,N_10752,N_10350);
xnor U11140 (N_11140,N_10564,N_10482);
or U11141 (N_11141,N_10567,N_10470);
nor U11142 (N_11142,N_10354,N_10700);
xor U11143 (N_11143,N_10376,N_10593);
xnor U11144 (N_11144,N_10716,N_10566);
nand U11145 (N_11145,N_10575,N_10555);
xor U11146 (N_11146,N_10403,N_10407);
nor U11147 (N_11147,N_10490,N_10690);
xnor U11148 (N_11148,N_10278,N_10532);
nor U11149 (N_11149,N_10347,N_10380);
nor U11150 (N_11150,N_10250,N_10593);
nand U11151 (N_11151,N_10611,N_10547);
or U11152 (N_11152,N_10298,N_10790);
nor U11153 (N_11153,N_10504,N_10553);
nand U11154 (N_11154,N_10227,N_10298);
and U11155 (N_11155,N_10645,N_10700);
or U11156 (N_11156,N_10326,N_10761);
and U11157 (N_11157,N_10470,N_10457);
and U11158 (N_11158,N_10329,N_10505);
nor U11159 (N_11159,N_10653,N_10741);
and U11160 (N_11160,N_10489,N_10400);
xnor U11161 (N_11161,N_10536,N_10379);
nand U11162 (N_11162,N_10248,N_10620);
nand U11163 (N_11163,N_10739,N_10310);
nor U11164 (N_11164,N_10263,N_10631);
xor U11165 (N_11165,N_10361,N_10316);
nor U11166 (N_11166,N_10310,N_10567);
xnor U11167 (N_11167,N_10500,N_10401);
xnor U11168 (N_11168,N_10274,N_10478);
xnor U11169 (N_11169,N_10366,N_10445);
xnor U11170 (N_11170,N_10325,N_10423);
nand U11171 (N_11171,N_10605,N_10698);
xnor U11172 (N_11172,N_10604,N_10765);
xor U11173 (N_11173,N_10419,N_10623);
xnor U11174 (N_11174,N_10386,N_10262);
xor U11175 (N_11175,N_10773,N_10771);
and U11176 (N_11176,N_10316,N_10552);
xor U11177 (N_11177,N_10317,N_10726);
and U11178 (N_11178,N_10597,N_10584);
xor U11179 (N_11179,N_10360,N_10763);
nand U11180 (N_11180,N_10424,N_10410);
nand U11181 (N_11181,N_10561,N_10353);
and U11182 (N_11182,N_10257,N_10427);
and U11183 (N_11183,N_10614,N_10491);
xor U11184 (N_11184,N_10210,N_10700);
nand U11185 (N_11185,N_10677,N_10333);
and U11186 (N_11186,N_10419,N_10528);
nor U11187 (N_11187,N_10556,N_10242);
nand U11188 (N_11188,N_10769,N_10719);
or U11189 (N_11189,N_10556,N_10435);
nor U11190 (N_11190,N_10512,N_10494);
and U11191 (N_11191,N_10618,N_10437);
nand U11192 (N_11192,N_10623,N_10227);
nor U11193 (N_11193,N_10453,N_10642);
nand U11194 (N_11194,N_10737,N_10699);
or U11195 (N_11195,N_10742,N_10389);
and U11196 (N_11196,N_10790,N_10524);
xor U11197 (N_11197,N_10769,N_10727);
and U11198 (N_11198,N_10234,N_10349);
nor U11199 (N_11199,N_10338,N_10794);
xor U11200 (N_11200,N_10622,N_10260);
or U11201 (N_11201,N_10585,N_10413);
and U11202 (N_11202,N_10522,N_10586);
nor U11203 (N_11203,N_10613,N_10369);
xnor U11204 (N_11204,N_10260,N_10581);
nor U11205 (N_11205,N_10550,N_10235);
and U11206 (N_11206,N_10508,N_10259);
nand U11207 (N_11207,N_10606,N_10601);
nand U11208 (N_11208,N_10306,N_10329);
and U11209 (N_11209,N_10504,N_10529);
xnor U11210 (N_11210,N_10272,N_10718);
or U11211 (N_11211,N_10351,N_10252);
nor U11212 (N_11212,N_10448,N_10376);
and U11213 (N_11213,N_10253,N_10220);
xor U11214 (N_11214,N_10709,N_10537);
nor U11215 (N_11215,N_10434,N_10409);
nand U11216 (N_11216,N_10433,N_10727);
nor U11217 (N_11217,N_10536,N_10402);
nand U11218 (N_11218,N_10428,N_10543);
nand U11219 (N_11219,N_10438,N_10359);
or U11220 (N_11220,N_10439,N_10619);
nand U11221 (N_11221,N_10771,N_10753);
nor U11222 (N_11222,N_10252,N_10733);
nor U11223 (N_11223,N_10369,N_10201);
and U11224 (N_11224,N_10269,N_10501);
and U11225 (N_11225,N_10377,N_10665);
xor U11226 (N_11226,N_10351,N_10278);
nand U11227 (N_11227,N_10635,N_10596);
nand U11228 (N_11228,N_10523,N_10622);
nor U11229 (N_11229,N_10738,N_10405);
nand U11230 (N_11230,N_10241,N_10460);
xor U11231 (N_11231,N_10374,N_10506);
xnor U11232 (N_11232,N_10262,N_10449);
or U11233 (N_11233,N_10609,N_10355);
nand U11234 (N_11234,N_10304,N_10514);
nor U11235 (N_11235,N_10372,N_10215);
nor U11236 (N_11236,N_10411,N_10384);
and U11237 (N_11237,N_10740,N_10559);
nor U11238 (N_11238,N_10561,N_10414);
and U11239 (N_11239,N_10640,N_10267);
nor U11240 (N_11240,N_10577,N_10383);
nor U11241 (N_11241,N_10655,N_10566);
or U11242 (N_11242,N_10434,N_10486);
nor U11243 (N_11243,N_10291,N_10311);
nand U11244 (N_11244,N_10420,N_10741);
nor U11245 (N_11245,N_10629,N_10348);
or U11246 (N_11246,N_10321,N_10703);
nor U11247 (N_11247,N_10200,N_10611);
or U11248 (N_11248,N_10469,N_10519);
and U11249 (N_11249,N_10210,N_10743);
xor U11250 (N_11250,N_10763,N_10258);
nor U11251 (N_11251,N_10229,N_10596);
nor U11252 (N_11252,N_10546,N_10661);
or U11253 (N_11253,N_10254,N_10269);
xor U11254 (N_11254,N_10752,N_10229);
and U11255 (N_11255,N_10456,N_10572);
nand U11256 (N_11256,N_10472,N_10362);
or U11257 (N_11257,N_10596,N_10763);
or U11258 (N_11258,N_10740,N_10773);
or U11259 (N_11259,N_10541,N_10483);
and U11260 (N_11260,N_10717,N_10703);
or U11261 (N_11261,N_10605,N_10341);
and U11262 (N_11262,N_10505,N_10303);
nand U11263 (N_11263,N_10783,N_10465);
xnor U11264 (N_11264,N_10758,N_10432);
nand U11265 (N_11265,N_10534,N_10465);
nor U11266 (N_11266,N_10660,N_10382);
or U11267 (N_11267,N_10542,N_10715);
and U11268 (N_11268,N_10734,N_10679);
or U11269 (N_11269,N_10444,N_10382);
and U11270 (N_11270,N_10757,N_10624);
nor U11271 (N_11271,N_10245,N_10623);
nor U11272 (N_11272,N_10537,N_10413);
nor U11273 (N_11273,N_10644,N_10289);
nor U11274 (N_11274,N_10670,N_10424);
nor U11275 (N_11275,N_10639,N_10350);
or U11276 (N_11276,N_10627,N_10505);
or U11277 (N_11277,N_10432,N_10507);
or U11278 (N_11278,N_10697,N_10525);
and U11279 (N_11279,N_10442,N_10235);
nor U11280 (N_11280,N_10346,N_10365);
and U11281 (N_11281,N_10352,N_10360);
xor U11282 (N_11282,N_10570,N_10413);
xor U11283 (N_11283,N_10637,N_10713);
xnor U11284 (N_11284,N_10403,N_10683);
nor U11285 (N_11285,N_10704,N_10608);
xor U11286 (N_11286,N_10550,N_10607);
and U11287 (N_11287,N_10459,N_10776);
nand U11288 (N_11288,N_10795,N_10322);
nor U11289 (N_11289,N_10512,N_10252);
nand U11290 (N_11290,N_10424,N_10573);
nor U11291 (N_11291,N_10363,N_10292);
nand U11292 (N_11292,N_10265,N_10411);
nand U11293 (N_11293,N_10262,N_10303);
or U11294 (N_11294,N_10256,N_10574);
or U11295 (N_11295,N_10624,N_10256);
nor U11296 (N_11296,N_10534,N_10691);
and U11297 (N_11297,N_10574,N_10255);
xor U11298 (N_11298,N_10253,N_10262);
xnor U11299 (N_11299,N_10750,N_10268);
and U11300 (N_11300,N_10268,N_10379);
or U11301 (N_11301,N_10625,N_10510);
nand U11302 (N_11302,N_10329,N_10799);
nand U11303 (N_11303,N_10328,N_10758);
and U11304 (N_11304,N_10792,N_10737);
or U11305 (N_11305,N_10484,N_10331);
xor U11306 (N_11306,N_10611,N_10204);
xor U11307 (N_11307,N_10628,N_10575);
and U11308 (N_11308,N_10344,N_10647);
and U11309 (N_11309,N_10553,N_10511);
and U11310 (N_11310,N_10764,N_10498);
nand U11311 (N_11311,N_10516,N_10251);
and U11312 (N_11312,N_10481,N_10271);
xnor U11313 (N_11313,N_10690,N_10739);
and U11314 (N_11314,N_10369,N_10690);
xor U11315 (N_11315,N_10556,N_10682);
xnor U11316 (N_11316,N_10310,N_10640);
xor U11317 (N_11317,N_10649,N_10658);
or U11318 (N_11318,N_10238,N_10362);
or U11319 (N_11319,N_10267,N_10242);
xor U11320 (N_11320,N_10251,N_10312);
xnor U11321 (N_11321,N_10656,N_10482);
nand U11322 (N_11322,N_10671,N_10213);
or U11323 (N_11323,N_10219,N_10351);
nor U11324 (N_11324,N_10265,N_10687);
nand U11325 (N_11325,N_10468,N_10223);
or U11326 (N_11326,N_10555,N_10420);
nor U11327 (N_11327,N_10630,N_10381);
and U11328 (N_11328,N_10616,N_10316);
or U11329 (N_11329,N_10755,N_10441);
nand U11330 (N_11330,N_10692,N_10467);
nor U11331 (N_11331,N_10701,N_10765);
nor U11332 (N_11332,N_10397,N_10550);
nor U11333 (N_11333,N_10417,N_10757);
or U11334 (N_11334,N_10246,N_10776);
nand U11335 (N_11335,N_10361,N_10742);
or U11336 (N_11336,N_10777,N_10453);
xor U11337 (N_11337,N_10707,N_10489);
xor U11338 (N_11338,N_10563,N_10522);
or U11339 (N_11339,N_10354,N_10404);
nor U11340 (N_11340,N_10351,N_10789);
and U11341 (N_11341,N_10478,N_10567);
nand U11342 (N_11342,N_10782,N_10229);
nand U11343 (N_11343,N_10508,N_10699);
nand U11344 (N_11344,N_10498,N_10676);
xnor U11345 (N_11345,N_10720,N_10453);
xor U11346 (N_11346,N_10482,N_10776);
or U11347 (N_11347,N_10326,N_10481);
nor U11348 (N_11348,N_10397,N_10400);
or U11349 (N_11349,N_10395,N_10377);
nor U11350 (N_11350,N_10344,N_10672);
xor U11351 (N_11351,N_10613,N_10742);
nand U11352 (N_11352,N_10478,N_10397);
and U11353 (N_11353,N_10428,N_10624);
nor U11354 (N_11354,N_10294,N_10464);
nor U11355 (N_11355,N_10370,N_10484);
xor U11356 (N_11356,N_10348,N_10402);
xnor U11357 (N_11357,N_10233,N_10713);
and U11358 (N_11358,N_10611,N_10219);
nand U11359 (N_11359,N_10683,N_10577);
xor U11360 (N_11360,N_10526,N_10366);
or U11361 (N_11361,N_10226,N_10567);
or U11362 (N_11362,N_10775,N_10441);
nor U11363 (N_11363,N_10666,N_10636);
xnor U11364 (N_11364,N_10663,N_10506);
nor U11365 (N_11365,N_10296,N_10470);
nor U11366 (N_11366,N_10654,N_10292);
and U11367 (N_11367,N_10245,N_10686);
nand U11368 (N_11368,N_10212,N_10727);
and U11369 (N_11369,N_10779,N_10493);
xnor U11370 (N_11370,N_10394,N_10408);
xor U11371 (N_11371,N_10446,N_10343);
xor U11372 (N_11372,N_10713,N_10474);
nand U11373 (N_11373,N_10233,N_10366);
or U11374 (N_11374,N_10431,N_10224);
and U11375 (N_11375,N_10483,N_10560);
or U11376 (N_11376,N_10476,N_10337);
xor U11377 (N_11377,N_10644,N_10640);
nand U11378 (N_11378,N_10233,N_10259);
and U11379 (N_11379,N_10365,N_10266);
nor U11380 (N_11380,N_10778,N_10353);
and U11381 (N_11381,N_10317,N_10770);
nor U11382 (N_11382,N_10700,N_10309);
xor U11383 (N_11383,N_10519,N_10790);
xor U11384 (N_11384,N_10700,N_10370);
nand U11385 (N_11385,N_10308,N_10774);
and U11386 (N_11386,N_10687,N_10756);
xor U11387 (N_11387,N_10628,N_10505);
nor U11388 (N_11388,N_10284,N_10217);
xor U11389 (N_11389,N_10741,N_10202);
or U11390 (N_11390,N_10515,N_10369);
xnor U11391 (N_11391,N_10581,N_10651);
nor U11392 (N_11392,N_10381,N_10246);
nand U11393 (N_11393,N_10464,N_10282);
xnor U11394 (N_11394,N_10471,N_10569);
xor U11395 (N_11395,N_10320,N_10593);
nand U11396 (N_11396,N_10463,N_10715);
and U11397 (N_11397,N_10750,N_10447);
nor U11398 (N_11398,N_10244,N_10726);
nor U11399 (N_11399,N_10391,N_10458);
or U11400 (N_11400,N_11162,N_11038);
and U11401 (N_11401,N_11090,N_11151);
and U11402 (N_11402,N_11023,N_10895);
xnor U11403 (N_11403,N_11129,N_11178);
or U11404 (N_11404,N_11369,N_11174);
nand U11405 (N_11405,N_11066,N_11045);
xor U11406 (N_11406,N_11095,N_11065);
nor U11407 (N_11407,N_10963,N_10846);
and U11408 (N_11408,N_11295,N_11398);
xor U11409 (N_11409,N_10847,N_11229);
and U11410 (N_11410,N_10925,N_10997);
and U11411 (N_11411,N_10862,N_11382);
or U11412 (N_11412,N_11137,N_11284);
nor U11413 (N_11413,N_11041,N_11141);
and U11414 (N_11414,N_11031,N_11275);
or U11415 (N_11415,N_11083,N_11088);
and U11416 (N_11416,N_11143,N_11245);
nor U11417 (N_11417,N_11225,N_10917);
xnor U11418 (N_11418,N_11384,N_10957);
nand U11419 (N_11419,N_10927,N_10878);
nor U11420 (N_11420,N_10866,N_10902);
and U11421 (N_11421,N_11020,N_11337);
xnor U11422 (N_11422,N_11061,N_11135);
xor U11423 (N_11423,N_11139,N_11293);
and U11424 (N_11424,N_10994,N_10800);
nor U11425 (N_11425,N_11358,N_11289);
and U11426 (N_11426,N_11113,N_11322);
or U11427 (N_11427,N_11222,N_11144);
and U11428 (N_11428,N_11030,N_10955);
and U11429 (N_11429,N_11013,N_11304);
nand U11430 (N_11430,N_10805,N_10836);
xor U11431 (N_11431,N_10833,N_10839);
or U11432 (N_11432,N_10907,N_11379);
nand U11433 (N_11433,N_11105,N_11334);
or U11434 (N_11434,N_11130,N_11299);
nor U11435 (N_11435,N_11303,N_11242);
nor U11436 (N_11436,N_11166,N_10851);
xor U11437 (N_11437,N_11138,N_11089);
nand U11438 (N_11438,N_11354,N_11274);
nor U11439 (N_11439,N_11282,N_10825);
nor U11440 (N_11440,N_11347,N_10841);
xor U11441 (N_11441,N_11048,N_11244);
xnor U11442 (N_11442,N_11216,N_11253);
nand U11443 (N_11443,N_11250,N_10937);
nand U11444 (N_11444,N_11291,N_11057);
or U11445 (N_11445,N_11211,N_11344);
xnor U11446 (N_11446,N_10983,N_11189);
xor U11447 (N_11447,N_11232,N_10988);
and U11448 (N_11448,N_11361,N_11165);
or U11449 (N_11449,N_11027,N_11318);
and U11450 (N_11450,N_11310,N_10956);
xnor U11451 (N_11451,N_11158,N_11373);
and U11452 (N_11452,N_11154,N_11161);
xor U11453 (N_11453,N_10934,N_10854);
or U11454 (N_11454,N_11306,N_11142);
nand U11455 (N_11455,N_11308,N_10940);
and U11456 (N_11456,N_11167,N_10831);
or U11457 (N_11457,N_10807,N_10962);
and U11458 (N_11458,N_11380,N_10813);
or U11459 (N_11459,N_11018,N_11012);
nor U11460 (N_11460,N_11281,N_11336);
nand U11461 (N_11461,N_11180,N_11351);
nand U11462 (N_11462,N_10979,N_11094);
nor U11463 (N_11463,N_11283,N_11163);
xnor U11464 (N_11464,N_10899,N_11022);
xor U11465 (N_11465,N_10816,N_11233);
and U11466 (N_11466,N_11194,N_11395);
xor U11467 (N_11467,N_11014,N_10929);
and U11468 (N_11468,N_11346,N_11079);
or U11469 (N_11469,N_11203,N_11058);
or U11470 (N_11470,N_11140,N_11333);
xnor U11471 (N_11471,N_11292,N_11285);
nor U11472 (N_11472,N_10920,N_10951);
or U11473 (N_11473,N_11146,N_11365);
and U11474 (N_11474,N_11301,N_11133);
and U11475 (N_11475,N_10844,N_10860);
xor U11476 (N_11476,N_11099,N_11348);
or U11477 (N_11477,N_11234,N_10885);
xnor U11478 (N_11478,N_10823,N_11390);
and U11479 (N_11479,N_11070,N_10973);
and U11480 (N_11480,N_11238,N_11312);
nor U11481 (N_11481,N_10911,N_11043);
nand U11482 (N_11482,N_11076,N_11069);
and U11483 (N_11483,N_11157,N_11325);
nor U11484 (N_11484,N_10879,N_10818);
or U11485 (N_11485,N_10887,N_11159);
nor U11486 (N_11486,N_10991,N_10923);
nor U11487 (N_11487,N_11145,N_11227);
or U11488 (N_11488,N_11075,N_11134);
or U11489 (N_11489,N_10830,N_11214);
xor U11490 (N_11490,N_10874,N_10810);
or U11491 (N_11491,N_10928,N_11341);
nor U11492 (N_11492,N_10910,N_11372);
nor U11493 (N_11493,N_11276,N_10974);
nor U11494 (N_11494,N_11032,N_10982);
nand U11495 (N_11495,N_10950,N_11055);
xor U11496 (N_11496,N_11188,N_11191);
nand U11497 (N_11497,N_11237,N_10814);
nand U11498 (N_11498,N_10972,N_11202);
nand U11499 (N_11499,N_10873,N_11086);
nand U11500 (N_11500,N_11085,N_11307);
or U11501 (N_11501,N_11082,N_11148);
nor U11502 (N_11502,N_11210,N_11241);
xnor U11503 (N_11503,N_11262,N_11338);
or U11504 (N_11504,N_11097,N_10971);
nor U11505 (N_11505,N_11224,N_11386);
or U11506 (N_11506,N_10900,N_10832);
or U11507 (N_11507,N_11215,N_11220);
xnor U11508 (N_11508,N_10890,N_10896);
and U11509 (N_11509,N_10998,N_10990);
nand U11510 (N_11510,N_10959,N_11316);
xor U11511 (N_11511,N_11399,N_10954);
and U11512 (N_11512,N_11153,N_11204);
and U11513 (N_11513,N_10898,N_10943);
xnor U11514 (N_11514,N_11201,N_10945);
or U11515 (N_11515,N_10931,N_10984);
nand U11516 (N_11516,N_10933,N_11231);
nand U11517 (N_11517,N_11251,N_11363);
nor U11518 (N_11518,N_11272,N_11117);
and U11519 (N_11519,N_11219,N_10861);
and U11520 (N_11520,N_11327,N_11235);
and U11521 (N_11521,N_10953,N_10965);
nor U11522 (N_11522,N_10952,N_11186);
or U11523 (N_11523,N_11212,N_11217);
nor U11524 (N_11524,N_10901,N_11156);
or U11525 (N_11525,N_11255,N_10882);
xor U11526 (N_11526,N_11261,N_11335);
nand U11527 (N_11527,N_11265,N_11100);
nor U11528 (N_11528,N_10888,N_11181);
nor U11529 (N_11529,N_10904,N_11039);
xor U11530 (N_11530,N_11190,N_11248);
nor U11531 (N_11531,N_11332,N_11008);
nand U11532 (N_11532,N_10801,N_10970);
nor U11533 (N_11533,N_11317,N_11277);
or U11534 (N_11534,N_11176,N_11199);
or U11535 (N_11535,N_11073,N_10803);
and U11536 (N_11536,N_11247,N_11315);
and U11537 (N_11537,N_10909,N_11209);
or U11538 (N_11538,N_10976,N_10916);
xnor U11539 (N_11539,N_11172,N_11192);
or U11540 (N_11540,N_11208,N_11102);
nor U11541 (N_11541,N_10822,N_10867);
and U11542 (N_11542,N_11371,N_11226);
and U11543 (N_11543,N_11213,N_10876);
and U11544 (N_11544,N_11391,N_11280);
xor U11545 (N_11545,N_11260,N_11147);
or U11546 (N_11546,N_10821,N_11021);
xor U11547 (N_11547,N_10829,N_10989);
or U11548 (N_11548,N_11087,N_10880);
or U11549 (N_11549,N_10961,N_10996);
nand U11550 (N_11550,N_10817,N_11125);
nand U11551 (N_11551,N_11356,N_11254);
and U11552 (N_11552,N_11297,N_11056);
nor U11553 (N_11553,N_10960,N_11124);
nand U11554 (N_11554,N_11360,N_11313);
nand U11555 (N_11555,N_11200,N_11004);
nand U11556 (N_11556,N_11271,N_11046);
xor U11557 (N_11557,N_11118,N_10838);
nor U11558 (N_11558,N_11394,N_11119);
xnor U11559 (N_11559,N_11331,N_11177);
xor U11560 (N_11560,N_10906,N_11108);
and U11561 (N_11561,N_11328,N_10981);
or U11562 (N_11562,N_11071,N_11196);
nor U11563 (N_11563,N_10824,N_11175);
and U11564 (N_11564,N_11267,N_10946);
and U11565 (N_11565,N_11121,N_11207);
xnor U11566 (N_11566,N_11050,N_11221);
and U11567 (N_11567,N_11128,N_10987);
or U11568 (N_11568,N_11064,N_11040);
nand U11569 (N_11569,N_11169,N_11270);
or U11570 (N_11570,N_11168,N_11003);
or U11571 (N_11571,N_11387,N_11001);
or U11572 (N_11572,N_11218,N_10889);
or U11573 (N_11573,N_11049,N_11002);
and U11574 (N_11574,N_11298,N_11246);
nor U11575 (N_11575,N_10992,N_10886);
or U11576 (N_11576,N_11296,N_11007);
and U11577 (N_11577,N_11042,N_11383);
xnor U11578 (N_11578,N_10850,N_10969);
or U11579 (N_11579,N_11198,N_11311);
nand U11580 (N_11580,N_11106,N_10881);
nor U11581 (N_11581,N_10967,N_11268);
nor U11582 (N_11582,N_10877,N_10912);
nand U11583 (N_11583,N_10827,N_11375);
nor U11584 (N_11584,N_10897,N_11170);
and U11585 (N_11585,N_11355,N_11112);
xor U11586 (N_11586,N_11343,N_11396);
nor U11587 (N_11587,N_11364,N_10935);
nand U11588 (N_11588,N_10930,N_11252);
or U11589 (N_11589,N_11026,N_11350);
nand U11590 (N_11590,N_11397,N_11366);
nand U11591 (N_11591,N_11388,N_11006);
nand U11592 (N_11592,N_11126,N_11015);
or U11593 (N_11593,N_11155,N_11193);
nor U11594 (N_11594,N_11152,N_10894);
nor U11595 (N_11595,N_10809,N_11179);
xor U11596 (N_11596,N_11047,N_10840);
or U11597 (N_11597,N_10905,N_10826);
xor U11598 (N_11598,N_11074,N_10871);
xnor U11599 (N_11599,N_11005,N_10819);
nand U11600 (N_11600,N_10865,N_11319);
xnor U11601 (N_11601,N_11036,N_11288);
nor U11602 (N_11602,N_11345,N_11326);
nand U11603 (N_11603,N_11302,N_11342);
and U11604 (N_11604,N_11025,N_11017);
nor U11605 (N_11605,N_10914,N_11269);
and U11606 (N_11606,N_11357,N_10995);
nor U11607 (N_11607,N_11362,N_10918);
nor U11608 (N_11608,N_10903,N_10913);
or U11609 (N_11609,N_10932,N_10986);
xor U11610 (N_11610,N_10837,N_11324);
nand U11611 (N_11611,N_10941,N_11349);
and U11612 (N_11612,N_10884,N_10947);
nor U11613 (N_11613,N_10863,N_11340);
or U11614 (N_11614,N_10948,N_11160);
nor U11615 (N_11615,N_11273,N_11309);
or U11616 (N_11616,N_11377,N_11393);
nand U11617 (N_11617,N_10980,N_10834);
or U11618 (N_11618,N_11329,N_11368);
nand U11619 (N_11619,N_11081,N_10820);
or U11620 (N_11620,N_11072,N_11239);
or U11621 (N_11621,N_11330,N_11367);
and U11622 (N_11622,N_11389,N_10845);
and U11623 (N_11623,N_11195,N_10869);
or U11624 (N_11624,N_10908,N_11374);
nor U11625 (N_11625,N_11037,N_11131);
or U11626 (N_11626,N_10958,N_11287);
nand U11627 (N_11627,N_10857,N_11392);
xnor U11628 (N_11628,N_10891,N_10842);
nor U11629 (N_11629,N_11183,N_11098);
or U11630 (N_11630,N_10843,N_11378);
or U11631 (N_11631,N_10922,N_10855);
xor U11632 (N_11632,N_11294,N_11062);
nor U11633 (N_11633,N_10864,N_11197);
and U11634 (N_11634,N_11104,N_11290);
xor U11635 (N_11635,N_10924,N_11060);
or U11636 (N_11636,N_11053,N_10938);
nand U11637 (N_11637,N_11096,N_11059);
or U11638 (N_11638,N_11256,N_10942);
nor U11639 (N_11639,N_10926,N_11051);
xor U11640 (N_11640,N_10872,N_11263);
and U11641 (N_11641,N_11249,N_10811);
xnor U11642 (N_11642,N_11205,N_11034);
nor U11643 (N_11643,N_10828,N_11052);
xor U11644 (N_11644,N_10892,N_11063);
nor U11645 (N_11645,N_11114,N_10875);
xor U11646 (N_11646,N_11000,N_11080);
nor U11647 (N_11647,N_11381,N_11352);
or U11648 (N_11648,N_10978,N_11019);
xor U11649 (N_11649,N_11092,N_11077);
or U11650 (N_11650,N_11068,N_11016);
xor U11651 (N_11651,N_11320,N_11044);
nand U11652 (N_11652,N_10848,N_10893);
xnor U11653 (N_11653,N_11084,N_11240);
xnor U11654 (N_11654,N_11136,N_11321);
nor U11655 (N_11655,N_11028,N_10919);
or U11656 (N_11656,N_10856,N_10921);
and U11657 (N_11657,N_11385,N_11228);
xor U11658 (N_11658,N_11109,N_10949);
or U11659 (N_11659,N_10804,N_10999);
or U11660 (N_11660,N_10849,N_11243);
or U11661 (N_11661,N_10936,N_10815);
or U11662 (N_11662,N_11111,N_11286);
and U11663 (N_11663,N_11353,N_10985);
xnor U11664 (N_11664,N_11259,N_10993);
and U11665 (N_11665,N_11173,N_11257);
nor U11666 (N_11666,N_11185,N_10966);
nor U11667 (N_11667,N_10868,N_10852);
or U11668 (N_11668,N_11115,N_10853);
or U11669 (N_11669,N_11033,N_11305);
and U11670 (N_11670,N_11278,N_11093);
and U11671 (N_11671,N_10835,N_11127);
or U11672 (N_11672,N_10806,N_11264);
xnor U11673 (N_11673,N_11054,N_10975);
or U11674 (N_11674,N_11101,N_11107);
nand U11675 (N_11675,N_10802,N_11011);
xnor U11676 (N_11676,N_10870,N_11132);
and U11677 (N_11677,N_11171,N_10858);
xor U11678 (N_11678,N_11149,N_11376);
and U11679 (N_11679,N_11236,N_11029);
or U11680 (N_11680,N_11323,N_11091);
and U11681 (N_11681,N_11258,N_11103);
nand U11682 (N_11682,N_10808,N_11164);
and U11683 (N_11683,N_11009,N_10968);
xor U11684 (N_11684,N_11339,N_11314);
or U11685 (N_11685,N_11122,N_11370);
nand U11686 (N_11686,N_11300,N_11024);
xnor U11687 (N_11687,N_11035,N_11266);
and U11688 (N_11688,N_11230,N_10883);
xor U11689 (N_11689,N_10977,N_10939);
or U11690 (N_11690,N_11120,N_11123);
nor U11691 (N_11691,N_11187,N_11150);
xor U11692 (N_11692,N_11078,N_11116);
nor U11693 (N_11693,N_10964,N_10944);
and U11694 (N_11694,N_10859,N_11279);
xnor U11695 (N_11695,N_10812,N_11206);
nand U11696 (N_11696,N_10915,N_11067);
and U11697 (N_11697,N_11182,N_11110);
nor U11698 (N_11698,N_11184,N_11010);
or U11699 (N_11699,N_11223,N_11359);
nand U11700 (N_11700,N_10944,N_11110);
and U11701 (N_11701,N_11360,N_11233);
and U11702 (N_11702,N_10868,N_10996);
nand U11703 (N_11703,N_10834,N_11314);
or U11704 (N_11704,N_10977,N_11010);
nor U11705 (N_11705,N_10913,N_11034);
or U11706 (N_11706,N_10867,N_11168);
and U11707 (N_11707,N_11356,N_11100);
nor U11708 (N_11708,N_10835,N_10867);
nand U11709 (N_11709,N_11390,N_11077);
xnor U11710 (N_11710,N_10810,N_11072);
or U11711 (N_11711,N_11074,N_11332);
and U11712 (N_11712,N_11154,N_11019);
xnor U11713 (N_11713,N_10865,N_11177);
nor U11714 (N_11714,N_11300,N_10880);
or U11715 (N_11715,N_11374,N_10853);
or U11716 (N_11716,N_10864,N_10865);
nand U11717 (N_11717,N_10807,N_11064);
nor U11718 (N_11718,N_11302,N_11071);
nand U11719 (N_11719,N_11130,N_11336);
and U11720 (N_11720,N_11193,N_11152);
nand U11721 (N_11721,N_11083,N_11267);
nor U11722 (N_11722,N_10998,N_10949);
and U11723 (N_11723,N_10885,N_11099);
or U11724 (N_11724,N_10964,N_10838);
nand U11725 (N_11725,N_11183,N_11259);
xor U11726 (N_11726,N_11084,N_10809);
or U11727 (N_11727,N_11194,N_11397);
nand U11728 (N_11728,N_11018,N_10865);
nand U11729 (N_11729,N_11354,N_10929);
or U11730 (N_11730,N_11226,N_11065);
nor U11731 (N_11731,N_10865,N_10912);
nand U11732 (N_11732,N_11224,N_11205);
and U11733 (N_11733,N_10920,N_10996);
and U11734 (N_11734,N_11097,N_10917);
and U11735 (N_11735,N_10873,N_11225);
nand U11736 (N_11736,N_10997,N_11226);
and U11737 (N_11737,N_11264,N_10820);
or U11738 (N_11738,N_10890,N_11025);
nor U11739 (N_11739,N_11072,N_11031);
and U11740 (N_11740,N_10809,N_10905);
or U11741 (N_11741,N_11241,N_11235);
nor U11742 (N_11742,N_11386,N_11359);
or U11743 (N_11743,N_11193,N_11239);
xor U11744 (N_11744,N_10806,N_11335);
or U11745 (N_11745,N_11283,N_11189);
and U11746 (N_11746,N_11240,N_10908);
xor U11747 (N_11747,N_11135,N_11251);
nor U11748 (N_11748,N_11218,N_10966);
and U11749 (N_11749,N_10892,N_11192);
or U11750 (N_11750,N_11223,N_11126);
xnor U11751 (N_11751,N_10931,N_11276);
or U11752 (N_11752,N_11095,N_11110);
or U11753 (N_11753,N_11130,N_11216);
nand U11754 (N_11754,N_11167,N_11057);
nand U11755 (N_11755,N_11233,N_11088);
xor U11756 (N_11756,N_11173,N_11008);
nor U11757 (N_11757,N_11241,N_11043);
xnor U11758 (N_11758,N_10967,N_11317);
nand U11759 (N_11759,N_11314,N_10979);
xnor U11760 (N_11760,N_11189,N_10890);
or U11761 (N_11761,N_11315,N_11238);
or U11762 (N_11762,N_11128,N_11362);
or U11763 (N_11763,N_10968,N_10879);
or U11764 (N_11764,N_11283,N_11083);
xnor U11765 (N_11765,N_11377,N_11339);
nand U11766 (N_11766,N_10862,N_10941);
nand U11767 (N_11767,N_11207,N_11185);
nand U11768 (N_11768,N_11316,N_11300);
or U11769 (N_11769,N_10939,N_10966);
and U11770 (N_11770,N_11059,N_11358);
nor U11771 (N_11771,N_11008,N_10874);
nand U11772 (N_11772,N_10971,N_10930);
nand U11773 (N_11773,N_11065,N_10814);
nand U11774 (N_11774,N_10868,N_11375);
xnor U11775 (N_11775,N_10952,N_11117);
nor U11776 (N_11776,N_10812,N_10824);
and U11777 (N_11777,N_11087,N_11061);
nor U11778 (N_11778,N_11105,N_11067);
nor U11779 (N_11779,N_10926,N_11178);
xor U11780 (N_11780,N_11068,N_11122);
xnor U11781 (N_11781,N_10900,N_11397);
and U11782 (N_11782,N_10825,N_11151);
xor U11783 (N_11783,N_11238,N_11221);
and U11784 (N_11784,N_11022,N_11333);
nor U11785 (N_11785,N_11222,N_10915);
and U11786 (N_11786,N_11175,N_11153);
nand U11787 (N_11787,N_11236,N_11072);
and U11788 (N_11788,N_11360,N_11175);
or U11789 (N_11789,N_11276,N_11289);
or U11790 (N_11790,N_11280,N_10996);
or U11791 (N_11791,N_11187,N_11164);
and U11792 (N_11792,N_10912,N_10821);
nand U11793 (N_11793,N_10813,N_10981);
and U11794 (N_11794,N_10896,N_10958);
nand U11795 (N_11795,N_10985,N_11299);
nor U11796 (N_11796,N_11292,N_11298);
nor U11797 (N_11797,N_11180,N_11242);
or U11798 (N_11798,N_11070,N_10963);
nand U11799 (N_11799,N_10823,N_11041);
nor U11800 (N_11800,N_11325,N_11067);
nand U11801 (N_11801,N_11216,N_11128);
nor U11802 (N_11802,N_11155,N_11355);
and U11803 (N_11803,N_10826,N_11341);
nor U11804 (N_11804,N_10912,N_11222);
and U11805 (N_11805,N_10868,N_11294);
xor U11806 (N_11806,N_10909,N_11387);
or U11807 (N_11807,N_11153,N_10967);
nand U11808 (N_11808,N_11256,N_11023);
nand U11809 (N_11809,N_10812,N_11317);
nor U11810 (N_11810,N_11071,N_11152);
or U11811 (N_11811,N_11042,N_10872);
xnor U11812 (N_11812,N_10922,N_11250);
nand U11813 (N_11813,N_10982,N_10827);
nor U11814 (N_11814,N_10960,N_11280);
nand U11815 (N_11815,N_11204,N_11284);
or U11816 (N_11816,N_10845,N_11070);
xor U11817 (N_11817,N_10841,N_11054);
nor U11818 (N_11818,N_11391,N_10947);
or U11819 (N_11819,N_11019,N_11033);
and U11820 (N_11820,N_11274,N_11132);
nand U11821 (N_11821,N_10861,N_10909);
or U11822 (N_11822,N_11180,N_10994);
nand U11823 (N_11823,N_10868,N_10895);
or U11824 (N_11824,N_11029,N_11101);
and U11825 (N_11825,N_11379,N_11164);
xor U11826 (N_11826,N_11300,N_11057);
or U11827 (N_11827,N_11191,N_10957);
xnor U11828 (N_11828,N_11165,N_10960);
nand U11829 (N_11829,N_10809,N_11251);
xnor U11830 (N_11830,N_11378,N_10809);
and U11831 (N_11831,N_11059,N_11158);
or U11832 (N_11832,N_11107,N_11104);
nor U11833 (N_11833,N_11278,N_11203);
nor U11834 (N_11834,N_11256,N_10946);
nor U11835 (N_11835,N_10809,N_11382);
nor U11836 (N_11836,N_11188,N_11173);
or U11837 (N_11837,N_11363,N_10834);
nand U11838 (N_11838,N_11122,N_11012);
xnor U11839 (N_11839,N_11185,N_11346);
nor U11840 (N_11840,N_11221,N_10847);
or U11841 (N_11841,N_11017,N_10899);
xnor U11842 (N_11842,N_10970,N_11368);
and U11843 (N_11843,N_10820,N_11357);
or U11844 (N_11844,N_11097,N_11245);
or U11845 (N_11845,N_11105,N_10831);
and U11846 (N_11846,N_11389,N_11246);
nor U11847 (N_11847,N_10932,N_11139);
nand U11848 (N_11848,N_10874,N_10867);
nand U11849 (N_11849,N_11183,N_10919);
and U11850 (N_11850,N_11373,N_11232);
nor U11851 (N_11851,N_11285,N_11388);
and U11852 (N_11852,N_10995,N_11128);
and U11853 (N_11853,N_10822,N_11226);
or U11854 (N_11854,N_10844,N_11383);
nor U11855 (N_11855,N_10859,N_11355);
xnor U11856 (N_11856,N_11374,N_11399);
and U11857 (N_11857,N_10992,N_10982);
nand U11858 (N_11858,N_10859,N_11337);
xnor U11859 (N_11859,N_10997,N_10859);
nor U11860 (N_11860,N_11394,N_10911);
or U11861 (N_11861,N_11084,N_11390);
or U11862 (N_11862,N_11288,N_11228);
nand U11863 (N_11863,N_11330,N_10966);
or U11864 (N_11864,N_11026,N_11024);
nand U11865 (N_11865,N_11071,N_11340);
and U11866 (N_11866,N_11370,N_10976);
xnor U11867 (N_11867,N_11040,N_11394);
nand U11868 (N_11868,N_11396,N_10916);
and U11869 (N_11869,N_10803,N_11054);
xor U11870 (N_11870,N_11005,N_11096);
nand U11871 (N_11871,N_10905,N_10883);
xnor U11872 (N_11872,N_10871,N_10899);
and U11873 (N_11873,N_11315,N_10809);
and U11874 (N_11874,N_10860,N_11388);
nor U11875 (N_11875,N_10958,N_11129);
xnor U11876 (N_11876,N_11167,N_10860);
nor U11877 (N_11877,N_10968,N_11055);
nand U11878 (N_11878,N_11203,N_11381);
nor U11879 (N_11879,N_11240,N_11171);
or U11880 (N_11880,N_11178,N_11227);
nor U11881 (N_11881,N_11197,N_11252);
and U11882 (N_11882,N_10828,N_11051);
and U11883 (N_11883,N_10958,N_11052);
or U11884 (N_11884,N_10919,N_11004);
nor U11885 (N_11885,N_10980,N_11325);
or U11886 (N_11886,N_11182,N_10958);
nand U11887 (N_11887,N_11366,N_10954);
nand U11888 (N_11888,N_11327,N_10985);
or U11889 (N_11889,N_11093,N_11088);
and U11890 (N_11890,N_11344,N_11249);
nor U11891 (N_11891,N_10907,N_10999);
nor U11892 (N_11892,N_10999,N_11258);
xor U11893 (N_11893,N_11254,N_11017);
or U11894 (N_11894,N_11303,N_10933);
and U11895 (N_11895,N_11219,N_10800);
nor U11896 (N_11896,N_11207,N_11189);
nor U11897 (N_11897,N_10941,N_11032);
nor U11898 (N_11898,N_11044,N_11369);
or U11899 (N_11899,N_10958,N_10904);
nand U11900 (N_11900,N_11390,N_10867);
and U11901 (N_11901,N_10963,N_11361);
or U11902 (N_11902,N_11066,N_11304);
and U11903 (N_11903,N_11242,N_10958);
and U11904 (N_11904,N_10974,N_11115);
nand U11905 (N_11905,N_11271,N_11260);
xor U11906 (N_11906,N_10888,N_11102);
xor U11907 (N_11907,N_11047,N_11334);
nor U11908 (N_11908,N_11032,N_11146);
nor U11909 (N_11909,N_11005,N_11028);
nand U11910 (N_11910,N_10841,N_10861);
nand U11911 (N_11911,N_10843,N_10996);
xnor U11912 (N_11912,N_11350,N_10854);
or U11913 (N_11913,N_11023,N_11058);
nand U11914 (N_11914,N_11080,N_10805);
nand U11915 (N_11915,N_11269,N_11059);
and U11916 (N_11916,N_10833,N_11370);
nand U11917 (N_11917,N_11059,N_11159);
xnor U11918 (N_11918,N_11279,N_10889);
xor U11919 (N_11919,N_10833,N_10804);
and U11920 (N_11920,N_11339,N_11176);
or U11921 (N_11921,N_11173,N_11236);
nand U11922 (N_11922,N_11311,N_11251);
and U11923 (N_11923,N_10850,N_11299);
or U11924 (N_11924,N_10989,N_11004);
nand U11925 (N_11925,N_11373,N_11324);
and U11926 (N_11926,N_11012,N_10975);
and U11927 (N_11927,N_11072,N_11068);
xor U11928 (N_11928,N_10946,N_11346);
and U11929 (N_11929,N_11270,N_10914);
nand U11930 (N_11930,N_10820,N_10824);
xnor U11931 (N_11931,N_11007,N_10858);
nor U11932 (N_11932,N_10825,N_11025);
xor U11933 (N_11933,N_10957,N_11393);
or U11934 (N_11934,N_11087,N_10906);
or U11935 (N_11935,N_10834,N_11367);
or U11936 (N_11936,N_10836,N_11226);
nand U11937 (N_11937,N_10909,N_10906);
or U11938 (N_11938,N_11020,N_10981);
and U11939 (N_11939,N_11316,N_11232);
xnor U11940 (N_11940,N_10988,N_11067);
nand U11941 (N_11941,N_11113,N_11390);
and U11942 (N_11942,N_11087,N_10828);
nand U11943 (N_11943,N_11306,N_11239);
xor U11944 (N_11944,N_10988,N_11198);
nor U11945 (N_11945,N_11137,N_11114);
nand U11946 (N_11946,N_10821,N_11316);
nor U11947 (N_11947,N_10902,N_11003);
nand U11948 (N_11948,N_11260,N_11306);
nor U11949 (N_11949,N_11249,N_11189);
xnor U11950 (N_11950,N_11346,N_11231);
and U11951 (N_11951,N_11171,N_11283);
nor U11952 (N_11952,N_11051,N_11162);
nor U11953 (N_11953,N_11158,N_11029);
and U11954 (N_11954,N_11325,N_11208);
xor U11955 (N_11955,N_11051,N_11347);
nor U11956 (N_11956,N_11102,N_11016);
xnor U11957 (N_11957,N_11197,N_10982);
and U11958 (N_11958,N_11159,N_11252);
nor U11959 (N_11959,N_10826,N_11349);
nor U11960 (N_11960,N_11385,N_11164);
and U11961 (N_11961,N_11237,N_11319);
xor U11962 (N_11962,N_10808,N_11310);
nand U11963 (N_11963,N_10870,N_10950);
nor U11964 (N_11964,N_10957,N_11045);
nand U11965 (N_11965,N_11062,N_11034);
xor U11966 (N_11966,N_11019,N_10953);
and U11967 (N_11967,N_11148,N_11293);
or U11968 (N_11968,N_11223,N_11242);
nand U11969 (N_11969,N_11029,N_11039);
nand U11970 (N_11970,N_11272,N_11350);
or U11971 (N_11971,N_11049,N_10998);
or U11972 (N_11972,N_11143,N_11219);
or U11973 (N_11973,N_11162,N_11056);
nand U11974 (N_11974,N_10934,N_10857);
or U11975 (N_11975,N_11214,N_10868);
or U11976 (N_11976,N_10970,N_10920);
or U11977 (N_11977,N_11385,N_10825);
or U11978 (N_11978,N_11223,N_11190);
xor U11979 (N_11979,N_11314,N_11049);
nor U11980 (N_11980,N_10800,N_11069);
and U11981 (N_11981,N_10987,N_11328);
nor U11982 (N_11982,N_11055,N_11188);
and U11983 (N_11983,N_11178,N_11109);
nand U11984 (N_11984,N_11303,N_11361);
xor U11985 (N_11985,N_11044,N_11159);
nand U11986 (N_11986,N_11239,N_10892);
or U11987 (N_11987,N_11348,N_11048);
nor U11988 (N_11988,N_10929,N_11313);
xnor U11989 (N_11989,N_10945,N_10936);
nor U11990 (N_11990,N_11227,N_11375);
nor U11991 (N_11991,N_10952,N_11075);
and U11992 (N_11992,N_11154,N_10956);
or U11993 (N_11993,N_10867,N_11251);
xor U11994 (N_11994,N_11388,N_11028);
nand U11995 (N_11995,N_10889,N_10862);
nand U11996 (N_11996,N_10933,N_11034);
or U11997 (N_11997,N_11091,N_10888);
xnor U11998 (N_11998,N_11292,N_11379);
xnor U11999 (N_11999,N_11290,N_11330);
xnor U12000 (N_12000,N_11798,N_11859);
nand U12001 (N_12001,N_11587,N_11541);
or U12002 (N_12002,N_11589,N_11494);
nand U12003 (N_12003,N_11847,N_11882);
nand U12004 (N_12004,N_11762,N_11921);
or U12005 (N_12005,N_11715,N_11567);
nand U12006 (N_12006,N_11414,N_11790);
nand U12007 (N_12007,N_11665,N_11938);
nand U12008 (N_12008,N_11875,N_11581);
or U12009 (N_12009,N_11559,N_11879);
nand U12010 (N_12010,N_11810,N_11582);
nand U12011 (N_12011,N_11677,N_11680);
xnor U12012 (N_12012,N_11966,N_11732);
nor U12013 (N_12013,N_11949,N_11770);
nand U12014 (N_12014,N_11603,N_11964);
xnor U12015 (N_12015,N_11661,N_11422);
xor U12016 (N_12016,N_11572,N_11924);
or U12017 (N_12017,N_11591,N_11459);
and U12018 (N_12018,N_11411,N_11534);
nor U12019 (N_12019,N_11473,N_11409);
nor U12020 (N_12020,N_11779,N_11830);
and U12021 (N_12021,N_11918,N_11638);
and U12022 (N_12022,N_11975,N_11834);
and U12023 (N_12023,N_11471,N_11520);
xnor U12024 (N_12024,N_11944,N_11728);
nand U12025 (N_12025,N_11961,N_11526);
or U12026 (N_12026,N_11963,N_11888);
nand U12027 (N_12027,N_11626,N_11740);
xor U12028 (N_12028,N_11537,N_11861);
or U12029 (N_12029,N_11495,N_11590);
and U12030 (N_12030,N_11605,N_11672);
xnor U12031 (N_12031,N_11687,N_11977);
or U12032 (N_12032,N_11693,N_11907);
and U12033 (N_12033,N_11768,N_11448);
xor U12034 (N_12034,N_11923,N_11983);
xnor U12035 (N_12035,N_11652,N_11931);
and U12036 (N_12036,N_11701,N_11857);
xor U12037 (N_12037,N_11992,N_11842);
nand U12038 (N_12038,N_11576,N_11998);
or U12039 (N_12039,N_11664,N_11926);
xnor U12040 (N_12040,N_11816,N_11507);
nand U12041 (N_12041,N_11848,N_11497);
or U12042 (N_12042,N_11408,N_11979);
nor U12043 (N_12043,N_11791,N_11633);
nand U12044 (N_12044,N_11438,N_11556);
nor U12045 (N_12045,N_11549,N_11630);
xor U12046 (N_12046,N_11838,N_11837);
and U12047 (N_12047,N_11872,N_11984);
or U12048 (N_12048,N_11855,N_11538);
xnor U12049 (N_12049,N_11464,N_11851);
xnor U12050 (N_12050,N_11955,N_11897);
or U12051 (N_12051,N_11500,N_11407);
nand U12052 (N_12052,N_11731,N_11906);
or U12053 (N_12053,N_11551,N_11472);
or U12054 (N_12054,N_11939,N_11825);
or U12055 (N_12055,N_11801,N_11694);
nand U12056 (N_12056,N_11917,N_11635);
or U12057 (N_12057,N_11719,N_11666);
nor U12058 (N_12058,N_11706,N_11609);
nand U12059 (N_12059,N_11583,N_11739);
xor U12060 (N_12060,N_11783,N_11795);
and U12061 (N_12061,N_11487,N_11807);
and U12062 (N_12062,N_11442,N_11533);
or U12063 (N_12063,N_11668,N_11584);
nand U12064 (N_12064,N_11451,N_11742);
and U12065 (N_12065,N_11714,N_11686);
xor U12066 (N_12066,N_11615,N_11824);
xnor U12067 (N_12067,N_11894,N_11458);
nand U12068 (N_12068,N_11593,N_11822);
or U12069 (N_12069,N_11622,N_11539);
nand U12070 (N_12070,N_11699,N_11829);
or U12071 (N_12071,N_11521,N_11936);
or U12072 (N_12072,N_11456,N_11821);
xor U12073 (N_12073,N_11692,N_11815);
or U12074 (N_12074,N_11493,N_11952);
and U12075 (N_12075,N_11475,N_11440);
or U12076 (N_12076,N_11889,N_11958);
nor U12077 (N_12077,N_11695,N_11419);
nor U12078 (N_12078,N_11702,N_11771);
and U12079 (N_12079,N_11483,N_11972);
xor U12080 (N_12080,N_11683,N_11647);
nor U12081 (N_12081,N_11571,N_11988);
nand U12082 (N_12082,N_11737,N_11913);
xor U12083 (N_12083,N_11654,N_11545);
nor U12084 (N_12084,N_11457,N_11928);
nand U12085 (N_12085,N_11621,N_11981);
nand U12086 (N_12086,N_11788,N_11579);
nand U12087 (N_12087,N_11707,N_11513);
nand U12088 (N_12088,N_11649,N_11951);
nor U12089 (N_12089,N_11767,N_11905);
nor U12090 (N_12090,N_11434,N_11772);
xor U12091 (N_12091,N_11712,N_11748);
or U12092 (N_12092,N_11887,N_11896);
xnor U12093 (N_12093,N_11523,N_11566);
nand U12094 (N_12094,N_11827,N_11515);
or U12095 (N_12095,N_11417,N_11508);
nor U12096 (N_12096,N_11789,N_11999);
xor U12097 (N_12097,N_11841,N_11540);
nand U12098 (N_12098,N_11580,N_11643);
xnor U12099 (N_12099,N_11718,N_11902);
xnor U12100 (N_12100,N_11929,N_11602);
or U12101 (N_12101,N_11900,N_11467);
xnor U12102 (N_12102,N_11480,N_11527);
or U12103 (N_12103,N_11849,N_11404);
xor U12104 (N_12104,N_11642,N_11890);
xnor U12105 (N_12105,N_11997,N_11685);
xor U12106 (N_12106,N_11738,N_11839);
or U12107 (N_12107,N_11836,N_11619);
and U12108 (N_12108,N_11820,N_11747);
and U12109 (N_12109,N_11563,N_11430);
nand U12110 (N_12110,N_11607,N_11753);
and U12111 (N_12111,N_11943,N_11852);
nand U12112 (N_12112,N_11736,N_11594);
nor U12113 (N_12113,N_11973,N_11794);
and U12114 (N_12114,N_11976,N_11778);
xnor U12115 (N_12115,N_11752,N_11443);
nor U12116 (N_12116,N_11991,N_11750);
nor U12117 (N_12117,N_11460,N_11751);
nor U12118 (N_12118,N_11802,N_11968);
and U12119 (N_12119,N_11546,N_11805);
nand U12120 (N_12120,N_11756,N_11780);
or U12121 (N_12121,N_11700,N_11624);
nor U12122 (N_12122,N_11477,N_11974);
nor U12123 (N_12123,N_11575,N_11877);
nor U12124 (N_12124,N_11588,N_11416);
or U12125 (N_12125,N_11560,N_11985);
nand U12126 (N_12126,N_11604,N_11444);
xor U12127 (N_12127,N_11421,N_11479);
and U12128 (N_12128,N_11755,N_11623);
and U12129 (N_12129,N_11793,N_11782);
xor U12130 (N_12130,N_11862,N_11501);
nand U12131 (N_12131,N_11696,N_11959);
or U12132 (N_12132,N_11452,N_11990);
nand U12133 (N_12133,N_11804,N_11598);
nand U12134 (N_12134,N_11843,N_11758);
or U12135 (N_12135,N_11530,N_11415);
xor U12136 (N_12136,N_11490,N_11558);
nand U12137 (N_12137,N_11858,N_11646);
and U12138 (N_12138,N_11403,N_11550);
xnor U12139 (N_12139,N_11504,N_11616);
nand U12140 (N_12140,N_11595,N_11965);
and U12141 (N_12141,N_11678,N_11450);
nor U12142 (N_12142,N_11697,N_11453);
nor U12143 (N_12143,N_11412,N_11568);
or U12144 (N_12144,N_11406,N_11811);
and U12145 (N_12145,N_11785,N_11818);
nor U12146 (N_12146,N_11760,N_11667);
or U12147 (N_12147,N_11611,N_11657);
xnor U12148 (N_12148,N_11759,N_11639);
and U12149 (N_12149,N_11812,N_11831);
and U12150 (N_12150,N_11846,N_11691);
or U12151 (N_12151,N_11627,N_11764);
xor U12152 (N_12152,N_11726,N_11925);
nor U12153 (N_12153,N_11514,N_11844);
xor U12154 (N_12154,N_11532,N_11987);
and U12155 (N_12155,N_11826,N_11993);
or U12156 (N_12156,N_11465,N_11916);
and U12157 (N_12157,N_11784,N_11437);
and U12158 (N_12158,N_11863,N_11424);
nand U12159 (N_12159,N_11431,N_11651);
nor U12160 (N_12160,N_11488,N_11787);
and U12161 (N_12161,N_11729,N_11865);
nand U12162 (N_12162,N_11734,N_11813);
xor U12163 (N_12163,N_11854,N_11806);
nor U12164 (N_12164,N_11553,N_11895);
and U12165 (N_12165,N_11721,N_11561);
nand U12166 (N_12166,N_11708,N_11565);
nor U12167 (N_12167,N_11915,N_11524);
nand U12168 (N_12168,N_11880,N_11876);
and U12169 (N_12169,N_11586,N_11542);
or U12170 (N_12170,N_11934,N_11727);
xor U12171 (N_12171,N_11632,N_11552);
nand U12172 (N_12172,N_11884,N_11569);
nand U12173 (N_12173,N_11625,N_11933);
nand U12174 (N_12174,N_11850,N_11620);
xor U12175 (N_12175,N_11942,N_11613);
nor U12176 (N_12176,N_11413,N_11946);
or U12177 (N_12177,N_11600,N_11585);
xor U12178 (N_12178,N_11903,N_11833);
nor U12179 (N_12179,N_11468,N_11645);
or U12180 (N_12180,N_11673,N_11948);
and U12181 (N_12181,N_11835,N_11786);
or U12182 (N_12182,N_11466,N_11423);
or U12183 (N_12183,N_11893,N_11484);
nor U12184 (N_12184,N_11814,N_11864);
nand U12185 (N_12185,N_11428,N_11447);
xor U12186 (N_12186,N_11935,N_11745);
nor U12187 (N_12187,N_11910,N_11891);
nor U12188 (N_12188,N_11525,N_11986);
nand U12189 (N_12189,N_11486,N_11631);
nand U12190 (N_12190,N_11743,N_11867);
or U12191 (N_12191,N_11769,N_11912);
xnor U12192 (N_12192,N_11474,N_11860);
nand U12193 (N_12193,N_11716,N_11761);
and U12194 (N_12194,N_11420,N_11445);
and U12195 (N_12195,N_11655,N_11796);
xnor U12196 (N_12196,N_11710,N_11754);
nand U12197 (N_12197,N_11911,N_11774);
nand U12198 (N_12198,N_11690,N_11644);
nand U12199 (N_12199,N_11883,N_11427);
nand U12200 (N_12200,N_11792,N_11711);
and U12201 (N_12201,N_11953,N_11868);
or U12202 (N_12202,N_11511,N_11809);
xor U12203 (N_12203,N_11596,N_11578);
or U12204 (N_12204,N_11410,N_11485);
and U12205 (N_12205,N_11722,N_11828);
xnor U12206 (N_12206,N_11512,N_11509);
or U12207 (N_12207,N_11717,N_11971);
and U12208 (N_12208,N_11989,N_11954);
nand U12209 (N_12209,N_11491,N_11724);
xnor U12210 (N_12210,N_11950,N_11922);
nand U12211 (N_12211,N_11544,N_11461);
nand U12212 (N_12212,N_11670,N_11777);
nand U12213 (N_12213,N_11522,N_11592);
nor U12214 (N_12214,N_11455,N_11940);
nor U12215 (N_12215,N_11597,N_11703);
and U12216 (N_12216,N_11531,N_11573);
nor U12217 (N_12217,N_11577,N_11817);
or U12218 (N_12218,N_11698,N_11684);
xor U12219 (N_12219,N_11557,N_11823);
nor U12220 (N_12220,N_11470,N_11874);
nand U12221 (N_12221,N_11709,N_11776);
nor U12222 (N_12222,N_11618,N_11648);
or U12223 (N_12223,N_11932,N_11658);
nor U12224 (N_12224,N_11969,N_11808);
nand U12225 (N_12225,N_11614,N_11519);
nor U12226 (N_12226,N_11505,N_11629);
nor U12227 (N_12227,N_11892,N_11775);
xnor U12228 (N_12228,N_11967,N_11898);
xor U12229 (N_12229,N_11555,N_11528);
or U12230 (N_12230,N_11489,N_11741);
nand U12231 (N_12231,N_11871,N_11446);
xnor U12232 (N_12232,N_11870,N_11634);
nor U12233 (N_12233,N_11640,N_11401);
nor U12234 (N_12234,N_11496,N_11994);
xnor U12235 (N_12235,N_11713,N_11919);
nand U12236 (N_12236,N_11636,N_11612);
and U12237 (N_12237,N_11886,N_11982);
xnor U12238 (N_12238,N_11679,N_11904);
nand U12239 (N_12239,N_11881,N_11650);
xnor U12240 (N_12240,N_11536,N_11773);
xor U12241 (N_12241,N_11766,N_11856);
and U12242 (N_12242,N_11425,N_11744);
or U12243 (N_12243,N_11995,N_11853);
or U12244 (N_12244,N_11462,N_11832);
or U12245 (N_12245,N_11405,N_11962);
nand U12246 (N_12246,N_11681,N_11562);
nor U12247 (N_12247,N_11869,N_11941);
or U12248 (N_12248,N_11720,N_11418);
nand U12249 (N_12249,N_11733,N_11518);
or U12250 (N_12250,N_11878,N_11749);
or U12251 (N_12251,N_11601,N_11476);
xor U12252 (N_12252,N_11840,N_11705);
or U12253 (N_12253,N_11502,N_11873);
xnor U12254 (N_12254,N_11937,N_11400);
or U12255 (N_12255,N_11960,N_11660);
and U12256 (N_12256,N_11803,N_11606);
and U12257 (N_12257,N_11980,N_11481);
nor U12258 (N_12258,N_11548,N_11449);
and U12259 (N_12259,N_11506,N_11503);
xor U12260 (N_12260,N_11757,N_11671);
nor U12261 (N_12261,N_11689,N_11432);
xor U12262 (N_12262,N_11516,N_11970);
and U12263 (N_12263,N_11996,N_11725);
nor U12264 (N_12264,N_11426,N_11441);
xnor U12265 (N_12265,N_11429,N_11662);
xor U12266 (N_12266,N_11763,N_11510);
or U12267 (N_12267,N_11899,N_11730);
xnor U12268 (N_12268,N_11535,N_11599);
nand U12269 (N_12269,N_11433,N_11439);
or U12270 (N_12270,N_11653,N_11800);
xor U12271 (N_12271,N_11735,N_11908);
xnor U12272 (N_12272,N_11463,N_11676);
nor U12273 (N_12273,N_11617,N_11608);
xor U12274 (N_12274,N_11704,N_11517);
or U12275 (N_12275,N_11947,N_11957);
or U12276 (N_12276,N_11628,N_11688);
or U12277 (N_12277,N_11920,N_11498);
and U12278 (N_12278,N_11765,N_11656);
nor U12279 (N_12279,N_11885,N_11570);
or U12280 (N_12280,N_11435,N_11564);
xnor U12281 (N_12281,N_11674,N_11547);
xnor U12282 (N_12282,N_11675,N_11799);
nand U12283 (N_12283,N_11492,N_11641);
nor U12284 (N_12284,N_11499,N_11543);
and U12285 (N_12285,N_11574,N_11682);
xnor U12286 (N_12286,N_11482,N_11781);
nor U12287 (N_12287,N_11436,N_11402);
xor U12288 (N_12288,N_11663,N_11554);
nor U12289 (N_12289,N_11845,N_11945);
nand U12290 (N_12290,N_11723,N_11469);
xor U12291 (N_12291,N_11659,N_11956);
and U12292 (N_12292,N_11819,N_11610);
nor U12293 (N_12293,N_11914,N_11746);
nor U12294 (N_12294,N_11637,N_11454);
and U12295 (N_12295,N_11529,N_11927);
and U12296 (N_12296,N_11978,N_11866);
nor U12297 (N_12297,N_11901,N_11669);
and U12298 (N_12298,N_11478,N_11930);
nand U12299 (N_12299,N_11909,N_11797);
nor U12300 (N_12300,N_11799,N_11885);
nor U12301 (N_12301,N_11898,N_11753);
or U12302 (N_12302,N_11934,N_11542);
or U12303 (N_12303,N_11858,N_11565);
nand U12304 (N_12304,N_11608,N_11719);
nor U12305 (N_12305,N_11647,N_11821);
nand U12306 (N_12306,N_11680,N_11587);
nand U12307 (N_12307,N_11597,N_11430);
nand U12308 (N_12308,N_11528,N_11885);
nand U12309 (N_12309,N_11930,N_11815);
nand U12310 (N_12310,N_11758,N_11974);
or U12311 (N_12311,N_11925,N_11932);
and U12312 (N_12312,N_11401,N_11636);
and U12313 (N_12313,N_11873,N_11884);
nand U12314 (N_12314,N_11714,N_11670);
nor U12315 (N_12315,N_11514,N_11912);
and U12316 (N_12316,N_11879,N_11931);
or U12317 (N_12317,N_11443,N_11847);
and U12318 (N_12318,N_11483,N_11848);
xnor U12319 (N_12319,N_11797,N_11716);
xnor U12320 (N_12320,N_11900,N_11682);
nor U12321 (N_12321,N_11790,N_11452);
nor U12322 (N_12322,N_11913,N_11587);
xor U12323 (N_12323,N_11781,N_11949);
nand U12324 (N_12324,N_11970,N_11770);
xnor U12325 (N_12325,N_11613,N_11466);
or U12326 (N_12326,N_11993,N_11972);
nor U12327 (N_12327,N_11742,N_11476);
nand U12328 (N_12328,N_11785,N_11956);
nor U12329 (N_12329,N_11439,N_11516);
and U12330 (N_12330,N_11566,N_11586);
or U12331 (N_12331,N_11419,N_11913);
or U12332 (N_12332,N_11737,N_11452);
xnor U12333 (N_12333,N_11626,N_11704);
nand U12334 (N_12334,N_11406,N_11790);
xor U12335 (N_12335,N_11663,N_11612);
or U12336 (N_12336,N_11947,N_11675);
xnor U12337 (N_12337,N_11738,N_11471);
xnor U12338 (N_12338,N_11534,N_11561);
nand U12339 (N_12339,N_11595,N_11474);
or U12340 (N_12340,N_11827,N_11420);
nand U12341 (N_12341,N_11473,N_11557);
nor U12342 (N_12342,N_11604,N_11442);
xnor U12343 (N_12343,N_11837,N_11991);
nand U12344 (N_12344,N_11508,N_11790);
nand U12345 (N_12345,N_11739,N_11921);
or U12346 (N_12346,N_11488,N_11566);
xor U12347 (N_12347,N_11756,N_11491);
and U12348 (N_12348,N_11900,N_11438);
nor U12349 (N_12349,N_11774,N_11981);
or U12350 (N_12350,N_11565,N_11787);
and U12351 (N_12351,N_11541,N_11807);
and U12352 (N_12352,N_11670,N_11550);
nor U12353 (N_12353,N_11862,N_11870);
nand U12354 (N_12354,N_11839,N_11873);
nand U12355 (N_12355,N_11765,N_11564);
or U12356 (N_12356,N_11486,N_11519);
or U12357 (N_12357,N_11741,N_11628);
nand U12358 (N_12358,N_11949,N_11719);
xor U12359 (N_12359,N_11674,N_11524);
nor U12360 (N_12360,N_11676,N_11752);
or U12361 (N_12361,N_11734,N_11798);
or U12362 (N_12362,N_11659,N_11873);
xor U12363 (N_12363,N_11523,N_11953);
or U12364 (N_12364,N_11876,N_11719);
nor U12365 (N_12365,N_11469,N_11893);
xor U12366 (N_12366,N_11822,N_11681);
nand U12367 (N_12367,N_11576,N_11602);
nand U12368 (N_12368,N_11781,N_11635);
xor U12369 (N_12369,N_11805,N_11917);
nand U12370 (N_12370,N_11497,N_11644);
and U12371 (N_12371,N_11515,N_11555);
or U12372 (N_12372,N_11722,N_11897);
or U12373 (N_12373,N_11552,N_11780);
xor U12374 (N_12374,N_11750,N_11774);
or U12375 (N_12375,N_11657,N_11445);
xor U12376 (N_12376,N_11667,N_11460);
xnor U12377 (N_12377,N_11427,N_11509);
or U12378 (N_12378,N_11524,N_11944);
nand U12379 (N_12379,N_11953,N_11707);
nor U12380 (N_12380,N_11808,N_11432);
nand U12381 (N_12381,N_11788,N_11873);
nand U12382 (N_12382,N_11806,N_11482);
nor U12383 (N_12383,N_11951,N_11410);
nand U12384 (N_12384,N_11628,N_11737);
nand U12385 (N_12385,N_11880,N_11620);
nor U12386 (N_12386,N_11555,N_11430);
and U12387 (N_12387,N_11719,N_11532);
or U12388 (N_12388,N_11988,N_11712);
nand U12389 (N_12389,N_11869,N_11825);
nand U12390 (N_12390,N_11964,N_11656);
xor U12391 (N_12391,N_11629,N_11428);
or U12392 (N_12392,N_11664,N_11921);
nor U12393 (N_12393,N_11999,N_11645);
nand U12394 (N_12394,N_11940,N_11631);
nor U12395 (N_12395,N_11983,N_11579);
xor U12396 (N_12396,N_11844,N_11588);
and U12397 (N_12397,N_11586,N_11971);
nor U12398 (N_12398,N_11870,N_11786);
nor U12399 (N_12399,N_11497,N_11875);
nand U12400 (N_12400,N_11781,N_11490);
xnor U12401 (N_12401,N_11419,N_11499);
nand U12402 (N_12402,N_11976,N_11973);
xnor U12403 (N_12403,N_11806,N_11855);
or U12404 (N_12404,N_11538,N_11727);
xor U12405 (N_12405,N_11687,N_11706);
xnor U12406 (N_12406,N_11793,N_11811);
or U12407 (N_12407,N_11538,N_11858);
xnor U12408 (N_12408,N_11766,N_11873);
or U12409 (N_12409,N_11940,N_11463);
xnor U12410 (N_12410,N_11719,N_11477);
and U12411 (N_12411,N_11438,N_11725);
nor U12412 (N_12412,N_11495,N_11512);
and U12413 (N_12413,N_11424,N_11927);
and U12414 (N_12414,N_11963,N_11729);
or U12415 (N_12415,N_11650,N_11432);
and U12416 (N_12416,N_11651,N_11533);
or U12417 (N_12417,N_11851,N_11658);
xnor U12418 (N_12418,N_11636,N_11425);
xnor U12419 (N_12419,N_11619,N_11812);
or U12420 (N_12420,N_11955,N_11607);
nand U12421 (N_12421,N_11472,N_11968);
and U12422 (N_12422,N_11621,N_11576);
nor U12423 (N_12423,N_11844,N_11930);
or U12424 (N_12424,N_11740,N_11596);
and U12425 (N_12425,N_11953,N_11846);
or U12426 (N_12426,N_11743,N_11721);
or U12427 (N_12427,N_11960,N_11418);
nor U12428 (N_12428,N_11927,N_11962);
nor U12429 (N_12429,N_11885,N_11993);
xor U12430 (N_12430,N_11754,N_11670);
nor U12431 (N_12431,N_11715,N_11446);
xnor U12432 (N_12432,N_11845,N_11463);
nor U12433 (N_12433,N_11851,N_11848);
nor U12434 (N_12434,N_11892,N_11407);
nand U12435 (N_12435,N_11510,N_11420);
or U12436 (N_12436,N_11528,N_11633);
xor U12437 (N_12437,N_11484,N_11932);
nand U12438 (N_12438,N_11747,N_11452);
and U12439 (N_12439,N_11493,N_11432);
xor U12440 (N_12440,N_11623,N_11465);
xnor U12441 (N_12441,N_11594,N_11857);
or U12442 (N_12442,N_11575,N_11529);
or U12443 (N_12443,N_11591,N_11509);
nor U12444 (N_12444,N_11446,N_11830);
nand U12445 (N_12445,N_11576,N_11788);
and U12446 (N_12446,N_11535,N_11690);
and U12447 (N_12447,N_11668,N_11459);
nor U12448 (N_12448,N_11547,N_11445);
nor U12449 (N_12449,N_11478,N_11444);
or U12450 (N_12450,N_11746,N_11703);
nand U12451 (N_12451,N_11891,N_11963);
and U12452 (N_12452,N_11656,N_11741);
and U12453 (N_12453,N_11998,N_11736);
nand U12454 (N_12454,N_11577,N_11508);
nand U12455 (N_12455,N_11811,N_11610);
or U12456 (N_12456,N_11666,N_11893);
nand U12457 (N_12457,N_11703,N_11971);
xnor U12458 (N_12458,N_11673,N_11949);
or U12459 (N_12459,N_11868,N_11473);
nor U12460 (N_12460,N_11459,N_11425);
nand U12461 (N_12461,N_11814,N_11473);
nand U12462 (N_12462,N_11757,N_11698);
xor U12463 (N_12463,N_11511,N_11810);
and U12464 (N_12464,N_11488,N_11733);
nor U12465 (N_12465,N_11503,N_11822);
xnor U12466 (N_12466,N_11728,N_11551);
or U12467 (N_12467,N_11441,N_11419);
nand U12468 (N_12468,N_11616,N_11638);
or U12469 (N_12469,N_11974,N_11686);
or U12470 (N_12470,N_11625,N_11527);
nand U12471 (N_12471,N_11539,N_11763);
nor U12472 (N_12472,N_11486,N_11456);
nand U12473 (N_12473,N_11948,N_11549);
or U12474 (N_12474,N_11773,N_11753);
nor U12475 (N_12475,N_11516,N_11758);
and U12476 (N_12476,N_11546,N_11737);
xor U12477 (N_12477,N_11489,N_11861);
nand U12478 (N_12478,N_11681,N_11664);
nand U12479 (N_12479,N_11447,N_11590);
nand U12480 (N_12480,N_11908,N_11610);
nand U12481 (N_12481,N_11845,N_11833);
xnor U12482 (N_12482,N_11922,N_11628);
nand U12483 (N_12483,N_11817,N_11813);
nor U12484 (N_12484,N_11603,N_11708);
and U12485 (N_12485,N_11834,N_11998);
nand U12486 (N_12486,N_11657,N_11476);
xor U12487 (N_12487,N_11722,N_11839);
nand U12488 (N_12488,N_11751,N_11659);
or U12489 (N_12489,N_11760,N_11673);
or U12490 (N_12490,N_11735,N_11931);
nor U12491 (N_12491,N_11484,N_11732);
and U12492 (N_12492,N_11468,N_11996);
nor U12493 (N_12493,N_11829,N_11498);
nor U12494 (N_12494,N_11698,N_11969);
xnor U12495 (N_12495,N_11513,N_11767);
or U12496 (N_12496,N_11726,N_11618);
nand U12497 (N_12497,N_11623,N_11431);
nand U12498 (N_12498,N_11964,N_11579);
xor U12499 (N_12499,N_11423,N_11995);
and U12500 (N_12500,N_11892,N_11731);
nand U12501 (N_12501,N_11457,N_11638);
nor U12502 (N_12502,N_11483,N_11663);
nand U12503 (N_12503,N_11610,N_11406);
nand U12504 (N_12504,N_11944,N_11938);
or U12505 (N_12505,N_11740,N_11486);
or U12506 (N_12506,N_11649,N_11624);
and U12507 (N_12507,N_11627,N_11895);
nand U12508 (N_12508,N_11561,N_11820);
or U12509 (N_12509,N_11565,N_11905);
nor U12510 (N_12510,N_11461,N_11581);
or U12511 (N_12511,N_11936,N_11990);
xnor U12512 (N_12512,N_11931,N_11483);
nor U12513 (N_12513,N_11954,N_11994);
and U12514 (N_12514,N_11427,N_11490);
nor U12515 (N_12515,N_11823,N_11625);
xor U12516 (N_12516,N_11957,N_11964);
and U12517 (N_12517,N_11795,N_11767);
nor U12518 (N_12518,N_11795,N_11645);
nor U12519 (N_12519,N_11739,N_11526);
and U12520 (N_12520,N_11983,N_11878);
nand U12521 (N_12521,N_11422,N_11494);
xor U12522 (N_12522,N_11860,N_11575);
xor U12523 (N_12523,N_11956,N_11616);
nor U12524 (N_12524,N_11700,N_11760);
and U12525 (N_12525,N_11822,N_11407);
and U12526 (N_12526,N_11916,N_11852);
or U12527 (N_12527,N_11976,N_11611);
and U12528 (N_12528,N_11735,N_11808);
xor U12529 (N_12529,N_11963,N_11432);
nor U12530 (N_12530,N_11486,N_11531);
nor U12531 (N_12531,N_11536,N_11858);
and U12532 (N_12532,N_11473,N_11628);
or U12533 (N_12533,N_11891,N_11729);
nor U12534 (N_12534,N_11997,N_11944);
xor U12535 (N_12535,N_11440,N_11744);
and U12536 (N_12536,N_11505,N_11514);
xor U12537 (N_12537,N_11554,N_11425);
and U12538 (N_12538,N_11750,N_11511);
xnor U12539 (N_12539,N_11451,N_11930);
xor U12540 (N_12540,N_11509,N_11522);
nand U12541 (N_12541,N_11926,N_11910);
and U12542 (N_12542,N_11662,N_11849);
nand U12543 (N_12543,N_11436,N_11923);
nor U12544 (N_12544,N_11593,N_11907);
or U12545 (N_12545,N_11727,N_11719);
nand U12546 (N_12546,N_11574,N_11765);
nor U12547 (N_12547,N_11832,N_11540);
or U12548 (N_12548,N_11660,N_11836);
or U12549 (N_12549,N_11802,N_11790);
xnor U12550 (N_12550,N_11639,N_11804);
and U12551 (N_12551,N_11742,N_11941);
nor U12552 (N_12552,N_11679,N_11767);
xor U12553 (N_12553,N_11557,N_11906);
nand U12554 (N_12554,N_11527,N_11782);
xnor U12555 (N_12555,N_11641,N_11621);
or U12556 (N_12556,N_11944,N_11439);
nor U12557 (N_12557,N_11631,N_11958);
nand U12558 (N_12558,N_11829,N_11591);
xor U12559 (N_12559,N_11467,N_11861);
and U12560 (N_12560,N_11806,N_11711);
xor U12561 (N_12561,N_11932,N_11954);
nor U12562 (N_12562,N_11897,N_11584);
and U12563 (N_12563,N_11768,N_11408);
nor U12564 (N_12564,N_11721,N_11690);
nand U12565 (N_12565,N_11614,N_11840);
nor U12566 (N_12566,N_11847,N_11992);
nand U12567 (N_12567,N_11631,N_11939);
or U12568 (N_12568,N_11912,N_11499);
nand U12569 (N_12569,N_11537,N_11579);
nand U12570 (N_12570,N_11783,N_11602);
nor U12571 (N_12571,N_11986,N_11837);
nand U12572 (N_12572,N_11679,N_11493);
nand U12573 (N_12573,N_11657,N_11407);
and U12574 (N_12574,N_11634,N_11941);
xnor U12575 (N_12575,N_11516,N_11560);
nand U12576 (N_12576,N_11974,N_11891);
and U12577 (N_12577,N_11542,N_11862);
nor U12578 (N_12578,N_11417,N_11548);
nor U12579 (N_12579,N_11704,N_11807);
or U12580 (N_12580,N_11874,N_11508);
nand U12581 (N_12581,N_11556,N_11863);
or U12582 (N_12582,N_11920,N_11901);
nand U12583 (N_12583,N_11626,N_11963);
nand U12584 (N_12584,N_11577,N_11513);
nand U12585 (N_12585,N_11773,N_11413);
or U12586 (N_12586,N_11841,N_11749);
nor U12587 (N_12587,N_11866,N_11609);
nand U12588 (N_12588,N_11990,N_11631);
nand U12589 (N_12589,N_11439,N_11626);
and U12590 (N_12590,N_11949,N_11845);
nor U12591 (N_12591,N_11629,N_11682);
or U12592 (N_12592,N_11466,N_11580);
nand U12593 (N_12593,N_11680,N_11718);
nand U12594 (N_12594,N_11477,N_11665);
or U12595 (N_12595,N_11413,N_11982);
nor U12596 (N_12596,N_11612,N_11580);
nor U12597 (N_12597,N_11619,N_11923);
xor U12598 (N_12598,N_11568,N_11910);
or U12599 (N_12599,N_11679,N_11428);
nand U12600 (N_12600,N_12289,N_12293);
or U12601 (N_12601,N_12000,N_12144);
xnor U12602 (N_12602,N_12128,N_12140);
or U12603 (N_12603,N_12409,N_12112);
nand U12604 (N_12604,N_12146,N_12416);
nor U12605 (N_12605,N_12545,N_12096);
nor U12606 (N_12606,N_12489,N_12386);
and U12607 (N_12607,N_12095,N_12257);
or U12608 (N_12608,N_12286,N_12404);
nor U12609 (N_12609,N_12408,N_12191);
or U12610 (N_12610,N_12371,N_12501);
nand U12611 (N_12611,N_12300,N_12283);
or U12612 (N_12612,N_12599,N_12256);
nand U12613 (N_12613,N_12124,N_12581);
nor U12614 (N_12614,N_12226,N_12249);
nor U12615 (N_12615,N_12434,N_12365);
and U12616 (N_12616,N_12524,N_12540);
nor U12617 (N_12617,N_12216,N_12041);
nand U12618 (N_12618,N_12102,N_12295);
or U12619 (N_12619,N_12573,N_12356);
xnor U12620 (N_12620,N_12443,N_12161);
xor U12621 (N_12621,N_12379,N_12267);
nand U12622 (N_12622,N_12305,N_12415);
and U12623 (N_12623,N_12506,N_12003);
nor U12624 (N_12624,N_12253,N_12264);
xnor U12625 (N_12625,N_12517,N_12413);
or U12626 (N_12626,N_12590,N_12263);
or U12627 (N_12627,N_12014,N_12232);
nand U12628 (N_12628,N_12131,N_12437);
and U12629 (N_12629,N_12205,N_12534);
and U12630 (N_12630,N_12453,N_12511);
nand U12631 (N_12631,N_12587,N_12569);
nand U12632 (N_12632,N_12065,N_12188);
xor U12633 (N_12633,N_12322,N_12036);
nand U12634 (N_12634,N_12233,N_12550);
and U12635 (N_12635,N_12548,N_12575);
xnor U12636 (N_12636,N_12173,N_12001);
nand U12637 (N_12637,N_12557,N_12228);
nand U12638 (N_12638,N_12230,N_12049);
xor U12639 (N_12639,N_12297,N_12209);
and U12640 (N_12640,N_12510,N_12227);
and U12641 (N_12641,N_12478,N_12598);
or U12642 (N_12642,N_12442,N_12594);
nand U12643 (N_12643,N_12178,N_12225);
nand U12644 (N_12644,N_12179,N_12250);
nor U12645 (N_12645,N_12298,N_12502);
nor U12646 (N_12646,N_12083,N_12183);
or U12647 (N_12647,N_12072,N_12012);
nor U12648 (N_12648,N_12113,N_12348);
xnor U12649 (N_12649,N_12077,N_12269);
nand U12650 (N_12650,N_12398,N_12156);
nor U12651 (N_12651,N_12115,N_12231);
and U12652 (N_12652,N_12568,N_12022);
nor U12653 (N_12653,N_12053,N_12523);
nor U12654 (N_12654,N_12536,N_12314);
nand U12655 (N_12655,N_12270,N_12273);
or U12656 (N_12656,N_12303,N_12337);
and U12657 (N_12657,N_12125,N_12410);
xnor U12658 (N_12658,N_12215,N_12375);
xnor U12659 (N_12659,N_12139,N_12084);
xnor U12660 (N_12660,N_12588,N_12308);
nor U12661 (N_12661,N_12358,N_12397);
or U12662 (N_12662,N_12496,N_12255);
or U12663 (N_12663,N_12234,N_12004);
xnor U12664 (N_12664,N_12103,N_12584);
xnor U12665 (N_12665,N_12060,N_12187);
nand U12666 (N_12666,N_12069,N_12207);
nand U12667 (N_12667,N_12252,N_12494);
nor U12668 (N_12668,N_12302,N_12352);
and U12669 (N_12669,N_12285,N_12407);
xnor U12670 (N_12670,N_12324,N_12164);
xnor U12671 (N_12671,N_12556,N_12149);
xnor U12672 (N_12672,N_12222,N_12242);
nand U12673 (N_12673,N_12132,N_12313);
xnor U12674 (N_12674,N_12197,N_12471);
nand U12675 (N_12675,N_12312,N_12218);
xor U12676 (N_12676,N_12591,N_12417);
and U12677 (N_12677,N_12533,N_12021);
or U12678 (N_12678,N_12210,N_12479);
nand U12679 (N_12679,N_12247,N_12214);
or U12680 (N_12680,N_12349,N_12526);
xor U12681 (N_12681,N_12520,N_12108);
and U12682 (N_12682,N_12359,N_12284);
nand U12683 (N_12683,N_12374,N_12236);
nand U12684 (N_12684,N_12428,N_12217);
nand U12685 (N_12685,N_12528,N_12384);
xor U12686 (N_12686,N_12552,N_12169);
xnor U12687 (N_12687,N_12450,N_12487);
xnor U12688 (N_12688,N_12159,N_12400);
and U12689 (N_12689,N_12596,N_12266);
nor U12690 (N_12690,N_12529,N_12332);
xor U12691 (N_12691,N_12045,N_12445);
or U12692 (N_12692,N_12372,N_12185);
and U12693 (N_12693,N_12032,N_12454);
xnor U12694 (N_12694,N_12050,N_12476);
and U12695 (N_12695,N_12422,N_12492);
or U12696 (N_12696,N_12504,N_12565);
xor U12697 (N_12697,N_12048,N_12505);
xor U12698 (N_12698,N_12465,N_12425);
and U12699 (N_12699,N_12200,N_12251);
or U12700 (N_12700,N_12190,N_12551);
and U12701 (N_12701,N_12593,N_12116);
xor U12702 (N_12702,N_12148,N_12490);
and U12703 (N_12703,N_12011,N_12497);
nand U12704 (N_12704,N_12175,N_12165);
nand U12705 (N_12705,N_12583,N_12005);
xor U12706 (N_12706,N_12491,N_12194);
nand U12707 (N_12707,N_12274,N_12061);
nor U12708 (N_12708,N_12448,N_12294);
nand U12709 (N_12709,N_12424,N_12592);
xor U12710 (N_12710,N_12589,N_12340);
xor U12711 (N_12711,N_12137,N_12064);
and U12712 (N_12712,N_12162,N_12595);
or U12713 (N_12713,N_12157,N_12109);
or U12714 (N_12714,N_12019,N_12553);
or U12715 (N_12715,N_12527,N_12241);
xor U12716 (N_12716,N_12304,N_12062);
xor U12717 (N_12717,N_12068,N_12512);
or U12718 (N_12718,N_12576,N_12421);
xnor U12719 (N_12719,N_12343,N_12086);
nor U12720 (N_12720,N_12515,N_12387);
or U12721 (N_12721,N_12299,N_12480);
xor U12722 (N_12722,N_12118,N_12455);
and U12723 (N_12723,N_12406,N_12531);
nor U12724 (N_12724,N_12571,N_12432);
nor U12725 (N_12725,N_12276,N_12029);
nor U12726 (N_12726,N_12093,N_12335);
nand U12727 (N_12727,N_12484,N_12025);
xor U12728 (N_12728,N_12017,N_12244);
and U12729 (N_12729,N_12182,N_12493);
or U12730 (N_12730,N_12213,N_12160);
nor U12731 (N_12731,N_12559,N_12399);
or U12732 (N_12732,N_12315,N_12122);
xor U12733 (N_12733,N_12039,N_12477);
nand U12734 (N_12734,N_12013,N_12525);
nand U12735 (N_12735,N_12354,N_12059);
xor U12736 (N_12736,N_12151,N_12171);
and U12737 (N_12737,N_12223,N_12212);
nand U12738 (N_12738,N_12024,N_12291);
nand U12739 (N_12739,N_12063,N_12586);
and U12740 (N_12740,N_12296,N_12431);
xnor U12741 (N_12741,N_12488,N_12037);
or U12742 (N_12742,N_12046,N_12288);
xor U12743 (N_12743,N_12094,N_12272);
nand U12744 (N_12744,N_12089,N_12259);
or U12745 (N_12745,N_12154,N_12562);
xor U12746 (N_12746,N_12206,N_12034);
nor U12747 (N_12747,N_12150,N_12073);
or U12748 (N_12748,N_12378,N_12180);
or U12749 (N_12749,N_12172,N_12135);
nor U12750 (N_12750,N_12100,N_12458);
nor U12751 (N_12751,N_12403,N_12129);
xor U12752 (N_12752,N_12339,N_12261);
nand U12753 (N_12753,N_12051,N_12331);
nand U12754 (N_12754,N_12088,N_12486);
or U12755 (N_12755,N_12360,N_12040);
xor U12756 (N_12756,N_12447,N_12396);
xor U12757 (N_12757,N_12016,N_12363);
nand U12758 (N_12758,N_12370,N_12317);
xor U12759 (N_12759,N_12390,N_12186);
or U12760 (N_12760,N_12380,N_12008);
and U12761 (N_12761,N_12326,N_12027);
or U12762 (N_12762,N_12546,N_12473);
nor U12763 (N_12763,N_12555,N_12208);
nand U12764 (N_12764,N_12333,N_12262);
xnor U12765 (N_12765,N_12318,N_12467);
nor U12766 (N_12766,N_12136,N_12463);
xor U12767 (N_12767,N_12071,N_12015);
nand U12768 (N_12768,N_12074,N_12110);
nand U12769 (N_12769,N_12133,N_12518);
nand U12770 (N_12770,N_12177,N_12203);
nand U12771 (N_12771,N_12010,N_12464);
nand U12772 (N_12772,N_12521,N_12138);
nand U12773 (N_12773,N_12355,N_12107);
nor U12774 (N_12774,N_12007,N_12485);
or U12775 (N_12775,N_12221,N_12147);
xnor U12776 (N_12776,N_12204,N_12460);
or U12777 (N_12777,N_12412,N_12211);
or U12778 (N_12778,N_12101,N_12309);
and U12779 (N_12779,N_12023,N_12566);
nand U12780 (N_12780,N_12405,N_12042);
and U12781 (N_12781,N_12092,N_12143);
and U12782 (N_12782,N_12351,N_12321);
and U12783 (N_12783,N_12306,N_12522);
xnor U12784 (N_12784,N_12342,N_12394);
or U12785 (N_12785,N_12373,N_12430);
nand U12786 (N_12786,N_12067,N_12325);
or U12787 (N_12787,N_12368,N_12411);
nand U12788 (N_12788,N_12574,N_12376);
or U12789 (N_12789,N_12224,N_12009);
xor U12790 (N_12790,N_12597,N_12091);
or U12791 (N_12791,N_12457,N_12462);
xnor U12792 (N_12792,N_12153,N_12483);
nor U12793 (N_12793,N_12393,N_12275);
or U12794 (N_12794,N_12130,N_12155);
or U12795 (N_12795,N_12449,N_12475);
and U12796 (N_12796,N_12176,N_12539);
nand U12797 (N_12797,N_12106,N_12391);
xor U12798 (N_12798,N_12420,N_12466);
or U12799 (N_12799,N_12423,N_12035);
and U12800 (N_12800,N_12530,N_12280);
xnor U12801 (N_12801,N_12082,N_12345);
or U12802 (N_12802,N_12469,N_12446);
xor U12803 (N_12803,N_12361,N_12018);
or U12804 (N_12804,N_12134,N_12195);
nand U12805 (N_12805,N_12006,N_12141);
nor U12806 (N_12806,N_12452,N_12369);
nor U12807 (N_12807,N_12117,N_12382);
nor U12808 (N_12808,N_12114,N_12519);
nand U12809 (N_12809,N_12508,N_12367);
and U12810 (N_12810,N_12543,N_12381);
nand U12811 (N_12811,N_12444,N_12500);
and U12812 (N_12812,N_12126,N_12170);
xnor U12813 (N_12813,N_12240,N_12085);
or U12814 (N_12814,N_12099,N_12090);
and U12815 (N_12815,N_12075,N_12585);
and U12816 (N_12816,N_12258,N_12026);
or U12817 (N_12817,N_12336,N_12254);
xnor U12818 (N_12818,N_12438,N_12043);
nor U12819 (N_12819,N_12353,N_12563);
or U12820 (N_12820,N_12123,N_12327);
or U12821 (N_12821,N_12119,N_12513);
xor U12822 (N_12822,N_12330,N_12028);
nand U12823 (N_12823,N_12181,N_12436);
and U12824 (N_12824,N_12451,N_12357);
or U12825 (N_12825,N_12482,N_12329);
and U12826 (N_12826,N_12544,N_12532);
and U12827 (N_12827,N_12271,N_12199);
nand U12828 (N_12828,N_12377,N_12057);
and U12829 (N_12829,N_12033,N_12503);
or U12830 (N_12830,N_12579,N_12547);
or U12831 (N_12831,N_12395,N_12310);
nand U12832 (N_12832,N_12388,N_12166);
xor U12833 (N_12833,N_12142,N_12538);
nand U12834 (N_12834,N_12426,N_12401);
and U12835 (N_12835,N_12248,N_12468);
or U12836 (N_12836,N_12564,N_12362);
xnor U12837 (N_12837,N_12239,N_12196);
nor U12838 (N_12838,N_12121,N_12030);
or U12839 (N_12839,N_12439,N_12389);
and U12840 (N_12840,N_12435,N_12441);
xor U12841 (N_12841,N_12198,N_12334);
or U12842 (N_12842,N_12054,N_12038);
and U12843 (N_12843,N_12056,N_12418);
nor U12844 (N_12844,N_12385,N_12268);
and U12845 (N_12845,N_12344,N_12078);
or U12846 (N_12846,N_12316,N_12572);
nand U12847 (N_12847,N_12350,N_12070);
nand U12848 (N_12848,N_12235,N_12535);
and U12849 (N_12849,N_12507,N_12537);
and U12850 (N_12850,N_12509,N_12481);
xor U12851 (N_12851,N_12260,N_12158);
nand U12852 (N_12852,N_12002,N_12097);
and U12853 (N_12853,N_12320,N_12301);
nor U12854 (N_12854,N_12052,N_12429);
or U12855 (N_12855,N_12338,N_12541);
nor U12856 (N_12856,N_12163,N_12328);
nand U12857 (N_12857,N_12554,N_12347);
or U12858 (N_12858,N_12495,N_12414);
nor U12859 (N_12859,N_12582,N_12229);
nand U12860 (N_12860,N_12577,N_12307);
and U12861 (N_12861,N_12364,N_12145);
nor U12862 (N_12862,N_12174,N_12542);
nand U12863 (N_12863,N_12219,N_12402);
nand U12864 (N_12864,N_12047,N_12104);
and U12865 (N_12865,N_12168,N_12238);
and U12866 (N_12866,N_12567,N_12201);
nand U12867 (N_12867,N_12580,N_12120);
and U12868 (N_12868,N_12277,N_12433);
nor U12869 (N_12869,N_12281,N_12079);
nand U12870 (N_12870,N_12514,N_12311);
or U12871 (N_12871,N_12127,N_12055);
nand U12872 (N_12872,N_12184,N_12472);
nor U12873 (N_12873,N_12570,N_12558);
nand U12874 (N_12874,N_12189,N_12578);
nand U12875 (N_12875,N_12323,N_12098);
or U12876 (N_12876,N_12044,N_12243);
nor U12877 (N_12877,N_12498,N_12341);
and U12878 (N_12878,N_12427,N_12105);
nand U12879 (N_12879,N_12237,N_12058);
nor U12880 (N_12880,N_12392,N_12474);
xnor U12881 (N_12881,N_12080,N_12076);
xnor U12882 (N_12882,N_12346,N_12282);
xor U12883 (N_12883,N_12549,N_12383);
nor U12884 (N_12884,N_12246,N_12292);
or U12885 (N_12885,N_12470,N_12278);
nand U12886 (N_12886,N_12192,N_12066);
nand U12887 (N_12887,N_12081,N_12319);
xor U12888 (N_12888,N_12440,N_12087);
nor U12889 (N_12889,N_12167,N_12031);
or U12890 (N_12890,N_12265,N_12560);
or U12891 (N_12891,N_12499,N_12020);
nand U12892 (N_12892,N_12459,N_12193);
nor U12893 (N_12893,N_12461,N_12220);
nand U12894 (N_12894,N_12456,N_12111);
nand U12895 (N_12895,N_12152,N_12245);
or U12896 (N_12896,N_12290,N_12516);
and U12897 (N_12897,N_12366,N_12279);
xnor U12898 (N_12898,N_12419,N_12561);
nor U12899 (N_12899,N_12202,N_12287);
nand U12900 (N_12900,N_12545,N_12568);
nor U12901 (N_12901,N_12275,N_12572);
nand U12902 (N_12902,N_12109,N_12048);
or U12903 (N_12903,N_12492,N_12311);
nand U12904 (N_12904,N_12093,N_12477);
xnor U12905 (N_12905,N_12285,N_12372);
xor U12906 (N_12906,N_12017,N_12039);
and U12907 (N_12907,N_12052,N_12501);
and U12908 (N_12908,N_12577,N_12540);
or U12909 (N_12909,N_12353,N_12541);
or U12910 (N_12910,N_12515,N_12283);
nand U12911 (N_12911,N_12373,N_12277);
xor U12912 (N_12912,N_12529,N_12271);
and U12913 (N_12913,N_12341,N_12485);
nand U12914 (N_12914,N_12231,N_12101);
and U12915 (N_12915,N_12076,N_12485);
or U12916 (N_12916,N_12079,N_12539);
nand U12917 (N_12917,N_12442,N_12014);
nor U12918 (N_12918,N_12193,N_12321);
and U12919 (N_12919,N_12172,N_12463);
and U12920 (N_12920,N_12477,N_12218);
xor U12921 (N_12921,N_12489,N_12490);
nor U12922 (N_12922,N_12446,N_12397);
and U12923 (N_12923,N_12559,N_12468);
nand U12924 (N_12924,N_12379,N_12056);
xnor U12925 (N_12925,N_12386,N_12596);
nand U12926 (N_12926,N_12045,N_12303);
xnor U12927 (N_12927,N_12549,N_12195);
xnor U12928 (N_12928,N_12051,N_12088);
nand U12929 (N_12929,N_12486,N_12084);
or U12930 (N_12930,N_12366,N_12196);
nor U12931 (N_12931,N_12561,N_12568);
or U12932 (N_12932,N_12106,N_12157);
xor U12933 (N_12933,N_12178,N_12528);
nand U12934 (N_12934,N_12369,N_12394);
and U12935 (N_12935,N_12103,N_12348);
xnor U12936 (N_12936,N_12336,N_12549);
nand U12937 (N_12937,N_12454,N_12236);
xnor U12938 (N_12938,N_12413,N_12479);
nor U12939 (N_12939,N_12357,N_12253);
nor U12940 (N_12940,N_12597,N_12219);
nor U12941 (N_12941,N_12361,N_12266);
nor U12942 (N_12942,N_12277,N_12166);
xnor U12943 (N_12943,N_12494,N_12316);
nor U12944 (N_12944,N_12307,N_12237);
and U12945 (N_12945,N_12569,N_12340);
nand U12946 (N_12946,N_12517,N_12143);
xor U12947 (N_12947,N_12392,N_12530);
and U12948 (N_12948,N_12177,N_12586);
xor U12949 (N_12949,N_12534,N_12562);
nand U12950 (N_12950,N_12492,N_12441);
xnor U12951 (N_12951,N_12557,N_12424);
and U12952 (N_12952,N_12134,N_12502);
nor U12953 (N_12953,N_12403,N_12574);
nand U12954 (N_12954,N_12027,N_12464);
and U12955 (N_12955,N_12476,N_12254);
or U12956 (N_12956,N_12189,N_12389);
or U12957 (N_12957,N_12183,N_12511);
nor U12958 (N_12958,N_12027,N_12286);
nor U12959 (N_12959,N_12457,N_12301);
and U12960 (N_12960,N_12566,N_12398);
nor U12961 (N_12961,N_12347,N_12352);
and U12962 (N_12962,N_12323,N_12540);
and U12963 (N_12963,N_12264,N_12588);
nand U12964 (N_12964,N_12347,N_12202);
nand U12965 (N_12965,N_12503,N_12485);
or U12966 (N_12966,N_12012,N_12003);
or U12967 (N_12967,N_12154,N_12519);
or U12968 (N_12968,N_12063,N_12490);
nor U12969 (N_12969,N_12253,N_12193);
nor U12970 (N_12970,N_12317,N_12103);
or U12971 (N_12971,N_12022,N_12322);
and U12972 (N_12972,N_12574,N_12375);
nand U12973 (N_12973,N_12373,N_12179);
nand U12974 (N_12974,N_12082,N_12052);
nor U12975 (N_12975,N_12162,N_12044);
nand U12976 (N_12976,N_12004,N_12113);
nor U12977 (N_12977,N_12484,N_12358);
nand U12978 (N_12978,N_12100,N_12076);
nand U12979 (N_12979,N_12547,N_12274);
nand U12980 (N_12980,N_12402,N_12146);
xnor U12981 (N_12981,N_12574,N_12517);
xnor U12982 (N_12982,N_12156,N_12128);
xor U12983 (N_12983,N_12552,N_12326);
and U12984 (N_12984,N_12403,N_12444);
or U12985 (N_12985,N_12165,N_12570);
xor U12986 (N_12986,N_12030,N_12411);
and U12987 (N_12987,N_12464,N_12533);
nand U12988 (N_12988,N_12573,N_12346);
nand U12989 (N_12989,N_12153,N_12468);
nand U12990 (N_12990,N_12390,N_12191);
xor U12991 (N_12991,N_12206,N_12211);
and U12992 (N_12992,N_12446,N_12502);
xor U12993 (N_12993,N_12017,N_12446);
nand U12994 (N_12994,N_12531,N_12079);
xor U12995 (N_12995,N_12432,N_12536);
nor U12996 (N_12996,N_12052,N_12482);
nand U12997 (N_12997,N_12510,N_12477);
or U12998 (N_12998,N_12183,N_12412);
and U12999 (N_12999,N_12213,N_12183);
and U13000 (N_13000,N_12137,N_12063);
nand U13001 (N_13001,N_12424,N_12076);
xor U13002 (N_13002,N_12430,N_12447);
and U13003 (N_13003,N_12538,N_12099);
xnor U13004 (N_13004,N_12349,N_12056);
nand U13005 (N_13005,N_12156,N_12203);
or U13006 (N_13006,N_12060,N_12547);
nand U13007 (N_13007,N_12365,N_12469);
or U13008 (N_13008,N_12056,N_12495);
nand U13009 (N_13009,N_12345,N_12286);
xnor U13010 (N_13010,N_12014,N_12195);
nand U13011 (N_13011,N_12361,N_12033);
nand U13012 (N_13012,N_12364,N_12570);
nand U13013 (N_13013,N_12109,N_12091);
nor U13014 (N_13014,N_12382,N_12221);
nand U13015 (N_13015,N_12203,N_12314);
nand U13016 (N_13016,N_12578,N_12452);
or U13017 (N_13017,N_12501,N_12209);
xnor U13018 (N_13018,N_12210,N_12016);
and U13019 (N_13019,N_12349,N_12454);
nand U13020 (N_13020,N_12136,N_12303);
or U13021 (N_13021,N_12243,N_12335);
xnor U13022 (N_13022,N_12308,N_12584);
xnor U13023 (N_13023,N_12433,N_12270);
nor U13024 (N_13024,N_12284,N_12407);
and U13025 (N_13025,N_12323,N_12531);
or U13026 (N_13026,N_12485,N_12448);
or U13027 (N_13027,N_12151,N_12271);
nor U13028 (N_13028,N_12553,N_12219);
nor U13029 (N_13029,N_12349,N_12479);
or U13030 (N_13030,N_12093,N_12323);
and U13031 (N_13031,N_12563,N_12438);
or U13032 (N_13032,N_12121,N_12098);
xnor U13033 (N_13033,N_12540,N_12532);
or U13034 (N_13034,N_12137,N_12148);
nor U13035 (N_13035,N_12234,N_12485);
nand U13036 (N_13036,N_12455,N_12576);
nor U13037 (N_13037,N_12493,N_12041);
and U13038 (N_13038,N_12314,N_12337);
and U13039 (N_13039,N_12526,N_12515);
and U13040 (N_13040,N_12481,N_12175);
and U13041 (N_13041,N_12138,N_12440);
nor U13042 (N_13042,N_12039,N_12178);
nand U13043 (N_13043,N_12169,N_12210);
or U13044 (N_13044,N_12137,N_12383);
nand U13045 (N_13045,N_12596,N_12427);
xor U13046 (N_13046,N_12356,N_12037);
nor U13047 (N_13047,N_12178,N_12515);
xnor U13048 (N_13048,N_12188,N_12240);
and U13049 (N_13049,N_12415,N_12587);
and U13050 (N_13050,N_12566,N_12505);
nor U13051 (N_13051,N_12298,N_12294);
nor U13052 (N_13052,N_12559,N_12180);
nor U13053 (N_13053,N_12425,N_12428);
nor U13054 (N_13054,N_12387,N_12554);
nor U13055 (N_13055,N_12583,N_12528);
and U13056 (N_13056,N_12597,N_12176);
or U13057 (N_13057,N_12136,N_12204);
and U13058 (N_13058,N_12035,N_12473);
or U13059 (N_13059,N_12297,N_12457);
nor U13060 (N_13060,N_12522,N_12594);
and U13061 (N_13061,N_12027,N_12541);
nor U13062 (N_13062,N_12446,N_12323);
nor U13063 (N_13063,N_12036,N_12471);
or U13064 (N_13064,N_12208,N_12387);
and U13065 (N_13065,N_12583,N_12288);
nand U13066 (N_13066,N_12231,N_12133);
nand U13067 (N_13067,N_12290,N_12386);
xor U13068 (N_13068,N_12339,N_12395);
nor U13069 (N_13069,N_12464,N_12426);
xor U13070 (N_13070,N_12218,N_12068);
nor U13071 (N_13071,N_12570,N_12124);
and U13072 (N_13072,N_12551,N_12126);
xnor U13073 (N_13073,N_12198,N_12219);
or U13074 (N_13074,N_12199,N_12459);
nand U13075 (N_13075,N_12151,N_12325);
and U13076 (N_13076,N_12543,N_12436);
xnor U13077 (N_13077,N_12598,N_12104);
and U13078 (N_13078,N_12365,N_12517);
nor U13079 (N_13079,N_12273,N_12539);
xnor U13080 (N_13080,N_12473,N_12028);
or U13081 (N_13081,N_12567,N_12146);
nand U13082 (N_13082,N_12295,N_12410);
nand U13083 (N_13083,N_12210,N_12507);
or U13084 (N_13084,N_12104,N_12464);
nor U13085 (N_13085,N_12430,N_12344);
or U13086 (N_13086,N_12562,N_12539);
nand U13087 (N_13087,N_12277,N_12464);
or U13088 (N_13088,N_12391,N_12053);
nand U13089 (N_13089,N_12411,N_12393);
and U13090 (N_13090,N_12433,N_12473);
and U13091 (N_13091,N_12579,N_12472);
nor U13092 (N_13092,N_12032,N_12068);
and U13093 (N_13093,N_12388,N_12422);
and U13094 (N_13094,N_12561,N_12032);
xor U13095 (N_13095,N_12373,N_12240);
nor U13096 (N_13096,N_12383,N_12392);
nor U13097 (N_13097,N_12302,N_12057);
nand U13098 (N_13098,N_12402,N_12424);
nor U13099 (N_13099,N_12357,N_12039);
or U13100 (N_13100,N_12199,N_12140);
nand U13101 (N_13101,N_12519,N_12479);
or U13102 (N_13102,N_12148,N_12525);
and U13103 (N_13103,N_12500,N_12306);
or U13104 (N_13104,N_12267,N_12031);
and U13105 (N_13105,N_12190,N_12482);
xnor U13106 (N_13106,N_12466,N_12159);
nor U13107 (N_13107,N_12134,N_12548);
and U13108 (N_13108,N_12532,N_12071);
nor U13109 (N_13109,N_12335,N_12119);
nand U13110 (N_13110,N_12225,N_12274);
nand U13111 (N_13111,N_12507,N_12079);
nand U13112 (N_13112,N_12262,N_12533);
and U13113 (N_13113,N_12291,N_12486);
nand U13114 (N_13114,N_12257,N_12319);
and U13115 (N_13115,N_12136,N_12231);
or U13116 (N_13116,N_12226,N_12443);
nor U13117 (N_13117,N_12390,N_12215);
and U13118 (N_13118,N_12066,N_12096);
nand U13119 (N_13119,N_12287,N_12551);
xor U13120 (N_13120,N_12057,N_12030);
nor U13121 (N_13121,N_12519,N_12021);
nor U13122 (N_13122,N_12217,N_12002);
nor U13123 (N_13123,N_12058,N_12416);
or U13124 (N_13124,N_12450,N_12341);
xor U13125 (N_13125,N_12241,N_12011);
xnor U13126 (N_13126,N_12393,N_12273);
and U13127 (N_13127,N_12088,N_12054);
xnor U13128 (N_13128,N_12358,N_12565);
or U13129 (N_13129,N_12133,N_12229);
nand U13130 (N_13130,N_12119,N_12416);
nand U13131 (N_13131,N_12012,N_12455);
nor U13132 (N_13132,N_12267,N_12089);
nand U13133 (N_13133,N_12025,N_12046);
xnor U13134 (N_13134,N_12315,N_12489);
nor U13135 (N_13135,N_12221,N_12550);
nor U13136 (N_13136,N_12363,N_12462);
nor U13137 (N_13137,N_12165,N_12076);
xor U13138 (N_13138,N_12475,N_12329);
xnor U13139 (N_13139,N_12078,N_12201);
nand U13140 (N_13140,N_12027,N_12457);
nor U13141 (N_13141,N_12075,N_12123);
xnor U13142 (N_13142,N_12446,N_12233);
or U13143 (N_13143,N_12403,N_12061);
nand U13144 (N_13144,N_12121,N_12223);
nor U13145 (N_13145,N_12388,N_12172);
xor U13146 (N_13146,N_12590,N_12034);
or U13147 (N_13147,N_12261,N_12569);
xor U13148 (N_13148,N_12087,N_12494);
nand U13149 (N_13149,N_12431,N_12061);
and U13150 (N_13150,N_12559,N_12487);
or U13151 (N_13151,N_12356,N_12286);
xnor U13152 (N_13152,N_12410,N_12423);
nor U13153 (N_13153,N_12011,N_12587);
and U13154 (N_13154,N_12393,N_12414);
and U13155 (N_13155,N_12415,N_12206);
nand U13156 (N_13156,N_12172,N_12309);
or U13157 (N_13157,N_12434,N_12171);
or U13158 (N_13158,N_12105,N_12520);
and U13159 (N_13159,N_12461,N_12355);
or U13160 (N_13160,N_12544,N_12190);
and U13161 (N_13161,N_12548,N_12159);
nand U13162 (N_13162,N_12340,N_12125);
xor U13163 (N_13163,N_12119,N_12372);
xor U13164 (N_13164,N_12494,N_12204);
or U13165 (N_13165,N_12472,N_12037);
nand U13166 (N_13166,N_12240,N_12325);
nand U13167 (N_13167,N_12052,N_12130);
xnor U13168 (N_13168,N_12471,N_12323);
or U13169 (N_13169,N_12395,N_12316);
nor U13170 (N_13170,N_12182,N_12029);
nand U13171 (N_13171,N_12166,N_12141);
and U13172 (N_13172,N_12097,N_12141);
xor U13173 (N_13173,N_12342,N_12415);
nor U13174 (N_13174,N_12320,N_12050);
or U13175 (N_13175,N_12206,N_12586);
and U13176 (N_13176,N_12462,N_12250);
nand U13177 (N_13177,N_12010,N_12366);
xor U13178 (N_13178,N_12375,N_12049);
or U13179 (N_13179,N_12286,N_12265);
xnor U13180 (N_13180,N_12139,N_12105);
xor U13181 (N_13181,N_12082,N_12105);
or U13182 (N_13182,N_12054,N_12123);
xor U13183 (N_13183,N_12204,N_12172);
or U13184 (N_13184,N_12215,N_12196);
and U13185 (N_13185,N_12107,N_12559);
nor U13186 (N_13186,N_12007,N_12427);
nand U13187 (N_13187,N_12371,N_12251);
nand U13188 (N_13188,N_12091,N_12585);
nor U13189 (N_13189,N_12222,N_12382);
or U13190 (N_13190,N_12054,N_12242);
and U13191 (N_13191,N_12453,N_12374);
nor U13192 (N_13192,N_12515,N_12579);
xor U13193 (N_13193,N_12405,N_12415);
nand U13194 (N_13194,N_12014,N_12174);
and U13195 (N_13195,N_12147,N_12059);
nand U13196 (N_13196,N_12445,N_12334);
nand U13197 (N_13197,N_12131,N_12111);
nand U13198 (N_13198,N_12504,N_12329);
nand U13199 (N_13199,N_12394,N_12490);
and U13200 (N_13200,N_13070,N_12705);
nand U13201 (N_13201,N_13041,N_12939);
and U13202 (N_13202,N_12855,N_13119);
and U13203 (N_13203,N_13181,N_12791);
nand U13204 (N_13204,N_13034,N_12806);
nand U13205 (N_13205,N_13071,N_13003);
xnor U13206 (N_13206,N_12815,N_12671);
or U13207 (N_13207,N_13144,N_12695);
and U13208 (N_13208,N_13199,N_12865);
nand U13209 (N_13209,N_12676,N_13150);
xor U13210 (N_13210,N_13006,N_13079);
xor U13211 (N_13211,N_12763,N_12930);
xnor U13212 (N_13212,N_12947,N_12692);
nor U13213 (N_13213,N_12785,N_13058);
xor U13214 (N_13214,N_13149,N_12708);
nand U13215 (N_13215,N_12822,N_13147);
nor U13216 (N_13216,N_12679,N_12683);
nand U13217 (N_13217,N_12736,N_12782);
or U13218 (N_13218,N_12819,N_12739);
and U13219 (N_13219,N_12602,N_13033);
and U13220 (N_13220,N_12788,N_12843);
nor U13221 (N_13221,N_12711,N_12801);
xor U13222 (N_13222,N_13010,N_12633);
and U13223 (N_13223,N_12710,N_13187);
nand U13224 (N_13224,N_12900,N_13168);
nand U13225 (N_13225,N_12878,N_12720);
nor U13226 (N_13226,N_13103,N_13108);
nor U13227 (N_13227,N_12625,N_12970);
nand U13228 (N_13228,N_12818,N_12870);
nor U13229 (N_13229,N_12767,N_12831);
or U13230 (N_13230,N_12879,N_12697);
and U13231 (N_13231,N_13189,N_12847);
xnor U13232 (N_13232,N_12761,N_12848);
or U13233 (N_13233,N_12615,N_12858);
xnor U13234 (N_13234,N_12724,N_12936);
xor U13235 (N_13235,N_12910,N_12614);
xor U13236 (N_13236,N_12616,N_12744);
nor U13237 (N_13237,N_12877,N_12601);
xnor U13238 (N_13238,N_12902,N_12707);
xnor U13239 (N_13239,N_13184,N_12639);
nand U13240 (N_13240,N_12700,N_12773);
and U13241 (N_13241,N_12712,N_13061);
or U13242 (N_13242,N_12716,N_13123);
and U13243 (N_13243,N_12898,N_12781);
or U13244 (N_13244,N_13073,N_13094);
xor U13245 (N_13245,N_12840,N_13105);
and U13246 (N_13246,N_12893,N_13170);
nand U13247 (N_13247,N_13171,N_13169);
nand U13248 (N_13248,N_12845,N_12757);
or U13249 (N_13249,N_12820,N_12914);
nor U13250 (N_13250,N_12717,N_12830);
nor U13251 (N_13251,N_12826,N_13101);
nor U13252 (N_13252,N_12926,N_12668);
nand U13253 (N_13253,N_12979,N_12608);
or U13254 (N_13254,N_12742,N_12938);
or U13255 (N_13255,N_12917,N_12886);
nor U13256 (N_13256,N_13057,N_12950);
xnor U13257 (N_13257,N_12646,N_12854);
and U13258 (N_13258,N_12637,N_13065);
and U13259 (N_13259,N_13087,N_12941);
nor U13260 (N_13260,N_13011,N_12632);
nand U13261 (N_13261,N_13091,N_13126);
or U13262 (N_13262,N_13163,N_13116);
nand U13263 (N_13263,N_12703,N_12772);
xnor U13264 (N_13264,N_12948,N_13114);
or U13265 (N_13265,N_13054,N_12940);
and U13266 (N_13266,N_13083,N_12783);
nand U13267 (N_13267,N_12644,N_12732);
or U13268 (N_13268,N_13014,N_12678);
nor U13269 (N_13269,N_12715,N_12817);
nand U13270 (N_13270,N_13066,N_12799);
nand U13271 (N_13271,N_12786,N_12984);
nor U13272 (N_13272,N_12856,N_12748);
nand U13273 (N_13273,N_12814,N_13102);
nand U13274 (N_13274,N_12857,N_12895);
xor U13275 (N_13275,N_12889,N_12699);
nor U13276 (N_13276,N_13148,N_12816);
nor U13277 (N_13277,N_12999,N_12760);
and U13278 (N_13278,N_12828,N_12961);
nor U13279 (N_13279,N_13172,N_12698);
and U13280 (N_13280,N_13160,N_12641);
or U13281 (N_13281,N_13132,N_13182);
nor U13282 (N_13282,N_12951,N_12643);
nand U13283 (N_13283,N_12628,N_12962);
and U13284 (N_13284,N_12880,N_12737);
and U13285 (N_13285,N_12796,N_13155);
xnor U13286 (N_13286,N_12829,N_12718);
and U13287 (N_13287,N_13064,N_12827);
nor U13288 (N_13288,N_12906,N_12762);
and U13289 (N_13289,N_13053,N_13027);
nor U13290 (N_13290,N_12967,N_12738);
nand U13291 (N_13291,N_12993,N_12807);
and U13292 (N_13292,N_12648,N_13085);
nand U13293 (N_13293,N_12627,N_12797);
xnor U13294 (N_13294,N_13096,N_12873);
nand U13295 (N_13295,N_12907,N_12811);
and U13296 (N_13296,N_12666,N_13137);
or U13297 (N_13297,N_12975,N_13019);
nand U13298 (N_13298,N_13020,N_13048);
nor U13299 (N_13299,N_12713,N_12623);
xnor U13300 (N_13300,N_12795,N_12645);
nand U13301 (N_13301,N_12909,N_13186);
and U13302 (N_13302,N_13042,N_12934);
and U13303 (N_13303,N_13175,N_12986);
nor U13304 (N_13304,N_13156,N_12613);
nand U13305 (N_13305,N_12618,N_12860);
xor U13306 (N_13306,N_13129,N_13145);
xor U13307 (N_13307,N_13029,N_12777);
and U13308 (N_13308,N_12721,N_13177);
nand U13309 (N_13309,N_12755,N_12964);
nor U13310 (N_13310,N_12851,N_12751);
nor U13311 (N_13311,N_12853,N_13174);
xor U13312 (N_13312,N_13060,N_13072);
or U13313 (N_13313,N_13043,N_12656);
and U13314 (N_13314,N_12978,N_12885);
nor U13315 (N_13315,N_12918,N_13035);
nand U13316 (N_13316,N_12802,N_12965);
xor U13317 (N_13317,N_12887,N_12908);
and U13318 (N_13318,N_13161,N_13122);
xor U13319 (N_13319,N_13075,N_12876);
nor U13320 (N_13320,N_13024,N_12912);
nand U13321 (N_13321,N_12691,N_12904);
and U13322 (N_13322,N_12704,N_12957);
and U13323 (N_13323,N_13179,N_12884);
or U13324 (N_13324,N_12674,N_12680);
nor U13325 (N_13325,N_12774,N_13153);
nor U13326 (N_13326,N_12946,N_12888);
nor U13327 (N_13327,N_13164,N_13197);
nor U13328 (N_13328,N_12607,N_12652);
xor U13329 (N_13329,N_13109,N_12714);
and U13330 (N_13330,N_13080,N_13157);
or U13331 (N_13331,N_12636,N_12684);
nand U13332 (N_13332,N_12734,N_12825);
nor U13333 (N_13333,N_12750,N_13110);
nand U13334 (N_13334,N_13045,N_13051);
xor U13335 (N_13335,N_12634,N_13022);
xnor U13336 (N_13336,N_12670,N_12741);
xnor U13337 (N_13337,N_12943,N_12745);
nor U13338 (N_13338,N_12874,N_13038);
nor U13339 (N_13339,N_12662,N_13067);
or U13340 (N_13340,N_12954,N_12976);
nand U13341 (N_13341,N_12821,N_12719);
or U13342 (N_13342,N_12842,N_12812);
nand U13343 (N_13343,N_12768,N_13192);
nor U13344 (N_13344,N_12881,N_12630);
and U13345 (N_13345,N_13159,N_13191);
nand U13346 (N_13346,N_12890,N_13124);
nor U13347 (N_13347,N_13097,N_12974);
xor U13348 (N_13348,N_12654,N_13000);
nand U13349 (N_13349,N_12706,N_13018);
xnor U13350 (N_13350,N_12769,N_13013);
and U13351 (N_13351,N_13046,N_12998);
xnor U13352 (N_13352,N_12973,N_12764);
xor U13353 (N_13353,N_12980,N_12832);
nand U13354 (N_13354,N_13076,N_13004);
xnor U13355 (N_13355,N_12977,N_13089);
and U13356 (N_13356,N_12932,N_13120);
xor U13357 (N_13357,N_13112,N_12701);
nor U13358 (N_13358,N_12663,N_13007);
and U13359 (N_13359,N_13069,N_12838);
nor U13360 (N_13360,N_12667,N_12921);
nor U13361 (N_13361,N_12651,N_13134);
xnor U13362 (N_13362,N_12911,N_13104);
and U13363 (N_13363,N_12677,N_13093);
and U13364 (N_13364,N_13040,N_12997);
nand U13365 (N_13365,N_12693,N_13026);
xor U13366 (N_13366,N_12937,N_13151);
and U13367 (N_13367,N_12754,N_12985);
xnor U13368 (N_13368,N_13183,N_12728);
xor U13369 (N_13369,N_12612,N_13056);
nand U13370 (N_13370,N_12624,N_13074);
nand U13371 (N_13371,N_12631,N_13030);
nor U13372 (N_13372,N_13090,N_13012);
nand U13373 (N_13373,N_12850,N_13190);
nand U13374 (N_13374,N_12622,N_12916);
nand U13375 (N_13375,N_13078,N_12733);
or U13376 (N_13376,N_12722,N_13081);
xor U13377 (N_13377,N_12871,N_13158);
xor U13378 (N_13378,N_13005,N_13052);
nor U13379 (N_13379,N_12657,N_12603);
nor U13380 (N_13380,N_12929,N_13127);
or U13381 (N_13381,N_12747,N_13195);
xnor U13382 (N_13382,N_12952,N_12730);
xnor U13383 (N_13383,N_12933,N_12746);
nand U13384 (N_13384,N_13165,N_13146);
or U13385 (N_13385,N_12619,N_13036);
xor U13386 (N_13386,N_12839,N_13082);
xnor U13387 (N_13387,N_12859,N_12923);
xor U13388 (N_13388,N_13128,N_12861);
xnor U13389 (N_13389,N_12600,N_13001);
nand U13390 (N_13390,N_12655,N_12846);
nand U13391 (N_13391,N_12694,N_12793);
nor U13392 (N_13392,N_12770,N_12659);
and U13393 (N_13393,N_12759,N_12661);
or U13394 (N_13394,N_13178,N_12605);
and U13395 (N_13395,N_12681,N_13032);
nor U13396 (N_13396,N_13176,N_12606);
xor U13397 (N_13397,N_13021,N_13121);
nand U13398 (N_13398,N_12949,N_13009);
or U13399 (N_13399,N_12731,N_12862);
xor U13400 (N_13400,N_12778,N_13111);
nand U13401 (N_13401,N_13050,N_13008);
nand U13402 (N_13402,N_13136,N_12901);
or U13403 (N_13403,N_12805,N_12685);
or U13404 (N_13404,N_12913,N_12726);
nor U13405 (N_13405,N_12905,N_12682);
xor U13406 (N_13406,N_13173,N_12798);
nand U13407 (N_13407,N_12992,N_13098);
nor U13408 (N_13408,N_12629,N_12779);
nand U13409 (N_13409,N_12647,N_12696);
or U13410 (N_13410,N_13115,N_13068);
nor U13411 (N_13411,N_13185,N_13141);
or U13412 (N_13412,N_12640,N_13194);
xor U13413 (N_13413,N_12813,N_12753);
nand U13414 (N_13414,N_12927,N_12924);
nor U13415 (N_13415,N_12686,N_12968);
nand U13416 (N_13416,N_13016,N_12665);
nand U13417 (N_13417,N_13028,N_12675);
xnor U13418 (N_13418,N_12789,N_12899);
or U13419 (N_13419,N_13167,N_13039);
xor U13420 (N_13420,N_12743,N_12702);
nand U13421 (N_13421,N_13100,N_12649);
xor U13422 (N_13422,N_13049,N_12990);
xnor U13423 (N_13423,N_12611,N_12928);
and U13424 (N_13424,N_12944,N_12664);
nand U13425 (N_13425,N_12823,N_12810);
nand U13426 (N_13426,N_12824,N_12960);
and U13427 (N_13427,N_12892,N_13154);
nor U13428 (N_13428,N_12635,N_13196);
nand U13429 (N_13429,N_12852,N_12610);
xnor U13430 (N_13430,N_12689,N_12653);
nor U13431 (N_13431,N_12864,N_12863);
nor U13432 (N_13432,N_13106,N_12638);
or U13433 (N_13433,N_12956,N_13193);
xor U13434 (N_13434,N_12844,N_13031);
nor U13435 (N_13435,N_13166,N_12919);
xor U13436 (N_13436,N_12800,N_13063);
nand U13437 (N_13437,N_12809,N_13139);
and U13438 (N_13438,N_12849,N_13152);
xnor U13439 (N_13439,N_12866,N_12687);
xor U13440 (N_13440,N_13143,N_12642);
or U13441 (N_13441,N_13017,N_12725);
or U13442 (N_13442,N_12896,N_12617);
nand U13443 (N_13443,N_12953,N_12891);
or U13444 (N_13444,N_12981,N_12867);
and U13445 (N_13445,N_12966,N_12727);
xor U13446 (N_13446,N_12942,N_12883);
and U13447 (N_13447,N_13130,N_12690);
nand U13448 (N_13448,N_12790,N_13086);
or U13449 (N_13449,N_13135,N_12897);
and U13450 (N_13450,N_13002,N_12784);
or U13451 (N_13451,N_12771,N_12982);
xnor U13452 (N_13452,N_12660,N_12766);
nor U13453 (N_13453,N_12780,N_13095);
xnor U13454 (N_13454,N_12740,N_13133);
xnor U13455 (N_13455,N_12776,N_13062);
xnor U13456 (N_13456,N_12672,N_12925);
or U13457 (N_13457,N_12729,N_12991);
nor U13458 (N_13458,N_12869,N_12749);
and U13459 (N_13459,N_12804,N_13180);
nand U13460 (N_13460,N_12994,N_12758);
xor U13461 (N_13461,N_12988,N_12835);
or U13462 (N_13462,N_12620,N_13125);
xnor U13463 (N_13463,N_12669,N_12837);
or U13464 (N_13464,N_12875,N_12621);
nor U13465 (N_13465,N_12872,N_13044);
xor U13466 (N_13466,N_12604,N_12723);
nor U13467 (N_13467,N_12792,N_13113);
nand U13468 (N_13468,N_13099,N_13023);
xor U13469 (N_13469,N_13059,N_12756);
or U13470 (N_13470,N_13092,N_12963);
xor U13471 (N_13471,N_12915,N_13138);
nor U13472 (N_13472,N_13188,N_12972);
and U13473 (N_13473,N_13131,N_12803);
and U13474 (N_13474,N_12920,N_12688);
xor U13475 (N_13475,N_12945,N_12922);
nand U13476 (N_13476,N_12836,N_12903);
nor U13477 (N_13477,N_13025,N_12969);
or U13478 (N_13478,N_12673,N_12609);
and U13479 (N_13479,N_13142,N_13140);
xor U13480 (N_13480,N_12955,N_12834);
nand U13481 (N_13481,N_12833,N_13037);
xnor U13482 (N_13482,N_13077,N_13107);
or U13483 (N_13483,N_12787,N_12794);
and U13484 (N_13484,N_13118,N_12971);
nand U13485 (N_13485,N_12626,N_13055);
nand U13486 (N_13486,N_12658,N_12894);
nand U13487 (N_13487,N_12735,N_12995);
and U13488 (N_13488,N_12996,N_12935);
nand U13489 (N_13489,N_12765,N_13047);
nor U13490 (N_13490,N_13015,N_12650);
nor U13491 (N_13491,N_13088,N_13162);
and U13492 (N_13492,N_12808,N_12775);
xor U13493 (N_13493,N_12983,N_12752);
and U13494 (N_13494,N_12931,N_12882);
or U13495 (N_13495,N_12841,N_13198);
nor U13496 (N_13496,N_13084,N_12958);
nand U13497 (N_13497,N_12987,N_12709);
and U13498 (N_13498,N_12989,N_12959);
or U13499 (N_13499,N_13117,N_12868);
xor U13500 (N_13500,N_12854,N_12873);
xnor U13501 (N_13501,N_13130,N_12665);
and U13502 (N_13502,N_12658,N_12687);
or U13503 (N_13503,N_13158,N_13144);
nand U13504 (N_13504,N_12945,N_13064);
nor U13505 (N_13505,N_13056,N_12605);
or U13506 (N_13506,N_13018,N_12982);
nor U13507 (N_13507,N_12878,N_13095);
or U13508 (N_13508,N_13068,N_12625);
and U13509 (N_13509,N_12989,N_12942);
or U13510 (N_13510,N_12614,N_12870);
or U13511 (N_13511,N_13010,N_13012);
and U13512 (N_13512,N_12943,N_13199);
xnor U13513 (N_13513,N_12736,N_12681);
nor U13514 (N_13514,N_12867,N_12978);
or U13515 (N_13515,N_12669,N_12656);
xnor U13516 (N_13516,N_12650,N_12764);
nand U13517 (N_13517,N_13063,N_13182);
or U13518 (N_13518,N_12617,N_12780);
or U13519 (N_13519,N_12782,N_13189);
nor U13520 (N_13520,N_13120,N_12760);
nand U13521 (N_13521,N_12985,N_13101);
or U13522 (N_13522,N_12887,N_12687);
or U13523 (N_13523,N_12758,N_12680);
nand U13524 (N_13524,N_13116,N_12787);
nand U13525 (N_13525,N_12908,N_12772);
and U13526 (N_13526,N_13041,N_12880);
nor U13527 (N_13527,N_12840,N_13134);
or U13528 (N_13528,N_12950,N_13009);
or U13529 (N_13529,N_12793,N_13181);
nand U13530 (N_13530,N_13178,N_13068);
xor U13531 (N_13531,N_12648,N_12646);
nor U13532 (N_13532,N_13092,N_12694);
or U13533 (N_13533,N_12757,N_12913);
nand U13534 (N_13534,N_12970,N_12806);
xnor U13535 (N_13535,N_12778,N_13133);
nand U13536 (N_13536,N_12701,N_12928);
nand U13537 (N_13537,N_12906,N_12892);
nand U13538 (N_13538,N_12656,N_12654);
and U13539 (N_13539,N_13121,N_12914);
xnor U13540 (N_13540,N_12719,N_12750);
nor U13541 (N_13541,N_12894,N_13150);
or U13542 (N_13542,N_13180,N_12802);
nand U13543 (N_13543,N_12944,N_12814);
nand U13544 (N_13544,N_12865,N_13175);
nor U13545 (N_13545,N_12892,N_12789);
and U13546 (N_13546,N_12635,N_13097);
or U13547 (N_13547,N_13175,N_12868);
and U13548 (N_13548,N_12749,N_13069);
nor U13549 (N_13549,N_12664,N_13091);
nand U13550 (N_13550,N_13132,N_12891);
nand U13551 (N_13551,N_12694,N_13124);
or U13552 (N_13552,N_13087,N_12830);
or U13553 (N_13553,N_13191,N_12829);
nor U13554 (N_13554,N_12758,N_12858);
and U13555 (N_13555,N_13127,N_12949);
and U13556 (N_13556,N_13010,N_12758);
or U13557 (N_13557,N_13015,N_13125);
nand U13558 (N_13558,N_12897,N_13190);
nor U13559 (N_13559,N_12871,N_12872);
nor U13560 (N_13560,N_12907,N_12911);
or U13561 (N_13561,N_12850,N_12950);
and U13562 (N_13562,N_13079,N_12950);
nand U13563 (N_13563,N_12753,N_13041);
nor U13564 (N_13564,N_12978,N_12880);
nand U13565 (N_13565,N_12635,N_13062);
or U13566 (N_13566,N_13074,N_12870);
and U13567 (N_13567,N_12827,N_13061);
nor U13568 (N_13568,N_12803,N_13178);
nand U13569 (N_13569,N_13101,N_12740);
or U13570 (N_13570,N_13111,N_13124);
or U13571 (N_13571,N_12824,N_13020);
xnor U13572 (N_13572,N_12658,N_13161);
and U13573 (N_13573,N_13153,N_12898);
xnor U13574 (N_13574,N_12754,N_12734);
and U13575 (N_13575,N_13195,N_12616);
xor U13576 (N_13576,N_12799,N_12632);
or U13577 (N_13577,N_12801,N_12979);
or U13578 (N_13578,N_13143,N_13060);
nor U13579 (N_13579,N_13154,N_12712);
and U13580 (N_13580,N_12889,N_12809);
nand U13581 (N_13581,N_13067,N_13032);
or U13582 (N_13582,N_12903,N_12710);
xnor U13583 (N_13583,N_13199,N_13022);
nand U13584 (N_13584,N_12898,N_13044);
or U13585 (N_13585,N_12718,N_13027);
xor U13586 (N_13586,N_13064,N_12732);
or U13587 (N_13587,N_12843,N_12936);
and U13588 (N_13588,N_12660,N_12637);
nand U13589 (N_13589,N_12979,N_13018);
or U13590 (N_13590,N_12941,N_12669);
nand U13591 (N_13591,N_12655,N_13011);
or U13592 (N_13592,N_13041,N_13139);
xnor U13593 (N_13593,N_13114,N_12789);
xor U13594 (N_13594,N_12610,N_12701);
xnor U13595 (N_13595,N_12873,N_13059);
or U13596 (N_13596,N_12814,N_13197);
nor U13597 (N_13597,N_12889,N_12876);
and U13598 (N_13598,N_12686,N_12605);
and U13599 (N_13599,N_12742,N_13045);
and U13600 (N_13600,N_13165,N_13046);
nor U13601 (N_13601,N_13003,N_12876);
and U13602 (N_13602,N_13041,N_12693);
nand U13603 (N_13603,N_12928,N_13041);
nor U13604 (N_13604,N_12763,N_12714);
xor U13605 (N_13605,N_13138,N_13083);
and U13606 (N_13606,N_12970,N_13151);
and U13607 (N_13607,N_12968,N_13161);
and U13608 (N_13608,N_12806,N_13016);
xor U13609 (N_13609,N_13121,N_13103);
nand U13610 (N_13610,N_12806,N_12743);
and U13611 (N_13611,N_13075,N_13049);
xor U13612 (N_13612,N_12839,N_12787);
or U13613 (N_13613,N_12902,N_12652);
nor U13614 (N_13614,N_12747,N_13134);
nor U13615 (N_13615,N_12985,N_13121);
nor U13616 (N_13616,N_12705,N_13161);
nor U13617 (N_13617,N_12877,N_12712);
or U13618 (N_13618,N_12628,N_12951);
nor U13619 (N_13619,N_12854,N_13188);
and U13620 (N_13620,N_13163,N_13111);
xnor U13621 (N_13621,N_12615,N_13184);
or U13622 (N_13622,N_12687,N_12642);
and U13623 (N_13623,N_12656,N_13036);
xnor U13624 (N_13624,N_12802,N_12824);
or U13625 (N_13625,N_13028,N_12909);
or U13626 (N_13626,N_12663,N_12889);
or U13627 (N_13627,N_12783,N_12643);
and U13628 (N_13628,N_13030,N_13034);
or U13629 (N_13629,N_12714,N_12693);
nand U13630 (N_13630,N_12824,N_12944);
or U13631 (N_13631,N_12727,N_12873);
nand U13632 (N_13632,N_12812,N_12884);
or U13633 (N_13633,N_12812,N_13002);
or U13634 (N_13634,N_12966,N_12659);
nor U13635 (N_13635,N_12984,N_12772);
and U13636 (N_13636,N_13097,N_13098);
nand U13637 (N_13637,N_12768,N_12972);
nand U13638 (N_13638,N_13146,N_12819);
or U13639 (N_13639,N_12944,N_12698);
xor U13640 (N_13640,N_12831,N_13144);
nand U13641 (N_13641,N_12830,N_12938);
nor U13642 (N_13642,N_12916,N_12771);
nor U13643 (N_13643,N_13005,N_12991);
nand U13644 (N_13644,N_13024,N_13104);
and U13645 (N_13645,N_12662,N_13111);
or U13646 (N_13646,N_12988,N_12609);
xnor U13647 (N_13647,N_12704,N_12622);
nor U13648 (N_13648,N_12711,N_13029);
and U13649 (N_13649,N_12952,N_12627);
nand U13650 (N_13650,N_12774,N_12677);
and U13651 (N_13651,N_12816,N_13163);
nand U13652 (N_13652,N_13108,N_12782);
or U13653 (N_13653,N_13104,N_12829);
nand U13654 (N_13654,N_12600,N_12612);
xnor U13655 (N_13655,N_13096,N_12710);
xor U13656 (N_13656,N_12785,N_12777);
nor U13657 (N_13657,N_12610,N_12617);
nand U13658 (N_13658,N_12824,N_13194);
xnor U13659 (N_13659,N_12871,N_12909);
nor U13660 (N_13660,N_12648,N_12611);
nand U13661 (N_13661,N_12853,N_12882);
or U13662 (N_13662,N_12958,N_12827);
or U13663 (N_13663,N_12998,N_12858);
or U13664 (N_13664,N_12907,N_12815);
nand U13665 (N_13665,N_13141,N_12732);
and U13666 (N_13666,N_12799,N_13106);
xnor U13667 (N_13667,N_12769,N_12860);
nand U13668 (N_13668,N_12682,N_12617);
nand U13669 (N_13669,N_12949,N_13020);
xor U13670 (N_13670,N_12651,N_12864);
nand U13671 (N_13671,N_12610,N_12861);
and U13672 (N_13672,N_12627,N_13154);
nor U13673 (N_13673,N_12986,N_12617);
nand U13674 (N_13674,N_13059,N_12894);
xnor U13675 (N_13675,N_12659,N_12911);
or U13676 (N_13676,N_12969,N_13030);
nand U13677 (N_13677,N_13184,N_13197);
xnor U13678 (N_13678,N_13145,N_12836);
or U13679 (N_13679,N_13095,N_12914);
nor U13680 (N_13680,N_12829,N_13067);
xnor U13681 (N_13681,N_13173,N_12635);
and U13682 (N_13682,N_13076,N_13049);
and U13683 (N_13683,N_12867,N_13012);
nor U13684 (N_13684,N_12666,N_12674);
or U13685 (N_13685,N_12940,N_13155);
xor U13686 (N_13686,N_12787,N_12654);
nor U13687 (N_13687,N_12907,N_12866);
nand U13688 (N_13688,N_12819,N_12812);
and U13689 (N_13689,N_12917,N_12692);
nand U13690 (N_13690,N_12739,N_12806);
and U13691 (N_13691,N_13186,N_12886);
nand U13692 (N_13692,N_12933,N_13051);
nor U13693 (N_13693,N_12936,N_12860);
nor U13694 (N_13694,N_12895,N_12985);
or U13695 (N_13695,N_12852,N_12913);
or U13696 (N_13696,N_12759,N_12794);
nand U13697 (N_13697,N_12650,N_12668);
and U13698 (N_13698,N_12733,N_13184);
or U13699 (N_13699,N_13190,N_12630);
xor U13700 (N_13700,N_12611,N_12655);
nor U13701 (N_13701,N_13021,N_12668);
nand U13702 (N_13702,N_13044,N_12930);
nand U13703 (N_13703,N_13059,N_12900);
xor U13704 (N_13704,N_12830,N_12802);
nor U13705 (N_13705,N_12612,N_12658);
xor U13706 (N_13706,N_12963,N_13188);
xnor U13707 (N_13707,N_13041,N_12616);
or U13708 (N_13708,N_13193,N_12867);
xor U13709 (N_13709,N_13129,N_13071);
nor U13710 (N_13710,N_12977,N_13097);
nor U13711 (N_13711,N_13116,N_13134);
xnor U13712 (N_13712,N_13098,N_13009);
or U13713 (N_13713,N_13128,N_13118);
xor U13714 (N_13714,N_12998,N_12965);
nor U13715 (N_13715,N_12684,N_12867);
or U13716 (N_13716,N_12870,N_13141);
or U13717 (N_13717,N_12996,N_13043);
nor U13718 (N_13718,N_13017,N_13163);
nand U13719 (N_13719,N_13033,N_12910);
or U13720 (N_13720,N_12881,N_12940);
nor U13721 (N_13721,N_12911,N_12967);
or U13722 (N_13722,N_12868,N_12601);
and U13723 (N_13723,N_12935,N_12717);
nand U13724 (N_13724,N_12959,N_12848);
or U13725 (N_13725,N_12830,N_12928);
nand U13726 (N_13726,N_13138,N_12950);
and U13727 (N_13727,N_12855,N_12924);
xnor U13728 (N_13728,N_13152,N_13192);
xnor U13729 (N_13729,N_12600,N_12978);
or U13730 (N_13730,N_12854,N_12815);
xnor U13731 (N_13731,N_13154,N_12921);
nor U13732 (N_13732,N_13101,N_12900);
nor U13733 (N_13733,N_13139,N_12770);
nand U13734 (N_13734,N_13042,N_13012);
xor U13735 (N_13735,N_12753,N_13109);
xnor U13736 (N_13736,N_12980,N_13161);
nand U13737 (N_13737,N_13182,N_12995);
nand U13738 (N_13738,N_12660,N_12687);
nand U13739 (N_13739,N_13022,N_12680);
and U13740 (N_13740,N_12869,N_12607);
nor U13741 (N_13741,N_12790,N_12917);
xor U13742 (N_13742,N_13082,N_12717);
xnor U13743 (N_13743,N_12699,N_12967);
nand U13744 (N_13744,N_12878,N_12831);
or U13745 (N_13745,N_13171,N_13070);
nor U13746 (N_13746,N_12631,N_13179);
or U13747 (N_13747,N_13001,N_13087);
xor U13748 (N_13748,N_12776,N_12916);
and U13749 (N_13749,N_12948,N_13039);
nor U13750 (N_13750,N_13170,N_13129);
or U13751 (N_13751,N_12950,N_13032);
xnor U13752 (N_13752,N_12691,N_12888);
nand U13753 (N_13753,N_12808,N_12770);
or U13754 (N_13754,N_13133,N_13087);
nand U13755 (N_13755,N_12705,N_12708);
xnor U13756 (N_13756,N_12848,N_12891);
xor U13757 (N_13757,N_13122,N_13149);
xnor U13758 (N_13758,N_13087,N_12761);
nand U13759 (N_13759,N_13185,N_12928);
or U13760 (N_13760,N_12882,N_12968);
xor U13761 (N_13761,N_12803,N_12766);
nor U13762 (N_13762,N_13076,N_13036);
and U13763 (N_13763,N_13173,N_12837);
nand U13764 (N_13764,N_13124,N_12942);
xor U13765 (N_13765,N_12866,N_12960);
or U13766 (N_13766,N_12727,N_12990);
and U13767 (N_13767,N_12892,N_12923);
nand U13768 (N_13768,N_12906,N_13129);
xnor U13769 (N_13769,N_12872,N_13184);
xnor U13770 (N_13770,N_12848,N_12612);
nand U13771 (N_13771,N_12611,N_13138);
and U13772 (N_13772,N_12691,N_13198);
nand U13773 (N_13773,N_13143,N_12689);
and U13774 (N_13774,N_12910,N_13117);
nor U13775 (N_13775,N_12840,N_12990);
and U13776 (N_13776,N_12633,N_12786);
or U13777 (N_13777,N_12752,N_12680);
or U13778 (N_13778,N_13002,N_12819);
nand U13779 (N_13779,N_12676,N_12633);
nor U13780 (N_13780,N_12894,N_12851);
or U13781 (N_13781,N_13072,N_12892);
nor U13782 (N_13782,N_12948,N_12775);
xnor U13783 (N_13783,N_12693,N_12736);
xor U13784 (N_13784,N_13185,N_13054);
nor U13785 (N_13785,N_12986,N_12920);
xor U13786 (N_13786,N_13039,N_13125);
and U13787 (N_13787,N_13118,N_12933);
or U13788 (N_13788,N_12772,N_12978);
and U13789 (N_13789,N_13061,N_13085);
nand U13790 (N_13790,N_12766,N_12600);
and U13791 (N_13791,N_13182,N_12931);
and U13792 (N_13792,N_12873,N_12761);
and U13793 (N_13793,N_12759,N_13039);
and U13794 (N_13794,N_13023,N_13162);
and U13795 (N_13795,N_12948,N_12994);
and U13796 (N_13796,N_12824,N_12891);
or U13797 (N_13797,N_12806,N_12945);
or U13798 (N_13798,N_12920,N_13103);
or U13799 (N_13799,N_12857,N_13137);
nor U13800 (N_13800,N_13747,N_13243);
or U13801 (N_13801,N_13498,N_13655);
or U13802 (N_13802,N_13669,N_13638);
or U13803 (N_13803,N_13579,N_13622);
nor U13804 (N_13804,N_13516,N_13640);
nor U13805 (N_13805,N_13678,N_13528);
nand U13806 (N_13806,N_13756,N_13418);
nand U13807 (N_13807,N_13580,N_13512);
and U13808 (N_13808,N_13455,N_13281);
nand U13809 (N_13809,N_13641,N_13203);
xor U13810 (N_13810,N_13362,N_13597);
nor U13811 (N_13811,N_13687,N_13639);
nor U13812 (N_13812,N_13371,N_13344);
or U13813 (N_13813,N_13269,N_13636);
xor U13814 (N_13814,N_13436,N_13340);
xnor U13815 (N_13815,N_13753,N_13754);
xnor U13816 (N_13816,N_13353,N_13306);
and U13817 (N_13817,N_13624,N_13534);
nand U13818 (N_13818,N_13331,N_13595);
nor U13819 (N_13819,N_13283,N_13410);
and U13820 (N_13820,N_13682,N_13521);
and U13821 (N_13821,N_13704,N_13642);
xor U13822 (N_13822,N_13529,N_13791);
and U13823 (N_13823,N_13329,N_13411);
nand U13824 (N_13824,N_13261,N_13322);
or U13825 (N_13825,N_13457,N_13231);
nand U13826 (N_13826,N_13746,N_13327);
nand U13827 (N_13827,N_13559,N_13279);
nor U13828 (N_13828,N_13317,N_13438);
and U13829 (N_13829,N_13648,N_13225);
nor U13830 (N_13830,N_13617,N_13675);
nor U13831 (N_13831,N_13369,N_13573);
nor U13832 (N_13832,N_13705,N_13337);
and U13833 (N_13833,N_13338,N_13471);
xnor U13834 (N_13834,N_13263,N_13275);
nand U13835 (N_13835,N_13771,N_13428);
nand U13836 (N_13836,N_13510,N_13702);
and U13837 (N_13837,N_13799,N_13793);
nor U13838 (N_13838,N_13776,N_13718);
nor U13839 (N_13839,N_13432,N_13672);
nor U13840 (N_13840,N_13554,N_13449);
nor U13841 (N_13841,N_13437,N_13752);
xor U13842 (N_13842,N_13764,N_13658);
or U13843 (N_13843,N_13538,N_13422);
nand U13844 (N_13844,N_13271,N_13242);
and U13845 (N_13845,N_13312,N_13465);
and U13846 (N_13846,N_13762,N_13213);
xnor U13847 (N_13847,N_13478,N_13551);
nand U13848 (N_13848,N_13208,N_13310);
and U13849 (N_13849,N_13740,N_13223);
or U13850 (N_13850,N_13739,N_13767);
nor U13851 (N_13851,N_13435,N_13433);
nand U13852 (N_13852,N_13325,N_13651);
xor U13853 (N_13853,N_13558,N_13526);
xnor U13854 (N_13854,N_13509,N_13377);
nand U13855 (N_13855,N_13626,N_13720);
nand U13856 (N_13856,N_13466,N_13241);
and U13857 (N_13857,N_13253,N_13605);
nor U13858 (N_13858,N_13772,N_13524);
nor U13859 (N_13859,N_13450,N_13204);
nor U13860 (N_13860,N_13616,N_13345);
and U13861 (N_13861,N_13205,N_13453);
or U13862 (N_13862,N_13691,N_13557);
nor U13863 (N_13863,N_13237,N_13659);
xor U13864 (N_13864,N_13259,N_13520);
nor U13865 (N_13865,N_13489,N_13211);
xor U13866 (N_13866,N_13630,N_13496);
or U13867 (N_13867,N_13603,N_13376);
and U13868 (N_13868,N_13488,N_13300);
nand U13869 (N_13869,N_13485,N_13599);
xor U13870 (N_13870,N_13715,N_13320);
xnor U13871 (N_13871,N_13459,N_13500);
nor U13872 (N_13872,N_13535,N_13236);
and U13873 (N_13873,N_13696,N_13710);
nor U13874 (N_13874,N_13571,N_13260);
and U13875 (N_13875,N_13610,N_13276);
or U13876 (N_13876,N_13224,N_13423);
or U13877 (N_13877,N_13350,N_13635);
xor U13878 (N_13878,N_13370,N_13222);
and U13879 (N_13879,N_13343,N_13692);
xnor U13880 (N_13880,N_13606,N_13654);
and U13881 (N_13881,N_13665,N_13592);
xnor U13882 (N_13882,N_13749,N_13722);
and U13883 (N_13883,N_13656,N_13620);
and U13884 (N_13884,N_13584,N_13447);
or U13885 (N_13885,N_13779,N_13293);
nor U13886 (N_13886,N_13701,N_13229);
xnor U13887 (N_13887,N_13266,N_13519);
nand U13888 (N_13888,N_13686,N_13618);
xor U13889 (N_13889,N_13598,N_13456);
or U13890 (N_13890,N_13246,N_13650);
nand U13891 (N_13891,N_13602,N_13484);
xnor U13892 (N_13892,N_13632,N_13378);
or U13893 (N_13893,N_13763,N_13416);
and U13894 (N_13894,N_13594,N_13609);
nand U13895 (N_13895,N_13738,N_13784);
nand U13896 (N_13896,N_13365,N_13566);
or U13897 (N_13897,N_13364,N_13613);
nand U13898 (N_13898,N_13219,N_13792);
and U13899 (N_13899,N_13462,N_13798);
and U13900 (N_13900,N_13412,N_13244);
xor U13901 (N_13901,N_13570,N_13522);
xor U13902 (N_13902,N_13318,N_13766);
and U13903 (N_13903,N_13273,N_13623);
nor U13904 (N_13904,N_13612,N_13321);
nand U13905 (N_13905,N_13759,N_13401);
nor U13906 (N_13906,N_13499,N_13444);
and U13907 (N_13907,N_13506,N_13716);
xnor U13908 (N_13908,N_13424,N_13288);
nand U13909 (N_13909,N_13742,N_13326);
nand U13910 (N_13910,N_13398,N_13730);
or U13911 (N_13911,N_13434,N_13287);
nand U13912 (N_13912,N_13707,N_13304);
or U13913 (N_13913,N_13482,N_13414);
or U13914 (N_13914,N_13479,N_13363);
and U13915 (N_13915,N_13341,N_13727);
and U13916 (N_13916,N_13218,N_13228);
nor U13917 (N_13917,N_13472,N_13569);
or U13918 (N_13918,N_13697,N_13296);
nor U13919 (N_13919,N_13706,N_13693);
and U13920 (N_13920,N_13247,N_13663);
xor U13921 (N_13921,N_13591,N_13307);
or U13922 (N_13922,N_13530,N_13240);
xor U13923 (N_13923,N_13770,N_13562);
nor U13924 (N_13924,N_13621,N_13700);
nor U13925 (N_13925,N_13585,N_13593);
or U13926 (N_13926,N_13789,N_13666);
nor U13927 (N_13927,N_13583,N_13421);
xnor U13928 (N_13928,N_13454,N_13653);
or U13929 (N_13929,N_13206,N_13564);
or U13930 (N_13930,N_13390,N_13335);
xor U13931 (N_13931,N_13785,N_13234);
and U13932 (N_13932,N_13731,N_13245);
xor U13933 (N_13933,N_13388,N_13387);
nor U13934 (N_13934,N_13212,N_13272);
nor U13935 (N_13935,N_13282,N_13588);
and U13936 (N_13936,N_13568,N_13607);
nor U13937 (N_13937,N_13695,N_13474);
nor U13938 (N_13938,N_13502,N_13572);
xnor U13939 (N_13939,N_13774,N_13575);
xnor U13940 (N_13940,N_13504,N_13647);
nand U13941 (N_13941,N_13513,N_13633);
xnor U13942 (N_13942,N_13761,N_13452);
nand U13943 (N_13943,N_13578,N_13589);
and U13944 (N_13944,N_13688,N_13525);
xnor U13945 (N_13945,N_13646,N_13743);
and U13946 (N_13946,N_13278,N_13460);
nor U13947 (N_13947,N_13501,N_13544);
nand U13948 (N_13948,N_13448,N_13409);
nand U13949 (N_13949,N_13230,N_13262);
nor U13950 (N_13950,N_13426,N_13332);
and U13951 (N_13951,N_13794,N_13417);
nor U13952 (N_13952,N_13728,N_13748);
or U13953 (N_13953,N_13375,N_13468);
or U13954 (N_13954,N_13667,N_13355);
or U13955 (N_13955,N_13649,N_13674);
or U13956 (N_13956,N_13662,N_13407);
xnor U13957 (N_13957,N_13539,N_13415);
or U13958 (N_13958,N_13797,N_13379);
and U13959 (N_13959,N_13627,N_13373);
or U13960 (N_13960,N_13209,N_13393);
xnor U13961 (N_13961,N_13406,N_13637);
or U13962 (N_13962,N_13419,N_13625);
or U13963 (N_13963,N_13291,N_13352);
nor U13964 (N_13964,N_13391,N_13565);
or U13965 (N_13965,N_13297,N_13795);
and U13966 (N_13966,N_13473,N_13685);
and U13967 (N_13967,N_13267,N_13323);
or U13968 (N_13968,N_13721,N_13541);
nor U13969 (N_13969,N_13671,N_13425);
nand U13970 (N_13970,N_13439,N_13475);
nor U13971 (N_13971,N_13790,N_13545);
and U13972 (N_13972,N_13250,N_13493);
or U13973 (N_13973,N_13392,N_13354);
and U13974 (N_13974,N_13429,N_13374);
xnor U13975 (N_13975,N_13221,N_13408);
nand U13976 (N_13976,N_13239,N_13470);
nor U13977 (N_13977,N_13295,N_13458);
and U13978 (N_13978,N_13596,N_13290);
or U13979 (N_13979,N_13760,N_13681);
nand U13980 (N_13980,N_13563,N_13305);
and U13981 (N_13981,N_13200,N_13333);
or U13982 (N_13982,N_13777,N_13301);
and U13983 (N_13983,N_13768,N_13342);
or U13984 (N_13984,N_13631,N_13395);
nand U13985 (N_13985,N_13531,N_13284);
xnor U13986 (N_13986,N_13280,N_13552);
xor U13987 (N_13987,N_13644,N_13645);
and U13988 (N_13988,N_13679,N_13628);
or U13989 (N_13989,N_13664,N_13389);
and U13990 (N_13990,N_13782,N_13490);
and U13991 (N_13991,N_13615,N_13258);
nand U13992 (N_13992,N_13315,N_13487);
and U13993 (N_13993,N_13336,N_13724);
and U13994 (N_13994,N_13733,N_13709);
xor U13995 (N_13995,N_13503,N_13586);
nand U13996 (N_13996,N_13492,N_13788);
nor U13997 (N_13997,N_13372,N_13382);
or U13998 (N_13998,N_13796,N_13548);
and U13999 (N_13999,N_13268,N_13289);
nand U14000 (N_14000,N_13590,N_13294);
or U14001 (N_14001,N_13608,N_13256);
and U14002 (N_14002,N_13677,N_13735);
xnor U14003 (N_14003,N_13351,N_13446);
and U14004 (N_14004,N_13311,N_13313);
nand U14005 (N_14005,N_13399,N_13238);
and U14006 (N_14006,N_13302,N_13201);
or U14007 (N_14007,N_13330,N_13634);
nand U14008 (N_14008,N_13361,N_13532);
xor U14009 (N_14009,N_13694,N_13712);
nand U14010 (N_14010,N_13546,N_13316);
nor U14011 (N_14011,N_13508,N_13385);
nor U14012 (N_14012,N_13339,N_13517);
nor U14013 (N_14013,N_13476,N_13334);
xnor U14014 (N_14014,N_13367,N_13614);
xor U14015 (N_14015,N_13582,N_13285);
or U14016 (N_14016,N_13758,N_13708);
and U14017 (N_14017,N_13619,N_13440);
nand U14018 (N_14018,N_13741,N_13477);
xor U14019 (N_14019,N_13540,N_13547);
and U14020 (N_14020,N_13726,N_13483);
xor U14021 (N_14021,N_13254,N_13381);
and U14022 (N_14022,N_13217,N_13673);
nor U14023 (N_14023,N_13576,N_13404);
xor U14024 (N_14024,N_13292,N_13783);
and U14025 (N_14025,N_13380,N_13308);
nor U14026 (N_14026,N_13543,N_13561);
and U14027 (N_14027,N_13358,N_13745);
and U14028 (N_14028,N_13577,N_13420);
nand U14029 (N_14029,N_13714,N_13486);
or U14030 (N_14030,N_13676,N_13441);
xor U14031 (N_14031,N_13781,N_13751);
xnor U14032 (N_14032,N_13734,N_13265);
or U14033 (N_14033,N_13397,N_13303);
nand U14034 (N_14034,N_13668,N_13553);
nand U14035 (N_14035,N_13732,N_13723);
nor U14036 (N_14036,N_13773,N_13765);
nor U14037 (N_14037,N_13233,N_13314);
nor U14038 (N_14038,N_13383,N_13549);
nand U14039 (N_14039,N_13348,N_13481);
xor U14040 (N_14040,N_13356,N_13386);
and U14041 (N_14041,N_13480,N_13207);
xor U14042 (N_14042,N_13220,N_13427);
nor U14043 (N_14043,N_13737,N_13443);
nand U14044 (N_14044,N_13347,N_13319);
or U14045 (N_14045,N_13787,N_13463);
nor U14046 (N_14046,N_13368,N_13270);
or U14047 (N_14047,N_13264,N_13680);
xor U14048 (N_14048,N_13309,N_13769);
and U14049 (N_14049,N_13725,N_13711);
xnor U14050 (N_14050,N_13515,N_13442);
xnor U14051 (N_14051,N_13683,N_13689);
nor U14052 (N_14052,N_13560,N_13366);
or U14053 (N_14053,N_13251,N_13775);
nor U14054 (N_14054,N_13384,N_13445);
and U14055 (N_14055,N_13467,N_13527);
and U14056 (N_14056,N_13713,N_13719);
and U14057 (N_14057,N_13717,N_13226);
nor U14058 (N_14058,N_13277,N_13232);
nand U14059 (N_14059,N_13349,N_13359);
nand U14060 (N_14060,N_13744,N_13214);
and U14061 (N_14061,N_13451,N_13587);
nand U14062 (N_14062,N_13657,N_13690);
nor U14063 (N_14063,N_13698,N_13523);
or U14064 (N_14064,N_13328,N_13215);
xor U14065 (N_14065,N_13643,N_13507);
nand U14066 (N_14066,N_13537,N_13413);
xor U14067 (N_14067,N_13567,N_13255);
and U14068 (N_14068,N_13661,N_13299);
xnor U14069 (N_14069,N_13518,N_13400);
nor U14070 (N_14070,N_13629,N_13430);
xor U14071 (N_14071,N_13511,N_13249);
nor U14072 (N_14072,N_13464,N_13699);
nor U14073 (N_14073,N_13461,N_13469);
and U14074 (N_14074,N_13778,N_13505);
nand U14075 (N_14075,N_13604,N_13574);
nand U14076 (N_14076,N_13216,N_13555);
nor U14077 (N_14077,N_13670,N_13514);
nor U14078 (N_14078,N_13495,N_13494);
or U14079 (N_14079,N_13403,N_13786);
xor U14080 (N_14080,N_13405,N_13298);
xor U14081 (N_14081,N_13703,N_13210);
or U14082 (N_14082,N_13274,N_13497);
and U14083 (N_14083,N_13431,N_13202);
nand U14084 (N_14084,N_13248,N_13360);
xor U14085 (N_14085,N_13252,N_13396);
nand U14086 (N_14086,N_13491,N_13581);
nor U14087 (N_14087,N_13402,N_13755);
and U14088 (N_14088,N_13257,N_13601);
and U14089 (N_14089,N_13357,N_13324);
nor U14090 (N_14090,N_13536,N_13660);
nand U14091 (N_14091,N_13757,N_13736);
nand U14092 (N_14092,N_13684,N_13600);
nand U14093 (N_14093,N_13542,N_13611);
nand U14094 (N_14094,N_13533,N_13394);
nand U14095 (N_14095,N_13550,N_13286);
xnor U14096 (N_14096,N_13227,N_13750);
xnor U14097 (N_14097,N_13346,N_13652);
or U14098 (N_14098,N_13235,N_13780);
nand U14099 (N_14099,N_13729,N_13556);
xor U14100 (N_14100,N_13716,N_13574);
xor U14101 (N_14101,N_13597,N_13232);
and U14102 (N_14102,N_13740,N_13229);
xnor U14103 (N_14103,N_13629,N_13291);
and U14104 (N_14104,N_13212,N_13799);
xnor U14105 (N_14105,N_13640,N_13207);
or U14106 (N_14106,N_13502,N_13778);
nand U14107 (N_14107,N_13427,N_13416);
nor U14108 (N_14108,N_13463,N_13320);
nor U14109 (N_14109,N_13589,N_13432);
nand U14110 (N_14110,N_13472,N_13565);
nor U14111 (N_14111,N_13799,N_13389);
nand U14112 (N_14112,N_13406,N_13582);
nor U14113 (N_14113,N_13744,N_13296);
or U14114 (N_14114,N_13370,N_13504);
nand U14115 (N_14115,N_13321,N_13416);
xnor U14116 (N_14116,N_13584,N_13391);
and U14117 (N_14117,N_13478,N_13597);
xnor U14118 (N_14118,N_13342,N_13373);
xor U14119 (N_14119,N_13690,N_13450);
nand U14120 (N_14120,N_13675,N_13463);
and U14121 (N_14121,N_13627,N_13423);
and U14122 (N_14122,N_13227,N_13346);
nand U14123 (N_14123,N_13277,N_13279);
xnor U14124 (N_14124,N_13240,N_13780);
xnor U14125 (N_14125,N_13389,N_13358);
nor U14126 (N_14126,N_13554,N_13433);
nor U14127 (N_14127,N_13387,N_13393);
nor U14128 (N_14128,N_13556,N_13777);
or U14129 (N_14129,N_13392,N_13448);
nor U14130 (N_14130,N_13679,N_13304);
or U14131 (N_14131,N_13213,N_13798);
nand U14132 (N_14132,N_13435,N_13790);
xor U14133 (N_14133,N_13424,N_13433);
and U14134 (N_14134,N_13519,N_13328);
xnor U14135 (N_14135,N_13283,N_13556);
xor U14136 (N_14136,N_13408,N_13351);
nand U14137 (N_14137,N_13406,N_13736);
xor U14138 (N_14138,N_13285,N_13574);
nor U14139 (N_14139,N_13672,N_13483);
or U14140 (N_14140,N_13499,N_13397);
nand U14141 (N_14141,N_13407,N_13730);
or U14142 (N_14142,N_13612,N_13224);
or U14143 (N_14143,N_13709,N_13265);
xnor U14144 (N_14144,N_13204,N_13598);
or U14145 (N_14145,N_13555,N_13488);
xor U14146 (N_14146,N_13754,N_13213);
and U14147 (N_14147,N_13666,N_13508);
and U14148 (N_14148,N_13529,N_13647);
nand U14149 (N_14149,N_13468,N_13339);
nor U14150 (N_14150,N_13441,N_13201);
nor U14151 (N_14151,N_13412,N_13628);
nor U14152 (N_14152,N_13424,N_13236);
or U14153 (N_14153,N_13330,N_13490);
and U14154 (N_14154,N_13237,N_13554);
and U14155 (N_14155,N_13469,N_13595);
xnor U14156 (N_14156,N_13328,N_13286);
or U14157 (N_14157,N_13237,N_13710);
nand U14158 (N_14158,N_13211,N_13799);
or U14159 (N_14159,N_13602,N_13621);
nor U14160 (N_14160,N_13597,N_13720);
xnor U14161 (N_14161,N_13677,N_13464);
or U14162 (N_14162,N_13588,N_13251);
xor U14163 (N_14163,N_13248,N_13455);
xnor U14164 (N_14164,N_13211,N_13643);
nand U14165 (N_14165,N_13627,N_13452);
nor U14166 (N_14166,N_13643,N_13274);
and U14167 (N_14167,N_13398,N_13320);
nor U14168 (N_14168,N_13528,N_13397);
and U14169 (N_14169,N_13483,N_13484);
xor U14170 (N_14170,N_13624,N_13208);
nand U14171 (N_14171,N_13335,N_13641);
or U14172 (N_14172,N_13672,N_13620);
nand U14173 (N_14173,N_13538,N_13490);
nand U14174 (N_14174,N_13398,N_13799);
nand U14175 (N_14175,N_13362,N_13745);
xor U14176 (N_14176,N_13223,N_13435);
or U14177 (N_14177,N_13573,N_13563);
nand U14178 (N_14178,N_13324,N_13790);
nor U14179 (N_14179,N_13278,N_13233);
nand U14180 (N_14180,N_13562,N_13675);
nor U14181 (N_14181,N_13294,N_13588);
and U14182 (N_14182,N_13751,N_13638);
nor U14183 (N_14183,N_13648,N_13785);
nand U14184 (N_14184,N_13728,N_13299);
nand U14185 (N_14185,N_13340,N_13235);
nand U14186 (N_14186,N_13635,N_13675);
nand U14187 (N_14187,N_13231,N_13332);
xor U14188 (N_14188,N_13646,N_13522);
and U14189 (N_14189,N_13481,N_13711);
nand U14190 (N_14190,N_13654,N_13456);
nor U14191 (N_14191,N_13468,N_13728);
and U14192 (N_14192,N_13209,N_13549);
nor U14193 (N_14193,N_13731,N_13564);
nor U14194 (N_14194,N_13363,N_13365);
and U14195 (N_14195,N_13260,N_13756);
or U14196 (N_14196,N_13309,N_13262);
nor U14197 (N_14197,N_13383,N_13323);
or U14198 (N_14198,N_13686,N_13684);
or U14199 (N_14199,N_13460,N_13680);
nor U14200 (N_14200,N_13328,N_13303);
nor U14201 (N_14201,N_13223,N_13687);
xor U14202 (N_14202,N_13651,N_13203);
nor U14203 (N_14203,N_13716,N_13345);
xnor U14204 (N_14204,N_13726,N_13569);
xnor U14205 (N_14205,N_13241,N_13333);
and U14206 (N_14206,N_13692,N_13342);
nor U14207 (N_14207,N_13206,N_13364);
or U14208 (N_14208,N_13355,N_13427);
xor U14209 (N_14209,N_13229,N_13662);
or U14210 (N_14210,N_13315,N_13291);
nand U14211 (N_14211,N_13532,N_13653);
nor U14212 (N_14212,N_13345,N_13504);
nand U14213 (N_14213,N_13454,N_13733);
or U14214 (N_14214,N_13585,N_13362);
and U14215 (N_14215,N_13769,N_13531);
nor U14216 (N_14216,N_13208,N_13569);
and U14217 (N_14217,N_13361,N_13479);
xor U14218 (N_14218,N_13299,N_13375);
or U14219 (N_14219,N_13654,N_13302);
or U14220 (N_14220,N_13624,N_13216);
xnor U14221 (N_14221,N_13494,N_13651);
or U14222 (N_14222,N_13530,N_13729);
nor U14223 (N_14223,N_13311,N_13690);
and U14224 (N_14224,N_13480,N_13229);
or U14225 (N_14225,N_13739,N_13428);
xnor U14226 (N_14226,N_13773,N_13367);
or U14227 (N_14227,N_13709,N_13590);
nor U14228 (N_14228,N_13604,N_13373);
nand U14229 (N_14229,N_13227,N_13336);
xor U14230 (N_14230,N_13428,N_13769);
nand U14231 (N_14231,N_13347,N_13783);
xnor U14232 (N_14232,N_13225,N_13726);
and U14233 (N_14233,N_13472,N_13202);
nor U14234 (N_14234,N_13672,N_13343);
nand U14235 (N_14235,N_13534,N_13218);
nor U14236 (N_14236,N_13526,N_13492);
nand U14237 (N_14237,N_13461,N_13257);
or U14238 (N_14238,N_13598,N_13443);
xnor U14239 (N_14239,N_13429,N_13377);
nand U14240 (N_14240,N_13368,N_13700);
and U14241 (N_14241,N_13718,N_13390);
and U14242 (N_14242,N_13654,N_13548);
or U14243 (N_14243,N_13451,N_13433);
nand U14244 (N_14244,N_13725,N_13691);
or U14245 (N_14245,N_13403,N_13214);
nor U14246 (N_14246,N_13473,N_13256);
xor U14247 (N_14247,N_13750,N_13448);
xnor U14248 (N_14248,N_13441,N_13538);
nor U14249 (N_14249,N_13535,N_13796);
nand U14250 (N_14250,N_13397,N_13286);
or U14251 (N_14251,N_13535,N_13219);
nand U14252 (N_14252,N_13775,N_13450);
nand U14253 (N_14253,N_13768,N_13649);
nor U14254 (N_14254,N_13631,N_13704);
nand U14255 (N_14255,N_13635,N_13490);
nor U14256 (N_14256,N_13285,N_13531);
or U14257 (N_14257,N_13640,N_13255);
xor U14258 (N_14258,N_13534,N_13260);
nor U14259 (N_14259,N_13744,N_13721);
xor U14260 (N_14260,N_13304,N_13486);
xor U14261 (N_14261,N_13227,N_13471);
nor U14262 (N_14262,N_13427,N_13324);
nand U14263 (N_14263,N_13347,N_13544);
and U14264 (N_14264,N_13231,N_13630);
and U14265 (N_14265,N_13485,N_13213);
and U14266 (N_14266,N_13398,N_13367);
and U14267 (N_14267,N_13283,N_13216);
nor U14268 (N_14268,N_13743,N_13783);
and U14269 (N_14269,N_13602,N_13489);
nand U14270 (N_14270,N_13250,N_13742);
nor U14271 (N_14271,N_13247,N_13433);
or U14272 (N_14272,N_13693,N_13277);
and U14273 (N_14273,N_13434,N_13312);
nor U14274 (N_14274,N_13344,N_13751);
and U14275 (N_14275,N_13247,N_13565);
and U14276 (N_14276,N_13335,N_13548);
nor U14277 (N_14277,N_13492,N_13725);
xnor U14278 (N_14278,N_13281,N_13389);
xor U14279 (N_14279,N_13795,N_13530);
or U14280 (N_14280,N_13343,N_13529);
xor U14281 (N_14281,N_13287,N_13368);
xor U14282 (N_14282,N_13793,N_13235);
xnor U14283 (N_14283,N_13701,N_13500);
and U14284 (N_14284,N_13741,N_13604);
nor U14285 (N_14285,N_13346,N_13584);
xor U14286 (N_14286,N_13353,N_13486);
and U14287 (N_14287,N_13437,N_13342);
or U14288 (N_14288,N_13283,N_13754);
xnor U14289 (N_14289,N_13359,N_13786);
and U14290 (N_14290,N_13264,N_13608);
nor U14291 (N_14291,N_13348,N_13464);
and U14292 (N_14292,N_13436,N_13799);
xnor U14293 (N_14293,N_13361,N_13231);
and U14294 (N_14294,N_13523,N_13635);
or U14295 (N_14295,N_13635,N_13433);
xor U14296 (N_14296,N_13783,N_13421);
xnor U14297 (N_14297,N_13446,N_13599);
nor U14298 (N_14298,N_13645,N_13290);
or U14299 (N_14299,N_13452,N_13623);
and U14300 (N_14300,N_13369,N_13572);
and U14301 (N_14301,N_13610,N_13608);
nand U14302 (N_14302,N_13315,N_13312);
and U14303 (N_14303,N_13226,N_13732);
nor U14304 (N_14304,N_13438,N_13296);
nand U14305 (N_14305,N_13651,N_13643);
nand U14306 (N_14306,N_13372,N_13747);
or U14307 (N_14307,N_13760,N_13688);
nand U14308 (N_14308,N_13775,N_13741);
and U14309 (N_14309,N_13371,N_13535);
nand U14310 (N_14310,N_13378,N_13428);
and U14311 (N_14311,N_13519,N_13677);
or U14312 (N_14312,N_13710,N_13249);
xor U14313 (N_14313,N_13235,N_13234);
or U14314 (N_14314,N_13381,N_13609);
nor U14315 (N_14315,N_13312,N_13657);
and U14316 (N_14316,N_13555,N_13738);
xor U14317 (N_14317,N_13382,N_13349);
or U14318 (N_14318,N_13303,N_13744);
or U14319 (N_14319,N_13512,N_13663);
and U14320 (N_14320,N_13217,N_13595);
and U14321 (N_14321,N_13464,N_13760);
and U14322 (N_14322,N_13636,N_13770);
nand U14323 (N_14323,N_13672,N_13731);
nand U14324 (N_14324,N_13542,N_13743);
nand U14325 (N_14325,N_13492,N_13763);
and U14326 (N_14326,N_13549,N_13658);
and U14327 (N_14327,N_13309,N_13390);
nand U14328 (N_14328,N_13361,N_13653);
xnor U14329 (N_14329,N_13535,N_13299);
or U14330 (N_14330,N_13714,N_13687);
or U14331 (N_14331,N_13532,N_13250);
nand U14332 (N_14332,N_13342,N_13737);
nand U14333 (N_14333,N_13545,N_13578);
nand U14334 (N_14334,N_13380,N_13391);
xor U14335 (N_14335,N_13376,N_13434);
nor U14336 (N_14336,N_13313,N_13487);
and U14337 (N_14337,N_13365,N_13544);
nand U14338 (N_14338,N_13635,N_13748);
nand U14339 (N_14339,N_13694,N_13687);
or U14340 (N_14340,N_13230,N_13780);
nor U14341 (N_14341,N_13300,N_13634);
xnor U14342 (N_14342,N_13687,N_13522);
and U14343 (N_14343,N_13210,N_13576);
or U14344 (N_14344,N_13614,N_13318);
nand U14345 (N_14345,N_13522,N_13708);
nor U14346 (N_14346,N_13327,N_13306);
and U14347 (N_14347,N_13246,N_13484);
xor U14348 (N_14348,N_13509,N_13641);
xnor U14349 (N_14349,N_13629,N_13221);
xor U14350 (N_14350,N_13353,N_13739);
and U14351 (N_14351,N_13497,N_13701);
xnor U14352 (N_14352,N_13660,N_13497);
or U14353 (N_14353,N_13568,N_13618);
and U14354 (N_14354,N_13255,N_13738);
nor U14355 (N_14355,N_13539,N_13323);
nand U14356 (N_14356,N_13440,N_13264);
and U14357 (N_14357,N_13311,N_13364);
or U14358 (N_14358,N_13229,N_13267);
and U14359 (N_14359,N_13269,N_13714);
nor U14360 (N_14360,N_13701,N_13289);
nor U14361 (N_14361,N_13243,N_13603);
nor U14362 (N_14362,N_13297,N_13764);
or U14363 (N_14363,N_13708,N_13710);
or U14364 (N_14364,N_13761,N_13300);
nor U14365 (N_14365,N_13358,N_13780);
nor U14366 (N_14366,N_13356,N_13516);
and U14367 (N_14367,N_13650,N_13417);
xor U14368 (N_14368,N_13277,N_13234);
xor U14369 (N_14369,N_13642,N_13639);
xnor U14370 (N_14370,N_13539,N_13337);
and U14371 (N_14371,N_13298,N_13234);
and U14372 (N_14372,N_13514,N_13723);
and U14373 (N_14373,N_13666,N_13672);
xor U14374 (N_14374,N_13525,N_13322);
xnor U14375 (N_14375,N_13235,N_13502);
or U14376 (N_14376,N_13647,N_13228);
nand U14377 (N_14377,N_13675,N_13513);
and U14378 (N_14378,N_13323,N_13638);
and U14379 (N_14379,N_13312,N_13536);
or U14380 (N_14380,N_13512,N_13496);
or U14381 (N_14381,N_13679,N_13688);
and U14382 (N_14382,N_13359,N_13476);
nand U14383 (N_14383,N_13646,N_13376);
nor U14384 (N_14384,N_13555,N_13683);
nor U14385 (N_14385,N_13282,N_13368);
and U14386 (N_14386,N_13679,N_13315);
nor U14387 (N_14387,N_13731,N_13642);
xor U14388 (N_14388,N_13574,N_13218);
or U14389 (N_14389,N_13706,N_13303);
nand U14390 (N_14390,N_13618,N_13217);
and U14391 (N_14391,N_13706,N_13537);
and U14392 (N_14392,N_13475,N_13324);
or U14393 (N_14393,N_13775,N_13436);
nor U14394 (N_14394,N_13416,N_13396);
or U14395 (N_14395,N_13515,N_13756);
xnor U14396 (N_14396,N_13339,N_13471);
nor U14397 (N_14397,N_13638,N_13604);
nor U14398 (N_14398,N_13329,N_13395);
and U14399 (N_14399,N_13691,N_13615);
nor U14400 (N_14400,N_13846,N_14009);
and U14401 (N_14401,N_14119,N_14080);
or U14402 (N_14402,N_13947,N_14382);
nand U14403 (N_14403,N_13820,N_14127);
nor U14404 (N_14404,N_14308,N_14170);
nand U14405 (N_14405,N_13868,N_13922);
and U14406 (N_14406,N_14181,N_13978);
and U14407 (N_14407,N_14018,N_14258);
nor U14408 (N_14408,N_13936,N_14034);
nor U14409 (N_14409,N_13861,N_13984);
or U14410 (N_14410,N_13896,N_14073);
nand U14411 (N_14411,N_14147,N_14326);
or U14412 (N_14412,N_14105,N_14068);
xnor U14413 (N_14413,N_13893,N_14261);
and U14414 (N_14414,N_14302,N_13812);
xor U14415 (N_14415,N_14341,N_14265);
and U14416 (N_14416,N_14145,N_13874);
and U14417 (N_14417,N_14083,N_14195);
and U14418 (N_14418,N_14107,N_14182);
and U14419 (N_14419,N_14140,N_13917);
and U14420 (N_14420,N_14059,N_14088);
or U14421 (N_14421,N_13892,N_14081);
nor U14422 (N_14422,N_14006,N_13924);
and U14423 (N_14423,N_14180,N_13901);
nor U14424 (N_14424,N_13958,N_14362);
xnor U14425 (N_14425,N_14190,N_14040);
nor U14426 (N_14426,N_14257,N_14279);
and U14427 (N_14427,N_14373,N_14358);
and U14428 (N_14428,N_14020,N_14293);
and U14429 (N_14429,N_13983,N_14204);
and U14430 (N_14430,N_14220,N_14309);
and U14431 (N_14431,N_14199,N_14032);
or U14432 (N_14432,N_13835,N_14215);
nor U14433 (N_14433,N_14281,N_13905);
or U14434 (N_14434,N_14229,N_14338);
and U14435 (N_14435,N_14003,N_14061);
and U14436 (N_14436,N_14267,N_14234);
nand U14437 (N_14437,N_14075,N_14323);
nand U14438 (N_14438,N_14393,N_14208);
or U14439 (N_14439,N_13939,N_13944);
xor U14440 (N_14440,N_14375,N_14026);
and U14441 (N_14441,N_13921,N_14198);
or U14442 (N_14442,N_14014,N_14352);
xnor U14443 (N_14443,N_13994,N_13957);
xnor U14444 (N_14444,N_14178,N_13990);
xor U14445 (N_14445,N_14386,N_13996);
and U14446 (N_14446,N_13884,N_14113);
nor U14447 (N_14447,N_14380,N_13910);
or U14448 (N_14448,N_14310,N_14078);
nor U14449 (N_14449,N_14089,N_13841);
xor U14450 (N_14450,N_14112,N_13928);
nor U14451 (N_14451,N_14254,N_13906);
and U14452 (N_14452,N_14146,N_13977);
nand U14453 (N_14453,N_14346,N_14044);
and U14454 (N_14454,N_13887,N_14028);
nor U14455 (N_14455,N_13992,N_13987);
nor U14456 (N_14456,N_13946,N_14251);
or U14457 (N_14457,N_14128,N_14202);
and U14458 (N_14458,N_14102,N_13980);
or U14459 (N_14459,N_14176,N_14217);
nand U14460 (N_14460,N_14158,N_13995);
or U14461 (N_14461,N_14163,N_14104);
nand U14462 (N_14462,N_14086,N_14085);
xnor U14463 (N_14463,N_14242,N_14387);
or U14464 (N_14464,N_14067,N_14304);
and U14465 (N_14465,N_13930,N_14397);
nand U14466 (N_14466,N_14005,N_14046);
nand U14467 (N_14467,N_14138,N_13937);
xor U14468 (N_14468,N_14360,N_14218);
xnor U14469 (N_14469,N_13927,N_14070);
nand U14470 (N_14470,N_13981,N_14038);
or U14471 (N_14471,N_13989,N_13899);
nor U14472 (N_14472,N_13900,N_14134);
nor U14473 (N_14473,N_14303,N_14364);
xnor U14474 (N_14474,N_13865,N_14206);
nand U14475 (N_14475,N_14063,N_14290);
and U14476 (N_14476,N_14270,N_14335);
and U14477 (N_14477,N_13911,N_13869);
or U14478 (N_14478,N_13801,N_14137);
or U14479 (N_14479,N_14057,N_14378);
nor U14480 (N_14480,N_13964,N_14318);
xor U14481 (N_14481,N_13898,N_14351);
and U14482 (N_14482,N_13961,N_14191);
xnor U14483 (N_14483,N_14277,N_14203);
nor U14484 (N_14484,N_13864,N_13822);
xnor U14485 (N_14485,N_14065,N_13926);
and U14486 (N_14486,N_13965,N_14150);
or U14487 (N_14487,N_14355,N_14363);
nand U14488 (N_14488,N_14224,N_14374);
or U14489 (N_14489,N_14300,N_13837);
nor U14490 (N_14490,N_14384,N_14148);
xor U14491 (N_14491,N_14256,N_13971);
xor U14492 (N_14492,N_13832,N_14371);
nand U14493 (N_14493,N_14350,N_14359);
nor U14494 (N_14494,N_13918,N_13807);
xnor U14495 (N_14495,N_14398,N_13806);
and U14496 (N_14496,N_13848,N_13942);
nand U14497 (N_14497,N_13976,N_14247);
nand U14498 (N_14498,N_14072,N_13954);
nand U14499 (N_14499,N_14297,N_13882);
nor U14500 (N_14500,N_14275,N_13979);
and U14501 (N_14501,N_14154,N_14389);
or U14502 (N_14502,N_13952,N_13867);
and U14503 (N_14503,N_14238,N_13870);
nand U14504 (N_14504,N_14269,N_13823);
nor U14505 (N_14505,N_14311,N_14337);
nor U14506 (N_14506,N_14201,N_14285);
and U14507 (N_14507,N_14062,N_13903);
and U14508 (N_14508,N_14010,N_14211);
and U14509 (N_14509,N_14047,N_14241);
or U14510 (N_14510,N_14214,N_14016);
and U14511 (N_14511,N_14216,N_13804);
nor U14512 (N_14512,N_14174,N_14159);
nand U14513 (N_14513,N_13935,N_14298);
xnor U14514 (N_14514,N_14268,N_14106);
xnor U14515 (N_14515,N_13862,N_13969);
and U14516 (N_14516,N_13830,N_14319);
or U14517 (N_14517,N_13850,N_14109);
and U14518 (N_14518,N_14339,N_14054);
nand U14519 (N_14519,N_14200,N_13919);
xor U14520 (N_14520,N_14381,N_14278);
nor U14521 (N_14521,N_13908,N_14344);
nand U14522 (N_14522,N_13960,N_14291);
nand U14523 (N_14523,N_13950,N_13816);
nor U14524 (N_14524,N_14282,N_14263);
nor U14525 (N_14525,N_13933,N_13821);
nor U14526 (N_14526,N_13886,N_13888);
and U14527 (N_14527,N_13889,N_14160);
or U14528 (N_14528,N_14132,N_14139);
nand U14529 (N_14529,N_14192,N_14029);
xor U14530 (N_14530,N_14342,N_14025);
nand U14531 (N_14531,N_14307,N_14325);
xnor U14532 (N_14532,N_13897,N_13834);
xor U14533 (N_14533,N_14022,N_13902);
or U14534 (N_14534,N_14253,N_14124);
nor U14535 (N_14535,N_14076,N_14015);
nand U14536 (N_14536,N_14316,N_14324);
xnor U14537 (N_14537,N_14356,N_14354);
and U14538 (N_14538,N_13866,N_14071);
xor U14539 (N_14539,N_13951,N_13829);
and U14540 (N_14540,N_14141,N_14144);
nor U14541 (N_14541,N_14157,N_13854);
xnor U14542 (N_14542,N_14121,N_13907);
or U14543 (N_14543,N_13998,N_14276);
nor U14544 (N_14544,N_13940,N_14092);
and U14545 (N_14545,N_14314,N_14294);
xor U14546 (N_14546,N_14168,N_14011);
or U14547 (N_14547,N_13938,N_14236);
xor U14548 (N_14548,N_13883,N_14255);
nor U14549 (N_14549,N_14260,N_14343);
or U14550 (N_14550,N_14090,N_14097);
xnor U14551 (N_14551,N_14264,N_14039);
xor U14552 (N_14552,N_14126,N_13934);
nor U14553 (N_14553,N_14021,N_14051);
xor U14554 (N_14554,N_14019,N_14329);
or U14555 (N_14555,N_13827,N_13851);
xnor U14556 (N_14556,N_13811,N_14252);
xor U14557 (N_14557,N_13988,N_14055);
nand U14558 (N_14558,N_14185,N_14120);
nand U14559 (N_14559,N_14000,N_14289);
nand U14560 (N_14560,N_14230,N_14095);
and U14561 (N_14561,N_14162,N_14212);
nand U14562 (N_14562,N_13879,N_14012);
nor U14563 (N_14563,N_14049,N_14196);
and U14564 (N_14564,N_13858,N_14379);
or U14565 (N_14565,N_14004,N_14131);
nand U14566 (N_14566,N_14322,N_13813);
nor U14567 (N_14567,N_13904,N_13982);
nand U14568 (N_14568,N_14093,N_13844);
or U14569 (N_14569,N_14395,N_14396);
nand U14570 (N_14570,N_13878,N_14328);
xnor U14571 (N_14571,N_14243,N_13912);
nor U14572 (N_14572,N_13941,N_14233);
nand U14573 (N_14573,N_14228,N_14287);
xor U14574 (N_14574,N_14272,N_14094);
and U14575 (N_14575,N_13973,N_14222);
or U14576 (N_14576,N_13929,N_13817);
nor U14577 (N_14577,N_14111,N_13856);
xnor U14578 (N_14578,N_14353,N_14262);
nand U14579 (N_14579,N_14052,N_14114);
nand U14580 (N_14580,N_13859,N_13920);
nand U14581 (N_14581,N_14245,N_14183);
and U14582 (N_14582,N_14171,N_14271);
nor U14583 (N_14583,N_14388,N_13819);
xor U14584 (N_14584,N_14266,N_14286);
nor U14585 (N_14585,N_14315,N_14048);
and U14586 (N_14586,N_14177,N_13809);
and U14587 (N_14587,N_14249,N_13860);
nor U14588 (N_14588,N_13909,N_14292);
or U14589 (N_14589,N_13831,N_13845);
nor U14590 (N_14590,N_14161,N_13839);
nand U14591 (N_14591,N_13842,N_14227);
or U14592 (N_14592,N_14226,N_13828);
and U14593 (N_14593,N_14349,N_14184);
nor U14594 (N_14594,N_14098,N_14060);
nor U14595 (N_14595,N_14017,N_13815);
or U14596 (N_14596,N_14152,N_14207);
or U14597 (N_14597,N_14041,N_14327);
nand U14598 (N_14598,N_14301,N_13852);
and U14599 (N_14599,N_13974,N_13853);
or U14600 (N_14600,N_13955,N_13914);
and U14601 (N_14601,N_14317,N_14099);
or U14602 (N_14602,N_13931,N_14074);
nor U14603 (N_14603,N_14125,N_13814);
xor U14604 (N_14604,N_14117,N_14035);
xor U14605 (N_14605,N_14295,N_13999);
nor U14606 (N_14606,N_14248,N_14246);
nand U14607 (N_14607,N_13833,N_13915);
xor U14608 (N_14608,N_13803,N_14084);
nor U14609 (N_14609,N_13962,N_13953);
or U14610 (N_14610,N_14340,N_14164);
nand U14611 (N_14611,N_13824,N_14232);
nor U14612 (N_14612,N_14205,N_14115);
xnor U14613 (N_14613,N_14066,N_14149);
xnor U14614 (N_14614,N_13932,N_14288);
nor U14615 (N_14615,N_13967,N_13838);
and U14616 (N_14616,N_14299,N_14188);
or U14617 (N_14617,N_14024,N_14219);
nand U14618 (N_14618,N_14077,N_14116);
nand U14619 (N_14619,N_14284,N_14053);
nor U14620 (N_14620,N_13836,N_14320);
and U14621 (N_14621,N_13948,N_13891);
nand U14622 (N_14622,N_14347,N_14331);
or U14623 (N_14623,N_14333,N_14091);
nand U14624 (N_14624,N_14033,N_13959);
nor U14625 (N_14625,N_14175,N_13968);
or U14626 (N_14626,N_14274,N_14332);
and U14627 (N_14627,N_13805,N_13877);
xnor U14628 (N_14628,N_14122,N_13881);
or U14629 (N_14629,N_13970,N_14280);
xnor U14630 (N_14630,N_14187,N_13855);
nor U14631 (N_14631,N_14151,N_14305);
nor U14632 (N_14632,N_13949,N_14377);
or U14633 (N_14633,N_14036,N_14330);
nand U14634 (N_14634,N_14365,N_14166);
nand U14635 (N_14635,N_13847,N_14259);
and U14636 (N_14636,N_14213,N_14167);
nand U14637 (N_14637,N_14399,N_14394);
and U14638 (N_14638,N_13956,N_14273);
and U14639 (N_14639,N_13843,N_13875);
nand U14640 (N_14640,N_13871,N_14334);
nor U14641 (N_14641,N_14096,N_13945);
and U14642 (N_14642,N_14156,N_14194);
or U14643 (N_14643,N_13997,N_14002);
nand U14644 (N_14644,N_14361,N_14345);
xor U14645 (N_14645,N_14013,N_13923);
xor U14646 (N_14646,N_14237,N_14186);
and U14647 (N_14647,N_14296,N_14133);
nand U14648 (N_14648,N_14129,N_13800);
nand U14649 (N_14649,N_14313,N_13890);
and U14650 (N_14650,N_14225,N_14110);
nand U14651 (N_14651,N_14143,N_14123);
nor U14652 (N_14652,N_14357,N_14042);
or U14653 (N_14653,N_14169,N_13925);
xnor U14654 (N_14654,N_14197,N_13876);
nor U14655 (N_14655,N_14058,N_13895);
xor U14656 (N_14656,N_14108,N_14008);
or U14657 (N_14657,N_14250,N_14221);
xnor U14658 (N_14658,N_13849,N_14142);
xor U14659 (N_14659,N_14372,N_13802);
or U14660 (N_14660,N_14189,N_13885);
and U14661 (N_14661,N_14101,N_14385);
nand U14662 (N_14662,N_14064,N_14179);
nand U14663 (N_14663,N_13894,N_14045);
xnor U14664 (N_14664,N_14173,N_13916);
nor U14665 (N_14665,N_14321,N_14235);
nand U14666 (N_14666,N_14239,N_14336);
nor U14667 (N_14667,N_14366,N_14136);
or U14668 (N_14668,N_14223,N_14370);
and U14669 (N_14669,N_14240,N_14348);
xor U14670 (N_14670,N_13826,N_14135);
or U14671 (N_14671,N_14390,N_13825);
or U14672 (N_14672,N_14031,N_14376);
xor U14673 (N_14673,N_14155,N_13986);
or U14674 (N_14674,N_13857,N_14079);
or U14675 (N_14675,N_14210,N_13840);
nor U14676 (N_14676,N_14118,N_13880);
xnor U14677 (N_14677,N_13943,N_14368);
and U14678 (N_14678,N_14392,N_14369);
nand U14679 (N_14679,N_14209,N_14367);
or U14680 (N_14680,N_14001,N_14069);
xnor U14681 (N_14681,N_14027,N_13963);
and U14682 (N_14682,N_13993,N_14306);
or U14683 (N_14683,N_13966,N_13975);
nor U14684 (N_14684,N_14153,N_13863);
nand U14685 (N_14685,N_13810,N_13972);
or U14686 (N_14686,N_14037,N_14100);
nand U14687 (N_14687,N_13985,N_14007);
nor U14688 (N_14688,N_13913,N_14043);
xor U14689 (N_14689,N_14103,N_14082);
nor U14690 (N_14690,N_14050,N_14165);
nor U14691 (N_14691,N_13808,N_14130);
and U14692 (N_14692,N_13872,N_14283);
and U14693 (N_14693,N_14172,N_14087);
and U14694 (N_14694,N_14023,N_14193);
or U14695 (N_14695,N_13991,N_13873);
nand U14696 (N_14696,N_14056,N_13818);
xor U14697 (N_14697,N_14030,N_14231);
xnor U14698 (N_14698,N_14391,N_14244);
and U14699 (N_14699,N_14383,N_14312);
nor U14700 (N_14700,N_14171,N_13836);
nor U14701 (N_14701,N_13929,N_13956);
nand U14702 (N_14702,N_14185,N_14228);
xor U14703 (N_14703,N_14376,N_14017);
nand U14704 (N_14704,N_13810,N_14023);
and U14705 (N_14705,N_14329,N_13973);
xnor U14706 (N_14706,N_13904,N_14113);
xor U14707 (N_14707,N_14321,N_13929);
or U14708 (N_14708,N_14397,N_14040);
nand U14709 (N_14709,N_14097,N_14065);
nor U14710 (N_14710,N_13959,N_14387);
nor U14711 (N_14711,N_14269,N_14165);
and U14712 (N_14712,N_14181,N_14302);
nand U14713 (N_14713,N_14344,N_14176);
and U14714 (N_14714,N_14315,N_14310);
or U14715 (N_14715,N_14392,N_14174);
xnor U14716 (N_14716,N_14108,N_13990);
nand U14717 (N_14717,N_13959,N_14346);
or U14718 (N_14718,N_14349,N_13884);
nor U14719 (N_14719,N_13800,N_14183);
xor U14720 (N_14720,N_14388,N_14166);
or U14721 (N_14721,N_13936,N_14371);
nor U14722 (N_14722,N_14092,N_13870);
nor U14723 (N_14723,N_14135,N_13858);
nand U14724 (N_14724,N_14398,N_14216);
xor U14725 (N_14725,N_14324,N_14180);
and U14726 (N_14726,N_14008,N_13898);
nand U14727 (N_14727,N_14129,N_14016);
xnor U14728 (N_14728,N_14103,N_14206);
xor U14729 (N_14729,N_14296,N_14327);
xor U14730 (N_14730,N_14025,N_14345);
nor U14731 (N_14731,N_14392,N_14393);
and U14732 (N_14732,N_14221,N_14043);
nor U14733 (N_14733,N_14344,N_14320);
and U14734 (N_14734,N_13943,N_14171);
nand U14735 (N_14735,N_14129,N_14137);
nor U14736 (N_14736,N_13842,N_14104);
nor U14737 (N_14737,N_14142,N_14276);
nor U14738 (N_14738,N_14339,N_14147);
and U14739 (N_14739,N_14308,N_13817);
nand U14740 (N_14740,N_14252,N_14284);
xnor U14741 (N_14741,N_14005,N_14337);
and U14742 (N_14742,N_14175,N_14119);
nand U14743 (N_14743,N_13970,N_14202);
nor U14744 (N_14744,N_13989,N_13923);
or U14745 (N_14745,N_13825,N_13840);
and U14746 (N_14746,N_13854,N_14295);
nand U14747 (N_14747,N_14140,N_14305);
and U14748 (N_14748,N_14327,N_14225);
nand U14749 (N_14749,N_14202,N_14264);
nor U14750 (N_14750,N_13939,N_14283);
nand U14751 (N_14751,N_14272,N_14343);
nor U14752 (N_14752,N_14363,N_14378);
xnor U14753 (N_14753,N_14036,N_14286);
and U14754 (N_14754,N_14036,N_13986);
nand U14755 (N_14755,N_13860,N_14312);
xor U14756 (N_14756,N_13885,N_14396);
and U14757 (N_14757,N_14046,N_14244);
nand U14758 (N_14758,N_14163,N_14135);
nand U14759 (N_14759,N_14246,N_14147);
nor U14760 (N_14760,N_14360,N_13993);
nand U14761 (N_14761,N_14255,N_14053);
or U14762 (N_14762,N_13982,N_14133);
nand U14763 (N_14763,N_14026,N_14148);
and U14764 (N_14764,N_14205,N_14011);
and U14765 (N_14765,N_13955,N_13939);
and U14766 (N_14766,N_14372,N_14230);
or U14767 (N_14767,N_14172,N_14352);
nor U14768 (N_14768,N_13822,N_14063);
xor U14769 (N_14769,N_13986,N_14245);
and U14770 (N_14770,N_14343,N_14132);
nor U14771 (N_14771,N_13903,N_13872);
and U14772 (N_14772,N_14381,N_14298);
or U14773 (N_14773,N_13970,N_14176);
and U14774 (N_14774,N_14085,N_13929);
xnor U14775 (N_14775,N_14184,N_14363);
and U14776 (N_14776,N_14128,N_13958);
nand U14777 (N_14777,N_14125,N_14143);
nand U14778 (N_14778,N_14367,N_14286);
nand U14779 (N_14779,N_13824,N_14156);
or U14780 (N_14780,N_14205,N_14066);
xor U14781 (N_14781,N_13829,N_14154);
nand U14782 (N_14782,N_14363,N_14117);
nand U14783 (N_14783,N_14342,N_13890);
xor U14784 (N_14784,N_14355,N_14127);
nor U14785 (N_14785,N_14360,N_13893);
or U14786 (N_14786,N_14397,N_14069);
nor U14787 (N_14787,N_14229,N_13834);
nor U14788 (N_14788,N_14106,N_14082);
nor U14789 (N_14789,N_14323,N_14267);
xnor U14790 (N_14790,N_14173,N_14018);
or U14791 (N_14791,N_14066,N_14085);
nor U14792 (N_14792,N_14307,N_14111);
xor U14793 (N_14793,N_13840,N_14279);
or U14794 (N_14794,N_14123,N_13824);
xor U14795 (N_14795,N_13970,N_14246);
xnor U14796 (N_14796,N_14307,N_14221);
nand U14797 (N_14797,N_13870,N_14013);
nand U14798 (N_14798,N_14190,N_14159);
or U14799 (N_14799,N_14202,N_13994);
nand U14800 (N_14800,N_14155,N_13917);
nor U14801 (N_14801,N_13820,N_14054);
nor U14802 (N_14802,N_14047,N_14104);
and U14803 (N_14803,N_13929,N_14098);
nor U14804 (N_14804,N_13866,N_14109);
or U14805 (N_14805,N_13988,N_14186);
nand U14806 (N_14806,N_13878,N_14038);
nand U14807 (N_14807,N_14065,N_13826);
or U14808 (N_14808,N_13953,N_14334);
nand U14809 (N_14809,N_14327,N_14365);
nor U14810 (N_14810,N_13936,N_14053);
xnor U14811 (N_14811,N_13877,N_14240);
and U14812 (N_14812,N_14153,N_13932);
nand U14813 (N_14813,N_13882,N_13952);
or U14814 (N_14814,N_14349,N_13977);
xor U14815 (N_14815,N_14082,N_14036);
xnor U14816 (N_14816,N_14142,N_14150);
nand U14817 (N_14817,N_14325,N_14258);
nor U14818 (N_14818,N_14002,N_14185);
xnor U14819 (N_14819,N_14067,N_13885);
nor U14820 (N_14820,N_13936,N_14220);
nor U14821 (N_14821,N_14063,N_13809);
and U14822 (N_14822,N_14253,N_13971);
nor U14823 (N_14823,N_14134,N_14278);
nand U14824 (N_14824,N_14286,N_13891);
or U14825 (N_14825,N_14344,N_14202);
and U14826 (N_14826,N_14207,N_14030);
and U14827 (N_14827,N_13913,N_14235);
xor U14828 (N_14828,N_14085,N_14194);
nand U14829 (N_14829,N_14339,N_14012);
nand U14830 (N_14830,N_13932,N_13975);
nand U14831 (N_14831,N_13810,N_13905);
or U14832 (N_14832,N_13830,N_14302);
or U14833 (N_14833,N_14105,N_14328);
xnor U14834 (N_14834,N_14246,N_14081);
and U14835 (N_14835,N_13833,N_14181);
and U14836 (N_14836,N_14162,N_14236);
and U14837 (N_14837,N_13910,N_13971);
or U14838 (N_14838,N_14198,N_14009);
nand U14839 (N_14839,N_14337,N_13839);
xor U14840 (N_14840,N_14314,N_14000);
or U14841 (N_14841,N_14173,N_14272);
nand U14842 (N_14842,N_13886,N_14214);
nor U14843 (N_14843,N_14162,N_14142);
xor U14844 (N_14844,N_14343,N_14308);
nor U14845 (N_14845,N_14143,N_14016);
or U14846 (N_14846,N_14283,N_13807);
or U14847 (N_14847,N_13803,N_14196);
nand U14848 (N_14848,N_14267,N_13881);
nand U14849 (N_14849,N_14396,N_13861);
and U14850 (N_14850,N_14150,N_14202);
or U14851 (N_14851,N_14282,N_14225);
or U14852 (N_14852,N_14221,N_14359);
nor U14853 (N_14853,N_13881,N_14369);
nor U14854 (N_14854,N_14229,N_14350);
xor U14855 (N_14855,N_14199,N_14248);
nor U14856 (N_14856,N_14160,N_13994);
nor U14857 (N_14857,N_13871,N_14176);
nor U14858 (N_14858,N_14223,N_14103);
or U14859 (N_14859,N_14144,N_14378);
and U14860 (N_14860,N_13946,N_14223);
and U14861 (N_14861,N_13992,N_13883);
xnor U14862 (N_14862,N_14316,N_13914);
xnor U14863 (N_14863,N_13878,N_14101);
nor U14864 (N_14864,N_14296,N_14078);
nor U14865 (N_14865,N_14063,N_13827);
xor U14866 (N_14866,N_14087,N_14325);
xnor U14867 (N_14867,N_14057,N_14284);
nand U14868 (N_14868,N_13988,N_13975);
xnor U14869 (N_14869,N_14105,N_14383);
nor U14870 (N_14870,N_13889,N_13846);
xnor U14871 (N_14871,N_14336,N_13901);
nand U14872 (N_14872,N_13816,N_14008);
and U14873 (N_14873,N_14223,N_14035);
xnor U14874 (N_14874,N_14056,N_13934);
xnor U14875 (N_14875,N_14063,N_13953);
nor U14876 (N_14876,N_14348,N_14354);
xnor U14877 (N_14877,N_14115,N_13854);
nand U14878 (N_14878,N_13955,N_14003);
and U14879 (N_14879,N_14289,N_13864);
nand U14880 (N_14880,N_14130,N_14161);
nor U14881 (N_14881,N_13928,N_14372);
or U14882 (N_14882,N_14124,N_13836);
nor U14883 (N_14883,N_14358,N_14208);
xnor U14884 (N_14884,N_13968,N_14145);
or U14885 (N_14885,N_14204,N_14207);
xnor U14886 (N_14886,N_14007,N_13855);
and U14887 (N_14887,N_14099,N_14041);
and U14888 (N_14888,N_13822,N_13949);
xor U14889 (N_14889,N_14357,N_13803);
or U14890 (N_14890,N_14223,N_14336);
nand U14891 (N_14891,N_13824,N_14136);
and U14892 (N_14892,N_14365,N_14359);
and U14893 (N_14893,N_14270,N_14331);
nand U14894 (N_14894,N_14210,N_13913);
nor U14895 (N_14895,N_13978,N_14101);
and U14896 (N_14896,N_13837,N_13918);
or U14897 (N_14897,N_14286,N_14053);
nand U14898 (N_14898,N_14303,N_13962);
and U14899 (N_14899,N_13803,N_14033);
xnor U14900 (N_14900,N_14010,N_13814);
or U14901 (N_14901,N_14067,N_14330);
xor U14902 (N_14902,N_14318,N_14105);
xnor U14903 (N_14903,N_14064,N_13983);
xor U14904 (N_14904,N_14110,N_13969);
nand U14905 (N_14905,N_13857,N_13982);
xnor U14906 (N_14906,N_13930,N_14305);
and U14907 (N_14907,N_14303,N_14105);
nor U14908 (N_14908,N_13961,N_14263);
xor U14909 (N_14909,N_14178,N_14360);
nor U14910 (N_14910,N_14366,N_13971);
and U14911 (N_14911,N_14094,N_14266);
nand U14912 (N_14912,N_14263,N_13805);
and U14913 (N_14913,N_14014,N_14230);
nand U14914 (N_14914,N_13862,N_13922);
or U14915 (N_14915,N_14302,N_14177);
xor U14916 (N_14916,N_13947,N_14272);
xor U14917 (N_14917,N_14280,N_14392);
or U14918 (N_14918,N_13892,N_13997);
and U14919 (N_14919,N_14097,N_13956);
or U14920 (N_14920,N_14171,N_13831);
xnor U14921 (N_14921,N_13853,N_13891);
and U14922 (N_14922,N_14150,N_14101);
xor U14923 (N_14923,N_13816,N_14253);
nand U14924 (N_14924,N_14157,N_14369);
nand U14925 (N_14925,N_14140,N_14180);
xor U14926 (N_14926,N_13920,N_13917);
and U14927 (N_14927,N_14212,N_14065);
nand U14928 (N_14928,N_14187,N_13842);
nor U14929 (N_14929,N_14384,N_13888);
and U14930 (N_14930,N_13917,N_14195);
and U14931 (N_14931,N_13914,N_13907);
and U14932 (N_14932,N_13988,N_14236);
or U14933 (N_14933,N_14327,N_14223);
and U14934 (N_14934,N_14164,N_13979);
nand U14935 (N_14935,N_14309,N_14181);
xor U14936 (N_14936,N_14188,N_14321);
or U14937 (N_14937,N_14277,N_14260);
nand U14938 (N_14938,N_14327,N_14120);
nor U14939 (N_14939,N_14346,N_13936);
nor U14940 (N_14940,N_14336,N_13942);
xnor U14941 (N_14941,N_14094,N_13837);
nor U14942 (N_14942,N_13930,N_14357);
nand U14943 (N_14943,N_13954,N_14021);
and U14944 (N_14944,N_14025,N_13831);
or U14945 (N_14945,N_13975,N_14290);
or U14946 (N_14946,N_14098,N_13953);
nand U14947 (N_14947,N_14012,N_14381);
xnor U14948 (N_14948,N_14010,N_14113);
nor U14949 (N_14949,N_14027,N_14197);
and U14950 (N_14950,N_14132,N_14257);
xor U14951 (N_14951,N_14194,N_14167);
nor U14952 (N_14952,N_13857,N_13824);
nand U14953 (N_14953,N_14054,N_14103);
nor U14954 (N_14954,N_14038,N_14302);
nor U14955 (N_14955,N_14187,N_13931);
xnor U14956 (N_14956,N_13962,N_14256);
xor U14957 (N_14957,N_14231,N_14073);
nor U14958 (N_14958,N_13921,N_14112);
xor U14959 (N_14959,N_14155,N_13831);
nand U14960 (N_14960,N_14134,N_14091);
or U14961 (N_14961,N_13930,N_14129);
or U14962 (N_14962,N_14029,N_14276);
and U14963 (N_14963,N_13821,N_13836);
or U14964 (N_14964,N_14189,N_13891);
and U14965 (N_14965,N_14349,N_13974);
nor U14966 (N_14966,N_13911,N_14230);
and U14967 (N_14967,N_14253,N_14223);
or U14968 (N_14968,N_14142,N_13969);
xnor U14969 (N_14969,N_14330,N_13818);
or U14970 (N_14970,N_14132,N_14381);
nor U14971 (N_14971,N_14276,N_14041);
nand U14972 (N_14972,N_13921,N_14328);
xor U14973 (N_14973,N_13997,N_13960);
nand U14974 (N_14974,N_14207,N_14250);
nor U14975 (N_14975,N_14336,N_13858);
xor U14976 (N_14976,N_13896,N_13865);
or U14977 (N_14977,N_14060,N_14314);
and U14978 (N_14978,N_14225,N_14024);
nand U14979 (N_14979,N_13893,N_14024);
or U14980 (N_14980,N_14137,N_14296);
nand U14981 (N_14981,N_13860,N_13902);
or U14982 (N_14982,N_13863,N_13987);
and U14983 (N_14983,N_13941,N_14002);
nor U14984 (N_14984,N_14198,N_14203);
or U14985 (N_14985,N_13861,N_14148);
nor U14986 (N_14986,N_14247,N_13952);
nand U14987 (N_14987,N_13984,N_13942);
and U14988 (N_14988,N_13822,N_14306);
or U14989 (N_14989,N_14042,N_14135);
nand U14990 (N_14990,N_14131,N_13980);
or U14991 (N_14991,N_14267,N_14097);
xor U14992 (N_14992,N_13822,N_14023);
xor U14993 (N_14993,N_14155,N_14107);
nand U14994 (N_14994,N_14050,N_13815);
nand U14995 (N_14995,N_13999,N_14232);
nor U14996 (N_14996,N_13811,N_14231);
or U14997 (N_14997,N_14110,N_13887);
nand U14998 (N_14998,N_14240,N_14250);
or U14999 (N_14999,N_14116,N_14080);
nand U15000 (N_15000,N_14913,N_14478);
nand U15001 (N_15001,N_14719,N_14867);
or U15002 (N_15002,N_14927,N_14653);
xnor U15003 (N_15003,N_14412,N_14556);
nor U15004 (N_15004,N_14744,N_14861);
xor U15005 (N_15005,N_14905,N_14696);
or U15006 (N_15006,N_14536,N_14651);
xor U15007 (N_15007,N_14843,N_14729);
xnor U15008 (N_15008,N_14438,N_14720);
xnor U15009 (N_15009,N_14740,N_14544);
nand U15010 (N_15010,N_14683,N_14659);
nand U15011 (N_15011,N_14496,N_14755);
nor U15012 (N_15012,N_14912,N_14992);
nor U15013 (N_15013,N_14917,N_14459);
or U15014 (N_15014,N_14858,N_14789);
nor U15015 (N_15015,N_14874,N_14838);
or U15016 (N_15016,N_14649,N_14797);
nand U15017 (N_15017,N_14497,N_14673);
nor U15018 (N_15018,N_14460,N_14884);
or U15019 (N_15019,N_14689,N_14569);
xnor U15020 (N_15020,N_14875,N_14699);
nand U15021 (N_15021,N_14507,N_14490);
and U15022 (N_15022,N_14816,N_14805);
or U15023 (N_15023,N_14603,N_14606);
nand U15024 (N_15024,N_14563,N_14523);
or U15025 (N_15025,N_14517,N_14648);
nand U15026 (N_15026,N_14510,N_14627);
xor U15027 (N_15027,N_14964,N_14535);
nand U15028 (N_15028,N_14582,N_14831);
nand U15029 (N_15029,N_14586,N_14423);
or U15030 (N_15030,N_14567,N_14574);
nand U15031 (N_15031,N_14531,N_14732);
nand U15032 (N_15032,N_14897,N_14773);
nand U15033 (N_15033,N_14753,N_14401);
xnor U15034 (N_15034,N_14770,N_14962);
nand U15035 (N_15035,N_14443,N_14887);
nand U15036 (N_15036,N_14489,N_14738);
nor U15037 (N_15037,N_14709,N_14849);
nand U15038 (N_15038,N_14585,N_14487);
nand U15039 (N_15039,N_14940,N_14982);
nor U15040 (N_15040,N_14868,N_14988);
and U15041 (N_15041,N_14522,N_14555);
nor U15042 (N_15042,N_14949,N_14617);
or U15043 (N_15043,N_14420,N_14519);
nor U15044 (N_15044,N_14691,N_14958);
and U15045 (N_15045,N_14652,N_14532);
nand U15046 (N_15046,N_14749,N_14469);
xor U15047 (N_15047,N_14939,N_14655);
xnor U15048 (N_15048,N_14971,N_14739);
and U15049 (N_15049,N_14752,N_14710);
nand U15050 (N_15050,N_14508,N_14952);
or U15051 (N_15051,N_14869,N_14641);
nand U15052 (N_15052,N_14981,N_14626);
nand U15053 (N_15053,N_14933,N_14860);
nand U15054 (N_15054,N_14456,N_14803);
and U15055 (N_15055,N_14424,N_14985);
nor U15056 (N_15056,N_14845,N_14801);
nor U15057 (N_15057,N_14724,N_14533);
or U15058 (N_15058,N_14785,N_14698);
or U15059 (N_15059,N_14560,N_14577);
nand U15060 (N_15060,N_14511,N_14764);
nor U15061 (N_15061,N_14421,N_14942);
xnor U15062 (N_15062,N_14414,N_14928);
and U15063 (N_15063,N_14473,N_14837);
xnor U15064 (N_15064,N_14904,N_14453);
xnor U15065 (N_15065,N_14468,N_14976);
xor U15066 (N_15066,N_14993,N_14754);
and U15067 (N_15067,N_14614,N_14591);
nand U15068 (N_15068,N_14442,N_14911);
xnor U15069 (N_15069,N_14483,N_14636);
or U15070 (N_15070,N_14945,N_14813);
nand U15071 (N_15071,N_14937,N_14891);
and U15072 (N_15072,N_14629,N_14778);
xnor U15073 (N_15073,N_14598,N_14712);
xor U15074 (N_15074,N_14642,N_14678);
xor U15075 (N_15075,N_14955,N_14656);
xor U15076 (N_15076,N_14650,N_14668);
nor U15077 (N_15077,N_14611,N_14704);
xor U15078 (N_15078,N_14824,N_14812);
xor U15079 (N_15079,N_14429,N_14640);
or U15080 (N_15080,N_14920,N_14925);
or U15081 (N_15081,N_14624,N_14736);
and U15082 (N_15082,N_14675,N_14903);
nand U15083 (N_15083,N_14944,N_14610);
and U15084 (N_15084,N_14883,N_14494);
or U15085 (N_15085,N_14609,N_14746);
nand U15086 (N_15086,N_14996,N_14514);
xor U15087 (N_15087,N_14408,N_14737);
xnor U15088 (N_15088,N_14714,N_14934);
nand U15089 (N_15089,N_14593,N_14743);
nand U15090 (N_15090,N_14440,N_14432);
and U15091 (N_15091,N_14758,N_14476);
or U15092 (N_15092,N_14500,N_14692);
nor U15093 (N_15093,N_14503,N_14924);
or U15094 (N_15094,N_14428,N_14763);
and U15095 (N_15095,N_14788,N_14674);
and U15096 (N_15096,N_14427,N_14597);
or U15097 (N_15097,N_14833,N_14879);
and U15098 (N_15098,N_14807,N_14757);
or U15099 (N_15099,N_14534,N_14774);
and U15100 (N_15100,N_14791,N_14465);
and U15101 (N_15101,N_14660,N_14618);
xor U15102 (N_15102,N_14454,N_14841);
or U15103 (N_15103,N_14926,N_14576);
nand U15104 (N_15104,N_14447,N_14956);
nand U15105 (N_15105,N_14422,N_14847);
and U15106 (N_15106,N_14592,N_14931);
xnor U15107 (N_15107,N_14516,N_14784);
xor U15108 (N_15108,N_14446,N_14747);
nand U15109 (N_15109,N_14644,N_14581);
or U15110 (N_15110,N_14608,N_14594);
nor U15111 (N_15111,N_14915,N_14681);
nor U15112 (N_15112,N_14458,N_14863);
and U15113 (N_15113,N_14679,N_14492);
or U15114 (N_15114,N_14589,N_14717);
or U15115 (N_15115,N_14495,N_14639);
and U15116 (N_15116,N_14471,N_14938);
xnor U15117 (N_15117,N_14530,N_14777);
and U15118 (N_15118,N_14413,N_14768);
or U15119 (N_15119,N_14596,N_14405);
or U15120 (N_15120,N_14526,N_14448);
nor U15121 (N_15121,N_14916,N_14584);
or U15122 (N_15122,N_14467,N_14799);
and U15123 (N_15123,N_14782,N_14781);
nand U15124 (N_15124,N_14703,N_14595);
or U15125 (N_15125,N_14557,N_14669);
nand U15126 (N_15126,N_14930,N_14987);
and U15127 (N_15127,N_14546,N_14578);
and U15128 (N_15128,N_14880,N_14735);
xor U15129 (N_15129,N_14866,N_14960);
nor U15130 (N_15130,N_14551,N_14607);
nor U15131 (N_15131,N_14549,N_14929);
and U15132 (N_15132,N_14646,N_14728);
nor U15133 (N_15133,N_14482,N_14452);
nor U15134 (N_15134,N_14707,N_14457);
and U15135 (N_15135,N_14829,N_14936);
or U15136 (N_15136,N_14579,N_14979);
and U15137 (N_15137,N_14525,N_14485);
xor U15138 (N_15138,N_14426,N_14750);
xnor U15139 (N_15139,N_14628,N_14463);
or U15140 (N_15140,N_14434,N_14910);
and U15141 (N_15141,N_14984,N_14695);
nor U15142 (N_15142,N_14435,N_14455);
or U15143 (N_15143,N_14715,N_14632);
xor U15144 (N_15144,N_14999,N_14643);
nand U15145 (N_15145,N_14889,N_14658);
and U15146 (N_15146,N_14721,N_14499);
and U15147 (N_15147,N_14769,N_14986);
nand U15148 (N_15148,N_14852,N_14767);
or U15149 (N_15149,N_14786,N_14705);
and U15150 (N_15150,N_14878,N_14436);
and U15151 (N_15151,N_14980,N_14590);
and U15152 (N_15152,N_14919,N_14765);
xor U15153 (N_15153,N_14561,N_14663);
nand U15154 (N_15154,N_14780,N_14848);
or U15155 (N_15155,N_14521,N_14825);
and U15156 (N_15156,N_14921,N_14951);
and U15157 (N_15157,N_14545,N_14893);
xnor U15158 (N_15158,N_14872,N_14991);
or U15159 (N_15159,N_14504,N_14621);
xor U15160 (N_15160,N_14711,N_14882);
or U15161 (N_15161,N_14842,N_14451);
nor U15162 (N_15162,N_14994,N_14548);
xnor U15163 (N_15163,N_14437,N_14898);
xnor U15164 (N_15164,N_14792,N_14954);
nand U15165 (N_15165,N_14515,N_14672);
xnor U15166 (N_15166,N_14961,N_14760);
nand U15167 (N_15167,N_14580,N_14706);
xor U15168 (N_15168,N_14409,N_14685);
or U15169 (N_15169,N_14832,N_14505);
xor U15170 (N_15170,N_14885,N_14725);
nor U15171 (N_15171,N_14493,N_14562);
or U15172 (N_15172,N_14851,N_14439);
or U15173 (N_15173,N_14795,N_14967);
nor U15174 (N_15174,N_14509,N_14989);
or U15175 (N_15175,N_14664,N_14620);
or U15176 (N_15176,N_14756,N_14701);
and U15177 (N_15177,N_14470,N_14968);
or U15178 (N_15178,N_14901,N_14821);
or U15179 (N_15179,N_14722,N_14430);
and U15180 (N_15180,N_14730,N_14759);
xnor U15181 (N_15181,N_14486,N_14498);
nor U15182 (N_15182,N_14894,N_14524);
xor U15183 (N_15183,N_14700,N_14550);
xnor U15184 (N_15184,N_14464,N_14957);
nor U15185 (N_15185,N_14941,N_14900);
xnor U15186 (N_15186,N_14990,N_14631);
and U15187 (N_15187,N_14793,N_14539);
and U15188 (N_15188,N_14932,N_14892);
and U15189 (N_15189,N_14873,N_14566);
nand U15190 (N_15190,N_14601,N_14572);
nor U15191 (N_15191,N_14416,N_14906);
nand U15192 (N_15192,N_14823,N_14977);
nand U15193 (N_15193,N_14479,N_14881);
and U15194 (N_15194,N_14818,N_14854);
xnor U15195 (N_15195,N_14625,N_14876);
and U15196 (N_15196,N_14775,N_14871);
nor U15197 (N_15197,N_14527,N_14766);
nor U15198 (N_15198,N_14619,N_14518);
and U15199 (N_15199,N_14425,N_14404);
or U15200 (N_15200,N_14857,N_14400);
nand U15201 (N_15201,N_14745,N_14441);
xor U15202 (N_15202,N_14846,N_14630);
nor U15203 (N_15203,N_14787,N_14612);
nor U15204 (N_15204,N_14896,N_14959);
nand U15205 (N_15205,N_14671,N_14822);
xnor U15206 (N_15206,N_14870,N_14776);
or U15207 (N_15207,N_14918,N_14512);
or U15208 (N_15208,N_14693,N_14761);
and U15209 (N_15209,N_14804,N_14573);
nand U15210 (N_15210,N_14839,N_14411);
or U15211 (N_15211,N_14575,N_14808);
and U15212 (N_15212,N_14410,N_14748);
nand U15213 (N_15213,N_14865,N_14907);
and U15214 (N_15214,N_14835,N_14802);
nor U15215 (N_15215,N_14817,N_14973);
nand U15216 (N_15216,N_14450,N_14613);
and U15217 (N_15217,N_14686,N_14998);
and U15218 (N_15218,N_14909,N_14461);
or U15219 (N_15219,N_14783,N_14682);
nand U15220 (N_15220,N_14946,N_14840);
nor U15221 (N_15221,N_14826,N_14723);
xor U15222 (N_15222,N_14798,N_14859);
nor U15223 (N_15223,N_14697,N_14815);
or U15224 (N_15224,N_14665,N_14419);
or U15225 (N_15225,N_14491,N_14657);
nand U15226 (N_15226,N_14742,N_14543);
and U15227 (N_15227,N_14661,N_14488);
or U15228 (N_15228,N_14472,N_14809);
xor U15229 (N_15229,N_14587,N_14694);
or U15230 (N_15230,N_14806,N_14947);
xor U15231 (N_15231,N_14734,N_14677);
and U15232 (N_15232,N_14864,N_14688);
nor U15233 (N_15233,N_14708,N_14948);
or U15234 (N_15234,N_14529,N_14850);
nor U15235 (N_15235,N_14666,N_14541);
nand U15236 (N_15236,N_14969,N_14983);
nor U15237 (N_15237,N_14637,N_14402);
nor U15238 (N_15238,N_14605,N_14751);
or U15239 (N_15239,N_14836,N_14475);
nand U15240 (N_15240,N_14856,N_14444);
and U15241 (N_15241,N_14474,N_14565);
xor U15242 (N_15242,N_14602,N_14604);
nand U15243 (N_15243,N_14713,N_14520);
and U15244 (N_15244,N_14953,N_14417);
xor U15245 (N_15245,N_14834,N_14895);
nand U15246 (N_15246,N_14552,N_14528);
xor U15247 (N_15247,N_14540,N_14501);
xnor U15248 (N_15248,N_14403,N_14687);
and U15249 (N_15249,N_14966,N_14814);
xor U15250 (N_15250,N_14771,N_14571);
and U15251 (N_15251,N_14433,N_14828);
and U15252 (N_15252,N_14477,N_14997);
and U15253 (N_15253,N_14726,N_14794);
or U15254 (N_15254,N_14600,N_14899);
or U15255 (N_15255,N_14796,N_14647);
nor U15256 (N_15256,N_14820,N_14676);
or U15257 (N_15257,N_14741,N_14588);
xor U15258 (N_15258,N_14513,N_14731);
xnor U15259 (N_15259,N_14623,N_14922);
and U15260 (N_15260,N_14547,N_14827);
and U15261 (N_15261,N_14727,N_14502);
xor U15262 (N_15262,N_14902,N_14690);
nor U15263 (N_15263,N_14633,N_14406);
and U15264 (N_15264,N_14418,N_14762);
nand U15265 (N_15265,N_14466,N_14407);
nor U15266 (N_15266,N_14638,N_14935);
nand U15267 (N_15267,N_14559,N_14667);
and U15268 (N_15268,N_14554,N_14877);
nand U15269 (N_15269,N_14680,N_14542);
nand U15270 (N_15270,N_14974,N_14564);
nand U15271 (N_15271,N_14844,N_14484);
xnor U15272 (N_15272,N_14662,N_14445);
and U15273 (N_15273,N_14570,N_14615);
nor U15274 (N_15274,N_14480,N_14645);
xor U15275 (N_15275,N_14599,N_14830);
nor U15276 (N_15276,N_14702,N_14811);
xor U15277 (N_15277,N_14972,N_14684);
or U15278 (N_15278,N_14800,N_14853);
xnor U15279 (N_15279,N_14950,N_14970);
or U15280 (N_15280,N_14583,N_14568);
nand U15281 (N_15281,N_14890,N_14779);
nor U15282 (N_15282,N_14888,N_14772);
xnor U15283 (N_15283,N_14718,N_14634);
nand U15284 (N_15284,N_14635,N_14943);
and U15285 (N_15285,N_14923,N_14431);
nor U15286 (N_15286,N_14819,N_14670);
and U15287 (N_15287,N_14965,N_14862);
xnor U15288 (N_15288,N_14538,N_14716);
or U15289 (N_15289,N_14616,N_14506);
nand U15290 (N_15290,N_14449,N_14914);
nor U15291 (N_15291,N_14963,N_14790);
nor U15292 (N_15292,N_14553,N_14995);
and U15293 (N_15293,N_14975,N_14978);
or U15294 (N_15294,N_14558,N_14622);
or U15295 (N_15295,N_14415,N_14908);
nor U15296 (N_15296,N_14886,N_14654);
nor U15297 (N_15297,N_14855,N_14462);
nor U15298 (N_15298,N_14481,N_14733);
nand U15299 (N_15299,N_14537,N_14810);
or U15300 (N_15300,N_14599,N_14851);
xor U15301 (N_15301,N_14569,N_14517);
nor U15302 (N_15302,N_14536,N_14633);
nand U15303 (N_15303,N_14462,N_14851);
or U15304 (N_15304,N_14981,N_14661);
or U15305 (N_15305,N_14916,N_14742);
and U15306 (N_15306,N_14515,N_14818);
nand U15307 (N_15307,N_14974,N_14478);
nand U15308 (N_15308,N_14704,N_14864);
nor U15309 (N_15309,N_14412,N_14474);
or U15310 (N_15310,N_14764,N_14794);
nand U15311 (N_15311,N_14743,N_14874);
nand U15312 (N_15312,N_14695,N_14451);
or U15313 (N_15313,N_14431,N_14670);
nand U15314 (N_15314,N_14681,N_14526);
or U15315 (N_15315,N_14977,N_14416);
nand U15316 (N_15316,N_14931,N_14447);
or U15317 (N_15317,N_14860,N_14885);
nor U15318 (N_15318,N_14860,N_14723);
nor U15319 (N_15319,N_14994,N_14855);
or U15320 (N_15320,N_14867,N_14623);
and U15321 (N_15321,N_14813,N_14764);
and U15322 (N_15322,N_14951,N_14440);
xor U15323 (N_15323,N_14894,N_14626);
nor U15324 (N_15324,N_14612,N_14674);
xor U15325 (N_15325,N_14937,N_14799);
and U15326 (N_15326,N_14458,N_14909);
nor U15327 (N_15327,N_14723,N_14837);
or U15328 (N_15328,N_14760,N_14635);
and U15329 (N_15329,N_14451,N_14935);
xnor U15330 (N_15330,N_14899,N_14421);
xor U15331 (N_15331,N_14641,N_14634);
and U15332 (N_15332,N_14790,N_14822);
nor U15333 (N_15333,N_14677,N_14909);
xor U15334 (N_15334,N_14469,N_14592);
nor U15335 (N_15335,N_14696,N_14839);
and U15336 (N_15336,N_14864,N_14752);
nor U15337 (N_15337,N_14641,N_14597);
xnor U15338 (N_15338,N_14471,N_14785);
nor U15339 (N_15339,N_14474,N_14797);
and U15340 (N_15340,N_14413,N_14558);
nor U15341 (N_15341,N_14979,N_14577);
or U15342 (N_15342,N_14582,N_14947);
or U15343 (N_15343,N_14634,N_14706);
nor U15344 (N_15344,N_14853,N_14857);
nor U15345 (N_15345,N_14949,N_14885);
or U15346 (N_15346,N_14768,N_14805);
xor U15347 (N_15347,N_14941,N_14605);
or U15348 (N_15348,N_14593,N_14420);
or U15349 (N_15349,N_14884,N_14755);
nand U15350 (N_15350,N_14807,N_14795);
nor U15351 (N_15351,N_14961,N_14755);
nor U15352 (N_15352,N_14718,N_14933);
or U15353 (N_15353,N_14454,N_14667);
nor U15354 (N_15354,N_14977,N_14964);
nor U15355 (N_15355,N_14818,N_14715);
nand U15356 (N_15356,N_14993,N_14727);
xnor U15357 (N_15357,N_14438,N_14952);
xnor U15358 (N_15358,N_14869,N_14945);
nand U15359 (N_15359,N_14428,N_14449);
and U15360 (N_15360,N_14946,N_14430);
or U15361 (N_15361,N_14654,N_14483);
or U15362 (N_15362,N_14775,N_14850);
nand U15363 (N_15363,N_14500,N_14878);
nand U15364 (N_15364,N_14528,N_14789);
or U15365 (N_15365,N_14957,N_14578);
xnor U15366 (N_15366,N_14532,N_14767);
xor U15367 (N_15367,N_14909,N_14518);
xnor U15368 (N_15368,N_14711,N_14660);
or U15369 (N_15369,N_14981,N_14745);
nor U15370 (N_15370,N_14406,N_14828);
nand U15371 (N_15371,N_14485,N_14616);
nand U15372 (N_15372,N_14422,N_14814);
and U15373 (N_15373,N_14840,N_14592);
or U15374 (N_15374,N_14649,N_14420);
and U15375 (N_15375,N_14470,N_14922);
xnor U15376 (N_15376,N_14466,N_14903);
nor U15377 (N_15377,N_14615,N_14847);
or U15378 (N_15378,N_14422,N_14568);
nor U15379 (N_15379,N_14579,N_14734);
nor U15380 (N_15380,N_14630,N_14863);
and U15381 (N_15381,N_14741,N_14827);
or U15382 (N_15382,N_14411,N_14825);
and U15383 (N_15383,N_14945,N_14421);
xnor U15384 (N_15384,N_14760,N_14411);
or U15385 (N_15385,N_14668,N_14654);
and U15386 (N_15386,N_14937,N_14793);
or U15387 (N_15387,N_14400,N_14716);
nand U15388 (N_15388,N_14617,N_14677);
nand U15389 (N_15389,N_14889,N_14809);
nor U15390 (N_15390,N_14417,N_14551);
or U15391 (N_15391,N_14540,N_14879);
nand U15392 (N_15392,N_14998,N_14487);
or U15393 (N_15393,N_14762,N_14401);
xnor U15394 (N_15394,N_14641,N_14620);
xor U15395 (N_15395,N_14415,N_14802);
nand U15396 (N_15396,N_14525,N_14496);
nor U15397 (N_15397,N_14924,N_14585);
nor U15398 (N_15398,N_14635,N_14764);
nor U15399 (N_15399,N_14522,N_14936);
and U15400 (N_15400,N_14941,N_14595);
nand U15401 (N_15401,N_14455,N_14932);
nand U15402 (N_15402,N_14406,N_14760);
nor U15403 (N_15403,N_14478,N_14986);
and U15404 (N_15404,N_14995,N_14434);
nand U15405 (N_15405,N_14828,N_14727);
or U15406 (N_15406,N_14938,N_14605);
nor U15407 (N_15407,N_14717,N_14401);
or U15408 (N_15408,N_14551,N_14984);
or U15409 (N_15409,N_14702,N_14916);
and U15410 (N_15410,N_14839,N_14420);
nand U15411 (N_15411,N_14586,N_14801);
or U15412 (N_15412,N_14627,N_14439);
and U15413 (N_15413,N_14743,N_14541);
or U15414 (N_15414,N_14530,N_14410);
xnor U15415 (N_15415,N_14401,N_14945);
xor U15416 (N_15416,N_14433,N_14941);
and U15417 (N_15417,N_14544,N_14814);
or U15418 (N_15418,N_14930,N_14875);
and U15419 (N_15419,N_14626,N_14451);
and U15420 (N_15420,N_14730,N_14936);
nand U15421 (N_15421,N_14411,N_14671);
and U15422 (N_15422,N_14487,N_14416);
nand U15423 (N_15423,N_14676,N_14906);
xor U15424 (N_15424,N_14816,N_14931);
xnor U15425 (N_15425,N_14776,N_14862);
nor U15426 (N_15426,N_14479,N_14931);
nand U15427 (N_15427,N_14495,N_14971);
nand U15428 (N_15428,N_14596,N_14498);
nand U15429 (N_15429,N_14423,N_14903);
or U15430 (N_15430,N_14434,N_14767);
nand U15431 (N_15431,N_14517,N_14771);
nand U15432 (N_15432,N_14905,N_14928);
xor U15433 (N_15433,N_14804,N_14794);
nor U15434 (N_15434,N_14460,N_14910);
and U15435 (N_15435,N_14990,N_14992);
nor U15436 (N_15436,N_14536,N_14719);
nand U15437 (N_15437,N_14664,N_14449);
nand U15438 (N_15438,N_14987,N_14558);
nand U15439 (N_15439,N_14437,N_14587);
xnor U15440 (N_15440,N_14575,N_14473);
nand U15441 (N_15441,N_14785,N_14934);
and U15442 (N_15442,N_14723,N_14531);
nor U15443 (N_15443,N_14469,N_14826);
and U15444 (N_15444,N_14435,N_14488);
nand U15445 (N_15445,N_14462,N_14459);
nand U15446 (N_15446,N_14614,N_14859);
or U15447 (N_15447,N_14855,N_14687);
nor U15448 (N_15448,N_14733,N_14441);
xor U15449 (N_15449,N_14760,N_14403);
or U15450 (N_15450,N_14834,N_14414);
nor U15451 (N_15451,N_14632,N_14888);
nor U15452 (N_15452,N_14480,N_14983);
nand U15453 (N_15453,N_14711,N_14811);
and U15454 (N_15454,N_14407,N_14950);
nor U15455 (N_15455,N_14609,N_14543);
nand U15456 (N_15456,N_14868,N_14594);
xnor U15457 (N_15457,N_14961,N_14582);
or U15458 (N_15458,N_14494,N_14492);
nor U15459 (N_15459,N_14704,N_14541);
or U15460 (N_15460,N_14541,N_14521);
xor U15461 (N_15461,N_14646,N_14723);
or U15462 (N_15462,N_14402,N_14534);
nand U15463 (N_15463,N_14451,N_14558);
or U15464 (N_15464,N_14751,N_14465);
or U15465 (N_15465,N_14965,N_14734);
or U15466 (N_15466,N_14419,N_14672);
nor U15467 (N_15467,N_14984,N_14783);
and U15468 (N_15468,N_14645,N_14774);
nor U15469 (N_15469,N_14766,N_14600);
or U15470 (N_15470,N_14464,N_14788);
or U15471 (N_15471,N_14994,N_14747);
xor U15472 (N_15472,N_14943,N_14920);
and U15473 (N_15473,N_14750,N_14747);
and U15474 (N_15474,N_14740,N_14599);
or U15475 (N_15475,N_14515,N_14744);
or U15476 (N_15476,N_14623,N_14755);
xnor U15477 (N_15477,N_14826,N_14562);
nand U15478 (N_15478,N_14862,N_14807);
and U15479 (N_15479,N_14800,N_14791);
and U15480 (N_15480,N_14806,N_14460);
or U15481 (N_15481,N_14484,N_14472);
and U15482 (N_15482,N_14699,N_14982);
and U15483 (N_15483,N_14570,N_14924);
and U15484 (N_15484,N_14978,N_14533);
nor U15485 (N_15485,N_14778,N_14734);
or U15486 (N_15486,N_14918,N_14464);
nand U15487 (N_15487,N_14608,N_14681);
xnor U15488 (N_15488,N_14513,N_14867);
nand U15489 (N_15489,N_14654,N_14960);
nor U15490 (N_15490,N_14726,N_14430);
nor U15491 (N_15491,N_14472,N_14945);
and U15492 (N_15492,N_14805,N_14728);
and U15493 (N_15493,N_14710,N_14690);
nand U15494 (N_15494,N_14758,N_14664);
and U15495 (N_15495,N_14875,N_14609);
and U15496 (N_15496,N_14942,N_14909);
and U15497 (N_15497,N_14954,N_14813);
nor U15498 (N_15498,N_14401,N_14731);
nand U15499 (N_15499,N_14940,N_14941);
or U15500 (N_15500,N_14481,N_14469);
nand U15501 (N_15501,N_14495,N_14612);
or U15502 (N_15502,N_14957,N_14739);
xnor U15503 (N_15503,N_14979,N_14827);
or U15504 (N_15504,N_14509,N_14493);
nor U15505 (N_15505,N_14763,N_14691);
xor U15506 (N_15506,N_14798,N_14432);
nor U15507 (N_15507,N_14566,N_14700);
nand U15508 (N_15508,N_14535,N_14653);
nor U15509 (N_15509,N_14725,N_14475);
nor U15510 (N_15510,N_14643,N_14880);
nor U15511 (N_15511,N_14831,N_14979);
and U15512 (N_15512,N_14441,N_14477);
or U15513 (N_15513,N_14893,N_14957);
xor U15514 (N_15514,N_14846,N_14446);
or U15515 (N_15515,N_14976,N_14938);
xnor U15516 (N_15516,N_14740,N_14834);
and U15517 (N_15517,N_14709,N_14527);
or U15518 (N_15518,N_14968,N_14787);
and U15519 (N_15519,N_14424,N_14812);
or U15520 (N_15520,N_14401,N_14585);
or U15521 (N_15521,N_14936,N_14894);
and U15522 (N_15522,N_14733,N_14783);
nor U15523 (N_15523,N_14565,N_14479);
nand U15524 (N_15524,N_14859,N_14664);
or U15525 (N_15525,N_14809,N_14825);
and U15526 (N_15526,N_14428,N_14916);
or U15527 (N_15527,N_14613,N_14769);
nand U15528 (N_15528,N_14515,N_14462);
nor U15529 (N_15529,N_14949,N_14543);
or U15530 (N_15530,N_14516,N_14957);
xor U15531 (N_15531,N_14454,N_14839);
or U15532 (N_15532,N_14627,N_14703);
or U15533 (N_15533,N_14631,N_14442);
nor U15534 (N_15534,N_14911,N_14512);
xnor U15535 (N_15535,N_14892,N_14459);
or U15536 (N_15536,N_14784,N_14722);
or U15537 (N_15537,N_14933,N_14954);
nand U15538 (N_15538,N_14497,N_14458);
nand U15539 (N_15539,N_14832,N_14512);
nand U15540 (N_15540,N_14949,N_14806);
and U15541 (N_15541,N_14847,N_14665);
or U15542 (N_15542,N_14722,N_14473);
xnor U15543 (N_15543,N_14479,N_14532);
and U15544 (N_15544,N_14691,N_14622);
nor U15545 (N_15545,N_14913,N_14582);
and U15546 (N_15546,N_14613,N_14993);
or U15547 (N_15547,N_14991,N_14727);
xor U15548 (N_15548,N_14731,N_14427);
nor U15549 (N_15549,N_14805,N_14523);
nor U15550 (N_15550,N_14613,N_14740);
nor U15551 (N_15551,N_14459,N_14440);
nor U15552 (N_15552,N_14415,N_14897);
or U15553 (N_15553,N_14834,N_14623);
or U15554 (N_15554,N_14701,N_14732);
or U15555 (N_15555,N_14958,N_14429);
and U15556 (N_15556,N_14942,N_14686);
xnor U15557 (N_15557,N_14591,N_14927);
or U15558 (N_15558,N_14690,N_14737);
and U15559 (N_15559,N_14857,N_14436);
nand U15560 (N_15560,N_14502,N_14736);
or U15561 (N_15561,N_14600,N_14865);
or U15562 (N_15562,N_14956,N_14860);
and U15563 (N_15563,N_14703,N_14700);
nor U15564 (N_15564,N_14447,N_14442);
and U15565 (N_15565,N_14758,N_14581);
nor U15566 (N_15566,N_14566,N_14477);
or U15567 (N_15567,N_14909,N_14434);
and U15568 (N_15568,N_14557,N_14429);
nand U15569 (N_15569,N_14486,N_14829);
and U15570 (N_15570,N_14790,N_14614);
or U15571 (N_15571,N_14780,N_14522);
xor U15572 (N_15572,N_14512,N_14438);
xor U15573 (N_15573,N_14750,N_14422);
nand U15574 (N_15574,N_14972,N_14749);
nor U15575 (N_15575,N_14724,N_14598);
nor U15576 (N_15576,N_14681,N_14528);
or U15577 (N_15577,N_14654,N_14721);
or U15578 (N_15578,N_14911,N_14858);
or U15579 (N_15579,N_14428,N_14464);
nand U15580 (N_15580,N_14870,N_14911);
nor U15581 (N_15581,N_14968,N_14941);
nor U15582 (N_15582,N_14501,N_14783);
and U15583 (N_15583,N_14410,N_14895);
xor U15584 (N_15584,N_14624,N_14499);
xnor U15585 (N_15585,N_14408,N_14404);
nor U15586 (N_15586,N_14496,N_14549);
or U15587 (N_15587,N_14516,N_14878);
nor U15588 (N_15588,N_14674,N_14464);
nor U15589 (N_15589,N_14700,N_14643);
or U15590 (N_15590,N_14904,N_14653);
xnor U15591 (N_15591,N_14485,N_14649);
nor U15592 (N_15592,N_14930,N_14653);
and U15593 (N_15593,N_14513,N_14418);
xnor U15594 (N_15594,N_14712,N_14817);
nor U15595 (N_15595,N_14668,N_14754);
or U15596 (N_15596,N_14976,N_14651);
nor U15597 (N_15597,N_14435,N_14482);
or U15598 (N_15598,N_14521,N_14910);
and U15599 (N_15599,N_14403,N_14692);
or U15600 (N_15600,N_15317,N_15392);
and U15601 (N_15601,N_15546,N_15112);
or U15602 (N_15602,N_15246,N_15327);
and U15603 (N_15603,N_15293,N_15589);
xor U15604 (N_15604,N_15396,N_15268);
or U15605 (N_15605,N_15563,N_15080);
xnor U15606 (N_15606,N_15348,N_15463);
or U15607 (N_15607,N_15130,N_15049);
xnor U15608 (N_15608,N_15524,N_15505);
and U15609 (N_15609,N_15264,N_15586);
and U15610 (N_15610,N_15275,N_15515);
and U15611 (N_15611,N_15141,N_15026);
xor U15612 (N_15612,N_15542,N_15371);
nor U15613 (N_15613,N_15552,N_15596);
and U15614 (N_15614,N_15222,N_15210);
or U15615 (N_15615,N_15322,N_15184);
or U15616 (N_15616,N_15598,N_15018);
or U15617 (N_15617,N_15226,N_15368);
nand U15618 (N_15618,N_15370,N_15543);
nand U15619 (N_15619,N_15223,N_15186);
nor U15620 (N_15620,N_15061,N_15167);
nand U15621 (N_15621,N_15104,N_15538);
nand U15622 (N_15622,N_15136,N_15235);
xor U15623 (N_15623,N_15206,N_15233);
or U15624 (N_15624,N_15056,N_15219);
and U15625 (N_15625,N_15457,N_15177);
or U15626 (N_15626,N_15060,N_15193);
and U15627 (N_15627,N_15415,N_15394);
or U15628 (N_15628,N_15431,N_15168);
nor U15629 (N_15629,N_15380,N_15227);
nor U15630 (N_15630,N_15428,N_15034);
nor U15631 (N_15631,N_15559,N_15137);
xor U15632 (N_15632,N_15000,N_15045);
and U15633 (N_15633,N_15169,N_15074);
and U15634 (N_15634,N_15465,N_15307);
and U15635 (N_15635,N_15148,N_15304);
and U15636 (N_15636,N_15551,N_15076);
or U15637 (N_15637,N_15084,N_15208);
nand U15638 (N_15638,N_15255,N_15331);
nor U15639 (N_15639,N_15520,N_15145);
or U15640 (N_15640,N_15570,N_15236);
or U15641 (N_15641,N_15260,N_15590);
or U15642 (N_15642,N_15452,N_15333);
xnor U15643 (N_15643,N_15135,N_15350);
xnor U15644 (N_15644,N_15161,N_15514);
xnor U15645 (N_15645,N_15464,N_15432);
nand U15646 (N_15646,N_15471,N_15288);
nand U15647 (N_15647,N_15292,N_15129);
nor U15648 (N_15648,N_15225,N_15162);
nand U15649 (N_15649,N_15351,N_15152);
or U15650 (N_15650,N_15593,N_15484);
or U15651 (N_15651,N_15578,N_15532);
nor U15652 (N_15652,N_15088,N_15439);
and U15653 (N_15653,N_15182,N_15065);
nor U15654 (N_15654,N_15154,N_15143);
nor U15655 (N_15655,N_15361,N_15277);
and U15656 (N_15656,N_15441,N_15442);
nand U15657 (N_15657,N_15533,N_15519);
xnor U15658 (N_15658,N_15384,N_15427);
xor U15659 (N_15659,N_15200,N_15339);
or U15660 (N_15660,N_15199,N_15165);
or U15661 (N_15661,N_15594,N_15021);
and U15662 (N_15662,N_15204,N_15248);
xor U15663 (N_15663,N_15382,N_15405);
xor U15664 (N_15664,N_15547,N_15330);
and U15665 (N_15665,N_15115,N_15599);
xnor U15666 (N_15666,N_15069,N_15151);
and U15667 (N_15667,N_15028,N_15466);
xor U15668 (N_15668,N_15114,N_15501);
or U15669 (N_15669,N_15353,N_15029);
or U15670 (N_15670,N_15269,N_15447);
and U15671 (N_15671,N_15566,N_15573);
or U15672 (N_15672,N_15079,N_15407);
nor U15673 (N_15673,N_15527,N_15530);
nor U15674 (N_15674,N_15244,N_15051);
nand U15675 (N_15675,N_15118,N_15521);
xor U15676 (N_15676,N_15138,N_15400);
nand U15677 (N_15677,N_15127,N_15075);
or U15678 (N_15678,N_15133,N_15095);
xnor U15679 (N_15679,N_15173,N_15580);
xnor U15680 (N_15680,N_15174,N_15240);
nor U15681 (N_15681,N_15592,N_15271);
nand U15682 (N_15682,N_15399,N_15078);
xor U15683 (N_15683,N_15425,N_15469);
or U15684 (N_15684,N_15356,N_15150);
nor U15685 (N_15685,N_15090,N_15013);
nand U15686 (N_15686,N_15247,N_15087);
xnor U15687 (N_15687,N_15446,N_15451);
or U15688 (N_15688,N_15047,N_15362);
and U15689 (N_15689,N_15040,N_15408);
nor U15690 (N_15690,N_15242,N_15057);
nor U15691 (N_15691,N_15276,N_15003);
and U15692 (N_15692,N_15209,N_15364);
xnor U15693 (N_15693,N_15387,N_15146);
xor U15694 (N_15694,N_15207,N_15403);
xor U15695 (N_15695,N_15468,N_15556);
nor U15696 (N_15696,N_15373,N_15241);
and U15697 (N_15697,N_15582,N_15218);
nand U15698 (N_15698,N_15153,N_15109);
and U15699 (N_15699,N_15259,N_15587);
nand U15700 (N_15700,N_15377,N_15429);
nand U15701 (N_15701,N_15190,N_15500);
or U15702 (N_15702,N_15094,N_15009);
nand U15703 (N_15703,N_15561,N_15478);
or U15704 (N_15704,N_15390,N_15585);
nor U15705 (N_15705,N_15054,N_15503);
or U15706 (N_15706,N_15103,N_15295);
and U15707 (N_15707,N_15323,N_15383);
nor U15708 (N_15708,N_15274,N_15316);
xnor U15709 (N_15709,N_15092,N_15335);
or U15710 (N_15710,N_15419,N_15261);
or U15711 (N_15711,N_15203,N_15495);
nand U15712 (N_15712,N_15488,N_15280);
nor U15713 (N_15713,N_15379,N_15041);
xor U15714 (N_15714,N_15300,N_15564);
nor U15715 (N_15715,N_15489,N_15569);
xor U15716 (N_15716,N_15588,N_15262);
or U15717 (N_15717,N_15024,N_15393);
xnor U15718 (N_15718,N_15416,N_15391);
or U15719 (N_15719,N_15343,N_15224);
nand U15720 (N_15720,N_15281,N_15250);
nor U15721 (N_15721,N_15212,N_15597);
nor U15722 (N_15722,N_15297,N_15097);
nor U15723 (N_15723,N_15196,N_15494);
or U15724 (N_15724,N_15073,N_15375);
nand U15725 (N_15725,N_15105,N_15461);
or U15726 (N_15726,N_15251,N_15321);
xor U15727 (N_15727,N_15517,N_15132);
nor U15728 (N_15728,N_15577,N_15395);
nand U15729 (N_15729,N_15315,N_15144);
and U15730 (N_15730,N_15002,N_15249);
nand U15731 (N_15731,N_15422,N_15512);
and U15732 (N_15732,N_15102,N_15411);
nor U15733 (N_15733,N_15459,N_15194);
and U15734 (N_15734,N_15077,N_15319);
nor U15735 (N_15735,N_15159,N_15306);
xor U15736 (N_15736,N_15336,N_15410);
or U15737 (N_15737,N_15285,N_15044);
and U15738 (N_15738,N_15091,N_15360);
nor U15739 (N_15739,N_15473,N_15560);
and U15740 (N_15740,N_15492,N_15272);
xnor U15741 (N_15741,N_15312,N_15001);
nor U15742 (N_15742,N_15301,N_15004);
and U15743 (N_15743,N_15243,N_15485);
xnor U15744 (N_15744,N_15365,N_15172);
xor U15745 (N_15745,N_15116,N_15499);
nand U15746 (N_15746,N_15456,N_15140);
nor U15747 (N_15747,N_15481,N_15011);
xnor U15748 (N_15748,N_15106,N_15359);
xnor U15749 (N_15749,N_15017,N_15420);
xor U15750 (N_15750,N_15309,N_15037);
and U15751 (N_15751,N_15205,N_15283);
nand U15752 (N_15752,N_15035,N_15438);
nand U15753 (N_15753,N_15433,N_15066);
and U15754 (N_15754,N_15064,N_15491);
xor U15755 (N_15755,N_15329,N_15014);
and U15756 (N_15756,N_15282,N_15213);
nor U15757 (N_15757,N_15413,N_15482);
and U15758 (N_15758,N_15089,N_15126);
xnor U15759 (N_15759,N_15231,N_15342);
and U15760 (N_15760,N_15591,N_15513);
xnor U15761 (N_15761,N_15526,N_15296);
or U15762 (N_15762,N_15449,N_15234);
nor U15763 (N_15763,N_15548,N_15358);
and U15764 (N_15764,N_15033,N_15349);
nand U15765 (N_15765,N_15541,N_15082);
or U15766 (N_15766,N_15254,N_15498);
or U15767 (N_15767,N_15458,N_15470);
nand U15768 (N_15768,N_15314,N_15022);
or U15769 (N_15769,N_15553,N_15313);
nand U15770 (N_15770,N_15445,N_15142);
nor U15771 (N_15771,N_15211,N_15099);
and U15772 (N_15772,N_15595,N_15052);
nor U15773 (N_15773,N_15038,N_15217);
nand U15774 (N_15774,N_15575,N_15120);
or U15775 (N_15775,N_15279,N_15472);
nor U15776 (N_15776,N_15302,N_15555);
nand U15777 (N_15777,N_15545,N_15020);
xor U15778 (N_15778,N_15518,N_15121);
xnor U15779 (N_15779,N_15531,N_15414);
xor U15780 (N_15780,N_15270,N_15324);
or U15781 (N_15781,N_15298,N_15549);
nor U15782 (N_15782,N_15171,N_15558);
or U15783 (N_15783,N_15523,N_15178);
xnor U15784 (N_15784,N_15156,N_15070);
or U15785 (N_15785,N_15253,N_15572);
nand U15786 (N_15786,N_15055,N_15185);
and U15787 (N_15787,N_15397,N_15273);
and U15788 (N_15788,N_15023,N_15557);
and U15789 (N_15789,N_15030,N_15032);
nor U15790 (N_15790,N_15238,N_15216);
and U15791 (N_15791,N_15048,N_15170);
nand U15792 (N_15792,N_15430,N_15110);
or U15793 (N_15793,N_15096,N_15423);
xor U15794 (N_15794,N_15344,N_15486);
nor U15795 (N_15795,N_15256,N_15477);
nand U15796 (N_15796,N_15181,N_15019);
nand U15797 (N_15797,N_15509,N_15529);
xnor U15798 (N_15798,N_15085,N_15012);
and U15799 (N_15799,N_15155,N_15550);
nor U15800 (N_15800,N_15506,N_15291);
xor U15801 (N_15801,N_15083,N_15567);
or U15802 (N_15802,N_15455,N_15487);
or U15803 (N_15803,N_15337,N_15122);
xnor U15804 (N_15804,N_15479,N_15474);
or U15805 (N_15805,N_15286,N_15576);
or U15806 (N_15806,N_15502,N_15025);
or U15807 (N_15807,N_15389,N_15149);
nand U15808 (N_15808,N_15245,N_15005);
and U15809 (N_15809,N_15139,N_15284);
nand U15810 (N_15810,N_15183,N_15202);
and U15811 (N_15811,N_15128,N_15436);
xor U15812 (N_15812,N_15239,N_15426);
xor U15813 (N_15813,N_15039,N_15453);
and U15814 (N_15814,N_15062,N_15230);
and U15815 (N_15815,N_15444,N_15435);
nor U15816 (N_15816,N_15418,N_15562);
or U15817 (N_15817,N_15326,N_15510);
and U15818 (N_15818,N_15355,N_15565);
nor U15819 (N_15819,N_15197,N_15374);
nand U15820 (N_15820,N_15320,N_15369);
xnor U15821 (N_15821,N_15376,N_15071);
nand U15822 (N_15822,N_15311,N_15113);
and U15823 (N_15823,N_15179,N_15310);
nor U15824 (N_15824,N_15583,N_15305);
and U15825 (N_15825,N_15581,N_15043);
xnor U15826 (N_15826,N_15584,N_15544);
nand U15827 (N_15827,N_15124,N_15493);
nor U15828 (N_15828,N_15540,N_15554);
nor U15829 (N_15829,N_15237,N_15053);
nor U15830 (N_15830,N_15328,N_15215);
nor U15831 (N_15831,N_15265,N_15462);
nand U15832 (N_15832,N_15163,N_15189);
or U15833 (N_15833,N_15042,N_15166);
nor U15834 (N_15834,N_15325,N_15192);
and U15835 (N_15835,N_15507,N_15160);
nand U15836 (N_15836,N_15525,N_15450);
xnor U15837 (N_15837,N_15434,N_15340);
nor U15838 (N_15838,N_15016,N_15357);
and U15839 (N_15839,N_15341,N_15508);
nor U15840 (N_15840,N_15406,N_15067);
or U15841 (N_15841,N_15006,N_15528);
and U15842 (N_15842,N_15579,N_15386);
nand U15843 (N_15843,N_15354,N_15497);
or U15844 (N_15844,N_15467,N_15409);
and U15845 (N_15845,N_15015,N_15220);
nor U15846 (N_15846,N_15367,N_15332);
nand U15847 (N_15847,N_15027,N_15345);
nor U15848 (N_15848,N_15201,N_15421);
xor U15849 (N_15849,N_15007,N_15093);
nor U15850 (N_15850,N_15278,N_15101);
nor U15851 (N_15851,N_15257,N_15537);
nor U15852 (N_15852,N_15440,N_15287);
xnor U15853 (N_15853,N_15195,N_15483);
and U15854 (N_15854,N_15125,N_15516);
nor U15855 (N_15855,N_15046,N_15347);
or U15856 (N_15856,N_15448,N_15263);
or U15857 (N_15857,N_15108,N_15378);
nor U15858 (N_15858,N_15198,N_15008);
nand U15859 (N_15859,N_15443,N_15031);
nor U15860 (N_15860,N_15058,N_15187);
xor U15861 (N_15861,N_15229,N_15147);
or U15862 (N_15862,N_15574,N_15111);
xnor U15863 (N_15863,N_15401,N_15119);
or U15864 (N_15864,N_15385,N_15098);
nor U15865 (N_15865,N_15496,N_15107);
xnor U15866 (N_15866,N_15571,N_15131);
or U15867 (N_15867,N_15402,N_15117);
or U15868 (N_15868,N_15050,N_15346);
nand U15869 (N_15869,N_15123,N_15476);
xnor U15870 (N_15870,N_15334,N_15511);
nand U15871 (N_15871,N_15010,N_15068);
nand U15872 (N_15872,N_15417,N_15258);
or U15873 (N_15873,N_15460,N_15164);
and U15874 (N_15874,N_15188,N_15475);
xor U15875 (N_15875,N_15252,N_15504);
or U15876 (N_15876,N_15299,N_15522);
xor U15877 (N_15877,N_15352,N_15176);
xor U15878 (N_15878,N_15388,N_15175);
or U15879 (N_15879,N_15191,N_15294);
nor U15880 (N_15880,N_15318,N_15536);
xnor U15881 (N_15881,N_15372,N_15158);
nor U15882 (N_15882,N_15100,N_15228);
xor U15883 (N_15883,N_15303,N_15308);
nand U15884 (N_15884,N_15063,N_15221);
and U15885 (N_15885,N_15134,N_15338);
nor U15886 (N_15886,N_15437,N_15454);
and U15887 (N_15887,N_15157,N_15412);
and U15888 (N_15888,N_15381,N_15036);
nand U15889 (N_15889,N_15363,N_15086);
nand U15890 (N_15890,N_15568,N_15404);
nand U15891 (N_15891,N_15180,N_15290);
nor U15892 (N_15892,N_15266,N_15424);
nand U15893 (N_15893,N_15398,N_15072);
xnor U15894 (N_15894,N_15535,N_15490);
nor U15895 (N_15895,N_15081,N_15366);
xor U15896 (N_15896,N_15539,N_15289);
or U15897 (N_15897,N_15232,N_15214);
and U15898 (N_15898,N_15059,N_15534);
and U15899 (N_15899,N_15267,N_15480);
nor U15900 (N_15900,N_15101,N_15221);
or U15901 (N_15901,N_15104,N_15227);
nand U15902 (N_15902,N_15437,N_15332);
xnor U15903 (N_15903,N_15076,N_15163);
or U15904 (N_15904,N_15314,N_15160);
nor U15905 (N_15905,N_15378,N_15489);
nor U15906 (N_15906,N_15213,N_15437);
nand U15907 (N_15907,N_15269,N_15337);
nor U15908 (N_15908,N_15005,N_15433);
nor U15909 (N_15909,N_15442,N_15289);
nand U15910 (N_15910,N_15412,N_15099);
nand U15911 (N_15911,N_15555,N_15485);
nand U15912 (N_15912,N_15155,N_15294);
or U15913 (N_15913,N_15288,N_15312);
or U15914 (N_15914,N_15179,N_15196);
nor U15915 (N_15915,N_15260,N_15099);
nor U15916 (N_15916,N_15081,N_15084);
nand U15917 (N_15917,N_15432,N_15312);
nor U15918 (N_15918,N_15568,N_15525);
and U15919 (N_15919,N_15381,N_15212);
nor U15920 (N_15920,N_15154,N_15499);
nand U15921 (N_15921,N_15366,N_15029);
xnor U15922 (N_15922,N_15375,N_15594);
or U15923 (N_15923,N_15030,N_15453);
nand U15924 (N_15924,N_15579,N_15176);
nor U15925 (N_15925,N_15206,N_15516);
nand U15926 (N_15926,N_15300,N_15106);
and U15927 (N_15927,N_15217,N_15545);
or U15928 (N_15928,N_15430,N_15580);
xor U15929 (N_15929,N_15007,N_15339);
or U15930 (N_15930,N_15291,N_15089);
xnor U15931 (N_15931,N_15436,N_15122);
nand U15932 (N_15932,N_15283,N_15048);
xnor U15933 (N_15933,N_15234,N_15253);
or U15934 (N_15934,N_15536,N_15174);
or U15935 (N_15935,N_15503,N_15437);
and U15936 (N_15936,N_15281,N_15303);
xor U15937 (N_15937,N_15022,N_15363);
and U15938 (N_15938,N_15229,N_15528);
or U15939 (N_15939,N_15570,N_15287);
and U15940 (N_15940,N_15587,N_15298);
xnor U15941 (N_15941,N_15573,N_15377);
or U15942 (N_15942,N_15019,N_15430);
or U15943 (N_15943,N_15522,N_15443);
nor U15944 (N_15944,N_15529,N_15199);
or U15945 (N_15945,N_15462,N_15329);
and U15946 (N_15946,N_15051,N_15242);
nand U15947 (N_15947,N_15512,N_15110);
xnor U15948 (N_15948,N_15206,N_15351);
nor U15949 (N_15949,N_15158,N_15526);
and U15950 (N_15950,N_15225,N_15335);
nor U15951 (N_15951,N_15327,N_15134);
or U15952 (N_15952,N_15481,N_15211);
nand U15953 (N_15953,N_15564,N_15136);
nand U15954 (N_15954,N_15325,N_15162);
nand U15955 (N_15955,N_15289,N_15449);
or U15956 (N_15956,N_15186,N_15484);
or U15957 (N_15957,N_15134,N_15104);
and U15958 (N_15958,N_15184,N_15398);
or U15959 (N_15959,N_15365,N_15268);
and U15960 (N_15960,N_15096,N_15283);
and U15961 (N_15961,N_15495,N_15278);
and U15962 (N_15962,N_15055,N_15334);
or U15963 (N_15963,N_15283,N_15454);
or U15964 (N_15964,N_15228,N_15285);
and U15965 (N_15965,N_15437,N_15455);
xnor U15966 (N_15966,N_15207,N_15529);
nand U15967 (N_15967,N_15040,N_15207);
xor U15968 (N_15968,N_15149,N_15048);
xnor U15969 (N_15969,N_15011,N_15378);
or U15970 (N_15970,N_15090,N_15263);
nor U15971 (N_15971,N_15566,N_15191);
and U15972 (N_15972,N_15165,N_15170);
xor U15973 (N_15973,N_15246,N_15140);
and U15974 (N_15974,N_15006,N_15336);
and U15975 (N_15975,N_15226,N_15552);
nand U15976 (N_15976,N_15009,N_15468);
or U15977 (N_15977,N_15018,N_15097);
nand U15978 (N_15978,N_15181,N_15093);
nor U15979 (N_15979,N_15492,N_15130);
or U15980 (N_15980,N_15077,N_15233);
nor U15981 (N_15981,N_15176,N_15348);
nor U15982 (N_15982,N_15587,N_15085);
xor U15983 (N_15983,N_15017,N_15463);
nand U15984 (N_15984,N_15195,N_15515);
or U15985 (N_15985,N_15569,N_15056);
nor U15986 (N_15986,N_15338,N_15318);
or U15987 (N_15987,N_15424,N_15383);
and U15988 (N_15988,N_15031,N_15573);
nor U15989 (N_15989,N_15296,N_15001);
xor U15990 (N_15990,N_15213,N_15336);
xnor U15991 (N_15991,N_15152,N_15096);
and U15992 (N_15992,N_15509,N_15124);
or U15993 (N_15993,N_15336,N_15285);
nor U15994 (N_15994,N_15443,N_15176);
xnor U15995 (N_15995,N_15247,N_15459);
xor U15996 (N_15996,N_15305,N_15331);
nand U15997 (N_15997,N_15134,N_15482);
or U15998 (N_15998,N_15163,N_15148);
and U15999 (N_15999,N_15311,N_15452);
nor U16000 (N_16000,N_15084,N_15484);
and U16001 (N_16001,N_15314,N_15327);
xnor U16002 (N_16002,N_15332,N_15009);
xnor U16003 (N_16003,N_15315,N_15146);
and U16004 (N_16004,N_15461,N_15230);
nor U16005 (N_16005,N_15497,N_15593);
nor U16006 (N_16006,N_15343,N_15416);
nand U16007 (N_16007,N_15204,N_15463);
xnor U16008 (N_16008,N_15221,N_15556);
nand U16009 (N_16009,N_15023,N_15244);
nor U16010 (N_16010,N_15434,N_15257);
nand U16011 (N_16011,N_15394,N_15350);
nand U16012 (N_16012,N_15393,N_15082);
and U16013 (N_16013,N_15532,N_15466);
nand U16014 (N_16014,N_15169,N_15519);
and U16015 (N_16015,N_15482,N_15323);
nor U16016 (N_16016,N_15352,N_15067);
nand U16017 (N_16017,N_15550,N_15446);
nor U16018 (N_16018,N_15512,N_15434);
or U16019 (N_16019,N_15359,N_15251);
or U16020 (N_16020,N_15570,N_15380);
and U16021 (N_16021,N_15450,N_15154);
and U16022 (N_16022,N_15117,N_15391);
and U16023 (N_16023,N_15344,N_15428);
and U16024 (N_16024,N_15058,N_15556);
and U16025 (N_16025,N_15473,N_15447);
nor U16026 (N_16026,N_15419,N_15091);
nand U16027 (N_16027,N_15585,N_15190);
and U16028 (N_16028,N_15038,N_15235);
nor U16029 (N_16029,N_15346,N_15360);
xnor U16030 (N_16030,N_15513,N_15306);
or U16031 (N_16031,N_15352,N_15338);
xor U16032 (N_16032,N_15200,N_15056);
nor U16033 (N_16033,N_15078,N_15018);
nor U16034 (N_16034,N_15409,N_15126);
nor U16035 (N_16035,N_15593,N_15185);
and U16036 (N_16036,N_15006,N_15427);
nor U16037 (N_16037,N_15292,N_15463);
nor U16038 (N_16038,N_15541,N_15422);
xnor U16039 (N_16039,N_15556,N_15039);
xnor U16040 (N_16040,N_15312,N_15401);
or U16041 (N_16041,N_15371,N_15408);
or U16042 (N_16042,N_15058,N_15054);
or U16043 (N_16043,N_15359,N_15311);
xor U16044 (N_16044,N_15399,N_15059);
xor U16045 (N_16045,N_15503,N_15247);
xnor U16046 (N_16046,N_15380,N_15015);
xor U16047 (N_16047,N_15487,N_15129);
xor U16048 (N_16048,N_15020,N_15059);
xor U16049 (N_16049,N_15301,N_15585);
and U16050 (N_16050,N_15410,N_15415);
or U16051 (N_16051,N_15475,N_15097);
nand U16052 (N_16052,N_15289,N_15017);
or U16053 (N_16053,N_15158,N_15073);
xnor U16054 (N_16054,N_15260,N_15359);
xnor U16055 (N_16055,N_15093,N_15564);
nor U16056 (N_16056,N_15479,N_15465);
nand U16057 (N_16057,N_15540,N_15457);
or U16058 (N_16058,N_15041,N_15088);
and U16059 (N_16059,N_15515,N_15537);
xor U16060 (N_16060,N_15374,N_15433);
xor U16061 (N_16061,N_15595,N_15074);
nand U16062 (N_16062,N_15186,N_15296);
and U16063 (N_16063,N_15055,N_15419);
and U16064 (N_16064,N_15212,N_15314);
nor U16065 (N_16065,N_15067,N_15526);
or U16066 (N_16066,N_15482,N_15118);
xor U16067 (N_16067,N_15483,N_15044);
nor U16068 (N_16068,N_15010,N_15072);
nand U16069 (N_16069,N_15570,N_15354);
or U16070 (N_16070,N_15459,N_15464);
and U16071 (N_16071,N_15164,N_15394);
and U16072 (N_16072,N_15579,N_15250);
nand U16073 (N_16073,N_15588,N_15273);
nand U16074 (N_16074,N_15362,N_15188);
nand U16075 (N_16075,N_15440,N_15486);
and U16076 (N_16076,N_15398,N_15490);
nand U16077 (N_16077,N_15105,N_15487);
and U16078 (N_16078,N_15221,N_15280);
xor U16079 (N_16079,N_15318,N_15558);
nor U16080 (N_16080,N_15169,N_15530);
or U16081 (N_16081,N_15155,N_15149);
and U16082 (N_16082,N_15585,N_15257);
and U16083 (N_16083,N_15271,N_15284);
and U16084 (N_16084,N_15123,N_15182);
nand U16085 (N_16085,N_15365,N_15547);
or U16086 (N_16086,N_15298,N_15330);
nor U16087 (N_16087,N_15468,N_15136);
or U16088 (N_16088,N_15522,N_15369);
xnor U16089 (N_16089,N_15168,N_15509);
and U16090 (N_16090,N_15218,N_15364);
and U16091 (N_16091,N_15057,N_15506);
and U16092 (N_16092,N_15067,N_15035);
xor U16093 (N_16093,N_15211,N_15190);
nor U16094 (N_16094,N_15495,N_15134);
and U16095 (N_16095,N_15097,N_15183);
nand U16096 (N_16096,N_15564,N_15232);
nand U16097 (N_16097,N_15129,N_15298);
xor U16098 (N_16098,N_15284,N_15436);
nor U16099 (N_16099,N_15050,N_15465);
nor U16100 (N_16100,N_15508,N_15326);
and U16101 (N_16101,N_15297,N_15448);
and U16102 (N_16102,N_15266,N_15359);
nand U16103 (N_16103,N_15199,N_15079);
nand U16104 (N_16104,N_15365,N_15516);
xor U16105 (N_16105,N_15003,N_15092);
nor U16106 (N_16106,N_15592,N_15575);
nand U16107 (N_16107,N_15102,N_15579);
or U16108 (N_16108,N_15492,N_15081);
and U16109 (N_16109,N_15598,N_15501);
nand U16110 (N_16110,N_15359,N_15585);
nand U16111 (N_16111,N_15289,N_15480);
or U16112 (N_16112,N_15311,N_15234);
nor U16113 (N_16113,N_15518,N_15515);
xor U16114 (N_16114,N_15124,N_15130);
and U16115 (N_16115,N_15186,N_15038);
xnor U16116 (N_16116,N_15228,N_15052);
or U16117 (N_16117,N_15223,N_15414);
or U16118 (N_16118,N_15018,N_15361);
nand U16119 (N_16119,N_15404,N_15375);
or U16120 (N_16120,N_15294,N_15065);
xnor U16121 (N_16121,N_15544,N_15207);
and U16122 (N_16122,N_15544,N_15360);
and U16123 (N_16123,N_15523,N_15545);
and U16124 (N_16124,N_15289,N_15580);
nor U16125 (N_16125,N_15311,N_15039);
nand U16126 (N_16126,N_15478,N_15292);
and U16127 (N_16127,N_15034,N_15581);
nor U16128 (N_16128,N_15136,N_15227);
nor U16129 (N_16129,N_15265,N_15190);
nor U16130 (N_16130,N_15592,N_15248);
and U16131 (N_16131,N_15186,N_15181);
nand U16132 (N_16132,N_15206,N_15484);
xnor U16133 (N_16133,N_15398,N_15327);
xor U16134 (N_16134,N_15368,N_15138);
or U16135 (N_16135,N_15586,N_15590);
and U16136 (N_16136,N_15245,N_15171);
xnor U16137 (N_16137,N_15321,N_15323);
or U16138 (N_16138,N_15387,N_15168);
xor U16139 (N_16139,N_15561,N_15149);
xnor U16140 (N_16140,N_15389,N_15216);
nor U16141 (N_16141,N_15540,N_15216);
nor U16142 (N_16142,N_15569,N_15166);
or U16143 (N_16143,N_15370,N_15446);
nor U16144 (N_16144,N_15093,N_15242);
and U16145 (N_16145,N_15102,N_15238);
or U16146 (N_16146,N_15506,N_15198);
nand U16147 (N_16147,N_15227,N_15029);
and U16148 (N_16148,N_15398,N_15015);
nor U16149 (N_16149,N_15045,N_15054);
or U16150 (N_16150,N_15030,N_15256);
xor U16151 (N_16151,N_15359,N_15037);
and U16152 (N_16152,N_15389,N_15044);
or U16153 (N_16153,N_15512,N_15227);
or U16154 (N_16154,N_15568,N_15528);
or U16155 (N_16155,N_15558,N_15412);
or U16156 (N_16156,N_15005,N_15428);
xnor U16157 (N_16157,N_15533,N_15472);
nand U16158 (N_16158,N_15109,N_15222);
xnor U16159 (N_16159,N_15178,N_15425);
nand U16160 (N_16160,N_15031,N_15495);
and U16161 (N_16161,N_15081,N_15314);
and U16162 (N_16162,N_15308,N_15319);
xor U16163 (N_16163,N_15314,N_15071);
nor U16164 (N_16164,N_15299,N_15451);
or U16165 (N_16165,N_15233,N_15216);
or U16166 (N_16166,N_15096,N_15421);
xnor U16167 (N_16167,N_15517,N_15288);
nor U16168 (N_16168,N_15267,N_15253);
nand U16169 (N_16169,N_15573,N_15078);
and U16170 (N_16170,N_15566,N_15521);
nor U16171 (N_16171,N_15492,N_15414);
xnor U16172 (N_16172,N_15323,N_15400);
nand U16173 (N_16173,N_15384,N_15234);
or U16174 (N_16174,N_15284,N_15463);
and U16175 (N_16175,N_15270,N_15348);
xor U16176 (N_16176,N_15111,N_15203);
and U16177 (N_16177,N_15135,N_15293);
nor U16178 (N_16178,N_15464,N_15234);
xor U16179 (N_16179,N_15203,N_15238);
and U16180 (N_16180,N_15106,N_15185);
nand U16181 (N_16181,N_15538,N_15334);
nand U16182 (N_16182,N_15477,N_15573);
nand U16183 (N_16183,N_15424,N_15077);
or U16184 (N_16184,N_15112,N_15174);
xor U16185 (N_16185,N_15435,N_15578);
nand U16186 (N_16186,N_15141,N_15588);
nand U16187 (N_16187,N_15356,N_15436);
nor U16188 (N_16188,N_15146,N_15504);
or U16189 (N_16189,N_15081,N_15257);
and U16190 (N_16190,N_15439,N_15005);
nor U16191 (N_16191,N_15242,N_15596);
and U16192 (N_16192,N_15200,N_15324);
xnor U16193 (N_16193,N_15165,N_15174);
nor U16194 (N_16194,N_15078,N_15258);
or U16195 (N_16195,N_15433,N_15197);
nand U16196 (N_16196,N_15191,N_15292);
nand U16197 (N_16197,N_15424,N_15001);
xor U16198 (N_16198,N_15212,N_15184);
nor U16199 (N_16199,N_15241,N_15410);
nor U16200 (N_16200,N_16125,N_15718);
nor U16201 (N_16201,N_16029,N_15762);
and U16202 (N_16202,N_16025,N_16196);
and U16203 (N_16203,N_15723,N_16011);
nand U16204 (N_16204,N_15659,N_15697);
nand U16205 (N_16205,N_15968,N_15800);
nor U16206 (N_16206,N_15758,N_16150);
and U16207 (N_16207,N_15747,N_15739);
or U16208 (N_16208,N_15828,N_16110);
nor U16209 (N_16209,N_15944,N_15716);
nor U16210 (N_16210,N_15887,N_15665);
and U16211 (N_16211,N_15662,N_15745);
and U16212 (N_16212,N_15982,N_16188);
nor U16213 (N_16213,N_15977,N_15640);
or U16214 (N_16214,N_16102,N_15954);
nor U16215 (N_16215,N_15965,N_15825);
and U16216 (N_16216,N_16006,N_15961);
and U16217 (N_16217,N_15600,N_16128);
and U16218 (N_16218,N_15811,N_15933);
nand U16219 (N_16219,N_15997,N_15724);
nand U16220 (N_16220,N_15930,N_16081);
and U16221 (N_16221,N_15787,N_15656);
xor U16222 (N_16222,N_15856,N_16065);
nand U16223 (N_16223,N_15689,N_16097);
xnor U16224 (N_16224,N_15920,N_15883);
nand U16225 (N_16225,N_15991,N_15637);
xnor U16226 (N_16226,N_15692,N_16005);
xor U16227 (N_16227,N_15975,N_15670);
or U16228 (N_16228,N_15629,N_16003);
nand U16229 (N_16229,N_16068,N_15704);
and U16230 (N_16230,N_16030,N_15885);
nor U16231 (N_16231,N_15831,N_15807);
or U16232 (N_16232,N_16108,N_16077);
nand U16233 (N_16233,N_15895,N_15868);
xnor U16234 (N_16234,N_16021,N_15642);
and U16235 (N_16235,N_16078,N_15632);
or U16236 (N_16236,N_15624,N_16140);
xnor U16237 (N_16237,N_16104,N_15789);
nor U16238 (N_16238,N_16000,N_15703);
xnor U16239 (N_16239,N_15879,N_15616);
xor U16240 (N_16240,N_16136,N_15936);
or U16241 (N_16241,N_15619,N_15748);
nand U16242 (N_16242,N_15668,N_15967);
and U16243 (N_16243,N_15791,N_16174);
nor U16244 (N_16244,N_16023,N_16126);
nor U16245 (N_16245,N_15765,N_15750);
xnor U16246 (N_16246,N_16033,N_16051);
nand U16247 (N_16247,N_15894,N_16020);
nand U16248 (N_16248,N_16056,N_15711);
xor U16249 (N_16249,N_16165,N_15666);
xnor U16250 (N_16250,N_15808,N_16139);
nand U16251 (N_16251,N_16083,N_15935);
and U16252 (N_16252,N_15925,N_15959);
or U16253 (N_16253,N_15706,N_16080);
nand U16254 (N_16254,N_16096,N_15679);
or U16255 (N_16255,N_15625,N_15976);
nand U16256 (N_16256,N_16154,N_16084);
or U16257 (N_16257,N_15648,N_15647);
and U16258 (N_16258,N_15804,N_15608);
nand U16259 (N_16259,N_16157,N_15915);
or U16260 (N_16260,N_15678,N_15881);
and U16261 (N_16261,N_15947,N_16058);
or U16262 (N_16262,N_15817,N_15966);
nor U16263 (N_16263,N_15902,N_15638);
xnor U16264 (N_16264,N_15712,N_15732);
or U16265 (N_16265,N_15777,N_16007);
and U16266 (N_16266,N_16131,N_15620);
and U16267 (N_16267,N_15633,N_15657);
nor U16268 (N_16268,N_15793,N_15859);
or U16269 (N_16269,N_16001,N_15972);
xor U16270 (N_16270,N_15645,N_15908);
and U16271 (N_16271,N_15676,N_15836);
or U16272 (N_16272,N_15761,N_16138);
and U16273 (N_16273,N_15612,N_15949);
nor U16274 (N_16274,N_16024,N_15864);
nor U16275 (N_16275,N_15722,N_16075);
nor U16276 (N_16276,N_15950,N_16141);
or U16277 (N_16277,N_15928,N_15960);
nand U16278 (N_16278,N_16124,N_15661);
or U16279 (N_16279,N_16060,N_16098);
and U16280 (N_16280,N_16090,N_15601);
xor U16281 (N_16281,N_16116,N_15698);
xnor U16282 (N_16282,N_15618,N_16105);
xor U16283 (N_16283,N_15771,N_16070);
or U16284 (N_16284,N_15713,N_15781);
or U16285 (N_16285,N_15896,N_15931);
nor U16286 (N_16286,N_15855,N_15844);
and U16287 (N_16287,N_15611,N_15847);
nor U16288 (N_16288,N_15820,N_15603);
and U16289 (N_16289,N_16019,N_15759);
and U16290 (N_16290,N_15801,N_15818);
and U16291 (N_16291,N_15866,N_15767);
nand U16292 (N_16292,N_15814,N_16197);
xnor U16293 (N_16293,N_16026,N_15622);
xor U16294 (N_16294,N_16153,N_15654);
or U16295 (N_16295,N_15687,N_15630);
and U16296 (N_16296,N_16155,N_16066);
nand U16297 (N_16297,N_15922,N_15742);
and U16298 (N_16298,N_16039,N_15770);
or U16299 (N_16299,N_16010,N_15970);
nor U16300 (N_16300,N_15727,N_15741);
nand U16301 (N_16301,N_15664,N_15663);
nor U16302 (N_16302,N_16179,N_15984);
and U16303 (N_16303,N_15606,N_15705);
xor U16304 (N_16304,N_15806,N_15918);
nor U16305 (N_16305,N_15822,N_15993);
or U16306 (N_16306,N_15812,N_16183);
nor U16307 (N_16307,N_15917,N_15614);
or U16308 (N_16308,N_15973,N_15851);
and U16309 (N_16309,N_15644,N_16107);
and U16310 (N_16310,N_15874,N_16144);
xor U16311 (N_16311,N_15821,N_15832);
nand U16312 (N_16312,N_16067,N_16008);
and U16313 (N_16313,N_15990,N_16017);
and U16314 (N_16314,N_15962,N_16094);
nor U16315 (N_16315,N_16135,N_15938);
nand U16316 (N_16316,N_15914,N_16162);
nor U16317 (N_16317,N_15901,N_15802);
or U16318 (N_16318,N_15652,N_16147);
or U16319 (N_16319,N_15730,N_16027);
or U16320 (N_16320,N_15833,N_16191);
nor U16321 (N_16321,N_16169,N_15751);
and U16322 (N_16322,N_15980,N_16132);
or U16323 (N_16323,N_15953,N_15913);
and U16324 (N_16324,N_15850,N_15726);
nand U16325 (N_16325,N_15904,N_16182);
nand U16326 (N_16326,N_15681,N_15686);
and U16327 (N_16327,N_15823,N_15658);
and U16328 (N_16328,N_16115,N_15744);
xor U16329 (N_16329,N_15969,N_16091);
xor U16330 (N_16330,N_15701,N_15702);
and U16331 (N_16331,N_15983,N_15636);
and U16332 (N_16332,N_15923,N_16168);
nor U16333 (N_16333,N_16148,N_15769);
nand U16334 (N_16334,N_15815,N_15840);
nor U16335 (N_16335,N_15941,N_15905);
or U16336 (N_16336,N_15872,N_15862);
and U16337 (N_16337,N_16171,N_16178);
or U16338 (N_16338,N_16073,N_15786);
xnor U16339 (N_16339,N_16002,N_16031);
or U16340 (N_16340,N_15852,N_15911);
and U16341 (N_16341,N_15841,N_15774);
or U16342 (N_16342,N_16103,N_16170);
and U16343 (N_16343,N_16164,N_16069);
nand U16344 (N_16344,N_16184,N_16134);
nand U16345 (N_16345,N_15845,N_15684);
xnor U16346 (N_16346,N_16161,N_16145);
nor U16347 (N_16347,N_16095,N_15796);
xor U16348 (N_16348,N_15688,N_15870);
and U16349 (N_16349,N_16137,N_15860);
or U16350 (N_16350,N_16028,N_16158);
nor U16351 (N_16351,N_15631,N_16160);
xnor U16352 (N_16352,N_15753,N_15888);
nand U16353 (N_16353,N_16038,N_15733);
nand U16354 (N_16354,N_16130,N_16185);
nor U16355 (N_16355,N_15671,N_15782);
nand U16356 (N_16356,N_15999,N_15617);
nor U16357 (N_16357,N_15754,N_15846);
nor U16358 (N_16358,N_16035,N_15707);
nand U16359 (N_16359,N_15998,N_15956);
and U16360 (N_16360,N_16055,N_15857);
nand U16361 (N_16361,N_15865,N_15871);
and U16362 (N_16362,N_16085,N_15788);
nor U16363 (N_16363,N_15790,N_15623);
nand U16364 (N_16364,N_15734,N_15783);
and U16365 (N_16365,N_16129,N_16166);
xnor U16366 (N_16366,N_15964,N_15942);
nand U16367 (N_16367,N_15854,N_15910);
xnor U16368 (N_16368,N_15715,N_15912);
nand U16369 (N_16369,N_15667,N_16152);
xnor U16370 (N_16370,N_15626,N_15867);
nand U16371 (N_16371,N_15880,N_15963);
or U16372 (N_16372,N_16052,N_15696);
nand U16373 (N_16373,N_15669,N_16177);
nor U16374 (N_16374,N_16199,N_15985);
xnor U16375 (N_16375,N_15834,N_15853);
nand U16376 (N_16376,N_16195,N_16194);
nand U16377 (N_16377,N_15763,N_15877);
nand U16378 (N_16378,N_16181,N_15699);
nand U16379 (N_16379,N_15987,N_16187);
xor U16380 (N_16380,N_16089,N_15641);
or U16381 (N_16381,N_16004,N_15627);
nor U16382 (N_16382,N_15604,N_15773);
and U16383 (N_16383,N_15752,N_15869);
and U16384 (N_16384,N_15924,N_15639);
xor U16385 (N_16385,N_16079,N_15610);
xnor U16386 (N_16386,N_16142,N_15609);
nor U16387 (N_16387,N_16120,N_15779);
nand U16388 (N_16388,N_15809,N_15735);
or U16389 (N_16389,N_15842,N_16071);
nand U16390 (N_16390,N_15628,N_15655);
nand U16391 (N_16391,N_15673,N_16054);
xnor U16392 (N_16392,N_15943,N_15738);
and U16393 (N_16393,N_16193,N_16032);
or U16394 (N_16394,N_16044,N_15937);
nor U16395 (N_16395,N_15810,N_16059);
xnor U16396 (N_16396,N_15660,N_16053);
xor U16397 (N_16397,N_16046,N_15772);
nand U16398 (N_16398,N_16087,N_15978);
or U16399 (N_16399,N_15757,N_15677);
nand U16400 (N_16400,N_16167,N_15940);
xnor U16401 (N_16401,N_16076,N_15996);
and U16402 (N_16402,N_15951,N_15602);
nor U16403 (N_16403,N_15675,N_15994);
nand U16404 (N_16404,N_16156,N_15775);
nand U16405 (N_16405,N_16012,N_15691);
or U16406 (N_16406,N_15974,N_16016);
xor U16407 (N_16407,N_15919,N_16114);
and U16408 (N_16408,N_16189,N_16180);
and U16409 (N_16409,N_16042,N_16041);
nand U16410 (N_16410,N_15607,N_15721);
and U16411 (N_16411,N_15892,N_16050);
nand U16412 (N_16412,N_15875,N_15683);
or U16413 (N_16413,N_15634,N_15934);
nand U16414 (N_16414,N_16092,N_15952);
nand U16415 (N_16415,N_16113,N_16034);
xor U16416 (N_16416,N_16018,N_16043);
xnor U16417 (N_16417,N_15899,N_15717);
nor U16418 (N_16418,N_15643,N_16037);
xor U16419 (N_16419,N_16122,N_15981);
or U16420 (N_16420,N_16151,N_15876);
nor U16421 (N_16421,N_15737,N_15893);
nand U16422 (N_16422,N_16149,N_16015);
and U16423 (N_16423,N_15605,N_15979);
and U16424 (N_16424,N_15766,N_15653);
nand U16425 (N_16425,N_15685,N_15635);
xor U16426 (N_16426,N_16048,N_15794);
nand U16427 (N_16427,N_15740,N_15890);
or U16428 (N_16428,N_15903,N_15816);
or U16429 (N_16429,N_15958,N_16106);
nor U16430 (N_16430,N_15824,N_16121);
and U16431 (N_16431,N_16036,N_15955);
nor U16432 (N_16432,N_15995,N_15768);
nor U16433 (N_16433,N_16123,N_16100);
or U16434 (N_16434,N_15693,N_15926);
nand U16435 (N_16435,N_15615,N_15674);
xor U16436 (N_16436,N_15848,N_15785);
nor U16437 (N_16437,N_15829,N_16063);
or U16438 (N_16438,N_15792,N_15805);
nand U16439 (N_16439,N_16099,N_16013);
nor U16440 (N_16440,N_16045,N_15819);
or U16441 (N_16441,N_15843,N_15700);
or U16442 (N_16442,N_16101,N_15946);
and U16443 (N_16443,N_16093,N_16062);
xor U16444 (N_16444,N_15708,N_16061);
xnor U16445 (N_16445,N_15743,N_16074);
nor U16446 (N_16446,N_15989,N_15646);
or U16447 (N_16447,N_16049,N_16143);
xor U16448 (N_16448,N_15971,N_16186);
xor U16449 (N_16449,N_15945,N_15755);
xor U16450 (N_16450,N_16146,N_15719);
xnor U16451 (N_16451,N_15651,N_16175);
xor U16452 (N_16452,N_15690,N_15731);
xnor U16453 (N_16453,N_15986,N_16109);
xor U16454 (N_16454,N_15898,N_16040);
and U16455 (N_16455,N_15988,N_16072);
nor U16456 (N_16456,N_16111,N_15695);
nor U16457 (N_16457,N_16088,N_16163);
and U16458 (N_16458,N_16119,N_16192);
or U16459 (N_16459,N_16064,N_15839);
nor U16460 (N_16460,N_15830,N_16127);
nand U16461 (N_16461,N_15797,N_15882);
xnor U16462 (N_16462,N_15921,N_15650);
nor U16463 (N_16463,N_15798,N_15873);
or U16464 (N_16464,N_15886,N_16198);
nand U16465 (N_16465,N_15714,N_16173);
and U16466 (N_16466,N_16112,N_15725);
and U16467 (N_16467,N_15672,N_15621);
and U16468 (N_16468,N_16086,N_15826);
xor U16469 (N_16469,N_15929,N_15889);
nand U16470 (N_16470,N_15760,N_15897);
nand U16471 (N_16471,N_15728,N_15861);
xnor U16472 (N_16472,N_15900,N_15710);
or U16473 (N_16473,N_15932,N_15709);
and U16474 (N_16474,N_15764,N_15957);
xnor U16475 (N_16475,N_16057,N_15613);
or U16476 (N_16476,N_15891,N_15776);
or U16477 (N_16477,N_15849,N_15827);
or U16478 (N_16478,N_16118,N_15784);
and U16479 (N_16479,N_15906,N_15838);
or U16480 (N_16480,N_15736,N_16190);
nand U16481 (N_16481,N_15909,N_16133);
nand U16482 (N_16482,N_15992,N_16047);
and U16483 (N_16483,N_15756,N_15927);
or U16484 (N_16484,N_16022,N_15720);
nor U16485 (N_16485,N_15729,N_16082);
or U16486 (N_16486,N_15749,N_15939);
and U16487 (N_16487,N_15813,N_15858);
and U16488 (N_16488,N_15907,N_15835);
nor U16489 (N_16489,N_15863,N_15778);
or U16490 (N_16490,N_16117,N_16014);
and U16491 (N_16491,N_15682,N_15948);
xor U16492 (N_16492,N_15795,N_15694);
xor U16493 (N_16493,N_15837,N_16176);
nor U16494 (N_16494,N_15780,N_16009);
xor U16495 (N_16495,N_15878,N_16172);
nor U16496 (N_16496,N_15916,N_16159);
and U16497 (N_16497,N_15746,N_15649);
xor U16498 (N_16498,N_15884,N_15799);
and U16499 (N_16499,N_15680,N_15803);
or U16500 (N_16500,N_16098,N_15824);
xor U16501 (N_16501,N_16032,N_15928);
or U16502 (N_16502,N_15964,N_15849);
or U16503 (N_16503,N_15906,N_16052);
xor U16504 (N_16504,N_15944,N_16193);
xnor U16505 (N_16505,N_16066,N_15755);
and U16506 (N_16506,N_15808,N_15880);
nand U16507 (N_16507,N_15666,N_16007);
and U16508 (N_16508,N_16024,N_15652);
xnor U16509 (N_16509,N_15873,N_15901);
and U16510 (N_16510,N_15687,N_15998);
and U16511 (N_16511,N_16160,N_15963);
or U16512 (N_16512,N_15713,N_15625);
nor U16513 (N_16513,N_15665,N_16128);
or U16514 (N_16514,N_16008,N_15825);
nand U16515 (N_16515,N_15916,N_15945);
and U16516 (N_16516,N_15611,N_16112);
nor U16517 (N_16517,N_15924,N_16198);
or U16518 (N_16518,N_16077,N_16093);
or U16519 (N_16519,N_15643,N_15638);
or U16520 (N_16520,N_16090,N_15968);
xnor U16521 (N_16521,N_16068,N_15907);
xor U16522 (N_16522,N_16020,N_15732);
xnor U16523 (N_16523,N_16080,N_15904);
and U16524 (N_16524,N_15842,N_15616);
nand U16525 (N_16525,N_16141,N_15921);
nand U16526 (N_16526,N_15931,N_15962);
xnor U16527 (N_16527,N_16177,N_15840);
nor U16528 (N_16528,N_16037,N_15685);
and U16529 (N_16529,N_15846,N_15876);
nor U16530 (N_16530,N_16053,N_15601);
xnor U16531 (N_16531,N_16153,N_15686);
and U16532 (N_16532,N_15698,N_15778);
xnor U16533 (N_16533,N_16180,N_15872);
nand U16534 (N_16534,N_15696,N_15633);
or U16535 (N_16535,N_16129,N_16169);
nand U16536 (N_16536,N_15933,N_16032);
xnor U16537 (N_16537,N_15752,N_16126);
nand U16538 (N_16538,N_15663,N_15780);
and U16539 (N_16539,N_16101,N_15980);
nor U16540 (N_16540,N_15864,N_16139);
xor U16541 (N_16541,N_16063,N_15752);
nand U16542 (N_16542,N_15703,N_15990);
nor U16543 (N_16543,N_15845,N_15778);
and U16544 (N_16544,N_16000,N_16025);
and U16545 (N_16545,N_16023,N_15752);
and U16546 (N_16546,N_16062,N_15994);
nand U16547 (N_16547,N_15892,N_15898);
xnor U16548 (N_16548,N_15949,N_15968);
or U16549 (N_16549,N_15753,N_15995);
or U16550 (N_16550,N_16023,N_15974);
or U16551 (N_16551,N_16087,N_16183);
nand U16552 (N_16552,N_15763,N_16026);
nor U16553 (N_16553,N_15805,N_15829);
or U16554 (N_16554,N_16090,N_15772);
nand U16555 (N_16555,N_16118,N_15759);
nand U16556 (N_16556,N_16071,N_15801);
or U16557 (N_16557,N_16165,N_15663);
nand U16558 (N_16558,N_16039,N_16038);
and U16559 (N_16559,N_16099,N_16120);
nor U16560 (N_16560,N_15642,N_15910);
or U16561 (N_16561,N_15691,N_15603);
nand U16562 (N_16562,N_15712,N_15840);
nor U16563 (N_16563,N_16024,N_15707);
and U16564 (N_16564,N_15655,N_16076);
nor U16565 (N_16565,N_16161,N_15754);
xnor U16566 (N_16566,N_15731,N_15692);
or U16567 (N_16567,N_16144,N_15768);
nand U16568 (N_16568,N_15905,N_15619);
and U16569 (N_16569,N_16188,N_15867);
xor U16570 (N_16570,N_15846,N_16049);
xor U16571 (N_16571,N_15675,N_15739);
nor U16572 (N_16572,N_15716,N_15833);
or U16573 (N_16573,N_15831,N_15682);
xnor U16574 (N_16574,N_15753,N_15856);
nor U16575 (N_16575,N_15810,N_16030);
or U16576 (N_16576,N_15848,N_15679);
or U16577 (N_16577,N_16121,N_16177);
nor U16578 (N_16578,N_15688,N_16076);
or U16579 (N_16579,N_15653,N_16026);
and U16580 (N_16580,N_15849,N_15795);
nor U16581 (N_16581,N_15615,N_16037);
xnor U16582 (N_16582,N_16160,N_15623);
nand U16583 (N_16583,N_16027,N_15937);
nor U16584 (N_16584,N_16002,N_15745);
nand U16585 (N_16585,N_15679,N_16086);
nor U16586 (N_16586,N_15947,N_15702);
xnor U16587 (N_16587,N_15669,N_16151);
and U16588 (N_16588,N_16169,N_15774);
nand U16589 (N_16589,N_16092,N_16058);
xor U16590 (N_16590,N_16174,N_15853);
and U16591 (N_16591,N_15646,N_15726);
xnor U16592 (N_16592,N_16186,N_15992);
or U16593 (N_16593,N_15904,N_15807);
xnor U16594 (N_16594,N_15819,N_15933);
xnor U16595 (N_16595,N_15795,N_16087);
nor U16596 (N_16596,N_15955,N_15636);
nor U16597 (N_16597,N_15954,N_15766);
nand U16598 (N_16598,N_15955,N_16197);
xnor U16599 (N_16599,N_16132,N_16040);
or U16600 (N_16600,N_15656,N_15642);
or U16601 (N_16601,N_15806,N_16086);
nand U16602 (N_16602,N_16183,N_16118);
nand U16603 (N_16603,N_15705,N_15904);
nand U16604 (N_16604,N_15867,N_15697);
and U16605 (N_16605,N_15904,N_15998);
nand U16606 (N_16606,N_16030,N_16183);
nor U16607 (N_16607,N_15840,N_15854);
nor U16608 (N_16608,N_16109,N_15727);
or U16609 (N_16609,N_15751,N_15869);
and U16610 (N_16610,N_16078,N_16060);
nor U16611 (N_16611,N_16199,N_16166);
xor U16612 (N_16612,N_16164,N_15832);
nor U16613 (N_16613,N_16137,N_15992);
and U16614 (N_16614,N_15950,N_16087);
and U16615 (N_16615,N_15641,N_15722);
and U16616 (N_16616,N_15783,N_16073);
nor U16617 (N_16617,N_15939,N_16073);
xor U16618 (N_16618,N_16084,N_15866);
xor U16619 (N_16619,N_15664,N_15774);
nor U16620 (N_16620,N_15998,N_16182);
and U16621 (N_16621,N_16018,N_15716);
xnor U16622 (N_16622,N_15939,N_16129);
or U16623 (N_16623,N_15959,N_15934);
nor U16624 (N_16624,N_16068,N_16185);
nand U16625 (N_16625,N_16132,N_16096);
and U16626 (N_16626,N_16111,N_15641);
nand U16627 (N_16627,N_16132,N_16139);
xor U16628 (N_16628,N_15752,N_15947);
or U16629 (N_16629,N_15996,N_16026);
nor U16630 (N_16630,N_16057,N_15810);
xnor U16631 (N_16631,N_15818,N_16158);
xor U16632 (N_16632,N_15899,N_16034);
xnor U16633 (N_16633,N_15824,N_15878);
nor U16634 (N_16634,N_16004,N_15791);
nand U16635 (N_16635,N_15739,N_15649);
or U16636 (N_16636,N_16033,N_15925);
nor U16637 (N_16637,N_15688,N_15723);
xnor U16638 (N_16638,N_16047,N_16074);
and U16639 (N_16639,N_15933,N_15728);
and U16640 (N_16640,N_15903,N_16199);
xor U16641 (N_16641,N_15658,N_15781);
or U16642 (N_16642,N_15628,N_16076);
and U16643 (N_16643,N_15661,N_16011);
xor U16644 (N_16644,N_15986,N_16182);
and U16645 (N_16645,N_16117,N_16011);
xor U16646 (N_16646,N_15631,N_15782);
or U16647 (N_16647,N_15762,N_15878);
xor U16648 (N_16648,N_15792,N_15633);
xor U16649 (N_16649,N_16184,N_15722);
xnor U16650 (N_16650,N_15776,N_16118);
or U16651 (N_16651,N_16036,N_15702);
nand U16652 (N_16652,N_15852,N_16131);
and U16653 (N_16653,N_16061,N_15813);
nor U16654 (N_16654,N_15719,N_16148);
or U16655 (N_16655,N_15797,N_16184);
and U16656 (N_16656,N_15817,N_16009);
nand U16657 (N_16657,N_15996,N_15981);
nand U16658 (N_16658,N_16098,N_15865);
nor U16659 (N_16659,N_16002,N_15797);
xor U16660 (N_16660,N_15606,N_16196);
or U16661 (N_16661,N_15983,N_15970);
or U16662 (N_16662,N_15829,N_15762);
nand U16663 (N_16663,N_16156,N_15921);
xor U16664 (N_16664,N_15871,N_15617);
xnor U16665 (N_16665,N_15709,N_15836);
or U16666 (N_16666,N_16081,N_16157);
nor U16667 (N_16667,N_16193,N_15709);
nor U16668 (N_16668,N_16150,N_15902);
nand U16669 (N_16669,N_15801,N_15724);
or U16670 (N_16670,N_15747,N_15629);
nand U16671 (N_16671,N_16016,N_16128);
or U16672 (N_16672,N_15736,N_15963);
or U16673 (N_16673,N_16006,N_15627);
xor U16674 (N_16674,N_15728,N_15655);
or U16675 (N_16675,N_15884,N_16183);
xor U16676 (N_16676,N_15813,N_15782);
or U16677 (N_16677,N_15720,N_15796);
or U16678 (N_16678,N_15855,N_16126);
xnor U16679 (N_16679,N_16030,N_15662);
nand U16680 (N_16680,N_16014,N_15926);
xor U16681 (N_16681,N_16180,N_15618);
and U16682 (N_16682,N_15867,N_16111);
xnor U16683 (N_16683,N_16143,N_16117);
or U16684 (N_16684,N_16130,N_15986);
and U16685 (N_16685,N_15901,N_15671);
or U16686 (N_16686,N_16077,N_16096);
nand U16687 (N_16687,N_15736,N_15907);
or U16688 (N_16688,N_15808,N_15942);
and U16689 (N_16689,N_15745,N_15946);
xor U16690 (N_16690,N_15758,N_15943);
nand U16691 (N_16691,N_16090,N_16020);
or U16692 (N_16692,N_16199,N_15819);
nand U16693 (N_16693,N_15855,N_15919);
or U16694 (N_16694,N_15915,N_16039);
and U16695 (N_16695,N_15637,N_16023);
xnor U16696 (N_16696,N_15928,N_16077);
and U16697 (N_16697,N_15683,N_15610);
nor U16698 (N_16698,N_15788,N_15745);
or U16699 (N_16699,N_15827,N_16123);
nor U16700 (N_16700,N_15696,N_15885);
or U16701 (N_16701,N_15797,N_15815);
nand U16702 (N_16702,N_15775,N_15975);
and U16703 (N_16703,N_15977,N_15756);
or U16704 (N_16704,N_15772,N_15635);
and U16705 (N_16705,N_16010,N_15891);
xor U16706 (N_16706,N_16171,N_16045);
xnor U16707 (N_16707,N_15962,N_15790);
xor U16708 (N_16708,N_15626,N_15652);
xor U16709 (N_16709,N_15606,N_16057);
nor U16710 (N_16710,N_16106,N_15918);
nand U16711 (N_16711,N_16036,N_15853);
nor U16712 (N_16712,N_15939,N_16198);
nand U16713 (N_16713,N_15997,N_15751);
nor U16714 (N_16714,N_16172,N_15692);
nor U16715 (N_16715,N_15615,N_15858);
and U16716 (N_16716,N_15686,N_15882);
nor U16717 (N_16717,N_16077,N_16176);
nand U16718 (N_16718,N_16157,N_16162);
xor U16719 (N_16719,N_16037,N_16199);
nor U16720 (N_16720,N_16126,N_16076);
xnor U16721 (N_16721,N_15971,N_15691);
xor U16722 (N_16722,N_15830,N_15855);
xor U16723 (N_16723,N_15923,N_15985);
nand U16724 (N_16724,N_16025,N_16044);
and U16725 (N_16725,N_15715,N_15778);
nor U16726 (N_16726,N_15975,N_16052);
and U16727 (N_16727,N_16040,N_15907);
xnor U16728 (N_16728,N_16009,N_15662);
xor U16729 (N_16729,N_15736,N_15704);
and U16730 (N_16730,N_16036,N_15676);
or U16731 (N_16731,N_16100,N_15659);
xnor U16732 (N_16732,N_16065,N_16156);
nor U16733 (N_16733,N_15673,N_16170);
nor U16734 (N_16734,N_15714,N_15792);
xnor U16735 (N_16735,N_15679,N_15689);
nand U16736 (N_16736,N_15914,N_16029);
nor U16737 (N_16737,N_16125,N_15654);
or U16738 (N_16738,N_15639,N_15781);
nand U16739 (N_16739,N_15607,N_15831);
nor U16740 (N_16740,N_15951,N_15777);
and U16741 (N_16741,N_15864,N_15859);
xnor U16742 (N_16742,N_15977,N_15841);
nand U16743 (N_16743,N_15930,N_15863);
or U16744 (N_16744,N_15752,N_15873);
and U16745 (N_16745,N_15937,N_15867);
nor U16746 (N_16746,N_15693,N_16135);
xor U16747 (N_16747,N_16071,N_16081);
and U16748 (N_16748,N_15941,N_15843);
or U16749 (N_16749,N_15783,N_15905);
nor U16750 (N_16750,N_15814,N_15854);
nand U16751 (N_16751,N_15840,N_15891);
xor U16752 (N_16752,N_15826,N_15638);
or U16753 (N_16753,N_15946,N_15966);
and U16754 (N_16754,N_15960,N_15702);
or U16755 (N_16755,N_15858,N_16074);
nand U16756 (N_16756,N_15677,N_16050);
nand U16757 (N_16757,N_15606,N_15961);
or U16758 (N_16758,N_15796,N_15625);
or U16759 (N_16759,N_15924,N_15873);
and U16760 (N_16760,N_16157,N_16037);
or U16761 (N_16761,N_15652,N_15988);
nor U16762 (N_16762,N_15877,N_16137);
nand U16763 (N_16763,N_16195,N_15935);
xor U16764 (N_16764,N_15633,N_15993);
nand U16765 (N_16765,N_15788,N_15677);
nor U16766 (N_16766,N_15749,N_16051);
nor U16767 (N_16767,N_16095,N_15947);
nor U16768 (N_16768,N_15730,N_15919);
nor U16769 (N_16769,N_15915,N_16162);
or U16770 (N_16770,N_16021,N_15662);
nor U16771 (N_16771,N_16197,N_15602);
xor U16772 (N_16772,N_15982,N_15614);
and U16773 (N_16773,N_15694,N_16155);
and U16774 (N_16774,N_15867,N_15931);
xor U16775 (N_16775,N_16021,N_15925);
xor U16776 (N_16776,N_15823,N_15607);
or U16777 (N_16777,N_15780,N_16052);
and U16778 (N_16778,N_16008,N_15903);
or U16779 (N_16779,N_15605,N_16161);
or U16780 (N_16780,N_15621,N_15865);
nor U16781 (N_16781,N_15901,N_15794);
and U16782 (N_16782,N_16177,N_16062);
or U16783 (N_16783,N_15629,N_16025);
nor U16784 (N_16784,N_16061,N_16190);
nand U16785 (N_16785,N_15643,N_15654);
nand U16786 (N_16786,N_15649,N_15712);
xor U16787 (N_16787,N_15887,N_16108);
xnor U16788 (N_16788,N_16083,N_16116);
nand U16789 (N_16789,N_16132,N_16080);
and U16790 (N_16790,N_15837,N_16072);
nor U16791 (N_16791,N_16152,N_15683);
nand U16792 (N_16792,N_15952,N_16054);
xor U16793 (N_16793,N_15680,N_15797);
nor U16794 (N_16794,N_15696,N_15873);
and U16795 (N_16795,N_15987,N_16099);
xnor U16796 (N_16796,N_15633,N_15644);
and U16797 (N_16797,N_16135,N_15786);
nand U16798 (N_16798,N_15632,N_15820);
xor U16799 (N_16799,N_15936,N_15636);
or U16800 (N_16800,N_16499,N_16236);
nand U16801 (N_16801,N_16474,N_16773);
nor U16802 (N_16802,N_16368,N_16456);
nand U16803 (N_16803,N_16653,N_16636);
xnor U16804 (N_16804,N_16615,N_16362);
and U16805 (N_16805,N_16520,N_16411);
or U16806 (N_16806,N_16736,N_16742);
and U16807 (N_16807,N_16464,N_16300);
xnor U16808 (N_16808,N_16533,N_16574);
and U16809 (N_16809,N_16758,N_16232);
nor U16810 (N_16810,N_16702,N_16457);
nor U16811 (N_16811,N_16295,N_16496);
xnor U16812 (N_16812,N_16685,N_16307);
xor U16813 (N_16813,N_16481,N_16652);
nand U16814 (N_16814,N_16339,N_16479);
or U16815 (N_16815,N_16647,N_16202);
nor U16816 (N_16816,N_16747,N_16248);
nand U16817 (N_16817,N_16738,N_16537);
or U16818 (N_16818,N_16353,N_16666);
nor U16819 (N_16819,N_16483,N_16347);
nand U16820 (N_16820,N_16719,N_16571);
or U16821 (N_16821,N_16741,N_16507);
nor U16822 (N_16822,N_16687,N_16560);
nand U16823 (N_16823,N_16777,N_16468);
xnor U16824 (N_16824,N_16315,N_16254);
nor U16825 (N_16825,N_16421,N_16782);
and U16826 (N_16826,N_16354,N_16548);
xnor U16827 (N_16827,N_16577,N_16342);
xnor U16828 (N_16828,N_16604,N_16612);
xor U16829 (N_16829,N_16428,N_16691);
nor U16830 (N_16830,N_16509,N_16267);
nor U16831 (N_16831,N_16429,N_16262);
nand U16832 (N_16832,N_16542,N_16563);
nor U16833 (N_16833,N_16203,N_16288);
or U16834 (N_16834,N_16480,N_16466);
nor U16835 (N_16835,N_16422,N_16397);
and U16836 (N_16836,N_16442,N_16382);
or U16837 (N_16837,N_16283,N_16238);
and U16838 (N_16838,N_16761,N_16601);
nand U16839 (N_16839,N_16768,N_16472);
xnor U16840 (N_16840,N_16780,N_16299);
nor U16841 (N_16841,N_16745,N_16331);
nor U16842 (N_16842,N_16335,N_16642);
nor U16843 (N_16843,N_16541,N_16301);
or U16844 (N_16844,N_16448,N_16408);
xor U16845 (N_16845,N_16746,N_16625);
nor U16846 (N_16846,N_16484,N_16273);
or U16847 (N_16847,N_16486,N_16561);
xor U16848 (N_16848,N_16623,N_16371);
or U16849 (N_16849,N_16569,N_16207);
nor U16850 (N_16850,N_16646,N_16692);
xnor U16851 (N_16851,N_16495,N_16407);
nor U16852 (N_16852,N_16280,N_16565);
and U16853 (N_16853,N_16516,N_16359);
or U16854 (N_16854,N_16200,N_16425);
and U16855 (N_16855,N_16416,N_16266);
nor U16856 (N_16856,N_16690,N_16799);
or U16857 (N_16857,N_16364,N_16640);
or U16858 (N_16858,N_16680,N_16440);
and U16859 (N_16859,N_16224,N_16222);
nand U16860 (N_16860,N_16629,N_16297);
xor U16861 (N_16861,N_16729,N_16659);
nand U16862 (N_16862,N_16667,N_16504);
nor U16863 (N_16863,N_16554,N_16792);
nand U16864 (N_16864,N_16336,N_16555);
and U16865 (N_16865,N_16239,N_16264);
nand U16866 (N_16866,N_16375,N_16521);
nor U16867 (N_16867,N_16304,N_16695);
xnor U16868 (N_16868,N_16547,N_16643);
or U16869 (N_16869,N_16631,N_16426);
xor U16870 (N_16870,N_16570,N_16274);
or U16871 (N_16871,N_16488,N_16501);
or U16872 (N_16872,N_16400,N_16344);
nor U16873 (N_16873,N_16796,N_16357);
or U16874 (N_16874,N_16510,N_16229);
or U16875 (N_16875,N_16662,N_16205);
nor U16876 (N_16876,N_16409,N_16517);
xnor U16877 (N_16877,N_16784,N_16700);
xor U16878 (N_16878,N_16461,N_16259);
nor U16879 (N_16879,N_16449,N_16597);
and U16880 (N_16880,N_16716,N_16211);
and U16881 (N_16881,N_16663,N_16797);
nand U16882 (N_16882,N_16306,N_16582);
nand U16883 (N_16883,N_16762,N_16506);
xor U16884 (N_16884,N_16734,N_16728);
and U16885 (N_16885,N_16291,N_16584);
or U16886 (N_16886,N_16220,N_16753);
or U16887 (N_16887,N_16715,N_16226);
xnor U16888 (N_16888,N_16379,N_16208);
nand U16889 (N_16889,N_16607,N_16697);
or U16890 (N_16890,N_16723,N_16223);
or U16891 (N_16891,N_16630,N_16525);
xnor U16892 (N_16892,N_16531,N_16522);
or U16893 (N_16893,N_16462,N_16390);
and U16894 (N_16894,N_16559,N_16219);
nor U16895 (N_16895,N_16743,N_16387);
nand U16896 (N_16896,N_16536,N_16550);
xor U16897 (N_16897,N_16242,N_16739);
and U16898 (N_16898,N_16500,N_16764);
nor U16899 (N_16899,N_16599,N_16543);
nor U16900 (N_16900,N_16535,N_16343);
xnor U16901 (N_16901,N_16576,N_16385);
nand U16902 (N_16902,N_16527,N_16437);
nor U16903 (N_16903,N_16632,N_16614);
nand U16904 (N_16904,N_16671,N_16323);
nand U16905 (N_16905,N_16706,N_16727);
nand U16906 (N_16906,N_16774,N_16286);
nand U16907 (N_16907,N_16600,N_16318);
nor U16908 (N_16908,N_16750,N_16699);
xnor U16909 (N_16909,N_16228,N_16707);
nand U16910 (N_16910,N_16586,N_16406);
nor U16911 (N_16911,N_16635,N_16538);
xnor U16912 (N_16912,N_16319,N_16658);
nand U16913 (N_16913,N_16427,N_16491);
and U16914 (N_16914,N_16245,N_16595);
nand U16915 (N_16915,N_16515,N_16776);
nor U16916 (N_16916,N_16534,N_16502);
nor U16917 (N_16917,N_16514,N_16641);
or U16918 (N_16918,N_16443,N_16730);
or U16919 (N_16919,N_16526,N_16377);
xor U16920 (N_16920,N_16591,N_16770);
or U16921 (N_16921,N_16268,N_16735);
nand U16922 (N_16922,N_16580,N_16621);
xor U16923 (N_16923,N_16369,N_16712);
and U16924 (N_16924,N_16476,N_16511);
xnor U16925 (N_16925,N_16322,N_16217);
nor U16926 (N_16926,N_16677,N_16261);
nor U16927 (N_16927,N_16260,N_16613);
xor U16928 (N_16928,N_16794,N_16287);
nor U16929 (N_16929,N_16320,N_16453);
nand U16930 (N_16930,N_16206,N_16405);
nand U16931 (N_16931,N_16392,N_16754);
or U16932 (N_16932,N_16469,N_16786);
nand U16933 (N_16933,N_16272,N_16290);
nand U16934 (N_16934,N_16608,N_16626);
and U16935 (N_16935,N_16572,N_16308);
and U16936 (N_16936,N_16765,N_16269);
nor U16937 (N_16937,N_16657,N_16749);
and U16938 (N_16938,N_16767,N_16455);
nor U16939 (N_16939,N_16714,N_16328);
or U16940 (N_16940,N_16415,N_16413);
and U16941 (N_16941,N_16670,N_16241);
or U16942 (N_16942,N_16310,N_16540);
xnor U16943 (N_16943,N_16675,N_16446);
nand U16944 (N_16944,N_16490,N_16498);
nor U16945 (N_16945,N_16684,N_16381);
nor U16946 (N_16946,N_16494,N_16669);
nor U16947 (N_16947,N_16436,N_16573);
and U16948 (N_16948,N_16265,N_16737);
nand U16949 (N_16949,N_16530,N_16656);
or U16950 (N_16950,N_16282,N_16513);
or U16951 (N_16951,N_16759,N_16255);
nor U16952 (N_16952,N_16789,N_16294);
nor U16953 (N_16953,N_16578,N_16549);
nor U16954 (N_16954,N_16590,N_16771);
or U16955 (N_16955,N_16284,N_16620);
and U16956 (N_16956,N_16309,N_16341);
xnor U16957 (N_16957,N_16709,N_16338);
and U16958 (N_16958,N_16419,N_16726);
nand U16959 (N_16959,N_16602,N_16645);
nand U16960 (N_16960,N_16326,N_16346);
and U16961 (N_16961,N_16451,N_16505);
xnor U16962 (N_16962,N_16311,N_16790);
xnor U16963 (N_16963,N_16606,N_16694);
nor U16964 (N_16964,N_16722,N_16470);
xor U16965 (N_16965,N_16492,N_16611);
or U16966 (N_16966,N_16785,N_16367);
and U16967 (N_16967,N_16412,N_16682);
nor U16968 (N_16968,N_16444,N_16445);
and U16969 (N_16969,N_16258,N_16334);
nand U16970 (N_16970,N_16356,N_16637);
nand U16971 (N_16971,N_16650,N_16683);
and U16972 (N_16972,N_16313,N_16439);
nor U16973 (N_16973,N_16383,N_16724);
nor U16974 (N_16974,N_16558,N_16566);
nand U16975 (N_16975,N_16235,N_16234);
and U16976 (N_16976,N_16363,N_16698);
and U16977 (N_16977,N_16708,N_16783);
xnor U16978 (N_16978,N_16546,N_16775);
or U16979 (N_16979,N_16497,N_16388);
and U16980 (N_16980,N_16589,N_16579);
and U16981 (N_16981,N_16788,N_16686);
xor U16982 (N_16982,N_16348,N_16372);
or U16983 (N_16983,N_16703,N_16325);
xnor U16984 (N_16984,N_16477,N_16760);
nor U16985 (N_16985,N_16250,N_16655);
nand U16986 (N_16986,N_16345,N_16660);
or U16987 (N_16987,N_16493,N_16370);
nor U16988 (N_16988,N_16434,N_16705);
nor U16989 (N_16989,N_16376,N_16281);
xor U16990 (N_16990,N_16303,N_16596);
xor U16991 (N_16991,N_16633,N_16246);
xnor U16992 (N_16992,N_16556,N_16401);
nand U16993 (N_16993,N_16624,N_16545);
nor U16994 (N_16994,N_16718,N_16450);
nor U16995 (N_16995,N_16213,N_16337);
or U16996 (N_16996,N_16373,N_16748);
and U16997 (N_16997,N_16733,N_16247);
nor U16998 (N_16998,N_16414,N_16523);
and U16999 (N_16999,N_16508,N_16316);
xor U17000 (N_17000,N_16679,N_16619);
and U17001 (N_17001,N_16251,N_16676);
nor U17002 (N_17002,N_16399,N_16678);
nand U17003 (N_17003,N_16581,N_16798);
xnor U17004 (N_17004,N_16243,N_16214);
nor U17005 (N_17005,N_16435,N_16240);
and U17006 (N_17006,N_16324,N_16503);
and U17007 (N_17007,N_16418,N_16380);
and U17008 (N_17008,N_16330,N_16417);
and U17009 (N_17009,N_16471,N_16271);
xor U17010 (N_17010,N_16627,N_16398);
xnor U17011 (N_17011,N_16512,N_16673);
nand U17012 (N_17012,N_16756,N_16321);
and U17013 (N_17013,N_16423,N_16402);
nor U17014 (N_17014,N_16215,N_16696);
xor U17015 (N_17015,N_16672,N_16616);
or U17016 (N_17016,N_16433,N_16487);
xor U17017 (N_17017,N_16787,N_16575);
nand U17018 (N_17018,N_16644,N_16755);
nor U17019 (N_17019,N_16252,N_16651);
nand U17020 (N_17020,N_16622,N_16277);
xor U17021 (N_17021,N_16568,N_16366);
and U17022 (N_17022,N_16779,N_16279);
nor U17023 (N_17023,N_16664,N_16327);
xnor U17024 (N_17024,N_16351,N_16225);
or U17025 (N_17025,N_16430,N_16285);
xnor U17026 (N_17026,N_16532,N_16751);
xnor U17027 (N_17027,N_16275,N_16389);
or U17028 (N_17028,N_16420,N_16257);
xor U17029 (N_17029,N_16218,N_16314);
xnor U17030 (N_17030,N_16465,N_16233);
nand U17031 (N_17031,N_16795,N_16447);
nand U17032 (N_17032,N_16278,N_16473);
nand U17033 (N_17033,N_16610,N_16772);
or U17034 (N_17034,N_16587,N_16216);
nand U17035 (N_17035,N_16365,N_16529);
nor U17036 (N_17036,N_16778,N_16441);
xnor U17037 (N_17037,N_16350,N_16432);
and U17038 (N_17038,N_16617,N_16384);
nand U17039 (N_17039,N_16693,N_16594);
xnor U17040 (N_17040,N_16231,N_16209);
nand U17041 (N_17041,N_16360,N_16791);
and U17042 (N_17042,N_16544,N_16552);
or U17043 (N_17043,N_16564,N_16585);
nor U17044 (N_17044,N_16438,N_16263);
and U17045 (N_17045,N_16567,N_16649);
and U17046 (N_17046,N_16654,N_16270);
nor U17047 (N_17047,N_16221,N_16204);
nand U17048 (N_17048,N_16475,N_16638);
and U17049 (N_17049,N_16391,N_16244);
xor U17050 (N_17050,N_16603,N_16352);
or U17051 (N_17051,N_16661,N_16732);
or U17052 (N_17052,N_16355,N_16769);
xor U17053 (N_17053,N_16332,N_16312);
and U17054 (N_17054,N_16539,N_16648);
xor U17055 (N_17055,N_16557,N_16394);
nor U17056 (N_17056,N_16374,N_16210);
nor U17057 (N_17057,N_16721,N_16634);
or U17058 (N_17058,N_16249,N_16458);
or U17059 (N_17059,N_16340,N_16256);
nor U17060 (N_17060,N_16296,N_16227);
or U17061 (N_17061,N_16378,N_16665);
and U17062 (N_17062,N_16276,N_16752);
and U17063 (N_17063,N_16395,N_16689);
nand U17064 (N_17064,N_16793,N_16553);
nor U17065 (N_17065,N_16292,N_16519);
nor U17066 (N_17066,N_16302,N_16551);
and U17067 (N_17067,N_16766,N_16403);
or U17068 (N_17068,N_16681,N_16358);
or U17069 (N_17069,N_16212,N_16528);
or U17070 (N_17070,N_16463,N_16720);
nor U17071 (N_17071,N_16452,N_16593);
or U17072 (N_17072,N_16237,N_16740);
xnor U17073 (N_17073,N_16361,N_16478);
and U17074 (N_17074,N_16489,N_16725);
xor U17075 (N_17075,N_16592,N_16710);
xnor U17076 (N_17076,N_16460,N_16396);
and U17077 (N_17077,N_16588,N_16609);
or U17078 (N_17078,N_16618,N_16781);
and U17079 (N_17079,N_16598,N_16298);
nor U17080 (N_17080,N_16393,N_16562);
or U17081 (N_17081,N_16467,N_16431);
nand U17082 (N_17082,N_16485,N_16524);
nor U17083 (N_17083,N_16583,N_16701);
nand U17084 (N_17084,N_16688,N_16763);
nand U17085 (N_17085,N_16711,N_16482);
xnor U17086 (N_17086,N_16386,N_16713);
or U17087 (N_17087,N_16757,N_16201);
nand U17088 (N_17088,N_16329,N_16605);
xor U17089 (N_17089,N_16293,N_16639);
and U17090 (N_17090,N_16253,N_16230);
nand U17091 (N_17091,N_16305,N_16704);
nand U17092 (N_17092,N_16628,N_16731);
nor U17093 (N_17093,N_16349,N_16410);
and U17094 (N_17094,N_16668,N_16744);
xnor U17095 (N_17095,N_16518,N_16404);
nand U17096 (N_17096,N_16333,N_16674);
or U17097 (N_17097,N_16459,N_16424);
xnor U17098 (N_17098,N_16454,N_16317);
nand U17099 (N_17099,N_16717,N_16289);
or U17100 (N_17100,N_16273,N_16365);
nor U17101 (N_17101,N_16212,N_16428);
nand U17102 (N_17102,N_16694,N_16711);
nor U17103 (N_17103,N_16525,N_16357);
and U17104 (N_17104,N_16372,N_16682);
nor U17105 (N_17105,N_16748,N_16238);
nor U17106 (N_17106,N_16766,N_16504);
nand U17107 (N_17107,N_16641,N_16233);
nor U17108 (N_17108,N_16406,N_16290);
xor U17109 (N_17109,N_16578,N_16393);
nor U17110 (N_17110,N_16541,N_16443);
xor U17111 (N_17111,N_16633,N_16748);
and U17112 (N_17112,N_16352,N_16551);
xor U17113 (N_17113,N_16460,N_16722);
nor U17114 (N_17114,N_16256,N_16649);
and U17115 (N_17115,N_16435,N_16453);
nor U17116 (N_17116,N_16618,N_16383);
xnor U17117 (N_17117,N_16481,N_16308);
nor U17118 (N_17118,N_16247,N_16386);
nand U17119 (N_17119,N_16532,N_16488);
or U17120 (N_17120,N_16580,N_16429);
and U17121 (N_17121,N_16565,N_16474);
and U17122 (N_17122,N_16738,N_16586);
nand U17123 (N_17123,N_16254,N_16212);
nor U17124 (N_17124,N_16346,N_16299);
nor U17125 (N_17125,N_16638,N_16569);
xnor U17126 (N_17126,N_16696,N_16381);
nand U17127 (N_17127,N_16678,N_16444);
or U17128 (N_17128,N_16455,N_16478);
or U17129 (N_17129,N_16446,N_16206);
xor U17130 (N_17130,N_16396,N_16661);
xor U17131 (N_17131,N_16342,N_16656);
nand U17132 (N_17132,N_16327,N_16790);
and U17133 (N_17133,N_16784,N_16586);
xnor U17134 (N_17134,N_16373,N_16353);
or U17135 (N_17135,N_16417,N_16580);
or U17136 (N_17136,N_16575,N_16667);
or U17137 (N_17137,N_16744,N_16394);
and U17138 (N_17138,N_16446,N_16387);
xnor U17139 (N_17139,N_16646,N_16732);
nand U17140 (N_17140,N_16738,N_16573);
or U17141 (N_17141,N_16719,N_16203);
xnor U17142 (N_17142,N_16501,N_16249);
xnor U17143 (N_17143,N_16730,N_16253);
and U17144 (N_17144,N_16510,N_16417);
and U17145 (N_17145,N_16437,N_16306);
or U17146 (N_17146,N_16328,N_16285);
or U17147 (N_17147,N_16699,N_16769);
xnor U17148 (N_17148,N_16243,N_16615);
and U17149 (N_17149,N_16574,N_16424);
xnor U17150 (N_17150,N_16532,N_16514);
or U17151 (N_17151,N_16432,N_16749);
nand U17152 (N_17152,N_16506,N_16419);
and U17153 (N_17153,N_16745,N_16773);
xor U17154 (N_17154,N_16475,N_16704);
nand U17155 (N_17155,N_16453,N_16580);
nor U17156 (N_17156,N_16765,N_16230);
nor U17157 (N_17157,N_16536,N_16408);
nand U17158 (N_17158,N_16315,N_16435);
and U17159 (N_17159,N_16697,N_16408);
or U17160 (N_17160,N_16351,N_16499);
nand U17161 (N_17161,N_16346,N_16745);
xnor U17162 (N_17162,N_16754,N_16419);
nor U17163 (N_17163,N_16651,N_16343);
or U17164 (N_17164,N_16671,N_16662);
nand U17165 (N_17165,N_16696,N_16255);
nor U17166 (N_17166,N_16787,N_16580);
and U17167 (N_17167,N_16271,N_16440);
and U17168 (N_17168,N_16570,N_16644);
xor U17169 (N_17169,N_16593,N_16584);
xor U17170 (N_17170,N_16788,N_16457);
and U17171 (N_17171,N_16718,N_16381);
and U17172 (N_17172,N_16742,N_16651);
nand U17173 (N_17173,N_16514,N_16577);
nand U17174 (N_17174,N_16431,N_16670);
nor U17175 (N_17175,N_16680,N_16420);
or U17176 (N_17176,N_16408,N_16296);
xor U17177 (N_17177,N_16600,N_16503);
and U17178 (N_17178,N_16557,N_16519);
or U17179 (N_17179,N_16676,N_16738);
nand U17180 (N_17180,N_16601,N_16399);
nor U17181 (N_17181,N_16352,N_16436);
and U17182 (N_17182,N_16421,N_16300);
or U17183 (N_17183,N_16780,N_16504);
xor U17184 (N_17184,N_16778,N_16785);
or U17185 (N_17185,N_16604,N_16637);
nand U17186 (N_17186,N_16223,N_16730);
and U17187 (N_17187,N_16555,N_16512);
xnor U17188 (N_17188,N_16720,N_16523);
nor U17189 (N_17189,N_16210,N_16732);
nor U17190 (N_17190,N_16571,N_16692);
xor U17191 (N_17191,N_16532,N_16364);
xnor U17192 (N_17192,N_16504,N_16728);
nor U17193 (N_17193,N_16511,N_16525);
xnor U17194 (N_17194,N_16447,N_16775);
xnor U17195 (N_17195,N_16738,N_16482);
nor U17196 (N_17196,N_16775,N_16791);
or U17197 (N_17197,N_16233,N_16494);
nand U17198 (N_17198,N_16418,N_16323);
xnor U17199 (N_17199,N_16337,N_16649);
nor U17200 (N_17200,N_16764,N_16251);
xor U17201 (N_17201,N_16319,N_16646);
xnor U17202 (N_17202,N_16211,N_16247);
or U17203 (N_17203,N_16256,N_16275);
or U17204 (N_17204,N_16592,N_16486);
and U17205 (N_17205,N_16287,N_16687);
and U17206 (N_17206,N_16335,N_16243);
xnor U17207 (N_17207,N_16670,N_16625);
or U17208 (N_17208,N_16620,N_16275);
xor U17209 (N_17209,N_16360,N_16342);
xnor U17210 (N_17210,N_16586,N_16663);
nor U17211 (N_17211,N_16733,N_16493);
nor U17212 (N_17212,N_16599,N_16300);
or U17213 (N_17213,N_16531,N_16363);
nand U17214 (N_17214,N_16226,N_16778);
nand U17215 (N_17215,N_16635,N_16533);
nand U17216 (N_17216,N_16297,N_16318);
xor U17217 (N_17217,N_16385,N_16338);
or U17218 (N_17218,N_16780,N_16302);
nand U17219 (N_17219,N_16209,N_16594);
and U17220 (N_17220,N_16656,N_16301);
nand U17221 (N_17221,N_16590,N_16417);
or U17222 (N_17222,N_16369,N_16491);
xor U17223 (N_17223,N_16592,N_16715);
nor U17224 (N_17224,N_16647,N_16237);
nor U17225 (N_17225,N_16475,N_16479);
xor U17226 (N_17226,N_16486,N_16487);
nor U17227 (N_17227,N_16545,N_16437);
xor U17228 (N_17228,N_16556,N_16335);
xor U17229 (N_17229,N_16739,N_16503);
xnor U17230 (N_17230,N_16433,N_16584);
nor U17231 (N_17231,N_16320,N_16263);
and U17232 (N_17232,N_16459,N_16616);
or U17233 (N_17233,N_16562,N_16467);
nand U17234 (N_17234,N_16631,N_16427);
or U17235 (N_17235,N_16344,N_16208);
xnor U17236 (N_17236,N_16408,N_16773);
nand U17237 (N_17237,N_16786,N_16411);
or U17238 (N_17238,N_16266,N_16337);
and U17239 (N_17239,N_16468,N_16605);
nor U17240 (N_17240,N_16577,N_16409);
nor U17241 (N_17241,N_16355,N_16309);
and U17242 (N_17242,N_16667,N_16389);
nor U17243 (N_17243,N_16546,N_16477);
or U17244 (N_17244,N_16523,N_16529);
nor U17245 (N_17245,N_16304,N_16787);
or U17246 (N_17246,N_16653,N_16377);
nand U17247 (N_17247,N_16330,N_16380);
or U17248 (N_17248,N_16682,N_16583);
and U17249 (N_17249,N_16698,N_16705);
nand U17250 (N_17250,N_16476,N_16251);
and U17251 (N_17251,N_16549,N_16455);
xor U17252 (N_17252,N_16735,N_16344);
xnor U17253 (N_17253,N_16722,N_16605);
nand U17254 (N_17254,N_16209,N_16317);
xor U17255 (N_17255,N_16593,N_16559);
and U17256 (N_17256,N_16707,N_16656);
and U17257 (N_17257,N_16540,N_16549);
nor U17258 (N_17258,N_16769,N_16596);
nor U17259 (N_17259,N_16287,N_16625);
and U17260 (N_17260,N_16742,N_16773);
nor U17261 (N_17261,N_16533,N_16720);
and U17262 (N_17262,N_16486,N_16431);
and U17263 (N_17263,N_16433,N_16497);
or U17264 (N_17264,N_16541,N_16775);
xor U17265 (N_17265,N_16788,N_16248);
nor U17266 (N_17266,N_16553,N_16317);
or U17267 (N_17267,N_16719,N_16701);
nand U17268 (N_17268,N_16634,N_16311);
nand U17269 (N_17269,N_16622,N_16575);
xnor U17270 (N_17270,N_16260,N_16564);
xnor U17271 (N_17271,N_16594,N_16635);
nand U17272 (N_17272,N_16353,N_16210);
xor U17273 (N_17273,N_16484,N_16350);
xor U17274 (N_17274,N_16386,N_16547);
and U17275 (N_17275,N_16271,N_16647);
xor U17276 (N_17276,N_16223,N_16739);
xnor U17277 (N_17277,N_16279,N_16208);
nand U17278 (N_17278,N_16585,N_16444);
nor U17279 (N_17279,N_16213,N_16427);
xor U17280 (N_17280,N_16791,N_16299);
and U17281 (N_17281,N_16484,N_16769);
and U17282 (N_17282,N_16504,N_16755);
nor U17283 (N_17283,N_16571,N_16478);
nor U17284 (N_17284,N_16615,N_16375);
or U17285 (N_17285,N_16293,N_16334);
nor U17286 (N_17286,N_16726,N_16693);
nand U17287 (N_17287,N_16771,N_16568);
xnor U17288 (N_17288,N_16552,N_16667);
nor U17289 (N_17289,N_16727,N_16254);
and U17290 (N_17290,N_16783,N_16391);
and U17291 (N_17291,N_16487,N_16594);
and U17292 (N_17292,N_16589,N_16326);
or U17293 (N_17293,N_16736,N_16766);
or U17294 (N_17294,N_16612,N_16773);
xor U17295 (N_17295,N_16420,N_16559);
or U17296 (N_17296,N_16328,N_16611);
or U17297 (N_17297,N_16354,N_16214);
and U17298 (N_17298,N_16399,N_16559);
and U17299 (N_17299,N_16309,N_16764);
or U17300 (N_17300,N_16599,N_16256);
or U17301 (N_17301,N_16267,N_16744);
and U17302 (N_17302,N_16460,N_16400);
and U17303 (N_17303,N_16387,N_16729);
or U17304 (N_17304,N_16482,N_16222);
or U17305 (N_17305,N_16275,N_16782);
nand U17306 (N_17306,N_16283,N_16391);
nor U17307 (N_17307,N_16445,N_16788);
xnor U17308 (N_17308,N_16511,N_16532);
nand U17309 (N_17309,N_16515,N_16576);
or U17310 (N_17310,N_16787,N_16453);
and U17311 (N_17311,N_16389,N_16636);
xor U17312 (N_17312,N_16213,N_16768);
nand U17313 (N_17313,N_16669,N_16795);
and U17314 (N_17314,N_16437,N_16652);
and U17315 (N_17315,N_16483,N_16666);
nand U17316 (N_17316,N_16725,N_16715);
xnor U17317 (N_17317,N_16673,N_16306);
or U17318 (N_17318,N_16462,N_16434);
nand U17319 (N_17319,N_16335,N_16492);
nand U17320 (N_17320,N_16391,N_16744);
nand U17321 (N_17321,N_16400,N_16749);
nand U17322 (N_17322,N_16729,N_16359);
and U17323 (N_17323,N_16552,N_16706);
and U17324 (N_17324,N_16445,N_16530);
or U17325 (N_17325,N_16423,N_16324);
xor U17326 (N_17326,N_16215,N_16444);
nor U17327 (N_17327,N_16763,N_16450);
xor U17328 (N_17328,N_16397,N_16200);
nand U17329 (N_17329,N_16415,N_16720);
nor U17330 (N_17330,N_16469,N_16732);
and U17331 (N_17331,N_16565,N_16607);
and U17332 (N_17332,N_16209,N_16679);
xnor U17333 (N_17333,N_16299,N_16660);
nor U17334 (N_17334,N_16241,N_16263);
and U17335 (N_17335,N_16612,N_16674);
nand U17336 (N_17336,N_16684,N_16707);
or U17337 (N_17337,N_16546,N_16595);
nand U17338 (N_17338,N_16689,N_16527);
and U17339 (N_17339,N_16792,N_16680);
and U17340 (N_17340,N_16701,N_16381);
nor U17341 (N_17341,N_16701,N_16278);
or U17342 (N_17342,N_16796,N_16669);
nor U17343 (N_17343,N_16374,N_16229);
or U17344 (N_17344,N_16738,N_16746);
xor U17345 (N_17345,N_16285,N_16344);
or U17346 (N_17346,N_16536,N_16432);
and U17347 (N_17347,N_16415,N_16629);
nand U17348 (N_17348,N_16381,N_16741);
nor U17349 (N_17349,N_16493,N_16628);
nor U17350 (N_17350,N_16492,N_16298);
or U17351 (N_17351,N_16501,N_16630);
or U17352 (N_17352,N_16661,N_16562);
or U17353 (N_17353,N_16206,N_16719);
xnor U17354 (N_17354,N_16490,N_16287);
xor U17355 (N_17355,N_16494,N_16585);
xnor U17356 (N_17356,N_16426,N_16574);
nor U17357 (N_17357,N_16281,N_16703);
xnor U17358 (N_17358,N_16585,N_16521);
nand U17359 (N_17359,N_16549,N_16697);
or U17360 (N_17360,N_16750,N_16744);
nand U17361 (N_17361,N_16652,N_16214);
or U17362 (N_17362,N_16778,N_16238);
or U17363 (N_17363,N_16350,N_16723);
nand U17364 (N_17364,N_16252,N_16611);
nand U17365 (N_17365,N_16216,N_16706);
nand U17366 (N_17366,N_16695,N_16433);
nand U17367 (N_17367,N_16616,N_16785);
nor U17368 (N_17368,N_16260,N_16448);
or U17369 (N_17369,N_16416,N_16758);
and U17370 (N_17370,N_16588,N_16388);
nor U17371 (N_17371,N_16388,N_16479);
and U17372 (N_17372,N_16288,N_16666);
nand U17373 (N_17373,N_16718,N_16468);
xnor U17374 (N_17374,N_16428,N_16404);
nand U17375 (N_17375,N_16362,N_16678);
xor U17376 (N_17376,N_16684,N_16606);
and U17377 (N_17377,N_16778,N_16777);
or U17378 (N_17378,N_16323,N_16622);
nand U17379 (N_17379,N_16682,N_16740);
and U17380 (N_17380,N_16649,N_16244);
nand U17381 (N_17381,N_16415,N_16470);
and U17382 (N_17382,N_16286,N_16397);
xor U17383 (N_17383,N_16669,N_16596);
nand U17384 (N_17384,N_16448,N_16498);
nor U17385 (N_17385,N_16496,N_16666);
and U17386 (N_17386,N_16693,N_16360);
nand U17387 (N_17387,N_16265,N_16440);
nand U17388 (N_17388,N_16375,N_16291);
nor U17389 (N_17389,N_16554,N_16508);
or U17390 (N_17390,N_16318,N_16407);
and U17391 (N_17391,N_16546,N_16498);
or U17392 (N_17392,N_16695,N_16528);
and U17393 (N_17393,N_16226,N_16231);
and U17394 (N_17394,N_16418,N_16690);
nand U17395 (N_17395,N_16403,N_16404);
nand U17396 (N_17396,N_16433,N_16686);
or U17397 (N_17397,N_16255,N_16663);
xor U17398 (N_17398,N_16299,N_16631);
or U17399 (N_17399,N_16644,N_16213);
nand U17400 (N_17400,N_16879,N_16827);
nand U17401 (N_17401,N_17304,N_17256);
xor U17402 (N_17402,N_17034,N_17270);
nand U17403 (N_17403,N_17220,N_16808);
nand U17404 (N_17404,N_17147,N_16815);
or U17405 (N_17405,N_17002,N_17262);
and U17406 (N_17406,N_17389,N_17377);
and U17407 (N_17407,N_17068,N_17066);
and U17408 (N_17408,N_17239,N_17072);
nor U17409 (N_17409,N_16968,N_16922);
and U17410 (N_17410,N_16969,N_17395);
xnor U17411 (N_17411,N_17014,N_17314);
or U17412 (N_17412,N_17114,N_16987);
nor U17413 (N_17413,N_16941,N_17214);
and U17414 (N_17414,N_17388,N_16932);
xnor U17415 (N_17415,N_17201,N_17298);
xnor U17416 (N_17416,N_16837,N_17120);
or U17417 (N_17417,N_17022,N_17370);
nor U17418 (N_17418,N_17382,N_17101);
and U17419 (N_17419,N_16954,N_17309);
and U17420 (N_17420,N_16972,N_17065);
xor U17421 (N_17421,N_17040,N_17087);
and U17422 (N_17422,N_17296,N_17209);
nor U17423 (N_17423,N_17153,N_17000);
nor U17424 (N_17424,N_17380,N_16908);
and U17425 (N_17425,N_17236,N_16807);
and U17426 (N_17426,N_17017,N_16855);
nand U17427 (N_17427,N_17045,N_17145);
or U17428 (N_17428,N_17108,N_17143);
or U17429 (N_17429,N_16848,N_16959);
or U17430 (N_17430,N_16897,N_17289);
or U17431 (N_17431,N_17356,N_17316);
nor U17432 (N_17432,N_16921,N_17267);
nor U17433 (N_17433,N_17302,N_16812);
xnor U17434 (N_17434,N_17275,N_17124);
xor U17435 (N_17435,N_17286,N_16814);
nand U17436 (N_17436,N_17182,N_17266);
and U17437 (N_17437,N_17190,N_17333);
xor U17438 (N_17438,N_17300,N_17225);
nor U17439 (N_17439,N_17295,N_17217);
or U17440 (N_17440,N_17037,N_16952);
or U17441 (N_17441,N_17144,N_17195);
or U17442 (N_17442,N_17176,N_17161);
nand U17443 (N_17443,N_17162,N_17142);
nor U17444 (N_17444,N_16974,N_17058);
nand U17445 (N_17445,N_17135,N_17131);
nor U17446 (N_17446,N_17028,N_16810);
xor U17447 (N_17447,N_16914,N_17375);
nand U17448 (N_17448,N_17369,N_16937);
nor U17449 (N_17449,N_17026,N_17320);
nor U17450 (N_17450,N_16945,N_16980);
and U17451 (N_17451,N_16940,N_17149);
or U17452 (N_17452,N_17328,N_17368);
or U17453 (N_17453,N_16989,N_17216);
nand U17454 (N_17454,N_17326,N_17310);
or U17455 (N_17455,N_17349,N_17245);
nor U17456 (N_17456,N_16834,N_17050);
xor U17457 (N_17457,N_17175,N_16833);
or U17458 (N_17458,N_17228,N_17129);
nand U17459 (N_17459,N_17152,N_17181);
nor U17460 (N_17460,N_17102,N_17027);
nand U17461 (N_17461,N_16894,N_16951);
xor U17462 (N_17462,N_17029,N_17252);
nand U17463 (N_17463,N_17079,N_17128);
xnor U17464 (N_17464,N_16900,N_16939);
and U17465 (N_17465,N_16902,N_16920);
xor U17466 (N_17466,N_17392,N_17387);
or U17467 (N_17467,N_17015,N_17139);
nand U17468 (N_17468,N_17242,N_16911);
xor U17469 (N_17469,N_17207,N_17018);
nand U17470 (N_17470,N_17154,N_17160);
nor U17471 (N_17471,N_17025,N_17170);
or U17472 (N_17472,N_16876,N_16956);
and U17473 (N_17473,N_17125,N_16806);
or U17474 (N_17474,N_17148,N_16963);
or U17475 (N_17475,N_17330,N_17339);
or U17476 (N_17476,N_17007,N_16899);
or U17477 (N_17477,N_16811,N_17321);
nor U17478 (N_17478,N_17200,N_17238);
nor U17479 (N_17479,N_17189,N_17227);
or U17480 (N_17480,N_16966,N_16846);
nor U17481 (N_17481,N_16817,N_17193);
nand U17482 (N_17482,N_16943,N_16985);
or U17483 (N_17483,N_16844,N_17350);
xnor U17484 (N_17484,N_17284,N_17095);
nand U17485 (N_17485,N_16988,N_16934);
nor U17486 (N_17486,N_16913,N_17036);
and U17487 (N_17487,N_16893,N_17071);
xnor U17488 (N_17488,N_16849,N_17011);
and U17489 (N_17489,N_17247,N_17269);
nand U17490 (N_17490,N_17010,N_17031);
nand U17491 (N_17491,N_16824,N_16975);
xor U17492 (N_17492,N_17255,N_17061);
nor U17493 (N_17493,N_17385,N_16884);
and U17494 (N_17494,N_16838,N_17042);
or U17495 (N_17495,N_17342,N_17064);
or U17496 (N_17496,N_17325,N_17276);
or U17497 (N_17497,N_16843,N_16878);
or U17498 (N_17498,N_17109,N_16821);
nor U17499 (N_17499,N_17273,N_16999);
xnor U17500 (N_17500,N_17136,N_17248);
xnor U17501 (N_17501,N_17005,N_16882);
nor U17502 (N_17502,N_16825,N_17244);
nor U17503 (N_17503,N_16829,N_17354);
nand U17504 (N_17504,N_17057,N_17035);
or U17505 (N_17505,N_17111,N_17078);
xnor U17506 (N_17506,N_16857,N_17218);
xor U17507 (N_17507,N_17106,N_16820);
nand U17508 (N_17508,N_16842,N_16978);
or U17509 (N_17509,N_17355,N_17331);
nor U17510 (N_17510,N_17063,N_17323);
nor U17511 (N_17511,N_17358,N_17223);
xor U17512 (N_17512,N_17197,N_17013);
nor U17513 (N_17513,N_17117,N_17023);
nor U17514 (N_17514,N_16930,N_16998);
nor U17515 (N_17515,N_17081,N_17317);
or U17516 (N_17516,N_17359,N_17279);
xor U17517 (N_17517,N_17059,N_17048);
and U17518 (N_17518,N_17032,N_17030);
xnor U17519 (N_17519,N_16991,N_17166);
nand U17520 (N_17520,N_17257,N_17287);
or U17521 (N_17521,N_17278,N_16986);
and U17522 (N_17522,N_17243,N_17096);
nor U17523 (N_17523,N_17335,N_17306);
and U17524 (N_17524,N_16979,N_17261);
or U17525 (N_17525,N_17047,N_17344);
xor U17526 (N_17526,N_16877,N_17232);
nor U17527 (N_17527,N_17092,N_17184);
nand U17528 (N_17528,N_17291,N_17250);
nand U17529 (N_17529,N_16868,N_17110);
and U17530 (N_17530,N_16931,N_17083);
and U17531 (N_17531,N_16905,N_17093);
xnor U17532 (N_17532,N_16892,N_17332);
nor U17533 (N_17533,N_17343,N_16896);
xnor U17534 (N_17534,N_17024,N_17240);
xor U17535 (N_17535,N_16936,N_16907);
xnor U17536 (N_17536,N_17126,N_17004);
xor U17537 (N_17537,N_16826,N_17060);
nand U17538 (N_17538,N_17386,N_17080);
or U17539 (N_17539,N_17288,N_16823);
nor U17540 (N_17540,N_17008,N_16990);
and U17541 (N_17541,N_17283,N_17215);
nand U17542 (N_17542,N_17378,N_17366);
nand U17543 (N_17543,N_17372,N_16935);
nor U17544 (N_17544,N_17222,N_17313);
or U17545 (N_17545,N_17196,N_16981);
nor U17546 (N_17546,N_16965,N_17324);
nor U17547 (N_17547,N_16906,N_16946);
xor U17548 (N_17548,N_16995,N_17353);
and U17549 (N_17549,N_17091,N_17089);
or U17550 (N_17550,N_17212,N_16866);
xnor U17551 (N_17551,N_16964,N_17177);
and U17552 (N_17552,N_17094,N_17163);
and U17553 (N_17553,N_17075,N_17169);
xor U17554 (N_17554,N_17351,N_16977);
or U17555 (N_17555,N_16867,N_16887);
xor U17556 (N_17556,N_17384,N_17338);
xnor U17557 (N_17557,N_16938,N_17088);
nor U17558 (N_17558,N_17246,N_17258);
and U17559 (N_17559,N_16996,N_17268);
and U17560 (N_17560,N_17186,N_16993);
nor U17561 (N_17561,N_16860,N_16872);
and U17562 (N_17562,N_17301,N_17103);
or U17563 (N_17563,N_16809,N_16927);
and U17564 (N_17564,N_17357,N_17188);
or U17565 (N_17565,N_16961,N_17318);
xnor U17566 (N_17566,N_17085,N_16851);
or U17567 (N_17567,N_16933,N_16865);
or U17568 (N_17568,N_17052,N_17006);
xor U17569 (N_17569,N_17345,N_17021);
nor U17570 (N_17570,N_17363,N_16863);
or U17571 (N_17571,N_17383,N_16830);
and U17572 (N_17572,N_17180,N_17107);
or U17573 (N_17573,N_17254,N_16929);
and U17574 (N_17574,N_17381,N_17155);
xor U17575 (N_17575,N_17046,N_16875);
xor U17576 (N_17576,N_16847,N_17168);
or U17577 (N_17577,N_17165,N_17334);
nor U17578 (N_17578,N_16973,N_17221);
xnor U17579 (N_17579,N_17192,N_16928);
and U17580 (N_17580,N_17077,N_17204);
or U17581 (N_17581,N_17230,N_16801);
or U17582 (N_17582,N_16955,N_17397);
xnor U17583 (N_17583,N_17082,N_17398);
and U17584 (N_17584,N_17271,N_16982);
nand U17585 (N_17585,N_17138,N_16828);
or U17586 (N_17586,N_17265,N_16871);
nor U17587 (N_17587,N_17293,N_17341);
or U17588 (N_17588,N_17098,N_17260);
nor U17589 (N_17589,N_16898,N_17185);
or U17590 (N_17590,N_17322,N_17253);
or U17591 (N_17591,N_17234,N_17062);
or U17592 (N_17592,N_17041,N_17167);
and U17593 (N_17593,N_16904,N_17157);
and U17594 (N_17594,N_16805,N_16850);
nand U17595 (N_17595,N_17127,N_17054);
and U17596 (N_17596,N_17116,N_16816);
and U17597 (N_17597,N_16992,N_16917);
or U17598 (N_17598,N_17150,N_17280);
xnor U17599 (N_17599,N_17235,N_17346);
and U17600 (N_17600,N_17376,N_17141);
xnor U17601 (N_17601,N_17019,N_16819);
nand U17602 (N_17602,N_17179,N_17074);
or U17603 (N_17603,N_17374,N_16891);
or U17604 (N_17604,N_16916,N_17277);
or U17605 (N_17605,N_17073,N_16802);
nor U17606 (N_17606,N_17274,N_17360);
nor U17607 (N_17607,N_16859,N_17105);
or U17608 (N_17608,N_16958,N_17053);
xor U17609 (N_17609,N_16912,N_16869);
nor U17610 (N_17610,N_17191,N_17249);
and U17611 (N_17611,N_17206,N_16861);
or U17612 (N_17612,N_16944,N_16924);
nand U17613 (N_17613,N_17122,N_17203);
or U17614 (N_17614,N_17224,N_17308);
or U17615 (N_17615,N_17361,N_16800);
nand U17616 (N_17616,N_16890,N_17208);
xnor U17617 (N_17617,N_17119,N_16854);
or U17618 (N_17618,N_17173,N_16957);
nand U17619 (N_17619,N_17329,N_17263);
and U17620 (N_17620,N_17140,N_16889);
or U17621 (N_17621,N_17132,N_16886);
or U17622 (N_17622,N_16983,N_17229);
nor U17623 (N_17623,N_16915,N_16839);
nor U17624 (N_17624,N_17039,N_16832);
nor U17625 (N_17625,N_16870,N_16895);
xor U17626 (N_17626,N_17210,N_17340);
nor U17627 (N_17627,N_16926,N_17202);
nor U17628 (N_17628,N_16910,N_17084);
nand U17629 (N_17629,N_17118,N_16918);
nand U17630 (N_17630,N_16881,N_17315);
and U17631 (N_17631,N_17146,N_17016);
xnor U17632 (N_17632,N_17159,N_17319);
xnor U17633 (N_17633,N_17151,N_17205);
nor U17634 (N_17634,N_17003,N_17373);
nand U17635 (N_17635,N_17049,N_17043);
nand U17636 (N_17636,N_17121,N_17158);
nor U17637 (N_17637,N_16942,N_17282);
and U17638 (N_17638,N_16804,N_17231);
nand U17639 (N_17639,N_17183,N_17038);
or U17640 (N_17640,N_17241,N_17307);
nor U17641 (N_17641,N_16836,N_17134);
nand U17642 (N_17642,N_16949,N_17113);
or U17643 (N_17643,N_16883,N_17367);
xnor U17644 (N_17644,N_17390,N_16947);
and U17645 (N_17645,N_17009,N_17393);
or U17646 (N_17646,N_17399,N_17090);
and U17647 (N_17647,N_16818,N_17104);
nand U17648 (N_17648,N_17194,N_17219);
or U17649 (N_17649,N_17379,N_16845);
nor U17650 (N_17650,N_17199,N_17281);
nor U17651 (N_17651,N_16971,N_17285);
and U17652 (N_17652,N_17211,N_17365);
and U17653 (N_17653,N_17264,N_17272);
and U17654 (N_17654,N_17137,N_17099);
and U17655 (N_17655,N_17051,N_17336);
or U17656 (N_17656,N_17178,N_17292);
xor U17657 (N_17657,N_17100,N_16853);
nor U17658 (N_17658,N_16858,N_17070);
nand U17659 (N_17659,N_16903,N_17371);
and U17660 (N_17660,N_17396,N_17187);
nor U17661 (N_17661,N_17312,N_17112);
and U17662 (N_17662,N_16953,N_17290);
nor U17663 (N_17663,N_17337,N_16835);
and U17664 (N_17664,N_17115,N_16841);
or U17665 (N_17665,N_17130,N_16948);
and U17666 (N_17666,N_17055,N_17123);
xor U17667 (N_17667,N_17174,N_17164);
nor U17668 (N_17668,N_17294,N_17352);
or U17669 (N_17669,N_16967,N_17076);
nand U17670 (N_17670,N_16901,N_16880);
or U17671 (N_17671,N_16885,N_16970);
nor U17672 (N_17672,N_16856,N_17226);
nand U17673 (N_17673,N_16888,N_16862);
nand U17674 (N_17674,N_17364,N_16909);
and U17675 (N_17675,N_16962,N_17133);
xor U17676 (N_17676,N_16874,N_17237);
nor U17677 (N_17677,N_16864,N_17348);
nor U17678 (N_17678,N_16831,N_17259);
and U17679 (N_17679,N_17251,N_17056);
nor U17680 (N_17680,N_16873,N_16925);
and U17681 (N_17681,N_16822,N_17086);
nor U17682 (N_17682,N_16976,N_17394);
or U17683 (N_17683,N_16803,N_17303);
and U17684 (N_17684,N_17044,N_17299);
nor U17685 (N_17685,N_17033,N_17069);
and U17686 (N_17686,N_17233,N_17305);
nor U17687 (N_17687,N_16950,N_17067);
nor U17688 (N_17688,N_17327,N_16813);
xor U17689 (N_17689,N_17391,N_17156);
or U17690 (N_17690,N_17012,N_16923);
or U17691 (N_17691,N_16919,N_16994);
xor U17692 (N_17692,N_17171,N_17311);
and U17693 (N_17693,N_17362,N_17297);
nor U17694 (N_17694,N_17213,N_17001);
nand U17695 (N_17695,N_17020,N_17347);
xnor U17696 (N_17696,N_17172,N_16997);
xor U17697 (N_17697,N_16960,N_17097);
nand U17698 (N_17698,N_17198,N_16984);
and U17699 (N_17699,N_16852,N_16840);
nor U17700 (N_17700,N_17077,N_17391);
and U17701 (N_17701,N_17043,N_17193);
or U17702 (N_17702,N_17114,N_16836);
nand U17703 (N_17703,N_16928,N_17318);
and U17704 (N_17704,N_17070,N_17230);
and U17705 (N_17705,N_16869,N_17053);
nor U17706 (N_17706,N_17134,N_16891);
and U17707 (N_17707,N_16838,N_17174);
nor U17708 (N_17708,N_17181,N_17106);
nor U17709 (N_17709,N_17301,N_16839);
nor U17710 (N_17710,N_17010,N_17032);
nor U17711 (N_17711,N_17202,N_17285);
nand U17712 (N_17712,N_16953,N_16827);
nand U17713 (N_17713,N_17336,N_17337);
or U17714 (N_17714,N_16822,N_17273);
nor U17715 (N_17715,N_17015,N_16934);
nor U17716 (N_17716,N_16808,N_17391);
nand U17717 (N_17717,N_17341,N_17313);
xnor U17718 (N_17718,N_17133,N_17243);
nor U17719 (N_17719,N_17192,N_17135);
and U17720 (N_17720,N_17191,N_16989);
or U17721 (N_17721,N_16903,N_17073);
or U17722 (N_17722,N_16838,N_17041);
nor U17723 (N_17723,N_16817,N_16981);
or U17724 (N_17724,N_16969,N_17321);
nand U17725 (N_17725,N_16984,N_17286);
or U17726 (N_17726,N_16985,N_16927);
or U17727 (N_17727,N_17131,N_17144);
and U17728 (N_17728,N_16949,N_17230);
nor U17729 (N_17729,N_17289,N_17123);
or U17730 (N_17730,N_17132,N_16810);
and U17731 (N_17731,N_17343,N_17093);
xnor U17732 (N_17732,N_17075,N_17353);
nand U17733 (N_17733,N_17313,N_17150);
xor U17734 (N_17734,N_16819,N_17054);
nor U17735 (N_17735,N_17038,N_17172);
nor U17736 (N_17736,N_17294,N_17227);
nor U17737 (N_17737,N_17276,N_17131);
nor U17738 (N_17738,N_16993,N_17058);
nand U17739 (N_17739,N_17230,N_16811);
and U17740 (N_17740,N_17199,N_17390);
nor U17741 (N_17741,N_17256,N_17029);
xor U17742 (N_17742,N_16941,N_17018);
nor U17743 (N_17743,N_16954,N_17348);
xnor U17744 (N_17744,N_17252,N_16919);
or U17745 (N_17745,N_17040,N_17341);
xnor U17746 (N_17746,N_17213,N_17335);
nand U17747 (N_17747,N_17112,N_17399);
or U17748 (N_17748,N_17252,N_17159);
or U17749 (N_17749,N_17140,N_17283);
and U17750 (N_17750,N_16910,N_17119);
or U17751 (N_17751,N_16863,N_16992);
nor U17752 (N_17752,N_17259,N_17366);
nor U17753 (N_17753,N_17208,N_17072);
xnor U17754 (N_17754,N_17021,N_17367);
xnor U17755 (N_17755,N_16864,N_17095);
or U17756 (N_17756,N_16933,N_17250);
or U17757 (N_17757,N_17123,N_17146);
and U17758 (N_17758,N_17001,N_16839);
and U17759 (N_17759,N_17152,N_16831);
nand U17760 (N_17760,N_17079,N_17384);
xnor U17761 (N_17761,N_16921,N_16977);
nor U17762 (N_17762,N_17070,N_17054);
nand U17763 (N_17763,N_17207,N_16829);
nand U17764 (N_17764,N_17237,N_17363);
xor U17765 (N_17765,N_17072,N_16804);
nand U17766 (N_17766,N_17137,N_17055);
or U17767 (N_17767,N_17354,N_16885);
xnor U17768 (N_17768,N_17012,N_16805);
xor U17769 (N_17769,N_17392,N_17046);
or U17770 (N_17770,N_16832,N_17222);
or U17771 (N_17771,N_17232,N_17253);
nand U17772 (N_17772,N_16848,N_17006);
nor U17773 (N_17773,N_17198,N_17297);
or U17774 (N_17774,N_16917,N_17089);
nand U17775 (N_17775,N_16827,N_16818);
xnor U17776 (N_17776,N_16972,N_17037);
or U17777 (N_17777,N_16982,N_16916);
nand U17778 (N_17778,N_17357,N_17246);
nand U17779 (N_17779,N_17229,N_17346);
nand U17780 (N_17780,N_16966,N_16945);
and U17781 (N_17781,N_17238,N_17250);
xor U17782 (N_17782,N_17073,N_17214);
and U17783 (N_17783,N_17387,N_17273);
xnor U17784 (N_17784,N_17046,N_17244);
nand U17785 (N_17785,N_17233,N_17214);
nor U17786 (N_17786,N_17254,N_17085);
and U17787 (N_17787,N_17086,N_16865);
nand U17788 (N_17788,N_17019,N_17002);
xnor U17789 (N_17789,N_17393,N_17047);
nor U17790 (N_17790,N_17237,N_17102);
nand U17791 (N_17791,N_17337,N_17153);
nand U17792 (N_17792,N_17057,N_17352);
nand U17793 (N_17793,N_17022,N_17049);
and U17794 (N_17794,N_17067,N_17104);
nor U17795 (N_17795,N_17011,N_17299);
nor U17796 (N_17796,N_17350,N_17177);
and U17797 (N_17797,N_17327,N_16963);
or U17798 (N_17798,N_16983,N_17304);
nor U17799 (N_17799,N_17313,N_16893);
nor U17800 (N_17800,N_16969,N_17135);
xnor U17801 (N_17801,N_17287,N_17123);
nor U17802 (N_17802,N_17032,N_17302);
xor U17803 (N_17803,N_16814,N_17356);
and U17804 (N_17804,N_17058,N_16832);
and U17805 (N_17805,N_16994,N_17138);
nand U17806 (N_17806,N_17252,N_16986);
xor U17807 (N_17807,N_16896,N_17334);
nand U17808 (N_17808,N_17023,N_17266);
or U17809 (N_17809,N_17041,N_17334);
and U17810 (N_17810,N_16876,N_16977);
nand U17811 (N_17811,N_17179,N_17300);
xor U17812 (N_17812,N_17051,N_17163);
xor U17813 (N_17813,N_17220,N_16877);
nand U17814 (N_17814,N_16986,N_16994);
and U17815 (N_17815,N_17317,N_16979);
and U17816 (N_17816,N_17233,N_17302);
and U17817 (N_17817,N_17251,N_17156);
nor U17818 (N_17818,N_17304,N_17247);
nor U17819 (N_17819,N_17247,N_17073);
or U17820 (N_17820,N_16876,N_17108);
and U17821 (N_17821,N_17095,N_16992);
nor U17822 (N_17822,N_17190,N_17140);
or U17823 (N_17823,N_17219,N_17021);
nand U17824 (N_17824,N_17368,N_16929);
nor U17825 (N_17825,N_17128,N_17026);
or U17826 (N_17826,N_17192,N_17319);
and U17827 (N_17827,N_16913,N_16822);
nor U17828 (N_17828,N_16936,N_16815);
or U17829 (N_17829,N_17303,N_17059);
xnor U17830 (N_17830,N_17095,N_17176);
nand U17831 (N_17831,N_17166,N_17280);
nor U17832 (N_17832,N_17152,N_17310);
or U17833 (N_17833,N_16993,N_17265);
nand U17834 (N_17834,N_16961,N_17214);
and U17835 (N_17835,N_17247,N_17123);
or U17836 (N_17836,N_17267,N_17362);
nand U17837 (N_17837,N_17245,N_16981);
nor U17838 (N_17838,N_17073,N_16817);
nand U17839 (N_17839,N_16857,N_17016);
or U17840 (N_17840,N_16858,N_17188);
and U17841 (N_17841,N_16908,N_17313);
or U17842 (N_17842,N_17198,N_17030);
and U17843 (N_17843,N_17209,N_16974);
and U17844 (N_17844,N_16893,N_16816);
and U17845 (N_17845,N_17137,N_17071);
nand U17846 (N_17846,N_17213,N_17239);
xor U17847 (N_17847,N_17206,N_16981);
xnor U17848 (N_17848,N_16997,N_17218);
and U17849 (N_17849,N_17058,N_17334);
nand U17850 (N_17850,N_17315,N_17092);
nand U17851 (N_17851,N_17058,N_16862);
xor U17852 (N_17852,N_17220,N_17103);
nand U17853 (N_17853,N_16854,N_17313);
xnor U17854 (N_17854,N_17169,N_17205);
or U17855 (N_17855,N_17384,N_16924);
xor U17856 (N_17856,N_17359,N_17352);
nor U17857 (N_17857,N_17102,N_17219);
nand U17858 (N_17858,N_17358,N_17276);
nor U17859 (N_17859,N_17287,N_17370);
or U17860 (N_17860,N_17348,N_17367);
xnor U17861 (N_17861,N_16903,N_16986);
nand U17862 (N_17862,N_17005,N_17361);
and U17863 (N_17863,N_17081,N_17393);
and U17864 (N_17864,N_17152,N_16808);
and U17865 (N_17865,N_17217,N_17267);
nor U17866 (N_17866,N_17318,N_16908);
nor U17867 (N_17867,N_16946,N_17332);
and U17868 (N_17868,N_17374,N_17362);
and U17869 (N_17869,N_17297,N_16927);
or U17870 (N_17870,N_17154,N_17369);
nand U17871 (N_17871,N_16862,N_17019);
xnor U17872 (N_17872,N_17201,N_17032);
nor U17873 (N_17873,N_17310,N_17099);
nor U17874 (N_17874,N_17073,N_17341);
nor U17875 (N_17875,N_17087,N_17312);
nand U17876 (N_17876,N_17376,N_17276);
or U17877 (N_17877,N_16933,N_17210);
nand U17878 (N_17878,N_16849,N_16840);
xor U17879 (N_17879,N_17388,N_17143);
nor U17880 (N_17880,N_17023,N_17066);
nor U17881 (N_17881,N_16960,N_17152);
and U17882 (N_17882,N_17145,N_16933);
nor U17883 (N_17883,N_17338,N_16983);
nor U17884 (N_17884,N_17372,N_17074);
nand U17885 (N_17885,N_17367,N_17315);
xor U17886 (N_17886,N_16829,N_17290);
and U17887 (N_17887,N_17303,N_17288);
or U17888 (N_17888,N_17349,N_16974);
and U17889 (N_17889,N_17034,N_16811);
nand U17890 (N_17890,N_17121,N_17311);
or U17891 (N_17891,N_16954,N_17263);
nand U17892 (N_17892,N_17301,N_17387);
xnor U17893 (N_17893,N_17281,N_16842);
xnor U17894 (N_17894,N_17310,N_17183);
xor U17895 (N_17895,N_17056,N_17285);
or U17896 (N_17896,N_17055,N_17374);
or U17897 (N_17897,N_17007,N_16941);
xor U17898 (N_17898,N_16936,N_17050);
nor U17899 (N_17899,N_17193,N_16905);
and U17900 (N_17900,N_16979,N_17231);
or U17901 (N_17901,N_17042,N_17056);
or U17902 (N_17902,N_16818,N_17291);
or U17903 (N_17903,N_17060,N_16842);
and U17904 (N_17904,N_16841,N_17365);
xnor U17905 (N_17905,N_17295,N_17106);
nor U17906 (N_17906,N_17355,N_16971);
and U17907 (N_17907,N_17037,N_17076);
xor U17908 (N_17908,N_17132,N_17196);
nor U17909 (N_17909,N_17127,N_17068);
xnor U17910 (N_17910,N_17135,N_16873);
xor U17911 (N_17911,N_16808,N_16841);
nand U17912 (N_17912,N_17157,N_17051);
nand U17913 (N_17913,N_17192,N_16944);
nor U17914 (N_17914,N_17310,N_16946);
nor U17915 (N_17915,N_17221,N_17314);
and U17916 (N_17916,N_16842,N_17231);
and U17917 (N_17917,N_17268,N_16905);
nor U17918 (N_17918,N_17352,N_17002);
and U17919 (N_17919,N_17106,N_17297);
and U17920 (N_17920,N_16826,N_17026);
xor U17921 (N_17921,N_17309,N_17026);
nor U17922 (N_17922,N_17121,N_17178);
nand U17923 (N_17923,N_16924,N_16807);
xnor U17924 (N_17924,N_16983,N_17177);
or U17925 (N_17925,N_16903,N_17044);
or U17926 (N_17926,N_17146,N_17091);
nor U17927 (N_17927,N_17208,N_16936);
nand U17928 (N_17928,N_17150,N_17394);
xnor U17929 (N_17929,N_17064,N_17311);
xor U17930 (N_17930,N_16812,N_17127);
or U17931 (N_17931,N_16811,N_16965);
or U17932 (N_17932,N_17084,N_16957);
nand U17933 (N_17933,N_16842,N_17328);
or U17934 (N_17934,N_17054,N_17344);
or U17935 (N_17935,N_16965,N_17022);
or U17936 (N_17936,N_17019,N_17133);
and U17937 (N_17937,N_17350,N_17392);
nand U17938 (N_17938,N_16992,N_16836);
and U17939 (N_17939,N_17322,N_16889);
nand U17940 (N_17940,N_17109,N_17354);
or U17941 (N_17941,N_16850,N_16820);
or U17942 (N_17942,N_17057,N_17159);
and U17943 (N_17943,N_16848,N_17075);
nand U17944 (N_17944,N_17132,N_16884);
xnor U17945 (N_17945,N_17238,N_17147);
xnor U17946 (N_17946,N_17221,N_17141);
and U17947 (N_17947,N_16896,N_16898);
nor U17948 (N_17948,N_16995,N_17133);
and U17949 (N_17949,N_17257,N_17134);
and U17950 (N_17950,N_17233,N_17296);
and U17951 (N_17951,N_17323,N_16831);
nand U17952 (N_17952,N_17076,N_17358);
or U17953 (N_17953,N_17208,N_17183);
and U17954 (N_17954,N_17386,N_17075);
nand U17955 (N_17955,N_17134,N_17029);
xor U17956 (N_17956,N_17186,N_17304);
nor U17957 (N_17957,N_17210,N_17241);
xor U17958 (N_17958,N_17294,N_17390);
xnor U17959 (N_17959,N_16913,N_17018);
xor U17960 (N_17960,N_17099,N_16901);
and U17961 (N_17961,N_17079,N_16898);
nand U17962 (N_17962,N_17340,N_17239);
nand U17963 (N_17963,N_17172,N_16843);
nand U17964 (N_17964,N_16890,N_17238);
xor U17965 (N_17965,N_17087,N_17202);
nor U17966 (N_17966,N_17268,N_17283);
xor U17967 (N_17967,N_17135,N_16917);
and U17968 (N_17968,N_17308,N_16970);
and U17969 (N_17969,N_16854,N_17210);
nor U17970 (N_17970,N_17085,N_17255);
and U17971 (N_17971,N_17035,N_16931);
or U17972 (N_17972,N_16899,N_17110);
xnor U17973 (N_17973,N_16889,N_17072);
or U17974 (N_17974,N_16880,N_17031);
and U17975 (N_17975,N_16839,N_17188);
nand U17976 (N_17976,N_17251,N_17348);
and U17977 (N_17977,N_16922,N_17316);
or U17978 (N_17978,N_16847,N_17077);
and U17979 (N_17979,N_17078,N_17202);
nand U17980 (N_17980,N_16864,N_17312);
xor U17981 (N_17981,N_16989,N_17026);
nand U17982 (N_17982,N_17304,N_17273);
nand U17983 (N_17983,N_17321,N_17303);
xor U17984 (N_17984,N_16872,N_17161);
or U17985 (N_17985,N_17095,N_16960);
or U17986 (N_17986,N_17260,N_17007);
and U17987 (N_17987,N_17307,N_16964);
and U17988 (N_17988,N_17384,N_16819);
nor U17989 (N_17989,N_17104,N_17177);
or U17990 (N_17990,N_17167,N_17002);
xnor U17991 (N_17991,N_17252,N_17342);
and U17992 (N_17992,N_16928,N_17039);
nand U17993 (N_17993,N_17300,N_17080);
nor U17994 (N_17994,N_17040,N_16918);
xnor U17995 (N_17995,N_17099,N_17320);
nand U17996 (N_17996,N_16980,N_17241);
nor U17997 (N_17997,N_16833,N_17274);
xnor U17998 (N_17998,N_17038,N_16910);
and U17999 (N_17999,N_17156,N_16854);
or U18000 (N_18000,N_17925,N_17721);
xor U18001 (N_18001,N_17496,N_17907);
nand U18002 (N_18002,N_17439,N_17586);
or U18003 (N_18003,N_17633,N_17477);
nand U18004 (N_18004,N_17951,N_17515);
nor U18005 (N_18005,N_17491,N_17433);
nor U18006 (N_18006,N_17603,N_17551);
xnor U18007 (N_18007,N_17738,N_17797);
nand U18008 (N_18008,N_17771,N_17632);
and U18009 (N_18009,N_17507,N_17517);
xor U18010 (N_18010,N_17548,N_17524);
nor U18011 (N_18011,N_17635,N_17823);
or U18012 (N_18012,N_17781,N_17802);
or U18013 (N_18013,N_17919,N_17564);
nand U18014 (N_18014,N_17735,N_17994);
nand U18015 (N_18015,N_17576,N_17931);
or U18016 (N_18016,N_17403,N_17930);
or U18017 (N_18017,N_17699,N_17530);
nor U18018 (N_18018,N_17875,N_17660);
xor U18019 (N_18019,N_17478,N_17813);
and U18020 (N_18020,N_17846,N_17655);
or U18021 (N_18021,N_17685,N_17918);
or U18022 (N_18022,N_17404,N_17844);
or U18023 (N_18023,N_17718,N_17816);
and U18024 (N_18024,N_17717,N_17670);
nor U18025 (N_18025,N_17622,N_17444);
xor U18026 (N_18026,N_17727,N_17619);
nand U18027 (N_18027,N_17973,N_17866);
nand U18028 (N_18028,N_17516,N_17805);
xnor U18029 (N_18029,N_17600,N_17522);
or U18030 (N_18030,N_17720,N_17833);
nor U18031 (N_18031,N_17598,N_17534);
and U18032 (N_18032,N_17452,N_17869);
nor U18033 (N_18033,N_17475,N_17443);
nor U18034 (N_18034,N_17687,N_17678);
and U18035 (N_18035,N_17894,N_17843);
nand U18036 (N_18036,N_17519,N_17476);
nand U18037 (N_18037,N_17957,N_17950);
nand U18038 (N_18038,N_17707,N_17725);
nor U18039 (N_18039,N_17594,N_17867);
and U18040 (N_18040,N_17640,N_17706);
and U18041 (N_18041,N_17750,N_17752);
and U18042 (N_18042,N_17856,N_17871);
and U18043 (N_18043,N_17803,N_17419);
xnor U18044 (N_18044,N_17520,N_17639);
and U18045 (N_18045,N_17913,N_17643);
or U18046 (N_18046,N_17641,N_17741);
nand U18047 (N_18047,N_17763,N_17479);
xor U18048 (N_18048,N_17512,N_17437);
or U18049 (N_18049,N_17722,N_17535);
nand U18050 (N_18050,N_17882,N_17588);
nor U18051 (N_18051,N_17523,N_17634);
or U18052 (N_18052,N_17665,N_17954);
xnor U18053 (N_18053,N_17703,N_17667);
nand U18054 (N_18054,N_17676,N_17458);
nor U18055 (N_18055,N_17502,N_17847);
nand U18056 (N_18056,N_17656,N_17653);
or U18057 (N_18057,N_17518,N_17447);
xnor U18058 (N_18058,N_17870,N_17784);
or U18059 (N_18059,N_17657,N_17956);
or U18060 (N_18060,N_17853,N_17506);
nand U18061 (N_18061,N_17441,N_17570);
and U18062 (N_18062,N_17465,N_17791);
or U18063 (N_18063,N_17495,N_17826);
nor U18064 (N_18064,N_17440,N_17932);
nor U18065 (N_18065,N_17609,N_17438);
nor U18066 (N_18066,N_17864,N_17448);
xor U18067 (N_18067,N_17769,N_17575);
xnor U18068 (N_18068,N_17605,N_17592);
or U18069 (N_18069,N_17645,N_17681);
and U18070 (N_18070,N_17662,N_17453);
nand U18071 (N_18071,N_17987,N_17577);
nor U18072 (N_18072,N_17415,N_17401);
nor U18073 (N_18073,N_17731,N_17877);
or U18074 (N_18074,N_17455,N_17786);
nand U18075 (N_18075,N_17513,N_17417);
nand U18076 (N_18076,N_17761,N_17568);
or U18077 (N_18077,N_17486,N_17400);
or U18078 (N_18078,N_17509,N_17531);
nor U18079 (N_18079,N_17481,N_17958);
nor U18080 (N_18080,N_17638,N_17658);
and U18081 (N_18081,N_17414,N_17546);
nand U18082 (N_18082,N_17471,N_17888);
or U18083 (N_18083,N_17528,N_17859);
and U18084 (N_18084,N_17514,N_17927);
nor U18085 (N_18085,N_17753,N_17792);
xor U18086 (N_18086,N_17719,N_17692);
nor U18087 (N_18087,N_17744,N_17664);
nand U18088 (N_18088,N_17916,N_17467);
and U18089 (N_18089,N_17412,N_17554);
and U18090 (N_18090,N_17601,N_17975);
and U18091 (N_18091,N_17651,N_17855);
and U18092 (N_18092,N_17505,N_17466);
xor U18093 (N_18093,N_17801,N_17745);
nand U18094 (N_18094,N_17830,N_17713);
xnor U18095 (N_18095,N_17608,N_17986);
nand U18096 (N_18096,N_17762,N_17759);
nor U18097 (N_18097,N_17860,N_17807);
nor U18098 (N_18098,N_17578,N_17972);
nor U18099 (N_18099,N_17616,N_17468);
or U18100 (N_18100,N_17914,N_17857);
xnor U18101 (N_18101,N_17470,N_17732);
and U18102 (N_18102,N_17760,N_17943);
or U18103 (N_18103,N_17607,N_17751);
xor U18104 (N_18104,N_17990,N_17945);
nand U18105 (N_18105,N_17566,N_17683);
xor U18106 (N_18106,N_17938,N_17572);
or U18107 (N_18107,N_17902,N_17911);
xor U18108 (N_18108,N_17937,N_17615);
or U18109 (N_18109,N_17898,N_17427);
or U18110 (N_18110,N_17776,N_17428);
nand U18111 (N_18111,N_17740,N_17899);
nor U18112 (N_18112,N_17777,N_17929);
or U18113 (N_18113,N_17672,N_17693);
nor U18114 (N_18114,N_17494,N_17689);
nand U18115 (N_18115,N_17891,N_17967);
or U18116 (N_18116,N_17739,N_17764);
nand U18117 (N_18117,N_17949,N_17818);
nor U18118 (N_18118,N_17828,N_17625);
nor U18119 (N_18119,N_17644,N_17984);
nor U18120 (N_18120,N_17728,N_17897);
xnor U18121 (N_18121,N_17964,N_17832);
xor U18122 (N_18122,N_17896,N_17454);
xor U18123 (N_18123,N_17538,N_17982);
nand U18124 (N_18124,N_17850,N_17593);
and U18125 (N_18125,N_17456,N_17880);
nand U18126 (N_18126,N_17749,N_17716);
or U18127 (N_18127,N_17473,N_17411);
xnor U18128 (N_18128,N_17980,N_17804);
or U18129 (N_18129,N_17827,N_17604);
nand U18130 (N_18130,N_17510,N_17695);
nand U18131 (N_18131,N_17539,N_17948);
or U18132 (N_18132,N_17773,N_17461);
nand U18133 (N_18133,N_17499,N_17557);
and U18134 (N_18134,N_17808,N_17410);
or U18135 (N_18135,N_17460,N_17574);
or U18136 (N_18136,N_17558,N_17445);
and U18137 (N_18137,N_17464,N_17977);
nand U18138 (N_18138,N_17733,N_17547);
nand U18139 (N_18139,N_17590,N_17597);
nor U18140 (N_18140,N_17583,N_17754);
or U18141 (N_18141,N_17878,N_17756);
nand U18142 (N_18142,N_17928,N_17571);
and U18143 (N_18143,N_17800,N_17407);
nand U18144 (N_18144,N_17862,N_17946);
xnor U18145 (N_18145,N_17734,N_17953);
xnor U18146 (N_18146,N_17966,N_17408);
nand U18147 (N_18147,N_17819,N_17431);
and U18148 (N_18148,N_17767,N_17527);
xnor U18149 (N_18149,N_17686,N_17999);
nor U18150 (N_18150,N_17936,N_17915);
or U18151 (N_18151,N_17924,N_17469);
and U18152 (N_18152,N_17831,N_17960);
xnor U18153 (N_18153,N_17874,N_17997);
xnor U18154 (N_18154,N_17965,N_17587);
nand U18155 (N_18155,N_17849,N_17562);
or U18156 (N_18156,N_17549,N_17650);
and U18157 (N_18157,N_17743,N_17556);
nand U18158 (N_18158,N_17611,N_17620);
nand U18159 (N_18159,N_17694,N_17446);
nor U18160 (N_18160,N_17774,N_17976);
nand U18161 (N_18161,N_17979,N_17544);
xor U18162 (N_18162,N_17947,N_17883);
nor U18163 (N_18163,N_17563,N_17579);
xnor U18164 (N_18164,N_17715,N_17941);
nand U18165 (N_18165,N_17785,N_17886);
or U18166 (N_18166,N_17796,N_17921);
and U18167 (N_18167,N_17591,N_17837);
or U18168 (N_18168,N_17698,N_17424);
and U18169 (N_18169,N_17559,N_17602);
or U18170 (N_18170,N_17508,N_17526);
nor U18171 (N_18171,N_17852,N_17906);
nand U18172 (N_18172,N_17910,N_17839);
nor U18173 (N_18173,N_17422,N_17712);
and U18174 (N_18174,N_17560,N_17962);
xnor U18175 (N_18175,N_17423,N_17810);
xor U18176 (N_18176,N_17669,N_17780);
nand U18177 (N_18177,N_17746,N_17736);
xnor U18178 (N_18178,N_17614,N_17459);
and U18179 (N_18179,N_17690,N_17868);
xnor U18180 (N_18180,N_17429,N_17895);
and U18181 (N_18181,N_17540,N_17908);
and U18182 (N_18182,N_17552,N_17606);
xor U18183 (N_18183,N_17790,N_17474);
and U18184 (N_18184,N_17617,N_17542);
nor U18185 (N_18185,N_17854,N_17498);
nor U18186 (N_18186,N_17696,N_17700);
and U18187 (N_18187,N_17865,N_17680);
nor U18188 (N_18188,N_17955,N_17425);
nor U18189 (N_18189,N_17580,N_17782);
xnor U18190 (N_18190,N_17613,N_17673);
nor U18191 (N_18191,N_17714,N_17770);
xor U18192 (N_18192,N_17532,N_17858);
nor U18193 (N_18193,N_17995,N_17783);
and U18194 (N_18194,N_17436,N_17890);
xnor U18195 (N_18195,N_17893,N_17942);
nor U18196 (N_18196,N_17820,N_17812);
nor U18197 (N_18197,N_17836,N_17684);
or U18198 (N_18198,N_17806,N_17472);
and U18199 (N_18199,N_17677,N_17905);
or U18200 (N_18200,N_17794,N_17497);
nor U18201 (N_18201,N_17450,N_17926);
xnor U18202 (N_18202,N_17585,N_17708);
nand U18203 (N_18203,N_17959,N_17789);
nor U18204 (N_18204,N_17485,N_17691);
and U18205 (N_18205,N_17900,N_17968);
or U18206 (N_18206,N_17838,N_17747);
nor U18207 (N_18207,N_17710,N_17674);
or U18208 (N_18208,N_17765,N_17726);
or U18209 (N_18209,N_17621,N_17565);
nand U18210 (N_18210,N_17503,N_17661);
or U18211 (N_18211,N_17876,N_17421);
and U18212 (N_18212,N_17969,N_17993);
xor U18213 (N_18213,N_17627,N_17406);
nand U18214 (N_18214,N_17861,N_17985);
and U18215 (N_18215,N_17541,N_17851);
and U18216 (N_18216,N_17996,N_17887);
or U18217 (N_18217,N_17755,N_17537);
and U18218 (N_18218,N_17920,N_17885);
nand U18219 (N_18219,N_17873,N_17817);
nand U18220 (N_18220,N_17775,N_17840);
and U18221 (N_18221,N_17841,N_17848);
nand U18222 (N_18222,N_17668,N_17798);
and U18223 (N_18223,N_17483,N_17405);
and U18224 (N_18224,N_17998,N_17724);
or U18225 (N_18225,N_17809,N_17647);
or U18226 (N_18226,N_17599,N_17659);
nand U18227 (N_18227,N_17500,N_17595);
and U18228 (N_18228,N_17729,N_17511);
xor U18229 (N_18229,N_17629,N_17567);
or U18230 (N_18230,N_17451,N_17663);
or U18231 (N_18231,N_17550,N_17766);
xor U18232 (N_18232,N_17799,N_17737);
and U18233 (N_18233,N_17788,N_17682);
nand U18234 (N_18234,N_17935,N_17487);
nand U18235 (N_18235,N_17493,N_17610);
or U18236 (N_18236,N_17702,N_17649);
and U18237 (N_18237,N_17845,N_17730);
or U18238 (N_18238,N_17795,N_17573);
nor U18239 (N_18239,N_17835,N_17418);
xnor U18240 (N_18240,N_17416,N_17778);
and U18241 (N_18241,N_17529,N_17757);
nor U18242 (N_18242,N_17654,N_17697);
nand U18243 (N_18243,N_17589,N_17909);
and U18244 (N_18244,N_17933,N_17675);
xor U18245 (N_18245,N_17628,N_17884);
and U18246 (N_18246,N_17904,N_17829);
and U18247 (N_18247,N_17889,N_17666);
nor U18248 (N_18248,N_17492,N_17709);
or U18249 (N_18249,N_17787,N_17779);
or U18250 (N_18250,N_17543,N_17811);
xor U18251 (N_18251,N_17630,N_17612);
xnor U18252 (N_18252,N_17569,N_17934);
xnor U18253 (N_18253,N_17923,N_17952);
nor U18254 (N_18254,N_17642,N_17912);
nor U18255 (N_18255,N_17521,N_17623);
nor U18256 (N_18256,N_17822,N_17992);
and U18257 (N_18257,N_17742,N_17705);
xnor U18258 (N_18258,N_17536,N_17978);
nor U18259 (N_18259,N_17704,N_17922);
nor U18260 (N_18260,N_17872,N_17501);
xnor U18261 (N_18261,N_17971,N_17903);
nand U18262 (N_18262,N_17974,N_17842);
nor U18263 (N_18263,N_17482,N_17701);
nor U18264 (N_18264,N_17723,N_17490);
nand U18265 (N_18265,N_17631,N_17626);
nand U18266 (N_18266,N_17462,N_17917);
nand U18267 (N_18267,N_17863,N_17545);
xor U18268 (N_18268,N_17793,N_17892);
or U18269 (N_18269,N_17409,N_17988);
and U18270 (N_18270,N_17480,N_17555);
or U18271 (N_18271,N_17434,N_17413);
and U18272 (N_18272,N_17636,N_17881);
or U18273 (N_18273,N_17768,N_17901);
nand U18274 (N_18274,N_17772,N_17679);
and U18275 (N_18275,N_17457,N_17940);
xor U18276 (N_18276,N_17646,N_17814);
xnor U18277 (N_18277,N_17970,N_17584);
xnor U18278 (N_18278,N_17671,N_17525);
and U18279 (N_18279,N_17981,N_17821);
xor U18280 (N_18280,N_17463,N_17533);
or U18281 (N_18281,N_17435,N_17989);
xor U18282 (N_18282,N_17825,N_17420);
nor U18283 (N_18283,N_17432,N_17504);
nor U18284 (N_18284,N_17624,N_17582);
and U18285 (N_18285,N_17402,N_17748);
or U18286 (N_18286,N_17488,N_17983);
nand U18287 (N_18287,N_17879,N_17939);
xnor U18288 (N_18288,N_17561,N_17815);
nand U18289 (N_18289,N_17944,N_17824);
and U18290 (N_18290,N_17430,N_17834);
nor U18291 (N_18291,N_17961,N_17596);
nand U18292 (N_18292,N_17426,N_17553);
or U18293 (N_18293,N_17758,N_17489);
xor U18294 (N_18294,N_17963,N_17581);
and U18295 (N_18295,N_17484,N_17991);
xor U18296 (N_18296,N_17449,N_17688);
nor U18297 (N_18297,N_17637,N_17442);
xor U18298 (N_18298,N_17618,N_17711);
xor U18299 (N_18299,N_17648,N_17652);
nand U18300 (N_18300,N_17932,N_17858);
nor U18301 (N_18301,N_17836,N_17632);
and U18302 (N_18302,N_17920,N_17466);
nand U18303 (N_18303,N_17856,N_17759);
nand U18304 (N_18304,N_17495,N_17588);
and U18305 (N_18305,N_17932,N_17619);
or U18306 (N_18306,N_17797,N_17852);
and U18307 (N_18307,N_17904,N_17891);
and U18308 (N_18308,N_17413,N_17857);
nand U18309 (N_18309,N_17992,N_17688);
nand U18310 (N_18310,N_17870,N_17739);
or U18311 (N_18311,N_17930,N_17777);
nor U18312 (N_18312,N_17470,N_17980);
and U18313 (N_18313,N_17620,N_17742);
nand U18314 (N_18314,N_17834,N_17421);
xor U18315 (N_18315,N_17630,N_17894);
nor U18316 (N_18316,N_17433,N_17635);
nor U18317 (N_18317,N_17683,N_17766);
nand U18318 (N_18318,N_17613,N_17878);
nand U18319 (N_18319,N_17644,N_17452);
xnor U18320 (N_18320,N_17584,N_17949);
and U18321 (N_18321,N_17901,N_17739);
or U18322 (N_18322,N_17657,N_17690);
nand U18323 (N_18323,N_17668,N_17725);
and U18324 (N_18324,N_17505,N_17899);
nor U18325 (N_18325,N_17534,N_17593);
nand U18326 (N_18326,N_17499,N_17596);
nor U18327 (N_18327,N_17494,N_17994);
and U18328 (N_18328,N_17706,N_17666);
or U18329 (N_18329,N_17681,N_17951);
or U18330 (N_18330,N_17789,N_17677);
or U18331 (N_18331,N_17582,N_17849);
xor U18332 (N_18332,N_17795,N_17539);
nor U18333 (N_18333,N_17979,N_17720);
nand U18334 (N_18334,N_17592,N_17940);
nand U18335 (N_18335,N_17670,N_17419);
and U18336 (N_18336,N_17624,N_17511);
nand U18337 (N_18337,N_17502,N_17423);
nor U18338 (N_18338,N_17756,N_17438);
nor U18339 (N_18339,N_17647,N_17944);
xnor U18340 (N_18340,N_17794,N_17927);
xor U18341 (N_18341,N_17506,N_17664);
or U18342 (N_18342,N_17734,N_17566);
or U18343 (N_18343,N_17677,N_17736);
nor U18344 (N_18344,N_17886,N_17723);
xor U18345 (N_18345,N_17656,N_17426);
or U18346 (N_18346,N_17833,N_17557);
nand U18347 (N_18347,N_17960,N_17666);
nand U18348 (N_18348,N_17906,N_17955);
and U18349 (N_18349,N_17497,N_17970);
and U18350 (N_18350,N_17477,N_17936);
nand U18351 (N_18351,N_17401,N_17928);
nand U18352 (N_18352,N_17874,N_17726);
nand U18353 (N_18353,N_17885,N_17537);
xor U18354 (N_18354,N_17750,N_17995);
nor U18355 (N_18355,N_17818,N_17723);
xor U18356 (N_18356,N_17842,N_17649);
nor U18357 (N_18357,N_17745,N_17589);
xnor U18358 (N_18358,N_17453,N_17690);
and U18359 (N_18359,N_17724,N_17715);
nor U18360 (N_18360,N_17536,N_17982);
xor U18361 (N_18361,N_17876,N_17933);
xor U18362 (N_18362,N_17918,N_17485);
and U18363 (N_18363,N_17945,N_17977);
nand U18364 (N_18364,N_17477,N_17600);
or U18365 (N_18365,N_17650,N_17541);
xnor U18366 (N_18366,N_17571,N_17435);
xor U18367 (N_18367,N_17695,N_17412);
and U18368 (N_18368,N_17528,N_17973);
and U18369 (N_18369,N_17832,N_17702);
and U18370 (N_18370,N_17967,N_17764);
nor U18371 (N_18371,N_17425,N_17728);
xor U18372 (N_18372,N_17900,N_17402);
or U18373 (N_18373,N_17535,N_17859);
or U18374 (N_18374,N_17661,N_17750);
nor U18375 (N_18375,N_17713,N_17825);
xnor U18376 (N_18376,N_17759,N_17461);
xor U18377 (N_18377,N_17419,N_17415);
nand U18378 (N_18378,N_17486,N_17802);
nor U18379 (N_18379,N_17997,N_17462);
nor U18380 (N_18380,N_17777,N_17825);
xnor U18381 (N_18381,N_17490,N_17630);
nand U18382 (N_18382,N_17489,N_17981);
xnor U18383 (N_18383,N_17518,N_17848);
nand U18384 (N_18384,N_17940,N_17954);
or U18385 (N_18385,N_17578,N_17924);
nand U18386 (N_18386,N_17936,N_17941);
or U18387 (N_18387,N_17453,N_17725);
and U18388 (N_18388,N_17405,N_17537);
nor U18389 (N_18389,N_17756,N_17735);
xnor U18390 (N_18390,N_17734,N_17563);
or U18391 (N_18391,N_17964,N_17732);
nand U18392 (N_18392,N_17513,N_17946);
nor U18393 (N_18393,N_17897,N_17947);
nor U18394 (N_18394,N_17858,N_17694);
nand U18395 (N_18395,N_17883,N_17542);
xnor U18396 (N_18396,N_17486,N_17510);
nand U18397 (N_18397,N_17733,N_17827);
xor U18398 (N_18398,N_17906,N_17772);
or U18399 (N_18399,N_17577,N_17982);
nand U18400 (N_18400,N_17453,N_17664);
or U18401 (N_18401,N_17775,N_17725);
xnor U18402 (N_18402,N_17882,N_17630);
nor U18403 (N_18403,N_17713,N_17952);
and U18404 (N_18404,N_17413,N_17637);
nand U18405 (N_18405,N_17617,N_17882);
xnor U18406 (N_18406,N_17525,N_17862);
xnor U18407 (N_18407,N_17456,N_17824);
xor U18408 (N_18408,N_17717,N_17908);
xnor U18409 (N_18409,N_17872,N_17467);
and U18410 (N_18410,N_17990,N_17562);
nor U18411 (N_18411,N_17525,N_17957);
nor U18412 (N_18412,N_17892,N_17781);
xor U18413 (N_18413,N_17456,N_17400);
or U18414 (N_18414,N_17780,N_17411);
xnor U18415 (N_18415,N_17979,N_17678);
or U18416 (N_18416,N_17643,N_17594);
nor U18417 (N_18417,N_17511,N_17996);
or U18418 (N_18418,N_17588,N_17547);
or U18419 (N_18419,N_17645,N_17611);
or U18420 (N_18420,N_17547,N_17623);
nand U18421 (N_18421,N_17997,N_17895);
and U18422 (N_18422,N_17960,N_17984);
nand U18423 (N_18423,N_17680,N_17896);
or U18424 (N_18424,N_17683,N_17892);
or U18425 (N_18425,N_17809,N_17856);
xor U18426 (N_18426,N_17789,N_17964);
xnor U18427 (N_18427,N_17413,N_17690);
or U18428 (N_18428,N_17809,N_17755);
or U18429 (N_18429,N_17585,N_17916);
nor U18430 (N_18430,N_17948,N_17921);
or U18431 (N_18431,N_17608,N_17467);
nor U18432 (N_18432,N_17927,N_17665);
xor U18433 (N_18433,N_17646,N_17747);
nor U18434 (N_18434,N_17474,N_17740);
nand U18435 (N_18435,N_17820,N_17489);
xor U18436 (N_18436,N_17836,N_17671);
xor U18437 (N_18437,N_17485,N_17503);
nand U18438 (N_18438,N_17663,N_17708);
xor U18439 (N_18439,N_17557,N_17664);
nor U18440 (N_18440,N_17918,N_17695);
xnor U18441 (N_18441,N_17402,N_17755);
nand U18442 (N_18442,N_17831,N_17914);
xnor U18443 (N_18443,N_17941,N_17537);
nor U18444 (N_18444,N_17742,N_17989);
or U18445 (N_18445,N_17858,N_17624);
or U18446 (N_18446,N_17611,N_17555);
nand U18447 (N_18447,N_17827,N_17922);
xor U18448 (N_18448,N_17628,N_17813);
or U18449 (N_18449,N_17864,N_17656);
or U18450 (N_18450,N_17753,N_17744);
nor U18451 (N_18451,N_17531,N_17780);
and U18452 (N_18452,N_17900,N_17413);
and U18453 (N_18453,N_17945,N_17860);
xnor U18454 (N_18454,N_17891,N_17459);
xnor U18455 (N_18455,N_17550,N_17783);
or U18456 (N_18456,N_17965,N_17739);
nor U18457 (N_18457,N_17534,N_17586);
or U18458 (N_18458,N_17496,N_17486);
nor U18459 (N_18459,N_17625,N_17691);
and U18460 (N_18460,N_17612,N_17800);
xor U18461 (N_18461,N_17844,N_17553);
xor U18462 (N_18462,N_17817,N_17608);
and U18463 (N_18463,N_17890,N_17404);
xnor U18464 (N_18464,N_17697,N_17956);
or U18465 (N_18465,N_17706,N_17860);
or U18466 (N_18466,N_17560,N_17720);
and U18467 (N_18467,N_17715,N_17862);
xnor U18468 (N_18468,N_17403,N_17400);
or U18469 (N_18469,N_17549,N_17732);
nand U18470 (N_18470,N_17743,N_17860);
and U18471 (N_18471,N_17618,N_17929);
nor U18472 (N_18472,N_17974,N_17833);
xor U18473 (N_18473,N_17985,N_17657);
and U18474 (N_18474,N_17446,N_17915);
or U18475 (N_18475,N_17924,N_17440);
and U18476 (N_18476,N_17809,N_17826);
and U18477 (N_18477,N_17693,N_17891);
nand U18478 (N_18478,N_17832,N_17719);
and U18479 (N_18479,N_17659,N_17540);
and U18480 (N_18480,N_17667,N_17912);
or U18481 (N_18481,N_17410,N_17692);
and U18482 (N_18482,N_17975,N_17626);
nand U18483 (N_18483,N_17619,N_17549);
and U18484 (N_18484,N_17714,N_17584);
and U18485 (N_18485,N_17495,N_17813);
xor U18486 (N_18486,N_17921,N_17588);
nand U18487 (N_18487,N_17493,N_17542);
nor U18488 (N_18488,N_17699,N_17603);
nor U18489 (N_18489,N_17468,N_17585);
nor U18490 (N_18490,N_17550,N_17808);
nor U18491 (N_18491,N_17766,N_17462);
nand U18492 (N_18492,N_17653,N_17799);
or U18493 (N_18493,N_17443,N_17899);
and U18494 (N_18494,N_17634,N_17766);
nor U18495 (N_18495,N_17997,N_17415);
xor U18496 (N_18496,N_17919,N_17981);
xor U18497 (N_18497,N_17652,N_17620);
nor U18498 (N_18498,N_17661,N_17906);
nor U18499 (N_18499,N_17403,N_17750);
xnor U18500 (N_18500,N_17851,N_17891);
or U18501 (N_18501,N_17905,N_17442);
nor U18502 (N_18502,N_17458,N_17745);
nand U18503 (N_18503,N_17622,N_17485);
or U18504 (N_18504,N_17621,N_17707);
nand U18505 (N_18505,N_17994,N_17590);
and U18506 (N_18506,N_17864,N_17890);
or U18507 (N_18507,N_17502,N_17441);
nand U18508 (N_18508,N_17952,N_17446);
or U18509 (N_18509,N_17496,N_17484);
xor U18510 (N_18510,N_17467,N_17588);
nand U18511 (N_18511,N_17803,N_17759);
nor U18512 (N_18512,N_17510,N_17432);
or U18513 (N_18513,N_17489,N_17711);
xnor U18514 (N_18514,N_17835,N_17430);
and U18515 (N_18515,N_17572,N_17579);
or U18516 (N_18516,N_17412,N_17418);
and U18517 (N_18517,N_17926,N_17683);
nor U18518 (N_18518,N_17658,N_17643);
nor U18519 (N_18519,N_17905,N_17491);
or U18520 (N_18520,N_17758,N_17637);
xnor U18521 (N_18521,N_17888,N_17423);
nor U18522 (N_18522,N_17895,N_17629);
or U18523 (N_18523,N_17925,N_17876);
xor U18524 (N_18524,N_17683,N_17838);
nand U18525 (N_18525,N_17742,N_17756);
nand U18526 (N_18526,N_17732,N_17910);
and U18527 (N_18527,N_17429,N_17823);
nand U18528 (N_18528,N_17469,N_17520);
xor U18529 (N_18529,N_17409,N_17589);
xor U18530 (N_18530,N_17615,N_17837);
xor U18531 (N_18531,N_17974,N_17769);
nand U18532 (N_18532,N_17469,N_17796);
nand U18533 (N_18533,N_17481,N_17842);
or U18534 (N_18534,N_17974,N_17647);
nand U18535 (N_18535,N_17806,N_17467);
and U18536 (N_18536,N_17647,N_17559);
and U18537 (N_18537,N_17596,N_17862);
nor U18538 (N_18538,N_17793,N_17983);
nand U18539 (N_18539,N_17716,N_17791);
or U18540 (N_18540,N_17470,N_17416);
or U18541 (N_18541,N_17534,N_17970);
xnor U18542 (N_18542,N_17688,N_17592);
nand U18543 (N_18543,N_17533,N_17544);
nor U18544 (N_18544,N_17686,N_17768);
and U18545 (N_18545,N_17956,N_17878);
xor U18546 (N_18546,N_17979,N_17523);
nor U18547 (N_18547,N_17982,N_17493);
nor U18548 (N_18548,N_17876,N_17949);
and U18549 (N_18549,N_17855,N_17481);
nor U18550 (N_18550,N_17962,N_17576);
nor U18551 (N_18551,N_17922,N_17719);
or U18552 (N_18552,N_17678,N_17884);
xnor U18553 (N_18553,N_17918,N_17434);
xnor U18554 (N_18554,N_17718,N_17995);
or U18555 (N_18555,N_17818,N_17781);
nand U18556 (N_18556,N_17838,N_17622);
nand U18557 (N_18557,N_17400,N_17947);
or U18558 (N_18558,N_17638,N_17403);
or U18559 (N_18559,N_17423,N_17400);
nand U18560 (N_18560,N_17719,N_17755);
nor U18561 (N_18561,N_17581,N_17599);
and U18562 (N_18562,N_17524,N_17972);
nor U18563 (N_18563,N_17451,N_17729);
xnor U18564 (N_18564,N_17778,N_17859);
nor U18565 (N_18565,N_17944,N_17403);
and U18566 (N_18566,N_17484,N_17417);
xor U18567 (N_18567,N_17951,N_17780);
and U18568 (N_18568,N_17803,N_17646);
nand U18569 (N_18569,N_17845,N_17534);
xnor U18570 (N_18570,N_17756,N_17625);
and U18571 (N_18571,N_17989,N_17772);
nor U18572 (N_18572,N_17802,N_17569);
nor U18573 (N_18573,N_17531,N_17957);
or U18574 (N_18574,N_17995,N_17519);
nand U18575 (N_18575,N_17957,N_17521);
or U18576 (N_18576,N_17977,N_17891);
or U18577 (N_18577,N_17902,N_17437);
and U18578 (N_18578,N_17509,N_17635);
and U18579 (N_18579,N_17691,N_17558);
nand U18580 (N_18580,N_17669,N_17622);
or U18581 (N_18581,N_17533,N_17782);
and U18582 (N_18582,N_17660,N_17812);
nor U18583 (N_18583,N_17474,N_17521);
and U18584 (N_18584,N_17952,N_17596);
and U18585 (N_18585,N_17422,N_17780);
or U18586 (N_18586,N_17402,N_17930);
nor U18587 (N_18587,N_17886,N_17904);
nand U18588 (N_18588,N_17788,N_17877);
and U18589 (N_18589,N_17954,N_17420);
xor U18590 (N_18590,N_17690,N_17925);
xor U18591 (N_18591,N_17568,N_17618);
nand U18592 (N_18592,N_17620,N_17677);
xor U18593 (N_18593,N_17451,N_17564);
or U18594 (N_18594,N_17550,N_17466);
and U18595 (N_18595,N_17946,N_17747);
nor U18596 (N_18596,N_17525,N_17868);
xnor U18597 (N_18597,N_17427,N_17609);
and U18598 (N_18598,N_17889,N_17418);
nor U18599 (N_18599,N_17568,N_17525);
and U18600 (N_18600,N_18038,N_18167);
xnor U18601 (N_18601,N_18111,N_18466);
and U18602 (N_18602,N_18109,N_18454);
nand U18603 (N_18603,N_18489,N_18455);
and U18604 (N_18604,N_18361,N_18305);
xnor U18605 (N_18605,N_18160,N_18042);
xor U18606 (N_18606,N_18108,N_18062);
and U18607 (N_18607,N_18512,N_18275);
xor U18608 (N_18608,N_18555,N_18403);
and U18609 (N_18609,N_18030,N_18198);
and U18610 (N_18610,N_18434,N_18479);
or U18611 (N_18611,N_18126,N_18084);
and U18612 (N_18612,N_18015,N_18067);
nor U18613 (N_18613,N_18319,N_18467);
and U18614 (N_18614,N_18289,N_18298);
nor U18615 (N_18615,N_18297,N_18285);
xor U18616 (N_18616,N_18511,N_18087);
xor U18617 (N_18617,N_18313,N_18472);
and U18618 (N_18618,N_18185,N_18291);
nor U18619 (N_18619,N_18175,N_18418);
nand U18620 (N_18620,N_18351,N_18035);
or U18621 (N_18621,N_18099,N_18047);
nand U18622 (N_18622,N_18274,N_18179);
nand U18623 (N_18623,N_18590,N_18352);
and U18624 (N_18624,N_18417,N_18329);
or U18625 (N_18625,N_18181,N_18071);
nand U18626 (N_18626,N_18483,N_18131);
nor U18627 (N_18627,N_18095,N_18471);
or U18628 (N_18628,N_18114,N_18475);
nand U18629 (N_18629,N_18252,N_18345);
and U18630 (N_18630,N_18120,N_18251);
nor U18631 (N_18631,N_18436,N_18036);
nand U18632 (N_18632,N_18468,N_18037);
and U18633 (N_18633,N_18428,N_18133);
or U18634 (N_18634,N_18562,N_18155);
and U18635 (N_18635,N_18498,N_18056);
nor U18636 (N_18636,N_18446,N_18094);
nor U18637 (N_18637,N_18384,N_18368);
nor U18638 (N_18638,N_18458,N_18584);
and U18639 (N_18639,N_18057,N_18162);
or U18640 (N_18640,N_18150,N_18494);
or U18641 (N_18641,N_18465,N_18052);
nor U18642 (N_18642,N_18541,N_18365);
or U18643 (N_18643,N_18140,N_18106);
nand U18644 (N_18644,N_18112,N_18441);
xor U18645 (N_18645,N_18238,N_18380);
nor U18646 (N_18646,N_18110,N_18320);
xnor U18647 (N_18647,N_18374,N_18533);
nor U18648 (N_18648,N_18206,N_18089);
nor U18649 (N_18649,N_18598,N_18060);
and U18650 (N_18650,N_18528,N_18088);
and U18651 (N_18651,N_18457,N_18557);
nor U18652 (N_18652,N_18515,N_18437);
nand U18653 (N_18653,N_18388,N_18199);
nand U18654 (N_18654,N_18576,N_18523);
nand U18655 (N_18655,N_18294,N_18383);
nor U18656 (N_18656,N_18544,N_18283);
nand U18657 (N_18657,N_18478,N_18407);
nor U18658 (N_18658,N_18264,N_18027);
and U18659 (N_18659,N_18082,N_18325);
or U18660 (N_18660,N_18213,N_18443);
and U18661 (N_18661,N_18081,N_18210);
nor U18662 (N_18662,N_18113,N_18396);
and U18663 (N_18663,N_18451,N_18002);
nand U18664 (N_18664,N_18547,N_18444);
and U18665 (N_18665,N_18172,N_18221);
xnor U18666 (N_18666,N_18408,N_18116);
or U18667 (N_18667,N_18265,N_18149);
xor U18668 (N_18668,N_18393,N_18013);
nor U18669 (N_18669,N_18018,N_18334);
xnor U18670 (N_18670,N_18044,N_18554);
xor U18671 (N_18671,N_18369,N_18163);
xor U18672 (N_18672,N_18281,N_18500);
xor U18673 (N_18673,N_18164,N_18566);
xnor U18674 (N_18674,N_18061,N_18245);
nand U18675 (N_18675,N_18226,N_18053);
nand U18676 (N_18676,N_18491,N_18177);
or U18677 (N_18677,N_18460,N_18415);
xnor U18678 (N_18678,N_18039,N_18214);
and U18679 (N_18679,N_18440,N_18370);
nand U18680 (N_18680,N_18241,N_18447);
nor U18681 (N_18681,N_18239,N_18518);
xor U18682 (N_18682,N_18247,N_18234);
nor U18683 (N_18683,N_18371,N_18197);
or U18684 (N_18684,N_18091,N_18019);
nand U18685 (N_18685,N_18017,N_18299);
or U18686 (N_18686,N_18190,N_18008);
nor U18687 (N_18687,N_18398,N_18492);
xnor U18688 (N_18688,N_18272,N_18355);
nor U18689 (N_18689,N_18308,N_18470);
xor U18690 (N_18690,N_18542,N_18293);
and U18691 (N_18691,N_18514,N_18553);
nand U18692 (N_18692,N_18020,N_18287);
nand U18693 (N_18693,N_18144,N_18263);
nor U18694 (N_18694,N_18461,N_18064);
or U18695 (N_18695,N_18323,N_18105);
xor U18696 (N_18696,N_18310,N_18201);
and U18697 (N_18697,N_18259,N_18349);
and U18698 (N_18698,N_18385,N_18069);
nor U18699 (N_18699,N_18159,N_18121);
and U18700 (N_18700,N_18335,N_18525);
nor U18701 (N_18701,N_18208,N_18249);
nor U18702 (N_18702,N_18326,N_18078);
nand U18703 (N_18703,N_18490,N_18519);
nor U18704 (N_18704,N_18191,N_18207);
or U18705 (N_18705,N_18059,N_18180);
nand U18706 (N_18706,N_18068,N_18049);
nor U18707 (N_18707,N_18040,N_18532);
xor U18708 (N_18708,N_18558,N_18550);
nand U18709 (N_18709,N_18507,N_18065);
xor U18710 (N_18710,N_18058,N_18166);
or U18711 (N_18711,N_18154,N_18250);
nand U18712 (N_18712,N_18083,N_18495);
and U18713 (N_18713,N_18477,N_18248);
or U18714 (N_18714,N_18389,N_18364);
or U18715 (N_18715,N_18222,N_18531);
or U18716 (N_18716,N_18410,N_18539);
and U18717 (N_18717,N_18151,N_18333);
nand U18718 (N_18718,N_18381,N_18025);
or U18719 (N_18719,N_18186,N_18304);
and U18720 (N_18720,N_18306,N_18168);
nor U18721 (N_18721,N_18445,N_18529);
and U18722 (N_18722,N_18493,N_18192);
xnor U18723 (N_18723,N_18358,N_18314);
and U18724 (N_18724,N_18288,N_18256);
nand U18725 (N_18725,N_18107,N_18045);
or U18726 (N_18726,N_18406,N_18536);
and U18727 (N_18727,N_18378,N_18397);
nand U18728 (N_18728,N_18543,N_18170);
xnor U18729 (N_18729,N_18327,N_18508);
and U18730 (N_18730,N_18004,N_18255);
xnor U18731 (N_18731,N_18591,N_18130);
or U18732 (N_18732,N_18473,N_18503);
or U18733 (N_18733,N_18506,N_18073);
nand U18734 (N_18734,N_18307,N_18100);
and U18735 (N_18735,N_18409,N_18520);
or U18736 (N_18736,N_18581,N_18548);
nand U18737 (N_18737,N_18429,N_18379);
nor U18738 (N_18738,N_18152,N_18330);
or U18739 (N_18739,N_18311,N_18141);
xnor U18740 (N_18740,N_18286,N_18537);
or U18741 (N_18741,N_18161,N_18411);
nand U18742 (N_18742,N_18359,N_18404);
and U18743 (N_18743,N_18273,N_18387);
or U18744 (N_18744,N_18243,N_18070);
and U18745 (N_18745,N_18597,N_18146);
xnor U18746 (N_18746,N_18295,N_18278);
nor U18747 (N_18747,N_18505,N_18413);
nor U18748 (N_18748,N_18101,N_18416);
and U18749 (N_18749,N_18344,N_18093);
and U18750 (N_18750,N_18549,N_18143);
and U18751 (N_18751,N_18439,N_18572);
or U18752 (N_18752,N_18309,N_18228);
xnor U18753 (N_18753,N_18302,N_18183);
xnor U18754 (N_18754,N_18196,N_18592);
nand U18755 (N_18755,N_18347,N_18033);
nand U18756 (N_18756,N_18136,N_18217);
or U18757 (N_18757,N_18579,N_18240);
nand U18758 (N_18758,N_18024,N_18211);
xor U18759 (N_18759,N_18484,N_18125);
and U18760 (N_18760,N_18194,N_18098);
or U18761 (N_18761,N_18414,N_18300);
or U18762 (N_18762,N_18405,N_18524);
nor U18763 (N_18763,N_18235,N_18189);
and U18764 (N_18764,N_18269,N_18337);
nand U18765 (N_18765,N_18595,N_18096);
xor U18766 (N_18766,N_18354,N_18236);
and U18767 (N_18767,N_18401,N_18296);
nand U18768 (N_18768,N_18317,N_18203);
and U18769 (N_18769,N_18209,N_18080);
and U18770 (N_18770,N_18315,N_18043);
or U18771 (N_18771,N_18254,N_18474);
or U18772 (N_18772,N_18032,N_18242);
xnor U18773 (N_18773,N_18123,N_18048);
and U18774 (N_18774,N_18261,N_18423);
and U18775 (N_18775,N_18450,N_18482);
xnor U18776 (N_18776,N_18430,N_18582);
nand U18777 (N_18777,N_18338,N_18090);
or U18778 (N_18778,N_18270,N_18501);
nor U18779 (N_18779,N_18362,N_18224);
nand U18780 (N_18780,N_18054,N_18076);
nand U18781 (N_18781,N_18118,N_18268);
or U18782 (N_18782,N_18014,N_18594);
nor U18783 (N_18783,N_18257,N_18431);
nor U18784 (N_18784,N_18200,N_18426);
nand U18785 (N_18785,N_18573,N_18469);
xnor U18786 (N_18786,N_18276,N_18427);
and U18787 (N_18787,N_18284,N_18570);
nand U18788 (N_18788,N_18092,N_18034);
nand U18789 (N_18789,N_18481,N_18559);
and U18790 (N_18790,N_18321,N_18022);
or U18791 (N_18791,N_18530,N_18202);
nand U18792 (N_18792,N_18322,N_18564);
xnor U18793 (N_18793,N_18367,N_18223);
or U18794 (N_18794,N_18551,N_18567);
nand U18795 (N_18795,N_18459,N_18363);
and U18796 (N_18796,N_18229,N_18328);
or U18797 (N_18797,N_18391,N_18051);
and U18798 (N_18798,N_18173,N_18497);
xnor U18799 (N_18799,N_18342,N_18124);
nand U18800 (N_18800,N_18253,N_18425);
xnor U18801 (N_18801,N_18122,N_18117);
or U18802 (N_18802,N_18055,N_18174);
and U18803 (N_18803,N_18341,N_18119);
and U18804 (N_18804,N_18586,N_18205);
nor U18805 (N_18805,N_18165,N_18237);
or U18806 (N_18806,N_18260,N_18233);
xnor U18807 (N_18807,N_18142,N_18016);
nor U18808 (N_18808,N_18448,N_18386);
xor U18809 (N_18809,N_18292,N_18563);
nor U18810 (N_18810,N_18282,N_18066);
nor U18811 (N_18811,N_18599,N_18516);
or U18812 (N_18812,N_18003,N_18504);
and U18813 (N_18813,N_18026,N_18277);
and U18814 (N_18814,N_18462,N_18464);
or U18815 (N_18815,N_18000,N_18097);
nand U18816 (N_18816,N_18128,N_18452);
nand U18817 (N_18817,N_18134,N_18225);
or U18818 (N_18818,N_18339,N_18230);
nand U18819 (N_18819,N_18546,N_18332);
xnor U18820 (N_18820,N_18578,N_18050);
xor U18821 (N_18821,N_18375,N_18279);
nand U18822 (N_18822,N_18395,N_18510);
and U18823 (N_18823,N_18178,N_18453);
or U18824 (N_18824,N_18589,N_18587);
xnor U18825 (N_18825,N_18266,N_18145);
and U18826 (N_18826,N_18422,N_18438);
xor U18827 (N_18827,N_18583,N_18139);
nor U18828 (N_18828,N_18487,N_18509);
or U18829 (N_18829,N_18392,N_18433);
nand U18830 (N_18830,N_18571,N_18496);
xnor U18831 (N_18831,N_18535,N_18227);
and U18832 (N_18832,N_18373,N_18331);
nor U18833 (N_18833,N_18577,N_18522);
nor U18834 (N_18834,N_18499,N_18588);
and U18835 (N_18835,N_18156,N_18449);
xor U18836 (N_18836,N_18005,N_18568);
and U18837 (N_18837,N_18021,N_18394);
nand U18838 (N_18838,N_18424,N_18115);
xnor U18839 (N_18839,N_18382,N_18480);
and U18840 (N_18840,N_18343,N_18246);
nand U18841 (N_18841,N_18290,N_18193);
nand U18842 (N_18842,N_18010,N_18012);
and U18843 (N_18843,N_18102,N_18486);
and U18844 (N_18844,N_18357,N_18527);
and U18845 (N_18845,N_18340,N_18360);
and U18846 (N_18846,N_18412,N_18075);
or U18847 (N_18847,N_18176,N_18138);
nand U18848 (N_18848,N_18561,N_18007);
and U18849 (N_18849,N_18215,N_18435);
xor U18850 (N_18850,N_18526,N_18216);
and U18851 (N_18851,N_18324,N_18153);
or U18852 (N_18852,N_18127,N_18596);
or U18853 (N_18853,N_18171,N_18104);
xnor U18854 (N_18854,N_18219,N_18377);
nand U18855 (N_18855,N_18376,N_18442);
or U18856 (N_18856,N_18301,N_18353);
and U18857 (N_18857,N_18318,N_18077);
nor U18858 (N_18858,N_18148,N_18187);
nand U18859 (N_18859,N_18346,N_18420);
nand U18860 (N_18860,N_18534,N_18072);
xor U18861 (N_18861,N_18169,N_18218);
nand U18862 (N_18862,N_18560,N_18063);
and U18863 (N_18863,N_18031,N_18262);
and U18864 (N_18864,N_18366,N_18220);
nor U18865 (N_18865,N_18132,N_18147);
nand U18866 (N_18866,N_18580,N_18188);
and U18867 (N_18867,N_18488,N_18485);
nor U18868 (N_18868,N_18129,N_18258);
and U18869 (N_18869,N_18552,N_18244);
nor U18870 (N_18870,N_18103,N_18517);
xor U18871 (N_18871,N_18271,N_18402);
nand U18872 (N_18872,N_18585,N_18348);
nand U18873 (N_18873,N_18350,N_18046);
xor U18874 (N_18874,N_18421,N_18267);
or U18875 (N_18875,N_18540,N_18432);
xor U18876 (N_18876,N_18009,N_18023);
and U18877 (N_18877,N_18336,N_18545);
or U18878 (N_18878,N_18157,N_18006);
nand U18879 (N_18879,N_18204,N_18312);
nand U18880 (N_18880,N_18028,N_18593);
or U18881 (N_18881,N_18399,N_18574);
nor U18882 (N_18882,N_18372,N_18195);
xor U18883 (N_18883,N_18041,N_18390);
nand U18884 (N_18884,N_18231,N_18556);
and U18885 (N_18885,N_18316,N_18513);
and U18886 (N_18886,N_18521,N_18182);
and U18887 (N_18887,N_18456,N_18280);
nor U18888 (N_18888,N_18400,N_18011);
or U18889 (N_18889,N_18419,N_18074);
or U18890 (N_18890,N_18001,N_18086);
nor U18891 (N_18891,N_18232,N_18079);
or U18892 (N_18892,N_18303,N_18569);
and U18893 (N_18893,N_18356,N_18029);
and U18894 (N_18894,N_18565,N_18184);
xnor U18895 (N_18895,N_18502,N_18212);
nor U18896 (N_18896,N_18137,N_18538);
and U18897 (N_18897,N_18158,N_18135);
nand U18898 (N_18898,N_18463,N_18085);
and U18899 (N_18899,N_18575,N_18476);
nor U18900 (N_18900,N_18597,N_18068);
nand U18901 (N_18901,N_18590,N_18103);
xor U18902 (N_18902,N_18357,N_18035);
nand U18903 (N_18903,N_18258,N_18325);
and U18904 (N_18904,N_18110,N_18325);
or U18905 (N_18905,N_18405,N_18217);
and U18906 (N_18906,N_18505,N_18308);
or U18907 (N_18907,N_18177,N_18557);
nand U18908 (N_18908,N_18250,N_18276);
nor U18909 (N_18909,N_18115,N_18450);
nand U18910 (N_18910,N_18244,N_18555);
xor U18911 (N_18911,N_18493,N_18149);
or U18912 (N_18912,N_18092,N_18161);
nor U18913 (N_18913,N_18521,N_18456);
xnor U18914 (N_18914,N_18571,N_18547);
xnor U18915 (N_18915,N_18248,N_18259);
nor U18916 (N_18916,N_18442,N_18382);
nor U18917 (N_18917,N_18333,N_18205);
xnor U18918 (N_18918,N_18438,N_18299);
xnor U18919 (N_18919,N_18549,N_18377);
nor U18920 (N_18920,N_18505,N_18091);
or U18921 (N_18921,N_18113,N_18262);
nand U18922 (N_18922,N_18267,N_18439);
nand U18923 (N_18923,N_18201,N_18087);
and U18924 (N_18924,N_18463,N_18280);
nand U18925 (N_18925,N_18278,N_18270);
nor U18926 (N_18926,N_18251,N_18432);
and U18927 (N_18927,N_18037,N_18320);
or U18928 (N_18928,N_18259,N_18251);
nand U18929 (N_18929,N_18104,N_18475);
xnor U18930 (N_18930,N_18388,N_18583);
nor U18931 (N_18931,N_18472,N_18103);
nor U18932 (N_18932,N_18175,N_18389);
nor U18933 (N_18933,N_18362,N_18092);
or U18934 (N_18934,N_18150,N_18466);
or U18935 (N_18935,N_18490,N_18271);
xnor U18936 (N_18936,N_18484,N_18395);
nand U18937 (N_18937,N_18550,N_18402);
xor U18938 (N_18938,N_18336,N_18547);
and U18939 (N_18939,N_18424,N_18005);
nand U18940 (N_18940,N_18558,N_18091);
and U18941 (N_18941,N_18409,N_18003);
nor U18942 (N_18942,N_18058,N_18024);
xor U18943 (N_18943,N_18225,N_18580);
or U18944 (N_18944,N_18372,N_18240);
nand U18945 (N_18945,N_18076,N_18239);
nor U18946 (N_18946,N_18284,N_18062);
and U18947 (N_18947,N_18487,N_18016);
or U18948 (N_18948,N_18448,N_18576);
xnor U18949 (N_18949,N_18060,N_18024);
nand U18950 (N_18950,N_18482,N_18262);
nand U18951 (N_18951,N_18542,N_18333);
nor U18952 (N_18952,N_18503,N_18463);
nor U18953 (N_18953,N_18034,N_18575);
nand U18954 (N_18954,N_18450,N_18439);
or U18955 (N_18955,N_18593,N_18013);
nor U18956 (N_18956,N_18431,N_18392);
and U18957 (N_18957,N_18456,N_18007);
nor U18958 (N_18958,N_18025,N_18090);
nor U18959 (N_18959,N_18593,N_18245);
nor U18960 (N_18960,N_18555,N_18289);
nand U18961 (N_18961,N_18015,N_18325);
nor U18962 (N_18962,N_18071,N_18019);
or U18963 (N_18963,N_18106,N_18574);
or U18964 (N_18964,N_18326,N_18131);
nor U18965 (N_18965,N_18011,N_18086);
and U18966 (N_18966,N_18211,N_18443);
and U18967 (N_18967,N_18288,N_18549);
and U18968 (N_18968,N_18274,N_18400);
nand U18969 (N_18969,N_18211,N_18130);
and U18970 (N_18970,N_18355,N_18025);
and U18971 (N_18971,N_18142,N_18405);
xnor U18972 (N_18972,N_18338,N_18200);
xnor U18973 (N_18973,N_18375,N_18042);
xor U18974 (N_18974,N_18520,N_18029);
nand U18975 (N_18975,N_18002,N_18368);
nor U18976 (N_18976,N_18290,N_18172);
nor U18977 (N_18977,N_18335,N_18480);
or U18978 (N_18978,N_18415,N_18428);
xor U18979 (N_18979,N_18008,N_18059);
nand U18980 (N_18980,N_18446,N_18079);
nand U18981 (N_18981,N_18059,N_18134);
or U18982 (N_18982,N_18393,N_18353);
and U18983 (N_18983,N_18066,N_18476);
nand U18984 (N_18984,N_18314,N_18289);
xnor U18985 (N_18985,N_18197,N_18007);
nor U18986 (N_18986,N_18116,N_18553);
nand U18987 (N_18987,N_18266,N_18537);
nand U18988 (N_18988,N_18156,N_18550);
and U18989 (N_18989,N_18235,N_18396);
xnor U18990 (N_18990,N_18429,N_18310);
and U18991 (N_18991,N_18086,N_18158);
xor U18992 (N_18992,N_18358,N_18091);
nor U18993 (N_18993,N_18425,N_18178);
and U18994 (N_18994,N_18445,N_18295);
nand U18995 (N_18995,N_18404,N_18182);
xnor U18996 (N_18996,N_18355,N_18400);
or U18997 (N_18997,N_18077,N_18371);
nand U18998 (N_18998,N_18461,N_18274);
or U18999 (N_18999,N_18505,N_18009);
and U19000 (N_19000,N_18220,N_18122);
nand U19001 (N_19001,N_18207,N_18363);
and U19002 (N_19002,N_18585,N_18231);
and U19003 (N_19003,N_18019,N_18334);
xnor U19004 (N_19004,N_18034,N_18192);
xnor U19005 (N_19005,N_18183,N_18448);
nand U19006 (N_19006,N_18229,N_18224);
nor U19007 (N_19007,N_18430,N_18566);
nand U19008 (N_19008,N_18539,N_18474);
or U19009 (N_19009,N_18143,N_18595);
xnor U19010 (N_19010,N_18079,N_18069);
or U19011 (N_19011,N_18027,N_18066);
nand U19012 (N_19012,N_18123,N_18370);
nor U19013 (N_19013,N_18535,N_18148);
nor U19014 (N_19014,N_18169,N_18368);
xor U19015 (N_19015,N_18564,N_18006);
xor U19016 (N_19016,N_18215,N_18317);
nand U19017 (N_19017,N_18457,N_18328);
nor U19018 (N_19018,N_18526,N_18553);
and U19019 (N_19019,N_18206,N_18080);
xor U19020 (N_19020,N_18036,N_18179);
nand U19021 (N_19021,N_18490,N_18401);
or U19022 (N_19022,N_18007,N_18091);
or U19023 (N_19023,N_18463,N_18533);
xnor U19024 (N_19024,N_18084,N_18156);
nor U19025 (N_19025,N_18402,N_18240);
and U19026 (N_19026,N_18502,N_18106);
xnor U19027 (N_19027,N_18036,N_18028);
and U19028 (N_19028,N_18316,N_18238);
nor U19029 (N_19029,N_18162,N_18105);
and U19030 (N_19030,N_18250,N_18236);
xor U19031 (N_19031,N_18399,N_18526);
or U19032 (N_19032,N_18259,N_18193);
or U19033 (N_19033,N_18154,N_18067);
nand U19034 (N_19034,N_18532,N_18365);
nand U19035 (N_19035,N_18204,N_18350);
and U19036 (N_19036,N_18250,N_18128);
xnor U19037 (N_19037,N_18399,N_18522);
and U19038 (N_19038,N_18063,N_18414);
nor U19039 (N_19039,N_18113,N_18148);
nand U19040 (N_19040,N_18269,N_18116);
nor U19041 (N_19041,N_18331,N_18070);
and U19042 (N_19042,N_18495,N_18405);
xnor U19043 (N_19043,N_18284,N_18286);
nand U19044 (N_19044,N_18336,N_18513);
nor U19045 (N_19045,N_18104,N_18300);
nor U19046 (N_19046,N_18401,N_18102);
xor U19047 (N_19047,N_18112,N_18423);
or U19048 (N_19048,N_18124,N_18594);
and U19049 (N_19049,N_18189,N_18464);
or U19050 (N_19050,N_18162,N_18581);
xor U19051 (N_19051,N_18378,N_18324);
and U19052 (N_19052,N_18537,N_18153);
nor U19053 (N_19053,N_18464,N_18598);
nand U19054 (N_19054,N_18346,N_18005);
and U19055 (N_19055,N_18530,N_18364);
nor U19056 (N_19056,N_18414,N_18570);
nor U19057 (N_19057,N_18551,N_18565);
and U19058 (N_19058,N_18593,N_18499);
nor U19059 (N_19059,N_18401,N_18224);
nor U19060 (N_19060,N_18272,N_18512);
xor U19061 (N_19061,N_18239,N_18403);
nand U19062 (N_19062,N_18425,N_18042);
and U19063 (N_19063,N_18014,N_18377);
xnor U19064 (N_19064,N_18496,N_18397);
and U19065 (N_19065,N_18453,N_18239);
xnor U19066 (N_19066,N_18167,N_18469);
or U19067 (N_19067,N_18387,N_18035);
xor U19068 (N_19068,N_18328,N_18361);
or U19069 (N_19069,N_18148,N_18200);
nor U19070 (N_19070,N_18088,N_18590);
xnor U19071 (N_19071,N_18298,N_18376);
and U19072 (N_19072,N_18268,N_18263);
nor U19073 (N_19073,N_18339,N_18027);
and U19074 (N_19074,N_18407,N_18271);
nor U19075 (N_19075,N_18454,N_18371);
xnor U19076 (N_19076,N_18042,N_18560);
nand U19077 (N_19077,N_18547,N_18032);
and U19078 (N_19078,N_18379,N_18320);
or U19079 (N_19079,N_18091,N_18186);
or U19080 (N_19080,N_18571,N_18355);
xnor U19081 (N_19081,N_18235,N_18164);
nor U19082 (N_19082,N_18316,N_18504);
or U19083 (N_19083,N_18374,N_18248);
nor U19084 (N_19084,N_18272,N_18537);
nor U19085 (N_19085,N_18550,N_18096);
or U19086 (N_19086,N_18158,N_18508);
nand U19087 (N_19087,N_18138,N_18097);
and U19088 (N_19088,N_18221,N_18176);
or U19089 (N_19089,N_18477,N_18148);
xor U19090 (N_19090,N_18228,N_18028);
and U19091 (N_19091,N_18116,N_18218);
xor U19092 (N_19092,N_18301,N_18355);
xnor U19093 (N_19093,N_18426,N_18501);
xor U19094 (N_19094,N_18301,N_18568);
or U19095 (N_19095,N_18310,N_18555);
nand U19096 (N_19096,N_18597,N_18149);
nand U19097 (N_19097,N_18096,N_18338);
or U19098 (N_19098,N_18597,N_18241);
and U19099 (N_19099,N_18228,N_18346);
or U19100 (N_19100,N_18157,N_18339);
nor U19101 (N_19101,N_18078,N_18370);
nand U19102 (N_19102,N_18303,N_18245);
or U19103 (N_19103,N_18573,N_18091);
nor U19104 (N_19104,N_18323,N_18480);
nor U19105 (N_19105,N_18128,N_18172);
nand U19106 (N_19106,N_18205,N_18274);
and U19107 (N_19107,N_18460,N_18242);
nand U19108 (N_19108,N_18173,N_18180);
nand U19109 (N_19109,N_18099,N_18471);
and U19110 (N_19110,N_18445,N_18510);
and U19111 (N_19111,N_18443,N_18205);
or U19112 (N_19112,N_18148,N_18422);
or U19113 (N_19113,N_18490,N_18354);
nor U19114 (N_19114,N_18553,N_18185);
and U19115 (N_19115,N_18322,N_18382);
nor U19116 (N_19116,N_18260,N_18513);
xor U19117 (N_19117,N_18034,N_18106);
and U19118 (N_19118,N_18062,N_18382);
xnor U19119 (N_19119,N_18376,N_18241);
or U19120 (N_19120,N_18490,N_18038);
and U19121 (N_19121,N_18531,N_18479);
nand U19122 (N_19122,N_18013,N_18586);
or U19123 (N_19123,N_18277,N_18131);
or U19124 (N_19124,N_18323,N_18369);
and U19125 (N_19125,N_18203,N_18344);
nor U19126 (N_19126,N_18508,N_18033);
and U19127 (N_19127,N_18154,N_18394);
nor U19128 (N_19128,N_18138,N_18203);
and U19129 (N_19129,N_18373,N_18254);
nand U19130 (N_19130,N_18443,N_18069);
xor U19131 (N_19131,N_18464,N_18548);
nand U19132 (N_19132,N_18426,N_18021);
and U19133 (N_19133,N_18267,N_18282);
nor U19134 (N_19134,N_18507,N_18455);
nand U19135 (N_19135,N_18235,N_18251);
xor U19136 (N_19136,N_18063,N_18131);
nor U19137 (N_19137,N_18513,N_18211);
or U19138 (N_19138,N_18315,N_18076);
nor U19139 (N_19139,N_18069,N_18463);
nand U19140 (N_19140,N_18046,N_18417);
xnor U19141 (N_19141,N_18117,N_18078);
nor U19142 (N_19142,N_18416,N_18357);
and U19143 (N_19143,N_18193,N_18262);
or U19144 (N_19144,N_18545,N_18513);
nand U19145 (N_19145,N_18259,N_18303);
nor U19146 (N_19146,N_18343,N_18424);
xnor U19147 (N_19147,N_18491,N_18031);
nor U19148 (N_19148,N_18542,N_18411);
and U19149 (N_19149,N_18338,N_18346);
and U19150 (N_19150,N_18172,N_18222);
and U19151 (N_19151,N_18492,N_18511);
or U19152 (N_19152,N_18101,N_18025);
or U19153 (N_19153,N_18151,N_18132);
nand U19154 (N_19154,N_18348,N_18008);
and U19155 (N_19155,N_18090,N_18441);
nand U19156 (N_19156,N_18552,N_18363);
xor U19157 (N_19157,N_18077,N_18146);
or U19158 (N_19158,N_18517,N_18385);
and U19159 (N_19159,N_18125,N_18111);
xnor U19160 (N_19160,N_18449,N_18211);
nand U19161 (N_19161,N_18252,N_18520);
nor U19162 (N_19162,N_18366,N_18208);
nor U19163 (N_19163,N_18501,N_18499);
xnor U19164 (N_19164,N_18538,N_18125);
xor U19165 (N_19165,N_18486,N_18403);
nand U19166 (N_19166,N_18384,N_18156);
and U19167 (N_19167,N_18251,N_18598);
nor U19168 (N_19168,N_18316,N_18334);
and U19169 (N_19169,N_18531,N_18559);
and U19170 (N_19170,N_18082,N_18438);
nand U19171 (N_19171,N_18417,N_18596);
xor U19172 (N_19172,N_18118,N_18312);
nand U19173 (N_19173,N_18089,N_18549);
and U19174 (N_19174,N_18234,N_18196);
or U19175 (N_19175,N_18054,N_18384);
xnor U19176 (N_19176,N_18436,N_18572);
and U19177 (N_19177,N_18041,N_18051);
nor U19178 (N_19178,N_18199,N_18138);
xnor U19179 (N_19179,N_18215,N_18473);
xnor U19180 (N_19180,N_18484,N_18354);
nand U19181 (N_19181,N_18247,N_18331);
nand U19182 (N_19182,N_18272,N_18500);
nand U19183 (N_19183,N_18074,N_18235);
or U19184 (N_19184,N_18557,N_18227);
or U19185 (N_19185,N_18281,N_18136);
or U19186 (N_19186,N_18278,N_18097);
and U19187 (N_19187,N_18409,N_18408);
and U19188 (N_19188,N_18437,N_18323);
nand U19189 (N_19189,N_18117,N_18223);
xnor U19190 (N_19190,N_18262,N_18170);
nor U19191 (N_19191,N_18302,N_18251);
and U19192 (N_19192,N_18244,N_18120);
xnor U19193 (N_19193,N_18423,N_18418);
and U19194 (N_19194,N_18407,N_18232);
xor U19195 (N_19195,N_18583,N_18094);
or U19196 (N_19196,N_18259,N_18014);
and U19197 (N_19197,N_18305,N_18348);
nor U19198 (N_19198,N_18499,N_18102);
or U19199 (N_19199,N_18275,N_18172);
and U19200 (N_19200,N_19168,N_18958);
and U19201 (N_19201,N_18815,N_18994);
nor U19202 (N_19202,N_18798,N_18953);
xor U19203 (N_19203,N_18904,N_18674);
nand U19204 (N_19204,N_19053,N_18842);
xor U19205 (N_19205,N_18949,N_19056);
nand U19206 (N_19206,N_18636,N_19100);
nor U19207 (N_19207,N_19070,N_19025);
and U19208 (N_19208,N_19038,N_19107);
and U19209 (N_19209,N_18708,N_18691);
nor U19210 (N_19210,N_18793,N_18903);
and U19211 (N_19211,N_18871,N_18847);
nor U19212 (N_19212,N_18955,N_18646);
and U19213 (N_19213,N_18931,N_18701);
nand U19214 (N_19214,N_19040,N_19089);
and U19215 (N_19215,N_19184,N_18688);
nand U19216 (N_19216,N_19095,N_19085);
and U19217 (N_19217,N_19193,N_18698);
nand U19218 (N_19218,N_18984,N_19088);
xor U19219 (N_19219,N_18826,N_19161);
xnor U19220 (N_19220,N_19047,N_18703);
and U19221 (N_19221,N_18620,N_18838);
nand U19222 (N_19222,N_18910,N_18684);
and U19223 (N_19223,N_18985,N_18977);
nand U19224 (N_19224,N_18754,N_19147);
or U19225 (N_19225,N_18868,N_18634);
nand U19226 (N_19226,N_18621,N_18801);
nor U19227 (N_19227,N_19041,N_18618);
and U19228 (N_19228,N_19083,N_19033);
nor U19229 (N_19229,N_19178,N_18655);
xnor U19230 (N_19230,N_18648,N_18612);
nor U19231 (N_19231,N_18813,N_18778);
nand U19232 (N_19232,N_18716,N_18865);
and U19233 (N_19233,N_18697,N_18809);
nor U19234 (N_19234,N_18600,N_18829);
xnor U19235 (N_19235,N_18998,N_18909);
or U19236 (N_19236,N_19113,N_18879);
nand U19237 (N_19237,N_18914,N_18605);
nor U19238 (N_19238,N_19014,N_19078);
nor U19239 (N_19239,N_19170,N_18745);
nor U19240 (N_19240,N_19004,N_18846);
and U19241 (N_19241,N_19103,N_18786);
or U19242 (N_19242,N_18643,N_18682);
nor U19243 (N_19243,N_19190,N_18719);
xnor U19244 (N_19244,N_19029,N_19062);
and U19245 (N_19245,N_18777,N_18905);
nand U19246 (N_19246,N_19188,N_18824);
nor U19247 (N_19247,N_18992,N_18650);
nand U19248 (N_19248,N_19013,N_18767);
xnor U19249 (N_19249,N_18653,N_19067);
nand U19250 (N_19250,N_18988,N_19198);
xor U19251 (N_19251,N_18952,N_18950);
nand U19252 (N_19252,N_19090,N_18819);
xnor U19253 (N_19253,N_18934,N_18869);
nand U19254 (N_19254,N_19151,N_18933);
xnor U19255 (N_19255,N_18746,N_19019);
nand U19256 (N_19256,N_18668,N_18916);
nor U19257 (N_19257,N_18918,N_18738);
and U19258 (N_19258,N_18792,N_18694);
nor U19259 (N_19259,N_18707,N_18687);
or U19260 (N_19260,N_19008,N_18610);
xor U19261 (N_19261,N_18844,N_19048);
xnor U19262 (N_19262,N_18639,N_19143);
nand U19263 (N_19263,N_18867,N_19139);
xor U19264 (N_19264,N_18928,N_18676);
xor U19265 (N_19265,N_19077,N_18835);
xor U19266 (N_19266,N_18751,N_18635);
nand U19267 (N_19267,N_19132,N_19102);
xnor U19268 (N_19268,N_19181,N_18893);
nand U19269 (N_19269,N_18802,N_19086);
or U19270 (N_19270,N_18656,N_19105);
and U19271 (N_19271,N_19141,N_19076);
xnor U19272 (N_19272,N_18706,N_18803);
nand U19273 (N_19273,N_18692,N_19064);
nor U19274 (N_19274,N_18756,N_18839);
and U19275 (N_19275,N_18690,N_19110);
xor U19276 (N_19276,N_19007,N_18836);
nor U19277 (N_19277,N_19060,N_19022);
and U19278 (N_19278,N_18900,N_18911);
or U19279 (N_19279,N_18947,N_18724);
or U19280 (N_19280,N_18946,N_19138);
and U19281 (N_19281,N_18741,N_18999);
xnor U19282 (N_19282,N_18915,N_18732);
xor U19283 (N_19283,N_18712,N_18885);
and U19284 (N_19284,N_19074,N_18622);
nand U19285 (N_19285,N_19012,N_18679);
and U19286 (N_19286,N_18886,N_18929);
and U19287 (N_19287,N_18660,N_18939);
nor U19288 (N_19288,N_18963,N_19032);
xnor U19289 (N_19289,N_18875,N_18616);
or U19290 (N_19290,N_18968,N_18833);
nor U19291 (N_19291,N_18628,N_19106);
xor U19292 (N_19292,N_19097,N_19093);
or U19293 (N_19293,N_19034,N_19119);
nand U19294 (N_19294,N_19058,N_19010);
nor U19295 (N_19295,N_19197,N_18727);
xor U19296 (N_19296,N_18830,N_18891);
and U19297 (N_19297,N_18919,N_18954);
nand U19298 (N_19298,N_18921,N_18810);
nand U19299 (N_19299,N_18689,N_18603);
and U19300 (N_19300,N_18657,N_19122);
xor U19301 (N_19301,N_19082,N_18742);
xnor U19302 (N_19302,N_19123,N_18852);
and U19303 (N_19303,N_19165,N_19146);
nand U19304 (N_19304,N_18884,N_19068);
nor U19305 (N_19305,N_18808,N_19015);
or U19306 (N_19306,N_19073,N_18630);
nor U19307 (N_19307,N_19155,N_19172);
or U19308 (N_19308,N_18848,N_19072);
nor U19309 (N_19309,N_19101,N_18644);
nand U19310 (N_19310,N_19098,N_18677);
nor U19311 (N_19311,N_18661,N_19133);
or U19312 (N_19312,N_19144,N_19081);
xor U19313 (N_19313,N_18617,N_18917);
nand U19314 (N_19314,N_18980,N_18669);
nand U19315 (N_19315,N_19160,N_18757);
nor U19316 (N_19316,N_18827,N_18974);
nand U19317 (N_19317,N_19071,N_18907);
xnor U19318 (N_19318,N_18753,N_18896);
nor U19319 (N_19319,N_18725,N_18787);
xor U19320 (N_19320,N_18944,N_18898);
and U19321 (N_19321,N_19057,N_18710);
xnor U19322 (N_19322,N_18744,N_19054);
or U19323 (N_19323,N_19176,N_19124);
nand U19324 (N_19324,N_18631,N_18731);
xnor U19325 (N_19325,N_18876,N_19063);
nor U19326 (N_19326,N_18748,N_19174);
xor U19327 (N_19327,N_18874,N_18723);
nand U19328 (N_19328,N_18685,N_19137);
and U19329 (N_19329,N_18990,N_18609);
xor U19330 (N_19330,N_18764,N_18695);
xor U19331 (N_19331,N_18762,N_18686);
nor U19332 (N_19332,N_18791,N_18627);
and U19333 (N_19333,N_19027,N_19135);
nor U19334 (N_19334,N_18780,N_19189);
nand U19335 (N_19335,N_19092,N_18888);
xor U19336 (N_19336,N_19125,N_19173);
nor U19337 (N_19337,N_18670,N_18986);
or U19338 (N_19338,N_19164,N_18926);
nor U19339 (N_19339,N_18770,N_19080);
xnor U19340 (N_19340,N_19052,N_18832);
xor U19341 (N_19341,N_18705,N_18795);
and U19342 (N_19342,N_19050,N_18659);
and U19343 (N_19343,N_18664,N_19163);
xor U19344 (N_19344,N_18602,N_19128);
xor U19345 (N_19345,N_19023,N_18774);
xnor U19346 (N_19346,N_18700,N_18800);
nand U19347 (N_19347,N_18925,N_18736);
and U19348 (N_19348,N_18814,N_18854);
xor U19349 (N_19349,N_19175,N_18902);
and U19350 (N_19350,N_18807,N_18632);
nor U19351 (N_19351,N_18820,N_18872);
xnor U19352 (N_19352,N_18964,N_18666);
nand U19353 (N_19353,N_19011,N_18972);
xor U19354 (N_19354,N_19145,N_18717);
nand U19355 (N_19355,N_19191,N_19169);
nor U19356 (N_19356,N_18675,N_18941);
nor U19357 (N_19357,N_18642,N_18702);
nand U19358 (N_19358,N_18709,N_18970);
and U19359 (N_19359,N_18995,N_18781);
xor U19360 (N_19360,N_18680,N_19131);
nor U19361 (N_19361,N_19003,N_18704);
and U19362 (N_19362,N_18878,N_18796);
nand U19363 (N_19363,N_18913,N_18726);
and U19364 (N_19364,N_18765,N_19179);
nand U19365 (N_19365,N_18611,N_19028);
nor U19366 (N_19366,N_18667,N_19127);
xor U19367 (N_19367,N_19115,N_18763);
xor U19368 (N_19368,N_18658,N_18637);
xnor U19369 (N_19369,N_18960,N_18883);
nand U19370 (N_19370,N_18651,N_19009);
nand U19371 (N_19371,N_18606,N_18663);
nor U19372 (N_19372,N_19142,N_19186);
nand U19373 (N_19373,N_18788,N_19157);
xnor U19374 (N_19374,N_18654,N_18923);
nand U19375 (N_19375,N_18969,N_19150);
or U19376 (N_19376,N_18811,N_18773);
and U19377 (N_19377,N_18671,N_18943);
and U19378 (N_19378,N_18750,N_18897);
or U19379 (N_19379,N_19199,N_18713);
and U19380 (N_19380,N_19035,N_18845);
or U19381 (N_19381,N_18942,N_18831);
xor U19382 (N_19382,N_19042,N_18849);
nor U19383 (N_19383,N_19031,N_19044);
or U19384 (N_19384,N_18956,N_18640);
xnor U19385 (N_19385,N_18747,N_18912);
nor U19386 (N_19386,N_19177,N_19171);
xor U19387 (N_19387,N_18873,N_19112);
xor U19388 (N_19388,N_18681,N_19020);
or U19389 (N_19389,N_19002,N_18937);
or U19390 (N_19390,N_18860,N_19126);
or U19391 (N_19391,N_19153,N_18743);
nand U19392 (N_19392,N_18957,N_18997);
nor U19393 (N_19393,N_18805,N_18850);
nor U19394 (N_19394,N_19005,N_18840);
nand U19395 (N_19395,N_18967,N_18901);
nand U19396 (N_19396,N_18823,N_18720);
nor U19397 (N_19397,N_19167,N_19030);
nor U19398 (N_19398,N_18734,N_18728);
or U19399 (N_19399,N_18673,N_18733);
nand U19400 (N_19400,N_19194,N_19111);
and U19401 (N_19401,N_19182,N_18932);
nor U19402 (N_19402,N_19136,N_18714);
xnor U19403 (N_19403,N_19116,N_18766);
or U19404 (N_19404,N_18938,N_18894);
xor U19405 (N_19405,N_18861,N_19069);
and U19406 (N_19406,N_18951,N_18899);
nand U19407 (N_19407,N_18785,N_18715);
xnor U19408 (N_19408,N_19051,N_19017);
or U19409 (N_19409,N_18794,N_18740);
nor U19410 (N_19410,N_18821,N_18906);
nor U19411 (N_19411,N_18856,N_18601);
nand U19412 (N_19412,N_18863,N_18779);
nand U19413 (N_19413,N_19140,N_18834);
or U19414 (N_19414,N_18859,N_18625);
xor U19415 (N_19415,N_18979,N_19024);
nand U19416 (N_19416,N_18790,N_18645);
and U19417 (N_19417,N_18678,N_19187);
or U19418 (N_19418,N_19183,N_18619);
or U19419 (N_19419,N_19043,N_18649);
and U19420 (N_19420,N_18908,N_18890);
nand U19421 (N_19421,N_18935,N_19156);
nor U19422 (N_19422,N_18604,N_18959);
and U19423 (N_19423,N_18799,N_18783);
or U19424 (N_19424,N_19001,N_18940);
xor U19425 (N_19425,N_19185,N_18749);
nand U19426 (N_19426,N_19099,N_19049);
xnor U19427 (N_19427,N_18936,N_19018);
nand U19428 (N_19428,N_19006,N_19159);
nor U19429 (N_19429,N_18978,N_19079);
or U19430 (N_19430,N_18945,N_18623);
nand U19431 (N_19431,N_19192,N_18927);
or U19432 (N_19432,N_18755,N_19026);
or U19433 (N_19433,N_18665,N_18760);
and U19434 (N_19434,N_18624,N_18672);
or U19435 (N_19435,N_18613,N_19094);
nor U19436 (N_19436,N_19055,N_19075);
nand U19437 (N_19437,N_19091,N_18930);
nand U19438 (N_19438,N_18696,N_18920);
or U19439 (N_19439,N_19154,N_19120);
or U19440 (N_19440,N_18818,N_18759);
nand U19441 (N_19441,N_18855,N_18895);
nand U19442 (N_19442,N_18718,N_19158);
and U19443 (N_19443,N_18966,N_18889);
nand U19444 (N_19444,N_18825,N_18922);
nand U19445 (N_19445,N_18973,N_18693);
and U19446 (N_19446,N_19045,N_18758);
nor U19447 (N_19447,N_19196,N_18647);
nand U19448 (N_19448,N_18699,N_18769);
and U19449 (N_19449,N_18993,N_19108);
xor U19450 (N_19450,N_18841,N_18948);
or U19451 (N_19451,N_18987,N_19021);
xor U19452 (N_19452,N_18761,N_19118);
or U19453 (N_19453,N_18828,N_18626);
nand U19454 (N_19454,N_18683,N_18768);
nand U19455 (N_19455,N_18638,N_18996);
and U19456 (N_19456,N_19117,N_18789);
or U19457 (N_19457,N_18982,N_19148);
nand U19458 (N_19458,N_18782,N_18662);
and U19459 (N_19459,N_18607,N_18729);
nor U19460 (N_19460,N_18641,N_19180);
nand U19461 (N_19461,N_18721,N_18843);
and U19462 (N_19462,N_18837,N_19166);
xnor U19463 (N_19463,N_18981,N_18615);
nor U19464 (N_19464,N_18971,N_19036);
and U19465 (N_19465,N_18784,N_18614);
and U19466 (N_19466,N_18887,N_18817);
or U19467 (N_19467,N_18739,N_18629);
or U19468 (N_19468,N_18816,N_18880);
and U19469 (N_19469,N_19195,N_18608);
nand U19470 (N_19470,N_18851,N_19046);
xnor U19471 (N_19471,N_18882,N_18771);
xor U19472 (N_19472,N_18752,N_18711);
nor U19473 (N_19473,N_18806,N_18822);
nand U19474 (N_19474,N_18877,N_18735);
and U19475 (N_19475,N_19087,N_19059);
or U19476 (N_19476,N_18730,N_18812);
or U19477 (N_19477,N_18737,N_18975);
or U19478 (N_19478,N_18989,N_19065);
nor U19479 (N_19479,N_18962,N_18857);
xor U19480 (N_19480,N_19149,N_18776);
and U19481 (N_19481,N_18961,N_19039);
nor U19482 (N_19482,N_18864,N_18633);
nand U19483 (N_19483,N_18870,N_18983);
xor U19484 (N_19484,N_19000,N_19129);
and U19485 (N_19485,N_18772,N_18991);
and U19486 (N_19486,N_18976,N_19114);
or U19487 (N_19487,N_18775,N_18797);
nor U19488 (N_19488,N_18862,N_19134);
xnor U19489 (N_19489,N_18652,N_19096);
nand U19490 (N_19490,N_19084,N_18924);
xnor U19491 (N_19491,N_19016,N_19037);
and U19492 (N_19492,N_18866,N_19061);
or U19493 (N_19493,N_18722,N_19109);
nor U19494 (N_19494,N_19130,N_19152);
or U19495 (N_19495,N_19066,N_18892);
xnor U19496 (N_19496,N_18881,N_18858);
and U19497 (N_19497,N_19121,N_18804);
xor U19498 (N_19498,N_18965,N_18853);
or U19499 (N_19499,N_19104,N_19162);
nand U19500 (N_19500,N_18875,N_19054);
nand U19501 (N_19501,N_18840,N_19037);
or U19502 (N_19502,N_19014,N_19004);
nand U19503 (N_19503,N_18667,N_19195);
nand U19504 (N_19504,N_18634,N_18968);
or U19505 (N_19505,N_19013,N_18857);
nand U19506 (N_19506,N_18725,N_19144);
xnor U19507 (N_19507,N_19008,N_19088);
or U19508 (N_19508,N_19002,N_19154);
and U19509 (N_19509,N_18851,N_18918);
nor U19510 (N_19510,N_18641,N_18637);
xor U19511 (N_19511,N_19007,N_18624);
and U19512 (N_19512,N_18934,N_18685);
nand U19513 (N_19513,N_18738,N_18912);
or U19514 (N_19514,N_18997,N_18755);
xor U19515 (N_19515,N_19086,N_19041);
or U19516 (N_19516,N_19016,N_19115);
and U19517 (N_19517,N_18638,N_18802);
nand U19518 (N_19518,N_18758,N_18788);
nand U19519 (N_19519,N_18938,N_18812);
nor U19520 (N_19520,N_19064,N_19129);
and U19521 (N_19521,N_18619,N_19065);
nor U19522 (N_19522,N_18993,N_18904);
xnor U19523 (N_19523,N_18861,N_19127);
and U19524 (N_19524,N_18805,N_18678);
or U19525 (N_19525,N_18938,N_18993);
and U19526 (N_19526,N_19191,N_18710);
nand U19527 (N_19527,N_19159,N_18839);
nor U19528 (N_19528,N_18923,N_19032);
xnor U19529 (N_19529,N_18960,N_18705);
nor U19530 (N_19530,N_18944,N_18706);
or U19531 (N_19531,N_18635,N_19154);
nand U19532 (N_19532,N_19023,N_18927);
and U19533 (N_19533,N_19144,N_18622);
xor U19534 (N_19534,N_18948,N_18686);
xnor U19535 (N_19535,N_18942,N_18873);
or U19536 (N_19536,N_19124,N_18883);
or U19537 (N_19537,N_19137,N_18777);
nor U19538 (N_19538,N_18992,N_19137);
nand U19539 (N_19539,N_19135,N_19031);
or U19540 (N_19540,N_18742,N_19120);
xor U19541 (N_19541,N_18950,N_19141);
nor U19542 (N_19542,N_18943,N_18659);
and U19543 (N_19543,N_19166,N_19109);
xor U19544 (N_19544,N_19047,N_18890);
xor U19545 (N_19545,N_19024,N_18654);
nand U19546 (N_19546,N_18755,N_19004);
or U19547 (N_19547,N_18976,N_19182);
or U19548 (N_19548,N_18613,N_18936);
nand U19549 (N_19549,N_18790,N_18857);
nor U19550 (N_19550,N_19039,N_18955);
nand U19551 (N_19551,N_18870,N_18722);
or U19552 (N_19552,N_18772,N_19168);
nor U19553 (N_19553,N_18881,N_18844);
and U19554 (N_19554,N_18962,N_19007);
or U19555 (N_19555,N_18919,N_18697);
or U19556 (N_19556,N_18961,N_18824);
and U19557 (N_19557,N_19153,N_18668);
and U19558 (N_19558,N_18773,N_18830);
nand U19559 (N_19559,N_18845,N_19028);
nor U19560 (N_19560,N_18724,N_18701);
nand U19561 (N_19561,N_18809,N_18953);
and U19562 (N_19562,N_18798,N_18721);
nor U19563 (N_19563,N_19097,N_19010);
nand U19564 (N_19564,N_18809,N_18695);
and U19565 (N_19565,N_19130,N_18726);
and U19566 (N_19566,N_18820,N_18844);
xnor U19567 (N_19567,N_18703,N_19012);
nor U19568 (N_19568,N_18650,N_18621);
and U19569 (N_19569,N_18608,N_18708);
or U19570 (N_19570,N_18918,N_19104);
nand U19571 (N_19571,N_18828,N_18850);
xor U19572 (N_19572,N_19045,N_18877);
nor U19573 (N_19573,N_18731,N_18670);
and U19574 (N_19574,N_18805,N_18875);
or U19575 (N_19575,N_18748,N_18673);
nor U19576 (N_19576,N_18904,N_18621);
xnor U19577 (N_19577,N_19086,N_18690);
nor U19578 (N_19578,N_19170,N_19179);
xor U19579 (N_19579,N_19167,N_18994);
xnor U19580 (N_19580,N_18606,N_18870);
or U19581 (N_19581,N_18840,N_18784);
nand U19582 (N_19582,N_18894,N_19071);
or U19583 (N_19583,N_18815,N_18955);
nand U19584 (N_19584,N_19174,N_19189);
xnor U19585 (N_19585,N_19190,N_18631);
nand U19586 (N_19586,N_18715,N_19187);
nor U19587 (N_19587,N_19087,N_18835);
nor U19588 (N_19588,N_19047,N_18902);
or U19589 (N_19589,N_18822,N_19038);
nor U19590 (N_19590,N_18715,N_19107);
xor U19591 (N_19591,N_19084,N_19160);
nor U19592 (N_19592,N_18764,N_18927);
or U19593 (N_19593,N_19150,N_19159);
and U19594 (N_19594,N_18829,N_18876);
xnor U19595 (N_19595,N_18747,N_18669);
and U19596 (N_19596,N_18776,N_18715);
and U19597 (N_19597,N_18877,N_18638);
nor U19598 (N_19598,N_18832,N_18779);
and U19599 (N_19599,N_18735,N_18994);
xnor U19600 (N_19600,N_18813,N_18851);
and U19601 (N_19601,N_19117,N_18979);
nand U19602 (N_19602,N_18974,N_18775);
xor U19603 (N_19603,N_18830,N_18980);
and U19604 (N_19604,N_18864,N_19113);
and U19605 (N_19605,N_18915,N_19036);
xnor U19606 (N_19606,N_19048,N_18714);
and U19607 (N_19607,N_18746,N_18970);
nor U19608 (N_19608,N_18952,N_19101);
nand U19609 (N_19609,N_18674,N_19115);
xor U19610 (N_19610,N_18691,N_18812);
and U19611 (N_19611,N_18879,N_19115);
xor U19612 (N_19612,N_19101,N_19152);
nor U19613 (N_19613,N_18796,N_18797);
or U19614 (N_19614,N_19066,N_18748);
nor U19615 (N_19615,N_19150,N_18660);
and U19616 (N_19616,N_19165,N_19057);
xnor U19617 (N_19617,N_18997,N_18808);
nor U19618 (N_19618,N_19156,N_18934);
nor U19619 (N_19619,N_18948,N_18949);
nand U19620 (N_19620,N_18643,N_18822);
or U19621 (N_19621,N_18666,N_18706);
xnor U19622 (N_19622,N_19165,N_18918);
or U19623 (N_19623,N_19176,N_19173);
xor U19624 (N_19624,N_19097,N_18762);
and U19625 (N_19625,N_19094,N_19006);
or U19626 (N_19626,N_18786,N_19108);
nor U19627 (N_19627,N_19199,N_18752);
or U19628 (N_19628,N_18719,N_18856);
or U19629 (N_19629,N_18616,N_19059);
xor U19630 (N_19630,N_18632,N_18951);
nand U19631 (N_19631,N_18691,N_18728);
and U19632 (N_19632,N_19099,N_18791);
nor U19633 (N_19633,N_18701,N_19111);
and U19634 (N_19634,N_19035,N_18749);
nand U19635 (N_19635,N_19090,N_19165);
or U19636 (N_19636,N_18852,N_18844);
nand U19637 (N_19637,N_18718,N_18639);
or U19638 (N_19638,N_18852,N_18939);
xnor U19639 (N_19639,N_18792,N_19173);
and U19640 (N_19640,N_18692,N_18828);
nand U19641 (N_19641,N_18805,N_18827);
nor U19642 (N_19642,N_18967,N_19005);
nor U19643 (N_19643,N_19172,N_18953);
nand U19644 (N_19644,N_19125,N_18607);
xor U19645 (N_19645,N_18867,N_18914);
nor U19646 (N_19646,N_18766,N_19139);
and U19647 (N_19647,N_19113,N_18923);
xor U19648 (N_19648,N_18753,N_18783);
nor U19649 (N_19649,N_18797,N_18914);
nor U19650 (N_19650,N_18880,N_19142);
nand U19651 (N_19651,N_18673,N_18807);
or U19652 (N_19652,N_19187,N_18969);
nor U19653 (N_19653,N_19111,N_19143);
nor U19654 (N_19654,N_18652,N_18830);
nand U19655 (N_19655,N_18774,N_19140);
nand U19656 (N_19656,N_18641,N_18636);
nor U19657 (N_19657,N_18655,N_19160);
and U19658 (N_19658,N_18800,N_18725);
nor U19659 (N_19659,N_19141,N_19186);
or U19660 (N_19660,N_18738,N_19161);
xnor U19661 (N_19661,N_18841,N_18804);
nand U19662 (N_19662,N_18916,N_18907);
and U19663 (N_19663,N_18769,N_18789);
nor U19664 (N_19664,N_18680,N_18750);
nor U19665 (N_19665,N_19094,N_18717);
and U19666 (N_19666,N_18612,N_18971);
or U19667 (N_19667,N_18735,N_18759);
nor U19668 (N_19668,N_18669,N_18967);
nand U19669 (N_19669,N_19121,N_18770);
xnor U19670 (N_19670,N_18648,N_18767);
xor U19671 (N_19671,N_19182,N_18630);
xor U19672 (N_19672,N_18795,N_19120);
and U19673 (N_19673,N_18807,N_18963);
or U19674 (N_19674,N_18686,N_18727);
xnor U19675 (N_19675,N_19198,N_19161);
nor U19676 (N_19676,N_18653,N_18754);
nor U19677 (N_19677,N_19052,N_18957);
nand U19678 (N_19678,N_18603,N_18628);
nor U19679 (N_19679,N_18673,N_18947);
xor U19680 (N_19680,N_18987,N_19074);
xor U19681 (N_19681,N_19049,N_18897);
xor U19682 (N_19682,N_18755,N_18766);
and U19683 (N_19683,N_18830,N_18756);
nor U19684 (N_19684,N_19099,N_19156);
nor U19685 (N_19685,N_18891,N_18962);
or U19686 (N_19686,N_18803,N_19077);
nand U19687 (N_19687,N_18860,N_18797);
xnor U19688 (N_19688,N_18956,N_18792);
and U19689 (N_19689,N_18992,N_19061);
nor U19690 (N_19690,N_18963,N_19115);
nand U19691 (N_19691,N_18893,N_18749);
and U19692 (N_19692,N_18990,N_18866);
xnor U19693 (N_19693,N_18790,N_18781);
nand U19694 (N_19694,N_18727,N_18644);
nor U19695 (N_19695,N_18955,N_18691);
nand U19696 (N_19696,N_18852,N_19000);
xor U19697 (N_19697,N_19173,N_19092);
nand U19698 (N_19698,N_18924,N_18694);
or U19699 (N_19699,N_19174,N_18710);
nand U19700 (N_19700,N_18805,N_18903);
and U19701 (N_19701,N_18994,N_18789);
nand U19702 (N_19702,N_18985,N_18909);
xnor U19703 (N_19703,N_18631,N_18891);
xnor U19704 (N_19704,N_18975,N_18718);
nand U19705 (N_19705,N_19092,N_18999);
and U19706 (N_19706,N_18894,N_18850);
xnor U19707 (N_19707,N_18694,N_18942);
and U19708 (N_19708,N_18845,N_18975);
xnor U19709 (N_19709,N_19056,N_19081);
or U19710 (N_19710,N_18944,N_18808);
xnor U19711 (N_19711,N_18644,N_19114);
or U19712 (N_19712,N_18939,N_18740);
and U19713 (N_19713,N_19183,N_18845);
nor U19714 (N_19714,N_18888,N_19076);
or U19715 (N_19715,N_18798,N_19176);
or U19716 (N_19716,N_19003,N_18759);
nand U19717 (N_19717,N_19017,N_18699);
and U19718 (N_19718,N_18704,N_18959);
nor U19719 (N_19719,N_18894,N_18616);
xor U19720 (N_19720,N_19092,N_18879);
nor U19721 (N_19721,N_19060,N_19007);
and U19722 (N_19722,N_18939,N_18698);
xnor U19723 (N_19723,N_19027,N_19199);
xor U19724 (N_19724,N_18972,N_18854);
nand U19725 (N_19725,N_18979,N_19103);
nand U19726 (N_19726,N_19004,N_18999);
nand U19727 (N_19727,N_19145,N_18672);
and U19728 (N_19728,N_18949,N_18712);
xor U19729 (N_19729,N_18825,N_19139);
or U19730 (N_19730,N_18759,N_18654);
nand U19731 (N_19731,N_18761,N_19065);
and U19732 (N_19732,N_19066,N_18727);
or U19733 (N_19733,N_19007,N_18731);
and U19734 (N_19734,N_18860,N_19188);
xor U19735 (N_19735,N_18995,N_18679);
and U19736 (N_19736,N_19116,N_18967);
and U19737 (N_19737,N_18907,N_18905);
nand U19738 (N_19738,N_19063,N_18836);
xor U19739 (N_19739,N_18956,N_18945);
xnor U19740 (N_19740,N_18786,N_19094);
nor U19741 (N_19741,N_18989,N_18935);
nand U19742 (N_19742,N_19009,N_19078);
nor U19743 (N_19743,N_19049,N_18673);
and U19744 (N_19744,N_18872,N_18797);
xor U19745 (N_19745,N_19126,N_18935);
nor U19746 (N_19746,N_19056,N_18851);
and U19747 (N_19747,N_18603,N_19158);
nor U19748 (N_19748,N_18770,N_18772);
nand U19749 (N_19749,N_19195,N_18630);
and U19750 (N_19750,N_18904,N_19122);
nor U19751 (N_19751,N_18719,N_18987);
and U19752 (N_19752,N_18961,N_18709);
nor U19753 (N_19753,N_19039,N_19001);
or U19754 (N_19754,N_18836,N_18636);
and U19755 (N_19755,N_19156,N_18615);
and U19756 (N_19756,N_19170,N_18903);
nor U19757 (N_19757,N_19186,N_19147);
and U19758 (N_19758,N_19135,N_18859);
and U19759 (N_19759,N_18993,N_18928);
nor U19760 (N_19760,N_19079,N_18979);
nand U19761 (N_19761,N_18724,N_18773);
or U19762 (N_19762,N_19031,N_18757);
or U19763 (N_19763,N_19137,N_18966);
nand U19764 (N_19764,N_18970,N_18729);
or U19765 (N_19765,N_19002,N_19011);
nor U19766 (N_19766,N_19047,N_18726);
nand U19767 (N_19767,N_18779,N_19109);
xnor U19768 (N_19768,N_18949,N_19060);
nand U19769 (N_19769,N_19126,N_18661);
nand U19770 (N_19770,N_19114,N_18950);
nand U19771 (N_19771,N_18809,N_19105);
or U19772 (N_19772,N_18990,N_19018);
nand U19773 (N_19773,N_18922,N_18663);
nand U19774 (N_19774,N_19039,N_19028);
xnor U19775 (N_19775,N_18677,N_19047);
nand U19776 (N_19776,N_19018,N_18639);
and U19777 (N_19777,N_18745,N_18839);
and U19778 (N_19778,N_18776,N_18739);
xnor U19779 (N_19779,N_18845,N_19180);
nand U19780 (N_19780,N_19119,N_18805);
or U19781 (N_19781,N_18987,N_18910);
xor U19782 (N_19782,N_18911,N_18798);
nor U19783 (N_19783,N_19067,N_19116);
and U19784 (N_19784,N_18980,N_19161);
or U19785 (N_19785,N_18702,N_19127);
nand U19786 (N_19786,N_19025,N_18867);
and U19787 (N_19787,N_19065,N_18641);
or U19788 (N_19788,N_18633,N_19188);
and U19789 (N_19789,N_19126,N_18714);
or U19790 (N_19790,N_19093,N_19152);
nor U19791 (N_19791,N_18735,N_19030);
nor U19792 (N_19792,N_18862,N_19105);
and U19793 (N_19793,N_19090,N_19142);
xor U19794 (N_19794,N_18952,N_18616);
xor U19795 (N_19795,N_18963,N_19148);
nand U19796 (N_19796,N_19120,N_19141);
nor U19797 (N_19797,N_18958,N_18921);
or U19798 (N_19798,N_19183,N_18818);
nand U19799 (N_19799,N_19029,N_18691);
xnor U19800 (N_19800,N_19586,N_19628);
nand U19801 (N_19801,N_19278,N_19773);
nor U19802 (N_19802,N_19347,N_19638);
or U19803 (N_19803,N_19287,N_19616);
and U19804 (N_19804,N_19564,N_19537);
nand U19805 (N_19805,N_19512,N_19511);
nand U19806 (N_19806,N_19262,N_19644);
and U19807 (N_19807,N_19459,N_19795);
and U19808 (N_19808,N_19217,N_19552);
nand U19809 (N_19809,N_19781,N_19595);
or U19810 (N_19810,N_19211,N_19715);
nor U19811 (N_19811,N_19466,N_19786);
xor U19812 (N_19812,N_19239,N_19708);
nand U19813 (N_19813,N_19357,N_19299);
and U19814 (N_19814,N_19770,N_19697);
nor U19815 (N_19815,N_19676,N_19584);
xor U19816 (N_19816,N_19585,N_19452);
nor U19817 (N_19817,N_19738,N_19279);
nand U19818 (N_19818,N_19291,N_19304);
nand U19819 (N_19819,N_19369,N_19551);
nor U19820 (N_19820,N_19640,N_19367);
or U19821 (N_19821,N_19707,N_19723);
or U19822 (N_19822,N_19328,N_19475);
xnor U19823 (N_19823,N_19501,N_19763);
xor U19824 (N_19824,N_19416,N_19513);
nand U19825 (N_19825,N_19794,N_19264);
nand U19826 (N_19826,N_19486,N_19493);
or U19827 (N_19827,N_19360,N_19393);
and U19828 (N_19828,N_19222,N_19611);
xor U19829 (N_19829,N_19253,N_19547);
xor U19830 (N_19830,N_19687,N_19752);
or U19831 (N_19831,N_19320,N_19303);
xnor U19832 (N_19832,N_19508,N_19449);
nor U19833 (N_19833,N_19724,N_19240);
xor U19834 (N_19834,N_19775,N_19319);
or U19835 (N_19835,N_19623,N_19353);
nand U19836 (N_19836,N_19308,N_19296);
and U19837 (N_19837,N_19376,N_19377);
or U19838 (N_19838,N_19577,N_19588);
nand U19839 (N_19839,N_19364,N_19338);
and U19840 (N_19840,N_19448,N_19218);
and U19841 (N_19841,N_19249,N_19271);
nor U19842 (N_19842,N_19206,N_19515);
and U19843 (N_19843,N_19418,N_19562);
nand U19844 (N_19844,N_19387,N_19548);
xor U19845 (N_19845,N_19720,N_19470);
and U19846 (N_19846,N_19432,N_19390);
and U19847 (N_19847,N_19354,N_19429);
nand U19848 (N_19848,N_19256,N_19471);
nor U19849 (N_19849,N_19578,N_19659);
xor U19850 (N_19850,N_19517,N_19326);
or U19851 (N_19851,N_19612,N_19231);
nor U19852 (N_19852,N_19229,N_19745);
nand U19853 (N_19853,N_19252,N_19245);
xor U19854 (N_19854,N_19604,N_19686);
or U19855 (N_19855,N_19767,N_19779);
or U19856 (N_19856,N_19587,N_19619);
and U19857 (N_19857,N_19384,N_19570);
nor U19858 (N_19858,N_19583,N_19386);
nor U19859 (N_19859,N_19784,N_19212);
nor U19860 (N_19860,N_19241,N_19593);
xor U19861 (N_19861,N_19358,N_19257);
nand U19862 (N_19862,N_19395,N_19651);
nor U19863 (N_19863,N_19567,N_19719);
or U19864 (N_19864,N_19589,N_19569);
xor U19865 (N_19865,N_19625,N_19591);
or U19866 (N_19866,N_19747,N_19737);
xnor U19867 (N_19867,N_19757,N_19624);
or U19868 (N_19868,N_19679,N_19546);
and U19869 (N_19869,N_19435,N_19388);
and U19870 (N_19870,N_19414,N_19348);
and U19871 (N_19871,N_19615,N_19778);
nand U19872 (N_19872,N_19527,N_19467);
nand U19873 (N_19873,N_19629,N_19661);
nor U19874 (N_19874,N_19341,N_19209);
xor U19875 (N_19875,N_19221,N_19251);
xor U19876 (N_19876,N_19441,N_19283);
or U19877 (N_19877,N_19433,N_19285);
nor U19878 (N_19878,N_19571,N_19460);
nor U19879 (N_19879,N_19572,N_19729);
and U19880 (N_19880,N_19702,N_19714);
or U19881 (N_19881,N_19635,N_19465);
xnor U19882 (N_19882,N_19323,N_19622);
or U19883 (N_19883,N_19743,N_19728);
nor U19884 (N_19884,N_19607,N_19764);
nand U19885 (N_19885,N_19292,N_19761);
xnor U19886 (N_19886,N_19339,N_19771);
or U19887 (N_19887,N_19334,N_19399);
xnor U19888 (N_19888,N_19247,N_19646);
and U19889 (N_19889,N_19506,N_19561);
nand U19890 (N_19890,N_19361,N_19497);
nand U19891 (N_19891,N_19553,N_19754);
nand U19892 (N_19892,N_19523,N_19489);
nand U19893 (N_19893,N_19538,N_19421);
nor U19894 (N_19894,N_19404,N_19270);
and U19895 (N_19895,N_19605,N_19760);
or U19896 (N_19896,N_19539,N_19768);
or U19897 (N_19897,N_19397,N_19243);
or U19898 (N_19898,N_19600,N_19237);
nand U19899 (N_19899,N_19407,N_19782);
nor U19900 (N_19900,N_19409,N_19575);
and U19901 (N_19901,N_19261,N_19396);
nor U19902 (N_19902,N_19727,N_19558);
nand U19903 (N_19903,N_19370,N_19579);
xnor U19904 (N_19904,N_19453,N_19718);
nand U19905 (N_19905,N_19330,N_19563);
nor U19906 (N_19906,N_19477,N_19699);
or U19907 (N_19907,N_19474,N_19685);
xnor U19908 (N_19908,N_19735,N_19688);
nor U19909 (N_19909,N_19742,N_19700);
or U19910 (N_19910,N_19736,N_19550);
nor U19911 (N_19911,N_19603,N_19372);
nand U19912 (N_19912,N_19254,N_19214);
or U19913 (N_19913,N_19568,N_19434);
xor U19914 (N_19914,N_19238,N_19533);
or U19915 (N_19915,N_19457,N_19312);
xor U19916 (N_19916,N_19650,N_19705);
nand U19917 (N_19917,N_19645,N_19281);
nand U19918 (N_19918,N_19260,N_19207);
nor U19919 (N_19919,N_19630,N_19648);
nor U19920 (N_19920,N_19496,N_19510);
nand U19921 (N_19921,N_19725,N_19290);
or U19922 (N_19922,N_19535,N_19574);
nand U19923 (N_19923,N_19200,N_19317);
xor U19924 (N_19924,N_19282,N_19236);
nand U19925 (N_19925,N_19385,N_19636);
xnor U19926 (N_19926,N_19632,N_19665);
or U19927 (N_19927,N_19300,N_19244);
and U19928 (N_19928,N_19419,N_19355);
nor U19929 (N_19929,N_19488,N_19626);
xor U19930 (N_19930,N_19242,N_19494);
nand U19931 (N_19931,N_19318,N_19487);
and U19932 (N_19932,N_19726,N_19520);
xnor U19933 (N_19933,N_19371,N_19706);
nor U19934 (N_19934,N_19202,N_19374);
or U19935 (N_19935,N_19541,N_19756);
nor U19936 (N_19936,N_19451,N_19566);
and U19937 (N_19937,N_19352,N_19504);
or U19938 (N_19938,N_19447,N_19618);
nor U19939 (N_19939,N_19614,N_19730);
nand U19940 (N_19940,N_19509,N_19280);
xnor U19941 (N_19941,N_19643,N_19744);
nor U19942 (N_19942,N_19792,N_19713);
nand U19943 (N_19943,N_19694,N_19704);
nand U19944 (N_19944,N_19524,N_19581);
and U19945 (N_19945,N_19712,N_19529);
or U19946 (N_19946,N_19701,N_19542);
nor U19947 (N_19947,N_19669,N_19456);
nand U19948 (N_19948,N_19289,N_19780);
nand U19949 (N_19949,N_19215,N_19762);
nand U19950 (N_19950,N_19798,N_19598);
xnor U19951 (N_19951,N_19464,N_19309);
nand U19952 (N_19952,N_19220,N_19205);
nor U19953 (N_19953,N_19536,N_19398);
nor U19954 (N_19954,N_19759,N_19329);
or U19955 (N_19955,N_19343,N_19682);
nand U19956 (N_19956,N_19311,N_19325);
and U19957 (N_19957,N_19674,N_19430);
or U19958 (N_19958,N_19673,N_19381);
or U19959 (N_19959,N_19208,N_19431);
xor U19960 (N_19960,N_19305,N_19655);
or U19961 (N_19961,N_19484,N_19482);
nand U19962 (N_19962,N_19362,N_19755);
nand U19963 (N_19963,N_19783,N_19746);
nor U19964 (N_19964,N_19753,N_19350);
xor U19965 (N_19965,N_19427,N_19442);
nor U19966 (N_19966,N_19365,N_19525);
nand U19967 (N_19967,N_19286,N_19733);
or U19968 (N_19968,N_19491,N_19345);
and U19969 (N_19969,N_19473,N_19382);
or U19970 (N_19970,N_19225,N_19662);
and U19971 (N_19971,N_19408,N_19633);
nor U19972 (N_19972,N_19789,N_19695);
and U19973 (N_19973,N_19333,N_19500);
or U19974 (N_19974,N_19269,N_19392);
or U19975 (N_19975,N_19313,N_19703);
nand U19976 (N_19976,N_19670,N_19543);
nand U19977 (N_19977,N_19394,N_19481);
or U19978 (N_19978,N_19652,N_19267);
xor U19979 (N_19979,N_19710,N_19306);
xnor U19980 (N_19980,N_19446,N_19749);
or U19981 (N_19981,N_19734,N_19666);
and U19982 (N_19982,N_19219,N_19250);
nand U19983 (N_19983,N_19379,N_19716);
xnor U19984 (N_19984,N_19693,N_19223);
or U19985 (N_19985,N_19692,N_19438);
nor U19986 (N_19986,N_19660,N_19498);
nor U19987 (N_19987,N_19480,N_19627);
nor U19988 (N_19988,N_19265,N_19246);
xnor U19989 (N_19989,N_19336,N_19573);
or U19990 (N_19990,N_19791,N_19307);
or U19991 (N_19991,N_19732,N_19696);
nor U19992 (N_19992,N_19596,N_19272);
nor U19993 (N_19993,N_19521,N_19437);
nor U19994 (N_19994,N_19678,N_19788);
nand U19995 (N_19995,N_19601,N_19594);
nand U19996 (N_19996,N_19556,N_19263);
nor U19997 (N_19997,N_19213,N_19423);
nor U19998 (N_19998,N_19210,N_19540);
and U19999 (N_19999,N_19351,N_19672);
or U20000 (N_20000,N_19439,N_19620);
and U20001 (N_20001,N_19503,N_19717);
or U20002 (N_20002,N_19366,N_19656);
and U20003 (N_20003,N_19462,N_19776);
nor U20004 (N_20004,N_19444,N_19314);
nor U20005 (N_20005,N_19302,N_19445);
xnor U20006 (N_20006,N_19531,N_19232);
xor U20007 (N_20007,N_19297,N_19224);
or U20008 (N_20008,N_19436,N_19649);
and U20009 (N_20009,N_19664,N_19293);
nor U20010 (N_20010,N_19400,N_19201);
or U20011 (N_20011,N_19258,N_19310);
and U20012 (N_20012,N_19606,N_19301);
nand U20013 (N_20013,N_19534,N_19766);
and U20014 (N_20014,N_19335,N_19799);
nand U20015 (N_20015,N_19274,N_19751);
nor U20016 (N_20016,N_19476,N_19544);
and U20017 (N_20017,N_19592,N_19647);
xnor U20018 (N_20018,N_19610,N_19599);
and U20019 (N_20019,N_19580,N_19417);
and U20020 (N_20020,N_19765,N_19411);
nand U20021 (N_20021,N_19479,N_19582);
or U20022 (N_20022,N_19565,N_19458);
and U20023 (N_20023,N_19275,N_19322);
nor U20024 (N_20024,N_19492,N_19631);
or U20025 (N_20025,N_19425,N_19653);
nor U20026 (N_20026,N_19602,N_19346);
nand U20027 (N_20027,N_19739,N_19657);
nand U20028 (N_20028,N_19402,N_19454);
or U20029 (N_20029,N_19327,N_19518);
nor U20030 (N_20030,N_19722,N_19359);
nand U20031 (N_20031,N_19294,N_19405);
and U20032 (N_20032,N_19472,N_19298);
xor U20033 (N_20033,N_19519,N_19495);
nor U20034 (N_20034,N_19389,N_19331);
and U20035 (N_20035,N_19363,N_19516);
nor U20036 (N_20036,N_19787,N_19268);
and U20037 (N_20037,N_19741,N_19758);
xor U20038 (N_20038,N_19502,N_19671);
nor U20039 (N_20039,N_19637,N_19691);
or U20040 (N_20040,N_19420,N_19680);
nor U20041 (N_20041,N_19227,N_19711);
nor U20042 (N_20042,N_19677,N_19681);
and U20043 (N_20043,N_19777,N_19774);
nand U20044 (N_20044,N_19424,N_19684);
nand U20045 (N_20045,N_19796,N_19259);
nor U20046 (N_20046,N_19549,N_19654);
or U20047 (N_20047,N_19545,N_19609);
nor U20048 (N_20048,N_19793,N_19391);
and U20049 (N_20049,N_19797,N_19276);
nor U20050 (N_20050,N_19590,N_19203);
and U20051 (N_20051,N_19380,N_19748);
or U20052 (N_20052,N_19443,N_19639);
and U20053 (N_20053,N_19514,N_19698);
and U20054 (N_20054,N_19455,N_19288);
nor U20055 (N_20055,N_19641,N_19234);
xor U20056 (N_20056,N_19613,N_19248);
xor U20057 (N_20057,N_19528,N_19344);
nand U20058 (N_20058,N_19337,N_19356);
and U20059 (N_20059,N_19406,N_19373);
or U20060 (N_20060,N_19422,N_19230);
and U20061 (N_20061,N_19634,N_19532);
or U20062 (N_20062,N_19277,N_19204);
nor U20063 (N_20063,N_19663,N_19530);
xnor U20064 (N_20064,N_19284,N_19576);
nor U20065 (N_20065,N_19216,N_19560);
xor U20066 (N_20066,N_19235,N_19555);
or U20067 (N_20067,N_19316,N_19709);
and U20068 (N_20068,N_19233,N_19772);
nor U20069 (N_20069,N_19490,N_19315);
nand U20070 (N_20070,N_19642,N_19675);
nand U20071 (N_20071,N_19378,N_19426);
or U20072 (N_20072,N_19505,N_19507);
nor U20073 (N_20073,N_19324,N_19295);
and U20074 (N_20074,N_19368,N_19769);
or U20075 (N_20075,N_19428,N_19273);
and U20076 (N_20076,N_19483,N_19321);
xor U20077 (N_20077,N_19440,N_19468);
and U20078 (N_20078,N_19340,N_19554);
and U20079 (N_20079,N_19790,N_19750);
nand U20080 (N_20080,N_19478,N_19485);
and U20081 (N_20081,N_19557,N_19597);
or U20082 (N_20082,N_19667,N_19689);
and U20083 (N_20083,N_19463,N_19375);
nor U20084 (N_20084,N_19469,N_19415);
nand U20085 (N_20085,N_19403,N_19413);
nor U20086 (N_20086,N_19410,N_19658);
or U20087 (N_20087,N_19226,N_19461);
or U20088 (N_20088,N_19450,N_19342);
nand U20089 (N_20089,N_19332,N_19412);
or U20090 (N_20090,N_19617,N_19401);
xor U20091 (N_20091,N_19526,N_19266);
nand U20092 (N_20092,N_19499,N_19721);
and U20093 (N_20093,N_19608,N_19228);
nor U20094 (N_20094,N_19785,N_19559);
nor U20095 (N_20095,N_19383,N_19522);
nand U20096 (N_20096,N_19668,N_19255);
nand U20097 (N_20097,N_19683,N_19621);
xnor U20098 (N_20098,N_19690,N_19740);
or U20099 (N_20099,N_19731,N_19349);
or U20100 (N_20100,N_19632,N_19394);
nand U20101 (N_20101,N_19755,N_19677);
and U20102 (N_20102,N_19532,N_19391);
and U20103 (N_20103,N_19474,N_19783);
or U20104 (N_20104,N_19356,N_19273);
nor U20105 (N_20105,N_19462,N_19760);
xnor U20106 (N_20106,N_19789,N_19779);
nand U20107 (N_20107,N_19595,N_19667);
and U20108 (N_20108,N_19729,N_19712);
xnor U20109 (N_20109,N_19614,N_19585);
or U20110 (N_20110,N_19248,N_19580);
nor U20111 (N_20111,N_19667,N_19588);
xor U20112 (N_20112,N_19776,N_19248);
xnor U20113 (N_20113,N_19496,N_19306);
or U20114 (N_20114,N_19419,N_19723);
nand U20115 (N_20115,N_19634,N_19290);
nor U20116 (N_20116,N_19509,N_19540);
and U20117 (N_20117,N_19265,N_19659);
nand U20118 (N_20118,N_19377,N_19260);
and U20119 (N_20119,N_19303,N_19423);
xnor U20120 (N_20120,N_19442,N_19628);
xnor U20121 (N_20121,N_19676,N_19767);
and U20122 (N_20122,N_19591,N_19416);
nor U20123 (N_20123,N_19740,N_19364);
xnor U20124 (N_20124,N_19281,N_19539);
and U20125 (N_20125,N_19488,N_19698);
or U20126 (N_20126,N_19398,N_19617);
xnor U20127 (N_20127,N_19521,N_19710);
nand U20128 (N_20128,N_19396,N_19680);
nor U20129 (N_20129,N_19236,N_19726);
nor U20130 (N_20130,N_19536,N_19437);
nor U20131 (N_20131,N_19799,N_19406);
nand U20132 (N_20132,N_19269,N_19429);
xnor U20133 (N_20133,N_19729,N_19746);
nor U20134 (N_20134,N_19730,N_19591);
and U20135 (N_20135,N_19646,N_19512);
or U20136 (N_20136,N_19364,N_19601);
or U20137 (N_20137,N_19615,N_19462);
or U20138 (N_20138,N_19458,N_19309);
and U20139 (N_20139,N_19213,N_19773);
nor U20140 (N_20140,N_19262,N_19457);
and U20141 (N_20141,N_19295,N_19757);
nand U20142 (N_20142,N_19637,N_19606);
nor U20143 (N_20143,N_19474,N_19490);
or U20144 (N_20144,N_19236,N_19222);
nand U20145 (N_20145,N_19745,N_19403);
nand U20146 (N_20146,N_19547,N_19244);
or U20147 (N_20147,N_19268,N_19376);
or U20148 (N_20148,N_19668,N_19321);
nand U20149 (N_20149,N_19504,N_19396);
xor U20150 (N_20150,N_19729,N_19507);
nor U20151 (N_20151,N_19507,N_19736);
nor U20152 (N_20152,N_19462,N_19494);
nor U20153 (N_20153,N_19217,N_19705);
nand U20154 (N_20154,N_19541,N_19393);
nand U20155 (N_20155,N_19348,N_19301);
nand U20156 (N_20156,N_19787,N_19306);
nand U20157 (N_20157,N_19656,N_19265);
and U20158 (N_20158,N_19705,N_19584);
nand U20159 (N_20159,N_19593,N_19493);
xnor U20160 (N_20160,N_19541,N_19450);
and U20161 (N_20161,N_19780,N_19396);
or U20162 (N_20162,N_19621,N_19331);
xnor U20163 (N_20163,N_19550,N_19433);
xor U20164 (N_20164,N_19586,N_19797);
or U20165 (N_20165,N_19578,N_19438);
nor U20166 (N_20166,N_19776,N_19211);
and U20167 (N_20167,N_19565,N_19718);
nor U20168 (N_20168,N_19513,N_19209);
nand U20169 (N_20169,N_19584,N_19718);
xnor U20170 (N_20170,N_19390,N_19220);
xor U20171 (N_20171,N_19560,N_19484);
and U20172 (N_20172,N_19539,N_19414);
and U20173 (N_20173,N_19259,N_19512);
and U20174 (N_20174,N_19263,N_19555);
nand U20175 (N_20175,N_19719,N_19404);
nand U20176 (N_20176,N_19439,N_19734);
nand U20177 (N_20177,N_19596,N_19610);
xor U20178 (N_20178,N_19641,N_19534);
nand U20179 (N_20179,N_19688,N_19732);
xor U20180 (N_20180,N_19284,N_19429);
xor U20181 (N_20181,N_19747,N_19497);
xor U20182 (N_20182,N_19399,N_19724);
nand U20183 (N_20183,N_19741,N_19670);
and U20184 (N_20184,N_19414,N_19496);
xnor U20185 (N_20185,N_19731,N_19723);
or U20186 (N_20186,N_19308,N_19568);
and U20187 (N_20187,N_19643,N_19758);
xnor U20188 (N_20188,N_19334,N_19248);
xnor U20189 (N_20189,N_19754,N_19225);
or U20190 (N_20190,N_19245,N_19766);
xor U20191 (N_20191,N_19289,N_19635);
nand U20192 (N_20192,N_19464,N_19683);
nand U20193 (N_20193,N_19238,N_19675);
xor U20194 (N_20194,N_19259,N_19642);
and U20195 (N_20195,N_19431,N_19552);
xor U20196 (N_20196,N_19743,N_19676);
nand U20197 (N_20197,N_19404,N_19712);
xor U20198 (N_20198,N_19519,N_19660);
nand U20199 (N_20199,N_19231,N_19312);
and U20200 (N_20200,N_19262,N_19590);
nor U20201 (N_20201,N_19201,N_19776);
nand U20202 (N_20202,N_19376,N_19764);
nor U20203 (N_20203,N_19638,N_19649);
and U20204 (N_20204,N_19571,N_19755);
xnor U20205 (N_20205,N_19687,N_19732);
and U20206 (N_20206,N_19533,N_19504);
nand U20207 (N_20207,N_19545,N_19418);
or U20208 (N_20208,N_19765,N_19246);
nor U20209 (N_20209,N_19535,N_19728);
nand U20210 (N_20210,N_19403,N_19218);
or U20211 (N_20211,N_19411,N_19519);
nor U20212 (N_20212,N_19724,N_19248);
xnor U20213 (N_20213,N_19729,N_19279);
and U20214 (N_20214,N_19547,N_19269);
xnor U20215 (N_20215,N_19271,N_19552);
nor U20216 (N_20216,N_19493,N_19609);
and U20217 (N_20217,N_19680,N_19631);
nor U20218 (N_20218,N_19615,N_19319);
nor U20219 (N_20219,N_19209,N_19661);
and U20220 (N_20220,N_19721,N_19248);
nand U20221 (N_20221,N_19791,N_19765);
xnor U20222 (N_20222,N_19446,N_19668);
xnor U20223 (N_20223,N_19698,N_19497);
xor U20224 (N_20224,N_19759,N_19429);
xnor U20225 (N_20225,N_19279,N_19349);
nor U20226 (N_20226,N_19736,N_19751);
nand U20227 (N_20227,N_19726,N_19343);
or U20228 (N_20228,N_19211,N_19728);
nor U20229 (N_20229,N_19440,N_19502);
xnor U20230 (N_20230,N_19769,N_19545);
and U20231 (N_20231,N_19474,N_19264);
xnor U20232 (N_20232,N_19238,N_19661);
nor U20233 (N_20233,N_19691,N_19363);
or U20234 (N_20234,N_19743,N_19301);
and U20235 (N_20235,N_19429,N_19635);
nor U20236 (N_20236,N_19743,N_19555);
nor U20237 (N_20237,N_19758,N_19688);
nand U20238 (N_20238,N_19451,N_19733);
nand U20239 (N_20239,N_19709,N_19542);
and U20240 (N_20240,N_19406,N_19363);
and U20241 (N_20241,N_19634,N_19742);
nand U20242 (N_20242,N_19640,N_19551);
xnor U20243 (N_20243,N_19227,N_19309);
nor U20244 (N_20244,N_19430,N_19216);
nand U20245 (N_20245,N_19628,N_19359);
and U20246 (N_20246,N_19710,N_19698);
nor U20247 (N_20247,N_19201,N_19223);
and U20248 (N_20248,N_19792,N_19652);
nand U20249 (N_20249,N_19351,N_19578);
and U20250 (N_20250,N_19633,N_19470);
nand U20251 (N_20251,N_19700,N_19441);
and U20252 (N_20252,N_19316,N_19213);
nand U20253 (N_20253,N_19628,N_19544);
xor U20254 (N_20254,N_19516,N_19756);
xnor U20255 (N_20255,N_19367,N_19290);
nor U20256 (N_20256,N_19762,N_19457);
or U20257 (N_20257,N_19201,N_19358);
and U20258 (N_20258,N_19339,N_19655);
or U20259 (N_20259,N_19544,N_19271);
or U20260 (N_20260,N_19799,N_19615);
nand U20261 (N_20261,N_19574,N_19618);
and U20262 (N_20262,N_19283,N_19765);
nand U20263 (N_20263,N_19790,N_19765);
xor U20264 (N_20264,N_19554,N_19683);
nor U20265 (N_20265,N_19497,N_19591);
xnor U20266 (N_20266,N_19346,N_19364);
or U20267 (N_20267,N_19700,N_19622);
nor U20268 (N_20268,N_19712,N_19786);
nand U20269 (N_20269,N_19655,N_19256);
or U20270 (N_20270,N_19608,N_19309);
xor U20271 (N_20271,N_19234,N_19493);
or U20272 (N_20272,N_19418,N_19583);
nand U20273 (N_20273,N_19268,N_19741);
nand U20274 (N_20274,N_19218,N_19548);
nand U20275 (N_20275,N_19522,N_19707);
and U20276 (N_20276,N_19326,N_19332);
and U20277 (N_20277,N_19560,N_19380);
nand U20278 (N_20278,N_19601,N_19665);
or U20279 (N_20279,N_19615,N_19257);
nand U20280 (N_20280,N_19458,N_19272);
nand U20281 (N_20281,N_19439,N_19374);
nor U20282 (N_20282,N_19384,N_19666);
or U20283 (N_20283,N_19734,N_19540);
and U20284 (N_20284,N_19660,N_19240);
and U20285 (N_20285,N_19767,N_19511);
nand U20286 (N_20286,N_19352,N_19747);
or U20287 (N_20287,N_19510,N_19681);
or U20288 (N_20288,N_19254,N_19502);
xnor U20289 (N_20289,N_19260,N_19395);
xnor U20290 (N_20290,N_19275,N_19786);
and U20291 (N_20291,N_19215,N_19450);
nand U20292 (N_20292,N_19394,N_19682);
nor U20293 (N_20293,N_19653,N_19271);
nor U20294 (N_20294,N_19339,N_19450);
or U20295 (N_20295,N_19451,N_19789);
nor U20296 (N_20296,N_19257,N_19577);
nor U20297 (N_20297,N_19757,N_19449);
nand U20298 (N_20298,N_19729,N_19776);
or U20299 (N_20299,N_19641,N_19693);
xnor U20300 (N_20300,N_19374,N_19310);
nand U20301 (N_20301,N_19557,N_19643);
nor U20302 (N_20302,N_19744,N_19559);
xnor U20303 (N_20303,N_19678,N_19776);
nor U20304 (N_20304,N_19651,N_19432);
nand U20305 (N_20305,N_19251,N_19378);
and U20306 (N_20306,N_19255,N_19324);
nand U20307 (N_20307,N_19627,N_19216);
nor U20308 (N_20308,N_19516,N_19254);
or U20309 (N_20309,N_19215,N_19448);
nor U20310 (N_20310,N_19776,N_19755);
nand U20311 (N_20311,N_19562,N_19288);
xnor U20312 (N_20312,N_19506,N_19289);
nand U20313 (N_20313,N_19350,N_19741);
nand U20314 (N_20314,N_19723,N_19398);
and U20315 (N_20315,N_19480,N_19459);
and U20316 (N_20316,N_19289,N_19503);
or U20317 (N_20317,N_19693,N_19769);
nand U20318 (N_20318,N_19204,N_19256);
nand U20319 (N_20319,N_19226,N_19675);
nor U20320 (N_20320,N_19404,N_19462);
and U20321 (N_20321,N_19457,N_19319);
and U20322 (N_20322,N_19463,N_19380);
nor U20323 (N_20323,N_19778,N_19376);
xor U20324 (N_20324,N_19714,N_19402);
xnor U20325 (N_20325,N_19787,N_19263);
xnor U20326 (N_20326,N_19512,N_19592);
nand U20327 (N_20327,N_19791,N_19404);
nand U20328 (N_20328,N_19561,N_19395);
or U20329 (N_20329,N_19750,N_19469);
nand U20330 (N_20330,N_19328,N_19655);
nand U20331 (N_20331,N_19450,N_19744);
or U20332 (N_20332,N_19641,N_19338);
or U20333 (N_20333,N_19607,N_19475);
or U20334 (N_20334,N_19296,N_19227);
or U20335 (N_20335,N_19776,N_19406);
nand U20336 (N_20336,N_19778,N_19478);
nand U20337 (N_20337,N_19662,N_19715);
xor U20338 (N_20338,N_19437,N_19760);
nand U20339 (N_20339,N_19540,N_19453);
nor U20340 (N_20340,N_19281,N_19458);
and U20341 (N_20341,N_19499,N_19779);
nand U20342 (N_20342,N_19586,N_19566);
nor U20343 (N_20343,N_19544,N_19515);
or U20344 (N_20344,N_19535,N_19679);
nor U20345 (N_20345,N_19412,N_19609);
nor U20346 (N_20346,N_19329,N_19262);
nor U20347 (N_20347,N_19794,N_19239);
and U20348 (N_20348,N_19444,N_19406);
nand U20349 (N_20349,N_19448,N_19525);
xor U20350 (N_20350,N_19789,N_19230);
nand U20351 (N_20351,N_19459,N_19441);
nor U20352 (N_20352,N_19410,N_19348);
or U20353 (N_20353,N_19705,N_19455);
xnor U20354 (N_20354,N_19603,N_19589);
xnor U20355 (N_20355,N_19238,N_19674);
or U20356 (N_20356,N_19675,N_19361);
nor U20357 (N_20357,N_19422,N_19725);
and U20358 (N_20358,N_19293,N_19373);
nor U20359 (N_20359,N_19707,N_19455);
xor U20360 (N_20360,N_19268,N_19679);
and U20361 (N_20361,N_19296,N_19336);
nor U20362 (N_20362,N_19401,N_19204);
nand U20363 (N_20363,N_19295,N_19231);
nand U20364 (N_20364,N_19571,N_19444);
or U20365 (N_20365,N_19788,N_19413);
or U20366 (N_20366,N_19292,N_19700);
nor U20367 (N_20367,N_19766,N_19473);
nor U20368 (N_20368,N_19795,N_19211);
or U20369 (N_20369,N_19615,N_19502);
nand U20370 (N_20370,N_19227,N_19467);
nand U20371 (N_20371,N_19293,N_19273);
or U20372 (N_20372,N_19696,N_19618);
nand U20373 (N_20373,N_19463,N_19715);
xor U20374 (N_20374,N_19432,N_19691);
or U20375 (N_20375,N_19420,N_19251);
nand U20376 (N_20376,N_19495,N_19647);
and U20377 (N_20377,N_19224,N_19598);
or U20378 (N_20378,N_19784,N_19569);
nor U20379 (N_20379,N_19612,N_19386);
or U20380 (N_20380,N_19480,N_19235);
nor U20381 (N_20381,N_19582,N_19214);
nand U20382 (N_20382,N_19229,N_19736);
xnor U20383 (N_20383,N_19352,N_19493);
xnor U20384 (N_20384,N_19521,N_19608);
and U20385 (N_20385,N_19765,N_19546);
or U20386 (N_20386,N_19252,N_19524);
nor U20387 (N_20387,N_19217,N_19283);
xor U20388 (N_20388,N_19487,N_19203);
nand U20389 (N_20389,N_19437,N_19640);
and U20390 (N_20390,N_19594,N_19418);
nor U20391 (N_20391,N_19523,N_19647);
and U20392 (N_20392,N_19547,N_19768);
or U20393 (N_20393,N_19540,N_19450);
nand U20394 (N_20394,N_19766,N_19518);
and U20395 (N_20395,N_19363,N_19546);
xnor U20396 (N_20396,N_19632,N_19713);
xnor U20397 (N_20397,N_19578,N_19464);
and U20398 (N_20398,N_19719,N_19222);
xor U20399 (N_20399,N_19539,N_19288);
and U20400 (N_20400,N_20177,N_19856);
xor U20401 (N_20401,N_19863,N_20370);
nand U20402 (N_20402,N_19809,N_19855);
and U20403 (N_20403,N_20198,N_19964);
or U20404 (N_20404,N_20331,N_20297);
or U20405 (N_20405,N_20244,N_20038);
nand U20406 (N_20406,N_20360,N_20340);
xnor U20407 (N_20407,N_20287,N_20067);
nand U20408 (N_20408,N_19847,N_19985);
nor U20409 (N_20409,N_19821,N_20023);
and U20410 (N_20410,N_19909,N_19858);
nand U20411 (N_20411,N_20006,N_20127);
or U20412 (N_20412,N_19984,N_20396);
xor U20413 (N_20413,N_20384,N_20211);
nand U20414 (N_20414,N_20276,N_20111);
nand U20415 (N_20415,N_20153,N_20356);
or U20416 (N_20416,N_20344,N_20274);
or U20417 (N_20417,N_20329,N_19830);
nand U20418 (N_20418,N_19944,N_20323);
nand U20419 (N_20419,N_20107,N_19945);
xnor U20420 (N_20420,N_19882,N_20029);
nand U20421 (N_20421,N_20358,N_19831);
or U20422 (N_20422,N_19921,N_20118);
xor U20423 (N_20423,N_20199,N_20052);
and U20424 (N_20424,N_19886,N_20366);
or U20425 (N_20425,N_20385,N_20005);
or U20426 (N_20426,N_20001,N_20306);
or U20427 (N_20427,N_20232,N_20392);
and U20428 (N_20428,N_20075,N_20255);
nor U20429 (N_20429,N_20129,N_20295);
or U20430 (N_20430,N_20395,N_20030);
and U20431 (N_20431,N_20321,N_19851);
and U20432 (N_20432,N_19829,N_19973);
and U20433 (N_20433,N_19881,N_19942);
or U20434 (N_20434,N_20182,N_20151);
nor U20435 (N_20435,N_19982,N_19865);
nor U20436 (N_20436,N_20156,N_19839);
or U20437 (N_20437,N_19998,N_20026);
nand U20438 (N_20438,N_20173,N_20221);
nor U20439 (N_20439,N_19841,N_20377);
nand U20440 (N_20440,N_20311,N_19864);
or U20441 (N_20441,N_20263,N_20109);
nor U20442 (N_20442,N_20234,N_20120);
or U20443 (N_20443,N_20355,N_20298);
xor U20444 (N_20444,N_19896,N_20175);
nand U20445 (N_20445,N_19903,N_19801);
xnor U20446 (N_20446,N_20246,N_20349);
and U20447 (N_20447,N_20167,N_19978);
nor U20448 (N_20448,N_20291,N_19980);
or U20449 (N_20449,N_20197,N_20378);
and U20450 (N_20450,N_19836,N_19954);
nor U20451 (N_20451,N_20205,N_19916);
and U20452 (N_20452,N_19806,N_20169);
or U20453 (N_20453,N_19871,N_20228);
and U20454 (N_20454,N_20288,N_20050);
nand U20455 (N_20455,N_19861,N_20243);
or U20456 (N_20456,N_20130,N_19956);
or U20457 (N_20457,N_19825,N_20119);
xor U20458 (N_20458,N_19827,N_19991);
nand U20459 (N_20459,N_19986,N_19877);
nor U20460 (N_20460,N_19887,N_20284);
nand U20461 (N_20461,N_19893,N_20210);
and U20462 (N_20462,N_19845,N_19884);
and U20463 (N_20463,N_19907,N_20148);
or U20464 (N_20464,N_19899,N_19835);
and U20465 (N_20465,N_20278,N_20047);
or U20466 (N_20466,N_20171,N_20270);
or U20467 (N_20467,N_20319,N_19930);
nand U20468 (N_20468,N_20230,N_19925);
nor U20469 (N_20469,N_20131,N_20055);
nand U20470 (N_20470,N_20213,N_19878);
xor U20471 (N_20471,N_20369,N_20231);
or U20472 (N_20472,N_19838,N_20147);
and U20473 (N_20473,N_20084,N_20086);
or U20474 (N_20474,N_20379,N_19940);
or U20475 (N_20475,N_20176,N_20240);
nor U20476 (N_20476,N_20304,N_20303);
nor U20477 (N_20477,N_19804,N_19805);
and U20478 (N_20478,N_19949,N_20172);
or U20479 (N_20479,N_20054,N_19815);
and U20480 (N_20480,N_19823,N_19876);
or U20481 (N_20481,N_20092,N_20196);
nor U20482 (N_20482,N_19912,N_20381);
nand U20483 (N_20483,N_20122,N_20053);
nor U20484 (N_20484,N_20114,N_20397);
xnor U20485 (N_20485,N_19832,N_20202);
or U20486 (N_20486,N_20324,N_20302);
or U20487 (N_20487,N_20218,N_19950);
nand U20488 (N_20488,N_19869,N_20040);
or U20489 (N_20489,N_19901,N_20179);
nor U20490 (N_20490,N_20194,N_20066);
and U20491 (N_20491,N_20007,N_20265);
nor U20492 (N_20492,N_19853,N_20165);
nor U20493 (N_20493,N_20168,N_20024);
or U20494 (N_20494,N_20383,N_20341);
xnor U20495 (N_20495,N_19946,N_20308);
nor U20496 (N_20496,N_20280,N_19852);
nor U20497 (N_20497,N_20162,N_20241);
xnor U20498 (N_20498,N_20330,N_19818);
nor U20499 (N_20499,N_20138,N_19943);
and U20500 (N_20500,N_20248,N_20154);
and U20501 (N_20501,N_20252,N_19834);
nor U20502 (N_20502,N_19933,N_20277);
xnor U20503 (N_20503,N_19898,N_20192);
xnor U20504 (N_20504,N_19977,N_19807);
or U20505 (N_20505,N_20335,N_19971);
nor U20506 (N_20506,N_19968,N_20368);
xor U20507 (N_20507,N_20032,N_20217);
or U20508 (N_20508,N_20065,N_20025);
nand U20509 (N_20509,N_20078,N_20388);
xnor U20510 (N_20510,N_20017,N_19873);
nand U20511 (N_20511,N_19974,N_20108);
nand U20512 (N_20512,N_20314,N_20002);
or U20513 (N_20513,N_20039,N_20170);
nand U20514 (N_20514,N_20071,N_19872);
xor U20515 (N_20515,N_20037,N_20019);
and U20516 (N_20516,N_20364,N_19868);
nand U20517 (N_20517,N_20031,N_20296);
nand U20518 (N_20518,N_20352,N_19953);
nand U20519 (N_20519,N_20375,N_20160);
xnor U20520 (N_20520,N_20088,N_20227);
and U20521 (N_20521,N_19867,N_20016);
nor U20522 (N_20522,N_20236,N_19824);
or U20523 (N_20523,N_20313,N_19892);
nand U20524 (N_20524,N_19965,N_19914);
nand U20525 (N_20525,N_19843,N_20262);
and U20526 (N_20526,N_20091,N_20376);
xor U20527 (N_20527,N_19883,N_20080);
nor U20528 (N_20528,N_20081,N_20100);
nand U20529 (N_20529,N_20336,N_20022);
nor U20530 (N_20530,N_19961,N_20027);
nand U20531 (N_20531,N_20000,N_20258);
and U20532 (N_20532,N_20159,N_20020);
xor U20533 (N_20533,N_19981,N_19890);
nand U20534 (N_20534,N_20203,N_19814);
and U20535 (N_20535,N_19939,N_20391);
xor U20536 (N_20536,N_19959,N_19811);
nor U20537 (N_20537,N_20191,N_19850);
nor U20538 (N_20538,N_20178,N_20134);
nor U20539 (N_20539,N_20099,N_20286);
or U20540 (N_20540,N_19894,N_19996);
xnor U20541 (N_20541,N_20103,N_20214);
nand U20542 (N_20542,N_19957,N_20174);
nor U20543 (N_20543,N_20294,N_20390);
and U20544 (N_20544,N_20184,N_20215);
and U20545 (N_20545,N_20056,N_19803);
and U20546 (N_20546,N_20018,N_20393);
nand U20547 (N_20547,N_19920,N_20097);
xnor U20548 (N_20548,N_20312,N_19888);
xnor U20549 (N_20549,N_19857,N_20036);
xnor U20550 (N_20550,N_19926,N_20189);
or U20551 (N_20551,N_19817,N_20328);
nor U20552 (N_20552,N_19849,N_20074);
and U20553 (N_20553,N_19862,N_20133);
and U20554 (N_20554,N_20326,N_20365);
nand U20555 (N_20555,N_20150,N_19922);
nand U20556 (N_20556,N_19951,N_20155);
or U20557 (N_20557,N_20290,N_20212);
or U20558 (N_20558,N_20141,N_19948);
nand U20559 (N_20559,N_20389,N_20094);
or U20560 (N_20560,N_20206,N_20220);
and U20561 (N_20561,N_20046,N_20117);
or U20562 (N_20562,N_20062,N_19975);
nor U20563 (N_20563,N_20116,N_20207);
or U20564 (N_20564,N_19812,N_20098);
and U20565 (N_20565,N_20110,N_20204);
and U20566 (N_20566,N_20282,N_20200);
and U20567 (N_20567,N_19875,N_19859);
nor U20568 (N_20568,N_20250,N_20193);
or U20569 (N_20569,N_20216,N_20301);
nand U20570 (N_20570,N_20157,N_20361);
nor U20571 (N_20571,N_20073,N_20112);
nand U20572 (N_20572,N_20051,N_20322);
or U20573 (N_20573,N_20043,N_19923);
or U20574 (N_20574,N_20354,N_20042);
and U20575 (N_20575,N_20337,N_20253);
nand U20576 (N_20576,N_20195,N_20223);
nand U20577 (N_20577,N_20013,N_20269);
and U20578 (N_20578,N_20180,N_20123);
xnor U20579 (N_20579,N_20229,N_19905);
and U20580 (N_20580,N_20093,N_20140);
xor U20581 (N_20581,N_20267,N_20143);
and U20582 (N_20582,N_20069,N_20342);
and U20583 (N_20583,N_19826,N_20096);
xor U20584 (N_20584,N_20316,N_20333);
or U20585 (N_20585,N_20224,N_20345);
or U20586 (N_20586,N_20318,N_20394);
and U20587 (N_20587,N_20310,N_20264);
and U20588 (N_20588,N_19902,N_19908);
nor U20589 (N_20589,N_20359,N_19937);
and U20590 (N_20590,N_19919,N_19990);
xnor U20591 (N_20591,N_19983,N_20187);
nand U20592 (N_20592,N_20257,N_19938);
and U20593 (N_20593,N_20315,N_20163);
nor U20594 (N_20594,N_20064,N_20079);
nor U20595 (N_20595,N_20095,N_20233);
nand U20596 (N_20596,N_20146,N_20374);
or U20597 (N_20597,N_20063,N_20219);
and U20598 (N_20598,N_20372,N_19960);
or U20599 (N_20599,N_20072,N_20279);
xnor U20600 (N_20600,N_19988,N_19987);
xnor U20601 (N_20601,N_20136,N_20259);
or U20602 (N_20602,N_20251,N_19935);
or U20603 (N_20603,N_19844,N_19989);
or U20604 (N_20604,N_20222,N_20382);
and U20605 (N_20605,N_20149,N_19879);
xnor U20606 (N_20606,N_20346,N_20083);
nor U20607 (N_20607,N_20371,N_20158);
and U20608 (N_20608,N_19917,N_20380);
nand U20609 (N_20609,N_19928,N_20077);
nand U20610 (N_20610,N_19816,N_19979);
or U20611 (N_20611,N_19870,N_20049);
nor U20612 (N_20612,N_20208,N_19885);
xor U20613 (N_20613,N_19936,N_20106);
and U20614 (N_20614,N_20033,N_20059);
xor U20615 (N_20615,N_19958,N_20285);
nand U20616 (N_20616,N_20239,N_20363);
and U20617 (N_20617,N_19952,N_19810);
and U20618 (N_20618,N_20237,N_20045);
xor U20619 (N_20619,N_20261,N_20003);
xnor U20620 (N_20620,N_19913,N_20028);
or U20621 (N_20621,N_20113,N_20087);
nand U20622 (N_20622,N_20044,N_19995);
or U20623 (N_20623,N_19889,N_19932);
nor U20624 (N_20624,N_19891,N_19822);
xnor U20625 (N_20625,N_20089,N_19941);
and U20626 (N_20626,N_20142,N_20254);
nor U20627 (N_20627,N_20128,N_20351);
xnor U20628 (N_20628,N_19904,N_19842);
and U20629 (N_20629,N_19915,N_20137);
nand U20630 (N_20630,N_19846,N_20293);
or U20631 (N_20631,N_20268,N_20161);
nor U20632 (N_20632,N_20034,N_20343);
or U20633 (N_20633,N_19874,N_20058);
and U20634 (N_20634,N_19963,N_20144);
xor U20635 (N_20635,N_20266,N_20009);
and U20636 (N_20636,N_19994,N_19929);
xor U20637 (N_20637,N_19906,N_19970);
and U20638 (N_20638,N_20090,N_19802);
or U20639 (N_20639,N_20362,N_20320);
nor U20640 (N_20640,N_20183,N_19808);
xor U20641 (N_20641,N_19800,N_20152);
nand U20642 (N_20642,N_20076,N_20225);
or U20643 (N_20643,N_20014,N_20102);
or U20644 (N_20644,N_20338,N_20386);
nor U20645 (N_20645,N_20008,N_19924);
or U20646 (N_20646,N_20048,N_20132);
nor U20647 (N_20647,N_19934,N_19927);
nor U20648 (N_20648,N_20373,N_20135);
xor U20649 (N_20649,N_19976,N_20188);
xnor U20650 (N_20650,N_19880,N_20299);
or U20651 (N_20651,N_20367,N_20387);
nor U20652 (N_20652,N_19997,N_19895);
and U20653 (N_20653,N_20357,N_20256);
xor U20654 (N_20654,N_19962,N_20347);
nor U20655 (N_20655,N_20300,N_19897);
nand U20656 (N_20656,N_20125,N_20260);
and U20657 (N_20657,N_19999,N_19910);
and U20658 (N_20658,N_20010,N_20325);
and U20659 (N_20659,N_19860,N_20101);
and U20660 (N_20660,N_19966,N_20115);
or U20661 (N_20661,N_20275,N_20104);
nor U20662 (N_20662,N_20035,N_20245);
nor U20663 (N_20663,N_20166,N_20070);
nor U20664 (N_20664,N_20350,N_20082);
xnor U20665 (N_20665,N_19955,N_20281);
nand U20666 (N_20666,N_20307,N_19828);
and U20667 (N_20667,N_20126,N_20249);
xor U20668 (N_20668,N_19947,N_20121);
nand U20669 (N_20669,N_20012,N_20353);
xnor U20670 (N_20670,N_20317,N_20057);
nor U20671 (N_20671,N_20209,N_19967);
xor U20672 (N_20672,N_20021,N_19854);
and U20673 (N_20673,N_20011,N_19918);
and U20674 (N_20674,N_20061,N_20272);
and U20675 (N_20675,N_20238,N_19931);
nor U20676 (N_20676,N_19833,N_20305);
nand U20677 (N_20677,N_19866,N_19972);
nand U20678 (N_20678,N_20348,N_20041);
or U20679 (N_20679,N_19819,N_19911);
nor U20680 (N_20680,N_20085,N_19848);
or U20681 (N_20681,N_19992,N_19840);
xor U20682 (N_20682,N_20004,N_20181);
and U20683 (N_20683,N_20124,N_19813);
and U20684 (N_20684,N_19969,N_20068);
xor U20685 (N_20685,N_20145,N_20332);
and U20686 (N_20686,N_20060,N_20247);
or U20687 (N_20687,N_20201,N_20242);
xnor U20688 (N_20688,N_20273,N_20015);
or U20689 (N_20689,N_19900,N_20334);
or U20690 (N_20690,N_20235,N_20190);
nand U20691 (N_20691,N_20226,N_20292);
nor U20692 (N_20692,N_20185,N_19993);
nand U20693 (N_20693,N_20399,N_20289);
or U20694 (N_20694,N_20105,N_20186);
xnor U20695 (N_20695,N_20398,N_19820);
xor U20696 (N_20696,N_20164,N_20339);
nand U20697 (N_20697,N_20309,N_19837);
nand U20698 (N_20698,N_20327,N_20271);
xnor U20699 (N_20699,N_20139,N_20283);
or U20700 (N_20700,N_19976,N_19999);
or U20701 (N_20701,N_20016,N_20096);
nor U20702 (N_20702,N_20174,N_20188);
and U20703 (N_20703,N_20354,N_20217);
xor U20704 (N_20704,N_19824,N_20389);
nand U20705 (N_20705,N_20228,N_19951);
and U20706 (N_20706,N_20374,N_20088);
nor U20707 (N_20707,N_20343,N_20061);
xnor U20708 (N_20708,N_19966,N_19866);
nor U20709 (N_20709,N_19994,N_19901);
and U20710 (N_20710,N_19807,N_19976);
nor U20711 (N_20711,N_20330,N_20245);
xor U20712 (N_20712,N_19939,N_19959);
nand U20713 (N_20713,N_19938,N_20087);
nor U20714 (N_20714,N_20279,N_20284);
nand U20715 (N_20715,N_20277,N_20075);
or U20716 (N_20716,N_20075,N_20133);
xor U20717 (N_20717,N_19848,N_20052);
or U20718 (N_20718,N_19984,N_19941);
nor U20719 (N_20719,N_20219,N_20031);
or U20720 (N_20720,N_20315,N_19897);
and U20721 (N_20721,N_19909,N_20205);
and U20722 (N_20722,N_19863,N_20073);
nand U20723 (N_20723,N_20161,N_20154);
nand U20724 (N_20724,N_20297,N_20145);
nor U20725 (N_20725,N_20178,N_20096);
nand U20726 (N_20726,N_20209,N_19916);
nor U20727 (N_20727,N_20193,N_19906);
nor U20728 (N_20728,N_19835,N_20128);
nor U20729 (N_20729,N_20258,N_20282);
nand U20730 (N_20730,N_20096,N_19918);
and U20731 (N_20731,N_20333,N_20062);
nor U20732 (N_20732,N_19959,N_19950);
or U20733 (N_20733,N_20031,N_19825);
xnor U20734 (N_20734,N_20000,N_20041);
xnor U20735 (N_20735,N_20184,N_20106);
xnor U20736 (N_20736,N_20226,N_20097);
nor U20737 (N_20737,N_19863,N_20198);
nand U20738 (N_20738,N_20233,N_20358);
xnor U20739 (N_20739,N_20328,N_20196);
nand U20740 (N_20740,N_20336,N_20268);
xor U20741 (N_20741,N_20060,N_20203);
nand U20742 (N_20742,N_19873,N_20197);
xnor U20743 (N_20743,N_20230,N_20125);
or U20744 (N_20744,N_20272,N_19974);
or U20745 (N_20745,N_20285,N_19828);
nor U20746 (N_20746,N_19985,N_20283);
nand U20747 (N_20747,N_20254,N_20271);
nor U20748 (N_20748,N_20277,N_20023);
xnor U20749 (N_20749,N_20276,N_20060);
nor U20750 (N_20750,N_20262,N_20146);
or U20751 (N_20751,N_20253,N_20094);
or U20752 (N_20752,N_19976,N_19993);
nand U20753 (N_20753,N_19880,N_20136);
or U20754 (N_20754,N_19938,N_20081);
nand U20755 (N_20755,N_20230,N_20274);
and U20756 (N_20756,N_19928,N_19991);
xor U20757 (N_20757,N_20081,N_19897);
nor U20758 (N_20758,N_19890,N_19881);
and U20759 (N_20759,N_19824,N_20118);
xor U20760 (N_20760,N_20399,N_19807);
and U20761 (N_20761,N_19909,N_19820);
nand U20762 (N_20762,N_20140,N_20248);
or U20763 (N_20763,N_20260,N_19994);
and U20764 (N_20764,N_20046,N_20064);
xor U20765 (N_20765,N_19842,N_20053);
nand U20766 (N_20766,N_20313,N_20168);
or U20767 (N_20767,N_19917,N_20269);
and U20768 (N_20768,N_20157,N_19969);
xnor U20769 (N_20769,N_19879,N_19957);
nor U20770 (N_20770,N_20330,N_20118);
and U20771 (N_20771,N_20040,N_19842);
and U20772 (N_20772,N_20385,N_20180);
or U20773 (N_20773,N_20124,N_19810);
nor U20774 (N_20774,N_19998,N_20391);
nor U20775 (N_20775,N_20252,N_19952);
nand U20776 (N_20776,N_19979,N_19914);
nor U20777 (N_20777,N_19837,N_19859);
or U20778 (N_20778,N_20361,N_20253);
xnor U20779 (N_20779,N_20278,N_20353);
xor U20780 (N_20780,N_19965,N_20283);
and U20781 (N_20781,N_20135,N_20030);
or U20782 (N_20782,N_20393,N_20337);
and U20783 (N_20783,N_19936,N_20205);
nand U20784 (N_20784,N_20038,N_20217);
nor U20785 (N_20785,N_20365,N_20185);
or U20786 (N_20786,N_19972,N_20215);
nand U20787 (N_20787,N_20307,N_20145);
or U20788 (N_20788,N_20190,N_20077);
nand U20789 (N_20789,N_20080,N_20226);
nor U20790 (N_20790,N_20178,N_20377);
xor U20791 (N_20791,N_20068,N_19965);
or U20792 (N_20792,N_20399,N_20205);
or U20793 (N_20793,N_19941,N_20239);
and U20794 (N_20794,N_20105,N_20249);
nand U20795 (N_20795,N_20220,N_20208);
and U20796 (N_20796,N_20264,N_19969);
nand U20797 (N_20797,N_20350,N_19868);
nor U20798 (N_20798,N_20398,N_19972);
xnor U20799 (N_20799,N_20262,N_20301);
nor U20800 (N_20800,N_20259,N_20047);
or U20801 (N_20801,N_20137,N_19899);
and U20802 (N_20802,N_20087,N_20228);
nand U20803 (N_20803,N_19852,N_19978);
nor U20804 (N_20804,N_20069,N_20150);
or U20805 (N_20805,N_19810,N_20267);
nor U20806 (N_20806,N_19865,N_19808);
nand U20807 (N_20807,N_19822,N_20330);
nand U20808 (N_20808,N_20217,N_19989);
nor U20809 (N_20809,N_20214,N_20043);
or U20810 (N_20810,N_20126,N_19992);
and U20811 (N_20811,N_20254,N_20319);
nand U20812 (N_20812,N_19922,N_20390);
and U20813 (N_20813,N_20060,N_20010);
and U20814 (N_20814,N_19855,N_20275);
nor U20815 (N_20815,N_20064,N_20347);
and U20816 (N_20816,N_19887,N_20151);
nor U20817 (N_20817,N_20320,N_19828);
and U20818 (N_20818,N_19881,N_20346);
xnor U20819 (N_20819,N_19832,N_19802);
xor U20820 (N_20820,N_20305,N_19842);
or U20821 (N_20821,N_20152,N_20325);
and U20822 (N_20822,N_20359,N_19813);
xnor U20823 (N_20823,N_20237,N_20372);
or U20824 (N_20824,N_20386,N_20092);
xor U20825 (N_20825,N_20258,N_20063);
and U20826 (N_20826,N_19922,N_20288);
nor U20827 (N_20827,N_20201,N_20061);
xnor U20828 (N_20828,N_20194,N_20142);
nand U20829 (N_20829,N_20041,N_20022);
xor U20830 (N_20830,N_19872,N_19852);
nor U20831 (N_20831,N_20268,N_19973);
or U20832 (N_20832,N_20292,N_20153);
and U20833 (N_20833,N_19828,N_20257);
and U20834 (N_20834,N_20352,N_20022);
nand U20835 (N_20835,N_20228,N_20390);
nor U20836 (N_20836,N_20235,N_19940);
nor U20837 (N_20837,N_19811,N_20283);
xnor U20838 (N_20838,N_20205,N_19896);
or U20839 (N_20839,N_20248,N_20024);
and U20840 (N_20840,N_20368,N_20263);
nand U20841 (N_20841,N_20327,N_20300);
xor U20842 (N_20842,N_20365,N_20044);
nand U20843 (N_20843,N_20118,N_19961);
xor U20844 (N_20844,N_20127,N_19842);
and U20845 (N_20845,N_20008,N_20233);
and U20846 (N_20846,N_20290,N_19920);
and U20847 (N_20847,N_20390,N_20062);
nor U20848 (N_20848,N_19946,N_20192);
or U20849 (N_20849,N_19870,N_20164);
xnor U20850 (N_20850,N_19833,N_19930);
nand U20851 (N_20851,N_19832,N_19923);
or U20852 (N_20852,N_20227,N_20321);
xor U20853 (N_20853,N_20232,N_20135);
or U20854 (N_20854,N_20000,N_20004);
nand U20855 (N_20855,N_20214,N_20187);
and U20856 (N_20856,N_20166,N_20185);
nor U20857 (N_20857,N_20175,N_19975);
xor U20858 (N_20858,N_20388,N_19827);
and U20859 (N_20859,N_19980,N_19835);
and U20860 (N_20860,N_19979,N_20367);
xor U20861 (N_20861,N_19815,N_20197);
nor U20862 (N_20862,N_20025,N_20339);
or U20863 (N_20863,N_20115,N_20122);
nand U20864 (N_20864,N_19998,N_19926);
nand U20865 (N_20865,N_19916,N_20158);
nand U20866 (N_20866,N_20384,N_20092);
and U20867 (N_20867,N_19903,N_20185);
or U20868 (N_20868,N_19887,N_20140);
xor U20869 (N_20869,N_19922,N_20082);
nor U20870 (N_20870,N_20018,N_20021);
and U20871 (N_20871,N_20021,N_20094);
xnor U20872 (N_20872,N_20329,N_19881);
xor U20873 (N_20873,N_19978,N_19844);
or U20874 (N_20874,N_19842,N_19824);
and U20875 (N_20875,N_19966,N_19886);
or U20876 (N_20876,N_19846,N_19999);
xnor U20877 (N_20877,N_19921,N_20357);
nand U20878 (N_20878,N_20047,N_19950);
nand U20879 (N_20879,N_20354,N_20053);
nor U20880 (N_20880,N_19898,N_20114);
xor U20881 (N_20881,N_20076,N_19951);
or U20882 (N_20882,N_20215,N_19994);
xor U20883 (N_20883,N_20277,N_20305);
nor U20884 (N_20884,N_20004,N_19882);
or U20885 (N_20885,N_20028,N_19813);
or U20886 (N_20886,N_19868,N_19953);
nor U20887 (N_20887,N_20317,N_19984);
and U20888 (N_20888,N_20028,N_19833);
nor U20889 (N_20889,N_19984,N_20218);
nand U20890 (N_20890,N_19834,N_20070);
nor U20891 (N_20891,N_20180,N_20102);
xor U20892 (N_20892,N_19975,N_19806);
and U20893 (N_20893,N_19906,N_20328);
nor U20894 (N_20894,N_19833,N_19838);
and U20895 (N_20895,N_20334,N_20194);
or U20896 (N_20896,N_20035,N_20363);
xnor U20897 (N_20897,N_20337,N_19875);
and U20898 (N_20898,N_20160,N_19850);
or U20899 (N_20899,N_20075,N_20178);
nor U20900 (N_20900,N_20040,N_20144);
or U20901 (N_20901,N_20048,N_19928);
nor U20902 (N_20902,N_20170,N_19942);
xor U20903 (N_20903,N_19961,N_19861);
and U20904 (N_20904,N_19980,N_19970);
and U20905 (N_20905,N_20372,N_20066);
and U20906 (N_20906,N_19916,N_20352);
nand U20907 (N_20907,N_20347,N_20166);
and U20908 (N_20908,N_19896,N_19959);
and U20909 (N_20909,N_20219,N_20267);
and U20910 (N_20910,N_20088,N_19843);
nand U20911 (N_20911,N_20199,N_20303);
xor U20912 (N_20912,N_20148,N_20340);
or U20913 (N_20913,N_19982,N_19917);
xnor U20914 (N_20914,N_20229,N_19836);
nand U20915 (N_20915,N_20319,N_19844);
xnor U20916 (N_20916,N_20045,N_20390);
nor U20917 (N_20917,N_20300,N_20251);
xnor U20918 (N_20918,N_20327,N_20165);
xor U20919 (N_20919,N_19925,N_20136);
nor U20920 (N_20920,N_20201,N_19855);
and U20921 (N_20921,N_19922,N_20231);
and U20922 (N_20922,N_20359,N_20199);
or U20923 (N_20923,N_19890,N_20286);
nand U20924 (N_20924,N_20069,N_20352);
nand U20925 (N_20925,N_19879,N_19979);
or U20926 (N_20926,N_19991,N_19923);
or U20927 (N_20927,N_20243,N_19947);
or U20928 (N_20928,N_20157,N_20129);
or U20929 (N_20929,N_19808,N_20179);
and U20930 (N_20930,N_20276,N_20050);
or U20931 (N_20931,N_19812,N_20184);
nor U20932 (N_20932,N_20167,N_20003);
and U20933 (N_20933,N_20117,N_20100);
or U20934 (N_20934,N_20218,N_20043);
nand U20935 (N_20935,N_20020,N_19925);
xor U20936 (N_20936,N_19839,N_19985);
nand U20937 (N_20937,N_19988,N_20285);
nor U20938 (N_20938,N_20295,N_19833);
and U20939 (N_20939,N_20053,N_20002);
nand U20940 (N_20940,N_20296,N_19954);
or U20941 (N_20941,N_20282,N_19969);
or U20942 (N_20942,N_20280,N_20398);
nor U20943 (N_20943,N_19828,N_20077);
or U20944 (N_20944,N_20098,N_19950);
and U20945 (N_20945,N_20279,N_20375);
nand U20946 (N_20946,N_19858,N_20291);
or U20947 (N_20947,N_20297,N_19949);
and U20948 (N_20948,N_20087,N_20280);
xor U20949 (N_20949,N_19950,N_20040);
or U20950 (N_20950,N_20399,N_20166);
xnor U20951 (N_20951,N_19886,N_20210);
xor U20952 (N_20952,N_19814,N_20127);
nand U20953 (N_20953,N_20317,N_20171);
nor U20954 (N_20954,N_19924,N_19986);
nor U20955 (N_20955,N_20330,N_19980);
or U20956 (N_20956,N_20141,N_20089);
xor U20957 (N_20957,N_20339,N_20066);
xnor U20958 (N_20958,N_19878,N_20177);
nor U20959 (N_20959,N_19918,N_20227);
and U20960 (N_20960,N_19999,N_19989);
nand U20961 (N_20961,N_20108,N_19872);
xnor U20962 (N_20962,N_19919,N_20025);
nor U20963 (N_20963,N_20353,N_19912);
or U20964 (N_20964,N_20310,N_20087);
xor U20965 (N_20965,N_20103,N_20372);
nor U20966 (N_20966,N_20074,N_20323);
nand U20967 (N_20967,N_20327,N_20040);
or U20968 (N_20968,N_20192,N_19874);
nor U20969 (N_20969,N_20149,N_19992);
xor U20970 (N_20970,N_20079,N_19953);
or U20971 (N_20971,N_20349,N_20253);
or U20972 (N_20972,N_19991,N_19959);
nand U20973 (N_20973,N_20317,N_20013);
xor U20974 (N_20974,N_19805,N_20023);
and U20975 (N_20975,N_19852,N_19993);
xnor U20976 (N_20976,N_19818,N_20362);
or U20977 (N_20977,N_20035,N_19939);
nor U20978 (N_20978,N_20238,N_20322);
xnor U20979 (N_20979,N_20309,N_19924);
nand U20980 (N_20980,N_20252,N_20017);
nand U20981 (N_20981,N_20365,N_19945);
nand U20982 (N_20982,N_20125,N_19836);
xnor U20983 (N_20983,N_20288,N_20143);
or U20984 (N_20984,N_19950,N_20378);
nand U20985 (N_20985,N_19946,N_20356);
or U20986 (N_20986,N_20184,N_20224);
or U20987 (N_20987,N_20305,N_20263);
and U20988 (N_20988,N_20306,N_20304);
nand U20989 (N_20989,N_20278,N_19839);
nor U20990 (N_20990,N_19867,N_19853);
nor U20991 (N_20991,N_19888,N_19839);
or U20992 (N_20992,N_20068,N_19956);
xor U20993 (N_20993,N_20181,N_20308);
and U20994 (N_20994,N_19960,N_20089);
nor U20995 (N_20995,N_19999,N_19960);
xnor U20996 (N_20996,N_20053,N_19892);
nand U20997 (N_20997,N_19916,N_20366);
or U20998 (N_20998,N_19805,N_19969);
or U20999 (N_20999,N_20048,N_20028);
and U21000 (N_21000,N_20817,N_20479);
nand U21001 (N_21001,N_20940,N_20975);
and U21002 (N_21002,N_20816,N_20652);
or U21003 (N_21003,N_20851,N_20427);
or U21004 (N_21004,N_20861,N_20482);
nor U21005 (N_21005,N_20574,N_20932);
nand U21006 (N_21006,N_20468,N_20909);
nor U21007 (N_21007,N_20737,N_20458);
and U21008 (N_21008,N_20442,N_20776);
or U21009 (N_21009,N_20749,N_20533);
or U21010 (N_21010,N_20834,N_20997);
or U21011 (N_21011,N_20467,N_20745);
xor U21012 (N_21012,N_20502,N_20720);
nand U21013 (N_21013,N_20838,N_20684);
xnor U21014 (N_21014,N_20639,N_20735);
and U21015 (N_21015,N_20551,N_20769);
xor U21016 (N_21016,N_20915,N_20724);
or U21017 (N_21017,N_20648,N_20739);
nand U21018 (N_21018,N_20582,N_20653);
and U21019 (N_21019,N_20741,N_20538);
xnor U21020 (N_21020,N_20992,N_20401);
nand U21021 (N_21021,N_20635,N_20417);
nor U21022 (N_21022,N_20564,N_20883);
xnor U21023 (N_21023,N_20733,N_20729);
xnor U21024 (N_21024,N_20498,N_20566);
nand U21025 (N_21025,N_20619,N_20865);
nor U21026 (N_21026,N_20873,N_20785);
xor U21027 (N_21027,N_20811,N_20887);
xnor U21028 (N_21028,N_20919,N_20877);
or U21029 (N_21029,N_20594,N_20882);
xor U21030 (N_21030,N_20476,N_20779);
nand U21031 (N_21031,N_20968,N_20478);
nor U21032 (N_21032,N_20872,N_20899);
nor U21033 (N_21033,N_20957,N_20660);
and U21034 (N_21034,N_20974,N_20777);
nor U21035 (N_21035,N_20444,N_20581);
xor U21036 (N_21036,N_20945,N_20807);
nand U21037 (N_21037,N_20634,N_20470);
xor U21038 (N_21038,N_20876,N_20740);
nor U21039 (N_21039,N_20762,N_20544);
nand U21040 (N_21040,N_20978,N_20512);
xnor U21041 (N_21041,N_20715,N_20840);
nor U21042 (N_21042,N_20774,N_20793);
and U21043 (N_21043,N_20555,N_20404);
nor U21044 (N_21044,N_20893,N_20434);
and U21045 (N_21045,N_20682,N_20505);
xnor U21046 (N_21046,N_20591,N_20493);
nor U21047 (N_21047,N_20959,N_20643);
xnor U21048 (N_21048,N_20681,N_20557);
nand U21049 (N_21049,N_20622,N_20641);
or U21050 (N_21050,N_20875,N_20515);
nor U21051 (N_21051,N_20924,N_20436);
and U21052 (N_21052,N_20925,N_20757);
nand U21053 (N_21053,N_20727,N_20979);
or U21054 (N_21054,N_20723,N_20462);
and U21055 (N_21055,N_20579,N_20441);
or U21056 (N_21056,N_20509,N_20988);
xnor U21057 (N_21057,N_20879,N_20751);
nor U21058 (N_21058,N_20839,N_20633);
xnor U21059 (N_21059,N_20714,N_20438);
nor U21060 (N_21060,N_20513,N_20752);
nand U21061 (N_21061,N_20416,N_20547);
or U21062 (N_21062,N_20411,N_20526);
and U21063 (N_21063,N_20750,N_20954);
nand U21064 (N_21064,N_20991,N_20593);
nor U21065 (N_21065,N_20577,N_20449);
and U21066 (N_21066,N_20772,N_20603);
xor U21067 (N_21067,N_20693,N_20699);
nand U21068 (N_21068,N_20791,N_20420);
and U21069 (N_21069,N_20624,N_20599);
or U21070 (N_21070,N_20530,N_20880);
nand U21071 (N_21071,N_20670,N_20709);
nor U21072 (N_21072,N_20613,N_20783);
nand U21073 (N_21073,N_20580,N_20929);
nand U21074 (N_21074,N_20927,N_20961);
nand U21075 (N_21075,N_20405,N_20952);
xnor U21076 (N_21076,N_20454,N_20632);
nor U21077 (N_21077,N_20523,N_20597);
or U21078 (N_21078,N_20463,N_20894);
nand U21079 (N_21079,N_20758,N_20665);
xnor U21080 (N_21080,N_20431,N_20782);
xor U21081 (N_21081,N_20428,N_20734);
nand U21082 (N_21082,N_20903,N_20548);
or U21083 (N_21083,N_20691,N_20938);
and U21084 (N_21084,N_20743,N_20522);
xnor U21085 (N_21085,N_20521,N_20447);
nand U21086 (N_21086,N_20525,N_20763);
or U21087 (N_21087,N_20799,N_20569);
nor U21088 (N_21088,N_20598,N_20765);
and U21089 (N_21089,N_20540,N_20874);
nor U21090 (N_21090,N_20748,N_20558);
and U21091 (N_21091,N_20747,N_20666);
nand U21092 (N_21092,N_20702,N_20687);
nor U21093 (N_21093,N_20814,N_20920);
or U21094 (N_21094,N_20955,N_20889);
nor U21095 (N_21095,N_20852,N_20946);
xor U21096 (N_21096,N_20725,N_20804);
and U21097 (N_21097,N_20705,N_20820);
nand U21098 (N_21098,N_20456,N_20517);
nor U21099 (N_21099,N_20808,N_20460);
xnor U21100 (N_21100,N_20706,N_20972);
or U21101 (N_21101,N_20833,N_20419);
xor U21102 (N_21102,N_20560,N_20572);
nand U21103 (N_21103,N_20402,N_20756);
or U21104 (N_21104,N_20717,N_20810);
nor U21105 (N_21105,N_20836,N_20649);
nand U21106 (N_21106,N_20996,N_20832);
nor U21107 (N_21107,N_20916,N_20913);
nor U21108 (N_21108,N_20778,N_20964);
nand U21109 (N_21109,N_20688,N_20895);
nor U21110 (N_21110,N_20592,N_20536);
xnor U21111 (N_21111,N_20926,N_20661);
xor U21112 (N_21112,N_20704,N_20918);
and U21113 (N_21113,N_20527,N_20472);
nor U21114 (N_21114,N_20870,N_20931);
nor U21115 (N_21115,N_20999,N_20443);
xor U21116 (N_21116,N_20654,N_20841);
or U21117 (N_21117,N_20892,N_20617);
nor U21118 (N_21118,N_20489,N_20537);
xor U21119 (N_21119,N_20923,N_20673);
and U21120 (N_21120,N_20475,N_20897);
and U21121 (N_21121,N_20503,N_20410);
xor U21122 (N_21122,N_20742,N_20678);
and U21123 (N_21123,N_20949,N_20656);
and U21124 (N_21124,N_20754,N_20849);
nand U21125 (N_21125,N_20484,N_20963);
nor U21126 (N_21126,N_20912,N_20738);
and U21127 (N_21127,N_20831,N_20614);
xnor U21128 (N_21128,N_20878,N_20828);
and U21129 (N_21129,N_20917,N_20668);
nor U21130 (N_21130,N_20939,N_20432);
nor U21131 (N_21131,N_20866,N_20983);
and U21132 (N_21132,N_20708,N_20585);
nand U21133 (N_21133,N_20590,N_20696);
or U21134 (N_21134,N_20473,N_20461);
or U21135 (N_21135,N_20822,N_20848);
or U21136 (N_21136,N_20575,N_20971);
xor U21137 (N_21137,N_20570,N_20636);
or U21138 (N_21138,N_20455,N_20850);
nor U21139 (N_21139,N_20768,N_20736);
or U21140 (N_21140,N_20845,N_20824);
nor U21141 (N_21141,N_20995,N_20683);
nand U21142 (N_21142,N_20511,N_20821);
nand U21143 (N_21143,N_20935,N_20722);
nand U21144 (N_21144,N_20960,N_20657);
nor U21145 (N_21145,N_20584,N_20623);
xor U21146 (N_21146,N_20885,N_20519);
xor U21147 (N_21147,N_20697,N_20900);
nor U21148 (N_21148,N_20773,N_20695);
or U21149 (N_21149,N_20825,N_20890);
nor U21150 (N_21150,N_20781,N_20869);
and U21151 (N_21151,N_20707,N_20789);
nor U21152 (N_21152,N_20914,N_20437);
and U21153 (N_21153,N_20507,N_20625);
xor U21154 (N_21154,N_20989,N_20790);
nand U21155 (N_21155,N_20618,N_20408);
xnor U21156 (N_21156,N_20847,N_20962);
or U21157 (N_21157,N_20674,N_20846);
nand U21158 (N_21158,N_20440,N_20888);
nor U21159 (N_21159,N_20567,N_20761);
xnor U21160 (N_21160,N_20857,N_20647);
or U21161 (N_21161,N_20541,N_20694);
nor U21162 (N_21162,N_20986,N_20837);
nand U21163 (N_21163,N_20587,N_20703);
nor U21164 (N_21164,N_20471,N_20545);
nor U21165 (N_21165,N_20504,N_20520);
xor U21166 (N_21166,N_20528,N_20531);
xor U21167 (N_21167,N_20928,N_20944);
and U21168 (N_21168,N_20711,N_20835);
nand U21169 (N_21169,N_20413,N_20800);
and U21170 (N_21170,N_20562,N_20829);
nor U21171 (N_21171,N_20607,N_20630);
nand U21172 (N_21172,N_20445,N_20794);
nand U21173 (N_21173,N_20514,N_20775);
and U21174 (N_21174,N_20856,N_20990);
xnor U21175 (N_21175,N_20430,N_20423);
nand U21176 (N_21176,N_20677,N_20898);
and U21177 (N_21177,N_20539,N_20663);
xor U21178 (N_21178,N_20422,N_20561);
nor U21179 (N_21179,N_20801,N_20465);
nand U21180 (N_21180,N_20549,N_20981);
nand U21181 (N_21181,N_20881,N_20780);
or U21182 (N_21182,N_20638,N_20951);
nand U21183 (N_21183,N_20662,N_20669);
nand U21184 (N_21184,N_20412,N_20956);
xnor U21185 (N_21185,N_20759,N_20676);
and U21186 (N_21186,N_20842,N_20813);
or U21187 (N_21187,N_20942,N_20604);
nor U21188 (N_21188,N_20469,N_20867);
xor U21189 (N_21189,N_20589,N_20586);
nand U21190 (N_21190,N_20609,N_20483);
and U21191 (N_21191,N_20980,N_20506);
and U21192 (N_21192,N_20690,N_20601);
nor U21193 (N_21193,N_20994,N_20855);
xnor U21194 (N_21194,N_20933,N_20910);
xnor U21195 (N_21195,N_20965,N_20823);
xor U21196 (N_21196,N_20853,N_20966);
nor U21197 (N_21197,N_20796,N_20827);
nand U21198 (N_21198,N_20770,N_20862);
or U21199 (N_21199,N_20786,N_20803);
or U21200 (N_21200,N_20516,N_20474);
and U21201 (N_21201,N_20680,N_20744);
xnor U21202 (N_21202,N_20921,N_20767);
nor U21203 (N_21203,N_20843,N_20985);
nor U21204 (N_21204,N_20610,N_20631);
nand U21205 (N_21205,N_20415,N_20712);
or U21206 (N_21206,N_20911,N_20930);
or U21207 (N_21207,N_20616,N_20795);
nand U21208 (N_21208,N_20701,N_20446);
xor U21209 (N_21209,N_20611,N_20760);
nand U21210 (N_21210,N_20859,N_20886);
xnor U21211 (N_21211,N_20571,N_20730);
or U21212 (N_21212,N_20937,N_20941);
xnor U21213 (N_21213,N_20675,N_20495);
and U21214 (N_21214,N_20439,N_20508);
nand U21215 (N_21215,N_20409,N_20578);
or U21216 (N_21216,N_20435,N_20573);
or U21217 (N_21217,N_20424,N_20896);
and U21218 (N_21218,N_20984,N_20826);
and U21219 (N_21219,N_20922,N_20732);
xor U21220 (N_21220,N_20595,N_20969);
and U21221 (N_21221,N_20477,N_20559);
nor U21222 (N_21222,N_20637,N_20906);
nor U21223 (N_21223,N_20970,N_20629);
or U21224 (N_21224,N_20905,N_20426);
or U21225 (N_21225,N_20973,N_20976);
nor U21226 (N_21226,N_20486,N_20863);
and U21227 (N_21227,N_20407,N_20884);
and U21228 (N_21228,N_20491,N_20908);
nor U21229 (N_21229,N_20858,N_20550);
or U21230 (N_21230,N_20543,N_20788);
and U21231 (N_21231,N_20953,N_20907);
and U21232 (N_21232,N_20644,N_20766);
and U21233 (N_21233,N_20689,N_20612);
nand U21234 (N_21234,N_20692,N_20819);
nor U21235 (N_21235,N_20718,N_20452);
and U21236 (N_21236,N_20967,N_20406);
xnor U21237 (N_21237,N_20868,N_20605);
and U21238 (N_21238,N_20998,N_20554);
and U21239 (N_21239,N_20529,N_20686);
or U21240 (N_21240,N_20563,N_20429);
nand U21241 (N_21241,N_20494,N_20400);
nand U21242 (N_21242,N_20787,N_20993);
nand U21243 (N_21243,N_20698,N_20719);
and U21244 (N_21244,N_20792,N_20710);
and U21245 (N_21245,N_20628,N_20606);
nand U21246 (N_21246,N_20421,N_20642);
xnor U21247 (N_21247,N_20453,N_20726);
and U21248 (N_21248,N_20576,N_20844);
and U21249 (N_21249,N_20871,N_20977);
nand U21250 (N_21250,N_20546,N_20679);
and U21251 (N_21251,N_20450,N_20501);
or U21252 (N_21252,N_20934,N_20685);
xnor U21253 (N_21253,N_20602,N_20830);
and U21254 (N_21254,N_20556,N_20403);
xnor U21255 (N_21255,N_20818,N_20466);
and U21256 (N_21256,N_20812,N_20626);
xor U21257 (N_21257,N_20753,N_20518);
and U21258 (N_21258,N_20542,N_20565);
nand U21259 (N_21259,N_20457,N_20568);
xnor U21260 (N_21260,N_20596,N_20784);
or U21261 (N_21261,N_20487,N_20721);
xor U21262 (N_21262,N_20448,N_20904);
nand U21263 (N_21263,N_20815,N_20948);
and U21264 (N_21264,N_20433,N_20553);
nor U21265 (N_21265,N_20987,N_20651);
nand U21266 (N_21266,N_20608,N_20510);
nand U21267 (N_21267,N_20659,N_20620);
nor U21268 (N_21268,N_20667,N_20615);
xnor U21269 (N_21269,N_20499,N_20672);
or U21270 (N_21270,N_20860,N_20583);
and U21271 (N_21271,N_20764,N_20459);
and U21272 (N_21272,N_20524,N_20809);
and U21273 (N_21273,N_20535,N_20600);
nand U21274 (N_21274,N_20947,N_20731);
nor U21275 (N_21275,N_20490,N_20798);
xnor U21276 (N_21276,N_20664,N_20902);
nand U21277 (N_21277,N_20728,N_20418);
nor U21278 (N_21278,N_20713,N_20797);
nor U21279 (N_21279,N_20500,N_20534);
xor U21280 (N_21280,N_20805,N_20943);
and U21281 (N_21281,N_20532,N_20982);
nand U21282 (N_21282,N_20627,N_20755);
or U21283 (N_21283,N_20646,N_20806);
nor U21284 (N_21284,N_20671,N_20650);
nor U21285 (N_21285,N_20802,N_20640);
nor U21286 (N_21286,N_20655,N_20936);
and U21287 (N_21287,N_20716,N_20891);
and U21288 (N_21288,N_20485,N_20854);
and U21289 (N_21289,N_20700,N_20958);
xnor U21290 (N_21290,N_20746,N_20658);
nor U21291 (N_21291,N_20864,N_20451);
or U21292 (N_21292,N_20496,N_20414);
nor U21293 (N_21293,N_20901,N_20425);
nand U21294 (N_21294,N_20480,N_20645);
nor U21295 (N_21295,N_20481,N_20552);
or U21296 (N_21296,N_20497,N_20950);
nand U21297 (N_21297,N_20621,N_20588);
or U21298 (N_21298,N_20492,N_20771);
or U21299 (N_21299,N_20488,N_20464);
xnor U21300 (N_21300,N_20424,N_20420);
or U21301 (N_21301,N_20784,N_20805);
and U21302 (N_21302,N_20791,N_20732);
xnor U21303 (N_21303,N_20405,N_20811);
xnor U21304 (N_21304,N_20848,N_20482);
nor U21305 (N_21305,N_20960,N_20405);
nand U21306 (N_21306,N_20644,N_20842);
nand U21307 (N_21307,N_20544,N_20464);
xor U21308 (N_21308,N_20682,N_20496);
xor U21309 (N_21309,N_20903,N_20465);
xor U21310 (N_21310,N_20877,N_20862);
xnor U21311 (N_21311,N_20846,N_20504);
nand U21312 (N_21312,N_20602,N_20536);
and U21313 (N_21313,N_20899,N_20468);
xnor U21314 (N_21314,N_20420,N_20461);
or U21315 (N_21315,N_20893,N_20941);
and U21316 (N_21316,N_20626,N_20765);
nor U21317 (N_21317,N_20663,N_20414);
nor U21318 (N_21318,N_20782,N_20426);
and U21319 (N_21319,N_20702,N_20731);
nand U21320 (N_21320,N_20657,N_20513);
nor U21321 (N_21321,N_20723,N_20985);
nand U21322 (N_21322,N_20631,N_20510);
nand U21323 (N_21323,N_20937,N_20879);
nand U21324 (N_21324,N_20419,N_20498);
or U21325 (N_21325,N_20482,N_20789);
nand U21326 (N_21326,N_20807,N_20735);
nand U21327 (N_21327,N_20707,N_20608);
nor U21328 (N_21328,N_20930,N_20661);
nor U21329 (N_21329,N_20443,N_20607);
xor U21330 (N_21330,N_20879,N_20596);
and U21331 (N_21331,N_20412,N_20683);
and U21332 (N_21332,N_20459,N_20593);
nor U21333 (N_21333,N_20932,N_20725);
or U21334 (N_21334,N_20853,N_20659);
xnor U21335 (N_21335,N_20803,N_20520);
nor U21336 (N_21336,N_20517,N_20927);
or U21337 (N_21337,N_20663,N_20823);
nor U21338 (N_21338,N_20846,N_20939);
and U21339 (N_21339,N_20432,N_20614);
or U21340 (N_21340,N_20860,N_20674);
or U21341 (N_21341,N_20423,N_20556);
and U21342 (N_21342,N_20465,N_20497);
nor U21343 (N_21343,N_20521,N_20788);
nor U21344 (N_21344,N_20951,N_20471);
nor U21345 (N_21345,N_20597,N_20475);
nand U21346 (N_21346,N_20876,N_20989);
nor U21347 (N_21347,N_20496,N_20963);
nand U21348 (N_21348,N_20647,N_20954);
nand U21349 (N_21349,N_20899,N_20592);
xnor U21350 (N_21350,N_20861,N_20442);
nand U21351 (N_21351,N_20541,N_20963);
and U21352 (N_21352,N_20429,N_20897);
nor U21353 (N_21353,N_20485,N_20633);
or U21354 (N_21354,N_20935,N_20423);
xor U21355 (N_21355,N_20517,N_20597);
and U21356 (N_21356,N_20674,N_20565);
xnor U21357 (N_21357,N_20578,N_20609);
nand U21358 (N_21358,N_20570,N_20836);
or U21359 (N_21359,N_20856,N_20554);
nand U21360 (N_21360,N_20658,N_20733);
or U21361 (N_21361,N_20438,N_20868);
nor U21362 (N_21362,N_20600,N_20881);
xor U21363 (N_21363,N_20873,N_20651);
nand U21364 (N_21364,N_20404,N_20525);
nand U21365 (N_21365,N_20489,N_20541);
nor U21366 (N_21366,N_20608,N_20850);
and U21367 (N_21367,N_20829,N_20685);
and U21368 (N_21368,N_20761,N_20609);
and U21369 (N_21369,N_20435,N_20525);
xor U21370 (N_21370,N_20700,N_20875);
and U21371 (N_21371,N_20662,N_20575);
or U21372 (N_21372,N_20467,N_20439);
or U21373 (N_21373,N_20730,N_20451);
nand U21374 (N_21374,N_20478,N_20658);
nor U21375 (N_21375,N_20674,N_20414);
nand U21376 (N_21376,N_20516,N_20800);
or U21377 (N_21377,N_20635,N_20969);
or U21378 (N_21378,N_20735,N_20979);
nand U21379 (N_21379,N_20462,N_20858);
nand U21380 (N_21380,N_20729,N_20460);
and U21381 (N_21381,N_20716,N_20469);
and U21382 (N_21382,N_20821,N_20901);
and U21383 (N_21383,N_20945,N_20775);
or U21384 (N_21384,N_20851,N_20799);
nand U21385 (N_21385,N_20806,N_20826);
nor U21386 (N_21386,N_20847,N_20840);
and U21387 (N_21387,N_20514,N_20497);
or U21388 (N_21388,N_20447,N_20564);
or U21389 (N_21389,N_20984,N_20993);
or U21390 (N_21390,N_20517,N_20905);
and U21391 (N_21391,N_20892,N_20638);
and U21392 (N_21392,N_20820,N_20781);
or U21393 (N_21393,N_20513,N_20674);
nand U21394 (N_21394,N_20551,N_20633);
and U21395 (N_21395,N_20483,N_20903);
or U21396 (N_21396,N_20838,N_20948);
xnor U21397 (N_21397,N_20509,N_20712);
nand U21398 (N_21398,N_20536,N_20917);
or U21399 (N_21399,N_20556,N_20733);
nor U21400 (N_21400,N_20947,N_20586);
and U21401 (N_21401,N_20596,N_20954);
nand U21402 (N_21402,N_20508,N_20702);
nand U21403 (N_21403,N_20569,N_20653);
or U21404 (N_21404,N_20446,N_20811);
xnor U21405 (N_21405,N_20940,N_20468);
and U21406 (N_21406,N_20845,N_20631);
nor U21407 (N_21407,N_20524,N_20864);
nand U21408 (N_21408,N_20920,N_20832);
xnor U21409 (N_21409,N_20629,N_20994);
nand U21410 (N_21410,N_20738,N_20881);
nand U21411 (N_21411,N_20570,N_20972);
nor U21412 (N_21412,N_20780,N_20591);
or U21413 (N_21413,N_20432,N_20519);
nand U21414 (N_21414,N_20473,N_20403);
nand U21415 (N_21415,N_20441,N_20891);
or U21416 (N_21416,N_20933,N_20459);
nor U21417 (N_21417,N_20499,N_20934);
nand U21418 (N_21418,N_20804,N_20947);
xor U21419 (N_21419,N_20456,N_20743);
or U21420 (N_21420,N_20823,N_20791);
nor U21421 (N_21421,N_20673,N_20516);
xnor U21422 (N_21422,N_20560,N_20999);
and U21423 (N_21423,N_20465,N_20850);
and U21424 (N_21424,N_20848,N_20965);
nand U21425 (N_21425,N_20936,N_20983);
or U21426 (N_21426,N_20884,N_20820);
nand U21427 (N_21427,N_20734,N_20522);
nor U21428 (N_21428,N_20907,N_20719);
or U21429 (N_21429,N_20946,N_20428);
xnor U21430 (N_21430,N_20596,N_20708);
and U21431 (N_21431,N_20990,N_20883);
nand U21432 (N_21432,N_20734,N_20545);
nor U21433 (N_21433,N_20637,N_20802);
and U21434 (N_21434,N_20924,N_20619);
and U21435 (N_21435,N_20473,N_20525);
nor U21436 (N_21436,N_20863,N_20555);
nand U21437 (N_21437,N_20500,N_20444);
xnor U21438 (N_21438,N_20988,N_20797);
nor U21439 (N_21439,N_20970,N_20468);
or U21440 (N_21440,N_20900,N_20969);
and U21441 (N_21441,N_20670,N_20968);
or U21442 (N_21442,N_20955,N_20574);
nor U21443 (N_21443,N_20423,N_20636);
and U21444 (N_21444,N_20761,N_20827);
and U21445 (N_21445,N_20896,N_20997);
nor U21446 (N_21446,N_20561,N_20835);
nor U21447 (N_21447,N_20431,N_20781);
or U21448 (N_21448,N_20444,N_20973);
nor U21449 (N_21449,N_20951,N_20838);
nor U21450 (N_21450,N_20563,N_20643);
nor U21451 (N_21451,N_20703,N_20503);
and U21452 (N_21452,N_20475,N_20777);
or U21453 (N_21453,N_20827,N_20786);
and U21454 (N_21454,N_20755,N_20956);
nand U21455 (N_21455,N_20499,N_20948);
xnor U21456 (N_21456,N_20407,N_20445);
xnor U21457 (N_21457,N_20762,N_20931);
nand U21458 (N_21458,N_20563,N_20879);
nand U21459 (N_21459,N_20854,N_20813);
and U21460 (N_21460,N_20742,N_20676);
nor U21461 (N_21461,N_20880,N_20420);
or U21462 (N_21462,N_20820,N_20740);
xor U21463 (N_21463,N_20413,N_20734);
and U21464 (N_21464,N_20693,N_20794);
and U21465 (N_21465,N_20910,N_20483);
and U21466 (N_21466,N_20955,N_20529);
nor U21467 (N_21467,N_20962,N_20787);
nor U21468 (N_21468,N_20621,N_20517);
and U21469 (N_21469,N_20935,N_20626);
or U21470 (N_21470,N_20789,N_20647);
nand U21471 (N_21471,N_20685,N_20924);
nor U21472 (N_21472,N_20822,N_20416);
or U21473 (N_21473,N_20404,N_20701);
xnor U21474 (N_21474,N_20433,N_20789);
nand U21475 (N_21475,N_20981,N_20628);
or U21476 (N_21476,N_20599,N_20835);
and U21477 (N_21477,N_20829,N_20775);
and U21478 (N_21478,N_20438,N_20841);
or U21479 (N_21479,N_20422,N_20920);
and U21480 (N_21480,N_20453,N_20732);
xor U21481 (N_21481,N_20478,N_20981);
nor U21482 (N_21482,N_20524,N_20852);
and U21483 (N_21483,N_20611,N_20788);
and U21484 (N_21484,N_20937,N_20424);
nor U21485 (N_21485,N_20818,N_20984);
or U21486 (N_21486,N_20679,N_20575);
nor U21487 (N_21487,N_20434,N_20623);
and U21488 (N_21488,N_20419,N_20735);
nand U21489 (N_21489,N_20972,N_20843);
and U21490 (N_21490,N_20880,N_20691);
nor U21491 (N_21491,N_20813,N_20457);
nand U21492 (N_21492,N_20973,N_20721);
nor U21493 (N_21493,N_20634,N_20449);
and U21494 (N_21494,N_20945,N_20938);
and U21495 (N_21495,N_20787,N_20640);
nor U21496 (N_21496,N_20981,N_20591);
and U21497 (N_21497,N_20473,N_20898);
and U21498 (N_21498,N_20658,N_20639);
nand U21499 (N_21499,N_20567,N_20446);
xor U21500 (N_21500,N_20936,N_20452);
or U21501 (N_21501,N_20401,N_20911);
nor U21502 (N_21502,N_20515,N_20761);
or U21503 (N_21503,N_20918,N_20550);
and U21504 (N_21504,N_20619,N_20585);
and U21505 (N_21505,N_20671,N_20825);
nand U21506 (N_21506,N_20801,N_20500);
or U21507 (N_21507,N_20640,N_20808);
xor U21508 (N_21508,N_20679,N_20641);
or U21509 (N_21509,N_20890,N_20701);
nand U21510 (N_21510,N_20557,N_20928);
or U21511 (N_21511,N_20562,N_20612);
nand U21512 (N_21512,N_20770,N_20646);
and U21513 (N_21513,N_20412,N_20847);
nand U21514 (N_21514,N_20632,N_20971);
nand U21515 (N_21515,N_20443,N_20853);
and U21516 (N_21516,N_20960,N_20600);
nand U21517 (N_21517,N_20879,N_20542);
xor U21518 (N_21518,N_20845,N_20453);
nand U21519 (N_21519,N_20427,N_20422);
and U21520 (N_21520,N_20855,N_20876);
xnor U21521 (N_21521,N_20810,N_20968);
or U21522 (N_21522,N_20938,N_20597);
nand U21523 (N_21523,N_20906,N_20699);
or U21524 (N_21524,N_20950,N_20996);
nor U21525 (N_21525,N_20852,N_20792);
nand U21526 (N_21526,N_20946,N_20676);
or U21527 (N_21527,N_20671,N_20922);
and U21528 (N_21528,N_20935,N_20526);
nor U21529 (N_21529,N_20403,N_20412);
xor U21530 (N_21530,N_20953,N_20855);
nor U21531 (N_21531,N_20553,N_20523);
and U21532 (N_21532,N_20605,N_20611);
nand U21533 (N_21533,N_20850,N_20426);
and U21534 (N_21534,N_20875,N_20952);
nand U21535 (N_21535,N_20561,N_20493);
nor U21536 (N_21536,N_20682,N_20830);
nor U21537 (N_21537,N_20773,N_20818);
nand U21538 (N_21538,N_20466,N_20859);
or U21539 (N_21539,N_20867,N_20562);
nand U21540 (N_21540,N_20487,N_20526);
nand U21541 (N_21541,N_20844,N_20803);
xor U21542 (N_21542,N_20612,N_20981);
and U21543 (N_21543,N_20518,N_20801);
xor U21544 (N_21544,N_20888,N_20679);
nand U21545 (N_21545,N_20524,N_20768);
xor U21546 (N_21546,N_20501,N_20532);
or U21547 (N_21547,N_20887,N_20699);
nor U21548 (N_21548,N_20518,N_20456);
nand U21549 (N_21549,N_20714,N_20826);
or U21550 (N_21550,N_20422,N_20768);
xor U21551 (N_21551,N_20840,N_20413);
or U21552 (N_21552,N_20863,N_20476);
and U21553 (N_21553,N_20582,N_20847);
and U21554 (N_21554,N_20561,N_20827);
and U21555 (N_21555,N_20963,N_20809);
nand U21556 (N_21556,N_20861,N_20715);
nand U21557 (N_21557,N_20405,N_20883);
or U21558 (N_21558,N_20828,N_20499);
nor U21559 (N_21559,N_20852,N_20418);
xor U21560 (N_21560,N_20944,N_20674);
nand U21561 (N_21561,N_20480,N_20846);
xnor U21562 (N_21562,N_20937,N_20465);
xnor U21563 (N_21563,N_20730,N_20470);
xor U21564 (N_21564,N_20607,N_20522);
nand U21565 (N_21565,N_20445,N_20916);
nand U21566 (N_21566,N_20484,N_20668);
or U21567 (N_21567,N_20746,N_20689);
nand U21568 (N_21568,N_20691,N_20855);
or U21569 (N_21569,N_20770,N_20736);
and U21570 (N_21570,N_20650,N_20928);
nor U21571 (N_21571,N_20764,N_20930);
nand U21572 (N_21572,N_20507,N_20957);
nand U21573 (N_21573,N_20514,N_20488);
and U21574 (N_21574,N_20430,N_20710);
xnor U21575 (N_21575,N_20420,N_20695);
nor U21576 (N_21576,N_20785,N_20664);
nor U21577 (N_21577,N_20768,N_20845);
nor U21578 (N_21578,N_20702,N_20854);
or U21579 (N_21579,N_20585,N_20832);
nor U21580 (N_21580,N_20702,N_20861);
and U21581 (N_21581,N_20981,N_20924);
or U21582 (N_21582,N_20809,N_20928);
xnor U21583 (N_21583,N_20829,N_20889);
nand U21584 (N_21584,N_20624,N_20738);
nand U21585 (N_21585,N_20770,N_20518);
and U21586 (N_21586,N_20577,N_20432);
nand U21587 (N_21587,N_20903,N_20961);
or U21588 (N_21588,N_20969,N_20640);
xor U21589 (N_21589,N_20736,N_20815);
xor U21590 (N_21590,N_20763,N_20490);
and U21591 (N_21591,N_20452,N_20917);
nand U21592 (N_21592,N_20952,N_20554);
xor U21593 (N_21593,N_20896,N_20609);
and U21594 (N_21594,N_20868,N_20488);
nor U21595 (N_21595,N_20858,N_20545);
or U21596 (N_21596,N_20497,N_20817);
and U21597 (N_21597,N_20719,N_20650);
xor U21598 (N_21598,N_20903,N_20966);
and U21599 (N_21599,N_20531,N_20703);
nand U21600 (N_21600,N_21376,N_21240);
nand U21601 (N_21601,N_21044,N_21232);
xor U21602 (N_21602,N_21496,N_21233);
or U21603 (N_21603,N_21526,N_21024);
and U21604 (N_21604,N_21192,N_21471);
nor U21605 (N_21605,N_21074,N_21482);
nor U21606 (N_21606,N_21151,N_21234);
or U21607 (N_21607,N_21082,N_21011);
xnor U21608 (N_21608,N_21014,N_21253);
nor U21609 (N_21609,N_21002,N_21169);
xnor U21610 (N_21610,N_21041,N_21593);
nor U21611 (N_21611,N_21590,N_21386);
or U21612 (N_21612,N_21182,N_21264);
and U21613 (N_21613,N_21245,N_21358);
nand U21614 (N_21614,N_21200,N_21202);
and U21615 (N_21615,N_21512,N_21267);
nor U21616 (N_21616,N_21388,N_21094);
and U21617 (N_21617,N_21341,N_21039);
nand U21618 (N_21618,N_21059,N_21159);
nand U21619 (N_21619,N_21069,N_21499);
and U21620 (N_21620,N_21438,N_21391);
and U21621 (N_21621,N_21345,N_21133);
nor U21622 (N_21622,N_21140,N_21164);
nor U21623 (N_21623,N_21291,N_21565);
or U21624 (N_21624,N_21516,N_21128);
nand U21625 (N_21625,N_21580,N_21073);
and U21626 (N_21626,N_21405,N_21543);
nor U21627 (N_21627,N_21038,N_21520);
nor U21628 (N_21628,N_21325,N_21181);
or U21629 (N_21629,N_21153,N_21235);
nor U21630 (N_21630,N_21582,N_21329);
nor U21631 (N_21631,N_21449,N_21020);
or U21632 (N_21632,N_21070,N_21150);
or U21633 (N_21633,N_21564,N_21005);
or U21634 (N_21634,N_21408,N_21502);
or U21635 (N_21635,N_21320,N_21436);
nand U21636 (N_21636,N_21442,N_21156);
and U21637 (N_21637,N_21268,N_21367);
or U21638 (N_21638,N_21052,N_21574);
or U21639 (N_21639,N_21224,N_21279);
or U21640 (N_21640,N_21415,N_21229);
xor U21641 (N_21641,N_21148,N_21461);
nand U21642 (N_21642,N_21395,N_21400);
and U21643 (N_21643,N_21101,N_21481);
nor U21644 (N_21644,N_21248,N_21554);
nor U21645 (N_21645,N_21061,N_21570);
and U21646 (N_21646,N_21191,N_21075);
or U21647 (N_21647,N_21326,N_21123);
and U21648 (N_21648,N_21095,N_21484);
nand U21649 (N_21649,N_21406,N_21212);
or U21650 (N_21650,N_21563,N_21403);
nand U21651 (N_21651,N_21342,N_21448);
and U21652 (N_21652,N_21165,N_21237);
xor U21653 (N_21653,N_21042,N_21102);
nand U21654 (N_21654,N_21383,N_21327);
xor U21655 (N_21655,N_21414,N_21284);
nor U21656 (N_21656,N_21349,N_21254);
and U21657 (N_21657,N_21218,N_21596);
and U21658 (N_21658,N_21431,N_21522);
nand U21659 (N_21659,N_21255,N_21302);
nor U21660 (N_21660,N_21258,N_21333);
and U21661 (N_21661,N_21247,N_21033);
or U21662 (N_21662,N_21043,N_21063);
xnor U21663 (N_21663,N_21353,N_21205);
nor U21664 (N_21664,N_21509,N_21010);
nor U21665 (N_21665,N_21385,N_21051);
and U21666 (N_21666,N_21372,N_21135);
nor U21667 (N_21667,N_21357,N_21060);
and U21668 (N_21668,N_21098,N_21534);
or U21669 (N_21669,N_21138,N_21146);
or U21670 (N_21670,N_21226,N_21348);
xnor U21671 (N_21671,N_21071,N_21318);
nor U21672 (N_21672,N_21223,N_21286);
nor U21673 (N_21673,N_21417,N_21167);
xnor U21674 (N_21674,N_21365,N_21027);
xor U21675 (N_21675,N_21242,N_21492);
and U21676 (N_21676,N_21425,N_21505);
nor U21677 (N_21677,N_21132,N_21297);
nand U21678 (N_21678,N_21065,N_21491);
and U21679 (N_21679,N_21572,N_21053);
xnor U21680 (N_21680,N_21322,N_21174);
or U21681 (N_21681,N_21187,N_21315);
nor U21682 (N_21682,N_21531,N_21462);
and U21683 (N_21683,N_21494,N_21422);
nand U21684 (N_21684,N_21289,N_21290);
xnor U21685 (N_21685,N_21556,N_21352);
xor U21686 (N_21686,N_21355,N_21077);
nor U21687 (N_21687,N_21036,N_21394);
xnor U21688 (N_21688,N_21519,N_21466);
or U21689 (N_21689,N_21274,N_21087);
nor U21690 (N_21690,N_21215,N_21547);
or U21691 (N_21691,N_21513,N_21458);
nor U21692 (N_21692,N_21433,N_21524);
and U21693 (N_21693,N_21592,N_21144);
nor U21694 (N_21694,N_21340,N_21006);
xnor U21695 (N_21695,N_21210,N_21529);
xor U21696 (N_21696,N_21149,N_21389);
nor U21697 (N_21697,N_21321,N_21343);
nor U21698 (N_21698,N_21195,N_21504);
xnor U21699 (N_21699,N_21430,N_21113);
nand U21700 (N_21700,N_21402,N_21177);
xor U21701 (N_21701,N_21562,N_21569);
and U21702 (N_21702,N_21147,N_21260);
nor U21703 (N_21703,N_21194,N_21118);
xnor U21704 (N_21704,N_21330,N_21441);
nand U21705 (N_21705,N_21045,N_21050);
nor U21706 (N_21706,N_21239,N_21366);
nand U21707 (N_21707,N_21532,N_21455);
nand U21708 (N_21708,N_21294,N_21595);
xnor U21709 (N_21709,N_21579,N_21546);
nor U21710 (N_21710,N_21567,N_21124);
xor U21711 (N_21711,N_21283,N_21185);
xor U21712 (N_21712,N_21518,N_21324);
nand U21713 (N_21713,N_21080,N_21300);
nand U21714 (N_21714,N_21206,N_21067);
xnor U21715 (N_21715,N_21281,N_21019);
or U21716 (N_21716,N_21046,N_21589);
nor U21717 (N_21717,N_21454,N_21236);
xnor U21718 (N_21718,N_21426,N_21266);
nor U21719 (N_21719,N_21477,N_21464);
nand U21720 (N_21720,N_21549,N_21213);
nor U21721 (N_21721,N_21566,N_21179);
nor U21722 (N_21722,N_21084,N_21017);
nor U21723 (N_21723,N_21419,N_21104);
and U21724 (N_21724,N_21457,N_21062);
and U21725 (N_21725,N_21335,N_21323);
nand U21726 (N_21726,N_21180,N_21064);
and U21727 (N_21727,N_21446,N_21081);
nor U21728 (N_21728,N_21152,N_21575);
nand U21729 (N_21729,N_21251,N_21424);
nor U21730 (N_21730,N_21500,N_21498);
or U21731 (N_21731,N_21557,N_21107);
xor U21732 (N_21732,N_21293,N_21023);
nor U21733 (N_21733,N_21409,N_21263);
xor U21734 (N_21734,N_21571,N_21404);
and U21735 (N_21735,N_21031,N_21003);
xnor U21736 (N_21736,N_21480,N_21004);
nor U21737 (N_21737,N_21009,N_21445);
nand U21738 (N_21738,N_21591,N_21558);
xnor U21739 (N_21739,N_21544,N_21136);
xnor U21740 (N_21740,N_21183,N_21497);
and U21741 (N_21741,N_21028,N_21392);
xor U21742 (N_21742,N_21427,N_21250);
nor U21743 (N_21743,N_21127,N_21256);
nand U21744 (N_21744,N_21598,N_21463);
and U21745 (N_21745,N_21285,N_21338);
xor U21746 (N_21746,N_21550,N_21162);
and U21747 (N_21747,N_21506,N_21114);
nor U21748 (N_21748,N_21129,N_21451);
xnor U21749 (N_21749,N_21271,N_21346);
nor U21750 (N_21750,N_21068,N_21577);
nor U21751 (N_21751,N_21396,N_21022);
or U21752 (N_21752,N_21282,N_21493);
or U21753 (N_21753,N_21334,N_21548);
and U21754 (N_21754,N_21197,N_21539);
and U21755 (N_21755,N_21288,N_21298);
nand U21756 (N_21756,N_21047,N_21198);
nand U21757 (N_21757,N_21261,N_21380);
and U21758 (N_21758,N_21048,N_21468);
nand U21759 (N_21759,N_21597,N_21581);
and U21760 (N_21760,N_21560,N_21190);
nor U21761 (N_21761,N_21021,N_21112);
and U21762 (N_21762,N_21201,N_21120);
or U21763 (N_21763,N_21576,N_21476);
and U21764 (N_21764,N_21428,N_21319);
and U21765 (N_21765,N_21373,N_21211);
and U21766 (N_21766,N_21317,N_21486);
xor U21767 (N_21767,N_21186,N_21533);
nor U21768 (N_21768,N_21407,N_21100);
or U21769 (N_21769,N_21540,N_21573);
nand U21770 (N_21770,N_21176,N_21054);
nor U21771 (N_21771,N_21528,N_21175);
and U21772 (N_21772,N_21125,N_21360);
and U21773 (N_21773,N_21375,N_21243);
and U21774 (N_21774,N_21410,N_21178);
nor U21775 (N_21775,N_21465,N_21078);
nor U21776 (N_21776,N_21561,N_21503);
nand U21777 (N_21777,N_21555,N_21363);
or U21778 (N_21778,N_21467,N_21055);
and U21779 (N_21779,N_21450,N_21154);
and U21780 (N_21780,N_21111,N_21244);
nand U21781 (N_21781,N_21586,N_21189);
or U21782 (N_21782,N_21475,N_21204);
nand U21783 (N_21783,N_21015,N_21025);
and U21784 (N_21784,N_21170,N_21137);
or U21785 (N_21785,N_21328,N_21155);
and U21786 (N_21786,N_21416,N_21246);
xnor U21787 (N_21787,N_21225,N_21578);
xor U21788 (N_21788,N_21331,N_21535);
xnor U21789 (N_21789,N_21277,N_21354);
or U21790 (N_21790,N_21032,N_21131);
xor U21791 (N_21791,N_21587,N_21018);
nand U21792 (N_21792,N_21305,N_21303);
xnor U21793 (N_21793,N_21368,N_21369);
nand U21794 (N_21794,N_21527,N_21280);
nand U21795 (N_21795,N_21272,N_21049);
and U21796 (N_21796,N_21143,N_21188);
nand U21797 (N_21797,N_21093,N_21435);
or U21798 (N_21798,N_21171,N_21103);
xor U21799 (N_21799,N_21311,N_21221);
or U21800 (N_21800,N_21099,N_21413);
nor U21801 (N_21801,N_21585,N_21142);
and U21802 (N_21802,N_21469,N_21121);
nor U21803 (N_21803,N_21460,N_21089);
nor U21804 (N_21804,N_21029,N_21083);
xor U21805 (N_21805,N_21085,N_21001);
and U21806 (N_21806,N_21130,N_21459);
or U21807 (N_21807,N_21310,N_21219);
and U21808 (N_21808,N_21057,N_21418);
and U21809 (N_21809,N_21013,N_21536);
nand U21810 (N_21810,N_21241,N_21096);
or U21811 (N_21811,N_21553,N_21537);
nand U21812 (N_21812,N_21259,N_21034);
and U21813 (N_21813,N_21452,N_21378);
and U21814 (N_21814,N_21072,N_21514);
nor U21815 (N_21815,N_21437,N_21270);
nand U21816 (N_21816,N_21420,N_21350);
and U21817 (N_21817,N_21091,N_21398);
nor U21818 (N_21818,N_21584,N_21116);
nor U21819 (N_21819,N_21440,N_21382);
nor U21820 (N_21820,N_21568,N_21551);
nor U21821 (N_21821,N_21227,N_21145);
nand U21822 (N_21822,N_21588,N_21485);
and U21823 (N_21823,N_21525,N_21040);
nand U21824 (N_21824,N_21347,N_21076);
nand U21825 (N_21825,N_21359,N_21088);
or U21826 (N_21826,N_21108,N_21401);
nand U21827 (N_21827,N_21412,N_21332);
nand U21828 (N_21828,N_21384,N_21545);
xor U21829 (N_21829,N_21056,N_21184);
nand U21830 (N_21830,N_21037,N_21278);
or U21831 (N_21831,N_21097,N_21434);
xnor U21832 (N_21832,N_21312,N_21301);
nor U21833 (N_21833,N_21399,N_21231);
nor U21834 (N_21834,N_21134,N_21207);
nand U21835 (N_21835,N_21110,N_21193);
and U21836 (N_21836,N_21411,N_21594);
and U21837 (N_21837,N_21292,N_21275);
xnor U21838 (N_21838,N_21379,N_21374);
nand U21839 (N_21839,N_21109,N_21361);
nand U21840 (N_21840,N_21390,N_21362);
nand U21841 (N_21841,N_21432,N_21035);
nor U21842 (N_21842,N_21308,N_21473);
xor U21843 (N_21843,N_21158,N_21447);
nand U21844 (N_21844,N_21453,N_21316);
or U21845 (N_21845,N_21356,N_21105);
or U21846 (N_21846,N_21008,N_21163);
and U21847 (N_21847,N_21474,N_21397);
or U21848 (N_21848,N_21429,N_21160);
and U21849 (N_21849,N_21269,N_21172);
nor U21850 (N_21850,N_21479,N_21472);
and U21851 (N_21851,N_21517,N_21443);
nand U21852 (N_21852,N_21220,N_21173);
nor U21853 (N_21853,N_21252,N_21530);
or U21854 (N_21854,N_21276,N_21287);
and U21855 (N_21855,N_21012,N_21086);
nand U21856 (N_21856,N_21216,N_21507);
nand U21857 (N_21857,N_21381,N_21339);
xnor U21858 (N_21858,N_21599,N_21214);
nand U21859 (N_21859,N_21344,N_21295);
xnor U21860 (N_21860,N_21166,N_21583);
and U21861 (N_21861,N_21304,N_21364);
or U21862 (N_21862,N_21296,N_21541);
or U21863 (N_21863,N_21122,N_21538);
nor U21864 (N_21864,N_21257,N_21314);
nand U21865 (N_21865,N_21141,N_21196);
or U21866 (N_21866,N_21523,N_21030);
nor U21867 (N_21867,N_21222,N_21501);
xor U21868 (N_21868,N_21115,N_21299);
xnor U21869 (N_21869,N_21092,N_21559);
nor U21870 (N_21870,N_21495,N_21007);
and U21871 (N_21871,N_21262,N_21079);
xor U21872 (N_21872,N_21106,N_21265);
or U21873 (N_21873,N_21273,N_21307);
or U21874 (N_21874,N_21306,N_21228);
nor U21875 (N_21875,N_21439,N_21090);
nand U21876 (N_21876,N_21456,N_21387);
and U21877 (N_21877,N_21168,N_21423);
nand U21878 (N_21878,N_21508,N_21487);
or U21879 (N_21879,N_21230,N_21238);
xor U21880 (N_21880,N_21199,N_21483);
nor U21881 (N_21881,N_21157,N_21309);
or U21882 (N_21882,N_21117,N_21470);
xnor U21883 (N_21883,N_21000,N_21478);
and U21884 (N_21884,N_21511,N_21249);
and U21885 (N_21885,N_21490,N_21119);
or U21886 (N_21886,N_21521,N_21489);
or U21887 (N_21887,N_21510,N_21058);
and U21888 (N_21888,N_21217,N_21026);
nand U21889 (N_21889,N_21421,N_21393);
or U21890 (N_21890,N_21488,N_21351);
or U21891 (N_21891,N_21161,N_21377);
or U21892 (N_21892,N_21552,N_21016);
and U21893 (N_21893,N_21444,N_21371);
or U21894 (N_21894,N_21337,N_21066);
or U21895 (N_21895,N_21203,N_21542);
nand U21896 (N_21896,N_21313,N_21209);
xor U21897 (N_21897,N_21370,N_21515);
and U21898 (N_21898,N_21336,N_21139);
and U21899 (N_21899,N_21208,N_21126);
xor U21900 (N_21900,N_21311,N_21055);
or U21901 (N_21901,N_21562,N_21275);
or U21902 (N_21902,N_21173,N_21503);
and U21903 (N_21903,N_21311,N_21220);
xnor U21904 (N_21904,N_21016,N_21146);
xnor U21905 (N_21905,N_21469,N_21219);
or U21906 (N_21906,N_21139,N_21295);
nand U21907 (N_21907,N_21185,N_21280);
nor U21908 (N_21908,N_21103,N_21091);
xnor U21909 (N_21909,N_21484,N_21405);
nand U21910 (N_21910,N_21066,N_21002);
xnor U21911 (N_21911,N_21162,N_21117);
nor U21912 (N_21912,N_21338,N_21521);
or U21913 (N_21913,N_21525,N_21277);
nor U21914 (N_21914,N_21156,N_21209);
nor U21915 (N_21915,N_21372,N_21112);
nor U21916 (N_21916,N_21095,N_21389);
and U21917 (N_21917,N_21218,N_21387);
nor U21918 (N_21918,N_21518,N_21426);
or U21919 (N_21919,N_21483,N_21001);
or U21920 (N_21920,N_21024,N_21054);
xor U21921 (N_21921,N_21192,N_21138);
or U21922 (N_21922,N_21371,N_21470);
nor U21923 (N_21923,N_21473,N_21204);
xor U21924 (N_21924,N_21306,N_21199);
nand U21925 (N_21925,N_21065,N_21465);
xnor U21926 (N_21926,N_21419,N_21449);
xnor U21927 (N_21927,N_21067,N_21036);
and U21928 (N_21928,N_21585,N_21058);
and U21929 (N_21929,N_21269,N_21410);
or U21930 (N_21930,N_21486,N_21017);
xor U21931 (N_21931,N_21506,N_21110);
nor U21932 (N_21932,N_21501,N_21509);
nand U21933 (N_21933,N_21347,N_21353);
and U21934 (N_21934,N_21061,N_21075);
nor U21935 (N_21935,N_21200,N_21434);
or U21936 (N_21936,N_21514,N_21183);
nand U21937 (N_21937,N_21445,N_21323);
xor U21938 (N_21938,N_21186,N_21538);
nor U21939 (N_21939,N_21452,N_21356);
nand U21940 (N_21940,N_21016,N_21299);
nor U21941 (N_21941,N_21508,N_21051);
and U21942 (N_21942,N_21420,N_21085);
xnor U21943 (N_21943,N_21446,N_21468);
nor U21944 (N_21944,N_21131,N_21270);
or U21945 (N_21945,N_21466,N_21474);
xor U21946 (N_21946,N_21139,N_21457);
nor U21947 (N_21947,N_21321,N_21146);
nand U21948 (N_21948,N_21355,N_21099);
and U21949 (N_21949,N_21250,N_21111);
and U21950 (N_21950,N_21019,N_21488);
nand U21951 (N_21951,N_21053,N_21078);
and U21952 (N_21952,N_21361,N_21067);
xor U21953 (N_21953,N_21179,N_21483);
and U21954 (N_21954,N_21056,N_21008);
xnor U21955 (N_21955,N_21498,N_21287);
xor U21956 (N_21956,N_21425,N_21454);
nand U21957 (N_21957,N_21155,N_21267);
or U21958 (N_21958,N_21319,N_21166);
and U21959 (N_21959,N_21528,N_21358);
and U21960 (N_21960,N_21324,N_21580);
and U21961 (N_21961,N_21202,N_21555);
xor U21962 (N_21962,N_21327,N_21429);
xor U21963 (N_21963,N_21564,N_21363);
or U21964 (N_21964,N_21323,N_21587);
and U21965 (N_21965,N_21006,N_21295);
or U21966 (N_21966,N_21366,N_21132);
and U21967 (N_21967,N_21448,N_21355);
or U21968 (N_21968,N_21067,N_21464);
nand U21969 (N_21969,N_21464,N_21352);
or U21970 (N_21970,N_21245,N_21173);
or U21971 (N_21971,N_21094,N_21483);
nor U21972 (N_21972,N_21301,N_21191);
or U21973 (N_21973,N_21413,N_21067);
nand U21974 (N_21974,N_21516,N_21321);
and U21975 (N_21975,N_21368,N_21555);
nor U21976 (N_21976,N_21112,N_21232);
xor U21977 (N_21977,N_21574,N_21473);
or U21978 (N_21978,N_21171,N_21487);
xnor U21979 (N_21979,N_21163,N_21475);
and U21980 (N_21980,N_21523,N_21590);
nor U21981 (N_21981,N_21581,N_21511);
xnor U21982 (N_21982,N_21188,N_21231);
and U21983 (N_21983,N_21320,N_21564);
xnor U21984 (N_21984,N_21463,N_21486);
and U21985 (N_21985,N_21599,N_21393);
and U21986 (N_21986,N_21041,N_21025);
nand U21987 (N_21987,N_21409,N_21167);
and U21988 (N_21988,N_21147,N_21166);
nand U21989 (N_21989,N_21354,N_21480);
xnor U21990 (N_21990,N_21512,N_21018);
nor U21991 (N_21991,N_21020,N_21065);
xor U21992 (N_21992,N_21017,N_21495);
xor U21993 (N_21993,N_21406,N_21280);
nor U21994 (N_21994,N_21500,N_21057);
nor U21995 (N_21995,N_21529,N_21376);
nor U21996 (N_21996,N_21494,N_21081);
or U21997 (N_21997,N_21485,N_21312);
nand U21998 (N_21998,N_21487,N_21303);
and U21999 (N_21999,N_21521,N_21045);
or U22000 (N_22000,N_21191,N_21215);
nand U22001 (N_22001,N_21213,N_21049);
or U22002 (N_22002,N_21219,N_21578);
xnor U22003 (N_22003,N_21499,N_21466);
nand U22004 (N_22004,N_21038,N_21281);
xnor U22005 (N_22005,N_21388,N_21083);
or U22006 (N_22006,N_21589,N_21379);
nor U22007 (N_22007,N_21337,N_21394);
xor U22008 (N_22008,N_21298,N_21088);
or U22009 (N_22009,N_21230,N_21216);
nand U22010 (N_22010,N_21326,N_21389);
xnor U22011 (N_22011,N_21019,N_21223);
or U22012 (N_22012,N_21572,N_21038);
xor U22013 (N_22013,N_21461,N_21355);
nand U22014 (N_22014,N_21518,N_21063);
xnor U22015 (N_22015,N_21186,N_21422);
or U22016 (N_22016,N_21030,N_21132);
nand U22017 (N_22017,N_21075,N_21148);
or U22018 (N_22018,N_21420,N_21472);
or U22019 (N_22019,N_21102,N_21421);
and U22020 (N_22020,N_21556,N_21215);
xnor U22021 (N_22021,N_21542,N_21415);
nand U22022 (N_22022,N_21299,N_21319);
nand U22023 (N_22023,N_21051,N_21549);
xor U22024 (N_22024,N_21026,N_21339);
nand U22025 (N_22025,N_21467,N_21327);
nor U22026 (N_22026,N_21352,N_21573);
or U22027 (N_22027,N_21231,N_21318);
nor U22028 (N_22028,N_21177,N_21491);
nor U22029 (N_22029,N_21067,N_21401);
nor U22030 (N_22030,N_21088,N_21028);
xnor U22031 (N_22031,N_21406,N_21266);
nand U22032 (N_22032,N_21404,N_21139);
nand U22033 (N_22033,N_21038,N_21330);
xor U22034 (N_22034,N_21094,N_21480);
or U22035 (N_22035,N_21561,N_21566);
xnor U22036 (N_22036,N_21345,N_21283);
nand U22037 (N_22037,N_21439,N_21013);
and U22038 (N_22038,N_21440,N_21433);
nor U22039 (N_22039,N_21018,N_21353);
nand U22040 (N_22040,N_21461,N_21275);
and U22041 (N_22041,N_21193,N_21175);
nand U22042 (N_22042,N_21222,N_21266);
and U22043 (N_22043,N_21585,N_21344);
nand U22044 (N_22044,N_21342,N_21254);
nand U22045 (N_22045,N_21439,N_21496);
or U22046 (N_22046,N_21238,N_21444);
xnor U22047 (N_22047,N_21454,N_21049);
nand U22048 (N_22048,N_21063,N_21228);
or U22049 (N_22049,N_21029,N_21542);
nand U22050 (N_22050,N_21284,N_21154);
xnor U22051 (N_22051,N_21069,N_21308);
or U22052 (N_22052,N_21593,N_21393);
xor U22053 (N_22053,N_21281,N_21121);
or U22054 (N_22054,N_21541,N_21181);
and U22055 (N_22055,N_21329,N_21337);
and U22056 (N_22056,N_21409,N_21364);
nor U22057 (N_22057,N_21388,N_21392);
nand U22058 (N_22058,N_21476,N_21318);
xnor U22059 (N_22059,N_21473,N_21272);
nor U22060 (N_22060,N_21095,N_21074);
and U22061 (N_22061,N_21571,N_21061);
nand U22062 (N_22062,N_21570,N_21451);
nand U22063 (N_22063,N_21524,N_21240);
and U22064 (N_22064,N_21042,N_21045);
nor U22065 (N_22065,N_21051,N_21239);
nor U22066 (N_22066,N_21187,N_21320);
and U22067 (N_22067,N_21310,N_21548);
nand U22068 (N_22068,N_21146,N_21238);
and U22069 (N_22069,N_21400,N_21125);
or U22070 (N_22070,N_21207,N_21356);
nor U22071 (N_22071,N_21256,N_21210);
nor U22072 (N_22072,N_21580,N_21526);
nor U22073 (N_22073,N_21240,N_21481);
or U22074 (N_22074,N_21316,N_21400);
nand U22075 (N_22075,N_21183,N_21196);
and U22076 (N_22076,N_21491,N_21019);
xnor U22077 (N_22077,N_21083,N_21499);
and U22078 (N_22078,N_21464,N_21271);
xor U22079 (N_22079,N_21231,N_21591);
xnor U22080 (N_22080,N_21242,N_21597);
nor U22081 (N_22081,N_21014,N_21225);
nand U22082 (N_22082,N_21566,N_21553);
xnor U22083 (N_22083,N_21097,N_21137);
or U22084 (N_22084,N_21543,N_21436);
or U22085 (N_22085,N_21421,N_21302);
nand U22086 (N_22086,N_21503,N_21115);
nor U22087 (N_22087,N_21297,N_21309);
and U22088 (N_22088,N_21413,N_21386);
xnor U22089 (N_22089,N_21375,N_21269);
or U22090 (N_22090,N_21414,N_21171);
nor U22091 (N_22091,N_21561,N_21554);
and U22092 (N_22092,N_21531,N_21265);
nor U22093 (N_22093,N_21161,N_21599);
nand U22094 (N_22094,N_21116,N_21353);
nand U22095 (N_22095,N_21412,N_21103);
and U22096 (N_22096,N_21256,N_21034);
and U22097 (N_22097,N_21585,N_21407);
nor U22098 (N_22098,N_21335,N_21189);
and U22099 (N_22099,N_21526,N_21014);
nand U22100 (N_22100,N_21244,N_21509);
nand U22101 (N_22101,N_21039,N_21246);
or U22102 (N_22102,N_21561,N_21164);
and U22103 (N_22103,N_21542,N_21153);
xnor U22104 (N_22104,N_21429,N_21409);
nand U22105 (N_22105,N_21022,N_21307);
nand U22106 (N_22106,N_21136,N_21225);
or U22107 (N_22107,N_21502,N_21128);
or U22108 (N_22108,N_21560,N_21064);
xor U22109 (N_22109,N_21345,N_21445);
xor U22110 (N_22110,N_21143,N_21033);
xnor U22111 (N_22111,N_21389,N_21016);
xnor U22112 (N_22112,N_21432,N_21471);
nor U22113 (N_22113,N_21264,N_21190);
nand U22114 (N_22114,N_21314,N_21350);
nor U22115 (N_22115,N_21552,N_21540);
or U22116 (N_22116,N_21432,N_21236);
or U22117 (N_22117,N_21128,N_21195);
xnor U22118 (N_22118,N_21284,N_21589);
or U22119 (N_22119,N_21516,N_21164);
nor U22120 (N_22120,N_21263,N_21485);
nand U22121 (N_22121,N_21217,N_21345);
and U22122 (N_22122,N_21017,N_21050);
xor U22123 (N_22123,N_21528,N_21173);
and U22124 (N_22124,N_21400,N_21218);
or U22125 (N_22125,N_21187,N_21301);
nor U22126 (N_22126,N_21330,N_21558);
xnor U22127 (N_22127,N_21435,N_21162);
nor U22128 (N_22128,N_21403,N_21018);
nand U22129 (N_22129,N_21532,N_21300);
xnor U22130 (N_22130,N_21304,N_21181);
nand U22131 (N_22131,N_21129,N_21425);
and U22132 (N_22132,N_21486,N_21182);
and U22133 (N_22133,N_21598,N_21099);
nor U22134 (N_22134,N_21033,N_21391);
nor U22135 (N_22135,N_21068,N_21563);
and U22136 (N_22136,N_21331,N_21055);
xor U22137 (N_22137,N_21170,N_21222);
nor U22138 (N_22138,N_21313,N_21026);
or U22139 (N_22139,N_21295,N_21045);
or U22140 (N_22140,N_21269,N_21422);
and U22141 (N_22141,N_21141,N_21193);
nor U22142 (N_22142,N_21004,N_21331);
xor U22143 (N_22143,N_21502,N_21181);
xnor U22144 (N_22144,N_21344,N_21198);
and U22145 (N_22145,N_21343,N_21101);
or U22146 (N_22146,N_21280,N_21337);
xnor U22147 (N_22147,N_21343,N_21125);
xor U22148 (N_22148,N_21529,N_21047);
or U22149 (N_22149,N_21410,N_21383);
or U22150 (N_22150,N_21074,N_21367);
nor U22151 (N_22151,N_21341,N_21202);
nor U22152 (N_22152,N_21389,N_21235);
nand U22153 (N_22153,N_21128,N_21577);
or U22154 (N_22154,N_21393,N_21578);
or U22155 (N_22155,N_21424,N_21065);
xor U22156 (N_22156,N_21461,N_21298);
or U22157 (N_22157,N_21401,N_21531);
or U22158 (N_22158,N_21344,N_21150);
nand U22159 (N_22159,N_21340,N_21446);
nand U22160 (N_22160,N_21589,N_21195);
nand U22161 (N_22161,N_21135,N_21113);
nand U22162 (N_22162,N_21590,N_21509);
xnor U22163 (N_22163,N_21438,N_21455);
nand U22164 (N_22164,N_21384,N_21215);
nor U22165 (N_22165,N_21025,N_21460);
or U22166 (N_22166,N_21066,N_21229);
nor U22167 (N_22167,N_21580,N_21181);
xnor U22168 (N_22168,N_21279,N_21190);
or U22169 (N_22169,N_21180,N_21577);
and U22170 (N_22170,N_21016,N_21326);
nor U22171 (N_22171,N_21156,N_21529);
nor U22172 (N_22172,N_21223,N_21578);
xnor U22173 (N_22173,N_21394,N_21099);
nand U22174 (N_22174,N_21193,N_21066);
or U22175 (N_22175,N_21239,N_21379);
nand U22176 (N_22176,N_21254,N_21220);
nor U22177 (N_22177,N_21550,N_21383);
or U22178 (N_22178,N_21026,N_21516);
xor U22179 (N_22179,N_21337,N_21070);
or U22180 (N_22180,N_21542,N_21221);
nor U22181 (N_22181,N_21011,N_21170);
nand U22182 (N_22182,N_21201,N_21423);
nand U22183 (N_22183,N_21375,N_21169);
and U22184 (N_22184,N_21207,N_21452);
or U22185 (N_22185,N_21471,N_21097);
xnor U22186 (N_22186,N_21507,N_21153);
or U22187 (N_22187,N_21455,N_21143);
nor U22188 (N_22188,N_21207,N_21466);
and U22189 (N_22189,N_21493,N_21497);
xnor U22190 (N_22190,N_21499,N_21434);
or U22191 (N_22191,N_21041,N_21061);
and U22192 (N_22192,N_21357,N_21149);
nor U22193 (N_22193,N_21522,N_21373);
xnor U22194 (N_22194,N_21290,N_21152);
or U22195 (N_22195,N_21468,N_21408);
nor U22196 (N_22196,N_21550,N_21067);
xor U22197 (N_22197,N_21509,N_21358);
or U22198 (N_22198,N_21053,N_21521);
or U22199 (N_22199,N_21182,N_21124);
xor U22200 (N_22200,N_22038,N_21867);
and U22201 (N_22201,N_22140,N_21664);
or U22202 (N_22202,N_22172,N_22144);
or U22203 (N_22203,N_21776,N_22195);
and U22204 (N_22204,N_21922,N_21904);
nor U22205 (N_22205,N_21782,N_22008);
xor U22206 (N_22206,N_21696,N_21972);
and U22207 (N_22207,N_22112,N_21953);
xnor U22208 (N_22208,N_21896,N_21766);
nor U22209 (N_22209,N_22198,N_21811);
xnor U22210 (N_22210,N_22013,N_22095);
and U22211 (N_22211,N_22128,N_21930);
xnor U22212 (N_22212,N_22145,N_21638);
nand U22213 (N_22213,N_21987,N_21851);
nand U22214 (N_22214,N_21626,N_21882);
and U22215 (N_22215,N_22066,N_22050);
or U22216 (N_22216,N_21752,N_22031);
xor U22217 (N_22217,N_21645,N_21715);
and U22218 (N_22218,N_21939,N_22016);
xor U22219 (N_22219,N_21886,N_22176);
or U22220 (N_22220,N_22025,N_22143);
and U22221 (N_22221,N_22097,N_22053);
and U22222 (N_22222,N_21880,N_22045);
nor U22223 (N_22223,N_22071,N_21614);
nand U22224 (N_22224,N_22147,N_21686);
and U22225 (N_22225,N_22076,N_21995);
nor U22226 (N_22226,N_22155,N_21672);
xor U22227 (N_22227,N_21746,N_21813);
and U22228 (N_22228,N_21670,N_21712);
nand U22229 (N_22229,N_22160,N_21908);
xor U22230 (N_22230,N_21871,N_21868);
or U22231 (N_22231,N_22075,N_21678);
nand U22232 (N_22232,N_21780,N_21679);
nand U22233 (N_22233,N_21846,N_21706);
xor U22234 (N_22234,N_22110,N_21666);
nor U22235 (N_22235,N_22019,N_22104);
nand U22236 (N_22236,N_21906,N_21753);
or U22237 (N_22237,N_22139,N_21762);
and U22238 (N_22238,N_22138,N_21899);
and U22239 (N_22239,N_21844,N_22191);
or U22240 (N_22240,N_22190,N_22062);
nand U22241 (N_22241,N_21903,N_21869);
nor U22242 (N_22242,N_22094,N_21817);
or U22243 (N_22243,N_22156,N_22065);
and U22244 (N_22244,N_22186,N_21719);
nor U22245 (N_22245,N_22010,N_21883);
and U22246 (N_22246,N_22039,N_21659);
nand U22247 (N_22247,N_21677,N_22153);
and U22248 (N_22248,N_22085,N_21769);
or U22249 (N_22249,N_22074,N_22126);
and U22250 (N_22250,N_22183,N_21876);
and U22251 (N_22251,N_21763,N_21718);
nor U22252 (N_22252,N_22079,N_21759);
nand U22253 (N_22253,N_21842,N_22026);
or U22254 (N_22254,N_22158,N_22057);
or U22255 (N_22255,N_21757,N_21612);
or U22256 (N_22256,N_21680,N_22103);
and U22257 (N_22257,N_22168,N_21892);
nor U22258 (N_22258,N_21747,N_21815);
nand U22259 (N_22259,N_21635,N_21702);
xor U22260 (N_22260,N_21803,N_21835);
xor U22261 (N_22261,N_21991,N_22020);
nand U22262 (N_22262,N_21893,N_21687);
xnor U22263 (N_22263,N_21605,N_21743);
xnor U22264 (N_22264,N_21826,N_22100);
nand U22265 (N_22265,N_21970,N_21713);
nor U22266 (N_22266,N_21681,N_22122);
and U22267 (N_22267,N_21839,N_21784);
and U22268 (N_22268,N_21971,N_21717);
xor U22269 (N_22269,N_21658,N_22180);
and U22270 (N_22270,N_21721,N_21938);
xnor U22271 (N_22271,N_22070,N_21996);
and U22272 (N_22272,N_21828,N_22119);
or U22273 (N_22273,N_21640,N_21733);
xnor U22274 (N_22274,N_22188,N_21969);
xor U22275 (N_22275,N_21671,N_21951);
or U22276 (N_22276,N_21796,N_21935);
or U22277 (N_22277,N_21631,N_21850);
nor U22278 (N_22278,N_21616,N_22197);
or U22279 (N_22279,N_21802,N_22022);
xor U22280 (N_22280,N_21642,N_21989);
nand U22281 (N_22281,N_21716,N_21806);
nor U22282 (N_22282,N_21646,N_21894);
and U22283 (N_22283,N_22012,N_22014);
nand U22284 (N_22284,N_21872,N_22108);
xnor U22285 (N_22285,N_21984,N_21841);
nor U22286 (N_22286,N_21755,N_21768);
xor U22287 (N_22287,N_21960,N_22090);
xnor U22288 (N_22288,N_22078,N_21629);
xnor U22289 (N_22289,N_22027,N_21760);
and U22290 (N_22290,N_21812,N_21600);
or U22291 (N_22291,N_21695,N_22196);
or U22292 (N_22292,N_21607,N_21699);
or U22293 (N_22293,N_21736,N_21750);
and U22294 (N_22294,N_21956,N_21902);
nor U22295 (N_22295,N_21667,N_21952);
and U22296 (N_22296,N_21929,N_21620);
nor U22297 (N_22297,N_22106,N_21810);
or U22298 (N_22298,N_21654,N_21853);
nand U22299 (N_22299,N_21915,N_21926);
nand U22300 (N_22300,N_21800,N_21805);
and U22301 (N_22301,N_21982,N_22157);
nand U22302 (N_22302,N_21669,N_21794);
and U22303 (N_22303,N_21820,N_21955);
and U22304 (N_22304,N_21829,N_21861);
nand U22305 (N_22305,N_22043,N_21824);
xnor U22306 (N_22306,N_22129,N_21613);
nor U22307 (N_22307,N_22134,N_22093);
and U22308 (N_22308,N_21986,N_22181);
and U22309 (N_22309,N_21676,N_22189);
xor U22310 (N_22310,N_21980,N_21931);
xnor U22311 (N_22311,N_22150,N_21879);
nor U22312 (N_22312,N_21675,N_22148);
xor U22313 (N_22313,N_22164,N_22179);
nor U22314 (N_22314,N_21916,N_22089);
or U22315 (N_22315,N_21637,N_21840);
nor U22316 (N_22316,N_21749,N_21847);
xor U22317 (N_22317,N_21804,N_21885);
or U22318 (N_22318,N_21891,N_22193);
and U22319 (N_22319,N_22064,N_21807);
or U22320 (N_22320,N_21641,N_21798);
and U22321 (N_22321,N_21632,N_21604);
and U22322 (N_22322,N_21725,N_22044);
and U22323 (N_22323,N_21808,N_21961);
nand U22324 (N_22324,N_22046,N_21801);
xnor U22325 (N_22325,N_22091,N_22033);
xor U22326 (N_22326,N_21979,N_22199);
and U22327 (N_22327,N_21799,N_21771);
or U22328 (N_22328,N_21773,N_21889);
xnor U22329 (N_22329,N_21857,N_21788);
nor U22330 (N_22330,N_21775,N_22000);
xnor U22331 (N_22331,N_22166,N_22009);
or U22332 (N_22332,N_21643,N_21774);
nor U22333 (N_22333,N_21742,N_21878);
nor U22334 (N_22334,N_21954,N_21981);
xnor U22335 (N_22335,N_21739,N_21787);
xor U22336 (N_22336,N_21709,N_22177);
nand U22337 (N_22337,N_22086,N_21625);
and U22338 (N_22338,N_21705,N_21647);
and U22339 (N_22339,N_21772,N_21884);
or U22340 (N_22340,N_21875,N_22021);
nor U22341 (N_22341,N_21897,N_21726);
and U22342 (N_22342,N_21785,N_21900);
and U22343 (N_22343,N_22133,N_21907);
and U22344 (N_22344,N_21724,N_21978);
xnor U22345 (N_22345,N_21966,N_21974);
nor U22346 (N_22346,N_21668,N_21852);
and U22347 (N_22347,N_21983,N_22137);
nand U22348 (N_22348,N_22167,N_22092);
xnor U22349 (N_22349,N_21649,N_21674);
or U22350 (N_22350,N_21873,N_22162);
xnor U22351 (N_22351,N_21823,N_21707);
or U22352 (N_22352,N_22120,N_21814);
nand U22353 (N_22353,N_21618,N_22081);
xnor U22354 (N_22354,N_22135,N_21837);
xor U22355 (N_22355,N_21700,N_21661);
nand U22356 (N_22356,N_22154,N_21656);
or U22357 (N_22357,N_21791,N_21834);
nand U22358 (N_22358,N_21633,N_22004);
nor U22359 (N_22359,N_21818,N_21624);
and U22360 (N_22360,N_21948,N_22011);
xor U22361 (N_22361,N_21601,N_21731);
nand U22362 (N_22362,N_22099,N_22109);
and U22363 (N_22363,N_21610,N_21919);
and U22364 (N_22364,N_21786,N_21636);
nor U22365 (N_22365,N_21693,N_21608);
nor U22366 (N_22366,N_21909,N_22114);
xnor U22367 (N_22367,N_21781,N_21660);
xor U22368 (N_22368,N_21941,N_22121);
and U22369 (N_22369,N_22015,N_22047);
nor U22370 (N_22370,N_21911,N_22132);
nand U22371 (N_22371,N_22141,N_22049);
xor U22372 (N_22372,N_21859,N_22151);
nand U22373 (N_22373,N_21682,N_21630);
or U22374 (N_22374,N_22058,N_22060);
nor U22375 (N_22375,N_21816,N_21890);
xor U22376 (N_22376,N_21964,N_21905);
nand U22377 (N_22377,N_22068,N_21827);
or U22378 (N_22378,N_21704,N_21959);
or U22379 (N_22379,N_22069,N_21862);
nor U22380 (N_22380,N_21698,N_22073);
nand U22381 (N_22381,N_21936,N_22037);
nor U22382 (N_22382,N_22107,N_22123);
and U22383 (N_22383,N_21934,N_22115);
and U22384 (N_22384,N_21925,N_21790);
nand U22385 (N_22385,N_21655,N_22127);
nor U22386 (N_22386,N_21606,N_21777);
nor U22387 (N_22387,N_21898,N_21783);
or U22388 (N_22388,N_21756,N_21740);
and U22389 (N_22389,N_21701,N_21703);
nor U22390 (N_22390,N_21877,N_22113);
and U22391 (N_22391,N_22059,N_21831);
xnor U22392 (N_22392,N_21628,N_21963);
nand U22393 (N_22393,N_22161,N_21663);
and U22394 (N_22394,N_22051,N_22175);
xor U22395 (N_22395,N_22149,N_22054);
or U22396 (N_22396,N_22152,N_22159);
or U22397 (N_22397,N_21792,N_21723);
nor U22398 (N_22398,N_21751,N_22005);
xnor U22399 (N_22399,N_22024,N_21967);
or U22400 (N_22400,N_22018,N_21830);
and U22401 (N_22401,N_21819,N_21838);
nand U22402 (N_22402,N_22174,N_21665);
and U22403 (N_22403,N_21990,N_21860);
xnor U22404 (N_22404,N_21732,N_22087);
xor U22405 (N_22405,N_21738,N_21843);
nor U22406 (N_22406,N_21692,N_21942);
and U22407 (N_22407,N_22178,N_21758);
nand U22408 (N_22408,N_21809,N_22096);
nand U22409 (N_22409,N_21789,N_22001);
xnor U22410 (N_22410,N_22056,N_21965);
nor U22411 (N_22411,N_21968,N_21727);
nand U22412 (N_22412,N_21688,N_21634);
or U22413 (N_22413,N_22146,N_22194);
or U22414 (N_22414,N_21694,N_21950);
nand U22415 (N_22415,N_22007,N_21945);
xnor U22416 (N_22416,N_21767,N_21683);
nor U22417 (N_22417,N_22136,N_21988);
and U22418 (N_22418,N_22105,N_22002);
xnor U22419 (N_22419,N_22030,N_22063);
or U22420 (N_22420,N_21895,N_22173);
nand U22421 (N_22421,N_21977,N_21985);
nor U22422 (N_22422,N_21833,N_21910);
or U22423 (N_22423,N_21914,N_21888);
xnor U22424 (N_22424,N_21822,N_21744);
or U22425 (N_22425,N_22171,N_21754);
nor U22426 (N_22426,N_21924,N_21741);
or U22427 (N_22427,N_21735,N_21691);
xor U22428 (N_22428,N_21650,N_21848);
and U22429 (N_22429,N_22040,N_22042);
and U22430 (N_22430,N_22023,N_21651);
nand U22431 (N_22431,N_22102,N_21918);
nor U22432 (N_22432,N_21611,N_21997);
and U22433 (N_22433,N_22118,N_21722);
nand U22434 (N_22434,N_22084,N_21958);
and U22435 (N_22435,N_22187,N_21623);
and U22436 (N_22436,N_21975,N_21881);
nor U22437 (N_22437,N_22142,N_21845);
nor U22438 (N_22438,N_21856,N_21998);
and U22439 (N_22439,N_22017,N_21615);
and U22440 (N_22440,N_21730,N_21684);
nand U22441 (N_22441,N_21887,N_22165);
and U22442 (N_22442,N_21825,N_22163);
and U22443 (N_22443,N_22124,N_22003);
xnor U22444 (N_22444,N_21764,N_21748);
nand U22445 (N_22445,N_21653,N_21689);
xor U22446 (N_22446,N_21947,N_22052);
nor U22447 (N_22447,N_21797,N_21648);
xnor U22448 (N_22448,N_22029,N_21943);
and U22449 (N_22449,N_21778,N_22125);
nand U22450 (N_22450,N_21609,N_21913);
and U22451 (N_22451,N_21933,N_22080);
nand U22452 (N_22452,N_22067,N_21836);
or U22453 (N_22453,N_21865,N_21793);
nand U22454 (N_22454,N_21923,N_21944);
xnor U22455 (N_22455,N_21602,N_21921);
or U22456 (N_22456,N_21940,N_22192);
xor U22457 (N_22457,N_21946,N_21729);
and U22458 (N_22458,N_21657,N_21999);
and U22459 (N_22459,N_21644,N_22088);
or U22460 (N_22460,N_21673,N_21870);
nand U22461 (N_22461,N_21779,N_21832);
xnor U22462 (N_22462,N_21973,N_21901);
and U22463 (N_22463,N_21603,N_21949);
or U22464 (N_22464,N_21690,N_21962);
or U22465 (N_22465,N_22055,N_21874);
xor U22466 (N_22466,N_21745,N_21854);
xnor U22467 (N_22467,N_22130,N_21697);
or U22468 (N_22468,N_21932,N_22169);
or U22469 (N_22469,N_21652,N_21863);
and U22470 (N_22470,N_21866,N_21619);
nor U22471 (N_22471,N_22131,N_21928);
nand U22472 (N_22472,N_21770,N_22101);
nand U22473 (N_22473,N_21849,N_22182);
or U22474 (N_22474,N_21992,N_22032);
or U22475 (N_22475,N_22006,N_22028);
nor U22476 (N_22476,N_21734,N_22035);
and U22477 (N_22477,N_21912,N_21821);
or U22478 (N_22478,N_21685,N_21617);
nor U22479 (N_22479,N_21937,N_22034);
and U22480 (N_22480,N_22116,N_21994);
or U22481 (N_22481,N_21957,N_21927);
or U22482 (N_22482,N_21621,N_21993);
xor U22483 (N_22483,N_21765,N_22117);
and U22484 (N_22484,N_21622,N_21795);
or U22485 (N_22485,N_22184,N_22072);
and U22486 (N_22486,N_22185,N_21976);
or U22487 (N_22487,N_22041,N_21761);
xnor U22488 (N_22488,N_21920,N_22111);
nor U22489 (N_22489,N_21737,N_22082);
nor U22490 (N_22490,N_21855,N_21711);
nor U22491 (N_22491,N_21662,N_22077);
nor U22492 (N_22492,N_21728,N_21714);
and U22493 (N_22493,N_22061,N_21710);
nor U22494 (N_22494,N_21917,N_21864);
nor U22495 (N_22495,N_21858,N_22083);
xor U22496 (N_22496,N_21627,N_21708);
xnor U22497 (N_22497,N_22048,N_21720);
and U22498 (N_22498,N_22098,N_22170);
and U22499 (N_22499,N_21639,N_22036);
and U22500 (N_22500,N_22130,N_21899);
and U22501 (N_22501,N_21843,N_22123);
xor U22502 (N_22502,N_21765,N_21829);
xnor U22503 (N_22503,N_21770,N_21837);
xnor U22504 (N_22504,N_22064,N_21758);
nand U22505 (N_22505,N_22113,N_21992);
xor U22506 (N_22506,N_21852,N_21997);
or U22507 (N_22507,N_21856,N_21640);
and U22508 (N_22508,N_22121,N_21857);
and U22509 (N_22509,N_22126,N_21831);
or U22510 (N_22510,N_21766,N_21610);
xnor U22511 (N_22511,N_21760,N_21703);
or U22512 (N_22512,N_22026,N_22157);
nor U22513 (N_22513,N_21728,N_21748);
nor U22514 (N_22514,N_21657,N_21866);
xor U22515 (N_22515,N_21952,N_21869);
or U22516 (N_22516,N_21820,N_21681);
and U22517 (N_22517,N_21908,N_22162);
nor U22518 (N_22518,N_22179,N_21911);
and U22519 (N_22519,N_21832,N_21929);
xnor U22520 (N_22520,N_21946,N_21810);
or U22521 (N_22521,N_21653,N_21825);
and U22522 (N_22522,N_21706,N_21843);
and U22523 (N_22523,N_22109,N_21917);
xor U22524 (N_22524,N_21781,N_21718);
nor U22525 (N_22525,N_22094,N_21637);
xnor U22526 (N_22526,N_21782,N_22143);
or U22527 (N_22527,N_21868,N_22132);
nor U22528 (N_22528,N_21943,N_22135);
and U22529 (N_22529,N_22123,N_21728);
and U22530 (N_22530,N_22021,N_21884);
or U22531 (N_22531,N_21793,N_21919);
xnor U22532 (N_22532,N_22122,N_21801);
xor U22533 (N_22533,N_21905,N_21846);
nor U22534 (N_22534,N_22102,N_21668);
and U22535 (N_22535,N_21625,N_21720);
or U22536 (N_22536,N_21626,N_21753);
nand U22537 (N_22537,N_21778,N_21917);
nor U22538 (N_22538,N_21997,N_21682);
and U22539 (N_22539,N_21711,N_21971);
nand U22540 (N_22540,N_21703,N_22135);
nor U22541 (N_22541,N_21795,N_22049);
nor U22542 (N_22542,N_21839,N_22026);
nor U22543 (N_22543,N_21851,N_21854);
or U22544 (N_22544,N_21671,N_21649);
or U22545 (N_22545,N_21738,N_21744);
nor U22546 (N_22546,N_22197,N_21674);
or U22547 (N_22547,N_21825,N_21615);
and U22548 (N_22548,N_21655,N_22017);
or U22549 (N_22549,N_22015,N_21745);
and U22550 (N_22550,N_21705,N_22009);
nor U22551 (N_22551,N_22172,N_22171);
nand U22552 (N_22552,N_22124,N_21943);
nor U22553 (N_22553,N_21605,N_21933);
and U22554 (N_22554,N_22068,N_21635);
nand U22555 (N_22555,N_21908,N_21755);
xnor U22556 (N_22556,N_21820,N_21942);
and U22557 (N_22557,N_22133,N_21837);
nand U22558 (N_22558,N_21647,N_22175);
or U22559 (N_22559,N_22163,N_21822);
and U22560 (N_22560,N_21963,N_21617);
xor U22561 (N_22561,N_22141,N_21863);
and U22562 (N_22562,N_21983,N_21863);
and U22563 (N_22563,N_21849,N_21833);
nand U22564 (N_22564,N_22111,N_22122);
nor U22565 (N_22565,N_21754,N_22008);
nand U22566 (N_22566,N_21777,N_22108);
nand U22567 (N_22567,N_22116,N_21762);
xor U22568 (N_22568,N_21669,N_22124);
and U22569 (N_22569,N_22036,N_21811);
or U22570 (N_22570,N_21822,N_22012);
nand U22571 (N_22571,N_21998,N_22033);
xor U22572 (N_22572,N_21884,N_21675);
or U22573 (N_22573,N_21788,N_21664);
nor U22574 (N_22574,N_21948,N_22194);
nor U22575 (N_22575,N_22068,N_21849);
xor U22576 (N_22576,N_21711,N_21951);
nor U22577 (N_22577,N_21837,N_21947);
nor U22578 (N_22578,N_22102,N_21641);
and U22579 (N_22579,N_22192,N_21770);
or U22580 (N_22580,N_21959,N_22015);
or U22581 (N_22581,N_21904,N_21921);
and U22582 (N_22582,N_21886,N_21629);
nand U22583 (N_22583,N_22048,N_21959);
xnor U22584 (N_22584,N_21716,N_22051);
nor U22585 (N_22585,N_22052,N_21736);
or U22586 (N_22586,N_21645,N_21986);
nand U22587 (N_22587,N_22138,N_22049);
xor U22588 (N_22588,N_21902,N_21697);
and U22589 (N_22589,N_22168,N_21737);
or U22590 (N_22590,N_21677,N_21877);
or U22591 (N_22591,N_21962,N_21895);
nor U22592 (N_22592,N_21873,N_21676);
or U22593 (N_22593,N_22149,N_21858);
nor U22594 (N_22594,N_21944,N_22082);
nor U22595 (N_22595,N_21777,N_21998);
or U22596 (N_22596,N_21816,N_22094);
xor U22597 (N_22597,N_22131,N_21797);
nor U22598 (N_22598,N_21618,N_21993);
and U22599 (N_22599,N_21696,N_21882);
nand U22600 (N_22600,N_21949,N_21614);
or U22601 (N_22601,N_21608,N_21842);
and U22602 (N_22602,N_22027,N_21725);
nor U22603 (N_22603,N_21830,N_21908);
nor U22604 (N_22604,N_21772,N_22030);
xnor U22605 (N_22605,N_21960,N_21889);
and U22606 (N_22606,N_21848,N_21680);
and U22607 (N_22607,N_22005,N_22183);
xnor U22608 (N_22608,N_21745,N_22149);
xor U22609 (N_22609,N_21913,N_22113);
and U22610 (N_22610,N_22125,N_22176);
or U22611 (N_22611,N_21850,N_21882);
and U22612 (N_22612,N_22124,N_21631);
or U22613 (N_22613,N_22146,N_21690);
nor U22614 (N_22614,N_22042,N_21819);
and U22615 (N_22615,N_21613,N_21855);
xor U22616 (N_22616,N_22044,N_21796);
or U22617 (N_22617,N_21972,N_22166);
nand U22618 (N_22618,N_21600,N_21623);
xnor U22619 (N_22619,N_21755,N_22129);
or U22620 (N_22620,N_21885,N_22014);
or U22621 (N_22621,N_21808,N_22067);
or U22622 (N_22622,N_21977,N_22156);
xnor U22623 (N_22623,N_22118,N_22006);
or U22624 (N_22624,N_21997,N_21748);
or U22625 (N_22625,N_21840,N_21949);
nor U22626 (N_22626,N_22142,N_22049);
xnor U22627 (N_22627,N_21773,N_21968);
or U22628 (N_22628,N_21946,N_21655);
and U22629 (N_22629,N_21656,N_22094);
nand U22630 (N_22630,N_21637,N_21863);
or U22631 (N_22631,N_22095,N_21956);
and U22632 (N_22632,N_22109,N_22179);
xnor U22633 (N_22633,N_22114,N_21860);
nor U22634 (N_22634,N_21816,N_22153);
and U22635 (N_22635,N_22104,N_21662);
xnor U22636 (N_22636,N_21809,N_21740);
nand U22637 (N_22637,N_21664,N_21934);
nor U22638 (N_22638,N_21920,N_21929);
nand U22639 (N_22639,N_21945,N_21767);
or U22640 (N_22640,N_21746,N_21678);
nand U22641 (N_22641,N_21910,N_21985);
nor U22642 (N_22642,N_21655,N_21687);
or U22643 (N_22643,N_21819,N_21882);
nand U22644 (N_22644,N_22075,N_21715);
nand U22645 (N_22645,N_21668,N_21632);
nand U22646 (N_22646,N_21784,N_21903);
nor U22647 (N_22647,N_21998,N_21938);
nor U22648 (N_22648,N_22046,N_21941);
or U22649 (N_22649,N_22145,N_21942);
and U22650 (N_22650,N_21806,N_21974);
nor U22651 (N_22651,N_22184,N_21833);
nor U22652 (N_22652,N_22089,N_22169);
and U22653 (N_22653,N_21790,N_22071);
nand U22654 (N_22654,N_22154,N_21934);
nor U22655 (N_22655,N_21890,N_22157);
or U22656 (N_22656,N_21741,N_22022);
and U22657 (N_22657,N_21764,N_22041);
and U22658 (N_22658,N_21994,N_22161);
nand U22659 (N_22659,N_22084,N_21766);
nand U22660 (N_22660,N_21943,N_21705);
nor U22661 (N_22661,N_21860,N_22028);
or U22662 (N_22662,N_21752,N_22117);
nand U22663 (N_22663,N_21864,N_21927);
and U22664 (N_22664,N_22095,N_21639);
and U22665 (N_22665,N_22039,N_21790);
nor U22666 (N_22666,N_21982,N_21762);
nor U22667 (N_22667,N_21727,N_21893);
nor U22668 (N_22668,N_21918,N_21626);
nand U22669 (N_22669,N_22081,N_22179);
nor U22670 (N_22670,N_22083,N_21715);
nor U22671 (N_22671,N_21864,N_22136);
and U22672 (N_22672,N_21842,N_22042);
or U22673 (N_22673,N_22195,N_21804);
nor U22674 (N_22674,N_21962,N_22191);
xnor U22675 (N_22675,N_22019,N_22011);
and U22676 (N_22676,N_21809,N_22049);
nand U22677 (N_22677,N_22116,N_21636);
nand U22678 (N_22678,N_21911,N_21828);
and U22679 (N_22679,N_22129,N_21890);
xnor U22680 (N_22680,N_21835,N_22158);
nand U22681 (N_22681,N_21907,N_21851);
or U22682 (N_22682,N_21980,N_21884);
nand U22683 (N_22683,N_22091,N_22034);
nor U22684 (N_22684,N_21922,N_21698);
xor U22685 (N_22685,N_21836,N_21647);
nand U22686 (N_22686,N_21787,N_21658);
or U22687 (N_22687,N_21786,N_21673);
xnor U22688 (N_22688,N_21886,N_22088);
xor U22689 (N_22689,N_21694,N_21688);
xor U22690 (N_22690,N_21699,N_21858);
or U22691 (N_22691,N_21909,N_21656);
nor U22692 (N_22692,N_22054,N_21918);
nand U22693 (N_22693,N_22002,N_22077);
and U22694 (N_22694,N_21814,N_22077);
or U22695 (N_22695,N_22047,N_21932);
or U22696 (N_22696,N_21798,N_21636);
nor U22697 (N_22697,N_21884,N_21792);
and U22698 (N_22698,N_22097,N_22094);
nor U22699 (N_22699,N_22146,N_21601);
and U22700 (N_22700,N_21644,N_21866);
and U22701 (N_22701,N_21873,N_22119);
and U22702 (N_22702,N_21946,N_21731);
xnor U22703 (N_22703,N_21927,N_22187);
xor U22704 (N_22704,N_22134,N_22138);
xnor U22705 (N_22705,N_21841,N_21990);
nand U22706 (N_22706,N_22187,N_22190);
nand U22707 (N_22707,N_22109,N_22053);
xor U22708 (N_22708,N_21617,N_21911);
nor U22709 (N_22709,N_21877,N_21818);
xor U22710 (N_22710,N_21634,N_21999);
xor U22711 (N_22711,N_22096,N_21877);
nand U22712 (N_22712,N_22003,N_22149);
xnor U22713 (N_22713,N_21888,N_21788);
nor U22714 (N_22714,N_21811,N_21620);
and U22715 (N_22715,N_21616,N_22009);
nand U22716 (N_22716,N_21957,N_22126);
xor U22717 (N_22717,N_21869,N_21897);
or U22718 (N_22718,N_21899,N_21968);
nor U22719 (N_22719,N_21661,N_22125);
nand U22720 (N_22720,N_22007,N_21797);
nor U22721 (N_22721,N_21993,N_21628);
or U22722 (N_22722,N_22177,N_22197);
xor U22723 (N_22723,N_21706,N_22183);
and U22724 (N_22724,N_22043,N_21835);
and U22725 (N_22725,N_22173,N_22175);
or U22726 (N_22726,N_21935,N_21743);
xor U22727 (N_22727,N_21723,N_22091);
nor U22728 (N_22728,N_21986,N_22066);
nand U22729 (N_22729,N_21819,N_21857);
or U22730 (N_22730,N_21873,N_21739);
xor U22731 (N_22731,N_22082,N_21928);
xor U22732 (N_22732,N_22118,N_22089);
nand U22733 (N_22733,N_21665,N_22034);
xnor U22734 (N_22734,N_21839,N_21733);
nor U22735 (N_22735,N_22176,N_21746);
and U22736 (N_22736,N_21804,N_21990);
or U22737 (N_22737,N_21672,N_21655);
or U22738 (N_22738,N_22007,N_22147);
and U22739 (N_22739,N_21872,N_22189);
nor U22740 (N_22740,N_22139,N_22060);
xnor U22741 (N_22741,N_21865,N_21786);
nand U22742 (N_22742,N_21634,N_21845);
or U22743 (N_22743,N_22054,N_21870);
and U22744 (N_22744,N_22154,N_21645);
xor U22745 (N_22745,N_22040,N_22045);
nor U22746 (N_22746,N_21707,N_22000);
and U22747 (N_22747,N_22098,N_21865);
nand U22748 (N_22748,N_22066,N_22136);
and U22749 (N_22749,N_21834,N_22095);
or U22750 (N_22750,N_21621,N_21927);
and U22751 (N_22751,N_21644,N_22071);
nor U22752 (N_22752,N_21836,N_21666);
nor U22753 (N_22753,N_21857,N_21924);
or U22754 (N_22754,N_21697,N_21856);
or U22755 (N_22755,N_21839,N_21626);
or U22756 (N_22756,N_21867,N_21753);
nor U22757 (N_22757,N_21889,N_22066);
xor U22758 (N_22758,N_21637,N_22170);
nor U22759 (N_22759,N_21789,N_21639);
xnor U22760 (N_22760,N_21991,N_21895);
nand U22761 (N_22761,N_22090,N_21650);
nand U22762 (N_22762,N_21728,N_22107);
and U22763 (N_22763,N_21930,N_21681);
and U22764 (N_22764,N_22152,N_21842);
xnor U22765 (N_22765,N_21916,N_22046);
and U22766 (N_22766,N_22010,N_21662);
xnor U22767 (N_22767,N_21884,N_21632);
or U22768 (N_22768,N_22069,N_21668);
nor U22769 (N_22769,N_21990,N_21604);
nand U22770 (N_22770,N_21729,N_22189);
xnor U22771 (N_22771,N_21934,N_21701);
or U22772 (N_22772,N_21990,N_21639);
nor U22773 (N_22773,N_21996,N_21880);
xnor U22774 (N_22774,N_21740,N_21826);
nand U22775 (N_22775,N_21994,N_21995);
nor U22776 (N_22776,N_21858,N_22101);
nand U22777 (N_22777,N_22076,N_21602);
nor U22778 (N_22778,N_21991,N_22098);
and U22779 (N_22779,N_21881,N_22194);
nand U22780 (N_22780,N_21670,N_21974);
nor U22781 (N_22781,N_21673,N_21942);
or U22782 (N_22782,N_21999,N_21842);
nand U22783 (N_22783,N_22118,N_21898);
xnor U22784 (N_22784,N_21969,N_22015);
xor U22785 (N_22785,N_21792,N_22049);
xor U22786 (N_22786,N_22146,N_21702);
xnor U22787 (N_22787,N_21634,N_21873);
nand U22788 (N_22788,N_21888,N_21989);
xor U22789 (N_22789,N_21786,N_21623);
or U22790 (N_22790,N_22195,N_21868);
nand U22791 (N_22791,N_21747,N_22113);
or U22792 (N_22792,N_21856,N_21838);
or U22793 (N_22793,N_22067,N_21834);
and U22794 (N_22794,N_21673,N_21901);
nand U22795 (N_22795,N_22056,N_21617);
and U22796 (N_22796,N_22033,N_21682);
or U22797 (N_22797,N_22032,N_21651);
or U22798 (N_22798,N_21667,N_22029);
xnor U22799 (N_22799,N_21998,N_21947);
nand U22800 (N_22800,N_22295,N_22652);
and U22801 (N_22801,N_22622,N_22748);
xor U22802 (N_22802,N_22441,N_22722);
xnor U22803 (N_22803,N_22342,N_22494);
nand U22804 (N_22804,N_22493,N_22485);
xnor U22805 (N_22805,N_22238,N_22796);
nor U22806 (N_22806,N_22336,N_22627);
nor U22807 (N_22807,N_22705,N_22793);
nor U22808 (N_22808,N_22603,N_22708);
nor U22809 (N_22809,N_22713,N_22791);
xnor U22810 (N_22810,N_22432,N_22241);
nor U22811 (N_22811,N_22205,N_22778);
and U22812 (N_22812,N_22512,N_22765);
xnor U22813 (N_22813,N_22224,N_22730);
and U22814 (N_22814,N_22332,N_22222);
or U22815 (N_22815,N_22741,N_22363);
and U22816 (N_22816,N_22264,N_22663);
xor U22817 (N_22817,N_22607,N_22479);
or U22818 (N_22818,N_22292,N_22357);
or U22819 (N_22819,N_22310,N_22235);
xnor U22820 (N_22820,N_22592,N_22661);
xor U22821 (N_22821,N_22434,N_22243);
nor U22822 (N_22822,N_22341,N_22377);
nand U22823 (N_22823,N_22714,N_22490);
and U22824 (N_22824,N_22369,N_22328);
nor U22825 (N_22825,N_22788,N_22526);
nand U22826 (N_22826,N_22385,N_22619);
or U22827 (N_22827,N_22448,N_22496);
xor U22828 (N_22828,N_22734,N_22431);
nand U22829 (N_22829,N_22305,N_22501);
nand U22830 (N_22830,N_22462,N_22777);
xor U22831 (N_22831,N_22384,N_22257);
or U22832 (N_22832,N_22306,N_22252);
xnor U22833 (N_22833,N_22206,N_22267);
or U22834 (N_22834,N_22260,N_22312);
nand U22835 (N_22835,N_22261,N_22633);
xnor U22836 (N_22836,N_22231,N_22263);
nand U22837 (N_22837,N_22348,N_22303);
or U22838 (N_22838,N_22254,N_22591);
and U22839 (N_22839,N_22474,N_22459);
xnor U22840 (N_22840,N_22737,N_22736);
or U22841 (N_22841,N_22239,N_22425);
nand U22842 (N_22842,N_22611,N_22707);
nand U22843 (N_22843,N_22350,N_22368);
or U22844 (N_22844,N_22686,N_22318);
and U22845 (N_22845,N_22287,N_22645);
or U22846 (N_22846,N_22745,N_22383);
nand U22847 (N_22847,N_22540,N_22609);
xor U22848 (N_22848,N_22691,N_22776);
and U22849 (N_22849,N_22402,N_22487);
nand U22850 (N_22850,N_22249,N_22687);
nor U22851 (N_22851,N_22314,N_22509);
and U22852 (N_22852,N_22207,N_22789);
nor U22853 (N_22853,N_22542,N_22209);
nor U22854 (N_22854,N_22416,N_22420);
and U22855 (N_22855,N_22760,N_22505);
and U22856 (N_22856,N_22309,N_22334);
nand U22857 (N_22857,N_22375,N_22770);
nand U22858 (N_22858,N_22571,N_22262);
or U22859 (N_22859,N_22772,N_22757);
or U22860 (N_22860,N_22221,N_22506);
or U22861 (N_22861,N_22654,N_22530);
nor U22862 (N_22862,N_22316,N_22297);
nand U22863 (N_22863,N_22213,N_22755);
or U22864 (N_22864,N_22531,N_22541);
or U22865 (N_22865,N_22629,N_22732);
or U22866 (N_22866,N_22701,N_22638);
and U22867 (N_22867,N_22492,N_22338);
xnor U22868 (N_22868,N_22331,N_22756);
nand U22869 (N_22869,N_22277,N_22658);
or U22870 (N_22870,N_22300,N_22411);
or U22871 (N_22871,N_22486,N_22565);
and U22872 (N_22872,N_22299,N_22408);
nor U22873 (N_22873,N_22573,N_22202);
xnor U22874 (N_22874,N_22449,N_22751);
xnor U22875 (N_22875,N_22397,N_22326);
or U22876 (N_22876,N_22259,N_22547);
or U22877 (N_22877,N_22698,N_22325);
and U22878 (N_22878,N_22696,N_22344);
and U22879 (N_22879,N_22229,N_22453);
nand U22880 (N_22880,N_22604,N_22747);
nand U22881 (N_22881,N_22394,N_22373);
or U22882 (N_22882,N_22475,N_22504);
xnor U22883 (N_22883,N_22739,N_22489);
or U22884 (N_22884,N_22409,N_22595);
or U22885 (N_22885,N_22483,N_22673);
nand U22886 (N_22886,N_22551,N_22232);
or U22887 (N_22887,N_22532,N_22216);
or U22888 (N_22888,N_22293,N_22616);
nand U22889 (N_22889,N_22343,N_22354);
and U22890 (N_22890,N_22218,N_22517);
xor U22891 (N_22891,N_22644,N_22525);
or U22892 (N_22892,N_22689,N_22403);
nor U22893 (N_22893,N_22270,N_22269);
nand U22894 (N_22894,N_22587,N_22700);
or U22895 (N_22895,N_22352,N_22330);
xnor U22896 (N_22896,N_22567,N_22337);
nor U22897 (N_22897,N_22641,N_22605);
and U22898 (N_22898,N_22726,N_22598);
or U22899 (N_22899,N_22217,N_22718);
and U22900 (N_22900,N_22214,N_22563);
xnor U22901 (N_22901,N_22539,N_22680);
and U22902 (N_22902,N_22301,N_22203);
xnor U22903 (N_22903,N_22323,N_22291);
nor U22904 (N_22904,N_22422,N_22313);
xnor U22905 (N_22905,N_22568,N_22647);
nand U22906 (N_22906,N_22750,N_22690);
nand U22907 (N_22907,N_22358,N_22455);
and U22908 (N_22908,N_22784,N_22290);
or U22909 (N_22909,N_22639,N_22400);
nor U22910 (N_22910,N_22543,N_22457);
xnor U22911 (N_22911,N_22444,N_22642);
and U22912 (N_22912,N_22401,N_22464);
xnor U22913 (N_22913,N_22398,N_22588);
xor U22914 (N_22914,N_22271,N_22781);
or U22915 (N_22915,N_22364,N_22439);
nor U22916 (N_22916,N_22681,N_22423);
or U22917 (N_22917,N_22307,N_22227);
and U22918 (N_22918,N_22201,N_22637);
or U22919 (N_22919,N_22589,N_22792);
xor U22920 (N_22920,N_22692,N_22365);
xnor U22921 (N_22921,N_22442,N_22549);
xor U22922 (N_22922,N_22507,N_22623);
nand U22923 (N_22923,N_22446,N_22552);
nor U22924 (N_22924,N_22215,N_22669);
nor U22925 (N_22925,N_22349,N_22586);
nand U22926 (N_22926,N_22766,N_22615);
and U22927 (N_22927,N_22665,N_22674);
nand U22928 (N_22928,N_22621,N_22664);
xnor U22929 (N_22929,N_22245,N_22631);
xnor U22930 (N_22930,N_22635,N_22582);
and U22931 (N_22931,N_22450,N_22790);
or U22932 (N_22932,N_22454,N_22225);
xor U22933 (N_22933,N_22676,N_22360);
nand U22934 (N_22934,N_22522,N_22780);
and U22935 (N_22935,N_22711,N_22570);
xor U22936 (N_22936,N_22728,N_22361);
and U22937 (N_22937,N_22347,N_22284);
nand U22938 (N_22938,N_22626,N_22799);
nor U22939 (N_22939,N_22721,N_22406);
nor U22940 (N_22940,N_22426,N_22302);
and U22941 (N_22941,N_22510,N_22561);
and U22942 (N_22942,N_22514,N_22666);
nor U22943 (N_22943,N_22733,N_22572);
or U22944 (N_22944,N_22678,N_22695);
xnor U22945 (N_22945,N_22304,N_22795);
or U22946 (N_22946,N_22610,N_22550);
xor U22947 (N_22947,N_22421,N_22283);
nand U22948 (N_22948,N_22743,N_22502);
and U22949 (N_22949,N_22559,N_22646);
and U22950 (N_22950,N_22240,N_22286);
nor U22951 (N_22951,N_22440,N_22590);
nand U22952 (N_22952,N_22579,N_22407);
nor U22953 (N_22953,N_22472,N_22508);
nand U22954 (N_22954,N_22768,N_22351);
nor U22955 (N_22955,N_22353,N_22655);
and U22956 (N_22956,N_22410,N_22497);
nor U22957 (N_22957,N_22702,N_22597);
or U22958 (N_22958,N_22473,N_22761);
and U22959 (N_22959,N_22537,N_22329);
nand U22960 (N_22960,N_22463,N_22767);
and U22961 (N_22961,N_22296,N_22576);
nand U22962 (N_22962,N_22771,N_22482);
nand U22963 (N_22963,N_22324,N_22211);
nor U22964 (N_22964,N_22320,N_22618);
nor U22965 (N_22965,N_22758,N_22534);
nand U22966 (N_22966,N_22560,N_22716);
and U22967 (N_22967,N_22613,N_22725);
nand U22968 (N_22968,N_22569,N_22548);
xnor U22969 (N_22969,N_22285,N_22258);
xnor U22970 (N_22970,N_22729,N_22220);
and U22971 (N_22971,N_22624,N_22787);
xnor U22972 (N_22972,N_22513,N_22581);
and U22973 (N_22973,N_22774,N_22500);
nor U22974 (N_22974,N_22226,N_22430);
nor U22975 (N_22975,N_22317,N_22578);
nand U22976 (N_22976,N_22451,N_22273);
and U22977 (N_22977,N_22461,N_22367);
and U22978 (N_22978,N_22608,N_22738);
and U22979 (N_22979,N_22685,N_22424);
nand U22980 (N_22980,N_22276,N_22387);
and U22981 (N_22981,N_22339,N_22556);
nand U22982 (N_22982,N_22436,N_22580);
nand U22983 (N_22983,N_22679,N_22744);
or U22984 (N_22984,N_22554,N_22632);
and U22985 (N_22985,N_22288,N_22251);
nand U22986 (N_22986,N_22404,N_22742);
nor U22987 (N_22987,N_22653,N_22694);
or U22988 (N_22988,N_22699,N_22763);
nor U22989 (N_22989,N_22566,N_22520);
xor U22990 (N_22990,N_22445,N_22280);
nand U22991 (N_22991,N_22391,N_22465);
xnor U22992 (N_22992,N_22200,N_22650);
xor U22993 (N_22993,N_22355,N_22753);
or U22994 (N_22994,N_22553,N_22672);
or U22995 (N_22995,N_22256,N_22390);
nor U22996 (N_22996,N_22278,N_22417);
nor U22997 (N_22997,N_22783,N_22319);
and U22998 (N_22998,N_22555,N_22706);
nand U22999 (N_22999,N_22519,N_22315);
and U23000 (N_23000,N_22242,N_22266);
and U23001 (N_23001,N_22333,N_22779);
or U23002 (N_23002,N_22533,N_22775);
or U23003 (N_23003,N_22557,N_22575);
xnor U23004 (N_23004,N_22460,N_22370);
xor U23005 (N_23005,N_22498,N_22544);
nand U23006 (N_23006,N_22412,N_22723);
nand U23007 (N_23007,N_22253,N_22298);
nand U23008 (N_23008,N_22628,N_22740);
xor U23009 (N_23009,N_22662,N_22727);
xnor U23010 (N_23010,N_22405,N_22670);
nand U23011 (N_23011,N_22683,N_22447);
nand U23012 (N_23012,N_22527,N_22389);
nor U23013 (N_23013,N_22456,N_22491);
nor U23014 (N_23014,N_22558,N_22746);
nand U23015 (N_23015,N_22643,N_22668);
xnor U23016 (N_23016,N_22602,N_22660);
nor U23017 (N_23017,N_22378,N_22798);
nand U23018 (N_23018,N_22709,N_22467);
and U23019 (N_23019,N_22396,N_22675);
xnor U23020 (N_23020,N_22428,N_22617);
or U23021 (N_23021,N_22515,N_22593);
xnor U23022 (N_23022,N_22419,N_22773);
or U23023 (N_23023,N_22393,N_22414);
or U23024 (N_23024,N_22667,N_22246);
xnor U23025 (N_23025,N_22562,N_22659);
nor U23026 (N_23026,N_22786,N_22268);
nand U23027 (N_23027,N_22599,N_22585);
nand U23028 (N_23028,N_22236,N_22371);
nor U23029 (N_23029,N_22495,N_22764);
and U23030 (N_23030,N_22247,N_22648);
or U23031 (N_23031,N_22470,N_22712);
nor U23032 (N_23032,N_22523,N_22794);
nor U23033 (N_23033,N_22469,N_22749);
and U23034 (N_23034,N_22308,N_22415);
nor U23035 (N_23035,N_22208,N_22596);
nand U23036 (N_23036,N_22265,N_22433);
nor U23037 (N_23037,N_22477,N_22468);
xor U23038 (N_23038,N_22335,N_22345);
nor U23039 (N_23039,N_22379,N_22503);
or U23040 (N_23040,N_22640,N_22584);
and U23041 (N_23041,N_22294,N_22356);
xnor U23042 (N_23042,N_22657,N_22374);
nand U23043 (N_23043,N_22471,N_22340);
and U23044 (N_23044,N_22762,N_22731);
xnor U23045 (N_23045,N_22656,N_22583);
or U23046 (N_23046,N_22372,N_22466);
nor U23047 (N_23047,N_22322,N_22545);
nand U23048 (N_23048,N_22594,N_22684);
xor U23049 (N_23049,N_22388,N_22429);
and U23050 (N_23050,N_22634,N_22476);
nand U23051 (N_23051,N_22219,N_22418);
and U23052 (N_23052,N_22359,N_22735);
and U23053 (N_23053,N_22289,N_22516);
xnor U23054 (N_23054,N_22272,N_22311);
xnor U23055 (N_23055,N_22577,N_22204);
xor U23056 (N_23056,N_22717,N_22480);
xor U23057 (N_23057,N_22250,N_22248);
or U23058 (N_23058,N_22443,N_22636);
nor U23059 (N_23059,N_22703,N_22230);
and U23060 (N_23060,N_22536,N_22435);
or U23061 (N_23061,N_22528,N_22710);
and U23062 (N_23062,N_22274,N_22228);
xnor U23063 (N_23063,N_22759,N_22321);
nand U23064 (N_23064,N_22529,N_22499);
xor U23065 (N_23065,N_22769,N_22521);
or U23066 (N_23066,N_22693,N_22399);
and U23067 (N_23067,N_22606,N_22518);
nand U23068 (N_23068,N_22614,N_22437);
nor U23069 (N_23069,N_22630,N_22382);
xor U23070 (N_23070,N_22386,N_22682);
nor U23071 (N_23071,N_22380,N_22327);
xnor U23072 (N_23072,N_22688,N_22376);
and U23073 (N_23073,N_22546,N_22210);
and U23074 (N_23074,N_22719,N_22237);
and U23075 (N_23075,N_22511,N_22715);
nand U23076 (N_23076,N_22478,N_22244);
and U23077 (N_23077,N_22724,N_22275);
or U23078 (N_23078,N_22395,N_22797);
nor U23079 (N_23079,N_22782,N_22234);
nor U23080 (N_23080,N_22413,N_22785);
nand U23081 (N_23081,N_22279,N_22704);
and U23082 (N_23082,N_22381,N_22255);
nand U23083 (N_23083,N_22600,N_22697);
or U23084 (N_23084,N_22481,N_22752);
nand U23085 (N_23085,N_22488,N_22677);
xnor U23086 (N_23086,N_22281,N_22212);
nand U23087 (N_23087,N_22458,N_22620);
nor U23088 (N_23088,N_22223,N_22427);
or U23089 (N_23089,N_22538,N_22720);
or U23090 (N_23090,N_22392,N_22535);
nand U23091 (N_23091,N_22574,N_22601);
nand U23092 (N_23092,N_22282,N_22754);
xnor U23093 (N_23093,N_22452,N_22362);
nand U23094 (N_23094,N_22233,N_22524);
and U23095 (N_23095,N_22564,N_22438);
and U23096 (N_23096,N_22484,N_22346);
xnor U23097 (N_23097,N_22625,N_22366);
xor U23098 (N_23098,N_22671,N_22651);
or U23099 (N_23099,N_22612,N_22649);
or U23100 (N_23100,N_22419,N_22576);
nand U23101 (N_23101,N_22249,N_22441);
or U23102 (N_23102,N_22274,N_22414);
and U23103 (N_23103,N_22573,N_22420);
nand U23104 (N_23104,N_22652,N_22364);
nor U23105 (N_23105,N_22337,N_22302);
or U23106 (N_23106,N_22474,N_22204);
and U23107 (N_23107,N_22408,N_22241);
nand U23108 (N_23108,N_22773,N_22657);
and U23109 (N_23109,N_22449,N_22633);
nor U23110 (N_23110,N_22328,N_22285);
and U23111 (N_23111,N_22708,N_22529);
xor U23112 (N_23112,N_22396,N_22428);
xnor U23113 (N_23113,N_22560,N_22400);
and U23114 (N_23114,N_22726,N_22506);
or U23115 (N_23115,N_22513,N_22524);
nand U23116 (N_23116,N_22598,N_22556);
nand U23117 (N_23117,N_22657,N_22402);
nor U23118 (N_23118,N_22532,N_22485);
nor U23119 (N_23119,N_22492,N_22362);
nand U23120 (N_23120,N_22498,N_22471);
nand U23121 (N_23121,N_22451,N_22721);
or U23122 (N_23122,N_22458,N_22481);
nand U23123 (N_23123,N_22355,N_22565);
nand U23124 (N_23124,N_22620,N_22421);
nor U23125 (N_23125,N_22407,N_22530);
and U23126 (N_23126,N_22575,N_22363);
xor U23127 (N_23127,N_22534,N_22730);
nor U23128 (N_23128,N_22405,N_22387);
and U23129 (N_23129,N_22663,N_22233);
xnor U23130 (N_23130,N_22507,N_22735);
and U23131 (N_23131,N_22350,N_22540);
nor U23132 (N_23132,N_22378,N_22394);
or U23133 (N_23133,N_22645,N_22407);
xnor U23134 (N_23134,N_22714,N_22767);
or U23135 (N_23135,N_22222,N_22659);
nor U23136 (N_23136,N_22259,N_22618);
nand U23137 (N_23137,N_22241,N_22687);
and U23138 (N_23138,N_22449,N_22434);
xor U23139 (N_23139,N_22275,N_22717);
nor U23140 (N_23140,N_22474,N_22361);
and U23141 (N_23141,N_22559,N_22664);
xor U23142 (N_23142,N_22558,N_22305);
xor U23143 (N_23143,N_22326,N_22741);
or U23144 (N_23144,N_22468,N_22312);
nand U23145 (N_23145,N_22398,N_22775);
xnor U23146 (N_23146,N_22771,N_22289);
xor U23147 (N_23147,N_22745,N_22207);
or U23148 (N_23148,N_22224,N_22617);
nand U23149 (N_23149,N_22728,N_22398);
or U23150 (N_23150,N_22567,N_22341);
or U23151 (N_23151,N_22778,N_22784);
or U23152 (N_23152,N_22684,N_22674);
nor U23153 (N_23153,N_22529,N_22301);
or U23154 (N_23154,N_22655,N_22688);
nand U23155 (N_23155,N_22240,N_22529);
or U23156 (N_23156,N_22639,N_22336);
or U23157 (N_23157,N_22549,N_22469);
xnor U23158 (N_23158,N_22533,N_22282);
or U23159 (N_23159,N_22756,N_22740);
nor U23160 (N_23160,N_22401,N_22350);
and U23161 (N_23161,N_22605,N_22556);
or U23162 (N_23162,N_22730,N_22647);
nor U23163 (N_23163,N_22669,N_22317);
xor U23164 (N_23164,N_22487,N_22523);
xnor U23165 (N_23165,N_22443,N_22742);
nor U23166 (N_23166,N_22440,N_22518);
nor U23167 (N_23167,N_22262,N_22690);
and U23168 (N_23168,N_22355,N_22220);
and U23169 (N_23169,N_22421,N_22672);
and U23170 (N_23170,N_22718,N_22201);
and U23171 (N_23171,N_22278,N_22717);
nand U23172 (N_23172,N_22210,N_22246);
nand U23173 (N_23173,N_22607,N_22413);
nor U23174 (N_23174,N_22619,N_22698);
or U23175 (N_23175,N_22612,N_22405);
xnor U23176 (N_23176,N_22293,N_22545);
and U23177 (N_23177,N_22451,N_22682);
xnor U23178 (N_23178,N_22309,N_22432);
xor U23179 (N_23179,N_22331,N_22460);
or U23180 (N_23180,N_22732,N_22535);
xor U23181 (N_23181,N_22266,N_22293);
and U23182 (N_23182,N_22665,N_22209);
xnor U23183 (N_23183,N_22418,N_22639);
nand U23184 (N_23184,N_22344,N_22607);
nand U23185 (N_23185,N_22239,N_22458);
or U23186 (N_23186,N_22239,N_22516);
xnor U23187 (N_23187,N_22445,N_22453);
xnor U23188 (N_23188,N_22271,N_22797);
or U23189 (N_23189,N_22543,N_22633);
nor U23190 (N_23190,N_22619,N_22363);
xnor U23191 (N_23191,N_22352,N_22341);
nor U23192 (N_23192,N_22408,N_22780);
nor U23193 (N_23193,N_22458,N_22582);
and U23194 (N_23194,N_22783,N_22231);
nand U23195 (N_23195,N_22545,N_22281);
nor U23196 (N_23196,N_22687,N_22232);
nand U23197 (N_23197,N_22294,N_22439);
nor U23198 (N_23198,N_22373,N_22676);
nor U23199 (N_23199,N_22573,N_22515);
and U23200 (N_23200,N_22690,N_22710);
and U23201 (N_23201,N_22272,N_22457);
or U23202 (N_23202,N_22742,N_22382);
xor U23203 (N_23203,N_22324,N_22249);
nor U23204 (N_23204,N_22304,N_22507);
nand U23205 (N_23205,N_22750,N_22480);
and U23206 (N_23206,N_22474,N_22390);
nand U23207 (N_23207,N_22710,N_22295);
nand U23208 (N_23208,N_22228,N_22507);
and U23209 (N_23209,N_22713,N_22303);
nor U23210 (N_23210,N_22262,N_22354);
or U23211 (N_23211,N_22581,N_22680);
nor U23212 (N_23212,N_22358,N_22243);
xor U23213 (N_23213,N_22686,N_22475);
or U23214 (N_23214,N_22746,N_22353);
or U23215 (N_23215,N_22791,N_22513);
or U23216 (N_23216,N_22743,N_22340);
and U23217 (N_23217,N_22388,N_22340);
xnor U23218 (N_23218,N_22499,N_22793);
and U23219 (N_23219,N_22227,N_22613);
or U23220 (N_23220,N_22208,N_22617);
and U23221 (N_23221,N_22730,N_22393);
nand U23222 (N_23222,N_22214,N_22474);
or U23223 (N_23223,N_22407,N_22511);
or U23224 (N_23224,N_22763,N_22446);
or U23225 (N_23225,N_22200,N_22472);
or U23226 (N_23226,N_22207,N_22288);
nand U23227 (N_23227,N_22428,N_22229);
or U23228 (N_23228,N_22243,N_22617);
xor U23229 (N_23229,N_22622,N_22523);
nand U23230 (N_23230,N_22302,N_22613);
and U23231 (N_23231,N_22594,N_22578);
nor U23232 (N_23232,N_22369,N_22300);
nor U23233 (N_23233,N_22593,N_22479);
and U23234 (N_23234,N_22718,N_22549);
and U23235 (N_23235,N_22367,N_22659);
xnor U23236 (N_23236,N_22465,N_22760);
or U23237 (N_23237,N_22737,N_22748);
or U23238 (N_23238,N_22607,N_22540);
xnor U23239 (N_23239,N_22615,N_22796);
xnor U23240 (N_23240,N_22207,N_22494);
nand U23241 (N_23241,N_22682,N_22511);
and U23242 (N_23242,N_22778,N_22659);
or U23243 (N_23243,N_22598,N_22411);
nor U23244 (N_23244,N_22397,N_22746);
or U23245 (N_23245,N_22718,N_22724);
or U23246 (N_23246,N_22613,N_22519);
nor U23247 (N_23247,N_22492,N_22516);
xor U23248 (N_23248,N_22586,N_22736);
nand U23249 (N_23249,N_22613,N_22683);
xnor U23250 (N_23250,N_22738,N_22649);
or U23251 (N_23251,N_22450,N_22366);
or U23252 (N_23252,N_22269,N_22258);
nand U23253 (N_23253,N_22773,N_22716);
or U23254 (N_23254,N_22725,N_22383);
nand U23255 (N_23255,N_22224,N_22498);
nand U23256 (N_23256,N_22348,N_22270);
or U23257 (N_23257,N_22218,N_22732);
and U23258 (N_23258,N_22618,N_22223);
nor U23259 (N_23259,N_22539,N_22623);
xor U23260 (N_23260,N_22381,N_22464);
xor U23261 (N_23261,N_22501,N_22626);
nor U23262 (N_23262,N_22532,N_22415);
or U23263 (N_23263,N_22297,N_22425);
nand U23264 (N_23264,N_22653,N_22417);
nor U23265 (N_23265,N_22615,N_22330);
xnor U23266 (N_23266,N_22597,N_22471);
nor U23267 (N_23267,N_22737,N_22790);
nand U23268 (N_23268,N_22468,N_22269);
and U23269 (N_23269,N_22526,N_22438);
and U23270 (N_23270,N_22792,N_22267);
xor U23271 (N_23271,N_22649,N_22797);
nor U23272 (N_23272,N_22441,N_22404);
xor U23273 (N_23273,N_22400,N_22350);
xnor U23274 (N_23274,N_22373,N_22686);
nor U23275 (N_23275,N_22584,N_22771);
nor U23276 (N_23276,N_22785,N_22713);
xor U23277 (N_23277,N_22475,N_22431);
or U23278 (N_23278,N_22256,N_22213);
nor U23279 (N_23279,N_22255,N_22627);
or U23280 (N_23280,N_22314,N_22550);
nand U23281 (N_23281,N_22769,N_22508);
and U23282 (N_23282,N_22412,N_22527);
nand U23283 (N_23283,N_22583,N_22425);
nor U23284 (N_23284,N_22650,N_22471);
nand U23285 (N_23285,N_22618,N_22497);
nor U23286 (N_23286,N_22726,N_22788);
nand U23287 (N_23287,N_22777,N_22607);
xor U23288 (N_23288,N_22705,N_22374);
and U23289 (N_23289,N_22641,N_22309);
xor U23290 (N_23290,N_22313,N_22524);
nor U23291 (N_23291,N_22621,N_22557);
and U23292 (N_23292,N_22600,N_22407);
xor U23293 (N_23293,N_22471,N_22463);
or U23294 (N_23294,N_22739,N_22210);
nor U23295 (N_23295,N_22761,N_22601);
nor U23296 (N_23296,N_22224,N_22408);
nor U23297 (N_23297,N_22240,N_22347);
nor U23298 (N_23298,N_22351,N_22385);
nor U23299 (N_23299,N_22602,N_22207);
and U23300 (N_23300,N_22447,N_22690);
xor U23301 (N_23301,N_22733,N_22261);
or U23302 (N_23302,N_22683,N_22503);
and U23303 (N_23303,N_22234,N_22510);
and U23304 (N_23304,N_22227,N_22540);
xnor U23305 (N_23305,N_22773,N_22369);
nor U23306 (N_23306,N_22549,N_22721);
and U23307 (N_23307,N_22403,N_22730);
or U23308 (N_23308,N_22257,N_22385);
xnor U23309 (N_23309,N_22682,N_22302);
and U23310 (N_23310,N_22468,N_22684);
or U23311 (N_23311,N_22595,N_22639);
and U23312 (N_23312,N_22229,N_22529);
and U23313 (N_23313,N_22415,N_22342);
or U23314 (N_23314,N_22228,N_22790);
nor U23315 (N_23315,N_22428,N_22365);
xnor U23316 (N_23316,N_22434,N_22242);
xnor U23317 (N_23317,N_22471,N_22571);
nand U23318 (N_23318,N_22579,N_22696);
and U23319 (N_23319,N_22611,N_22346);
or U23320 (N_23320,N_22287,N_22630);
nor U23321 (N_23321,N_22776,N_22666);
nand U23322 (N_23322,N_22338,N_22273);
xnor U23323 (N_23323,N_22698,N_22514);
nand U23324 (N_23324,N_22746,N_22334);
xnor U23325 (N_23325,N_22791,N_22702);
nand U23326 (N_23326,N_22405,N_22470);
nand U23327 (N_23327,N_22479,N_22651);
xor U23328 (N_23328,N_22398,N_22201);
nor U23329 (N_23329,N_22434,N_22245);
xnor U23330 (N_23330,N_22730,N_22218);
xnor U23331 (N_23331,N_22420,N_22545);
and U23332 (N_23332,N_22267,N_22244);
nand U23333 (N_23333,N_22739,N_22652);
and U23334 (N_23334,N_22641,N_22482);
nand U23335 (N_23335,N_22711,N_22539);
nor U23336 (N_23336,N_22380,N_22204);
or U23337 (N_23337,N_22750,N_22719);
nand U23338 (N_23338,N_22203,N_22519);
nand U23339 (N_23339,N_22708,N_22775);
xnor U23340 (N_23340,N_22290,N_22515);
xnor U23341 (N_23341,N_22264,N_22504);
xnor U23342 (N_23342,N_22613,N_22537);
xnor U23343 (N_23343,N_22433,N_22624);
nand U23344 (N_23344,N_22412,N_22451);
nor U23345 (N_23345,N_22238,N_22209);
or U23346 (N_23346,N_22655,N_22212);
and U23347 (N_23347,N_22227,N_22645);
nor U23348 (N_23348,N_22404,N_22453);
and U23349 (N_23349,N_22642,N_22776);
xnor U23350 (N_23350,N_22679,N_22793);
xnor U23351 (N_23351,N_22231,N_22506);
nand U23352 (N_23352,N_22798,N_22232);
xor U23353 (N_23353,N_22773,N_22236);
nor U23354 (N_23354,N_22220,N_22486);
nand U23355 (N_23355,N_22773,N_22550);
nor U23356 (N_23356,N_22454,N_22781);
or U23357 (N_23357,N_22202,N_22582);
or U23358 (N_23358,N_22445,N_22369);
or U23359 (N_23359,N_22290,N_22734);
or U23360 (N_23360,N_22643,N_22526);
and U23361 (N_23361,N_22780,N_22620);
nor U23362 (N_23362,N_22500,N_22610);
and U23363 (N_23363,N_22254,N_22297);
nand U23364 (N_23364,N_22351,N_22389);
nand U23365 (N_23365,N_22216,N_22446);
or U23366 (N_23366,N_22546,N_22486);
nand U23367 (N_23367,N_22230,N_22295);
xor U23368 (N_23368,N_22446,N_22205);
or U23369 (N_23369,N_22308,N_22301);
and U23370 (N_23370,N_22634,N_22542);
nand U23371 (N_23371,N_22241,N_22558);
and U23372 (N_23372,N_22726,N_22264);
nand U23373 (N_23373,N_22717,N_22508);
and U23374 (N_23374,N_22469,N_22435);
nand U23375 (N_23375,N_22750,N_22629);
nor U23376 (N_23376,N_22354,N_22783);
nor U23377 (N_23377,N_22744,N_22317);
and U23378 (N_23378,N_22422,N_22629);
nand U23379 (N_23379,N_22784,N_22470);
or U23380 (N_23380,N_22608,N_22344);
and U23381 (N_23381,N_22490,N_22455);
or U23382 (N_23382,N_22459,N_22546);
nor U23383 (N_23383,N_22501,N_22547);
nand U23384 (N_23384,N_22479,N_22207);
nor U23385 (N_23385,N_22324,N_22359);
xnor U23386 (N_23386,N_22569,N_22706);
or U23387 (N_23387,N_22280,N_22426);
nand U23388 (N_23388,N_22248,N_22473);
or U23389 (N_23389,N_22541,N_22451);
xnor U23390 (N_23390,N_22522,N_22641);
and U23391 (N_23391,N_22329,N_22688);
and U23392 (N_23392,N_22331,N_22582);
xor U23393 (N_23393,N_22467,N_22575);
or U23394 (N_23394,N_22517,N_22271);
or U23395 (N_23395,N_22227,N_22421);
nor U23396 (N_23396,N_22241,N_22743);
nand U23397 (N_23397,N_22792,N_22540);
nand U23398 (N_23398,N_22628,N_22579);
or U23399 (N_23399,N_22420,N_22258);
nand U23400 (N_23400,N_23186,N_22978);
and U23401 (N_23401,N_22881,N_23165);
nand U23402 (N_23402,N_22885,N_23244);
xnor U23403 (N_23403,N_22846,N_23080);
or U23404 (N_23404,N_22803,N_23271);
and U23405 (N_23405,N_23129,N_23290);
xnor U23406 (N_23406,N_23176,N_23172);
and U23407 (N_23407,N_23027,N_23230);
or U23408 (N_23408,N_22998,N_22853);
nand U23409 (N_23409,N_22955,N_23082);
xor U23410 (N_23410,N_23277,N_23157);
or U23411 (N_23411,N_22960,N_22989);
xnor U23412 (N_23412,N_23064,N_23335);
and U23413 (N_23413,N_23096,N_23378);
nand U23414 (N_23414,N_22999,N_23089);
or U23415 (N_23415,N_23357,N_23353);
or U23416 (N_23416,N_22805,N_23133);
or U23417 (N_23417,N_23048,N_23368);
nand U23418 (N_23418,N_22867,N_23159);
nor U23419 (N_23419,N_23017,N_22858);
nand U23420 (N_23420,N_22876,N_23022);
nor U23421 (N_23421,N_23019,N_22893);
or U23422 (N_23422,N_23264,N_23347);
nor U23423 (N_23423,N_23262,N_22877);
or U23424 (N_23424,N_22872,N_23209);
and U23425 (N_23425,N_22828,N_23320);
or U23426 (N_23426,N_23128,N_22954);
and U23427 (N_23427,N_22871,N_23010);
or U23428 (N_23428,N_22890,N_23091);
nor U23429 (N_23429,N_22952,N_23310);
nor U23430 (N_23430,N_23203,N_23374);
xor U23431 (N_23431,N_22825,N_22953);
nand U23432 (N_23432,N_23325,N_23332);
nor U23433 (N_23433,N_23306,N_23126);
nor U23434 (N_23434,N_23127,N_22949);
nor U23435 (N_23435,N_23311,N_22830);
and U23436 (N_23436,N_23339,N_22892);
and U23437 (N_23437,N_23340,N_23235);
or U23438 (N_23438,N_23168,N_23386);
nor U23439 (N_23439,N_23196,N_23000);
xnor U23440 (N_23440,N_22884,N_22941);
nand U23441 (N_23441,N_22986,N_23355);
or U23442 (N_23442,N_22880,N_23121);
xor U23443 (N_23443,N_23143,N_22951);
and U23444 (N_23444,N_23314,N_23087);
xor U23445 (N_23445,N_22966,N_23372);
nand U23446 (N_23446,N_23327,N_22970);
xnor U23447 (N_23447,N_23063,N_23026);
nand U23448 (N_23448,N_22808,N_22901);
xor U23449 (N_23449,N_22802,N_22963);
nand U23450 (N_23450,N_23212,N_23289);
nand U23451 (N_23451,N_22866,N_23315);
or U23452 (N_23452,N_23199,N_23072);
xnor U23453 (N_23453,N_23173,N_22943);
nand U23454 (N_23454,N_23214,N_23057);
nand U23455 (N_23455,N_23399,N_22856);
xor U23456 (N_23456,N_23398,N_23276);
and U23457 (N_23457,N_23058,N_23253);
xnor U23458 (N_23458,N_23329,N_23179);
nor U23459 (N_23459,N_22944,N_23042);
or U23460 (N_23460,N_23393,N_23097);
and U23461 (N_23461,N_23170,N_23066);
xor U23462 (N_23462,N_23316,N_23202);
and U23463 (N_23463,N_23052,N_23060);
nand U23464 (N_23464,N_23260,N_23389);
and U23465 (N_23465,N_23115,N_22940);
nor U23466 (N_23466,N_23261,N_22860);
and U23467 (N_23467,N_23132,N_23308);
nand U23468 (N_23468,N_22815,N_22979);
and U23469 (N_23469,N_23231,N_23137);
and U23470 (N_23470,N_23365,N_22980);
or U23471 (N_23471,N_23041,N_23274);
and U23472 (N_23472,N_22813,N_23153);
nor U23473 (N_23473,N_23321,N_23148);
xnor U23474 (N_23474,N_22827,N_22801);
nand U23475 (N_23475,N_23191,N_23216);
nand U23476 (N_23476,N_22844,N_23384);
xor U23477 (N_23477,N_23160,N_23319);
or U23478 (N_23478,N_23279,N_23180);
xor U23479 (N_23479,N_23349,N_23013);
nor U23480 (N_23480,N_22982,N_22950);
nand U23481 (N_23481,N_23283,N_23050);
or U23482 (N_23482,N_22821,N_22946);
xnor U23483 (N_23483,N_22983,N_23217);
nand U23484 (N_23484,N_23004,N_23292);
and U23485 (N_23485,N_23051,N_22995);
nor U23486 (N_23486,N_22865,N_22832);
and U23487 (N_23487,N_22873,N_22956);
xor U23488 (N_23488,N_22967,N_23356);
nand U23489 (N_23489,N_22948,N_23229);
xor U23490 (N_23490,N_23171,N_22826);
xnor U23491 (N_23491,N_23198,N_22900);
and U23492 (N_23492,N_23123,N_23268);
and U23493 (N_23493,N_22863,N_23140);
xor U23494 (N_23494,N_23003,N_23341);
or U23495 (N_23495,N_23193,N_22907);
xnor U23496 (N_23496,N_23032,N_23323);
or U23497 (N_23497,N_23237,N_23383);
or U23498 (N_23498,N_23093,N_23059);
xor U23499 (N_23499,N_23055,N_22929);
xor U23500 (N_23500,N_22994,N_23364);
nor U23501 (N_23501,N_23256,N_23005);
xor U23502 (N_23502,N_23366,N_22973);
nor U23503 (N_23503,N_23102,N_23287);
nand U23504 (N_23504,N_22809,N_22938);
nor U23505 (N_23505,N_22895,N_23360);
or U23506 (N_23506,N_23088,N_22820);
or U23507 (N_23507,N_23324,N_23269);
nand U23508 (N_23508,N_22862,N_23252);
nand U23509 (N_23509,N_23358,N_23305);
nor U23510 (N_23510,N_23293,N_23309);
xor U23511 (N_23511,N_23039,N_23070);
nor U23512 (N_23512,N_23213,N_23164);
nand U23513 (N_23513,N_23377,N_22987);
and U23514 (N_23514,N_23385,N_22906);
nor U23515 (N_23515,N_23344,N_22812);
nor U23516 (N_23516,N_22857,N_23238);
and U23517 (N_23517,N_23257,N_22918);
or U23518 (N_23518,N_23151,N_22945);
xnor U23519 (N_23519,N_23215,N_22928);
or U23520 (N_23520,N_23286,N_23313);
nand U23521 (N_23521,N_23381,N_22972);
and U23522 (N_23522,N_23391,N_23034);
xnor U23523 (N_23523,N_23336,N_22975);
nor U23524 (N_23524,N_23208,N_22930);
nand U23525 (N_23525,N_23382,N_23330);
xnor U23526 (N_23526,N_23352,N_23219);
nand U23527 (N_23527,N_22915,N_23190);
nor U23528 (N_23528,N_23023,N_23317);
nor U23529 (N_23529,N_22855,N_23071);
or U23530 (N_23530,N_23192,N_23337);
nor U23531 (N_23531,N_23395,N_22990);
nand U23532 (N_23532,N_22839,N_22819);
nor U23533 (N_23533,N_22958,N_23134);
and U23534 (N_23534,N_23387,N_23218);
nor U23535 (N_23535,N_23099,N_22947);
xnor U23536 (N_23536,N_23079,N_23018);
or U23537 (N_23537,N_22854,N_23035);
xnor U23538 (N_23538,N_22838,N_22869);
nor U23539 (N_23539,N_23343,N_22902);
nand U23540 (N_23540,N_23009,N_23144);
nor U23541 (N_23541,N_23025,N_22816);
xor U23542 (N_23542,N_23396,N_23243);
xor U23543 (N_23543,N_23254,N_23334);
nor U23544 (N_23544,N_22957,N_23001);
or U23545 (N_23545,N_22926,N_23118);
nand U23546 (N_23546,N_22879,N_22977);
nand U23547 (N_23547,N_23105,N_22886);
nand U23548 (N_23548,N_22868,N_23187);
nor U23549 (N_23549,N_23224,N_22984);
nor U23550 (N_23550,N_23136,N_23322);
or U23551 (N_23551,N_23275,N_23211);
xor U23552 (N_23552,N_22914,N_23351);
xnor U23553 (N_23553,N_22837,N_22905);
nor U23554 (N_23554,N_22852,N_22919);
or U23555 (N_23555,N_23012,N_23234);
nand U23556 (N_23556,N_23006,N_22996);
or U23557 (N_23557,N_22814,N_23040);
and U23558 (N_23558,N_22997,N_22847);
nand U23559 (N_23559,N_23284,N_22903);
or U23560 (N_23560,N_23037,N_22933);
or U23561 (N_23561,N_22840,N_23201);
and U23562 (N_23562,N_23247,N_23109);
and U23563 (N_23563,N_22883,N_22806);
or U23564 (N_23564,N_23369,N_22848);
xnor U23565 (N_23565,N_23220,N_22937);
or U23566 (N_23566,N_23074,N_23248);
nand U23567 (N_23567,N_23104,N_22925);
nor U23568 (N_23568,N_23114,N_23146);
xnor U23569 (N_23569,N_23295,N_23255);
nand U23570 (N_23570,N_22969,N_23141);
and U23571 (N_23571,N_22991,N_22912);
xnor U23572 (N_23572,N_23086,N_23388);
xnor U23573 (N_23573,N_23204,N_23065);
nor U23574 (N_23574,N_22836,N_23246);
nor U23575 (N_23575,N_23241,N_22913);
or U23576 (N_23576,N_23033,N_23150);
and U23577 (N_23577,N_22807,N_23119);
and U23578 (N_23578,N_23043,N_23302);
or U23579 (N_23579,N_22824,N_23328);
xnor U23580 (N_23580,N_23110,N_23103);
nor U23581 (N_23581,N_23236,N_23166);
xor U23582 (N_23582,N_23038,N_22908);
and U23583 (N_23583,N_23162,N_23259);
nor U23584 (N_23584,N_23232,N_23200);
nor U23585 (N_23585,N_22896,N_22845);
or U23586 (N_23586,N_22942,N_22935);
xor U23587 (N_23587,N_22992,N_23116);
nand U23588 (N_23588,N_23251,N_23210);
xnor U23589 (N_23589,N_22899,N_23263);
and U23590 (N_23590,N_23167,N_23107);
nand U23591 (N_23591,N_23270,N_22974);
nor U23592 (N_23592,N_23194,N_23076);
nand U23593 (N_23593,N_22894,N_22817);
xnor U23594 (N_23594,N_22887,N_23177);
nor U23595 (N_23595,N_23161,N_22916);
or U23596 (N_23596,N_23233,N_23394);
nand U23597 (N_23597,N_23297,N_23081);
xnor U23598 (N_23598,N_22921,N_23067);
xor U23599 (N_23599,N_23338,N_23124);
and U23600 (N_23600,N_22843,N_23185);
or U23601 (N_23601,N_23367,N_22859);
xor U23602 (N_23602,N_23195,N_22924);
xnor U23603 (N_23603,N_23285,N_23296);
xnor U23604 (N_23604,N_23142,N_22841);
nor U23605 (N_23605,N_23112,N_23007);
xnor U23606 (N_23606,N_22818,N_23183);
nand U23607 (N_23607,N_23101,N_22861);
xnor U23608 (N_23608,N_23345,N_23073);
nor U23609 (N_23609,N_23045,N_23350);
nor U23610 (N_23610,N_22864,N_23371);
nand U23611 (N_23611,N_23375,N_23359);
nand U23612 (N_23612,N_23113,N_23361);
or U23613 (N_23613,N_23265,N_22931);
or U23614 (N_23614,N_23282,N_23291);
and U23615 (N_23615,N_22976,N_23226);
nand U23616 (N_23616,N_23028,N_23331);
and U23617 (N_23617,N_23207,N_23333);
xor U23618 (N_23618,N_22968,N_23300);
xor U23619 (N_23619,N_23249,N_22804);
nor U23620 (N_23620,N_23174,N_23002);
and U23621 (N_23621,N_23380,N_22875);
nand U23622 (N_23622,N_22927,N_23069);
nor U23623 (N_23623,N_22874,N_23149);
xnor U23624 (N_23624,N_23239,N_23354);
nor U23625 (N_23625,N_22842,N_23301);
nand U23626 (N_23626,N_23008,N_23280);
xor U23627 (N_23627,N_23266,N_23342);
xor U23628 (N_23628,N_23188,N_23077);
nor U23629 (N_23629,N_23181,N_23288);
or U23630 (N_23630,N_22870,N_23139);
nand U23631 (N_23631,N_23147,N_23130);
xor U23632 (N_23632,N_23131,N_23135);
nor U23633 (N_23633,N_23250,N_23054);
xor U23634 (N_23634,N_22923,N_23307);
or U23635 (N_23635,N_23222,N_23154);
or U23636 (N_23636,N_23011,N_22889);
or U23637 (N_23637,N_23175,N_23303);
or U23638 (N_23638,N_23245,N_23021);
xnor U23639 (N_23639,N_22934,N_22964);
nor U23640 (N_23640,N_23182,N_22829);
and U23641 (N_23641,N_22898,N_22800);
nand U23642 (N_23642,N_23084,N_23049);
or U23643 (N_23643,N_22897,N_23397);
or U23644 (N_23644,N_23145,N_23016);
xor U23645 (N_23645,N_23390,N_23029);
xor U23646 (N_23646,N_23163,N_22811);
xor U23647 (N_23647,N_23206,N_23221);
xor U23648 (N_23648,N_22833,N_22810);
nand U23649 (N_23649,N_22835,N_22822);
or U23650 (N_23650,N_23111,N_23083);
and U23651 (N_23651,N_23158,N_23169);
nor U23652 (N_23652,N_22985,N_22831);
and U23653 (N_23653,N_23346,N_22910);
or U23654 (N_23654,N_23294,N_23100);
or U23655 (N_23655,N_23078,N_23281);
xnor U23656 (N_23656,N_23014,N_23095);
xor U23657 (N_23657,N_23152,N_23122);
or U23658 (N_23658,N_22849,N_23036);
or U23659 (N_23659,N_23120,N_22961);
or U23660 (N_23660,N_22936,N_23242);
xor U23661 (N_23661,N_23098,N_23184);
nor U23662 (N_23662,N_23178,N_23068);
nand U23663 (N_23663,N_23273,N_22981);
or U23664 (N_23664,N_23085,N_23298);
or U23665 (N_23665,N_22939,N_23318);
or U23666 (N_23666,N_23205,N_23108);
nor U23667 (N_23667,N_22959,N_23392);
and U23668 (N_23668,N_23228,N_23125);
nand U23669 (N_23669,N_23376,N_22993);
nand U23670 (N_23670,N_22971,N_23056);
nor U23671 (N_23671,N_23225,N_23024);
or U23672 (N_23672,N_22891,N_23312);
xnor U23673 (N_23673,N_23047,N_23075);
xor U23674 (N_23674,N_23197,N_23348);
or U23675 (N_23675,N_22911,N_23090);
nand U23676 (N_23676,N_23094,N_22904);
and U23677 (N_23677,N_23092,N_23053);
or U23678 (N_23678,N_23156,N_23031);
xor U23679 (N_23679,N_23363,N_22823);
or U23680 (N_23680,N_22850,N_22851);
and U23681 (N_23681,N_23189,N_23240);
xnor U23682 (N_23682,N_22888,N_22932);
or U23683 (N_23683,N_23278,N_23046);
nand U23684 (N_23684,N_23138,N_23379);
or U23685 (N_23685,N_23362,N_22909);
and U23686 (N_23686,N_23015,N_23326);
or U23687 (N_23687,N_22882,N_22922);
nor U23688 (N_23688,N_23227,N_22920);
nand U23689 (N_23689,N_23267,N_23155);
nor U23690 (N_23690,N_22962,N_22965);
nand U23691 (N_23691,N_22834,N_23117);
nor U23692 (N_23692,N_22917,N_23373);
xor U23693 (N_23693,N_23061,N_22878);
xor U23694 (N_23694,N_23370,N_23030);
or U23695 (N_23695,N_23044,N_23258);
nor U23696 (N_23696,N_22988,N_23272);
xnor U23697 (N_23697,N_23062,N_23106);
xor U23698 (N_23698,N_23299,N_23304);
xor U23699 (N_23699,N_23020,N_23223);
nand U23700 (N_23700,N_23284,N_23150);
and U23701 (N_23701,N_23117,N_22940);
or U23702 (N_23702,N_22874,N_22808);
xnor U23703 (N_23703,N_23003,N_23170);
and U23704 (N_23704,N_22905,N_23395);
xor U23705 (N_23705,N_23013,N_23104);
or U23706 (N_23706,N_22876,N_23114);
nor U23707 (N_23707,N_22863,N_23351);
nor U23708 (N_23708,N_23287,N_23148);
nand U23709 (N_23709,N_23095,N_22913);
xnor U23710 (N_23710,N_23330,N_23058);
nand U23711 (N_23711,N_22859,N_23284);
or U23712 (N_23712,N_23218,N_23196);
and U23713 (N_23713,N_23280,N_22926);
xor U23714 (N_23714,N_23113,N_23130);
xnor U23715 (N_23715,N_22861,N_23383);
nor U23716 (N_23716,N_22879,N_23035);
and U23717 (N_23717,N_22827,N_22935);
and U23718 (N_23718,N_22952,N_23150);
nand U23719 (N_23719,N_23149,N_22947);
xor U23720 (N_23720,N_23258,N_23164);
or U23721 (N_23721,N_22910,N_23162);
and U23722 (N_23722,N_23052,N_23091);
xor U23723 (N_23723,N_23141,N_22872);
xor U23724 (N_23724,N_23396,N_23140);
xnor U23725 (N_23725,N_22945,N_22915);
and U23726 (N_23726,N_23187,N_23159);
xnor U23727 (N_23727,N_23266,N_22844);
nand U23728 (N_23728,N_22984,N_22944);
nand U23729 (N_23729,N_22922,N_22866);
or U23730 (N_23730,N_22959,N_22814);
or U23731 (N_23731,N_23088,N_23353);
or U23732 (N_23732,N_22926,N_23167);
xnor U23733 (N_23733,N_23193,N_23391);
and U23734 (N_23734,N_23345,N_23042);
nand U23735 (N_23735,N_23273,N_23211);
xor U23736 (N_23736,N_23202,N_23179);
or U23737 (N_23737,N_22899,N_22897);
xnor U23738 (N_23738,N_22948,N_22949);
xnor U23739 (N_23739,N_22889,N_22906);
or U23740 (N_23740,N_22929,N_23331);
xor U23741 (N_23741,N_23298,N_23374);
or U23742 (N_23742,N_23180,N_23396);
nor U23743 (N_23743,N_23266,N_23091);
or U23744 (N_23744,N_22834,N_23066);
or U23745 (N_23745,N_22802,N_23094);
or U23746 (N_23746,N_22984,N_23379);
or U23747 (N_23747,N_23151,N_23175);
nand U23748 (N_23748,N_23021,N_23298);
or U23749 (N_23749,N_23120,N_22905);
xnor U23750 (N_23750,N_23012,N_22873);
xnor U23751 (N_23751,N_23052,N_23135);
nor U23752 (N_23752,N_22908,N_23373);
or U23753 (N_23753,N_22854,N_22963);
or U23754 (N_23754,N_23309,N_22813);
xnor U23755 (N_23755,N_22865,N_23377);
nand U23756 (N_23756,N_22981,N_23006);
nand U23757 (N_23757,N_23101,N_22930);
nor U23758 (N_23758,N_23196,N_22824);
nor U23759 (N_23759,N_23317,N_23269);
and U23760 (N_23760,N_23223,N_23025);
and U23761 (N_23761,N_23290,N_23291);
nor U23762 (N_23762,N_23141,N_23319);
and U23763 (N_23763,N_22955,N_23013);
nor U23764 (N_23764,N_23174,N_23176);
and U23765 (N_23765,N_22896,N_23274);
or U23766 (N_23766,N_22976,N_22905);
xnor U23767 (N_23767,N_22802,N_23079);
and U23768 (N_23768,N_23148,N_22832);
or U23769 (N_23769,N_23243,N_23277);
or U23770 (N_23770,N_23226,N_23159);
or U23771 (N_23771,N_22989,N_23177);
and U23772 (N_23772,N_23191,N_22850);
and U23773 (N_23773,N_23138,N_23082);
nand U23774 (N_23774,N_23009,N_23140);
or U23775 (N_23775,N_23003,N_23037);
xnor U23776 (N_23776,N_22803,N_23341);
nor U23777 (N_23777,N_22802,N_23362);
nor U23778 (N_23778,N_23238,N_23298);
nor U23779 (N_23779,N_22868,N_22840);
or U23780 (N_23780,N_23221,N_22808);
or U23781 (N_23781,N_23059,N_23158);
xnor U23782 (N_23782,N_22827,N_22841);
and U23783 (N_23783,N_22954,N_22869);
xnor U23784 (N_23784,N_23314,N_23080);
xnor U23785 (N_23785,N_23359,N_22852);
xnor U23786 (N_23786,N_23123,N_22999);
xnor U23787 (N_23787,N_22806,N_22897);
nor U23788 (N_23788,N_23215,N_23348);
nand U23789 (N_23789,N_23234,N_23241);
nor U23790 (N_23790,N_23092,N_23363);
nand U23791 (N_23791,N_23234,N_23108);
xnor U23792 (N_23792,N_23087,N_22827);
nor U23793 (N_23793,N_22970,N_23150);
nor U23794 (N_23794,N_23249,N_23033);
xnor U23795 (N_23795,N_22813,N_23198);
or U23796 (N_23796,N_23078,N_23030);
and U23797 (N_23797,N_22844,N_23113);
xor U23798 (N_23798,N_23311,N_23397);
xor U23799 (N_23799,N_23009,N_23339);
nor U23800 (N_23800,N_23279,N_23278);
xnor U23801 (N_23801,N_22886,N_22948);
xnor U23802 (N_23802,N_22993,N_22950);
nor U23803 (N_23803,N_22996,N_22917);
or U23804 (N_23804,N_23349,N_22824);
nor U23805 (N_23805,N_22949,N_23257);
or U23806 (N_23806,N_23302,N_22820);
nor U23807 (N_23807,N_23037,N_22940);
nand U23808 (N_23808,N_23257,N_23252);
or U23809 (N_23809,N_23222,N_22824);
nor U23810 (N_23810,N_22889,N_22922);
nor U23811 (N_23811,N_23002,N_23104);
nand U23812 (N_23812,N_22883,N_23199);
nand U23813 (N_23813,N_22879,N_22852);
nor U23814 (N_23814,N_23055,N_23247);
nor U23815 (N_23815,N_23333,N_23059);
nor U23816 (N_23816,N_23110,N_23229);
nand U23817 (N_23817,N_23396,N_23385);
nand U23818 (N_23818,N_22966,N_23336);
xor U23819 (N_23819,N_22956,N_22937);
or U23820 (N_23820,N_23126,N_22920);
xnor U23821 (N_23821,N_23015,N_23053);
nor U23822 (N_23822,N_23363,N_23182);
nor U23823 (N_23823,N_23354,N_23351);
nand U23824 (N_23824,N_23149,N_23202);
and U23825 (N_23825,N_23319,N_23237);
nand U23826 (N_23826,N_23343,N_23320);
and U23827 (N_23827,N_23018,N_23314);
and U23828 (N_23828,N_23364,N_23217);
and U23829 (N_23829,N_23070,N_23304);
or U23830 (N_23830,N_23171,N_22855);
and U23831 (N_23831,N_22926,N_23152);
nand U23832 (N_23832,N_23298,N_23317);
nand U23833 (N_23833,N_23047,N_23312);
xnor U23834 (N_23834,N_22989,N_23057);
nand U23835 (N_23835,N_23340,N_23112);
nor U23836 (N_23836,N_22851,N_23160);
xor U23837 (N_23837,N_22984,N_23041);
xor U23838 (N_23838,N_22933,N_22837);
nand U23839 (N_23839,N_22910,N_23047);
nand U23840 (N_23840,N_23000,N_23031);
nand U23841 (N_23841,N_22988,N_23225);
xor U23842 (N_23842,N_23097,N_23149);
xnor U23843 (N_23843,N_23230,N_23205);
nor U23844 (N_23844,N_22991,N_23070);
nor U23845 (N_23845,N_23073,N_23006);
nand U23846 (N_23846,N_23041,N_22914);
nor U23847 (N_23847,N_22912,N_22862);
xnor U23848 (N_23848,N_22834,N_22866);
nand U23849 (N_23849,N_22890,N_22812);
or U23850 (N_23850,N_23323,N_23085);
and U23851 (N_23851,N_22858,N_23139);
nor U23852 (N_23852,N_22997,N_23338);
nand U23853 (N_23853,N_23227,N_23394);
or U23854 (N_23854,N_23163,N_22910);
xor U23855 (N_23855,N_23185,N_22853);
nand U23856 (N_23856,N_23109,N_23165);
nand U23857 (N_23857,N_23181,N_23074);
and U23858 (N_23858,N_22911,N_23140);
xnor U23859 (N_23859,N_23071,N_23398);
nor U23860 (N_23860,N_23136,N_22839);
and U23861 (N_23861,N_22890,N_22979);
nor U23862 (N_23862,N_23080,N_22904);
nor U23863 (N_23863,N_23060,N_23372);
or U23864 (N_23864,N_22819,N_23213);
or U23865 (N_23865,N_22900,N_22837);
xnor U23866 (N_23866,N_22981,N_23053);
and U23867 (N_23867,N_23287,N_23064);
and U23868 (N_23868,N_22863,N_23125);
nand U23869 (N_23869,N_23362,N_23263);
or U23870 (N_23870,N_23379,N_23001);
or U23871 (N_23871,N_23124,N_23259);
xnor U23872 (N_23872,N_22898,N_23286);
nor U23873 (N_23873,N_23235,N_22890);
xor U23874 (N_23874,N_23095,N_23252);
nand U23875 (N_23875,N_22807,N_22989);
nand U23876 (N_23876,N_22855,N_23067);
and U23877 (N_23877,N_22816,N_22817);
nand U23878 (N_23878,N_22844,N_23273);
or U23879 (N_23879,N_23281,N_23306);
xnor U23880 (N_23880,N_23187,N_23034);
and U23881 (N_23881,N_23061,N_23049);
or U23882 (N_23882,N_23139,N_23320);
xnor U23883 (N_23883,N_22898,N_23071);
or U23884 (N_23884,N_22912,N_23216);
or U23885 (N_23885,N_22938,N_22873);
nor U23886 (N_23886,N_23209,N_23354);
xor U23887 (N_23887,N_23199,N_23148);
or U23888 (N_23888,N_23338,N_23388);
nor U23889 (N_23889,N_23134,N_23266);
xor U23890 (N_23890,N_22947,N_23226);
nor U23891 (N_23891,N_23347,N_23114);
nor U23892 (N_23892,N_23265,N_22865);
nor U23893 (N_23893,N_22816,N_23057);
xnor U23894 (N_23894,N_23134,N_23160);
and U23895 (N_23895,N_23074,N_23333);
nand U23896 (N_23896,N_23149,N_23255);
or U23897 (N_23897,N_22947,N_23300);
and U23898 (N_23898,N_22863,N_23176);
xnor U23899 (N_23899,N_23215,N_22814);
nor U23900 (N_23900,N_22997,N_23001);
nor U23901 (N_23901,N_23168,N_23319);
nor U23902 (N_23902,N_23268,N_23366);
or U23903 (N_23903,N_23357,N_23081);
and U23904 (N_23904,N_23197,N_23216);
and U23905 (N_23905,N_22977,N_22832);
or U23906 (N_23906,N_23072,N_23152);
nor U23907 (N_23907,N_22911,N_23121);
and U23908 (N_23908,N_22920,N_23328);
nor U23909 (N_23909,N_23226,N_23234);
xor U23910 (N_23910,N_23054,N_22949);
nor U23911 (N_23911,N_22997,N_23297);
xor U23912 (N_23912,N_22811,N_23159);
or U23913 (N_23913,N_22843,N_23034);
and U23914 (N_23914,N_23052,N_23191);
xor U23915 (N_23915,N_23359,N_23079);
and U23916 (N_23916,N_23291,N_23025);
or U23917 (N_23917,N_23127,N_22976);
and U23918 (N_23918,N_23146,N_23248);
or U23919 (N_23919,N_22824,N_23233);
nor U23920 (N_23920,N_23124,N_23019);
xnor U23921 (N_23921,N_23153,N_22831);
and U23922 (N_23922,N_22943,N_23195);
nor U23923 (N_23923,N_23129,N_23202);
or U23924 (N_23924,N_23347,N_23076);
nor U23925 (N_23925,N_23080,N_23275);
nand U23926 (N_23926,N_23320,N_23002);
xor U23927 (N_23927,N_23023,N_23043);
nand U23928 (N_23928,N_23366,N_22907);
and U23929 (N_23929,N_23019,N_23183);
nand U23930 (N_23930,N_23308,N_23131);
or U23931 (N_23931,N_23151,N_23319);
or U23932 (N_23932,N_23376,N_22937);
or U23933 (N_23933,N_23012,N_23282);
or U23934 (N_23934,N_23215,N_23052);
nor U23935 (N_23935,N_22988,N_23078);
or U23936 (N_23936,N_23243,N_23373);
xnor U23937 (N_23937,N_22846,N_22993);
nor U23938 (N_23938,N_23282,N_22939);
nor U23939 (N_23939,N_23384,N_23047);
and U23940 (N_23940,N_23294,N_23025);
nand U23941 (N_23941,N_23240,N_23177);
xnor U23942 (N_23942,N_22809,N_22834);
and U23943 (N_23943,N_23369,N_23333);
and U23944 (N_23944,N_23223,N_22946);
and U23945 (N_23945,N_22996,N_23008);
and U23946 (N_23946,N_23324,N_23138);
and U23947 (N_23947,N_22872,N_23104);
or U23948 (N_23948,N_22928,N_23184);
and U23949 (N_23949,N_23052,N_23356);
and U23950 (N_23950,N_23380,N_23137);
xnor U23951 (N_23951,N_22929,N_22990);
and U23952 (N_23952,N_22998,N_22917);
or U23953 (N_23953,N_23383,N_23309);
and U23954 (N_23954,N_22983,N_23336);
or U23955 (N_23955,N_23214,N_23306);
and U23956 (N_23956,N_23119,N_23321);
nand U23957 (N_23957,N_23206,N_23025);
xnor U23958 (N_23958,N_23280,N_23366);
and U23959 (N_23959,N_22944,N_23090);
and U23960 (N_23960,N_23218,N_23142);
xor U23961 (N_23961,N_23238,N_23025);
or U23962 (N_23962,N_22971,N_23271);
xnor U23963 (N_23963,N_23076,N_23215);
and U23964 (N_23964,N_23262,N_22868);
xnor U23965 (N_23965,N_23020,N_23361);
nor U23966 (N_23966,N_23137,N_23136);
and U23967 (N_23967,N_23324,N_23207);
nand U23968 (N_23968,N_22824,N_23039);
nand U23969 (N_23969,N_23050,N_23262);
nand U23970 (N_23970,N_22989,N_22914);
and U23971 (N_23971,N_22896,N_23363);
or U23972 (N_23972,N_23394,N_23358);
xnor U23973 (N_23973,N_22992,N_22833);
xor U23974 (N_23974,N_22974,N_22869);
or U23975 (N_23975,N_23070,N_23134);
or U23976 (N_23976,N_23132,N_23330);
and U23977 (N_23977,N_23108,N_23369);
or U23978 (N_23978,N_22882,N_23158);
and U23979 (N_23979,N_23377,N_23339);
nor U23980 (N_23980,N_23204,N_23013);
and U23981 (N_23981,N_22827,N_23229);
nor U23982 (N_23982,N_23310,N_23304);
and U23983 (N_23983,N_23142,N_23196);
and U23984 (N_23984,N_23353,N_22816);
nor U23985 (N_23985,N_23247,N_23063);
xnor U23986 (N_23986,N_23186,N_23139);
xnor U23987 (N_23987,N_22986,N_23090);
or U23988 (N_23988,N_23018,N_22803);
and U23989 (N_23989,N_22833,N_22919);
xor U23990 (N_23990,N_23384,N_23101);
xor U23991 (N_23991,N_23209,N_23109);
xnor U23992 (N_23992,N_23119,N_22923);
nand U23993 (N_23993,N_22891,N_22838);
xnor U23994 (N_23994,N_23393,N_23094);
and U23995 (N_23995,N_23017,N_23367);
and U23996 (N_23996,N_23003,N_22904);
and U23997 (N_23997,N_23247,N_23361);
xnor U23998 (N_23998,N_22958,N_22894);
nor U23999 (N_23999,N_22940,N_22920);
and U24000 (N_24000,N_23408,N_23744);
xnor U24001 (N_24001,N_23675,N_23583);
and U24002 (N_24002,N_23779,N_23891);
and U24003 (N_24003,N_23963,N_23411);
and U24004 (N_24004,N_23814,N_23867);
and U24005 (N_24005,N_23679,N_23949);
nand U24006 (N_24006,N_23993,N_23685);
xnor U24007 (N_24007,N_23809,N_23912);
nor U24008 (N_24008,N_23656,N_23995);
nand U24009 (N_24009,N_23506,N_23954);
nand U24010 (N_24010,N_23777,N_23775);
and U24011 (N_24011,N_23860,N_23498);
and U24012 (N_24012,N_23601,N_23973);
xor U24013 (N_24013,N_23765,N_23482);
and U24014 (N_24014,N_23519,N_23629);
xnor U24015 (N_24015,N_23405,N_23572);
nand U24016 (N_24016,N_23738,N_23933);
nand U24017 (N_24017,N_23714,N_23757);
nand U24018 (N_24018,N_23403,N_23707);
nor U24019 (N_24019,N_23609,N_23946);
nand U24020 (N_24020,N_23903,N_23795);
and U24021 (N_24021,N_23828,N_23546);
nand U24022 (N_24022,N_23691,N_23931);
and U24023 (N_24023,N_23771,N_23712);
nor U24024 (N_24024,N_23762,N_23663);
xor U24025 (N_24025,N_23450,N_23502);
nor U24026 (N_24026,N_23945,N_23430);
and U24027 (N_24027,N_23585,N_23441);
and U24028 (N_24028,N_23821,N_23892);
or U24029 (N_24029,N_23819,N_23513);
or U24030 (N_24030,N_23574,N_23471);
nor U24031 (N_24031,N_23454,N_23735);
nor U24032 (N_24032,N_23812,N_23829);
nor U24033 (N_24033,N_23889,N_23541);
xor U24034 (N_24034,N_23756,N_23568);
nor U24035 (N_24035,N_23758,N_23863);
and U24036 (N_24036,N_23528,N_23565);
nand U24037 (N_24037,N_23811,N_23416);
nand U24038 (N_24038,N_23780,N_23409);
or U24039 (N_24039,N_23831,N_23717);
or U24040 (N_24040,N_23970,N_23976);
or U24041 (N_24041,N_23670,N_23570);
nor U24042 (N_24042,N_23564,N_23861);
nor U24043 (N_24043,N_23996,N_23822);
nor U24044 (N_24044,N_23567,N_23603);
nor U24045 (N_24045,N_23415,N_23681);
or U24046 (N_24046,N_23900,N_23718);
nand U24047 (N_24047,N_23739,N_23635);
nor U24048 (N_24048,N_23888,N_23847);
nand U24049 (N_24049,N_23941,N_23952);
xor U24050 (N_24050,N_23404,N_23590);
nor U24051 (N_24051,N_23545,N_23916);
nor U24052 (N_24052,N_23790,N_23875);
or U24053 (N_24053,N_23763,N_23488);
or U24054 (N_24054,N_23470,N_23543);
and U24055 (N_24055,N_23742,N_23447);
and U24056 (N_24056,N_23436,N_23508);
nand U24057 (N_24057,N_23852,N_23817);
or U24058 (N_24058,N_23997,N_23424);
nand U24059 (N_24059,N_23885,N_23604);
xor U24060 (N_24060,N_23522,N_23840);
or U24061 (N_24061,N_23858,N_23682);
or U24062 (N_24062,N_23666,N_23526);
xnor U24063 (N_24063,N_23540,N_23461);
nor U24064 (N_24064,N_23710,N_23702);
or U24065 (N_24065,N_23808,N_23674);
xor U24066 (N_24066,N_23689,N_23703);
xor U24067 (N_24067,N_23524,N_23910);
and U24068 (N_24068,N_23451,N_23457);
and U24069 (N_24069,N_23878,N_23898);
or U24070 (N_24070,N_23928,N_23708);
xor U24071 (N_24071,N_23466,N_23641);
and U24072 (N_24072,N_23417,N_23669);
or U24073 (N_24073,N_23715,N_23854);
nor U24074 (N_24074,N_23975,N_23605);
or U24075 (N_24075,N_23726,N_23838);
xnor U24076 (N_24076,N_23772,N_23648);
and U24077 (N_24077,N_23535,N_23620);
and U24078 (N_24078,N_23581,N_23458);
nor U24079 (N_24079,N_23706,N_23614);
xnor U24080 (N_24080,N_23673,N_23848);
xor U24081 (N_24081,N_23723,N_23951);
or U24082 (N_24082,N_23406,N_23741);
and U24083 (N_24083,N_23445,N_23789);
nor U24084 (N_24084,N_23607,N_23944);
nor U24085 (N_24085,N_23783,N_23899);
nand U24086 (N_24086,N_23991,N_23504);
and U24087 (N_24087,N_23753,N_23971);
xor U24088 (N_24088,N_23988,N_23833);
xnor U24089 (N_24089,N_23495,N_23489);
and U24090 (N_24090,N_23523,N_23705);
nand U24091 (N_24091,N_23980,N_23839);
and U24092 (N_24092,N_23948,N_23732);
xnor U24093 (N_24093,N_23571,N_23761);
nor U24094 (N_24094,N_23425,N_23815);
or U24095 (N_24095,N_23734,N_23768);
or U24096 (N_24096,N_23781,N_23982);
nand U24097 (N_24097,N_23802,N_23719);
xnor U24098 (N_24098,N_23624,N_23446);
nand U24099 (N_24099,N_23449,N_23677);
or U24100 (N_24100,N_23643,N_23992);
nand U24101 (N_24101,N_23709,N_23942);
and U24102 (N_24102,N_23479,N_23544);
nor U24103 (N_24103,N_23902,N_23467);
or U24104 (N_24104,N_23953,N_23909);
or U24105 (N_24105,N_23501,N_23750);
nand U24106 (N_24106,N_23872,N_23754);
nor U24107 (N_24107,N_23429,N_23667);
xor U24108 (N_24108,N_23619,N_23859);
nor U24109 (N_24109,N_23977,N_23419);
nand U24110 (N_24110,N_23936,N_23748);
or U24111 (N_24111,N_23805,N_23455);
xnor U24112 (N_24112,N_23562,N_23960);
nor U24113 (N_24113,N_23751,N_23713);
nor U24114 (N_24114,N_23615,N_23925);
or U24115 (N_24115,N_23444,N_23786);
and U24116 (N_24116,N_23917,N_23743);
or U24117 (N_24117,N_23464,N_23651);
xor U24118 (N_24118,N_23695,N_23746);
and U24119 (N_24119,N_23979,N_23548);
xor U24120 (N_24120,N_23499,N_23456);
nand U24121 (N_24121,N_23935,N_23862);
or U24122 (N_24122,N_23955,N_23422);
nand U24123 (N_24123,N_23600,N_23553);
nor U24124 (N_24124,N_23532,N_23402);
nor U24125 (N_24125,N_23968,N_23428);
and U24126 (N_24126,N_23573,N_23906);
and U24127 (N_24127,N_23920,N_23640);
or U24128 (N_24128,N_23883,N_23652);
nand U24129 (N_24129,N_23791,N_23989);
or U24130 (N_24130,N_23593,N_23496);
xnor U24131 (N_24131,N_23832,N_23964);
xor U24132 (N_24132,N_23533,N_23400);
and U24133 (N_24133,N_23427,N_23694);
or U24134 (N_24134,N_23810,N_23664);
and U24135 (N_24135,N_23438,N_23655);
xnor U24136 (N_24136,N_23555,N_23820);
or U24137 (N_24137,N_23881,N_23686);
xor U24138 (N_24138,N_23797,N_23999);
nor U24139 (N_24139,N_23764,N_23550);
xor U24140 (N_24140,N_23922,N_23853);
nor U24141 (N_24141,N_23630,N_23850);
nor U24142 (N_24142,N_23632,N_23577);
nand U24143 (N_24143,N_23653,N_23967);
nand U24144 (N_24144,N_23517,N_23788);
or U24145 (N_24145,N_23990,N_23806);
nor U24146 (N_24146,N_23589,N_23401);
nor U24147 (N_24147,N_23827,N_23475);
nand U24148 (N_24148,N_23729,N_23646);
nor U24149 (N_24149,N_23986,N_23816);
xnor U24150 (N_24150,N_23678,N_23722);
and U24151 (N_24151,N_23700,N_23760);
xnor U24152 (N_24152,N_23837,N_23659);
xor U24153 (N_24153,N_23974,N_23904);
nor U24154 (N_24154,N_23873,N_23684);
xnor U24155 (N_24155,N_23895,N_23687);
nor U24156 (N_24156,N_23494,N_23650);
nor U24157 (N_24157,N_23759,N_23901);
nor U24158 (N_24158,N_23972,N_23957);
nand U24159 (N_24159,N_23824,N_23534);
nor U24160 (N_24160,N_23937,N_23721);
and U24161 (N_24161,N_23616,N_23849);
nand U24162 (N_24162,N_23793,N_23884);
nor U24163 (N_24163,N_23493,N_23418);
nor U24164 (N_24164,N_23561,N_23658);
and U24165 (N_24165,N_23897,N_23531);
xnor U24166 (N_24166,N_23490,N_23410);
nand U24167 (N_24167,N_23591,N_23530);
and U24168 (N_24168,N_23592,N_23939);
nand U24169 (N_24169,N_23654,N_23563);
xor U24170 (N_24170,N_23556,N_23639);
nor U24171 (N_24171,N_23453,N_23907);
or U24172 (N_24172,N_23688,N_23420);
or U24173 (N_24173,N_23575,N_23552);
and U24174 (N_24174,N_23882,N_23716);
nor U24175 (N_24175,N_23637,N_23433);
nand U24176 (N_24176,N_23938,N_23825);
and U24177 (N_24177,N_23927,N_23520);
and U24178 (N_24178,N_23537,N_23423);
nor U24179 (N_24179,N_23978,N_23911);
xnor U24180 (N_24180,N_23452,N_23484);
or U24181 (N_24181,N_23497,N_23886);
nand U24182 (N_24182,N_23855,N_23800);
nor U24183 (N_24183,N_23638,N_23787);
nand U24184 (N_24184,N_23966,N_23736);
xor U24185 (N_24185,N_23576,N_23435);
and U24186 (N_24186,N_23440,N_23894);
nor U24187 (N_24187,N_23893,N_23767);
nand U24188 (N_24188,N_23584,N_23961);
nor U24189 (N_24189,N_23985,N_23740);
and U24190 (N_24190,N_23460,N_23492);
or U24191 (N_24191,N_23836,N_23472);
or U24192 (N_24192,N_23518,N_23459);
and U24193 (N_24193,N_23940,N_23514);
or U24194 (N_24194,N_23926,N_23958);
or U24195 (N_24195,N_23769,N_23965);
nor U24196 (N_24196,N_23803,N_23554);
xnor U24197 (N_24197,N_23529,N_23476);
nor U24198 (N_24198,N_23680,N_23704);
xor U24199 (N_24199,N_23625,N_23558);
or U24200 (N_24200,N_23984,N_23595);
and U24201 (N_24201,N_23865,N_23602);
and U24202 (N_24202,N_23644,N_23645);
and U24203 (N_24203,N_23676,N_23657);
nor U24204 (N_24204,N_23807,N_23510);
nor U24205 (N_24205,N_23627,N_23994);
and U24206 (N_24206,N_23693,N_23606);
nor U24207 (N_24207,N_23857,N_23823);
nand U24208 (N_24208,N_23835,N_23798);
nand U24209 (N_24209,N_23801,N_23724);
or U24210 (N_24210,N_23439,N_23621);
or U24211 (N_24211,N_23804,N_23662);
nand U24212 (N_24212,N_23921,N_23880);
nand U24213 (N_24213,N_23956,N_23412);
or U24214 (N_24214,N_23516,N_23943);
and U24215 (N_24215,N_23536,N_23597);
xnor U24216 (N_24216,N_23887,N_23870);
nor U24217 (N_24217,N_23580,N_23711);
nor U24218 (N_24218,N_23642,N_23500);
nor U24219 (N_24219,N_23842,N_23813);
and U24220 (N_24220,N_23784,N_23628);
xnor U24221 (N_24221,N_23915,N_23549);
xor U24222 (N_24222,N_23720,N_23586);
nor U24223 (N_24223,N_23505,N_23923);
nor U24224 (N_24224,N_23622,N_23618);
nor U24225 (N_24225,N_23843,N_23962);
nand U24226 (N_24226,N_23818,N_23737);
and U24227 (N_24227,N_23442,N_23913);
or U24228 (N_24228,N_23871,N_23846);
and U24229 (N_24229,N_23566,N_23551);
xor U24230 (N_24230,N_23696,N_23733);
xnor U24231 (N_24231,N_23698,N_23557);
or U24232 (N_24232,N_23559,N_23692);
nand U24233 (N_24233,N_23727,N_23969);
and U24234 (N_24234,N_23672,N_23611);
or U24235 (N_24235,N_23539,N_23437);
xnor U24236 (N_24236,N_23649,N_23668);
nand U24237 (N_24237,N_23728,N_23699);
xnor U24238 (N_24238,N_23876,N_23799);
or U24239 (N_24239,N_23547,N_23623);
and U24240 (N_24240,N_23463,N_23918);
nand U24241 (N_24241,N_23599,N_23491);
nor U24242 (N_24242,N_23527,N_23485);
and U24243 (N_24243,N_23697,N_23512);
nor U24244 (N_24244,N_23594,N_23959);
nand U24245 (N_24245,N_23773,N_23874);
or U24246 (N_24246,N_23414,N_23851);
nor U24247 (N_24247,N_23785,N_23830);
xor U24248 (N_24248,N_23864,N_23478);
and U24249 (N_24249,N_23587,N_23929);
nand U24250 (N_24250,N_23998,N_23745);
or U24251 (N_24251,N_23770,N_23774);
xnor U24252 (N_24252,N_23776,N_23766);
nor U24253 (N_24253,N_23613,N_23596);
nand U24254 (N_24254,N_23486,N_23612);
or U24255 (N_24255,N_23462,N_23542);
nor U24256 (N_24256,N_23987,N_23503);
xor U24257 (N_24257,N_23469,N_23868);
nor U24258 (N_24258,N_23511,N_23731);
nor U24259 (N_24259,N_23582,N_23578);
xnor U24260 (N_24260,N_23473,N_23636);
and U24261 (N_24261,N_23661,N_23671);
xnor U24262 (N_24262,N_23730,N_23896);
or U24263 (N_24263,N_23480,N_23690);
nand U24264 (N_24264,N_23919,N_23487);
and U24265 (N_24265,N_23483,N_23569);
and U24266 (N_24266,N_23755,N_23579);
and U24267 (N_24267,N_23477,N_23908);
nor U24268 (N_24268,N_23468,N_23782);
or U24269 (N_24269,N_23905,N_23890);
nand U24270 (N_24270,N_23434,N_23507);
nor U24271 (N_24271,N_23826,N_23725);
or U24272 (N_24272,N_23794,N_23856);
xor U24273 (N_24273,N_23465,N_23869);
and U24274 (N_24274,N_23509,N_23749);
and U24275 (N_24275,N_23481,N_23413);
nor U24276 (N_24276,N_23841,N_23914);
xor U24277 (N_24277,N_23515,N_23443);
xor U24278 (N_24278,N_23633,N_23834);
or U24279 (N_24279,N_23796,N_23474);
nor U24280 (N_24280,N_23407,N_23924);
and U24281 (N_24281,N_23631,N_23950);
and U24282 (N_24282,N_23634,N_23747);
xor U24283 (N_24283,N_23521,N_23934);
nand U24284 (N_24284,N_23610,N_23426);
or U24285 (N_24285,N_23845,N_23448);
nor U24286 (N_24286,N_23932,N_23981);
and U24287 (N_24287,N_23626,N_23538);
nand U24288 (N_24288,N_23525,N_23431);
and U24289 (N_24289,N_23877,N_23844);
or U24290 (N_24290,N_23617,N_23947);
and U24291 (N_24291,N_23660,N_23752);
nand U24292 (N_24292,N_23866,N_23792);
xor U24293 (N_24293,N_23421,N_23608);
nand U24294 (N_24294,N_23647,N_23665);
or U24295 (N_24295,N_23879,N_23701);
and U24296 (N_24296,N_23930,N_23983);
nor U24297 (N_24297,N_23683,N_23598);
nand U24298 (N_24298,N_23432,N_23560);
xor U24299 (N_24299,N_23778,N_23588);
nor U24300 (N_24300,N_23402,N_23949);
xor U24301 (N_24301,N_23589,N_23615);
or U24302 (N_24302,N_23901,N_23652);
or U24303 (N_24303,N_23663,N_23773);
and U24304 (N_24304,N_23579,N_23603);
xor U24305 (N_24305,N_23404,N_23911);
nor U24306 (N_24306,N_23822,N_23675);
and U24307 (N_24307,N_23950,N_23654);
or U24308 (N_24308,N_23987,N_23578);
or U24309 (N_24309,N_23963,N_23936);
xor U24310 (N_24310,N_23435,N_23757);
nor U24311 (N_24311,N_23989,N_23501);
and U24312 (N_24312,N_23847,N_23940);
or U24313 (N_24313,N_23533,N_23817);
nor U24314 (N_24314,N_23878,N_23976);
or U24315 (N_24315,N_23935,N_23769);
xor U24316 (N_24316,N_23517,N_23745);
nor U24317 (N_24317,N_23504,N_23563);
and U24318 (N_24318,N_23684,N_23574);
nand U24319 (N_24319,N_23713,N_23421);
nor U24320 (N_24320,N_23918,N_23756);
or U24321 (N_24321,N_23963,N_23591);
or U24322 (N_24322,N_23902,N_23727);
nor U24323 (N_24323,N_23983,N_23799);
nand U24324 (N_24324,N_23994,N_23987);
or U24325 (N_24325,N_23838,N_23713);
nor U24326 (N_24326,N_23491,N_23506);
nand U24327 (N_24327,N_23420,N_23843);
nor U24328 (N_24328,N_23511,N_23445);
and U24329 (N_24329,N_23657,N_23848);
or U24330 (N_24330,N_23818,N_23734);
nand U24331 (N_24331,N_23797,N_23488);
and U24332 (N_24332,N_23863,N_23862);
or U24333 (N_24333,N_23580,N_23528);
nor U24334 (N_24334,N_23737,N_23847);
nand U24335 (N_24335,N_23542,N_23951);
or U24336 (N_24336,N_23456,N_23540);
and U24337 (N_24337,N_23702,N_23473);
nand U24338 (N_24338,N_23849,N_23900);
nor U24339 (N_24339,N_23979,N_23571);
nand U24340 (N_24340,N_23868,N_23522);
and U24341 (N_24341,N_23697,N_23490);
xor U24342 (N_24342,N_23732,N_23723);
nand U24343 (N_24343,N_23982,N_23921);
or U24344 (N_24344,N_23684,N_23605);
xor U24345 (N_24345,N_23789,N_23775);
nor U24346 (N_24346,N_23899,N_23721);
nand U24347 (N_24347,N_23545,N_23453);
nor U24348 (N_24348,N_23492,N_23552);
nor U24349 (N_24349,N_23927,N_23428);
or U24350 (N_24350,N_23655,N_23792);
xnor U24351 (N_24351,N_23606,N_23704);
and U24352 (N_24352,N_23556,N_23864);
or U24353 (N_24353,N_23857,N_23412);
nor U24354 (N_24354,N_23893,N_23588);
xor U24355 (N_24355,N_23565,N_23437);
or U24356 (N_24356,N_23908,N_23790);
xor U24357 (N_24357,N_23811,N_23700);
and U24358 (N_24358,N_23619,N_23551);
nand U24359 (N_24359,N_23597,N_23467);
nand U24360 (N_24360,N_23952,N_23980);
xor U24361 (N_24361,N_23533,N_23901);
xnor U24362 (N_24362,N_23904,N_23921);
nand U24363 (N_24363,N_23941,N_23436);
nor U24364 (N_24364,N_23533,N_23611);
nor U24365 (N_24365,N_23673,N_23970);
and U24366 (N_24366,N_23978,N_23719);
or U24367 (N_24367,N_23797,N_23430);
and U24368 (N_24368,N_23750,N_23700);
nand U24369 (N_24369,N_23456,N_23998);
nor U24370 (N_24370,N_23947,N_23998);
nor U24371 (N_24371,N_23859,N_23498);
and U24372 (N_24372,N_23703,N_23593);
nor U24373 (N_24373,N_23927,N_23967);
and U24374 (N_24374,N_23697,N_23795);
nand U24375 (N_24375,N_23774,N_23597);
nor U24376 (N_24376,N_23896,N_23506);
or U24377 (N_24377,N_23646,N_23829);
and U24378 (N_24378,N_23733,N_23407);
nand U24379 (N_24379,N_23474,N_23544);
nor U24380 (N_24380,N_23462,N_23913);
or U24381 (N_24381,N_23688,N_23721);
and U24382 (N_24382,N_23625,N_23431);
xor U24383 (N_24383,N_23718,N_23638);
and U24384 (N_24384,N_23709,N_23636);
nor U24385 (N_24385,N_23443,N_23847);
xor U24386 (N_24386,N_23606,N_23949);
xnor U24387 (N_24387,N_23823,N_23622);
and U24388 (N_24388,N_23874,N_23682);
xor U24389 (N_24389,N_23731,N_23720);
and U24390 (N_24390,N_23997,N_23903);
nand U24391 (N_24391,N_23615,N_23960);
or U24392 (N_24392,N_23712,N_23814);
nand U24393 (N_24393,N_23525,N_23608);
nor U24394 (N_24394,N_23986,N_23871);
and U24395 (N_24395,N_23585,N_23746);
nand U24396 (N_24396,N_23741,N_23994);
xor U24397 (N_24397,N_23756,N_23662);
or U24398 (N_24398,N_23806,N_23428);
xnor U24399 (N_24399,N_23510,N_23927);
nor U24400 (N_24400,N_23752,N_23725);
xor U24401 (N_24401,N_23643,N_23745);
nor U24402 (N_24402,N_23705,N_23673);
or U24403 (N_24403,N_23730,N_23940);
xnor U24404 (N_24404,N_23705,N_23447);
nand U24405 (N_24405,N_23677,N_23680);
nor U24406 (N_24406,N_23602,N_23767);
xor U24407 (N_24407,N_23530,N_23508);
or U24408 (N_24408,N_23775,N_23672);
or U24409 (N_24409,N_23426,N_23509);
and U24410 (N_24410,N_23413,N_23692);
xnor U24411 (N_24411,N_23492,N_23931);
nand U24412 (N_24412,N_23540,N_23620);
and U24413 (N_24413,N_23649,N_23569);
or U24414 (N_24414,N_23674,N_23521);
nor U24415 (N_24415,N_23951,N_23563);
xnor U24416 (N_24416,N_23633,N_23654);
nor U24417 (N_24417,N_23492,N_23495);
nor U24418 (N_24418,N_23627,N_23456);
nand U24419 (N_24419,N_23985,N_23960);
xor U24420 (N_24420,N_23614,N_23796);
nor U24421 (N_24421,N_23832,N_23944);
and U24422 (N_24422,N_23641,N_23922);
or U24423 (N_24423,N_23841,N_23559);
xor U24424 (N_24424,N_23520,N_23518);
nand U24425 (N_24425,N_23730,N_23491);
and U24426 (N_24426,N_23852,N_23962);
nor U24427 (N_24427,N_23632,N_23979);
xnor U24428 (N_24428,N_23563,N_23737);
xnor U24429 (N_24429,N_23584,N_23537);
or U24430 (N_24430,N_23842,N_23894);
nor U24431 (N_24431,N_23870,N_23909);
nor U24432 (N_24432,N_23993,N_23736);
or U24433 (N_24433,N_23678,N_23476);
or U24434 (N_24434,N_23547,N_23589);
nand U24435 (N_24435,N_23433,N_23408);
and U24436 (N_24436,N_23844,N_23791);
nand U24437 (N_24437,N_23466,N_23489);
xnor U24438 (N_24438,N_23531,N_23542);
nor U24439 (N_24439,N_23818,N_23751);
xnor U24440 (N_24440,N_23558,N_23591);
nand U24441 (N_24441,N_23444,N_23951);
xnor U24442 (N_24442,N_23845,N_23843);
xnor U24443 (N_24443,N_23418,N_23476);
nor U24444 (N_24444,N_23682,N_23593);
xnor U24445 (N_24445,N_23644,N_23610);
nand U24446 (N_24446,N_23574,N_23647);
xor U24447 (N_24447,N_23833,N_23648);
xor U24448 (N_24448,N_23742,N_23409);
nand U24449 (N_24449,N_23406,N_23976);
or U24450 (N_24450,N_23855,N_23870);
and U24451 (N_24451,N_23616,N_23700);
nor U24452 (N_24452,N_23646,N_23579);
nand U24453 (N_24453,N_23568,N_23592);
or U24454 (N_24454,N_23942,N_23731);
nor U24455 (N_24455,N_23805,N_23825);
nand U24456 (N_24456,N_23449,N_23609);
or U24457 (N_24457,N_23528,N_23573);
or U24458 (N_24458,N_23769,N_23736);
nand U24459 (N_24459,N_23977,N_23882);
xnor U24460 (N_24460,N_23432,N_23822);
and U24461 (N_24461,N_23804,N_23668);
and U24462 (N_24462,N_23736,N_23541);
nand U24463 (N_24463,N_23871,N_23483);
xnor U24464 (N_24464,N_23955,N_23819);
or U24465 (N_24465,N_23884,N_23734);
xnor U24466 (N_24466,N_23795,N_23819);
or U24467 (N_24467,N_23750,N_23483);
nand U24468 (N_24468,N_23825,N_23537);
or U24469 (N_24469,N_23474,N_23449);
nand U24470 (N_24470,N_23562,N_23687);
nand U24471 (N_24471,N_23801,N_23822);
and U24472 (N_24472,N_23696,N_23929);
or U24473 (N_24473,N_23772,N_23463);
xnor U24474 (N_24474,N_23594,N_23469);
nor U24475 (N_24475,N_23968,N_23706);
nor U24476 (N_24476,N_23410,N_23597);
or U24477 (N_24477,N_23433,N_23817);
or U24478 (N_24478,N_23466,N_23481);
nand U24479 (N_24479,N_23739,N_23768);
nor U24480 (N_24480,N_23680,N_23637);
or U24481 (N_24481,N_23477,N_23459);
nor U24482 (N_24482,N_23418,N_23425);
or U24483 (N_24483,N_23977,N_23755);
nand U24484 (N_24484,N_23975,N_23749);
and U24485 (N_24485,N_23877,N_23482);
nand U24486 (N_24486,N_23737,N_23529);
nand U24487 (N_24487,N_23617,N_23819);
or U24488 (N_24488,N_23520,N_23739);
nand U24489 (N_24489,N_23940,N_23484);
nor U24490 (N_24490,N_23708,N_23889);
nand U24491 (N_24491,N_23761,N_23995);
nor U24492 (N_24492,N_23832,N_23513);
xnor U24493 (N_24493,N_23993,N_23595);
and U24494 (N_24494,N_23795,N_23563);
xnor U24495 (N_24495,N_23793,N_23969);
and U24496 (N_24496,N_23873,N_23522);
xnor U24497 (N_24497,N_23639,N_23501);
xor U24498 (N_24498,N_23458,N_23727);
xnor U24499 (N_24499,N_23996,N_23849);
or U24500 (N_24500,N_23987,N_23753);
xor U24501 (N_24501,N_23974,N_23419);
nor U24502 (N_24502,N_23584,N_23895);
or U24503 (N_24503,N_23595,N_23990);
or U24504 (N_24504,N_23868,N_23900);
nand U24505 (N_24505,N_23859,N_23600);
nand U24506 (N_24506,N_23559,N_23954);
nand U24507 (N_24507,N_23646,N_23480);
and U24508 (N_24508,N_23805,N_23562);
and U24509 (N_24509,N_23712,N_23899);
nand U24510 (N_24510,N_23900,N_23565);
nand U24511 (N_24511,N_23490,N_23658);
and U24512 (N_24512,N_23639,N_23483);
xnor U24513 (N_24513,N_23517,N_23917);
xnor U24514 (N_24514,N_23621,N_23513);
xor U24515 (N_24515,N_23965,N_23633);
nor U24516 (N_24516,N_23400,N_23855);
xor U24517 (N_24517,N_23546,N_23799);
nor U24518 (N_24518,N_23836,N_23599);
nand U24519 (N_24519,N_23439,N_23551);
or U24520 (N_24520,N_23435,N_23763);
xnor U24521 (N_24521,N_23557,N_23760);
xor U24522 (N_24522,N_23498,N_23436);
nor U24523 (N_24523,N_23935,N_23623);
nand U24524 (N_24524,N_23873,N_23542);
nand U24525 (N_24525,N_23914,N_23884);
or U24526 (N_24526,N_23728,N_23533);
nor U24527 (N_24527,N_23534,N_23904);
nand U24528 (N_24528,N_23516,N_23956);
xor U24529 (N_24529,N_23802,N_23508);
and U24530 (N_24530,N_23776,N_23490);
and U24531 (N_24531,N_23762,N_23626);
nand U24532 (N_24532,N_23774,N_23809);
xor U24533 (N_24533,N_23987,N_23705);
xnor U24534 (N_24534,N_23647,N_23769);
xnor U24535 (N_24535,N_23790,N_23526);
or U24536 (N_24536,N_23671,N_23939);
and U24537 (N_24537,N_23750,N_23908);
nor U24538 (N_24538,N_23874,N_23426);
nor U24539 (N_24539,N_23646,N_23845);
and U24540 (N_24540,N_23915,N_23778);
xor U24541 (N_24541,N_23493,N_23805);
or U24542 (N_24542,N_23925,N_23733);
and U24543 (N_24543,N_23815,N_23755);
nor U24544 (N_24544,N_23674,N_23949);
xor U24545 (N_24545,N_23819,N_23646);
or U24546 (N_24546,N_23612,N_23813);
or U24547 (N_24547,N_23680,N_23621);
nand U24548 (N_24548,N_23851,N_23866);
nor U24549 (N_24549,N_23966,N_23994);
xnor U24550 (N_24550,N_23579,N_23963);
or U24551 (N_24551,N_23864,N_23535);
nor U24552 (N_24552,N_23493,N_23740);
nor U24553 (N_24553,N_23448,N_23695);
nand U24554 (N_24554,N_23402,N_23996);
and U24555 (N_24555,N_23891,N_23458);
xnor U24556 (N_24556,N_23560,N_23706);
or U24557 (N_24557,N_23676,N_23609);
or U24558 (N_24558,N_23864,N_23947);
and U24559 (N_24559,N_23997,N_23630);
nand U24560 (N_24560,N_23529,N_23777);
and U24561 (N_24561,N_23472,N_23676);
xor U24562 (N_24562,N_23880,N_23620);
nand U24563 (N_24563,N_23754,N_23644);
nor U24564 (N_24564,N_23880,N_23581);
or U24565 (N_24565,N_23728,N_23514);
nand U24566 (N_24566,N_23706,N_23504);
or U24567 (N_24567,N_23943,N_23913);
or U24568 (N_24568,N_23812,N_23482);
or U24569 (N_24569,N_23810,N_23841);
xnor U24570 (N_24570,N_23685,N_23737);
and U24571 (N_24571,N_23412,N_23456);
xnor U24572 (N_24572,N_23556,N_23696);
xor U24573 (N_24573,N_23852,N_23448);
xnor U24574 (N_24574,N_23533,N_23884);
or U24575 (N_24575,N_23630,N_23836);
xnor U24576 (N_24576,N_23964,N_23566);
nor U24577 (N_24577,N_23551,N_23658);
xnor U24578 (N_24578,N_23504,N_23553);
or U24579 (N_24579,N_23477,N_23751);
and U24580 (N_24580,N_23930,N_23514);
nor U24581 (N_24581,N_23541,N_23647);
nand U24582 (N_24582,N_23657,N_23699);
and U24583 (N_24583,N_23463,N_23936);
nand U24584 (N_24584,N_23564,N_23906);
and U24585 (N_24585,N_23873,N_23779);
xor U24586 (N_24586,N_23826,N_23767);
or U24587 (N_24587,N_23454,N_23845);
or U24588 (N_24588,N_23836,N_23898);
nor U24589 (N_24589,N_23639,N_23765);
nand U24590 (N_24590,N_23897,N_23818);
and U24591 (N_24591,N_23497,N_23528);
nand U24592 (N_24592,N_23993,N_23727);
xor U24593 (N_24593,N_23615,N_23553);
xnor U24594 (N_24594,N_23888,N_23640);
nand U24595 (N_24595,N_23717,N_23648);
nor U24596 (N_24596,N_23751,N_23813);
nor U24597 (N_24597,N_23425,N_23818);
nor U24598 (N_24598,N_23600,N_23619);
or U24599 (N_24599,N_23463,N_23792);
or U24600 (N_24600,N_24186,N_24154);
and U24601 (N_24601,N_24098,N_24380);
and U24602 (N_24602,N_24353,N_24320);
nand U24603 (N_24603,N_24296,N_24252);
or U24604 (N_24604,N_24257,N_24493);
and U24605 (N_24605,N_24286,N_24454);
or U24606 (N_24606,N_24197,N_24254);
xor U24607 (N_24607,N_24335,N_24152);
and U24608 (N_24608,N_24275,N_24025);
xnor U24609 (N_24609,N_24149,N_24094);
nor U24610 (N_24610,N_24321,N_24356);
nor U24611 (N_24611,N_24040,N_24531);
nor U24612 (N_24612,N_24176,N_24234);
and U24613 (N_24613,N_24375,N_24045);
and U24614 (N_24614,N_24279,N_24036);
nand U24615 (N_24615,N_24247,N_24245);
xnor U24616 (N_24616,N_24444,N_24563);
nand U24617 (N_24617,N_24537,N_24579);
or U24618 (N_24618,N_24136,N_24050);
or U24619 (N_24619,N_24478,N_24410);
xor U24620 (N_24620,N_24561,N_24293);
xnor U24621 (N_24621,N_24417,N_24528);
or U24622 (N_24622,N_24346,N_24474);
or U24623 (N_24623,N_24333,N_24250);
or U24624 (N_24624,N_24280,N_24158);
and U24625 (N_24625,N_24242,N_24143);
nor U24626 (N_24626,N_24379,N_24522);
and U24627 (N_24627,N_24300,N_24438);
nor U24628 (N_24628,N_24093,N_24437);
or U24629 (N_24629,N_24457,N_24559);
or U24630 (N_24630,N_24473,N_24418);
nand U24631 (N_24631,N_24381,N_24080);
nand U24632 (N_24632,N_24494,N_24170);
nor U24633 (N_24633,N_24448,N_24549);
or U24634 (N_24634,N_24368,N_24273);
nand U24635 (N_24635,N_24387,N_24396);
nor U24636 (N_24636,N_24187,N_24255);
or U24637 (N_24637,N_24433,N_24239);
nand U24638 (N_24638,N_24081,N_24403);
and U24639 (N_24639,N_24586,N_24486);
nor U24640 (N_24640,N_24503,N_24466);
or U24641 (N_24641,N_24012,N_24434);
nor U24642 (N_24642,N_24316,N_24551);
nand U24643 (N_24643,N_24035,N_24392);
nor U24644 (N_24644,N_24006,N_24569);
nand U24645 (N_24645,N_24395,N_24496);
or U24646 (N_24646,N_24340,N_24244);
xnor U24647 (N_24647,N_24538,N_24483);
or U24648 (N_24648,N_24424,N_24355);
and U24649 (N_24649,N_24156,N_24347);
nor U24650 (N_24650,N_24598,N_24352);
or U24651 (N_24651,N_24520,N_24270);
xnor U24652 (N_24652,N_24043,N_24521);
nand U24653 (N_24653,N_24595,N_24406);
nand U24654 (N_24654,N_24568,N_24363);
nor U24655 (N_24655,N_24066,N_24146);
and U24656 (N_24656,N_24120,N_24189);
xor U24657 (N_24657,N_24104,N_24177);
or U24658 (N_24658,N_24558,N_24384);
xor U24659 (N_24659,N_24402,N_24204);
and U24660 (N_24660,N_24307,N_24552);
or U24661 (N_24661,N_24211,N_24481);
xor U24662 (N_24662,N_24557,N_24354);
and U24663 (N_24663,N_24308,N_24578);
and U24664 (N_24664,N_24505,N_24231);
xor U24665 (N_24665,N_24000,N_24210);
nand U24666 (N_24666,N_24205,N_24342);
nor U24667 (N_24667,N_24084,N_24086);
or U24668 (N_24668,N_24126,N_24472);
xnor U24669 (N_24669,N_24562,N_24400);
and U24670 (N_24670,N_24208,N_24470);
nor U24671 (N_24671,N_24023,N_24370);
nand U24672 (N_24672,N_24243,N_24128);
and U24673 (N_24673,N_24408,N_24113);
nor U24674 (N_24674,N_24476,N_24180);
and U24675 (N_24675,N_24553,N_24580);
nand U24676 (N_24676,N_24348,N_24222);
xnor U24677 (N_24677,N_24100,N_24367);
and U24678 (N_24678,N_24570,N_24310);
nand U24679 (N_24679,N_24574,N_24449);
xnor U24680 (N_24680,N_24060,N_24376);
xor U24681 (N_24681,N_24504,N_24461);
or U24682 (N_24682,N_24053,N_24052);
or U24683 (N_24683,N_24423,N_24223);
or U24684 (N_24684,N_24193,N_24447);
xnor U24685 (N_24685,N_24394,N_24039);
and U24686 (N_24686,N_24338,N_24261);
nor U24687 (N_24687,N_24021,N_24185);
nand U24688 (N_24688,N_24018,N_24218);
and U24689 (N_24689,N_24059,N_24124);
or U24690 (N_24690,N_24389,N_24305);
xor U24691 (N_24691,N_24309,N_24322);
nor U24692 (N_24692,N_24369,N_24219);
and U24693 (N_24693,N_24482,N_24067);
nor U24694 (N_24694,N_24390,N_24539);
or U24695 (N_24695,N_24150,N_24217);
or U24696 (N_24696,N_24366,N_24372);
nor U24697 (N_24697,N_24287,N_24191);
xnor U24698 (N_24698,N_24589,N_24421);
nor U24699 (N_24699,N_24290,N_24031);
xor U24700 (N_24700,N_24456,N_24329);
nor U24701 (N_24701,N_24401,N_24141);
and U24702 (N_24702,N_24272,N_24238);
nand U24703 (N_24703,N_24215,N_24230);
nand U24704 (N_24704,N_24464,N_24164);
and U24705 (N_24705,N_24529,N_24121);
and U24706 (N_24706,N_24118,N_24485);
nand U24707 (N_24707,N_24014,N_24502);
and U24708 (N_24708,N_24029,N_24214);
and U24709 (N_24709,N_24301,N_24440);
nor U24710 (N_24710,N_24249,N_24324);
nand U24711 (N_24711,N_24548,N_24334);
nand U24712 (N_24712,N_24077,N_24543);
xor U24713 (N_24713,N_24587,N_24107);
nor U24714 (N_24714,N_24571,N_24047);
nor U24715 (N_24715,N_24148,N_24489);
xnor U24716 (N_24716,N_24479,N_24016);
nand U24717 (N_24717,N_24532,N_24005);
and U24718 (N_24718,N_24109,N_24122);
nand U24719 (N_24719,N_24393,N_24079);
and U24720 (N_24720,N_24398,N_24055);
xor U24721 (N_24721,N_24030,N_24248);
xor U24722 (N_24722,N_24588,N_24056);
nand U24723 (N_24723,N_24144,N_24477);
xnor U24724 (N_24724,N_24344,N_24350);
or U24725 (N_24725,N_24303,N_24337);
nand U24726 (N_24726,N_24452,N_24397);
or U24727 (N_24727,N_24560,N_24169);
nand U24728 (N_24728,N_24034,N_24510);
nor U24729 (N_24729,N_24003,N_24178);
nand U24730 (N_24730,N_24110,N_24265);
xnor U24731 (N_24731,N_24592,N_24419);
and U24732 (N_24732,N_24063,N_24179);
xnor U24733 (N_24733,N_24202,N_24357);
or U24734 (N_24734,N_24413,N_24446);
and U24735 (N_24735,N_24330,N_24546);
nor U24736 (N_24736,N_24581,N_24585);
nand U24737 (N_24737,N_24127,N_24371);
nor U24738 (N_24738,N_24256,N_24001);
or U24739 (N_24739,N_24475,N_24508);
and U24740 (N_24740,N_24313,N_24135);
nor U24741 (N_24741,N_24534,N_24276);
or U24742 (N_24742,N_24577,N_24274);
or U24743 (N_24743,N_24314,N_24200);
nor U24744 (N_24744,N_24129,N_24042);
nand U24745 (N_24745,N_24572,N_24069);
and U24746 (N_24746,N_24054,N_24108);
nor U24747 (N_24747,N_24591,N_24147);
and U24748 (N_24748,N_24099,N_24339);
nor U24749 (N_24749,N_24140,N_24299);
and U24750 (N_24750,N_24407,N_24530);
nor U24751 (N_24751,N_24385,N_24564);
or U24752 (N_24752,N_24192,N_24341);
nor U24753 (N_24753,N_24498,N_24360);
nor U24754 (N_24754,N_24058,N_24159);
and U24755 (N_24755,N_24114,N_24594);
and U24756 (N_24756,N_24554,N_24317);
and U24757 (N_24757,N_24227,N_24221);
or U24758 (N_24758,N_24511,N_24007);
and U24759 (N_24759,N_24377,N_24328);
xor U24760 (N_24760,N_24453,N_24203);
or U24761 (N_24761,N_24311,N_24288);
nand U24762 (N_24762,N_24028,N_24541);
and U24763 (N_24763,N_24240,N_24318);
and U24764 (N_24764,N_24495,N_24237);
or U24765 (N_24765,N_24388,N_24213);
or U24766 (N_24766,N_24291,N_24491);
or U24767 (N_24767,N_24289,N_24173);
and U24768 (N_24768,N_24471,N_24188);
or U24769 (N_24769,N_24343,N_24088);
xor U24770 (N_24770,N_24233,N_24183);
and U24771 (N_24771,N_24480,N_24365);
nor U24772 (N_24772,N_24116,N_24282);
nand U24773 (N_24773,N_24171,N_24246);
and U24774 (N_24774,N_24451,N_24409);
or U24775 (N_24775,N_24404,N_24106);
nor U24776 (N_24776,N_24445,N_24302);
nand U24777 (N_24777,N_24130,N_24263);
nor U24778 (N_24778,N_24096,N_24499);
xnor U24779 (N_24779,N_24165,N_24160);
and U24780 (N_24780,N_24362,N_24326);
xnor U24781 (N_24781,N_24573,N_24506);
xnor U24782 (N_24782,N_24414,N_24269);
nor U24783 (N_24783,N_24155,N_24184);
and U24784 (N_24784,N_24073,N_24582);
xnor U24785 (N_24785,N_24467,N_24181);
nor U24786 (N_24786,N_24102,N_24199);
or U24787 (N_24787,N_24226,N_24051);
nor U24788 (N_24788,N_24209,N_24294);
nand U24789 (N_24789,N_24224,N_24236);
nor U24790 (N_24790,N_24450,N_24142);
or U24791 (N_24791,N_24374,N_24095);
nand U24792 (N_24792,N_24415,N_24364);
and U24793 (N_24793,N_24206,N_24323);
xnor U24794 (N_24794,N_24429,N_24443);
xor U24795 (N_24795,N_24312,N_24439);
xor U24796 (N_24796,N_24391,N_24190);
nor U24797 (N_24797,N_24523,N_24004);
and U24798 (N_24798,N_24484,N_24138);
and U24799 (N_24799,N_24576,N_24207);
or U24800 (N_24800,N_24253,N_24426);
xnor U24801 (N_24801,N_24258,N_24596);
nor U24802 (N_24802,N_24022,N_24420);
nand U24803 (N_24803,N_24358,N_24009);
nor U24804 (N_24804,N_24458,N_24331);
and U24805 (N_24805,N_24068,N_24026);
and U24806 (N_24806,N_24351,N_24412);
xnor U24807 (N_24807,N_24441,N_24516);
nor U24808 (N_24808,N_24442,N_24597);
and U24809 (N_24809,N_24566,N_24168);
nor U24810 (N_24810,N_24545,N_24327);
or U24811 (N_24811,N_24512,N_24405);
and U24812 (N_24812,N_24262,N_24011);
or U24813 (N_24813,N_24500,N_24555);
nor U24814 (N_24814,N_24260,N_24195);
or U24815 (N_24815,N_24399,N_24278);
or U24816 (N_24816,N_24460,N_24044);
nand U24817 (N_24817,N_24097,N_24432);
nor U24818 (N_24818,N_24386,N_24599);
and U24819 (N_24819,N_24332,N_24198);
xnor U24820 (N_24820,N_24048,N_24137);
xnor U24821 (N_24821,N_24174,N_24065);
xor U24822 (N_24822,N_24550,N_24083);
xor U24823 (N_24823,N_24487,N_24085);
and U24824 (N_24824,N_24513,N_24153);
xnor U24825 (N_24825,N_24057,N_24216);
xnor U24826 (N_24826,N_24062,N_24325);
xor U24827 (N_24827,N_24527,N_24315);
nor U24828 (N_24828,N_24072,N_24519);
nor U24829 (N_24829,N_24336,N_24235);
xnor U24830 (N_24830,N_24172,N_24020);
nand U24831 (N_24831,N_24593,N_24431);
or U24832 (N_24832,N_24515,N_24071);
xnor U24833 (N_24833,N_24525,N_24359);
nor U24834 (N_24834,N_24092,N_24076);
nor U24835 (N_24835,N_24038,N_24468);
nand U24836 (N_24836,N_24281,N_24087);
and U24837 (N_24837,N_24161,N_24465);
or U24838 (N_24838,N_24268,N_24266);
or U24839 (N_24839,N_24567,N_24536);
and U24840 (N_24840,N_24017,N_24382);
or U24841 (N_24841,N_24070,N_24166);
xor U24842 (N_24842,N_24583,N_24427);
xor U24843 (N_24843,N_24112,N_24490);
or U24844 (N_24844,N_24383,N_24212);
and U24845 (N_24845,N_24533,N_24251);
nor U24846 (N_24846,N_24378,N_24037);
xnor U24847 (N_24847,N_24285,N_24132);
xnor U24848 (N_24848,N_24229,N_24319);
nand U24849 (N_24849,N_24074,N_24133);
xnor U24850 (N_24850,N_24232,N_24497);
or U24851 (N_24851,N_24027,N_24078);
xnor U24852 (N_24852,N_24526,N_24416);
and U24853 (N_24853,N_24123,N_24061);
xor U24854 (N_24854,N_24535,N_24139);
nand U24855 (N_24855,N_24013,N_24162);
nor U24856 (N_24856,N_24411,N_24225);
nor U24857 (N_24857,N_24151,N_24101);
nor U24858 (N_24858,N_24196,N_24544);
nand U24859 (N_24859,N_24241,N_24175);
or U24860 (N_24860,N_24157,N_24090);
nor U24861 (N_24861,N_24194,N_24119);
nor U24862 (N_24862,N_24264,N_24008);
nor U24863 (N_24863,N_24469,N_24145);
nor U24864 (N_24864,N_24117,N_24514);
or U24865 (N_24865,N_24297,N_24492);
xor U24866 (N_24866,N_24345,N_24488);
nand U24867 (N_24867,N_24306,N_24111);
and U24868 (N_24868,N_24304,N_24033);
nor U24869 (N_24869,N_24134,N_24015);
nand U24870 (N_24870,N_24032,N_24349);
xor U24871 (N_24871,N_24459,N_24428);
and U24872 (N_24872,N_24019,N_24540);
or U24873 (N_24873,N_24565,N_24298);
nor U24874 (N_24874,N_24590,N_24501);
and U24875 (N_24875,N_24046,N_24518);
xor U24876 (N_24876,N_24259,N_24267);
or U24877 (N_24877,N_24271,N_24435);
xor U24878 (N_24878,N_24002,N_24201);
and U24879 (N_24879,N_24064,N_24584);
and U24880 (N_24880,N_24507,N_24517);
xnor U24881 (N_24881,N_24115,N_24455);
xnor U24882 (N_24882,N_24373,N_24091);
or U24883 (N_24883,N_24167,N_24361);
and U24884 (N_24884,N_24125,N_24283);
nor U24885 (N_24885,N_24422,N_24509);
and U24886 (N_24886,N_24089,N_24105);
xnor U24887 (N_24887,N_24542,N_24292);
xnor U24888 (N_24888,N_24462,N_24041);
nor U24889 (N_24889,N_24436,N_24075);
nor U24890 (N_24890,N_24049,N_24103);
nand U24891 (N_24891,N_24220,N_24010);
and U24892 (N_24892,N_24024,N_24228);
and U24893 (N_24893,N_24430,N_24524);
xnor U24894 (N_24894,N_24284,N_24463);
nand U24895 (N_24895,N_24556,N_24182);
nand U24896 (N_24896,N_24082,N_24163);
nor U24897 (N_24897,N_24575,N_24425);
or U24898 (N_24898,N_24295,N_24547);
or U24899 (N_24899,N_24277,N_24131);
nand U24900 (N_24900,N_24550,N_24002);
or U24901 (N_24901,N_24319,N_24483);
and U24902 (N_24902,N_24245,N_24053);
xor U24903 (N_24903,N_24239,N_24392);
nor U24904 (N_24904,N_24451,N_24562);
and U24905 (N_24905,N_24511,N_24181);
nor U24906 (N_24906,N_24069,N_24124);
nand U24907 (N_24907,N_24470,N_24364);
nor U24908 (N_24908,N_24098,N_24007);
nor U24909 (N_24909,N_24532,N_24381);
xnor U24910 (N_24910,N_24004,N_24241);
or U24911 (N_24911,N_24035,N_24452);
nor U24912 (N_24912,N_24200,N_24417);
or U24913 (N_24913,N_24587,N_24070);
nor U24914 (N_24914,N_24230,N_24532);
xor U24915 (N_24915,N_24413,N_24115);
xnor U24916 (N_24916,N_24409,N_24584);
nand U24917 (N_24917,N_24216,N_24205);
xor U24918 (N_24918,N_24384,N_24397);
and U24919 (N_24919,N_24185,N_24251);
nor U24920 (N_24920,N_24227,N_24224);
xor U24921 (N_24921,N_24095,N_24525);
nand U24922 (N_24922,N_24039,N_24246);
and U24923 (N_24923,N_24056,N_24014);
or U24924 (N_24924,N_24120,N_24510);
nor U24925 (N_24925,N_24216,N_24593);
xor U24926 (N_24926,N_24113,N_24359);
or U24927 (N_24927,N_24094,N_24539);
or U24928 (N_24928,N_24055,N_24192);
or U24929 (N_24929,N_24547,N_24270);
nor U24930 (N_24930,N_24068,N_24599);
nand U24931 (N_24931,N_24334,N_24059);
or U24932 (N_24932,N_24252,N_24294);
nor U24933 (N_24933,N_24112,N_24450);
nand U24934 (N_24934,N_24468,N_24205);
or U24935 (N_24935,N_24536,N_24258);
or U24936 (N_24936,N_24123,N_24176);
nand U24937 (N_24937,N_24435,N_24185);
or U24938 (N_24938,N_24389,N_24452);
nor U24939 (N_24939,N_24195,N_24430);
and U24940 (N_24940,N_24156,N_24294);
nand U24941 (N_24941,N_24464,N_24308);
xnor U24942 (N_24942,N_24357,N_24147);
or U24943 (N_24943,N_24318,N_24180);
and U24944 (N_24944,N_24460,N_24351);
and U24945 (N_24945,N_24528,N_24317);
xor U24946 (N_24946,N_24207,N_24492);
nor U24947 (N_24947,N_24309,N_24325);
or U24948 (N_24948,N_24466,N_24215);
nor U24949 (N_24949,N_24346,N_24507);
nand U24950 (N_24950,N_24083,N_24535);
and U24951 (N_24951,N_24100,N_24434);
nand U24952 (N_24952,N_24385,N_24102);
nor U24953 (N_24953,N_24041,N_24544);
nand U24954 (N_24954,N_24162,N_24117);
xor U24955 (N_24955,N_24015,N_24586);
and U24956 (N_24956,N_24306,N_24399);
nor U24957 (N_24957,N_24155,N_24134);
nand U24958 (N_24958,N_24491,N_24563);
nor U24959 (N_24959,N_24568,N_24111);
nand U24960 (N_24960,N_24503,N_24463);
nor U24961 (N_24961,N_24020,N_24359);
and U24962 (N_24962,N_24158,N_24580);
and U24963 (N_24963,N_24399,N_24043);
xor U24964 (N_24964,N_24209,N_24481);
or U24965 (N_24965,N_24563,N_24588);
or U24966 (N_24966,N_24308,N_24013);
nand U24967 (N_24967,N_24268,N_24587);
xor U24968 (N_24968,N_24383,N_24381);
xor U24969 (N_24969,N_24392,N_24320);
or U24970 (N_24970,N_24554,N_24181);
nor U24971 (N_24971,N_24553,N_24242);
and U24972 (N_24972,N_24458,N_24325);
nand U24973 (N_24973,N_24510,N_24452);
nand U24974 (N_24974,N_24397,N_24369);
nand U24975 (N_24975,N_24417,N_24361);
nor U24976 (N_24976,N_24339,N_24588);
xnor U24977 (N_24977,N_24594,N_24167);
xor U24978 (N_24978,N_24297,N_24115);
and U24979 (N_24979,N_24350,N_24031);
nor U24980 (N_24980,N_24047,N_24453);
or U24981 (N_24981,N_24394,N_24525);
nand U24982 (N_24982,N_24404,N_24087);
nand U24983 (N_24983,N_24006,N_24098);
and U24984 (N_24984,N_24076,N_24575);
nand U24985 (N_24985,N_24375,N_24585);
xnor U24986 (N_24986,N_24444,N_24026);
nor U24987 (N_24987,N_24196,N_24432);
nor U24988 (N_24988,N_24142,N_24462);
nor U24989 (N_24989,N_24539,N_24215);
nand U24990 (N_24990,N_24180,N_24134);
nand U24991 (N_24991,N_24293,N_24143);
and U24992 (N_24992,N_24101,N_24086);
and U24993 (N_24993,N_24335,N_24547);
and U24994 (N_24994,N_24342,N_24139);
or U24995 (N_24995,N_24464,N_24112);
nor U24996 (N_24996,N_24151,N_24530);
or U24997 (N_24997,N_24449,N_24288);
and U24998 (N_24998,N_24295,N_24246);
nand U24999 (N_24999,N_24079,N_24398);
or U25000 (N_25000,N_24411,N_24455);
xor U25001 (N_25001,N_24530,N_24433);
xor U25002 (N_25002,N_24199,N_24569);
xor U25003 (N_25003,N_24221,N_24378);
or U25004 (N_25004,N_24421,N_24249);
xnor U25005 (N_25005,N_24398,N_24583);
nor U25006 (N_25006,N_24562,N_24514);
nand U25007 (N_25007,N_24195,N_24000);
or U25008 (N_25008,N_24423,N_24298);
nand U25009 (N_25009,N_24215,N_24447);
or U25010 (N_25010,N_24452,N_24048);
nor U25011 (N_25011,N_24350,N_24516);
nand U25012 (N_25012,N_24096,N_24570);
nor U25013 (N_25013,N_24071,N_24411);
and U25014 (N_25014,N_24000,N_24045);
nor U25015 (N_25015,N_24537,N_24347);
or U25016 (N_25016,N_24366,N_24415);
and U25017 (N_25017,N_24288,N_24043);
xnor U25018 (N_25018,N_24163,N_24296);
nor U25019 (N_25019,N_24261,N_24508);
nor U25020 (N_25020,N_24342,N_24107);
xnor U25021 (N_25021,N_24534,N_24175);
nor U25022 (N_25022,N_24402,N_24035);
nand U25023 (N_25023,N_24181,N_24558);
nand U25024 (N_25024,N_24102,N_24418);
nor U25025 (N_25025,N_24224,N_24379);
nand U25026 (N_25026,N_24230,N_24249);
xor U25027 (N_25027,N_24205,N_24287);
and U25028 (N_25028,N_24011,N_24325);
nand U25029 (N_25029,N_24213,N_24220);
nor U25030 (N_25030,N_24271,N_24485);
nor U25031 (N_25031,N_24214,N_24117);
and U25032 (N_25032,N_24187,N_24389);
or U25033 (N_25033,N_24595,N_24039);
and U25034 (N_25034,N_24466,N_24527);
or U25035 (N_25035,N_24205,N_24158);
nor U25036 (N_25036,N_24548,N_24012);
xnor U25037 (N_25037,N_24139,N_24522);
xnor U25038 (N_25038,N_24260,N_24554);
nand U25039 (N_25039,N_24574,N_24302);
and U25040 (N_25040,N_24049,N_24223);
or U25041 (N_25041,N_24495,N_24070);
and U25042 (N_25042,N_24036,N_24033);
nor U25043 (N_25043,N_24193,N_24355);
xnor U25044 (N_25044,N_24473,N_24470);
and U25045 (N_25045,N_24142,N_24018);
nand U25046 (N_25046,N_24101,N_24542);
xnor U25047 (N_25047,N_24520,N_24001);
xnor U25048 (N_25048,N_24489,N_24384);
xor U25049 (N_25049,N_24101,N_24529);
xor U25050 (N_25050,N_24331,N_24380);
nor U25051 (N_25051,N_24513,N_24505);
nand U25052 (N_25052,N_24497,N_24397);
or U25053 (N_25053,N_24593,N_24059);
nor U25054 (N_25054,N_24296,N_24468);
xnor U25055 (N_25055,N_24077,N_24132);
and U25056 (N_25056,N_24518,N_24184);
or U25057 (N_25057,N_24439,N_24010);
and U25058 (N_25058,N_24182,N_24126);
xnor U25059 (N_25059,N_24289,N_24047);
xnor U25060 (N_25060,N_24497,N_24387);
nor U25061 (N_25061,N_24324,N_24450);
nand U25062 (N_25062,N_24599,N_24590);
and U25063 (N_25063,N_24519,N_24051);
nor U25064 (N_25064,N_24067,N_24405);
and U25065 (N_25065,N_24183,N_24361);
xor U25066 (N_25066,N_24236,N_24330);
xnor U25067 (N_25067,N_24274,N_24060);
xnor U25068 (N_25068,N_24279,N_24269);
xnor U25069 (N_25069,N_24439,N_24296);
xor U25070 (N_25070,N_24285,N_24381);
nand U25071 (N_25071,N_24318,N_24201);
nand U25072 (N_25072,N_24062,N_24027);
and U25073 (N_25073,N_24435,N_24282);
xor U25074 (N_25074,N_24056,N_24012);
and U25075 (N_25075,N_24091,N_24200);
nor U25076 (N_25076,N_24323,N_24044);
and U25077 (N_25077,N_24330,N_24328);
and U25078 (N_25078,N_24588,N_24538);
or U25079 (N_25079,N_24464,N_24384);
and U25080 (N_25080,N_24544,N_24536);
and U25081 (N_25081,N_24379,N_24007);
nand U25082 (N_25082,N_24058,N_24276);
xor U25083 (N_25083,N_24419,N_24587);
xnor U25084 (N_25084,N_24575,N_24123);
nor U25085 (N_25085,N_24292,N_24370);
nor U25086 (N_25086,N_24476,N_24224);
nor U25087 (N_25087,N_24578,N_24368);
xnor U25088 (N_25088,N_24151,N_24238);
xor U25089 (N_25089,N_24294,N_24113);
nand U25090 (N_25090,N_24288,N_24335);
and U25091 (N_25091,N_24394,N_24148);
and U25092 (N_25092,N_24488,N_24565);
or U25093 (N_25093,N_24388,N_24009);
nor U25094 (N_25094,N_24149,N_24289);
or U25095 (N_25095,N_24110,N_24301);
nand U25096 (N_25096,N_24147,N_24570);
nor U25097 (N_25097,N_24049,N_24394);
or U25098 (N_25098,N_24514,N_24282);
nand U25099 (N_25099,N_24522,N_24036);
and U25100 (N_25100,N_24339,N_24137);
nor U25101 (N_25101,N_24119,N_24291);
and U25102 (N_25102,N_24297,N_24283);
nand U25103 (N_25103,N_24570,N_24465);
xnor U25104 (N_25104,N_24487,N_24538);
nor U25105 (N_25105,N_24336,N_24393);
nand U25106 (N_25106,N_24342,N_24029);
and U25107 (N_25107,N_24010,N_24230);
nand U25108 (N_25108,N_24417,N_24102);
nand U25109 (N_25109,N_24586,N_24559);
xor U25110 (N_25110,N_24198,N_24156);
xnor U25111 (N_25111,N_24399,N_24064);
xnor U25112 (N_25112,N_24374,N_24414);
nor U25113 (N_25113,N_24348,N_24130);
or U25114 (N_25114,N_24565,N_24301);
and U25115 (N_25115,N_24169,N_24223);
nor U25116 (N_25116,N_24200,N_24418);
or U25117 (N_25117,N_24564,N_24466);
nand U25118 (N_25118,N_24095,N_24092);
or U25119 (N_25119,N_24043,N_24542);
or U25120 (N_25120,N_24519,N_24531);
or U25121 (N_25121,N_24466,N_24591);
nor U25122 (N_25122,N_24113,N_24330);
or U25123 (N_25123,N_24182,N_24153);
or U25124 (N_25124,N_24201,N_24541);
nor U25125 (N_25125,N_24324,N_24063);
xnor U25126 (N_25126,N_24360,N_24410);
or U25127 (N_25127,N_24213,N_24319);
or U25128 (N_25128,N_24222,N_24089);
xnor U25129 (N_25129,N_24258,N_24288);
and U25130 (N_25130,N_24066,N_24556);
nor U25131 (N_25131,N_24203,N_24298);
nor U25132 (N_25132,N_24394,N_24434);
and U25133 (N_25133,N_24060,N_24188);
nor U25134 (N_25134,N_24053,N_24100);
nor U25135 (N_25135,N_24252,N_24390);
and U25136 (N_25136,N_24034,N_24511);
or U25137 (N_25137,N_24465,N_24403);
or U25138 (N_25138,N_24142,N_24442);
and U25139 (N_25139,N_24398,N_24047);
nor U25140 (N_25140,N_24507,N_24009);
and U25141 (N_25141,N_24433,N_24387);
xor U25142 (N_25142,N_24275,N_24579);
xnor U25143 (N_25143,N_24446,N_24390);
and U25144 (N_25144,N_24111,N_24389);
nand U25145 (N_25145,N_24057,N_24515);
or U25146 (N_25146,N_24595,N_24190);
nand U25147 (N_25147,N_24274,N_24396);
and U25148 (N_25148,N_24020,N_24478);
nor U25149 (N_25149,N_24475,N_24181);
and U25150 (N_25150,N_24099,N_24175);
xnor U25151 (N_25151,N_24591,N_24363);
nor U25152 (N_25152,N_24186,N_24590);
or U25153 (N_25153,N_24100,N_24563);
xor U25154 (N_25154,N_24068,N_24140);
or U25155 (N_25155,N_24028,N_24354);
or U25156 (N_25156,N_24222,N_24363);
xor U25157 (N_25157,N_24509,N_24094);
nor U25158 (N_25158,N_24308,N_24520);
and U25159 (N_25159,N_24549,N_24300);
nand U25160 (N_25160,N_24155,N_24497);
and U25161 (N_25161,N_24162,N_24110);
nor U25162 (N_25162,N_24414,N_24127);
xnor U25163 (N_25163,N_24456,N_24135);
nand U25164 (N_25164,N_24381,N_24074);
or U25165 (N_25165,N_24107,N_24044);
or U25166 (N_25166,N_24121,N_24118);
xnor U25167 (N_25167,N_24431,N_24383);
or U25168 (N_25168,N_24451,N_24478);
nor U25169 (N_25169,N_24509,N_24162);
nor U25170 (N_25170,N_24041,N_24403);
nor U25171 (N_25171,N_24349,N_24589);
and U25172 (N_25172,N_24232,N_24253);
nor U25173 (N_25173,N_24365,N_24228);
or U25174 (N_25174,N_24355,N_24142);
nand U25175 (N_25175,N_24577,N_24190);
xnor U25176 (N_25176,N_24214,N_24169);
and U25177 (N_25177,N_24422,N_24429);
or U25178 (N_25178,N_24087,N_24252);
xnor U25179 (N_25179,N_24396,N_24253);
or U25180 (N_25180,N_24327,N_24319);
nor U25181 (N_25181,N_24527,N_24035);
xor U25182 (N_25182,N_24166,N_24544);
nor U25183 (N_25183,N_24038,N_24549);
nor U25184 (N_25184,N_24133,N_24057);
xnor U25185 (N_25185,N_24512,N_24138);
and U25186 (N_25186,N_24352,N_24277);
and U25187 (N_25187,N_24300,N_24574);
nand U25188 (N_25188,N_24139,N_24037);
or U25189 (N_25189,N_24194,N_24251);
nand U25190 (N_25190,N_24107,N_24353);
nor U25191 (N_25191,N_24106,N_24530);
nor U25192 (N_25192,N_24587,N_24050);
nand U25193 (N_25193,N_24146,N_24175);
or U25194 (N_25194,N_24192,N_24178);
and U25195 (N_25195,N_24313,N_24443);
nand U25196 (N_25196,N_24072,N_24116);
and U25197 (N_25197,N_24415,N_24402);
and U25198 (N_25198,N_24329,N_24291);
nor U25199 (N_25199,N_24524,N_24194);
and U25200 (N_25200,N_24616,N_24816);
xor U25201 (N_25201,N_24728,N_24743);
xnor U25202 (N_25202,N_25095,N_25138);
nand U25203 (N_25203,N_24978,N_25183);
or U25204 (N_25204,N_24957,N_25034);
or U25205 (N_25205,N_24929,N_24736);
or U25206 (N_25206,N_25067,N_24760);
xnor U25207 (N_25207,N_24658,N_25037);
and U25208 (N_25208,N_24697,N_24864);
or U25209 (N_25209,N_24913,N_24730);
and U25210 (N_25210,N_24639,N_24802);
or U25211 (N_25211,N_25115,N_25197);
and U25212 (N_25212,N_25004,N_24909);
xnor U25213 (N_25213,N_24877,N_24608);
nand U25214 (N_25214,N_24763,N_25098);
or U25215 (N_25215,N_24750,N_25056);
and U25216 (N_25216,N_24718,N_25167);
xnor U25217 (N_25217,N_24725,N_24949);
and U25218 (N_25218,N_24969,N_24894);
nand U25219 (N_25219,N_25005,N_24838);
nor U25220 (N_25220,N_24719,N_25099);
and U25221 (N_25221,N_24903,N_24994);
xnor U25222 (N_25222,N_24635,N_24706);
xor U25223 (N_25223,N_24773,N_24920);
and U25224 (N_25224,N_24902,N_24840);
or U25225 (N_25225,N_24704,N_24765);
xor U25226 (N_25226,N_24601,N_25178);
nor U25227 (N_25227,N_24729,N_25134);
and U25228 (N_25228,N_25150,N_24636);
nor U25229 (N_25229,N_24711,N_25033);
nor U25230 (N_25230,N_24629,N_25137);
xor U25231 (N_25231,N_24649,N_25124);
xnor U25232 (N_25232,N_25113,N_24684);
nor U25233 (N_25233,N_24812,N_24866);
nor U25234 (N_25234,N_24678,N_24795);
nor U25235 (N_25235,N_24695,N_24680);
nor U25236 (N_25236,N_24785,N_25045);
nor U25237 (N_25237,N_25076,N_24828);
nand U25238 (N_25238,N_24609,N_25032);
or U25239 (N_25239,N_25157,N_25184);
xnor U25240 (N_25240,N_24674,N_25070);
nor U25241 (N_25241,N_24955,N_25130);
xnor U25242 (N_25242,N_24991,N_25109);
and U25243 (N_25243,N_24713,N_25008);
nor U25244 (N_25244,N_24921,N_25194);
or U25245 (N_25245,N_25125,N_25039);
nor U25246 (N_25246,N_25019,N_25191);
nand U25247 (N_25247,N_24858,N_25164);
and U25248 (N_25248,N_24982,N_24893);
xor U25249 (N_25249,N_24746,N_24822);
nand U25250 (N_25250,N_25022,N_24790);
nor U25251 (N_25251,N_24664,N_24880);
xnor U25252 (N_25252,N_24694,N_25000);
nand U25253 (N_25253,N_24979,N_25187);
nand U25254 (N_25254,N_24624,N_24737);
and U25255 (N_25255,N_24634,N_25020);
nand U25256 (N_25256,N_24830,N_24650);
nor U25257 (N_25257,N_24954,N_24977);
and U25258 (N_25258,N_24683,N_24853);
nor U25259 (N_25259,N_24871,N_24708);
or U25260 (N_25260,N_25176,N_25141);
xor U25261 (N_25261,N_24915,N_25041);
and U25262 (N_25262,N_25112,N_24881);
xor U25263 (N_25263,N_24848,N_24861);
nor U25264 (N_25264,N_25116,N_24603);
nor U25265 (N_25265,N_24745,N_25144);
nand U25266 (N_25266,N_25043,N_24803);
nand U25267 (N_25267,N_25096,N_24663);
nor U25268 (N_25268,N_25085,N_24827);
xnor U25269 (N_25269,N_25010,N_25162);
or U25270 (N_25270,N_24772,N_24922);
nor U25271 (N_25271,N_24723,N_24889);
nand U25272 (N_25272,N_24888,N_24999);
or U25273 (N_25273,N_24749,N_25123);
xor U25274 (N_25274,N_24669,N_25003);
or U25275 (N_25275,N_24897,N_24852);
nand U25276 (N_25276,N_24699,N_24679);
xor U25277 (N_25277,N_24644,N_24927);
nor U25278 (N_25278,N_25089,N_25110);
nor U25279 (N_25279,N_24914,N_24835);
or U25280 (N_25280,N_24910,N_24778);
nand U25281 (N_25281,N_24726,N_25073);
nand U25282 (N_25282,N_24739,N_24863);
or U25283 (N_25283,N_24899,N_25016);
or U25284 (N_25284,N_24740,N_24990);
and U25285 (N_25285,N_24618,N_24985);
nand U25286 (N_25286,N_25151,N_24892);
nand U25287 (N_25287,N_25092,N_24924);
nand U25288 (N_25288,N_24885,N_24604);
and U25289 (N_25289,N_24916,N_24700);
xor U25290 (N_25290,N_24950,N_24811);
nand U25291 (N_25291,N_25047,N_25105);
xor U25292 (N_25292,N_24770,N_25168);
nand U25293 (N_25293,N_25177,N_24904);
xnor U25294 (N_25294,N_24661,N_24926);
nor U25295 (N_25295,N_24630,N_24967);
and U25296 (N_25296,N_24813,N_24753);
nor U25297 (N_25297,N_25155,N_24829);
xor U25298 (N_25298,N_25195,N_24841);
and U25299 (N_25299,N_25148,N_24686);
nand U25300 (N_25300,N_24698,N_25060);
nor U25301 (N_25301,N_24947,N_24670);
or U25302 (N_25302,N_24952,N_24896);
and U25303 (N_25303,N_25158,N_24756);
nor U25304 (N_25304,N_24807,N_24797);
and U25305 (N_25305,N_24855,N_24878);
nor U25306 (N_25306,N_24677,N_24843);
or U25307 (N_25307,N_24972,N_24755);
or U25308 (N_25308,N_24958,N_24821);
or U25309 (N_25309,N_24685,N_25101);
nand U25310 (N_25310,N_25017,N_25011);
nand U25311 (N_25311,N_24944,N_24675);
or U25312 (N_25312,N_24987,N_24646);
and U25313 (N_25313,N_25147,N_24655);
or U25314 (N_25314,N_24776,N_24938);
nor U25315 (N_25315,N_25103,N_24891);
and U25316 (N_25316,N_24932,N_24814);
or U25317 (N_25317,N_24945,N_24784);
and U25318 (N_25318,N_25055,N_25044);
nand U25319 (N_25319,N_25031,N_25080);
xor U25320 (N_25320,N_25097,N_24605);
and U25321 (N_25321,N_25111,N_24879);
and U25322 (N_25322,N_24622,N_25030);
xor U25323 (N_25323,N_24724,N_25106);
nand U25324 (N_25324,N_24810,N_24825);
xnor U25325 (N_25325,N_24867,N_25093);
xor U25326 (N_25326,N_25153,N_24959);
and U25327 (N_25327,N_24942,N_24839);
and U25328 (N_25328,N_25025,N_25078);
nand U25329 (N_25329,N_24602,N_25023);
nand U25330 (N_25330,N_24925,N_24721);
or U25331 (N_25331,N_24870,N_24850);
or U25332 (N_25332,N_24672,N_25028);
or U25333 (N_25333,N_24611,N_25007);
xnor U25334 (N_25334,N_25169,N_24846);
and U25335 (N_25335,N_25050,N_24984);
and U25336 (N_25336,N_25174,N_24826);
nor U25337 (N_25337,N_24710,N_25122);
and U25338 (N_25338,N_24691,N_24742);
xor U25339 (N_25339,N_25058,N_24961);
or U25340 (N_25340,N_24845,N_25036);
or U25341 (N_25341,N_24633,N_24953);
xnor U25342 (N_25342,N_25118,N_24948);
xnor U25343 (N_25343,N_24720,N_24627);
xor U25344 (N_25344,N_24992,N_25090);
nand U25345 (N_25345,N_24615,N_24872);
nor U25346 (N_25346,N_24901,N_25139);
xor U25347 (N_25347,N_24906,N_24844);
or U25348 (N_25348,N_24671,N_24714);
or U25349 (N_25349,N_24715,N_24662);
and U25350 (N_25350,N_25152,N_24783);
nor U25351 (N_25351,N_24895,N_24780);
nand U25352 (N_25352,N_24762,N_24707);
nor U25353 (N_25353,N_25042,N_24918);
nor U25354 (N_25354,N_25057,N_24873);
nor U25355 (N_25355,N_25142,N_25027);
or U25356 (N_25356,N_24777,N_24693);
nand U25357 (N_25357,N_24923,N_25015);
nor U25358 (N_25358,N_24779,N_25040);
xor U25359 (N_25359,N_24817,N_25018);
nor U25360 (N_25360,N_24791,N_25029);
xor U25361 (N_25361,N_24875,N_25066);
and U25362 (N_25362,N_24641,N_24976);
nand U25363 (N_25363,N_24789,N_25171);
xor U25364 (N_25364,N_24761,N_24966);
xnor U25365 (N_25365,N_25062,N_24874);
nand U25366 (N_25366,N_24744,N_24939);
and U25367 (N_25367,N_24625,N_25046);
nor U25368 (N_25368,N_24722,N_24823);
nand U25369 (N_25369,N_24676,N_25006);
nand U25370 (N_25370,N_25013,N_25143);
and U25371 (N_25371,N_24653,N_25129);
or U25372 (N_25372,N_25038,N_24796);
nor U25373 (N_25373,N_24883,N_24717);
or U25374 (N_25374,N_24884,N_24887);
xnor U25375 (N_25375,N_25074,N_24775);
and U25376 (N_25376,N_24727,N_25069);
nand U25377 (N_25377,N_24696,N_24665);
xnor U25378 (N_25378,N_24933,N_24645);
nand U25379 (N_25379,N_24619,N_25064);
xnor U25380 (N_25380,N_24820,N_24824);
or U25381 (N_25381,N_24660,N_25082);
and U25382 (N_25382,N_24687,N_24692);
nand U25383 (N_25383,N_25052,N_25170);
nor U25384 (N_25384,N_24632,N_25145);
nor U25385 (N_25385,N_25001,N_24659);
xor U25386 (N_25386,N_24962,N_25135);
or U25387 (N_25387,N_25075,N_24862);
nor U25388 (N_25388,N_24754,N_24734);
xnor U25389 (N_25389,N_24876,N_24788);
nand U25390 (N_25390,N_24983,N_25181);
nand U25391 (N_25391,N_25012,N_25108);
xnor U25392 (N_25392,N_24620,N_24651);
xor U25393 (N_25393,N_24988,N_25014);
nand U25394 (N_25394,N_25172,N_25163);
xor U25395 (N_25395,N_25132,N_25068);
or U25396 (N_25396,N_24856,N_24946);
or U25397 (N_25397,N_24751,N_25182);
and U25398 (N_25398,N_24607,N_24794);
nand U25399 (N_25399,N_24836,N_25081);
xor U25400 (N_25400,N_24690,N_24793);
or U25401 (N_25401,N_24654,N_24865);
nand U25402 (N_25402,N_25024,N_24703);
xor U25403 (N_25403,N_25149,N_24617);
and U25404 (N_25404,N_24936,N_24640);
and U25405 (N_25405,N_25035,N_24767);
xor U25406 (N_25406,N_24831,N_24648);
or U25407 (N_25407,N_24613,N_25053);
xor U25408 (N_25408,N_24682,N_24732);
or U25409 (N_25409,N_24980,N_24857);
nand U25410 (N_25410,N_24781,N_24689);
xor U25411 (N_25411,N_24995,N_24766);
and U25412 (N_25412,N_24782,N_24759);
nor U25413 (N_25413,N_24786,N_25084);
xnor U25414 (N_25414,N_24774,N_24940);
nor U25415 (N_25415,N_24800,N_25117);
nor U25416 (N_25416,N_24974,N_24673);
and U25417 (N_25417,N_24842,N_24935);
nor U25418 (N_25418,N_24809,N_25065);
xnor U25419 (N_25419,N_25059,N_24834);
or U25420 (N_25420,N_24804,N_24768);
nor U25421 (N_25421,N_25083,N_24801);
and U25422 (N_25422,N_24981,N_24642);
xnor U25423 (N_25423,N_24657,N_24621);
nor U25424 (N_25424,N_25127,N_24747);
nor U25425 (N_25425,N_25100,N_24965);
or U25426 (N_25426,N_24963,N_24928);
or U25427 (N_25427,N_24837,N_24993);
and U25428 (N_25428,N_25166,N_25193);
nand U25429 (N_25429,N_24638,N_24712);
or U25430 (N_25430,N_25088,N_25049);
nor U25431 (N_25431,N_24631,N_24764);
or U25432 (N_25432,N_25175,N_24818);
or U25433 (N_25433,N_24805,N_24702);
or U25434 (N_25434,N_24833,N_24849);
nand U25435 (N_25435,N_24911,N_25173);
nand U25436 (N_25436,N_25156,N_24986);
and U25437 (N_25437,N_24968,N_24733);
or U25438 (N_25438,N_24907,N_24931);
or U25439 (N_25439,N_25009,N_25189);
nand U25440 (N_25440,N_24905,N_25063);
or U25441 (N_25441,N_25192,N_25119);
or U25442 (N_25442,N_24943,N_24930);
nand U25443 (N_25443,N_24757,N_25087);
xnor U25444 (N_25444,N_25185,N_24643);
nor U25445 (N_25445,N_25021,N_24851);
or U25446 (N_25446,N_24900,N_24647);
or U25447 (N_25447,N_24623,N_25159);
xor U25448 (N_25448,N_24792,N_24917);
and U25449 (N_25449,N_25114,N_24941);
and U25450 (N_25450,N_25199,N_25104);
nand U25451 (N_25451,N_25198,N_25165);
nand U25452 (N_25452,N_25131,N_24919);
and U25453 (N_25453,N_24758,N_24701);
xnor U25454 (N_25454,N_25077,N_24890);
xor U25455 (N_25455,N_24626,N_24668);
or U25456 (N_25456,N_24815,N_25140);
nand U25457 (N_25457,N_24799,N_24898);
nor U25458 (N_25458,N_24612,N_25188);
xor U25459 (N_25459,N_25136,N_24748);
nand U25460 (N_25460,N_24656,N_25121);
or U25461 (N_25461,N_24652,N_25160);
xor U25462 (N_25462,N_24996,N_25051);
or U25463 (N_25463,N_24868,N_25190);
and U25464 (N_25464,N_24964,N_25128);
xnor U25465 (N_25465,N_25094,N_24666);
nor U25466 (N_25466,N_25120,N_24735);
xor U25467 (N_25467,N_24752,N_25146);
nand U25468 (N_25468,N_24614,N_24882);
or U25469 (N_25469,N_24859,N_25133);
or U25470 (N_25470,N_24771,N_24860);
nand U25471 (N_25471,N_24934,N_24989);
xor U25472 (N_25472,N_24847,N_24681);
xor U25473 (N_25473,N_24806,N_24998);
xor U25474 (N_25474,N_24667,N_24628);
or U25475 (N_25475,N_24832,N_25002);
xnor U25476 (N_25476,N_24600,N_24738);
nand U25477 (N_25477,N_24606,N_24951);
nor U25478 (N_25478,N_24688,N_24610);
nand U25479 (N_25479,N_25086,N_24937);
or U25480 (N_25480,N_25054,N_24741);
and U25481 (N_25481,N_25126,N_24769);
and U25482 (N_25482,N_24975,N_24854);
and U25483 (N_25483,N_25180,N_25026);
or U25484 (N_25484,N_24798,N_25061);
xnor U25485 (N_25485,N_25154,N_25091);
or U25486 (N_25486,N_24705,N_24787);
nand U25487 (N_25487,N_25102,N_25107);
or U25488 (N_25488,N_24637,N_24956);
nor U25489 (N_25489,N_25072,N_25179);
or U25490 (N_25490,N_25071,N_24886);
and U25491 (N_25491,N_25196,N_24973);
nand U25492 (N_25492,N_24912,N_24716);
or U25493 (N_25493,N_24819,N_24997);
xnor U25494 (N_25494,N_25161,N_25079);
xnor U25495 (N_25495,N_24869,N_25186);
nand U25496 (N_25496,N_24731,N_24908);
nand U25497 (N_25497,N_24970,N_24971);
or U25498 (N_25498,N_25048,N_24709);
and U25499 (N_25499,N_24808,N_24960);
or U25500 (N_25500,N_25079,N_25089);
and U25501 (N_25501,N_24816,N_25142);
xnor U25502 (N_25502,N_25189,N_24781);
nor U25503 (N_25503,N_24966,N_25134);
and U25504 (N_25504,N_25047,N_24834);
and U25505 (N_25505,N_24619,N_24730);
nand U25506 (N_25506,N_24740,N_24728);
nand U25507 (N_25507,N_25011,N_25131);
and U25508 (N_25508,N_24670,N_24964);
and U25509 (N_25509,N_25111,N_25107);
and U25510 (N_25510,N_24777,N_24908);
or U25511 (N_25511,N_25074,N_25068);
xnor U25512 (N_25512,N_24795,N_24734);
and U25513 (N_25513,N_25147,N_24651);
or U25514 (N_25514,N_24906,N_25060);
nor U25515 (N_25515,N_24992,N_24736);
nand U25516 (N_25516,N_24924,N_25109);
or U25517 (N_25517,N_24928,N_25136);
xnor U25518 (N_25518,N_24649,N_25046);
xnor U25519 (N_25519,N_25181,N_24822);
nand U25520 (N_25520,N_24986,N_25142);
or U25521 (N_25521,N_25199,N_24908);
and U25522 (N_25522,N_25049,N_25135);
and U25523 (N_25523,N_24918,N_24885);
xnor U25524 (N_25524,N_24957,N_24633);
nor U25525 (N_25525,N_24998,N_24896);
nand U25526 (N_25526,N_24937,N_25122);
xor U25527 (N_25527,N_24755,N_24620);
nand U25528 (N_25528,N_24606,N_24749);
or U25529 (N_25529,N_24980,N_24760);
nand U25530 (N_25530,N_25197,N_25125);
nand U25531 (N_25531,N_25008,N_24896);
and U25532 (N_25532,N_24869,N_24685);
or U25533 (N_25533,N_24968,N_24818);
xnor U25534 (N_25534,N_25153,N_24730);
and U25535 (N_25535,N_25003,N_24812);
nand U25536 (N_25536,N_24757,N_24715);
xnor U25537 (N_25537,N_24692,N_24671);
or U25538 (N_25538,N_24891,N_24744);
and U25539 (N_25539,N_24686,N_24772);
and U25540 (N_25540,N_24947,N_24749);
nand U25541 (N_25541,N_24961,N_24811);
nand U25542 (N_25542,N_24767,N_24967);
and U25543 (N_25543,N_24614,N_24674);
nand U25544 (N_25544,N_25160,N_24903);
and U25545 (N_25545,N_24802,N_25173);
nor U25546 (N_25546,N_25173,N_24693);
and U25547 (N_25547,N_24673,N_25032);
xor U25548 (N_25548,N_25106,N_24888);
nor U25549 (N_25549,N_24843,N_25094);
nor U25550 (N_25550,N_25133,N_24733);
and U25551 (N_25551,N_24738,N_25173);
or U25552 (N_25552,N_24824,N_24836);
xnor U25553 (N_25553,N_25054,N_25140);
nand U25554 (N_25554,N_24750,N_24757);
nor U25555 (N_25555,N_24691,N_25072);
nor U25556 (N_25556,N_25077,N_24601);
or U25557 (N_25557,N_25030,N_24798);
or U25558 (N_25558,N_24846,N_24835);
nor U25559 (N_25559,N_24743,N_24834);
or U25560 (N_25560,N_24824,N_24988);
or U25561 (N_25561,N_24842,N_24771);
xor U25562 (N_25562,N_24737,N_24678);
and U25563 (N_25563,N_25071,N_25146);
and U25564 (N_25564,N_24815,N_24870);
or U25565 (N_25565,N_24928,N_24975);
xnor U25566 (N_25566,N_25166,N_24703);
and U25567 (N_25567,N_24964,N_24783);
xor U25568 (N_25568,N_24887,N_24881);
xor U25569 (N_25569,N_24692,N_25184);
xor U25570 (N_25570,N_25120,N_25058);
xor U25571 (N_25571,N_25020,N_24858);
xor U25572 (N_25572,N_25106,N_24985);
nor U25573 (N_25573,N_24695,N_24849);
and U25574 (N_25574,N_24601,N_24967);
nor U25575 (N_25575,N_25156,N_24891);
or U25576 (N_25576,N_24883,N_24996);
nor U25577 (N_25577,N_24871,N_24684);
and U25578 (N_25578,N_24740,N_25047);
xor U25579 (N_25579,N_25123,N_25006);
nand U25580 (N_25580,N_25180,N_24785);
or U25581 (N_25581,N_25169,N_25017);
nand U25582 (N_25582,N_24818,N_24837);
nor U25583 (N_25583,N_24819,N_25193);
or U25584 (N_25584,N_24694,N_24672);
or U25585 (N_25585,N_24962,N_24818);
xnor U25586 (N_25586,N_25009,N_24654);
and U25587 (N_25587,N_24745,N_25163);
and U25588 (N_25588,N_24769,N_24956);
nor U25589 (N_25589,N_24943,N_24840);
nand U25590 (N_25590,N_25065,N_24650);
nand U25591 (N_25591,N_25033,N_24674);
or U25592 (N_25592,N_24684,N_25199);
and U25593 (N_25593,N_24623,N_25035);
nand U25594 (N_25594,N_24929,N_24831);
and U25595 (N_25595,N_24813,N_25090);
xnor U25596 (N_25596,N_24811,N_24631);
nor U25597 (N_25597,N_25191,N_24850);
xor U25598 (N_25598,N_25141,N_25170);
xor U25599 (N_25599,N_24840,N_24643);
nand U25600 (N_25600,N_24608,N_25064);
nand U25601 (N_25601,N_25150,N_24743);
and U25602 (N_25602,N_25101,N_24674);
and U25603 (N_25603,N_24652,N_25067);
and U25604 (N_25604,N_25045,N_24910);
and U25605 (N_25605,N_25113,N_24856);
nor U25606 (N_25606,N_24988,N_24798);
or U25607 (N_25607,N_24676,N_24837);
nand U25608 (N_25608,N_24803,N_25118);
or U25609 (N_25609,N_24959,N_24634);
xnor U25610 (N_25610,N_25000,N_24880);
xor U25611 (N_25611,N_24847,N_24866);
or U25612 (N_25612,N_24610,N_24946);
and U25613 (N_25613,N_25134,N_24735);
and U25614 (N_25614,N_24784,N_24944);
or U25615 (N_25615,N_24870,N_25041);
nand U25616 (N_25616,N_24723,N_24997);
nor U25617 (N_25617,N_24827,N_24700);
and U25618 (N_25618,N_24655,N_24941);
nor U25619 (N_25619,N_25106,N_25092);
or U25620 (N_25620,N_24813,N_25052);
xor U25621 (N_25621,N_25099,N_25195);
or U25622 (N_25622,N_24832,N_24823);
and U25623 (N_25623,N_25099,N_24873);
or U25624 (N_25624,N_24988,N_24699);
or U25625 (N_25625,N_25107,N_25042);
and U25626 (N_25626,N_25011,N_25042);
or U25627 (N_25627,N_25057,N_24976);
xor U25628 (N_25628,N_25172,N_24861);
and U25629 (N_25629,N_24817,N_24772);
xor U25630 (N_25630,N_25000,N_24858);
nand U25631 (N_25631,N_24616,N_24683);
nand U25632 (N_25632,N_24649,N_25056);
xnor U25633 (N_25633,N_24677,N_25011);
or U25634 (N_25634,N_24783,N_25085);
nor U25635 (N_25635,N_24666,N_25052);
xor U25636 (N_25636,N_24607,N_24657);
nand U25637 (N_25637,N_24874,N_24953);
nor U25638 (N_25638,N_24961,N_24709);
xnor U25639 (N_25639,N_25039,N_25071);
and U25640 (N_25640,N_24934,N_24687);
and U25641 (N_25641,N_24924,N_25128);
nor U25642 (N_25642,N_24938,N_24636);
nand U25643 (N_25643,N_25184,N_25148);
or U25644 (N_25644,N_25061,N_24674);
xor U25645 (N_25645,N_24671,N_25130);
nor U25646 (N_25646,N_24824,N_25055);
xnor U25647 (N_25647,N_25129,N_25032);
xnor U25648 (N_25648,N_25191,N_24738);
xnor U25649 (N_25649,N_24804,N_24799);
or U25650 (N_25650,N_25072,N_24884);
or U25651 (N_25651,N_24629,N_24660);
nand U25652 (N_25652,N_24751,N_24631);
or U25653 (N_25653,N_25087,N_24641);
nor U25654 (N_25654,N_24649,N_25095);
and U25655 (N_25655,N_25080,N_25198);
nand U25656 (N_25656,N_25141,N_25188);
or U25657 (N_25657,N_24791,N_24890);
nor U25658 (N_25658,N_25026,N_24639);
and U25659 (N_25659,N_25014,N_24954);
nand U25660 (N_25660,N_24747,N_24936);
xnor U25661 (N_25661,N_25015,N_24865);
nor U25662 (N_25662,N_24904,N_25134);
xor U25663 (N_25663,N_24665,N_24852);
or U25664 (N_25664,N_24944,N_25109);
xnor U25665 (N_25665,N_25178,N_25054);
xnor U25666 (N_25666,N_25091,N_24857);
and U25667 (N_25667,N_25165,N_25040);
xnor U25668 (N_25668,N_24844,N_25093);
xor U25669 (N_25669,N_25088,N_25007);
xnor U25670 (N_25670,N_25038,N_24853);
xnor U25671 (N_25671,N_25125,N_25184);
or U25672 (N_25672,N_25022,N_25055);
or U25673 (N_25673,N_25116,N_24926);
xor U25674 (N_25674,N_24681,N_24622);
xnor U25675 (N_25675,N_25187,N_24804);
xnor U25676 (N_25676,N_25101,N_25031);
nand U25677 (N_25677,N_24917,N_25015);
nand U25678 (N_25678,N_25155,N_25146);
and U25679 (N_25679,N_25051,N_25071);
or U25680 (N_25680,N_24666,N_24811);
nor U25681 (N_25681,N_24652,N_25031);
nand U25682 (N_25682,N_24843,N_24657);
nor U25683 (N_25683,N_24842,N_25061);
nand U25684 (N_25684,N_25126,N_24663);
nor U25685 (N_25685,N_24737,N_24956);
nand U25686 (N_25686,N_24808,N_24896);
or U25687 (N_25687,N_25103,N_24737);
and U25688 (N_25688,N_25127,N_24913);
or U25689 (N_25689,N_24681,N_24846);
or U25690 (N_25690,N_24756,N_24929);
nor U25691 (N_25691,N_25107,N_25179);
nor U25692 (N_25692,N_24799,N_24635);
nand U25693 (N_25693,N_24628,N_25004);
or U25694 (N_25694,N_25053,N_24828);
nor U25695 (N_25695,N_24900,N_24984);
nand U25696 (N_25696,N_24699,N_25050);
and U25697 (N_25697,N_24760,N_24729);
and U25698 (N_25698,N_24879,N_24823);
and U25699 (N_25699,N_24771,N_25005);
or U25700 (N_25700,N_24628,N_24623);
nor U25701 (N_25701,N_25159,N_24733);
or U25702 (N_25702,N_25015,N_24626);
nor U25703 (N_25703,N_24741,N_25164);
xor U25704 (N_25704,N_24971,N_24731);
nor U25705 (N_25705,N_25011,N_24990);
or U25706 (N_25706,N_24952,N_24698);
nor U25707 (N_25707,N_24745,N_25130);
or U25708 (N_25708,N_25142,N_24976);
nand U25709 (N_25709,N_25197,N_24995);
nand U25710 (N_25710,N_25063,N_24663);
and U25711 (N_25711,N_24811,N_24608);
and U25712 (N_25712,N_24606,N_24724);
nand U25713 (N_25713,N_25026,N_24684);
nor U25714 (N_25714,N_24945,N_24899);
and U25715 (N_25715,N_25154,N_24756);
nor U25716 (N_25716,N_24623,N_24666);
nor U25717 (N_25717,N_24900,N_25077);
nand U25718 (N_25718,N_25167,N_24884);
and U25719 (N_25719,N_24717,N_24720);
or U25720 (N_25720,N_25182,N_24700);
xor U25721 (N_25721,N_24625,N_25027);
or U25722 (N_25722,N_25021,N_24681);
nand U25723 (N_25723,N_25084,N_25170);
or U25724 (N_25724,N_24839,N_25184);
nor U25725 (N_25725,N_24930,N_24698);
and U25726 (N_25726,N_24932,N_24607);
xnor U25727 (N_25727,N_24614,N_24985);
nand U25728 (N_25728,N_25002,N_25083);
nand U25729 (N_25729,N_24764,N_24650);
or U25730 (N_25730,N_24755,N_25171);
nor U25731 (N_25731,N_25168,N_24741);
and U25732 (N_25732,N_25007,N_24918);
xor U25733 (N_25733,N_24994,N_24667);
and U25734 (N_25734,N_24969,N_25104);
nand U25735 (N_25735,N_25062,N_24699);
or U25736 (N_25736,N_25153,N_24901);
nand U25737 (N_25737,N_24913,N_24938);
nor U25738 (N_25738,N_24986,N_24997);
nand U25739 (N_25739,N_25037,N_25170);
nor U25740 (N_25740,N_24631,N_25124);
and U25741 (N_25741,N_25178,N_24752);
xnor U25742 (N_25742,N_24858,N_24786);
or U25743 (N_25743,N_24983,N_24763);
nand U25744 (N_25744,N_25000,N_25072);
or U25745 (N_25745,N_25018,N_24907);
nor U25746 (N_25746,N_24621,N_24788);
or U25747 (N_25747,N_24721,N_25128);
nor U25748 (N_25748,N_24833,N_24604);
nor U25749 (N_25749,N_24916,N_24897);
xor U25750 (N_25750,N_24730,N_24798);
and U25751 (N_25751,N_24689,N_24973);
nand U25752 (N_25752,N_24639,N_25199);
nand U25753 (N_25753,N_25051,N_24909);
nor U25754 (N_25754,N_25122,N_24738);
or U25755 (N_25755,N_24690,N_24935);
and U25756 (N_25756,N_24810,N_24919);
and U25757 (N_25757,N_25059,N_25161);
and U25758 (N_25758,N_25026,N_25107);
nand U25759 (N_25759,N_24970,N_24663);
and U25760 (N_25760,N_24705,N_24655);
xnor U25761 (N_25761,N_24671,N_24908);
nand U25762 (N_25762,N_24610,N_25068);
or U25763 (N_25763,N_25036,N_24895);
xnor U25764 (N_25764,N_24648,N_24815);
nand U25765 (N_25765,N_25135,N_25012);
nand U25766 (N_25766,N_24950,N_25045);
xor U25767 (N_25767,N_24917,N_24729);
and U25768 (N_25768,N_24675,N_25060);
or U25769 (N_25769,N_24894,N_24869);
nor U25770 (N_25770,N_24707,N_24813);
nand U25771 (N_25771,N_24664,N_24897);
and U25772 (N_25772,N_25090,N_24932);
nand U25773 (N_25773,N_24677,N_24754);
and U25774 (N_25774,N_25061,N_24695);
nand U25775 (N_25775,N_24667,N_24899);
xnor U25776 (N_25776,N_24698,N_24782);
or U25777 (N_25777,N_24835,N_25162);
nand U25778 (N_25778,N_24889,N_24623);
nor U25779 (N_25779,N_24899,N_24828);
or U25780 (N_25780,N_25028,N_24739);
and U25781 (N_25781,N_25164,N_24988);
or U25782 (N_25782,N_24888,N_25063);
and U25783 (N_25783,N_25025,N_25104);
and U25784 (N_25784,N_25073,N_25124);
or U25785 (N_25785,N_24609,N_25114);
xor U25786 (N_25786,N_24778,N_25074);
nand U25787 (N_25787,N_24761,N_24748);
nor U25788 (N_25788,N_25175,N_24738);
and U25789 (N_25789,N_24607,N_24890);
xnor U25790 (N_25790,N_24976,N_24798);
and U25791 (N_25791,N_25152,N_24750);
or U25792 (N_25792,N_24817,N_24864);
or U25793 (N_25793,N_25135,N_24916);
or U25794 (N_25794,N_24779,N_24762);
nor U25795 (N_25795,N_24926,N_24973);
and U25796 (N_25796,N_24720,N_24882);
xor U25797 (N_25797,N_24963,N_25118);
nor U25798 (N_25798,N_25108,N_25027);
nand U25799 (N_25799,N_24956,N_25116);
nand U25800 (N_25800,N_25387,N_25226);
xnor U25801 (N_25801,N_25748,N_25672);
or U25802 (N_25802,N_25573,N_25345);
nor U25803 (N_25803,N_25293,N_25424);
or U25804 (N_25804,N_25227,N_25671);
nor U25805 (N_25805,N_25596,N_25792);
and U25806 (N_25806,N_25525,N_25500);
nand U25807 (N_25807,N_25605,N_25410);
nand U25808 (N_25808,N_25702,N_25287);
or U25809 (N_25809,N_25750,N_25408);
nand U25810 (N_25810,N_25550,N_25274);
and U25811 (N_25811,N_25552,N_25647);
nand U25812 (N_25812,N_25568,N_25349);
and U25813 (N_25813,N_25768,N_25343);
nand U25814 (N_25814,N_25639,N_25317);
nor U25815 (N_25815,N_25609,N_25288);
and U25816 (N_25816,N_25228,N_25704);
nor U25817 (N_25817,N_25480,N_25431);
nand U25818 (N_25818,N_25784,N_25764);
nand U25819 (N_25819,N_25608,N_25323);
xor U25820 (N_25820,N_25307,N_25320);
or U25821 (N_25821,N_25273,N_25300);
nor U25822 (N_25822,N_25236,N_25218);
or U25823 (N_25823,N_25232,N_25225);
nor U25824 (N_25824,N_25423,N_25360);
xnor U25825 (N_25825,N_25467,N_25717);
xor U25826 (N_25826,N_25591,N_25520);
and U25827 (N_25827,N_25673,N_25694);
nand U25828 (N_25828,N_25312,N_25347);
or U25829 (N_25829,N_25526,N_25649);
or U25830 (N_25830,N_25466,N_25384);
or U25831 (N_25831,N_25305,N_25318);
xnor U25832 (N_25832,N_25429,N_25632);
xor U25833 (N_25833,N_25462,N_25353);
or U25834 (N_25834,N_25205,N_25494);
xnor U25835 (N_25835,N_25558,N_25701);
nor U25836 (N_25836,N_25442,N_25635);
nor U25837 (N_25837,N_25269,N_25278);
nor U25838 (N_25838,N_25346,N_25470);
or U25839 (N_25839,N_25251,N_25235);
nor U25840 (N_25840,N_25391,N_25627);
xnor U25841 (N_25841,N_25545,N_25556);
or U25842 (N_25842,N_25219,N_25371);
nand U25843 (N_25843,N_25242,N_25561);
nand U25844 (N_25844,N_25714,N_25341);
xnor U25845 (N_25845,N_25386,N_25711);
nand U25846 (N_25846,N_25450,N_25683);
xor U25847 (N_25847,N_25449,N_25432);
or U25848 (N_25848,N_25472,N_25245);
and U25849 (N_25849,N_25641,N_25490);
nor U25850 (N_25850,N_25652,N_25689);
xor U25851 (N_25851,N_25372,N_25460);
nand U25852 (N_25852,N_25644,N_25769);
xnor U25853 (N_25853,N_25590,N_25565);
nand U25854 (N_25854,N_25262,N_25517);
or U25855 (N_25855,N_25439,N_25741);
xor U25856 (N_25856,N_25633,N_25531);
nand U25857 (N_25857,N_25624,N_25686);
or U25858 (N_25858,N_25660,N_25452);
xnor U25859 (N_25859,N_25420,N_25640);
nor U25860 (N_25860,N_25402,N_25709);
or U25861 (N_25861,N_25752,N_25497);
or U25862 (N_25862,N_25504,N_25285);
nand U25863 (N_25863,N_25326,N_25729);
nand U25864 (N_25864,N_25571,N_25428);
nor U25865 (N_25865,N_25283,N_25398);
and U25866 (N_25866,N_25453,N_25648);
nand U25867 (N_25867,N_25316,N_25418);
xor U25868 (N_25868,N_25629,N_25230);
nor U25869 (N_25869,N_25370,N_25512);
nor U25870 (N_25870,N_25625,N_25478);
nand U25871 (N_25871,N_25679,N_25322);
nor U25872 (N_25872,N_25352,N_25443);
xor U25873 (N_25873,N_25335,N_25518);
nor U25874 (N_25874,N_25770,N_25730);
and U25875 (N_25875,N_25537,N_25581);
or U25876 (N_25876,N_25476,N_25619);
nand U25877 (N_25877,N_25592,N_25297);
nand U25878 (N_25878,N_25749,N_25603);
nand U25879 (N_25879,N_25529,N_25761);
xnor U25880 (N_25880,N_25503,N_25407);
or U25881 (N_25881,N_25358,N_25210);
nand U25882 (N_25882,N_25725,N_25664);
xor U25883 (N_25883,N_25330,N_25502);
or U25884 (N_25884,N_25738,N_25691);
nand U25885 (N_25885,N_25782,N_25217);
and U25886 (N_25886,N_25454,N_25459);
or U25887 (N_25887,N_25206,N_25618);
nor U25888 (N_25888,N_25224,N_25576);
nor U25889 (N_25889,N_25308,N_25744);
and U25890 (N_25890,N_25507,N_25435);
xor U25891 (N_25891,N_25303,N_25703);
or U25892 (N_25892,N_25456,N_25755);
and U25893 (N_25893,N_25549,N_25563);
and U25894 (N_25894,N_25286,N_25298);
nor U25895 (N_25895,N_25250,N_25238);
xor U25896 (N_25896,N_25421,N_25572);
and U25897 (N_25897,N_25374,N_25464);
nand U25898 (N_25898,N_25394,N_25299);
xor U25899 (N_25899,N_25306,N_25515);
nand U25900 (N_25900,N_25513,N_25739);
xnor U25901 (N_25901,N_25787,N_25687);
nor U25902 (N_25902,N_25661,N_25674);
nand U25903 (N_25903,N_25400,N_25636);
nand U25904 (N_25904,N_25570,N_25742);
xnor U25905 (N_25905,N_25366,N_25684);
nand U25906 (N_25906,N_25357,N_25212);
or U25907 (N_25907,N_25759,N_25241);
nand U25908 (N_25908,N_25613,N_25413);
or U25909 (N_25909,N_25446,N_25789);
nand U25910 (N_25910,N_25434,N_25348);
xnor U25911 (N_25911,N_25646,N_25390);
nor U25912 (N_25912,N_25659,N_25707);
or U25913 (N_25913,N_25302,N_25301);
xor U25914 (N_25914,N_25417,N_25536);
xor U25915 (N_25915,N_25488,N_25699);
xnor U25916 (N_25916,N_25597,N_25796);
and U25917 (N_25917,N_25756,N_25240);
nor U25918 (N_25918,N_25334,N_25389);
or U25919 (N_25919,N_25319,N_25261);
nor U25920 (N_25920,N_25700,N_25268);
xnor U25921 (N_25921,N_25766,N_25746);
nand U25922 (N_25922,N_25747,N_25498);
and U25923 (N_25923,N_25406,N_25753);
nor U25924 (N_25924,N_25211,N_25356);
nand U25925 (N_25925,N_25482,N_25680);
and U25926 (N_25926,N_25243,N_25380);
or U25927 (N_25927,N_25617,N_25767);
nand U25928 (N_25928,N_25578,N_25783);
xor U25929 (N_25929,N_25560,N_25339);
xnor U25930 (N_25930,N_25458,N_25595);
and U25931 (N_25931,N_25781,N_25233);
or U25932 (N_25932,N_25760,N_25296);
nand U25933 (N_25933,N_25533,N_25506);
nor U25934 (N_25934,N_25511,N_25495);
or U25935 (N_25935,N_25559,N_25541);
xnor U25936 (N_25936,N_25361,N_25655);
nand U25937 (N_25937,N_25519,N_25788);
nand U25938 (N_25938,N_25209,N_25487);
or U25939 (N_25939,N_25698,N_25732);
nor U25940 (N_25940,N_25682,N_25542);
nor U25941 (N_25941,N_25751,N_25414);
nor U25942 (N_25942,N_25258,N_25292);
or U25943 (N_25943,N_25202,N_25315);
xnor U25944 (N_25944,N_25530,N_25611);
nand U25945 (N_25945,N_25696,N_25589);
nand U25946 (N_25946,N_25416,N_25364);
nor U25947 (N_25947,N_25653,N_25441);
xnor U25948 (N_25948,N_25797,N_25604);
and U25949 (N_25949,N_25616,N_25638);
nand U25950 (N_25950,N_25681,N_25379);
or U25951 (N_25951,N_25486,N_25489);
and U25952 (N_25952,N_25378,N_25575);
xnor U25953 (N_25953,N_25247,N_25675);
and U25954 (N_25954,N_25440,N_25314);
or U25955 (N_25955,N_25257,N_25721);
nor U25956 (N_25956,N_25492,N_25623);
xor U25957 (N_25957,N_25468,N_25282);
or U25958 (N_25958,N_25567,N_25279);
nand U25959 (N_25959,N_25600,N_25309);
or U25960 (N_25960,N_25369,N_25777);
and U25961 (N_25961,N_25255,N_25779);
or U25962 (N_25962,N_25397,N_25514);
xnor U25963 (N_25963,N_25272,N_25667);
and U25964 (N_25964,N_25620,N_25215);
or U25965 (N_25965,N_25697,N_25271);
nand U25966 (N_25966,N_25601,N_25637);
or U25967 (N_25967,N_25291,N_25445);
or U25968 (N_25968,N_25425,N_25252);
nand U25969 (N_25969,N_25485,N_25580);
nor U25970 (N_25970,N_25548,N_25264);
or U25971 (N_25971,N_25728,N_25733);
xnor U25972 (N_25972,N_25794,N_25231);
xnor U25973 (N_25973,N_25574,N_25362);
nand U25974 (N_25974,N_25634,N_25213);
or U25975 (N_25975,N_25260,N_25522);
xnor U25976 (N_25976,N_25535,N_25471);
nor U25977 (N_25977,N_25685,N_25773);
nand U25978 (N_25978,N_25656,N_25363);
and U25979 (N_25979,N_25284,N_25493);
xnor U25980 (N_25980,N_25289,N_25583);
xnor U25981 (N_25981,N_25628,N_25336);
xor U25982 (N_25982,N_25695,N_25277);
or U25983 (N_25983,N_25534,N_25795);
or U25984 (N_25984,N_25731,N_25216);
and U25985 (N_25985,N_25771,N_25722);
or U25986 (N_25986,N_25598,N_25376);
xor U25987 (N_25987,N_25793,N_25607);
or U25988 (N_25988,N_25313,N_25239);
or U25989 (N_25989,N_25724,N_25333);
and U25990 (N_25990,N_25621,N_25355);
xnor U25991 (N_25991,N_25281,N_25203);
xor U25992 (N_25992,N_25393,N_25785);
nand U25993 (N_25993,N_25708,N_25762);
nand U25994 (N_25994,N_25311,N_25246);
nor U25995 (N_25995,N_25521,N_25474);
or U25996 (N_25996,N_25594,N_25321);
nand U25997 (N_25997,N_25373,N_25223);
and U25998 (N_25998,N_25610,N_25587);
xor U25999 (N_25999,N_25713,N_25329);
nand U26000 (N_26000,N_25643,N_25463);
nand U26001 (N_26001,N_25582,N_25658);
and U26002 (N_26002,N_25350,N_25381);
and U26003 (N_26003,N_25564,N_25200);
xnor U26004 (N_26004,N_25479,N_25754);
nand U26005 (N_26005,N_25505,N_25249);
and U26006 (N_26006,N_25715,N_25668);
xnor U26007 (N_26007,N_25662,N_25786);
nor U26008 (N_26008,N_25448,N_25477);
or U26009 (N_26009,N_25774,N_25676);
xor U26010 (N_26010,N_25222,N_25557);
or U26011 (N_26011,N_25651,N_25383);
or U26012 (N_26012,N_25584,N_25745);
nand U26013 (N_26013,N_25392,N_25776);
and U26014 (N_26014,N_25265,N_25555);
or U26015 (N_26015,N_25433,N_25527);
and U26016 (N_26016,N_25221,N_25688);
and U26017 (N_26017,N_25327,N_25275);
nor U26018 (N_26018,N_25365,N_25538);
nor U26019 (N_26019,N_25775,N_25426);
or U26020 (N_26020,N_25422,N_25665);
or U26021 (N_26021,N_25602,N_25670);
xnor U26022 (N_26022,N_25726,N_25528);
or U26023 (N_26023,N_25798,N_25396);
nand U26024 (N_26024,N_25263,N_25267);
nor U26025 (N_26025,N_25657,N_25692);
or U26026 (N_26026,N_25229,N_25510);
and U26027 (N_26027,N_25208,N_25516);
nand U26028 (N_26028,N_25310,N_25340);
xor U26029 (N_26029,N_25585,N_25220);
or U26030 (N_26030,N_25447,N_25588);
xnor U26031 (N_26031,N_25642,N_25735);
nand U26032 (N_26032,N_25399,N_25690);
xor U26033 (N_26033,N_25204,N_25654);
nor U26034 (N_26034,N_25677,N_25693);
or U26035 (N_26035,N_25451,N_25606);
nor U26036 (N_26036,N_25214,N_25259);
xnor U26037 (N_26037,N_25412,N_25740);
and U26038 (N_26038,N_25743,N_25645);
and U26039 (N_26039,N_25405,N_25475);
xnor U26040 (N_26040,N_25562,N_25566);
nor U26041 (N_26041,N_25351,N_25388);
xor U26042 (N_26042,N_25579,N_25551);
xnor U26043 (N_26043,N_25248,N_25473);
and U26044 (N_26044,N_25615,N_25234);
xor U26045 (N_26045,N_25778,N_25201);
and U26046 (N_26046,N_25415,N_25780);
nor U26047 (N_26047,N_25444,N_25716);
nor U26048 (N_26048,N_25622,N_25469);
xnor U26049 (N_26049,N_25501,N_25403);
nor U26050 (N_26050,N_25544,N_25553);
nand U26051 (N_26051,N_25569,N_25280);
xor U26052 (N_26052,N_25719,N_25705);
or U26053 (N_26053,N_25496,N_25491);
or U26054 (N_26054,N_25457,N_25461);
nand U26055 (N_26055,N_25710,N_25546);
nor U26056 (N_26056,N_25437,N_25539);
xnor U26057 (N_26057,N_25266,N_25723);
nand U26058 (N_26058,N_25484,N_25626);
xnor U26059 (N_26059,N_25254,N_25331);
nand U26060 (N_26060,N_25367,N_25455);
nand U26061 (N_26061,N_25509,N_25790);
or U26062 (N_26062,N_25436,N_25324);
or U26063 (N_26063,N_25395,N_25385);
or U26064 (N_26064,N_25409,N_25253);
nor U26065 (N_26065,N_25547,N_25543);
nand U26066 (N_26066,N_25799,N_25337);
or U26067 (N_26067,N_25354,N_25524);
nand U26068 (N_26068,N_25382,N_25359);
xor U26069 (N_26069,N_25772,N_25465);
nor U26070 (N_26070,N_25481,N_25294);
nand U26071 (N_26071,N_25290,N_25207);
or U26072 (N_26072,N_25295,N_25720);
or U26073 (N_26073,N_25758,N_25344);
xnor U26074 (N_26074,N_25411,N_25237);
xnor U26075 (N_26075,N_25430,N_25631);
nand U26076 (N_26076,N_25763,N_25666);
nand U26077 (N_26077,N_25669,N_25325);
nand U26078 (N_26078,N_25523,N_25678);
nor U26079 (N_26079,N_25338,N_25368);
nor U26080 (N_26080,N_25599,N_25377);
nor U26081 (N_26081,N_25404,N_25427);
and U26082 (N_26082,N_25734,N_25499);
and U26083 (N_26083,N_25532,N_25737);
and U26084 (N_26084,N_25718,N_25593);
nand U26085 (N_26085,N_25612,N_25342);
and U26086 (N_26086,N_25375,N_25706);
or U26087 (N_26087,N_25419,N_25256);
nand U26088 (N_26088,N_25332,N_25554);
nor U26089 (N_26089,N_25586,N_25276);
nand U26090 (N_26090,N_25244,N_25540);
and U26091 (N_26091,N_25650,N_25508);
or U26092 (N_26092,N_25791,N_25483);
nand U26093 (N_26093,N_25438,N_25736);
or U26094 (N_26094,N_25614,N_25270);
and U26095 (N_26095,N_25765,N_25630);
and U26096 (N_26096,N_25757,N_25663);
nand U26097 (N_26097,N_25328,N_25727);
or U26098 (N_26098,N_25577,N_25304);
nor U26099 (N_26099,N_25712,N_25401);
xnor U26100 (N_26100,N_25213,N_25548);
and U26101 (N_26101,N_25429,N_25508);
and U26102 (N_26102,N_25262,N_25236);
and U26103 (N_26103,N_25253,N_25574);
and U26104 (N_26104,N_25503,N_25394);
nand U26105 (N_26105,N_25434,N_25554);
or U26106 (N_26106,N_25529,N_25203);
or U26107 (N_26107,N_25216,N_25243);
nand U26108 (N_26108,N_25385,N_25294);
and U26109 (N_26109,N_25790,N_25652);
xor U26110 (N_26110,N_25227,N_25657);
or U26111 (N_26111,N_25783,N_25201);
nor U26112 (N_26112,N_25608,N_25382);
or U26113 (N_26113,N_25251,N_25249);
nor U26114 (N_26114,N_25786,N_25208);
xnor U26115 (N_26115,N_25516,N_25755);
and U26116 (N_26116,N_25585,N_25313);
nor U26117 (N_26117,N_25715,N_25645);
and U26118 (N_26118,N_25797,N_25774);
nand U26119 (N_26119,N_25329,N_25626);
xor U26120 (N_26120,N_25480,N_25325);
or U26121 (N_26121,N_25456,N_25642);
nor U26122 (N_26122,N_25761,N_25462);
nand U26123 (N_26123,N_25753,N_25512);
xor U26124 (N_26124,N_25604,N_25741);
xor U26125 (N_26125,N_25516,N_25586);
nor U26126 (N_26126,N_25377,N_25573);
or U26127 (N_26127,N_25785,N_25247);
nor U26128 (N_26128,N_25757,N_25772);
nand U26129 (N_26129,N_25604,N_25312);
or U26130 (N_26130,N_25676,N_25568);
nor U26131 (N_26131,N_25298,N_25307);
nor U26132 (N_26132,N_25613,N_25407);
nor U26133 (N_26133,N_25351,N_25355);
xnor U26134 (N_26134,N_25593,N_25716);
nor U26135 (N_26135,N_25395,N_25275);
nor U26136 (N_26136,N_25783,N_25369);
or U26137 (N_26137,N_25628,N_25247);
nor U26138 (N_26138,N_25681,N_25706);
and U26139 (N_26139,N_25333,N_25229);
xor U26140 (N_26140,N_25307,N_25347);
nor U26141 (N_26141,N_25326,N_25769);
nand U26142 (N_26142,N_25323,N_25553);
xor U26143 (N_26143,N_25409,N_25376);
xor U26144 (N_26144,N_25559,N_25680);
and U26145 (N_26145,N_25465,N_25339);
xor U26146 (N_26146,N_25423,N_25637);
or U26147 (N_26147,N_25259,N_25257);
xor U26148 (N_26148,N_25755,N_25391);
xor U26149 (N_26149,N_25736,N_25308);
nor U26150 (N_26150,N_25607,N_25323);
nor U26151 (N_26151,N_25432,N_25412);
nand U26152 (N_26152,N_25263,N_25273);
and U26153 (N_26153,N_25768,N_25234);
and U26154 (N_26154,N_25671,N_25255);
nand U26155 (N_26155,N_25607,N_25542);
nand U26156 (N_26156,N_25392,N_25551);
and U26157 (N_26157,N_25293,N_25704);
nor U26158 (N_26158,N_25730,N_25523);
and U26159 (N_26159,N_25509,N_25783);
xor U26160 (N_26160,N_25385,N_25552);
nand U26161 (N_26161,N_25417,N_25332);
nand U26162 (N_26162,N_25536,N_25754);
xnor U26163 (N_26163,N_25691,N_25709);
nor U26164 (N_26164,N_25279,N_25537);
nand U26165 (N_26165,N_25444,N_25375);
nand U26166 (N_26166,N_25705,N_25514);
nor U26167 (N_26167,N_25774,N_25710);
xor U26168 (N_26168,N_25234,N_25469);
or U26169 (N_26169,N_25674,N_25301);
or U26170 (N_26170,N_25651,N_25664);
and U26171 (N_26171,N_25630,N_25625);
xnor U26172 (N_26172,N_25443,N_25427);
or U26173 (N_26173,N_25541,N_25793);
nor U26174 (N_26174,N_25236,N_25765);
and U26175 (N_26175,N_25400,N_25782);
and U26176 (N_26176,N_25428,N_25654);
or U26177 (N_26177,N_25581,N_25579);
nand U26178 (N_26178,N_25277,N_25405);
nor U26179 (N_26179,N_25636,N_25550);
xnor U26180 (N_26180,N_25399,N_25363);
nor U26181 (N_26181,N_25252,N_25236);
and U26182 (N_26182,N_25709,N_25334);
nor U26183 (N_26183,N_25565,N_25783);
or U26184 (N_26184,N_25316,N_25704);
and U26185 (N_26185,N_25217,N_25576);
or U26186 (N_26186,N_25758,N_25317);
or U26187 (N_26187,N_25209,N_25235);
or U26188 (N_26188,N_25786,N_25216);
nand U26189 (N_26189,N_25404,N_25288);
nor U26190 (N_26190,N_25357,N_25234);
xnor U26191 (N_26191,N_25317,N_25554);
nand U26192 (N_26192,N_25374,N_25599);
nand U26193 (N_26193,N_25408,N_25534);
nor U26194 (N_26194,N_25454,N_25479);
xnor U26195 (N_26195,N_25574,N_25747);
nand U26196 (N_26196,N_25525,N_25300);
nor U26197 (N_26197,N_25345,N_25647);
xnor U26198 (N_26198,N_25724,N_25649);
xnor U26199 (N_26199,N_25564,N_25213);
xnor U26200 (N_26200,N_25594,N_25201);
and U26201 (N_26201,N_25770,N_25576);
and U26202 (N_26202,N_25419,N_25585);
nand U26203 (N_26203,N_25424,N_25462);
xor U26204 (N_26204,N_25348,N_25564);
or U26205 (N_26205,N_25381,N_25234);
xor U26206 (N_26206,N_25633,N_25648);
and U26207 (N_26207,N_25387,N_25284);
or U26208 (N_26208,N_25428,N_25223);
nor U26209 (N_26209,N_25523,N_25560);
and U26210 (N_26210,N_25295,N_25320);
xor U26211 (N_26211,N_25206,N_25353);
nand U26212 (N_26212,N_25367,N_25622);
nor U26213 (N_26213,N_25579,N_25698);
and U26214 (N_26214,N_25483,N_25588);
and U26215 (N_26215,N_25585,N_25525);
and U26216 (N_26216,N_25232,N_25515);
nand U26217 (N_26217,N_25226,N_25204);
or U26218 (N_26218,N_25658,N_25538);
nand U26219 (N_26219,N_25629,N_25483);
nand U26220 (N_26220,N_25585,N_25634);
xor U26221 (N_26221,N_25580,N_25669);
nor U26222 (N_26222,N_25730,N_25541);
and U26223 (N_26223,N_25431,N_25398);
nand U26224 (N_26224,N_25366,N_25347);
nand U26225 (N_26225,N_25362,N_25419);
nor U26226 (N_26226,N_25298,N_25375);
xor U26227 (N_26227,N_25615,N_25237);
xor U26228 (N_26228,N_25354,N_25390);
and U26229 (N_26229,N_25561,N_25609);
xnor U26230 (N_26230,N_25459,N_25589);
xnor U26231 (N_26231,N_25552,N_25702);
and U26232 (N_26232,N_25575,N_25456);
or U26233 (N_26233,N_25557,N_25512);
nor U26234 (N_26234,N_25473,N_25491);
and U26235 (N_26235,N_25706,N_25597);
and U26236 (N_26236,N_25773,N_25536);
xor U26237 (N_26237,N_25451,N_25360);
nor U26238 (N_26238,N_25599,N_25438);
nand U26239 (N_26239,N_25677,N_25481);
xnor U26240 (N_26240,N_25289,N_25374);
xnor U26241 (N_26241,N_25333,N_25676);
xor U26242 (N_26242,N_25747,N_25450);
or U26243 (N_26243,N_25736,N_25618);
nor U26244 (N_26244,N_25767,N_25446);
or U26245 (N_26245,N_25385,N_25397);
or U26246 (N_26246,N_25598,N_25751);
and U26247 (N_26247,N_25407,N_25669);
xnor U26248 (N_26248,N_25617,N_25691);
and U26249 (N_26249,N_25233,N_25329);
nand U26250 (N_26250,N_25459,N_25260);
nand U26251 (N_26251,N_25655,N_25550);
xor U26252 (N_26252,N_25438,N_25733);
and U26253 (N_26253,N_25624,N_25358);
nand U26254 (N_26254,N_25505,N_25545);
and U26255 (N_26255,N_25489,N_25231);
nor U26256 (N_26256,N_25724,N_25653);
nor U26257 (N_26257,N_25451,N_25785);
and U26258 (N_26258,N_25505,N_25264);
nand U26259 (N_26259,N_25316,N_25298);
or U26260 (N_26260,N_25353,N_25243);
or U26261 (N_26261,N_25465,N_25701);
and U26262 (N_26262,N_25729,N_25338);
xor U26263 (N_26263,N_25541,N_25330);
nor U26264 (N_26264,N_25628,N_25299);
and U26265 (N_26265,N_25459,N_25554);
xnor U26266 (N_26266,N_25697,N_25427);
nor U26267 (N_26267,N_25314,N_25634);
nand U26268 (N_26268,N_25648,N_25320);
or U26269 (N_26269,N_25703,N_25312);
xnor U26270 (N_26270,N_25427,N_25562);
or U26271 (N_26271,N_25758,N_25390);
xnor U26272 (N_26272,N_25549,N_25290);
or U26273 (N_26273,N_25397,N_25791);
and U26274 (N_26274,N_25265,N_25724);
and U26275 (N_26275,N_25465,N_25633);
and U26276 (N_26276,N_25652,N_25584);
xor U26277 (N_26277,N_25249,N_25210);
or U26278 (N_26278,N_25575,N_25614);
nor U26279 (N_26279,N_25491,N_25714);
xor U26280 (N_26280,N_25758,N_25639);
nor U26281 (N_26281,N_25555,N_25232);
or U26282 (N_26282,N_25394,N_25293);
nor U26283 (N_26283,N_25485,N_25767);
or U26284 (N_26284,N_25438,N_25794);
xnor U26285 (N_26285,N_25217,N_25506);
xor U26286 (N_26286,N_25323,N_25252);
nand U26287 (N_26287,N_25381,N_25679);
or U26288 (N_26288,N_25216,N_25398);
xnor U26289 (N_26289,N_25390,N_25338);
nand U26290 (N_26290,N_25590,N_25278);
nand U26291 (N_26291,N_25740,N_25289);
nand U26292 (N_26292,N_25275,N_25610);
nor U26293 (N_26293,N_25742,N_25787);
xnor U26294 (N_26294,N_25600,N_25517);
and U26295 (N_26295,N_25567,N_25696);
nand U26296 (N_26296,N_25317,N_25265);
nor U26297 (N_26297,N_25348,N_25600);
nor U26298 (N_26298,N_25611,N_25672);
nand U26299 (N_26299,N_25220,N_25404);
nor U26300 (N_26300,N_25414,N_25709);
nand U26301 (N_26301,N_25614,N_25387);
nor U26302 (N_26302,N_25631,N_25745);
and U26303 (N_26303,N_25528,N_25329);
nor U26304 (N_26304,N_25350,N_25457);
xnor U26305 (N_26305,N_25317,N_25771);
xor U26306 (N_26306,N_25566,N_25392);
xnor U26307 (N_26307,N_25408,N_25345);
nor U26308 (N_26308,N_25432,N_25361);
or U26309 (N_26309,N_25253,N_25358);
or U26310 (N_26310,N_25374,N_25213);
and U26311 (N_26311,N_25477,N_25615);
and U26312 (N_26312,N_25798,N_25462);
or U26313 (N_26313,N_25290,N_25651);
xor U26314 (N_26314,N_25610,N_25302);
and U26315 (N_26315,N_25389,N_25635);
nand U26316 (N_26316,N_25275,N_25483);
xor U26317 (N_26317,N_25430,N_25205);
nand U26318 (N_26318,N_25286,N_25462);
nand U26319 (N_26319,N_25214,N_25594);
and U26320 (N_26320,N_25385,N_25564);
and U26321 (N_26321,N_25692,N_25616);
nand U26322 (N_26322,N_25382,N_25595);
xnor U26323 (N_26323,N_25617,N_25238);
nor U26324 (N_26324,N_25207,N_25695);
nand U26325 (N_26325,N_25431,N_25512);
and U26326 (N_26326,N_25725,N_25350);
and U26327 (N_26327,N_25631,N_25569);
and U26328 (N_26328,N_25285,N_25513);
or U26329 (N_26329,N_25457,N_25570);
or U26330 (N_26330,N_25346,N_25635);
xor U26331 (N_26331,N_25522,N_25640);
nor U26332 (N_26332,N_25259,N_25274);
or U26333 (N_26333,N_25648,N_25418);
or U26334 (N_26334,N_25431,N_25348);
and U26335 (N_26335,N_25694,N_25369);
xor U26336 (N_26336,N_25542,N_25481);
nor U26337 (N_26337,N_25505,N_25575);
nand U26338 (N_26338,N_25556,N_25770);
xnor U26339 (N_26339,N_25617,N_25591);
xnor U26340 (N_26340,N_25446,N_25729);
and U26341 (N_26341,N_25683,N_25417);
nor U26342 (N_26342,N_25700,N_25317);
nand U26343 (N_26343,N_25604,N_25520);
nor U26344 (N_26344,N_25501,N_25344);
nand U26345 (N_26345,N_25758,N_25325);
nor U26346 (N_26346,N_25733,N_25359);
xnor U26347 (N_26347,N_25749,N_25376);
or U26348 (N_26348,N_25265,N_25534);
or U26349 (N_26349,N_25509,N_25296);
and U26350 (N_26350,N_25200,N_25570);
and U26351 (N_26351,N_25328,N_25469);
nand U26352 (N_26352,N_25626,N_25544);
and U26353 (N_26353,N_25279,N_25339);
xor U26354 (N_26354,N_25690,N_25311);
xnor U26355 (N_26355,N_25617,N_25235);
nor U26356 (N_26356,N_25208,N_25641);
nor U26357 (N_26357,N_25593,N_25234);
nand U26358 (N_26358,N_25356,N_25694);
nand U26359 (N_26359,N_25327,N_25630);
xnor U26360 (N_26360,N_25347,N_25299);
xnor U26361 (N_26361,N_25730,N_25564);
xor U26362 (N_26362,N_25706,N_25622);
nor U26363 (N_26363,N_25613,N_25288);
or U26364 (N_26364,N_25741,N_25715);
nor U26365 (N_26365,N_25543,N_25312);
nor U26366 (N_26366,N_25301,N_25348);
xnor U26367 (N_26367,N_25429,N_25247);
xor U26368 (N_26368,N_25289,N_25491);
xor U26369 (N_26369,N_25234,N_25585);
nand U26370 (N_26370,N_25215,N_25736);
or U26371 (N_26371,N_25583,N_25481);
nand U26372 (N_26372,N_25528,N_25539);
xnor U26373 (N_26373,N_25272,N_25762);
or U26374 (N_26374,N_25785,N_25523);
nand U26375 (N_26375,N_25647,N_25506);
xor U26376 (N_26376,N_25745,N_25458);
xnor U26377 (N_26377,N_25225,N_25586);
or U26378 (N_26378,N_25254,N_25461);
nand U26379 (N_26379,N_25385,N_25575);
nand U26380 (N_26380,N_25462,N_25491);
xnor U26381 (N_26381,N_25471,N_25422);
nor U26382 (N_26382,N_25264,N_25716);
nor U26383 (N_26383,N_25386,N_25406);
or U26384 (N_26384,N_25290,N_25514);
or U26385 (N_26385,N_25676,N_25769);
nand U26386 (N_26386,N_25384,N_25530);
or U26387 (N_26387,N_25350,N_25640);
nand U26388 (N_26388,N_25640,N_25298);
nor U26389 (N_26389,N_25445,N_25356);
and U26390 (N_26390,N_25761,N_25657);
or U26391 (N_26391,N_25450,N_25236);
xor U26392 (N_26392,N_25761,N_25400);
xnor U26393 (N_26393,N_25627,N_25217);
or U26394 (N_26394,N_25479,N_25612);
and U26395 (N_26395,N_25242,N_25705);
and U26396 (N_26396,N_25736,N_25302);
nand U26397 (N_26397,N_25276,N_25557);
xnor U26398 (N_26398,N_25706,N_25240);
or U26399 (N_26399,N_25578,N_25503);
or U26400 (N_26400,N_26125,N_26345);
and U26401 (N_26401,N_26235,N_26129);
nor U26402 (N_26402,N_26295,N_25814);
xnor U26403 (N_26403,N_26180,N_26124);
xor U26404 (N_26404,N_26261,N_26111);
or U26405 (N_26405,N_25960,N_26285);
nor U26406 (N_26406,N_26387,N_25949);
nor U26407 (N_26407,N_26341,N_25815);
or U26408 (N_26408,N_26205,N_26234);
and U26409 (N_26409,N_26031,N_26242);
nor U26410 (N_26410,N_26147,N_26077);
xor U26411 (N_26411,N_25942,N_25989);
or U26412 (N_26412,N_25947,N_26184);
xor U26413 (N_26413,N_25857,N_26193);
and U26414 (N_26414,N_25958,N_26231);
and U26415 (N_26415,N_26136,N_26220);
xnor U26416 (N_26416,N_26130,N_26068);
xor U26417 (N_26417,N_26300,N_26064);
xor U26418 (N_26418,N_26066,N_26095);
nor U26419 (N_26419,N_26099,N_26097);
nand U26420 (N_26420,N_25931,N_26360);
nor U26421 (N_26421,N_26380,N_26358);
xor U26422 (N_26422,N_25850,N_26286);
nor U26423 (N_26423,N_25856,N_26128);
nor U26424 (N_26424,N_26011,N_26094);
or U26425 (N_26425,N_26185,N_26246);
nand U26426 (N_26426,N_26154,N_26116);
nor U26427 (N_26427,N_26119,N_26354);
and U26428 (N_26428,N_25811,N_26148);
or U26429 (N_26429,N_26227,N_26103);
nand U26430 (N_26430,N_26115,N_25859);
and U26431 (N_26431,N_26229,N_26023);
or U26432 (N_26432,N_26336,N_26056);
xnor U26433 (N_26433,N_26057,N_26118);
nand U26434 (N_26434,N_26054,N_26112);
and U26435 (N_26435,N_26046,N_26212);
xor U26436 (N_26436,N_26014,N_26133);
or U26437 (N_26437,N_26313,N_26203);
xnor U26438 (N_26438,N_26319,N_25844);
xnor U26439 (N_26439,N_26135,N_26196);
nand U26440 (N_26440,N_26101,N_25955);
nor U26441 (N_26441,N_25914,N_25800);
or U26442 (N_26442,N_26252,N_26140);
or U26443 (N_26443,N_26236,N_25943);
xnor U26444 (N_26444,N_26176,N_26038);
or U26445 (N_26445,N_26204,N_25847);
xnor U26446 (N_26446,N_25801,N_26330);
xnor U26447 (N_26447,N_26157,N_25845);
xnor U26448 (N_26448,N_26131,N_26343);
or U26449 (N_26449,N_26257,N_25889);
and U26450 (N_26450,N_26039,N_26164);
or U26451 (N_26451,N_26312,N_26108);
nand U26452 (N_26452,N_26379,N_26316);
or U26453 (N_26453,N_25918,N_25839);
or U26454 (N_26454,N_26017,N_26183);
nor U26455 (N_26455,N_26156,N_26155);
xor U26456 (N_26456,N_26211,N_26069);
nand U26457 (N_26457,N_26318,N_25997);
or U26458 (N_26458,N_25954,N_25974);
nor U26459 (N_26459,N_25988,N_26262);
or U26460 (N_26460,N_26320,N_26375);
nor U26461 (N_26461,N_26144,N_26059);
nand U26462 (N_26462,N_26292,N_26134);
xor U26463 (N_26463,N_25925,N_26092);
xor U26464 (N_26464,N_26329,N_26090);
nor U26465 (N_26465,N_26363,N_26350);
xor U26466 (N_26466,N_26137,N_26141);
and U26467 (N_26467,N_26289,N_26171);
xor U26468 (N_26468,N_26160,N_26338);
nand U26469 (N_26469,N_26009,N_26047);
and U26470 (N_26470,N_26361,N_26079);
xor U26471 (N_26471,N_26273,N_26091);
xor U26472 (N_26472,N_26248,N_26041);
nor U26473 (N_26473,N_25902,N_25977);
nor U26474 (N_26474,N_26332,N_26163);
and U26475 (N_26475,N_25933,N_25895);
nand U26476 (N_26476,N_26226,N_26384);
nand U26477 (N_26477,N_25817,N_25904);
xor U26478 (N_26478,N_26310,N_26333);
nand U26479 (N_26479,N_26007,N_25872);
xor U26480 (N_26480,N_26051,N_26238);
xnor U26481 (N_26481,N_26207,N_25978);
or U26482 (N_26482,N_25877,N_26269);
nand U26483 (N_26483,N_26277,N_26049);
or U26484 (N_26484,N_26357,N_25951);
or U26485 (N_26485,N_26355,N_25948);
nor U26486 (N_26486,N_26278,N_26142);
nand U26487 (N_26487,N_25881,N_26087);
or U26488 (N_26488,N_26394,N_25831);
nor U26489 (N_26489,N_26325,N_26383);
nand U26490 (N_26490,N_25963,N_25897);
and U26491 (N_26491,N_26048,N_25874);
nand U26492 (N_26492,N_25803,N_26388);
nand U26493 (N_26493,N_26399,N_26071);
or U26494 (N_26494,N_25972,N_25980);
nand U26495 (N_26495,N_26398,N_26178);
xor U26496 (N_26496,N_26143,N_25910);
or U26497 (N_26497,N_26194,N_26233);
or U26498 (N_26498,N_25990,N_25998);
nand U26499 (N_26499,N_26058,N_26179);
xor U26500 (N_26500,N_25810,N_26121);
or U26501 (N_26501,N_25905,N_26139);
and U26502 (N_26502,N_26377,N_26224);
and U26503 (N_26503,N_25861,N_25827);
or U26504 (N_26504,N_25940,N_26372);
nand U26505 (N_26505,N_26020,N_26065);
nor U26506 (N_26506,N_26362,N_25808);
and U26507 (N_26507,N_26279,N_25858);
nand U26508 (N_26508,N_26188,N_26282);
nand U26509 (N_26509,N_26003,N_26368);
nand U26510 (N_26510,N_26168,N_26067);
xnor U26511 (N_26511,N_25982,N_26018);
and U26512 (N_26512,N_25876,N_26309);
and U26513 (N_26513,N_26335,N_26053);
or U26514 (N_26514,N_26022,N_25934);
nor U26515 (N_26515,N_26166,N_25860);
nor U26516 (N_26516,N_26264,N_26382);
or U26517 (N_26517,N_26214,N_26305);
nand U26518 (N_26518,N_26240,N_25991);
xnor U26519 (N_26519,N_25953,N_26173);
and U26520 (N_26520,N_25921,N_26352);
nand U26521 (N_26521,N_26237,N_25941);
and U26522 (N_26522,N_25888,N_25926);
xnor U26523 (N_26523,N_26271,N_26311);
xor U26524 (N_26524,N_26146,N_25986);
and U26525 (N_26525,N_26367,N_26322);
or U26526 (N_26526,N_26317,N_25944);
or U26527 (N_26527,N_26082,N_26202);
nand U26528 (N_26528,N_26192,N_26026);
nor U26529 (N_26529,N_26089,N_26102);
nand U26530 (N_26530,N_26172,N_26274);
nand U26531 (N_26531,N_26169,N_25984);
or U26532 (N_26532,N_26323,N_26307);
and U26533 (N_26533,N_26288,N_26113);
and U26534 (N_26534,N_25824,N_26037);
and U26535 (N_26535,N_25936,N_26258);
or U26536 (N_26536,N_25883,N_25959);
nor U26537 (N_26537,N_25821,N_25832);
nand U26538 (N_26538,N_26221,N_26138);
nand U26539 (N_26539,N_25976,N_25983);
xor U26540 (N_26540,N_26199,N_26019);
or U26541 (N_26541,N_26050,N_25923);
nand U26542 (N_26542,N_26063,N_26287);
nand U26543 (N_26543,N_26344,N_26025);
and U26544 (N_26544,N_26356,N_25915);
or U26545 (N_26545,N_26189,N_26086);
and U26546 (N_26546,N_26337,N_26085);
nor U26547 (N_26547,N_26013,N_26396);
and U26548 (N_26548,N_25884,N_25927);
and U26549 (N_26549,N_25891,N_26251);
nand U26550 (N_26550,N_26353,N_26359);
xnor U26551 (N_26551,N_26104,N_26346);
or U26552 (N_26552,N_25946,N_26216);
and U26553 (N_26553,N_26072,N_25994);
nand U26554 (N_26554,N_26306,N_26215);
nand U26555 (N_26555,N_26392,N_26109);
or U26556 (N_26556,N_25967,N_26145);
and U26557 (N_26557,N_26161,N_26210);
xnor U26558 (N_26558,N_25968,N_25819);
nand U26559 (N_26559,N_26008,N_26348);
and U26560 (N_26560,N_26206,N_26078);
xor U26561 (N_26561,N_26244,N_25820);
and U26562 (N_26562,N_25855,N_26098);
or U26563 (N_26563,N_25893,N_25909);
or U26564 (N_26564,N_26106,N_26324);
and U26565 (N_26565,N_26120,N_26021);
xor U26566 (N_26566,N_25818,N_26107);
and U26567 (N_26567,N_25912,N_26123);
nor U26568 (N_26568,N_25842,N_26364);
xnor U26569 (N_26569,N_26314,N_26159);
or U26570 (N_26570,N_26393,N_25939);
nor U26571 (N_26571,N_26281,N_26239);
nor U26572 (N_26572,N_25836,N_25826);
or U26573 (N_26573,N_25981,N_25894);
and U26574 (N_26574,N_26061,N_25837);
nor U26575 (N_26575,N_26030,N_26042);
xor U26576 (N_26576,N_25813,N_25825);
and U26577 (N_26577,N_25999,N_25922);
xnor U26578 (N_26578,N_26076,N_26397);
nand U26579 (N_26579,N_25829,N_25885);
and U26580 (N_26580,N_26122,N_26339);
xnor U26581 (N_26581,N_26186,N_25805);
nor U26582 (N_26582,N_26075,N_26044);
xor U26583 (N_26583,N_25812,N_26386);
nor U26584 (N_26584,N_26187,N_25966);
and U26585 (N_26585,N_25880,N_25864);
nand U26586 (N_26586,N_25961,N_25870);
nor U26587 (N_26587,N_26293,N_26303);
xor U26588 (N_26588,N_25804,N_26218);
or U26589 (N_26589,N_26084,N_26035);
nand U26590 (N_26590,N_25892,N_25971);
and U26591 (N_26591,N_26016,N_26126);
xor U26592 (N_26592,N_26223,N_25848);
and U26593 (N_26593,N_26028,N_26254);
or U26594 (N_26594,N_26340,N_25950);
or U26595 (N_26595,N_25957,N_26055);
and U26596 (N_26596,N_26149,N_25962);
or U26597 (N_26597,N_26073,N_25873);
and U26598 (N_26598,N_25830,N_25928);
xor U26599 (N_26599,N_26225,N_26297);
and U26600 (N_26600,N_25913,N_26391);
xor U26601 (N_26601,N_26032,N_26284);
nor U26602 (N_26602,N_26191,N_25979);
nor U26603 (N_26603,N_26280,N_26342);
nor U26604 (N_26604,N_26291,N_25816);
or U26605 (N_26605,N_26243,N_26152);
nor U26606 (N_26606,N_25935,N_26083);
or U26607 (N_26607,N_25866,N_25996);
nand U26608 (N_26608,N_26177,N_26001);
nand U26609 (N_26609,N_26249,N_26381);
and U26610 (N_26610,N_26250,N_26209);
or U26611 (N_26611,N_26158,N_26181);
or U26612 (N_26612,N_26256,N_26349);
nor U26613 (N_26613,N_26081,N_25882);
nand U26614 (N_26614,N_26331,N_26114);
and U26615 (N_26615,N_25901,N_26190);
nor U26616 (N_26616,N_26040,N_25840);
nand U26617 (N_26617,N_25841,N_26245);
and U26618 (N_26618,N_26217,N_26000);
xnor U26619 (N_26619,N_25863,N_26005);
nand U26620 (N_26620,N_25956,N_26230);
and U26621 (N_26621,N_26389,N_25865);
or U26622 (N_26622,N_26365,N_26270);
and U26623 (N_26623,N_26298,N_26010);
nand U26624 (N_26624,N_26347,N_26027);
nor U26625 (N_26625,N_26308,N_26167);
nand U26626 (N_26626,N_25993,N_26219);
nand U26627 (N_26627,N_25930,N_26299);
and U26628 (N_26628,N_25992,N_26110);
nand U26629 (N_26629,N_26296,N_25908);
and U26630 (N_26630,N_25973,N_26247);
or U26631 (N_26631,N_26132,N_26029);
xnor U26632 (N_26632,N_26033,N_25806);
xor U26633 (N_26633,N_26060,N_26117);
or U26634 (N_26634,N_25890,N_25965);
or U26635 (N_26635,N_25900,N_26222);
and U26636 (N_26636,N_26150,N_26200);
nor U26637 (N_26637,N_26376,N_25838);
or U26638 (N_26638,N_25867,N_25929);
nand U26639 (N_26639,N_25906,N_25851);
and U26640 (N_26640,N_26294,N_25987);
xor U26641 (N_26641,N_25833,N_25969);
or U26642 (N_26642,N_25834,N_26267);
or U26643 (N_26643,N_25809,N_26321);
xnor U26644 (N_26644,N_26265,N_25869);
and U26645 (N_26645,N_25970,N_25896);
nand U26646 (N_26646,N_26174,N_25924);
xnor U26647 (N_26647,N_25995,N_25862);
nor U26648 (N_26648,N_26370,N_25852);
nand U26649 (N_26649,N_25879,N_26232);
nand U26650 (N_26650,N_26198,N_25907);
and U26651 (N_26651,N_26328,N_26283);
nor U26652 (N_26652,N_26062,N_26395);
xnor U26653 (N_26653,N_26276,N_26070);
and U26654 (N_26654,N_26045,N_25916);
xnor U26655 (N_26655,N_26385,N_25846);
xnor U26656 (N_26656,N_26260,N_25886);
nand U26657 (N_26657,N_25964,N_26228);
or U26658 (N_26658,N_26096,N_26182);
and U26659 (N_26659,N_26213,N_26201);
nand U26660 (N_26660,N_26170,N_26052);
and U26661 (N_26661,N_26351,N_26366);
or U26662 (N_26662,N_26074,N_25854);
or U26663 (N_26663,N_26105,N_26100);
xnor U26664 (N_26664,N_25899,N_25878);
and U26665 (N_26665,N_26259,N_26012);
xnor U26666 (N_26666,N_25932,N_26327);
nand U26667 (N_26667,N_25938,N_26275);
nand U26668 (N_26668,N_26127,N_26374);
xnor U26669 (N_26669,N_26290,N_26263);
nor U26670 (N_26670,N_26315,N_26015);
nor U26671 (N_26671,N_26304,N_26301);
nor U26672 (N_26672,N_26253,N_26151);
nand U26673 (N_26673,N_26002,N_25828);
xor U26674 (N_26674,N_26268,N_25849);
nand U26675 (N_26675,N_26165,N_26334);
or U26676 (N_26676,N_26266,N_25871);
and U26677 (N_26677,N_25975,N_25822);
nand U26678 (N_26678,N_26093,N_26080);
or U26679 (N_26679,N_26034,N_25911);
or U26680 (N_26680,N_26153,N_25903);
nand U26681 (N_26681,N_25898,N_25945);
or U26682 (N_26682,N_25920,N_25985);
or U26683 (N_26683,N_26272,N_25868);
xor U26684 (N_26684,N_25917,N_26036);
nor U26685 (N_26685,N_26378,N_26043);
nor U26686 (N_26686,N_26302,N_26024);
and U26687 (N_26687,N_26162,N_25919);
and U26688 (N_26688,N_25835,N_25807);
nor U26689 (N_26689,N_25853,N_26326);
and U26690 (N_26690,N_26241,N_26175);
nor U26691 (N_26691,N_25952,N_26208);
nand U26692 (N_26692,N_26195,N_26371);
nand U26693 (N_26693,N_25875,N_26369);
nor U26694 (N_26694,N_25887,N_25843);
and U26695 (N_26695,N_26006,N_26088);
or U26696 (N_26696,N_26255,N_25823);
nor U26697 (N_26697,N_26373,N_26004);
nand U26698 (N_26698,N_25802,N_25937);
nor U26699 (N_26699,N_26390,N_26197);
and U26700 (N_26700,N_25832,N_26000);
or U26701 (N_26701,N_26047,N_25997);
xor U26702 (N_26702,N_25919,N_25920);
or U26703 (N_26703,N_26169,N_26170);
or U26704 (N_26704,N_26252,N_25986);
and U26705 (N_26705,N_25854,N_26019);
and U26706 (N_26706,N_25872,N_25997);
or U26707 (N_26707,N_25962,N_25900);
xor U26708 (N_26708,N_26220,N_26272);
nor U26709 (N_26709,N_25982,N_26374);
and U26710 (N_26710,N_25984,N_26036);
or U26711 (N_26711,N_26215,N_26235);
nand U26712 (N_26712,N_25849,N_26133);
or U26713 (N_26713,N_26284,N_26116);
nand U26714 (N_26714,N_26261,N_26087);
or U26715 (N_26715,N_26084,N_26110);
nor U26716 (N_26716,N_26036,N_26211);
or U26717 (N_26717,N_25992,N_26298);
or U26718 (N_26718,N_26000,N_25886);
nand U26719 (N_26719,N_26280,N_26021);
or U26720 (N_26720,N_25863,N_26385);
xnor U26721 (N_26721,N_26062,N_26187);
nor U26722 (N_26722,N_26060,N_26187);
and U26723 (N_26723,N_26222,N_26133);
or U26724 (N_26724,N_25951,N_26295);
xnor U26725 (N_26725,N_26188,N_26146);
and U26726 (N_26726,N_26255,N_25930);
nor U26727 (N_26727,N_26283,N_25891);
nor U26728 (N_26728,N_26183,N_25836);
xor U26729 (N_26729,N_26226,N_26110);
nand U26730 (N_26730,N_26262,N_26040);
or U26731 (N_26731,N_26081,N_25942);
or U26732 (N_26732,N_26089,N_26042);
or U26733 (N_26733,N_26061,N_26122);
nand U26734 (N_26734,N_26248,N_26219);
or U26735 (N_26735,N_25845,N_26345);
nand U26736 (N_26736,N_26026,N_25841);
xor U26737 (N_26737,N_26376,N_26373);
nor U26738 (N_26738,N_25940,N_26218);
nand U26739 (N_26739,N_26258,N_26272);
nand U26740 (N_26740,N_26101,N_25870);
or U26741 (N_26741,N_26069,N_26114);
nand U26742 (N_26742,N_25802,N_26004);
xnor U26743 (N_26743,N_26063,N_26163);
nor U26744 (N_26744,N_26077,N_25910);
and U26745 (N_26745,N_26155,N_26150);
nor U26746 (N_26746,N_26159,N_25817);
xnor U26747 (N_26747,N_25841,N_25994);
and U26748 (N_26748,N_26353,N_25818);
xnor U26749 (N_26749,N_25983,N_26097);
nor U26750 (N_26750,N_26182,N_26145);
and U26751 (N_26751,N_25878,N_26059);
nand U26752 (N_26752,N_25836,N_26331);
and U26753 (N_26753,N_26047,N_26300);
or U26754 (N_26754,N_26004,N_26314);
or U26755 (N_26755,N_25902,N_26026);
xor U26756 (N_26756,N_26287,N_25866);
nor U26757 (N_26757,N_26338,N_26157);
xnor U26758 (N_26758,N_26399,N_25906);
xnor U26759 (N_26759,N_25877,N_26135);
xor U26760 (N_26760,N_26268,N_26363);
xnor U26761 (N_26761,N_26245,N_26171);
xor U26762 (N_26762,N_25819,N_25863);
nand U26763 (N_26763,N_26327,N_26198);
nand U26764 (N_26764,N_25840,N_26340);
or U26765 (N_26765,N_25964,N_25801);
xor U26766 (N_26766,N_26147,N_25982);
xnor U26767 (N_26767,N_25921,N_26311);
or U26768 (N_26768,N_26187,N_25917);
nor U26769 (N_26769,N_25824,N_25913);
and U26770 (N_26770,N_25849,N_26187);
or U26771 (N_26771,N_26340,N_26290);
or U26772 (N_26772,N_25903,N_26384);
nor U26773 (N_26773,N_26185,N_26368);
nor U26774 (N_26774,N_25836,N_25819);
nor U26775 (N_26775,N_26304,N_25828);
nand U26776 (N_26776,N_26348,N_26346);
nand U26777 (N_26777,N_25910,N_26013);
and U26778 (N_26778,N_25979,N_25838);
xor U26779 (N_26779,N_26125,N_25920);
nand U26780 (N_26780,N_26108,N_25960);
or U26781 (N_26781,N_26169,N_25846);
nand U26782 (N_26782,N_26004,N_26273);
nor U26783 (N_26783,N_26141,N_26233);
or U26784 (N_26784,N_25986,N_26199);
nor U26785 (N_26785,N_26156,N_25916);
xnor U26786 (N_26786,N_26197,N_26058);
or U26787 (N_26787,N_25864,N_26356);
nand U26788 (N_26788,N_25960,N_26380);
and U26789 (N_26789,N_25926,N_26054);
xnor U26790 (N_26790,N_26322,N_26080);
or U26791 (N_26791,N_25868,N_25900);
or U26792 (N_26792,N_26029,N_25924);
xnor U26793 (N_26793,N_25863,N_26061);
nor U26794 (N_26794,N_25906,N_25928);
nor U26795 (N_26795,N_26123,N_25902);
nor U26796 (N_26796,N_26094,N_26071);
nor U26797 (N_26797,N_26251,N_26310);
or U26798 (N_26798,N_25864,N_26070);
nor U26799 (N_26799,N_26027,N_26096);
nor U26800 (N_26800,N_26098,N_26306);
or U26801 (N_26801,N_26009,N_25844);
and U26802 (N_26802,N_26117,N_26325);
or U26803 (N_26803,N_26233,N_26033);
xor U26804 (N_26804,N_26038,N_26115);
or U26805 (N_26805,N_26162,N_25833);
or U26806 (N_26806,N_25944,N_26042);
xnor U26807 (N_26807,N_26053,N_25933);
or U26808 (N_26808,N_25945,N_26036);
and U26809 (N_26809,N_25942,N_25870);
nor U26810 (N_26810,N_26294,N_25959);
nand U26811 (N_26811,N_26342,N_26198);
nand U26812 (N_26812,N_26140,N_25820);
and U26813 (N_26813,N_26089,N_25945);
nor U26814 (N_26814,N_25870,N_26035);
and U26815 (N_26815,N_26107,N_25950);
nand U26816 (N_26816,N_26035,N_26223);
or U26817 (N_26817,N_26155,N_26315);
nor U26818 (N_26818,N_26019,N_26385);
nor U26819 (N_26819,N_26003,N_26050);
and U26820 (N_26820,N_25833,N_26297);
xor U26821 (N_26821,N_26311,N_26041);
nand U26822 (N_26822,N_26172,N_26191);
and U26823 (N_26823,N_26123,N_26154);
nor U26824 (N_26824,N_26344,N_25940);
nor U26825 (N_26825,N_25974,N_25887);
nand U26826 (N_26826,N_25885,N_26111);
nor U26827 (N_26827,N_25901,N_26302);
or U26828 (N_26828,N_26170,N_26224);
and U26829 (N_26829,N_26394,N_26250);
nor U26830 (N_26830,N_26157,N_26035);
or U26831 (N_26831,N_25918,N_26210);
and U26832 (N_26832,N_26275,N_26057);
and U26833 (N_26833,N_25864,N_25894);
and U26834 (N_26834,N_25959,N_26265);
or U26835 (N_26835,N_26020,N_26125);
or U26836 (N_26836,N_25860,N_25904);
or U26837 (N_26837,N_26285,N_26170);
and U26838 (N_26838,N_25903,N_25947);
nor U26839 (N_26839,N_26328,N_26045);
or U26840 (N_26840,N_26303,N_26275);
xor U26841 (N_26841,N_25957,N_25800);
nor U26842 (N_26842,N_26055,N_26116);
and U26843 (N_26843,N_26311,N_25865);
nor U26844 (N_26844,N_26240,N_26293);
xor U26845 (N_26845,N_26143,N_26118);
and U26846 (N_26846,N_26095,N_25956);
xnor U26847 (N_26847,N_26106,N_26292);
nand U26848 (N_26848,N_26222,N_25835);
and U26849 (N_26849,N_25987,N_25956);
nand U26850 (N_26850,N_25875,N_26308);
and U26851 (N_26851,N_26102,N_26227);
or U26852 (N_26852,N_26119,N_25921);
or U26853 (N_26853,N_26383,N_26163);
and U26854 (N_26854,N_26053,N_26180);
and U26855 (N_26855,N_26200,N_25982);
xnor U26856 (N_26856,N_25987,N_26248);
nand U26857 (N_26857,N_25919,N_25962);
xnor U26858 (N_26858,N_26120,N_26381);
or U26859 (N_26859,N_25807,N_26219);
nand U26860 (N_26860,N_26125,N_25873);
and U26861 (N_26861,N_25967,N_26374);
or U26862 (N_26862,N_26021,N_25803);
nor U26863 (N_26863,N_26014,N_26168);
or U26864 (N_26864,N_26025,N_26028);
nor U26865 (N_26865,N_26261,N_25889);
xnor U26866 (N_26866,N_26218,N_26035);
and U26867 (N_26867,N_25826,N_25988);
nand U26868 (N_26868,N_25879,N_26032);
xor U26869 (N_26869,N_26228,N_26396);
xnor U26870 (N_26870,N_26016,N_26394);
xor U26871 (N_26871,N_25913,N_25979);
or U26872 (N_26872,N_25838,N_26306);
or U26873 (N_26873,N_26186,N_26315);
xnor U26874 (N_26874,N_25958,N_25954);
and U26875 (N_26875,N_26092,N_25824);
xnor U26876 (N_26876,N_26234,N_26096);
and U26877 (N_26877,N_26208,N_25903);
and U26878 (N_26878,N_26257,N_26315);
and U26879 (N_26879,N_26134,N_25827);
or U26880 (N_26880,N_25879,N_26117);
or U26881 (N_26881,N_26205,N_25947);
nor U26882 (N_26882,N_25857,N_26289);
and U26883 (N_26883,N_26041,N_26389);
xnor U26884 (N_26884,N_26173,N_25822);
and U26885 (N_26885,N_25952,N_26151);
and U26886 (N_26886,N_26219,N_26107);
nand U26887 (N_26887,N_26228,N_26361);
nor U26888 (N_26888,N_25821,N_26328);
and U26889 (N_26889,N_26242,N_25817);
nor U26890 (N_26890,N_25955,N_25921);
xor U26891 (N_26891,N_26272,N_25960);
or U26892 (N_26892,N_26191,N_25943);
xor U26893 (N_26893,N_25937,N_25875);
or U26894 (N_26894,N_25916,N_26114);
and U26895 (N_26895,N_26337,N_26025);
nand U26896 (N_26896,N_26224,N_26207);
xor U26897 (N_26897,N_26166,N_26136);
xor U26898 (N_26898,N_26011,N_25955);
and U26899 (N_26899,N_26110,N_26271);
and U26900 (N_26900,N_25941,N_26274);
xnor U26901 (N_26901,N_26205,N_26042);
nor U26902 (N_26902,N_26008,N_26292);
and U26903 (N_26903,N_25893,N_25933);
nor U26904 (N_26904,N_26292,N_26254);
nand U26905 (N_26905,N_26378,N_26339);
and U26906 (N_26906,N_26165,N_26214);
nor U26907 (N_26907,N_26098,N_26007);
nand U26908 (N_26908,N_25863,N_26325);
and U26909 (N_26909,N_26160,N_25821);
xor U26910 (N_26910,N_25935,N_26394);
and U26911 (N_26911,N_26137,N_25954);
and U26912 (N_26912,N_25913,N_25919);
xor U26913 (N_26913,N_26185,N_26149);
nand U26914 (N_26914,N_26193,N_25897);
and U26915 (N_26915,N_25953,N_26350);
nand U26916 (N_26916,N_25970,N_26229);
nor U26917 (N_26917,N_26023,N_26108);
and U26918 (N_26918,N_26015,N_26038);
nand U26919 (N_26919,N_25847,N_25809);
or U26920 (N_26920,N_26044,N_26155);
xnor U26921 (N_26921,N_26273,N_26274);
or U26922 (N_26922,N_26268,N_26235);
nor U26923 (N_26923,N_26075,N_26271);
xor U26924 (N_26924,N_26313,N_26074);
nand U26925 (N_26925,N_26300,N_25855);
and U26926 (N_26926,N_26391,N_26018);
and U26927 (N_26927,N_26113,N_26130);
and U26928 (N_26928,N_25968,N_26190);
nand U26929 (N_26929,N_26156,N_26336);
and U26930 (N_26930,N_25920,N_25842);
and U26931 (N_26931,N_26057,N_25841);
xor U26932 (N_26932,N_26235,N_26282);
or U26933 (N_26933,N_26016,N_26141);
nor U26934 (N_26934,N_26190,N_25818);
or U26935 (N_26935,N_25806,N_26252);
and U26936 (N_26936,N_26289,N_25980);
or U26937 (N_26937,N_25953,N_25991);
and U26938 (N_26938,N_25890,N_25819);
and U26939 (N_26939,N_26111,N_26351);
nor U26940 (N_26940,N_26123,N_26167);
xor U26941 (N_26941,N_26221,N_26126);
nand U26942 (N_26942,N_25807,N_25814);
or U26943 (N_26943,N_25906,N_26088);
nor U26944 (N_26944,N_26079,N_25859);
nor U26945 (N_26945,N_26389,N_25888);
nand U26946 (N_26946,N_26292,N_26347);
and U26947 (N_26947,N_26375,N_26202);
or U26948 (N_26948,N_26263,N_25819);
or U26949 (N_26949,N_26392,N_25920);
nor U26950 (N_26950,N_26207,N_25976);
or U26951 (N_26951,N_26271,N_26047);
nor U26952 (N_26952,N_26020,N_25900);
and U26953 (N_26953,N_25846,N_26106);
nor U26954 (N_26954,N_26166,N_25867);
nor U26955 (N_26955,N_25924,N_26293);
and U26956 (N_26956,N_25930,N_26295);
xnor U26957 (N_26957,N_26034,N_25839);
xnor U26958 (N_26958,N_26094,N_25880);
or U26959 (N_26959,N_25967,N_26087);
or U26960 (N_26960,N_26225,N_26375);
nor U26961 (N_26961,N_25815,N_26387);
xor U26962 (N_26962,N_25997,N_25862);
and U26963 (N_26963,N_25837,N_25905);
xor U26964 (N_26964,N_26361,N_25802);
or U26965 (N_26965,N_26338,N_25801);
and U26966 (N_26966,N_26327,N_26374);
or U26967 (N_26967,N_26246,N_26051);
and U26968 (N_26968,N_25888,N_25962);
xnor U26969 (N_26969,N_25990,N_26172);
nor U26970 (N_26970,N_26000,N_26236);
or U26971 (N_26971,N_25812,N_26205);
nor U26972 (N_26972,N_26055,N_25820);
nor U26973 (N_26973,N_26367,N_26151);
and U26974 (N_26974,N_25813,N_26105);
or U26975 (N_26975,N_25877,N_25962);
and U26976 (N_26976,N_26305,N_26010);
or U26977 (N_26977,N_26285,N_26340);
nor U26978 (N_26978,N_25977,N_26070);
xor U26979 (N_26979,N_26139,N_26212);
nand U26980 (N_26980,N_25931,N_26179);
xor U26981 (N_26981,N_26311,N_26396);
xnor U26982 (N_26982,N_26183,N_25840);
or U26983 (N_26983,N_26153,N_26173);
nor U26984 (N_26984,N_26031,N_25828);
and U26985 (N_26985,N_25923,N_25869);
nor U26986 (N_26986,N_26287,N_26269);
and U26987 (N_26987,N_26199,N_26316);
nor U26988 (N_26988,N_25844,N_25802);
nor U26989 (N_26989,N_26305,N_25980);
nor U26990 (N_26990,N_26141,N_26048);
or U26991 (N_26991,N_26037,N_26207);
nor U26992 (N_26992,N_26352,N_26148);
nand U26993 (N_26993,N_26348,N_26178);
and U26994 (N_26994,N_26210,N_25993);
and U26995 (N_26995,N_26179,N_25905);
or U26996 (N_26996,N_26005,N_26248);
and U26997 (N_26997,N_26235,N_26389);
xnor U26998 (N_26998,N_25881,N_26027);
nor U26999 (N_26999,N_26132,N_26021);
nand U27000 (N_27000,N_26786,N_26754);
or U27001 (N_27001,N_26416,N_26675);
and U27002 (N_27002,N_26809,N_26855);
and U27003 (N_27003,N_26716,N_26918);
xnor U27004 (N_27004,N_26775,N_26839);
xnor U27005 (N_27005,N_26993,N_26963);
nor U27006 (N_27006,N_26653,N_26593);
and U27007 (N_27007,N_26686,N_26605);
xnor U27008 (N_27008,N_26457,N_26475);
and U27009 (N_27009,N_26897,N_26769);
nand U27010 (N_27010,N_26739,N_26537);
xor U27011 (N_27011,N_26538,N_26471);
xor U27012 (N_27012,N_26922,N_26917);
nor U27013 (N_27013,N_26735,N_26817);
nand U27014 (N_27014,N_26934,N_26900);
nand U27015 (N_27015,N_26893,N_26927);
xnor U27016 (N_27016,N_26911,N_26752);
or U27017 (N_27017,N_26969,N_26847);
or U27018 (N_27018,N_26550,N_26854);
and U27019 (N_27019,N_26522,N_26955);
nand U27020 (N_27020,N_26808,N_26743);
or U27021 (N_27021,N_26683,N_26936);
nand U27022 (N_27022,N_26999,N_26602);
nor U27023 (N_27023,N_26821,N_26564);
and U27024 (N_27024,N_26878,N_26852);
nand U27025 (N_27025,N_26598,N_26534);
xor U27026 (N_27026,N_26453,N_26723);
and U27027 (N_27027,N_26884,N_26826);
nand U27028 (N_27028,N_26626,N_26915);
nor U27029 (N_27029,N_26780,N_26555);
nand U27030 (N_27030,N_26532,N_26456);
and U27031 (N_27031,N_26460,N_26757);
nand U27032 (N_27032,N_26882,N_26539);
xor U27033 (N_27033,N_26742,N_26877);
nand U27034 (N_27034,N_26549,N_26766);
xnor U27035 (N_27035,N_26488,N_26570);
nand U27036 (N_27036,N_26436,N_26748);
or U27037 (N_27037,N_26482,N_26493);
xor U27038 (N_27038,N_26941,N_26853);
and U27039 (N_27039,N_26466,N_26709);
and U27040 (N_27040,N_26793,N_26873);
nor U27041 (N_27041,N_26740,N_26584);
nand U27042 (N_27042,N_26650,N_26422);
xor U27043 (N_27043,N_26664,N_26872);
nand U27044 (N_27044,N_26901,N_26556);
nor U27045 (N_27045,N_26458,N_26518);
and U27046 (N_27046,N_26846,N_26880);
xor U27047 (N_27047,N_26985,N_26656);
and U27048 (N_27048,N_26601,N_26498);
or U27049 (N_27049,N_26960,N_26486);
and U27050 (N_27050,N_26797,N_26816);
or U27051 (N_27051,N_26926,N_26618);
nand U27052 (N_27052,N_26856,N_26685);
xor U27053 (N_27053,N_26542,N_26505);
nand U27054 (N_27054,N_26541,N_26851);
and U27055 (N_27055,N_26508,N_26724);
nand U27056 (N_27056,N_26659,N_26992);
xor U27057 (N_27057,N_26545,N_26703);
xnor U27058 (N_27058,N_26421,N_26528);
xor U27059 (N_27059,N_26613,N_26527);
nor U27060 (N_27060,N_26708,N_26758);
nand U27061 (N_27061,N_26502,N_26595);
nand U27062 (N_27062,N_26417,N_26753);
nor U27063 (N_27063,N_26699,N_26414);
or U27064 (N_27064,N_26449,N_26863);
or U27065 (N_27065,N_26660,N_26712);
nand U27066 (N_27066,N_26507,N_26599);
nor U27067 (N_27067,N_26476,N_26516);
or U27068 (N_27068,N_26696,N_26459);
nor U27069 (N_27069,N_26432,N_26828);
or U27070 (N_27070,N_26731,N_26710);
or U27071 (N_27071,N_26480,N_26760);
or U27072 (N_27072,N_26940,N_26672);
and U27073 (N_27073,N_26904,N_26619);
xnor U27074 (N_27074,N_26481,N_26563);
nor U27075 (N_27075,N_26446,N_26485);
or U27076 (N_27076,N_26947,N_26778);
nand U27077 (N_27077,N_26407,N_26818);
nand U27078 (N_27078,N_26573,N_26634);
nor U27079 (N_27079,N_26764,N_26939);
nor U27080 (N_27080,N_26666,N_26409);
and U27081 (N_27081,N_26833,N_26945);
nand U27082 (N_27082,N_26574,N_26806);
nand U27083 (N_27083,N_26881,N_26772);
nand U27084 (N_27084,N_26864,N_26657);
or U27085 (N_27085,N_26491,N_26495);
or U27086 (N_27086,N_26937,N_26623);
and U27087 (N_27087,N_26500,N_26569);
and U27088 (N_27088,N_26938,N_26535);
xor U27089 (N_27089,N_26596,N_26559);
xor U27090 (N_27090,N_26720,N_26694);
or U27091 (N_27091,N_26981,N_26603);
or U27092 (N_27092,N_26916,N_26718);
xnor U27093 (N_27093,N_26787,N_26943);
nand U27094 (N_27094,N_26803,N_26636);
nor U27095 (N_27095,N_26651,N_26698);
and U27096 (N_27096,N_26933,N_26445);
or U27097 (N_27097,N_26568,N_26942);
xnor U27098 (N_27098,N_26631,N_26746);
xnor U27099 (N_27099,N_26438,N_26715);
and U27100 (N_27100,N_26580,N_26565);
xnor U27101 (N_27101,N_26761,N_26474);
nor U27102 (N_27102,N_26519,N_26649);
nor U27103 (N_27103,N_26827,N_26661);
nor U27104 (N_27104,N_26845,N_26857);
nand U27105 (N_27105,N_26707,N_26713);
xor U27106 (N_27106,N_26467,N_26891);
xnor U27107 (N_27107,N_26865,N_26702);
xnor U27108 (N_27108,N_26967,N_26452);
nand U27109 (N_27109,N_26540,N_26734);
xor U27110 (N_27110,N_26774,N_26907);
and U27111 (N_27111,N_26807,N_26455);
and U27112 (N_27112,N_26905,N_26406);
or U27113 (N_27113,N_26597,N_26487);
nor U27114 (N_27114,N_26795,N_26948);
nand U27115 (N_27115,N_26861,N_26990);
or U27116 (N_27116,N_26987,N_26577);
xor U27117 (N_27117,N_26517,N_26871);
nand U27118 (N_27118,N_26469,N_26444);
or U27119 (N_27119,N_26984,N_26697);
nor U27120 (N_27120,N_26420,N_26544);
nand U27121 (N_27121,N_26658,N_26970);
xor U27122 (N_27122,N_26405,N_26621);
nand U27123 (N_27123,N_26705,N_26430);
nor U27124 (N_27124,N_26768,N_26737);
and U27125 (N_27125,N_26701,N_26957);
and U27126 (N_27126,N_26804,N_26511);
or U27127 (N_27127,N_26607,N_26567);
xnor U27128 (N_27128,N_26441,N_26501);
nand U27129 (N_27129,N_26678,N_26779);
xor U27130 (N_27130,N_26831,N_26503);
nor U27131 (N_27131,N_26971,N_26426);
or U27132 (N_27132,N_26763,N_26874);
nand U27133 (N_27133,N_26526,N_26546);
nand U27134 (N_27134,N_26810,N_26935);
and U27135 (N_27135,N_26591,N_26682);
nor U27136 (N_27136,N_26552,N_26730);
xnor U27137 (N_27137,N_26662,N_26729);
xnor U27138 (N_27138,N_26886,N_26914);
nor U27139 (N_27139,N_26468,N_26642);
nor U27140 (N_27140,N_26510,N_26732);
or U27141 (N_27141,N_26627,N_26980);
or U27142 (N_27142,N_26465,N_26755);
nand U27143 (N_27143,N_26801,N_26860);
and U27144 (N_27144,N_26814,N_26403);
nor U27145 (N_27145,N_26972,N_26654);
and U27146 (N_27146,N_26749,N_26944);
nand U27147 (N_27147,N_26473,N_26687);
nor U27148 (N_27148,N_26461,N_26840);
or U27149 (N_27149,N_26625,N_26923);
nor U27150 (N_27150,N_26677,N_26805);
and U27151 (N_27151,N_26974,N_26684);
and U27152 (N_27152,N_26490,N_26896);
nor U27153 (N_27153,N_26913,N_26431);
and U27154 (N_27154,N_26428,N_26885);
xor U27155 (N_27155,N_26830,N_26448);
nor U27156 (N_27156,N_26747,N_26609);
nor U27157 (N_27157,N_26998,N_26796);
or U27158 (N_27158,N_26585,N_26859);
nor U27159 (N_27159,N_26433,N_26910);
xnor U27160 (N_27160,N_26496,N_26524);
xor U27161 (N_27161,N_26437,N_26930);
or U27162 (N_27162,N_26892,N_26557);
nor U27163 (N_27163,N_26566,N_26628);
and U27164 (N_27164,N_26722,N_26714);
xor U27165 (N_27165,N_26733,N_26695);
nor U27166 (N_27166,N_26690,N_26889);
nor U27167 (N_27167,N_26615,N_26590);
xnor U27168 (N_27168,N_26640,N_26838);
nand U27169 (N_27169,N_26425,N_26866);
nand U27170 (N_27170,N_26842,N_26652);
and U27171 (N_27171,N_26727,N_26523);
nand U27172 (N_27172,N_26671,N_26767);
or U27173 (N_27173,N_26515,N_26946);
and U27174 (N_27174,N_26783,N_26589);
nor U27175 (N_27175,N_26921,N_26909);
nor U27176 (N_27176,N_26961,N_26711);
or U27177 (N_27177,N_26858,N_26400);
and U27178 (N_27178,N_26844,N_26558);
nor U27179 (N_27179,N_26875,N_26560);
or U27180 (N_27180,N_26782,N_26899);
nor U27181 (N_27181,N_26908,N_26588);
xnor U27182 (N_27182,N_26484,N_26792);
nand U27183 (N_27183,N_26439,N_26647);
xor U27184 (N_27184,N_26463,N_26781);
and U27185 (N_27185,N_26949,N_26529);
or U27186 (N_27186,N_26520,N_26610);
xnor U27187 (N_27187,N_26410,N_26953);
or U27188 (N_27188,N_26788,N_26408);
and U27189 (N_27189,N_26464,N_26401);
nor U27190 (N_27190,N_26419,N_26995);
nand U27191 (N_27191,N_26415,N_26632);
nor U27192 (N_27192,N_26835,N_26789);
or U27193 (N_27193,N_26543,N_26614);
or U27194 (N_27194,N_26841,N_26587);
nand U27195 (N_27195,N_26888,N_26950);
nand U27196 (N_27196,N_26721,N_26429);
and U27197 (N_27197,N_26620,N_26962);
nand U27198 (N_27198,N_26513,N_26834);
nor U27199 (N_27199,N_26777,N_26454);
or U27200 (N_27200,N_26867,N_26669);
nor U27201 (N_27201,N_26771,N_26876);
xnor U27202 (N_27202,N_26784,N_26622);
nand U27203 (N_27203,N_26726,N_26820);
nand U27204 (N_27204,N_26676,N_26443);
nand U27205 (N_27205,N_26679,N_26616);
and U27206 (N_27206,N_26706,N_26689);
or U27207 (N_27207,N_26756,N_26478);
nor U27208 (N_27208,N_26988,N_26423);
nand U27209 (N_27209,N_26979,N_26612);
and U27210 (N_27210,N_26802,N_26402);
nand U27211 (N_27211,N_26837,N_26608);
xnor U27212 (N_27212,N_26906,N_26581);
xnor U27213 (N_27213,N_26725,N_26521);
and U27214 (N_27214,N_26499,N_26509);
or U27215 (N_27215,N_26750,N_26819);
nor U27216 (N_27216,N_26954,N_26968);
and U27217 (N_27217,N_26579,N_26667);
nor U27218 (N_27218,N_26850,N_26773);
or U27219 (N_27219,N_26604,N_26643);
nor U27220 (N_27220,N_26790,N_26572);
or U27221 (N_27221,N_26673,N_26890);
nor U27222 (N_27222,N_26424,N_26479);
or U27223 (N_27223,N_26870,N_26794);
and U27224 (N_27224,N_26575,N_26829);
xnor U27225 (N_27225,N_26964,N_26849);
nor U27226 (N_27226,N_26770,N_26606);
nand U27227 (N_27227,N_26418,N_26655);
nand U27228 (N_27228,N_26751,N_26929);
nand U27229 (N_27229,N_26822,N_26670);
nor U27230 (N_27230,N_26548,N_26447);
xnor U27231 (N_27231,N_26586,N_26629);
nor U27232 (N_27232,N_26412,N_26951);
and U27233 (N_27233,N_26648,N_26561);
and U27234 (N_27234,N_26531,N_26932);
and U27235 (N_27235,N_26411,N_26959);
and U27236 (N_27236,N_26435,N_26958);
nand U27237 (N_27237,N_26646,N_26427);
xnor U27238 (N_27238,N_26492,N_26404);
and U27239 (N_27239,N_26977,N_26719);
nor U27240 (N_27240,N_26728,N_26641);
nor U27241 (N_27241,N_26530,N_26989);
or U27242 (N_27242,N_26952,N_26639);
or U27243 (N_27243,N_26688,N_26894);
xnor U27244 (N_27244,N_26451,N_26553);
or U27245 (N_27245,N_26920,N_26887);
nor U27246 (N_27246,N_26738,N_26832);
or U27247 (N_27247,N_26978,N_26895);
nand U27248 (N_27248,N_26630,N_26592);
nor U27249 (N_27249,N_26848,N_26879);
nand U27250 (N_27250,N_26966,N_26462);
or U27251 (N_27251,N_26681,N_26497);
xnor U27252 (N_27252,N_26434,N_26996);
and U27253 (N_27253,N_26843,N_26925);
xnor U27254 (N_27254,N_26717,N_26862);
nor U27255 (N_27255,N_26973,N_26692);
xor U27256 (N_27256,N_26975,N_26825);
nor U27257 (N_27257,N_26815,N_26997);
nand U27258 (N_27258,N_26504,N_26869);
nor U27259 (N_27259,N_26562,N_26413);
nor U27260 (N_27260,N_26536,N_26547);
xnor U27261 (N_27261,N_26551,N_26635);
or U27262 (N_27262,N_26798,N_26442);
or U27263 (N_27263,N_26440,N_26624);
nand U27264 (N_27264,N_26594,N_26644);
and U27265 (N_27265,N_26665,N_26483);
nand U27266 (N_27266,N_26762,N_26898);
and U27267 (N_27267,N_26868,N_26883);
xor U27268 (N_27268,N_26617,N_26533);
and U27269 (N_27269,N_26986,N_26903);
and U27270 (N_27270,N_26489,N_26776);
and U27271 (N_27271,N_26704,N_26811);
xnor U27272 (N_27272,N_26700,N_26812);
xor U27273 (N_27273,N_26791,N_26741);
or U27274 (N_27274,N_26924,N_26674);
and U27275 (N_27275,N_26668,N_26450);
xnor U27276 (N_27276,N_26680,N_26823);
xnor U27277 (N_27277,N_26836,N_26745);
xor U27278 (N_27278,N_26799,N_26512);
nand U27279 (N_27279,N_26965,N_26514);
xnor U27280 (N_27280,N_26824,N_26611);
xor U27281 (N_27281,N_26813,N_26638);
or U27282 (N_27282,N_26800,N_26902);
nor U27283 (N_27283,N_26956,N_26765);
nor U27284 (N_27284,N_26494,N_26576);
and U27285 (N_27285,N_26571,N_26982);
nor U27286 (N_27286,N_26633,N_26983);
nand U27287 (N_27287,N_26637,N_26994);
and U27288 (N_27288,N_26600,N_26744);
xor U27289 (N_27289,N_26578,N_26554);
nand U27290 (N_27290,N_26583,N_26693);
and U27291 (N_27291,N_26976,N_26477);
nor U27292 (N_27292,N_26785,N_26691);
and U27293 (N_27293,N_26919,N_26470);
nor U27294 (N_27294,N_26582,N_26506);
and U27295 (N_27295,N_26928,N_26931);
nand U27296 (N_27296,N_26991,N_26472);
or U27297 (N_27297,N_26759,N_26912);
or U27298 (N_27298,N_26663,N_26525);
or U27299 (N_27299,N_26736,N_26645);
and U27300 (N_27300,N_26656,N_26607);
nand U27301 (N_27301,N_26641,N_26674);
or U27302 (N_27302,N_26880,N_26596);
nand U27303 (N_27303,N_26957,N_26411);
xnor U27304 (N_27304,N_26830,N_26532);
nor U27305 (N_27305,N_26960,N_26434);
or U27306 (N_27306,N_26594,N_26851);
xor U27307 (N_27307,N_26424,N_26665);
or U27308 (N_27308,N_26953,N_26848);
nand U27309 (N_27309,N_26729,N_26974);
nor U27310 (N_27310,N_26951,N_26833);
nor U27311 (N_27311,N_26934,N_26879);
and U27312 (N_27312,N_26554,N_26820);
nand U27313 (N_27313,N_26523,N_26903);
nand U27314 (N_27314,N_26950,N_26796);
xnor U27315 (N_27315,N_26429,N_26882);
nor U27316 (N_27316,N_26505,N_26418);
xnor U27317 (N_27317,N_26907,N_26867);
or U27318 (N_27318,N_26436,N_26609);
or U27319 (N_27319,N_26696,N_26643);
nand U27320 (N_27320,N_26542,N_26965);
and U27321 (N_27321,N_26523,N_26886);
or U27322 (N_27322,N_26797,N_26579);
nand U27323 (N_27323,N_26827,N_26496);
xnor U27324 (N_27324,N_26577,N_26957);
and U27325 (N_27325,N_26568,N_26762);
xnor U27326 (N_27326,N_26837,N_26610);
xnor U27327 (N_27327,N_26947,N_26600);
or U27328 (N_27328,N_26489,N_26841);
nor U27329 (N_27329,N_26720,N_26979);
nand U27330 (N_27330,N_26559,N_26969);
nand U27331 (N_27331,N_26511,N_26510);
and U27332 (N_27332,N_26494,N_26552);
nor U27333 (N_27333,N_26469,N_26594);
nand U27334 (N_27334,N_26645,N_26852);
and U27335 (N_27335,N_26762,N_26818);
or U27336 (N_27336,N_26420,N_26749);
nor U27337 (N_27337,N_26998,N_26890);
nand U27338 (N_27338,N_26432,N_26727);
nand U27339 (N_27339,N_26642,N_26910);
nand U27340 (N_27340,N_26891,N_26541);
nor U27341 (N_27341,N_26915,N_26969);
and U27342 (N_27342,N_26516,N_26623);
nand U27343 (N_27343,N_26571,N_26751);
or U27344 (N_27344,N_26597,N_26400);
nor U27345 (N_27345,N_26729,N_26726);
and U27346 (N_27346,N_26885,N_26730);
nand U27347 (N_27347,N_26567,N_26722);
xor U27348 (N_27348,N_26992,N_26643);
xor U27349 (N_27349,N_26524,N_26577);
and U27350 (N_27350,N_26877,N_26840);
xor U27351 (N_27351,N_26841,N_26452);
nand U27352 (N_27352,N_26513,N_26540);
xor U27353 (N_27353,N_26789,N_26462);
nand U27354 (N_27354,N_26810,N_26532);
nor U27355 (N_27355,N_26455,N_26613);
nor U27356 (N_27356,N_26926,N_26850);
and U27357 (N_27357,N_26529,N_26824);
nand U27358 (N_27358,N_26770,N_26956);
or U27359 (N_27359,N_26581,N_26627);
and U27360 (N_27360,N_26595,N_26873);
or U27361 (N_27361,N_26556,N_26559);
or U27362 (N_27362,N_26425,N_26864);
nor U27363 (N_27363,N_26474,N_26682);
xor U27364 (N_27364,N_26432,N_26895);
and U27365 (N_27365,N_26506,N_26700);
or U27366 (N_27366,N_26970,N_26488);
and U27367 (N_27367,N_26405,N_26731);
and U27368 (N_27368,N_26986,N_26961);
nor U27369 (N_27369,N_26769,N_26645);
or U27370 (N_27370,N_26976,N_26730);
nand U27371 (N_27371,N_26626,N_26610);
xor U27372 (N_27372,N_26771,N_26521);
or U27373 (N_27373,N_26635,N_26982);
or U27374 (N_27374,N_26464,N_26676);
nand U27375 (N_27375,N_26810,N_26977);
xnor U27376 (N_27376,N_26838,N_26624);
xor U27377 (N_27377,N_26888,N_26481);
xnor U27378 (N_27378,N_26955,N_26548);
and U27379 (N_27379,N_26733,N_26829);
and U27380 (N_27380,N_26798,N_26522);
xor U27381 (N_27381,N_26813,N_26825);
or U27382 (N_27382,N_26516,N_26706);
or U27383 (N_27383,N_26920,N_26416);
nand U27384 (N_27384,N_26912,N_26747);
nor U27385 (N_27385,N_26504,N_26664);
nor U27386 (N_27386,N_26506,N_26754);
nand U27387 (N_27387,N_26576,N_26870);
nand U27388 (N_27388,N_26538,N_26621);
and U27389 (N_27389,N_26569,N_26571);
xnor U27390 (N_27390,N_26648,N_26604);
and U27391 (N_27391,N_26672,N_26774);
or U27392 (N_27392,N_26776,N_26805);
or U27393 (N_27393,N_26656,N_26707);
and U27394 (N_27394,N_26650,N_26870);
nor U27395 (N_27395,N_26919,N_26986);
and U27396 (N_27396,N_26627,N_26851);
nand U27397 (N_27397,N_26976,N_26481);
and U27398 (N_27398,N_26798,N_26803);
nor U27399 (N_27399,N_26506,N_26697);
nand U27400 (N_27400,N_26932,N_26586);
nand U27401 (N_27401,N_26537,N_26407);
or U27402 (N_27402,N_26673,N_26601);
nor U27403 (N_27403,N_26543,N_26836);
xnor U27404 (N_27404,N_26412,N_26997);
nor U27405 (N_27405,N_26802,N_26949);
or U27406 (N_27406,N_26566,N_26696);
and U27407 (N_27407,N_26404,N_26777);
nor U27408 (N_27408,N_26852,N_26922);
and U27409 (N_27409,N_26627,N_26696);
and U27410 (N_27410,N_26791,N_26712);
xor U27411 (N_27411,N_26650,N_26575);
nand U27412 (N_27412,N_26581,N_26576);
or U27413 (N_27413,N_26959,N_26710);
nand U27414 (N_27414,N_26833,N_26500);
nor U27415 (N_27415,N_26724,N_26438);
nor U27416 (N_27416,N_26743,N_26653);
and U27417 (N_27417,N_26628,N_26511);
xnor U27418 (N_27418,N_26414,N_26910);
nand U27419 (N_27419,N_26585,N_26584);
and U27420 (N_27420,N_26424,N_26439);
nor U27421 (N_27421,N_26698,N_26709);
nor U27422 (N_27422,N_26623,N_26786);
xnor U27423 (N_27423,N_26876,N_26984);
and U27424 (N_27424,N_26912,N_26562);
xor U27425 (N_27425,N_26862,N_26914);
nand U27426 (N_27426,N_26536,N_26962);
nor U27427 (N_27427,N_26814,N_26561);
and U27428 (N_27428,N_26952,N_26922);
or U27429 (N_27429,N_26555,N_26947);
nor U27430 (N_27430,N_26506,N_26402);
xnor U27431 (N_27431,N_26908,N_26953);
nand U27432 (N_27432,N_26997,N_26497);
and U27433 (N_27433,N_26672,N_26629);
nand U27434 (N_27434,N_26561,N_26741);
and U27435 (N_27435,N_26734,N_26747);
or U27436 (N_27436,N_26943,N_26703);
or U27437 (N_27437,N_26541,N_26896);
nor U27438 (N_27438,N_26926,N_26486);
nand U27439 (N_27439,N_26944,N_26820);
nor U27440 (N_27440,N_26648,N_26922);
and U27441 (N_27441,N_26608,N_26605);
nor U27442 (N_27442,N_26871,N_26590);
and U27443 (N_27443,N_26702,N_26569);
nor U27444 (N_27444,N_26656,N_26445);
and U27445 (N_27445,N_26887,N_26703);
and U27446 (N_27446,N_26716,N_26890);
nor U27447 (N_27447,N_26703,N_26714);
nor U27448 (N_27448,N_26630,N_26595);
and U27449 (N_27449,N_26525,N_26424);
nor U27450 (N_27450,N_26675,N_26422);
nand U27451 (N_27451,N_26408,N_26726);
xor U27452 (N_27452,N_26749,N_26720);
or U27453 (N_27453,N_26705,N_26804);
and U27454 (N_27454,N_26826,N_26653);
and U27455 (N_27455,N_26958,N_26918);
or U27456 (N_27456,N_26557,N_26847);
or U27457 (N_27457,N_26573,N_26884);
and U27458 (N_27458,N_26629,N_26929);
and U27459 (N_27459,N_26686,N_26620);
xnor U27460 (N_27460,N_26587,N_26838);
xor U27461 (N_27461,N_26404,N_26718);
nand U27462 (N_27462,N_26729,N_26562);
and U27463 (N_27463,N_26605,N_26634);
and U27464 (N_27464,N_26401,N_26930);
nand U27465 (N_27465,N_26895,N_26666);
and U27466 (N_27466,N_26824,N_26699);
or U27467 (N_27467,N_26813,N_26618);
nand U27468 (N_27468,N_26410,N_26813);
xnor U27469 (N_27469,N_26447,N_26589);
nor U27470 (N_27470,N_26929,N_26774);
or U27471 (N_27471,N_26721,N_26586);
and U27472 (N_27472,N_26583,N_26868);
xnor U27473 (N_27473,N_26948,N_26542);
nand U27474 (N_27474,N_26609,N_26921);
xnor U27475 (N_27475,N_26495,N_26786);
xnor U27476 (N_27476,N_26521,N_26537);
nand U27477 (N_27477,N_26593,N_26704);
or U27478 (N_27478,N_26556,N_26758);
or U27479 (N_27479,N_26479,N_26730);
nor U27480 (N_27480,N_26865,N_26610);
or U27481 (N_27481,N_26869,N_26428);
xor U27482 (N_27482,N_26848,N_26512);
xnor U27483 (N_27483,N_26999,N_26828);
or U27484 (N_27484,N_26767,N_26829);
or U27485 (N_27485,N_26506,N_26984);
nand U27486 (N_27486,N_26880,N_26657);
or U27487 (N_27487,N_26511,N_26649);
and U27488 (N_27488,N_26774,N_26597);
and U27489 (N_27489,N_26994,N_26550);
nor U27490 (N_27490,N_26645,N_26600);
and U27491 (N_27491,N_26887,N_26491);
nor U27492 (N_27492,N_26776,N_26539);
xor U27493 (N_27493,N_26609,N_26716);
or U27494 (N_27494,N_26537,N_26621);
and U27495 (N_27495,N_26532,N_26841);
or U27496 (N_27496,N_26736,N_26573);
xor U27497 (N_27497,N_26837,N_26753);
and U27498 (N_27498,N_26763,N_26978);
xnor U27499 (N_27499,N_26943,N_26637);
nor U27500 (N_27500,N_26429,N_26991);
or U27501 (N_27501,N_26638,N_26511);
or U27502 (N_27502,N_26945,N_26598);
nor U27503 (N_27503,N_26493,N_26835);
xor U27504 (N_27504,N_26550,N_26873);
nor U27505 (N_27505,N_26623,N_26983);
xor U27506 (N_27506,N_26967,N_26617);
and U27507 (N_27507,N_26764,N_26590);
xor U27508 (N_27508,N_26618,N_26410);
and U27509 (N_27509,N_26573,N_26458);
or U27510 (N_27510,N_26674,N_26748);
xnor U27511 (N_27511,N_26970,N_26961);
and U27512 (N_27512,N_26632,N_26970);
or U27513 (N_27513,N_26507,N_26944);
or U27514 (N_27514,N_26605,N_26457);
nand U27515 (N_27515,N_26748,N_26586);
nor U27516 (N_27516,N_26827,N_26797);
or U27517 (N_27517,N_26948,N_26477);
nor U27518 (N_27518,N_26911,N_26429);
or U27519 (N_27519,N_26585,N_26519);
nand U27520 (N_27520,N_26635,N_26607);
nand U27521 (N_27521,N_26428,N_26834);
nor U27522 (N_27522,N_26764,N_26736);
xor U27523 (N_27523,N_26813,N_26698);
and U27524 (N_27524,N_26525,N_26511);
or U27525 (N_27525,N_26583,N_26422);
and U27526 (N_27526,N_26775,N_26711);
xnor U27527 (N_27527,N_26731,N_26451);
xor U27528 (N_27528,N_26806,N_26632);
or U27529 (N_27529,N_26690,N_26628);
or U27530 (N_27530,N_26946,N_26442);
xnor U27531 (N_27531,N_26528,N_26747);
nor U27532 (N_27532,N_26567,N_26773);
xnor U27533 (N_27533,N_26621,N_26743);
xor U27534 (N_27534,N_26988,N_26404);
or U27535 (N_27535,N_26838,N_26823);
nor U27536 (N_27536,N_26508,N_26598);
or U27537 (N_27537,N_26751,N_26642);
or U27538 (N_27538,N_26874,N_26925);
xnor U27539 (N_27539,N_26873,N_26927);
nand U27540 (N_27540,N_26909,N_26512);
nor U27541 (N_27541,N_26578,N_26920);
xnor U27542 (N_27542,N_26418,N_26756);
nand U27543 (N_27543,N_26479,N_26565);
xnor U27544 (N_27544,N_26975,N_26778);
nand U27545 (N_27545,N_26625,N_26797);
and U27546 (N_27546,N_26557,N_26887);
and U27547 (N_27547,N_26588,N_26735);
and U27548 (N_27548,N_26871,N_26698);
nand U27549 (N_27549,N_26670,N_26789);
xnor U27550 (N_27550,N_26650,N_26531);
nor U27551 (N_27551,N_26502,N_26443);
nand U27552 (N_27552,N_26577,N_26560);
nor U27553 (N_27553,N_26924,N_26902);
xor U27554 (N_27554,N_26417,N_26446);
xor U27555 (N_27555,N_26601,N_26492);
or U27556 (N_27556,N_26852,N_26687);
and U27557 (N_27557,N_26568,N_26991);
nor U27558 (N_27558,N_26720,N_26952);
nor U27559 (N_27559,N_26473,N_26800);
nand U27560 (N_27560,N_26870,N_26598);
and U27561 (N_27561,N_26572,N_26543);
and U27562 (N_27562,N_26507,N_26461);
xor U27563 (N_27563,N_26742,N_26941);
and U27564 (N_27564,N_26896,N_26682);
and U27565 (N_27565,N_26422,N_26817);
nor U27566 (N_27566,N_26424,N_26815);
xnor U27567 (N_27567,N_26665,N_26421);
nor U27568 (N_27568,N_26629,N_26420);
or U27569 (N_27569,N_26854,N_26934);
nand U27570 (N_27570,N_26552,N_26682);
and U27571 (N_27571,N_26963,N_26840);
or U27572 (N_27572,N_26483,N_26584);
and U27573 (N_27573,N_26650,N_26884);
xor U27574 (N_27574,N_26841,N_26842);
nand U27575 (N_27575,N_26737,N_26918);
xnor U27576 (N_27576,N_26562,N_26502);
xnor U27577 (N_27577,N_26638,N_26948);
nand U27578 (N_27578,N_26485,N_26472);
xor U27579 (N_27579,N_26805,N_26828);
xor U27580 (N_27580,N_26769,N_26753);
nor U27581 (N_27581,N_26780,N_26471);
or U27582 (N_27582,N_26665,N_26609);
nor U27583 (N_27583,N_26822,N_26422);
nand U27584 (N_27584,N_26976,N_26638);
nand U27585 (N_27585,N_26893,N_26515);
xor U27586 (N_27586,N_26746,N_26899);
nand U27587 (N_27587,N_26995,N_26647);
and U27588 (N_27588,N_26635,N_26586);
and U27589 (N_27589,N_26775,N_26621);
and U27590 (N_27590,N_26751,N_26821);
or U27591 (N_27591,N_26754,N_26966);
nand U27592 (N_27592,N_26984,N_26459);
nor U27593 (N_27593,N_26552,N_26847);
nor U27594 (N_27594,N_26554,N_26894);
and U27595 (N_27595,N_26779,N_26806);
nor U27596 (N_27596,N_26722,N_26896);
xor U27597 (N_27597,N_26598,N_26691);
nor U27598 (N_27598,N_26474,N_26478);
and U27599 (N_27599,N_26880,N_26701);
and U27600 (N_27600,N_27499,N_27388);
xnor U27601 (N_27601,N_27469,N_27332);
and U27602 (N_27602,N_27501,N_27472);
or U27603 (N_27603,N_27155,N_27431);
or U27604 (N_27604,N_27416,N_27081);
xnor U27605 (N_27605,N_27485,N_27230);
nor U27606 (N_27606,N_27584,N_27364);
and U27607 (N_27607,N_27234,N_27170);
and U27608 (N_27608,N_27118,N_27504);
nand U27609 (N_27609,N_27454,N_27082);
xnor U27610 (N_27610,N_27362,N_27140);
nand U27611 (N_27611,N_27309,N_27196);
nor U27612 (N_27612,N_27453,N_27080);
and U27613 (N_27613,N_27411,N_27449);
xnor U27614 (N_27614,N_27069,N_27053);
or U27615 (N_27615,N_27523,N_27237);
and U27616 (N_27616,N_27206,N_27199);
xor U27617 (N_27617,N_27022,N_27011);
and U27618 (N_27618,N_27437,N_27542);
nand U27619 (N_27619,N_27361,N_27208);
and U27620 (N_27620,N_27113,N_27027);
xor U27621 (N_27621,N_27198,N_27597);
and U27622 (N_27622,N_27083,N_27566);
or U27623 (N_27623,N_27127,N_27514);
xor U27624 (N_27624,N_27316,N_27333);
xor U27625 (N_27625,N_27079,N_27164);
and U27626 (N_27626,N_27508,N_27233);
nand U27627 (N_27627,N_27572,N_27112);
nor U27628 (N_27628,N_27176,N_27313);
and U27629 (N_27629,N_27355,N_27008);
or U27630 (N_27630,N_27009,N_27246);
nand U27631 (N_27631,N_27518,N_27178);
nor U27632 (N_27632,N_27274,N_27447);
xor U27633 (N_27633,N_27488,N_27038);
and U27634 (N_27634,N_27184,N_27486);
or U27635 (N_27635,N_27301,N_27075);
or U27636 (N_27636,N_27271,N_27497);
nand U27637 (N_27637,N_27205,N_27281);
nand U27638 (N_27638,N_27494,N_27458);
nor U27639 (N_27639,N_27489,N_27231);
and U27640 (N_27640,N_27573,N_27434);
and U27641 (N_27641,N_27399,N_27585);
xor U27642 (N_27642,N_27255,N_27269);
nand U27643 (N_27643,N_27282,N_27369);
xnor U27644 (N_27644,N_27560,N_27293);
or U27645 (N_27645,N_27496,N_27010);
nand U27646 (N_27646,N_27438,N_27120);
nand U27647 (N_27647,N_27302,N_27219);
or U27648 (N_27648,N_27180,N_27330);
xnor U27649 (N_27649,N_27517,N_27142);
nand U27650 (N_27650,N_27122,N_27145);
nor U27651 (N_27651,N_27159,N_27479);
xor U27652 (N_27652,N_27070,N_27457);
and U27653 (N_27653,N_27529,N_27522);
nand U27654 (N_27654,N_27032,N_27419);
xor U27655 (N_27655,N_27322,N_27304);
nor U27656 (N_27656,N_27390,N_27539);
and U27657 (N_27657,N_27280,N_27352);
and U27658 (N_27658,N_27202,N_27135);
nor U27659 (N_27659,N_27534,N_27561);
and U27660 (N_27660,N_27295,N_27284);
and U27661 (N_27661,N_27288,N_27065);
and U27662 (N_27662,N_27014,N_27250);
nor U27663 (N_27663,N_27287,N_27100);
nor U27664 (N_27664,N_27341,N_27446);
and U27665 (N_27665,N_27130,N_27144);
or U27666 (N_27666,N_27181,N_27161);
nor U27667 (N_27667,N_27521,N_27049);
or U27668 (N_27668,N_27063,N_27487);
and U27669 (N_27669,N_27136,N_27448);
nor U27670 (N_27670,N_27252,N_27039);
xor U27671 (N_27671,N_27041,N_27592);
xnor U27672 (N_27672,N_27156,N_27051);
and U27673 (N_27673,N_27154,N_27263);
nor U27674 (N_27674,N_27096,N_27241);
nor U27675 (N_27675,N_27299,N_27591);
or U27676 (N_27676,N_27466,N_27347);
xor U27677 (N_27677,N_27109,N_27267);
nor U27678 (N_27678,N_27456,N_27172);
nor U27679 (N_27679,N_27297,N_27318);
nor U27680 (N_27680,N_27290,N_27021);
nor U27681 (N_27681,N_27405,N_27005);
and U27682 (N_27682,N_27503,N_27509);
nor U27683 (N_27683,N_27106,N_27013);
nand U27684 (N_27684,N_27210,N_27110);
nand U27685 (N_27685,N_27450,N_27580);
or U27686 (N_27686,N_27427,N_27244);
nor U27687 (N_27687,N_27356,N_27593);
and U27688 (N_27688,N_27387,N_27305);
nor U27689 (N_27689,N_27569,N_27365);
or U27690 (N_27690,N_27442,N_27149);
xor U27691 (N_27691,N_27168,N_27354);
nand U27692 (N_27692,N_27344,N_27368);
nor U27693 (N_27693,N_27191,N_27259);
and U27694 (N_27694,N_27088,N_27391);
nand U27695 (N_27695,N_27484,N_27286);
or U27696 (N_27696,N_27559,N_27311);
and U27697 (N_27697,N_27470,N_27382);
and U27698 (N_27698,N_27220,N_27495);
and U27699 (N_27699,N_27372,N_27308);
xor U27700 (N_27700,N_27045,N_27264);
xor U27701 (N_27701,N_27526,N_27239);
nor U27702 (N_27702,N_27498,N_27047);
xor U27703 (N_27703,N_27463,N_27462);
xor U27704 (N_27704,N_27307,N_27242);
and U27705 (N_27705,N_27533,N_27519);
or U27706 (N_27706,N_27071,N_27058);
or U27707 (N_27707,N_27327,N_27098);
nor U27708 (N_27708,N_27429,N_27378);
xor U27709 (N_27709,N_27160,N_27317);
nand U27710 (N_27710,N_27186,N_27420);
xor U27711 (N_27711,N_27260,N_27424);
and U27712 (N_27712,N_27595,N_27238);
nand U27713 (N_27713,N_27028,N_27235);
or U27714 (N_27714,N_27474,N_27175);
xnor U27715 (N_27715,N_27003,N_27015);
nand U27716 (N_27716,N_27275,N_27451);
nor U27717 (N_27717,N_27257,N_27520);
nor U27718 (N_27718,N_27035,N_27314);
or U27719 (N_27719,N_27089,N_27349);
xnor U27720 (N_27720,N_27360,N_27444);
and U27721 (N_27721,N_27012,N_27565);
and U27722 (N_27722,N_27553,N_27016);
nand U27723 (N_27723,N_27422,N_27408);
and U27724 (N_27724,N_27084,N_27243);
and U27725 (N_27725,N_27590,N_27473);
nand U27726 (N_27726,N_27248,N_27465);
nor U27727 (N_27727,N_27440,N_27029);
xnor U27728 (N_27728,N_27090,N_27306);
nand U27729 (N_27729,N_27342,N_27087);
and U27730 (N_27730,N_27139,N_27066);
and U27731 (N_27731,N_27421,N_27568);
or U27732 (N_27732,N_27169,N_27173);
and U27733 (N_27733,N_27006,N_27435);
nor U27734 (N_27734,N_27535,N_27328);
and U27735 (N_27735,N_27548,N_27174);
or U27736 (N_27736,N_27085,N_27092);
xnor U27737 (N_27737,N_27564,N_27150);
or U27738 (N_27738,N_27190,N_27228);
or U27739 (N_27739,N_27126,N_27194);
or U27740 (N_27740,N_27443,N_27214);
nand U27741 (N_27741,N_27108,N_27377);
nand U27742 (N_27742,N_27544,N_27131);
nor U27743 (N_27743,N_27555,N_27067);
or U27744 (N_27744,N_27031,N_27549);
or U27745 (N_27745,N_27037,N_27213);
and U27746 (N_27746,N_27338,N_27315);
xor U27747 (N_27747,N_27157,N_27400);
nor U27748 (N_27748,N_27409,N_27337);
nand U27749 (N_27749,N_27077,N_27207);
nor U27750 (N_27750,N_27059,N_27477);
nor U27751 (N_27751,N_27283,N_27211);
and U27752 (N_27752,N_27289,N_27107);
nand U27753 (N_27753,N_27325,N_27414);
nor U27754 (N_27754,N_27543,N_27201);
and U27755 (N_27755,N_27133,N_27137);
nand U27756 (N_27756,N_27581,N_27562);
xnor U27757 (N_27757,N_27183,N_27598);
xor U27758 (N_27758,N_27367,N_27430);
nand U27759 (N_27759,N_27064,N_27506);
nand U27760 (N_27760,N_27551,N_27024);
and U27761 (N_27761,N_27188,N_27273);
nand U27762 (N_27762,N_27143,N_27587);
nor U27763 (N_27763,N_27510,N_27326);
and U27764 (N_27764,N_27261,N_27547);
xor U27765 (N_27765,N_27074,N_27373);
xnor U27766 (N_27766,N_27018,N_27123);
or U27767 (N_27767,N_27423,N_27445);
nor U27768 (N_27768,N_27203,N_27303);
nor U27769 (N_27769,N_27165,N_27556);
or U27770 (N_27770,N_27114,N_27329);
xor U27771 (N_27771,N_27236,N_27558);
nor U27772 (N_27772,N_27227,N_27044);
nand U27773 (N_27773,N_27483,N_27531);
and U27774 (N_27774,N_27393,N_27339);
or U27775 (N_27775,N_27030,N_27153);
nor U27776 (N_27776,N_27397,N_27417);
or U27777 (N_27777,N_27348,N_27002);
or U27778 (N_27778,N_27036,N_27189);
nor U27779 (N_27779,N_27386,N_27358);
xor U27780 (N_27780,N_27247,N_27586);
nand U27781 (N_27781,N_27223,N_27343);
or U27782 (N_27782,N_27285,N_27040);
nand U27783 (N_27783,N_27515,N_27398);
xor U27784 (N_27784,N_27455,N_27312);
and U27785 (N_27785,N_27141,N_27020);
or U27786 (N_27786,N_27046,N_27412);
and U27787 (N_27787,N_27138,N_27589);
or U27788 (N_27788,N_27374,N_27033);
and U27789 (N_27789,N_27072,N_27345);
xnor U27790 (N_27790,N_27251,N_27125);
and U27791 (N_27791,N_27166,N_27425);
nand U27792 (N_27792,N_27117,N_27093);
nor U27793 (N_27793,N_27406,N_27277);
nor U27794 (N_27794,N_27209,N_27103);
and U27795 (N_27795,N_27357,N_27262);
or U27796 (N_27796,N_27091,N_27232);
nand U27797 (N_27797,N_27415,N_27433);
nand U27798 (N_27798,N_27000,N_27596);
nor U27799 (N_27799,N_27389,N_27121);
nand U27800 (N_27800,N_27187,N_27384);
or U27801 (N_27801,N_27383,N_27432);
or U27802 (N_27802,N_27554,N_27512);
nor U27803 (N_27803,N_27528,N_27102);
nand U27804 (N_27804,N_27217,N_27407);
xor U27805 (N_27805,N_27200,N_27490);
nor U27806 (N_27806,N_27363,N_27516);
nor U27807 (N_27807,N_27530,N_27550);
nor U27808 (N_27808,N_27197,N_27500);
xnor U27809 (N_27809,N_27245,N_27158);
nand U27810 (N_27810,N_27436,N_27350);
xnor U27811 (N_27811,N_27101,N_27061);
or U27812 (N_27812,N_27278,N_27163);
xnor U27813 (N_27813,N_27146,N_27502);
xor U27814 (N_27814,N_27124,N_27319);
and U27815 (N_27815,N_27418,N_27300);
nor U27816 (N_27816,N_27078,N_27105);
and U27817 (N_27817,N_27478,N_27375);
nand U27818 (N_27818,N_27294,N_27195);
xnor U27819 (N_27819,N_27588,N_27578);
nand U27820 (N_27820,N_27480,N_27221);
nor U27821 (N_27821,N_27353,N_27104);
nor U27822 (N_27822,N_27268,N_27583);
nand U27823 (N_27823,N_27476,N_27545);
nor U27824 (N_27824,N_27291,N_27379);
nor U27825 (N_27825,N_27310,N_27320);
xor U27826 (N_27826,N_27240,N_27111);
nor U27827 (N_27827,N_27525,N_27073);
nand U27828 (N_27828,N_27475,N_27552);
xnor U27829 (N_27829,N_27222,N_27225);
nand U27830 (N_27830,N_27570,N_27298);
nand U27831 (N_27831,N_27296,N_27116);
and U27832 (N_27832,N_27048,N_27218);
xnor U27833 (N_27833,N_27467,N_27380);
or U27834 (N_27834,N_27270,N_27253);
and U27835 (N_27835,N_27594,N_27538);
and U27836 (N_27836,N_27471,N_27050);
and U27837 (N_27837,N_27292,N_27042);
nand U27838 (N_27838,N_27086,N_27019);
nor U27839 (N_27839,N_27511,N_27055);
nand U27840 (N_27840,N_27056,N_27152);
xor U27841 (N_27841,N_27401,N_27043);
or U27842 (N_27842,N_27321,N_27216);
xor U27843 (N_27843,N_27575,N_27540);
and U27844 (N_27844,N_27574,N_27057);
xor U27845 (N_27845,N_27441,N_27428);
xnor U27846 (N_27846,N_27576,N_27371);
nand U27847 (N_27847,N_27335,N_27537);
and U27848 (N_27848,N_27505,N_27054);
nor U27849 (N_27849,N_27541,N_27258);
nor U27850 (N_27850,N_27004,N_27052);
and U27851 (N_27851,N_27148,N_27266);
nor U27852 (N_27852,N_27171,N_27177);
and U27853 (N_27853,N_27359,N_27095);
nand U27854 (N_27854,N_27452,N_27464);
and U27855 (N_27855,N_27394,N_27094);
or U27856 (N_27856,N_27481,N_27162);
xor U27857 (N_27857,N_27215,N_27439);
nor U27858 (N_27858,N_27212,N_27226);
and U27859 (N_27859,N_27062,N_27147);
or U27860 (N_27860,N_27323,N_27491);
nor U27861 (N_27861,N_27492,N_27119);
or U27862 (N_27862,N_27579,N_27324);
xor U27863 (N_27863,N_27132,N_27192);
nand U27864 (N_27864,N_27395,N_27507);
nand U27865 (N_27865,N_27402,N_27128);
and U27866 (N_27866,N_27346,N_27571);
and U27867 (N_27867,N_27527,N_27224);
xnor U27868 (N_27868,N_27577,N_27193);
xnor U27869 (N_27869,N_27134,N_27025);
nand U27870 (N_27870,N_27396,N_27340);
nand U27871 (N_27871,N_27582,N_27392);
or U27872 (N_27872,N_27256,N_27254);
nand U27873 (N_27873,N_27460,N_27536);
or U27874 (N_27874,N_27026,N_27076);
nor U27875 (N_27875,N_27336,N_27182);
nor U27876 (N_27876,N_27185,N_27461);
nand U27877 (N_27877,N_27115,N_27524);
nand U27878 (N_27878,N_27410,N_27279);
nor U27879 (N_27879,N_27007,N_27532);
xnor U27880 (N_27880,N_27129,N_27493);
or U27881 (N_27881,N_27563,N_27099);
nor U27882 (N_27882,N_27381,N_27017);
nor U27883 (N_27883,N_27167,N_27265);
nand U27884 (N_27884,N_27334,N_27567);
or U27885 (N_27885,N_27403,N_27276);
or U27886 (N_27886,N_27413,N_27272);
or U27887 (N_27887,N_27034,N_27097);
or U27888 (N_27888,N_27023,N_27599);
and U27889 (N_27889,N_27331,N_27557);
xor U27890 (N_27890,N_27060,N_27513);
nor U27891 (N_27891,N_27404,N_27204);
nor U27892 (N_27892,N_27376,N_27179);
or U27893 (N_27893,N_27426,N_27229);
xnor U27894 (N_27894,N_27366,N_27459);
or U27895 (N_27895,N_27001,N_27249);
nand U27896 (N_27896,N_27482,N_27468);
and U27897 (N_27897,N_27351,N_27385);
nand U27898 (N_27898,N_27151,N_27370);
or U27899 (N_27899,N_27546,N_27068);
xnor U27900 (N_27900,N_27481,N_27101);
xnor U27901 (N_27901,N_27476,N_27130);
or U27902 (N_27902,N_27413,N_27551);
or U27903 (N_27903,N_27596,N_27313);
nand U27904 (N_27904,N_27331,N_27061);
nand U27905 (N_27905,N_27334,N_27099);
and U27906 (N_27906,N_27173,N_27441);
nand U27907 (N_27907,N_27479,N_27126);
or U27908 (N_27908,N_27366,N_27492);
and U27909 (N_27909,N_27545,N_27535);
nand U27910 (N_27910,N_27019,N_27532);
nor U27911 (N_27911,N_27205,N_27318);
nor U27912 (N_27912,N_27547,N_27137);
and U27913 (N_27913,N_27568,N_27457);
nand U27914 (N_27914,N_27546,N_27557);
nor U27915 (N_27915,N_27162,N_27205);
nand U27916 (N_27916,N_27029,N_27578);
xor U27917 (N_27917,N_27071,N_27183);
or U27918 (N_27918,N_27131,N_27169);
nand U27919 (N_27919,N_27415,N_27485);
or U27920 (N_27920,N_27267,N_27251);
nand U27921 (N_27921,N_27562,N_27384);
or U27922 (N_27922,N_27316,N_27449);
nor U27923 (N_27923,N_27141,N_27209);
xnor U27924 (N_27924,N_27275,N_27560);
or U27925 (N_27925,N_27531,N_27266);
or U27926 (N_27926,N_27514,N_27136);
and U27927 (N_27927,N_27217,N_27518);
xnor U27928 (N_27928,N_27365,N_27068);
or U27929 (N_27929,N_27286,N_27596);
or U27930 (N_27930,N_27340,N_27056);
xnor U27931 (N_27931,N_27234,N_27148);
or U27932 (N_27932,N_27257,N_27332);
nand U27933 (N_27933,N_27458,N_27579);
or U27934 (N_27934,N_27372,N_27266);
or U27935 (N_27935,N_27455,N_27186);
nand U27936 (N_27936,N_27359,N_27078);
or U27937 (N_27937,N_27539,N_27373);
nor U27938 (N_27938,N_27194,N_27576);
nor U27939 (N_27939,N_27405,N_27409);
or U27940 (N_27940,N_27254,N_27571);
nand U27941 (N_27941,N_27498,N_27017);
or U27942 (N_27942,N_27223,N_27396);
nor U27943 (N_27943,N_27421,N_27025);
nand U27944 (N_27944,N_27061,N_27478);
xnor U27945 (N_27945,N_27286,N_27470);
and U27946 (N_27946,N_27207,N_27197);
xor U27947 (N_27947,N_27563,N_27259);
or U27948 (N_27948,N_27295,N_27538);
nand U27949 (N_27949,N_27579,N_27015);
or U27950 (N_27950,N_27310,N_27298);
nand U27951 (N_27951,N_27321,N_27401);
or U27952 (N_27952,N_27181,N_27477);
xnor U27953 (N_27953,N_27436,N_27249);
or U27954 (N_27954,N_27322,N_27365);
nor U27955 (N_27955,N_27461,N_27334);
xnor U27956 (N_27956,N_27098,N_27152);
xnor U27957 (N_27957,N_27191,N_27064);
nor U27958 (N_27958,N_27367,N_27219);
nor U27959 (N_27959,N_27542,N_27420);
and U27960 (N_27960,N_27179,N_27505);
and U27961 (N_27961,N_27168,N_27557);
and U27962 (N_27962,N_27540,N_27537);
and U27963 (N_27963,N_27364,N_27386);
and U27964 (N_27964,N_27496,N_27596);
or U27965 (N_27965,N_27515,N_27557);
or U27966 (N_27966,N_27549,N_27482);
nor U27967 (N_27967,N_27024,N_27150);
nand U27968 (N_27968,N_27479,N_27338);
nor U27969 (N_27969,N_27218,N_27299);
or U27970 (N_27970,N_27102,N_27449);
nor U27971 (N_27971,N_27371,N_27556);
nand U27972 (N_27972,N_27408,N_27273);
and U27973 (N_27973,N_27341,N_27047);
and U27974 (N_27974,N_27531,N_27507);
nor U27975 (N_27975,N_27143,N_27461);
and U27976 (N_27976,N_27128,N_27414);
nor U27977 (N_27977,N_27454,N_27507);
or U27978 (N_27978,N_27589,N_27253);
and U27979 (N_27979,N_27059,N_27420);
nand U27980 (N_27980,N_27060,N_27211);
and U27981 (N_27981,N_27556,N_27019);
nor U27982 (N_27982,N_27205,N_27129);
and U27983 (N_27983,N_27146,N_27426);
and U27984 (N_27984,N_27360,N_27099);
or U27985 (N_27985,N_27573,N_27302);
xor U27986 (N_27986,N_27135,N_27196);
and U27987 (N_27987,N_27298,N_27260);
nand U27988 (N_27988,N_27555,N_27540);
or U27989 (N_27989,N_27069,N_27300);
and U27990 (N_27990,N_27183,N_27141);
xnor U27991 (N_27991,N_27185,N_27597);
xnor U27992 (N_27992,N_27548,N_27324);
or U27993 (N_27993,N_27415,N_27012);
xnor U27994 (N_27994,N_27090,N_27166);
nor U27995 (N_27995,N_27488,N_27299);
and U27996 (N_27996,N_27412,N_27099);
and U27997 (N_27997,N_27511,N_27052);
and U27998 (N_27998,N_27112,N_27117);
and U27999 (N_27999,N_27320,N_27486);
and U28000 (N_28000,N_27407,N_27556);
nor U28001 (N_28001,N_27056,N_27352);
xor U28002 (N_28002,N_27177,N_27221);
nand U28003 (N_28003,N_27019,N_27442);
and U28004 (N_28004,N_27102,N_27448);
or U28005 (N_28005,N_27390,N_27069);
nor U28006 (N_28006,N_27436,N_27340);
nand U28007 (N_28007,N_27090,N_27171);
and U28008 (N_28008,N_27422,N_27257);
nand U28009 (N_28009,N_27538,N_27313);
or U28010 (N_28010,N_27033,N_27026);
and U28011 (N_28011,N_27240,N_27040);
nand U28012 (N_28012,N_27031,N_27597);
or U28013 (N_28013,N_27405,N_27002);
or U28014 (N_28014,N_27285,N_27120);
or U28015 (N_28015,N_27300,N_27410);
or U28016 (N_28016,N_27299,N_27236);
and U28017 (N_28017,N_27392,N_27589);
nor U28018 (N_28018,N_27492,N_27408);
nand U28019 (N_28019,N_27319,N_27301);
nor U28020 (N_28020,N_27340,N_27324);
xnor U28021 (N_28021,N_27513,N_27117);
nor U28022 (N_28022,N_27141,N_27573);
nand U28023 (N_28023,N_27214,N_27500);
nor U28024 (N_28024,N_27591,N_27322);
xor U28025 (N_28025,N_27502,N_27124);
or U28026 (N_28026,N_27164,N_27209);
xor U28027 (N_28027,N_27450,N_27083);
nor U28028 (N_28028,N_27541,N_27288);
and U28029 (N_28029,N_27271,N_27586);
or U28030 (N_28030,N_27282,N_27527);
or U28031 (N_28031,N_27564,N_27388);
and U28032 (N_28032,N_27578,N_27137);
and U28033 (N_28033,N_27253,N_27229);
and U28034 (N_28034,N_27190,N_27068);
and U28035 (N_28035,N_27368,N_27189);
or U28036 (N_28036,N_27255,N_27552);
nor U28037 (N_28037,N_27543,N_27482);
nor U28038 (N_28038,N_27384,N_27540);
nor U28039 (N_28039,N_27102,N_27361);
or U28040 (N_28040,N_27272,N_27017);
and U28041 (N_28041,N_27421,N_27418);
nor U28042 (N_28042,N_27359,N_27003);
and U28043 (N_28043,N_27430,N_27516);
nand U28044 (N_28044,N_27398,N_27418);
nor U28045 (N_28045,N_27466,N_27299);
nor U28046 (N_28046,N_27074,N_27404);
and U28047 (N_28047,N_27048,N_27148);
xor U28048 (N_28048,N_27446,N_27319);
or U28049 (N_28049,N_27355,N_27289);
or U28050 (N_28050,N_27095,N_27586);
nor U28051 (N_28051,N_27110,N_27339);
xnor U28052 (N_28052,N_27013,N_27426);
xor U28053 (N_28053,N_27068,N_27470);
or U28054 (N_28054,N_27210,N_27576);
nor U28055 (N_28055,N_27450,N_27007);
xor U28056 (N_28056,N_27114,N_27026);
or U28057 (N_28057,N_27420,N_27196);
and U28058 (N_28058,N_27115,N_27369);
and U28059 (N_28059,N_27124,N_27508);
or U28060 (N_28060,N_27248,N_27045);
nor U28061 (N_28061,N_27501,N_27111);
nand U28062 (N_28062,N_27244,N_27373);
nand U28063 (N_28063,N_27050,N_27047);
nand U28064 (N_28064,N_27072,N_27421);
xor U28065 (N_28065,N_27476,N_27158);
nand U28066 (N_28066,N_27137,N_27441);
or U28067 (N_28067,N_27012,N_27178);
nor U28068 (N_28068,N_27020,N_27142);
or U28069 (N_28069,N_27013,N_27098);
nand U28070 (N_28070,N_27327,N_27141);
nor U28071 (N_28071,N_27248,N_27178);
nor U28072 (N_28072,N_27443,N_27449);
xnor U28073 (N_28073,N_27553,N_27532);
nand U28074 (N_28074,N_27387,N_27588);
xnor U28075 (N_28075,N_27244,N_27502);
nor U28076 (N_28076,N_27471,N_27494);
or U28077 (N_28077,N_27312,N_27347);
xor U28078 (N_28078,N_27287,N_27108);
nand U28079 (N_28079,N_27583,N_27324);
nor U28080 (N_28080,N_27378,N_27367);
xor U28081 (N_28081,N_27277,N_27339);
or U28082 (N_28082,N_27508,N_27195);
or U28083 (N_28083,N_27275,N_27127);
nand U28084 (N_28084,N_27009,N_27207);
xor U28085 (N_28085,N_27462,N_27566);
or U28086 (N_28086,N_27193,N_27368);
and U28087 (N_28087,N_27119,N_27140);
or U28088 (N_28088,N_27585,N_27021);
nand U28089 (N_28089,N_27113,N_27218);
xor U28090 (N_28090,N_27532,N_27387);
nand U28091 (N_28091,N_27392,N_27154);
nor U28092 (N_28092,N_27140,N_27222);
xor U28093 (N_28093,N_27539,N_27352);
nand U28094 (N_28094,N_27333,N_27355);
nand U28095 (N_28095,N_27315,N_27033);
nor U28096 (N_28096,N_27335,N_27302);
nor U28097 (N_28097,N_27339,N_27480);
nor U28098 (N_28098,N_27573,N_27099);
and U28099 (N_28099,N_27581,N_27248);
and U28100 (N_28100,N_27026,N_27420);
xnor U28101 (N_28101,N_27454,N_27595);
or U28102 (N_28102,N_27241,N_27511);
or U28103 (N_28103,N_27258,N_27475);
nand U28104 (N_28104,N_27411,N_27344);
or U28105 (N_28105,N_27293,N_27241);
and U28106 (N_28106,N_27095,N_27165);
or U28107 (N_28107,N_27287,N_27113);
or U28108 (N_28108,N_27241,N_27194);
nor U28109 (N_28109,N_27557,N_27390);
or U28110 (N_28110,N_27285,N_27137);
or U28111 (N_28111,N_27295,N_27597);
and U28112 (N_28112,N_27283,N_27467);
nand U28113 (N_28113,N_27580,N_27511);
nand U28114 (N_28114,N_27399,N_27369);
or U28115 (N_28115,N_27504,N_27093);
or U28116 (N_28116,N_27179,N_27478);
nor U28117 (N_28117,N_27288,N_27437);
nand U28118 (N_28118,N_27351,N_27210);
nand U28119 (N_28119,N_27418,N_27593);
xnor U28120 (N_28120,N_27036,N_27574);
xor U28121 (N_28121,N_27499,N_27221);
nor U28122 (N_28122,N_27589,N_27497);
nor U28123 (N_28123,N_27084,N_27235);
nand U28124 (N_28124,N_27041,N_27076);
and U28125 (N_28125,N_27199,N_27020);
nand U28126 (N_28126,N_27013,N_27595);
nand U28127 (N_28127,N_27133,N_27357);
or U28128 (N_28128,N_27449,N_27429);
nand U28129 (N_28129,N_27254,N_27005);
xor U28130 (N_28130,N_27068,N_27224);
nor U28131 (N_28131,N_27163,N_27106);
nand U28132 (N_28132,N_27126,N_27467);
and U28133 (N_28133,N_27076,N_27570);
nor U28134 (N_28134,N_27495,N_27570);
and U28135 (N_28135,N_27583,N_27448);
xnor U28136 (N_28136,N_27405,N_27266);
nand U28137 (N_28137,N_27554,N_27264);
xor U28138 (N_28138,N_27234,N_27418);
and U28139 (N_28139,N_27337,N_27260);
and U28140 (N_28140,N_27428,N_27399);
and U28141 (N_28141,N_27363,N_27288);
nor U28142 (N_28142,N_27368,N_27146);
nand U28143 (N_28143,N_27347,N_27367);
nor U28144 (N_28144,N_27175,N_27150);
nor U28145 (N_28145,N_27069,N_27587);
nand U28146 (N_28146,N_27360,N_27598);
or U28147 (N_28147,N_27023,N_27484);
nor U28148 (N_28148,N_27325,N_27473);
xnor U28149 (N_28149,N_27465,N_27467);
nor U28150 (N_28150,N_27150,N_27114);
and U28151 (N_28151,N_27345,N_27161);
xnor U28152 (N_28152,N_27472,N_27585);
and U28153 (N_28153,N_27459,N_27302);
nand U28154 (N_28154,N_27154,N_27267);
nor U28155 (N_28155,N_27299,N_27546);
nand U28156 (N_28156,N_27488,N_27094);
nand U28157 (N_28157,N_27150,N_27375);
xnor U28158 (N_28158,N_27012,N_27194);
nor U28159 (N_28159,N_27308,N_27596);
xor U28160 (N_28160,N_27172,N_27139);
and U28161 (N_28161,N_27215,N_27054);
and U28162 (N_28162,N_27174,N_27342);
nor U28163 (N_28163,N_27466,N_27187);
and U28164 (N_28164,N_27280,N_27231);
and U28165 (N_28165,N_27286,N_27215);
nand U28166 (N_28166,N_27029,N_27292);
or U28167 (N_28167,N_27095,N_27070);
nand U28168 (N_28168,N_27446,N_27336);
nand U28169 (N_28169,N_27180,N_27195);
xor U28170 (N_28170,N_27144,N_27181);
xnor U28171 (N_28171,N_27083,N_27254);
nor U28172 (N_28172,N_27292,N_27137);
nor U28173 (N_28173,N_27577,N_27056);
xor U28174 (N_28174,N_27122,N_27213);
nand U28175 (N_28175,N_27059,N_27291);
nor U28176 (N_28176,N_27146,N_27113);
xnor U28177 (N_28177,N_27569,N_27053);
nand U28178 (N_28178,N_27088,N_27096);
xnor U28179 (N_28179,N_27408,N_27047);
or U28180 (N_28180,N_27311,N_27183);
nand U28181 (N_28181,N_27178,N_27220);
and U28182 (N_28182,N_27524,N_27435);
and U28183 (N_28183,N_27454,N_27151);
and U28184 (N_28184,N_27332,N_27384);
nor U28185 (N_28185,N_27461,N_27332);
nor U28186 (N_28186,N_27577,N_27117);
nand U28187 (N_28187,N_27274,N_27319);
nor U28188 (N_28188,N_27354,N_27063);
xnor U28189 (N_28189,N_27525,N_27199);
and U28190 (N_28190,N_27598,N_27184);
nand U28191 (N_28191,N_27255,N_27010);
or U28192 (N_28192,N_27562,N_27152);
xor U28193 (N_28193,N_27446,N_27092);
nor U28194 (N_28194,N_27014,N_27534);
xor U28195 (N_28195,N_27393,N_27260);
xor U28196 (N_28196,N_27024,N_27566);
and U28197 (N_28197,N_27092,N_27027);
nand U28198 (N_28198,N_27556,N_27048);
xor U28199 (N_28199,N_27068,N_27333);
nand U28200 (N_28200,N_27868,N_27642);
or U28201 (N_28201,N_28104,N_28134);
nor U28202 (N_28202,N_27869,N_28149);
or U28203 (N_28203,N_27653,N_27749);
or U28204 (N_28204,N_27841,N_27704);
xnor U28205 (N_28205,N_27644,N_27662);
nand U28206 (N_28206,N_27787,N_27742);
and U28207 (N_28207,N_27702,N_28084);
and U28208 (N_28208,N_27772,N_27615);
nand U28209 (N_28209,N_28004,N_28012);
and U28210 (N_28210,N_27832,N_27935);
xnor U28211 (N_28211,N_28066,N_27923);
xnor U28212 (N_28212,N_28140,N_27915);
or U28213 (N_28213,N_27974,N_28197);
nand U28214 (N_28214,N_27760,N_28015);
nor U28215 (N_28215,N_28169,N_27754);
or U28216 (N_28216,N_28037,N_28038);
nor U28217 (N_28217,N_28135,N_27689);
and U28218 (N_28218,N_27831,N_27724);
nor U28219 (N_28219,N_27850,N_27759);
nor U28220 (N_28220,N_28009,N_27784);
nand U28221 (N_28221,N_28050,N_28046);
and U28222 (N_28222,N_27898,N_27778);
and U28223 (N_28223,N_27911,N_27984);
nor U28224 (N_28224,N_27985,N_28101);
xnor U28225 (N_28225,N_27649,N_28166);
nor U28226 (N_28226,N_28044,N_27849);
nand U28227 (N_28227,N_27703,N_28001);
or U28228 (N_28228,N_27908,N_27848);
and U28229 (N_28229,N_28145,N_27651);
and U28230 (N_28230,N_27757,N_28087);
or U28231 (N_28231,N_27957,N_27639);
xor U28232 (N_28232,N_28040,N_28157);
xnor U28233 (N_28233,N_28088,N_27794);
or U28234 (N_28234,N_27840,N_27876);
xnor U28235 (N_28235,N_27620,N_27942);
xor U28236 (N_28236,N_28177,N_27780);
xnor U28237 (N_28237,N_28144,N_28010);
xor U28238 (N_28238,N_27862,N_27874);
and U28239 (N_28239,N_28195,N_28143);
and U28240 (N_28240,N_27808,N_28022);
nor U28241 (N_28241,N_27924,N_27687);
xor U28242 (N_28242,N_27830,N_27654);
xor U28243 (N_28243,N_27885,N_27939);
xor U28244 (N_28244,N_27796,N_27765);
and U28245 (N_28245,N_28178,N_27652);
and U28246 (N_28246,N_28071,N_28192);
nor U28247 (N_28247,N_28198,N_28196);
xor U28248 (N_28248,N_27920,N_27695);
nor U28249 (N_28249,N_27902,N_27810);
nand U28250 (N_28250,N_27975,N_27916);
xnor U28251 (N_28251,N_28152,N_27931);
nand U28252 (N_28252,N_28128,N_27851);
nor U28253 (N_28253,N_28094,N_27999);
nand U28254 (N_28254,N_27956,N_28077);
xor U28255 (N_28255,N_27774,N_27725);
and U28256 (N_28256,N_27616,N_27606);
nand U28257 (N_28257,N_27827,N_27886);
nor U28258 (N_28258,N_27839,N_28172);
and U28259 (N_28259,N_28091,N_27755);
xnor U28260 (N_28260,N_27601,N_27640);
nor U28261 (N_28261,N_28051,N_28173);
or U28262 (N_28262,N_28163,N_28043);
nand U28263 (N_28263,N_27979,N_27681);
xnor U28264 (N_28264,N_28019,N_27896);
nor U28265 (N_28265,N_28139,N_27610);
and U28266 (N_28266,N_27990,N_27867);
nand U28267 (N_28267,N_27801,N_27962);
and U28268 (N_28268,N_27903,N_27929);
nand U28269 (N_28269,N_27613,N_27762);
nand U28270 (N_28270,N_28119,N_27680);
nand U28271 (N_28271,N_28083,N_27803);
or U28272 (N_28272,N_27980,N_27641);
and U28273 (N_28273,N_27927,N_28093);
nand U28274 (N_28274,N_28112,N_27970);
or U28275 (N_28275,N_28158,N_27629);
or U28276 (N_28276,N_27743,N_28186);
or U28277 (N_28277,N_27806,N_27953);
and U28278 (N_28278,N_27822,N_28058);
nor U28279 (N_28279,N_27709,N_28183);
xor U28280 (N_28280,N_27633,N_28095);
nor U28281 (N_28281,N_28164,N_28098);
or U28282 (N_28282,N_28124,N_27878);
nor U28283 (N_28283,N_27873,N_27661);
or U28284 (N_28284,N_27861,N_27945);
and U28285 (N_28285,N_27779,N_28185);
nor U28286 (N_28286,N_28030,N_27845);
and U28287 (N_28287,N_28137,N_28026);
nand U28288 (N_28288,N_28054,N_27855);
and U28289 (N_28289,N_27993,N_28193);
or U28290 (N_28290,N_28146,N_28007);
or U28291 (N_28291,N_27864,N_27701);
nor U28292 (N_28292,N_27734,N_27852);
xnor U28293 (N_28293,N_27946,N_28133);
nor U28294 (N_28294,N_28153,N_27952);
and U28295 (N_28295,N_27968,N_27628);
and U28296 (N_28296,N_27837,N_28102);
nand U28297 (N_28297,N_27688,N_27786);
nand U28298 (N_28298,N_27949,N_27752);
nor U28299 (N_28299,N_28125,N_28118);
and U28300 (N_28300,N_28089,N_27705);
or U28301 (N_28301,N_27722,N_28086);
xnor U28302 (N_28302,N_27948,N_27947);
or U28303 (N_28303,N_27731,N_28148);
nand U28304 (N_28304,N_27895,N_28041);
xor U28305 (N_28305,N_27727,N_28069);
xnor U28306 (N_28306,N_27775,N_27815);
or U28307 (N_28307,N_27904,N_27892);
xnor U28308 (N_28308,N_28179,N_27614);
nor U28309 (N_28309,N_27789,N_27671);
xnor U28310 (N_28310,N_27684,N_28132);
nor U28311 (N_28311,N_27820,N_28073);
nand U28312 (N_28312,N_27604,N_27693);
or U28313 (N_28313,N_27624,N_27826);
or U28314 (N_28314,N_27863,N_28053);
xnor U28315 (N_28315,N_27977,N_27901);
nand U28316 (N_28316,N_27676,N_28078);
xnor U28317 (N_28317,N_28070,N_27730);
xnor U28318 (N_28318,N_27991,N_28106);
nor U28319 (N_28319,N_27881,N_27951);
xor U28320 (N_28320,N_27781,N_27744);
and U28321 (N_28321,N_27802,N_27685);
or U28322 (N_28322,N_28018,N_27618);
nor U28323 (N_28323,N_27891,N_28047);
nand U28324 (N_28324,N_27738,N_27768);
nor U28325 (N_28325,N_28020,N_27632);
or U28326 (N_28326,N_27713,N_27737);
nand U28327 (N_28327,N_27710,N_27978);
nor U28328 (N_28328,N_27871,N_27894);
nor U28329 (N_28329,N_28082,N_27995);
nand U28330 (N_28330,N_27888,N_28151);
and U28331 (N_28331,N_28068,N_27686);
nand U28332 (N_28332,N_27699,N_28055);
nor U28333 (N_28333,N_27976,N_27795);
xor U28334 (N_28334,N_27989,N_27748);
nand U28335 (N_28335,N_27833,N_27865);
or U28336 (N_28336,N_27807,N_28168);
nor U28337 (N_28337,N_28029,N_27720);
nor U28338 (N_28338,N_27797,N_27660);
and U28339 (N_28339,N_27967,N_28110);
nor U28340 (N_28340,N_27859,N_28079);
nor U28341 (N_28341,N_27858,N_27809);
nor U28342 (N_28342,N_28108,N_27636);
xor U28343 (N_28343,N_28011,N_27773);
and U28344 (N_28344,N_28033,N_27758);
or U28345 (N_28345,N_27843,N_28080);
or U28346 (N_28346,N_27740,N_28031);
nand U28347 (N_28347,N_27994,N_28167);
and U28348 (N_28348,N_27630,N_27691);
nor U28349 (N_28349,N_27756,N_28107);
nand U28350 (N_28350,N_27971,N_27791);
xnor U28351 (N_28351,N_28121,N_27608);
nand U28352 (N_28352,N_28190,N_27792);
and U28353 (N_28353,N_28131,N_27712);
nor U28354 (N_28354,N_27969,N_27623);
or U28355 (N_28355,N_27783,N_28103);
and U28356 (N_28356,N_28052,N_27696);
and U28357 (N_28357,N_28142,N_27626);
nor U28358 (N_28358,N_27764,N_28187);
nor U28359 (N_28359,N_28016,N_27925);
xor U28360 (N_28360,N_27657,N_27860);
nand U28361 (N_28361,N_27659,N_27926);
and U28362 (N_28362,N_27782,N_27893);
or U28363 (N_28363,N_28136,N_27958);
xnor U28364 (N_28364,N_27847,N_27882);
nand U28365 (N_28365,N_27741,N_27866);
or U28366 (N_28366,N_27655,N_27824);
nand U28367 (N_28367,N_28174,N_28072);
xnor U28368 (N_28368,N_28141,N_28024);
or U28369 (N_28369,N_27761,N_27918);
nor U28370 (N_28370,N_27645,N_27668);
nor U28371 (N_28371,N_27825,N_28162);
and U28372 (N_28372,N_27943,N_28059);
nand U28373 (N_28373,N_28000,N_28159);
or U28374 (N_28374,N_27692,N_28042);
or U28375 (N_28375,N_27900,N_27816);
or U28376 (N_28376,N_27955,N_27828);
and U28377 (N_28377,N_27637,N_27880);
nor U28378 (N_28378,N_27932,N_27798);
nand U28379 (N_28379,N_28156,N_27997);
or U28380 (N_28380,N_27732,N_28048);
and U28381 (N_28381,N_27872,N_27718);
nor U28382 (N_28382,N_28180,N_28075);
xnor U28383 (N_28383,N_27788,N_27631);
nand U28384 (N_28384,N_27934,N_27763);
or U28385 (N_28385,N_27887,N_27635);
or U28386 (N_28386,N_28130,N_27853);
nand U28387 (N_28387,N_27811,N_28032);
nand U28388 (N_28388,N_27733,N_28126);
and U28389 (N_28389,N_28199,N_27996);
nor U28390 (N_28390,N_27634,N_27875);
and U28391 (N_28391,N_27964,N_27607);
and U28392 (N_28392,N_27711,N_27921);
or U28393 (N_28393,N_28189,N_27805);
or U28394 (N_28394,N_27966,N_27981);
and U28395 (N_28395,N_27890,N_27650);
or U28396 (N_28396,N_28006,N_28002);
xnor U28397 (N_28397,N_28165,N_27821);
xnor U28398 (N_28398,N_27667,N_27658);
nor U28399 (N_28399,N_27646,N_27690);
and U28400 (N_28400,N_28074,N_28116);
nor U28401 (N_28401,N_28194,N_27954);
nand U28402 (N_28402,N_27603,N_27884);
or U28403 (N_28403,N_27619,N_27913);
or U28404 (N_28404,N_28013,N_28155);
nand U28405 (N_28405,N_27877,N_28064);
nand U28406 (N_28406,N_28115,N_27998);
xnor U28407 (N_28407,N_27656,N_28063);
or U28408 (N_28408,N_27941,N_27679);
or U28409 (N_28409,N_27627,N_28176);
nand U28410 (N_28410,N_27917,N_28138);
or U28411 (N_28411,N_28100,N_27972);
nand U28412 (N_28412,N_28109,N_27829);
nand U28413 (N_28413,N_27836,N_28096);
xnor U28414 (N_28414,N_28036,N_27870);
or U28415 (N_28415,N_27889,N_27670);
or U28416 (N_28416,N_27625,N_27910);
xor U28417 (N_28417,N_27897,N_28160);
xnor U28418 (N_28418,N_27683,N_28171);
xnor U28419 (N_28419,N_27602,N_27987);
nor U28420 (N_28420,N_27983,N_27677);
nor U28421 (N_28421,N_27643,N_27856);
or U28422 (N_28422,N_28092,N_27906);
and U28423 (N_28423,N_27817,N_27766);
and U28424 (N_28424,N_28023,N_27747);
or U28425 (N_28425,N_27682,N_27750);
xnor U28426 (N_28426,N_27694,N_28150);
nor U28427 (N_28427,N_27919,N_27771);
nand U28428 (N_28428,N_27936,N_27767);
and U28429 (N_28429,N_27930,N_27799);
or U28430 (N_28430,N_27770,N_27665);
and U28431 (N_28431,N_27899,N_28127);
and U28432 (N_28432,N_27961,N_28017);
xor U28433 (N_28433,N_27735,N_27736);
nand U28434 (N_28434,N_27960,N_28097);
and U28435 (N_28435,N_28049,N_28175);
nor U28436 (N_28436,N_28028,N_28129);
nand U28437 (N_28437,N_27838,N_28045);
xor U28438 (N_28438,N_27726,N_27664);
and U28439 (N_28439,N_27813,N_28014);
nand U28440 (N_28440,N_28188,N_27835);
xnor U28441 (N_28441,N_28067,N_28123);
and U28442 (N_28442,N_27800,N_27719);
and U28443 (N_28443,N_27950,N_27940);
and U28444 (N_28444,N_27600,N_28057);
or U28445 (N_28445,N_28035,N_27973);
nand U28446 (N_28446,N_28056,N_28147);
and U28447 (N_28447,N_28034,N_27793);
xor U28448 (N_28448,N_28027,N_27746);
nand U28449 (N_28449,N_28113,N_28005);
nor U28450 (N_28450,N_27729,N_27988);
xor U28451 (N_28451,N_28021,N_27716);
or U28452 (N_28452,N_27938,N_27905);
or U28453 (N_28453,N_27612,N_28182);
or U28454 (N_28454,N_28025,N_27922);
nor U28455 (N_28455,N_27609,N_28099);
nor U28456 (N_28456,N_28008,N_27818);
nor U28457 (N_28457,N_27673,N_27697);
nor U28458 (N_28458,N_27982,N_28065);
xor U28459 (N_28459,N_27721,N_28122);
nand U28460 (N_28460,N_27672,N_27714);
nor U28461 (N_28461,N_27647,N_27777);
nor U28462 (N_28462,N_27728,N_28003);
and U28463 (N_28463,N_28060,N_27854);
or U28464 (N_28464,N_27819,N_27804);
or U28465 (N_28465,N_27790,N_27717);
and U28466 (N_28466,N_27776,N_27605);
nor U28467 (N_28467,N_28170,N_28184);
nor U28468 (N_28468,N_28105,N_27959);
or U28469 (N_28469,N_28181,N_27883);
xnor U28470 (N_28470,N_27638,N_27944);
nor U28471 (N_28471,N_27907,N_27617);
and U28472 (N_28472,N_27909,N_28076);
nand U28473 (N_28473,N_27611,N_28117);
xor U28474 (N_28474,N_27769,N_28161);
and U28475 (N_28475,N_27992,N_27842);
nand U28476 (N_28476,N_27663,N_27823);
nand U28477 (N_28477,N_28114,N_27834);
or U28478 (N_28478,N_27933,N_28090);
nor U28479 (N_28479,N_28154,N_28120);
nor U28480 (N_28480,N_28062,N_27785);
xnor U28481 (N_28481,N_27912,N_28085);
xor U28482 (N_28482,N_27739,N_27879);
and U28483 (N_28483,N_27708,N_27914);
or U28484 (N_28484,N_27814,N_27666);
xnor U28485 (N_28485,N_27857,N_27928);
and U28486 (N_28486,N_27715,N_27700);
xor U28487 (N_28487,N_27986,N_28111);
or U28488 (N_28488,N_27675,N_27622);
xor U28489 (N_28489,N_27745,N_27751);
or U28490 (N_28490,N_27844,N_27621);
or U28491 (N_28491,N_27648,N_28081);
or U28492 (N_28492,N_27723,N_27753);
xor U28493 (N_28493,N_27669,N_27963);
nand U28494 (N_28494,N_27812,N_27707);
and U28495 (N_28495,N_27698,N_28191);
and U28496 (N_28496,N_27706,N_27674);
nor U28497 (N_28497,N_27846,N_27678);
nor U28498 (N_28498,N_28039,N_28061);
nor U28499 (N_28499,N_27965,N_27937);
nor U28500 (N_28500,N_27922,N_27931);
and U28501 (N_28501,N_27956,N_27959);
and U28502 (N_28502,N_27883,N_28061);
xor U28503 (N_28503,N_27618,N_28047);
nand U28504 (N_28504,N_28076,N_27992);
nor U28505 (N_28505,N_27965,N_28126);
nor U28506 (N_28506,N_28188,N_28038);
or U28507 (N_28507,N_28025,N_27987);
nor U28508 (N_28508,N_27875,N_27937);
nand U28509 (N_28509,N_27769,N_27833);
xnor U28510 (N_28510,N_28188,N_27779);
and U28511 (N_28511,N_27642,N_28007);
and U28512 (N_28512,N_28054,N_27853);
nor U28513 (N_28513,N_27915,N_27981);
and U28514 (N_28514,N_27949,N_28077);
and U28515 (N_28515,N_27607,N_27657);
xor U28516 (N_28516,N_27862,N_27829);
or U28517 (N_28517,N_28133,N_28096);
or U28518 (N_28518,N_27712,N_27800);
nor U28519 (N_28519,N_27639,N_27675);
or U28520 (N_28520,N_28188,N_27618);
nand U28521 (N_28521,N_27742,N_27924);
or U28522 (N_28522,N_28116,N_27999);
nand U28523 (N_28523,N_27896,N_28194);
nor U28524 (N_28524,N_27927,N_28188);
nand U28525 (N_28525,N_27636,N_27675);
nand U28526 (N_28526,N_28089,N_28005);
or U28527 (N_28527,N_28139,N_27819);
nand U28528 (N_28528,N_27921,N_27767);
xor U28529 (N_28529,N_28049,N_27823);
nor U28530 (N_28530,N_27641,N_27696);
nand U28531 (N_28531,N_27910,N_28145);
nand U28532 (N_28532,N_27789,N_28075);
and U28533 (N_28533,N_27742,N_28029);
nor U28534 (N_28534,N_28182,N_27675);
or U28535 (N_28535,N_27659,N_27922);
xnor U28536 (N_28536,N_27812,N_28047);
xnor U28537 (N_28537,N_27900,N_27899);
or U28538 (N_28538,N_28085,N_28124);
or U28539 (N_28539,N_27917,N_28173);
nand U28540 (N_28540,N_27783,N_28133);
and U28541 (N_28541,N_28127,N_27724);
nand U28542 (N_28542,N_27699,N_27875);
and U28543 (N_28543,N_27925,N_27830);
xor U28544 (N_28544,N_27702,N_27606);
nand U28545 (N_28545,N_28183,N_27859);
or U28546 (N_28546,N_27812,N_28185);
and U28547 (N_28547,N_27721,N_28059);
xor U28548 (N_28548,N_27899,N_28031);
nand U28549 (N_28549,N_28106,N_27811);
nand U28550 (N_28550,N_27683,N_27784);
xor U28551 (N_28551,N_27715,N_27645);
and U28552 (N_28552,N_27785,N_27799);
nand U28553 (N_28553,N_27892,N_27619);
xor U28554 (N_28554,N_28045,N_28151);
nand U28555 (N_28555,N_27728,N_27671);
nand U28556 (N_28556,N_27850,N_27768);
nor U28557 (N_28557,N_27987,N_27977);
nand U28558 (N_28558,N_28024,N_27682);
or U28559 (N_28559,N_27851,N_27911);
nor U28560 (N_28560,N_28079,N_28154);
nor U28561 (N_28561,N_28092,N_28118);
nor U28562 (N_28562,N_27807,N_27976);
nor U28563 (N_28563,N_27923,N_27960);
nor U28564 (N_28564,N_27775,N_27994);
and U28565 (N_28565,N_27634,N_27697);
nor U28566 (N_28566,N_27912,N_28190);
xor U28567 (N_28567,N_27719,N_27622);
nor U28568 (N_28568,N_27772,N_27676);
nand U28569 (N_28569,N_27798,N_27843);
nor U28570 (N_28570,N_28145,N_27883);
nor U28571 (N_28571,N_28175,N_27687);
or U28572 (N_28572,N_27966,N_27964);
or U28573 (N_28573,N_27928,N_27640);
and U28574 (N_28574,N_27700,N_27849);
and U28575 (N_28575,N_27992,N_27949);
nand U28576 (N_28576,N_27863,N_28088);
xnor U28577 (N_28577,N_28093,N_28146);
or U28578 (N_28578,N_28152,N_27652);
xnor U28579 (N_28579,N_27769,N_27659);
or U28580 (N_28580,N_27873,N_27660);
or U28581 (N_28581,N_27839,N_27936);
xor U28582 (N_28582,N_27626,N_27875);
and U28583 (N_28583,N_28094,N_27863);
nor U28584 (N_28584,N_28194,N_27931);
or U28585 (N_28585,N_28199,N_28163);
nor U28586 (N_28586,N_28029,N_28159);
or U28587 (N_28587,N_28158,N_27725);
or U28588 (N_28588,N_27695,N_27988);
nor U28589 (N_28589,N_27653,N_28094);
or U28590 (N_28590,N_28029,N_28013);
or U28591 (N_28591,N_27881,N_27896);
and U28592 (N_28592,N_28028,N_27999);
nor U28593 (N_28593,N_27711,N_28115);
and U28594 (N_28594,N_27966,N_27802);
xnor U28595 (N_28595,N_28175,N_27657);
and U28596 (N_28596,N_27857,N_27923);
nor U28597 (N_28597,N_28176,N_27689);
or U28598 (N_28598,N_27714,N_28155);
xnor U28599 (N_28599,N_27764,N_27941);
or U28600 (N_28600,N_28057,N_27627);
nor U28601 (N_28601,N_27860,N_27730);
xnor U28602 (N_28602,N_28010,N_27691);
nand U28603 (N_28603,N_27739,N_27689);
nand U28604 (N_28604,N_27622,N_27616);
and U28605 (N_28605,N_27975,N_27912);
or U28606 (N_28606,N_28195,N_28075);
nor U28607 (N_28607,N_28108,N_27657);
or U28608 (N_28608,N_27609,N_28041);
or U28609 (N_28609,N_27625,N_28068);
xnor U28610 (N_28610,N_27737,N_27750);
nor U28611 (N_28611,N_28175,N_28068);
nand U28612 (N_28612,N_27671,N_27604);
nand U28613 (N_28613,N_28080,N_27659);
xor U28614 (N_28614,N_27811,N_27938);
or U28615 (N_28615,N_27980,N_27856);
xnor U28616 (N_28616,N_27652,N_27638);
nand U28617 (N_28617,N_27679,N_28197);
or U28618 (N_28618,N_27784,N_28168);
nand U28619 (N_28619,N_27844,N_27614);
and U28620 (N_28620,N_27949,N_27723);
and U28621 (N_28621,N_27973,N_28028);
and U28622 (N_28622,N_27789,N_27691);
nor U28623 (N_28623,N_28155,N_27731);
and U28624 (N_28624,N_27808,N_28024);
nor U28625 (N_28625,N_27837,N_27624);
nor U28626 (N_28626,N_27833,N_28180);
xnor U28627 (N_28627,N_28021,N_27945);
or U28628 (N_28628,N_27907,N_27930);
xor U28629 (N_28629,N_27930,N_27719);
xnor U28630 (N_28630,N_28116,N_27726);
or U28631 (N_28631,N_28039,N_28135);
xor U28632 (N_28632,N_27611,N_28146);
or U28633 (N_28633,N_27698,N_27694);
and U28634 (N_28634,N_27865,N_27747);
nor U28635 (N_28635,N_28131,N_27648);
or U28636 (N_28636,N_27714,N_28194);
nor U28637 (N_28637,N_27652,N_27931);
and U28638 (N_28638,N_27836,N_27930);
and U28639 (N_28639,N_28178,N_28033);
and U28640 (N_28640,N_27678,N_28138);
and U28641 (N_28641,N_28193,N_27703);
nand U28642 (N_28642,N_27732,N_28167);
xor U28643 (N_28643,N_27963,N_27668);
and U28644 (N_28644,N_27765,N_28006);
and U28645 (N_28645,N_27733,N_27817);
and U28646 (N_28646,N_28142,N_28155);
nor U28647 (N_28647,N_27936,N_28014);
nor U28648 (N_28648,N_27954,N_27682);
xnor U28649 (N_28649,N_28171,N_27647);
nand U28650 (N_28650,N_27835,N_27615);
nand U28651 (N_28651,N_28097,N_27965);
or U28652 (N_28652,N_28107,N_28120);
nor U28653 (N_28653,N_28118,N_28008);
and U28654 (N_28654,N_27890,N_28193);
and U28655 (N_28655,N_27694,N_27748);
xnor U28656 (N_28656,N_27823,N_27710);
or U28657 (N_28657,N_27942,N_27969);
nand U28658 (N_28658,N_28131,N_27957);
xnor U28659 (N_28659,N_27729,N_27871);
xnor U28660 (N_28660,N_28078,N_27826);
nor U28661 (N_28661,N_27980,N_28128);
nand U28662 (N_28662,N_27837,N_27770);
xnor U28663 (N_28663,N_27708,N_28165);
nand U28664 (N_28664,N_28115,N_28010);
and U28665 (N_28665,N_27711,N_27992);
or U28666 (N_28666,N_27930,N_27782);
nand U28667 (N_28667,N_28020,N_28065);
nor U28668 (N_28668,N_28174,N_27657);
nor U28669 (N_28669,N_27776,N_27677);
and U28670 (N_28670,N_28147,N_27989);
or U28671 (N_28671,N_27703,N_28018);
nor U28672 (N_28672,N_27904,N_27910);
nor U28673 (N_28673,N_27732,N_27774);
or U28674 (N_28674,N_27611,N_27882);
or U28675 (N_28675,N_27701,N_28029);
nand U28676 (N_28676,N_27957,N_27750);
or U28677 (N_28677,N_28140,N_27971);
xnor U28678 (N_28678,N_27659,N_27984);
nand U28679 (N_28679,N_27817,N_28041);
nand U28680 (N_28680,N_27797,N_27698);
or U28681 (N_28681,N_27972,N_28117);
nand U28682 (N_28682,N_27841,N_27955);
nand U28683 (N_28683,N_28113,N_27954);
nand U28684 (N_28684,N_27956,N_27910);
nor U28685 (N_28685,N_28176,N_27967);
nor U28686 (N_28686,N_28116,N_27847);
nor U28687 (N_28687,N_28167,N_28100);
and U28688 (N_28688,N_27756,N_27913);
xor U28689 (N_28689,N_28057,N_27653);
xnor U28690 (N_28690,N_28118,N_28024);
and U28691 (N_28691,N_27717,N_27925);
xnor U28692 (N_28692,N_27683,N_27793);
or U28693 (N_28693,N_27994,N_28128);
xnor U28694 (N_28694,N_27912,N_28176);
and U28695 (N_28695,N_27749,N_28072);
and U28696 (N_28696,N_27979,N_28159);
xnor U28697 (N_28697,N_27876,N_27788);
nor U28698 (N_28698,N_27898,N_27964);
nor U28699 (N_28699,N_27870,N_27632);
xnor U28700 (N_28700,N_27721,N_27793);
xnor U28701 (N_28701,N_28015,N_27745);
nand U28702 (N_28702,N_28090,N_27772);
nor U28703 (N_28703,N_28143,N_27974);
and U28704 (N_28704,N_27820,N_27646);
nor U28705 (N_28705,N_27809,N_28031);
nor U28706 (N_28706,N_27648,N_27734);
or U28707 (N_28707,N_28193,N_28112);
or U28708 (N_28708,N_27957,N_27901);
or U28709 (N_28709,N_28095,N_28108);
or U28710 (N_28710,N_27794,N_28144);
nand U28711 (N_28711,N_27724,N_27686);
and U28712 (N_28712,N_27659,N_28129);
and U28713 (N_28713,N_27692,N_27650);
or U28714 (N_28714,N_27926,N_27609);
xor U28715 (N_28715,N_27826,N_27706);
nand U28716 (N_28716,N_28162,N_27901);
nand U28717 (N_28717,N_28080,N_27609);
nand U28718 (N_28718,N_27827,N_28199);
nand U28719 (N_28719,N_27923,N_27767);
nand U28720 (N_28720,N_28024,N_27713);
and U28721 (N_28721,N_27816,N_27734);
nor U28722 (N_28722,N_28081,N_27979);
nand U28723 (N_28723,N_27893,N_27622);
and U28724 (N_28724,N_27700,N_28002);
or U28725 (N_28725,N_28154,N_28014);
or U28726 (N_28726,N_28142,N_27676);
nand U28727 (N_28727,N_27982,N_27957);
nor U28728 (N_28728,N_27900,N_28121);
nand U28729 (N_28729,N_27859,N_27884);
nor U28730 (N_28730,N_27712,N_27983);
xor U28731 (N_28731,N_28153,N_27760);
and U28732 (N_28732,N_28120,N_28189);
nand U28733 (N_28733,N_27943,N_27801);
nand U28734 (N_28734,N_28021,N_27640);
xor U28735 (N_28735,N_28179,N_28175);
xor U28736 (N_28736,N_27794,N_27840);
nor U28737 (N_28737,N_27702,N_27730);
xnor U28738 (N_28738,N_27892,N_28055);
and U28739 (N_28739,N_27788,N_27855);
or U28740 (N_28740,N_27631,N_27866);
nand U28741 (N_28741,N_27891,N_27832);
and U28742 (N_28742,N_27618,N_27653);
nor U28743 (N_28743,N_28063,N_27729);
nand U28744 (N_28744,N_27737,N_28160);
nand U28745 (N_28745,N_27783,N_28067);
nand U28746 (N_28746,N_28055,N_28005);
and U28747 (N_28747,N_27758,N_28046);
or U28748 (N_28748,N_27664,N_28037);
nor U28749 (N_28749,N_28190,N_28092);
or U28750 (N_28750,N_28128,N_27628);
nand U28751 (N_28751,N_27852,N_27611);
and U28752 (N_28752,N_27635,N_28050);
or U28753 (N_28753,N_27999,N_27865);
and U28754 (N_28754,N_27667,N_27780);
nor U28755 (N_28755,N_28093,N_27912);
or U28756 (N_28756,N_27838,N_27848);
xor U28757 (N_28757,N_27735,N_28122);
and U28758 (N_28758,N_27864,N_27985);
or U28759 (N_28759,N_27998,N_28130);
nand U28760 (N_28760,N_28030,N_27832);
and U28761 (N_28761,N_27895,N_28045);
or U28762 (N_28762,N_27843,N_27777);
nor U28763 (N_28763,N_28006,N_27712);
and U28764 (N_28764,N_27750,N_27649);
and U28765 (N_28765,N_27865,N_27963);
nor U28766 (N_28766,N_27758,N_27738);
and U28767 (N_28767,N_27992,N_27871);
xnor U28768 (N_28768,N_28089,N_28006);
nand U28769 (N_28769,N_27695,N_27657);
nor U28770 (N_28770,N_27709,N_28126);
and U28771 (N_28771,N_27622,N_27642);
nand U28772 (N_28772,N_27688,N_28147);
nand U28773 (N_28773,N_28161,N_28067);
or U28774 (N_28774,N_28037,N_27756);
or U28775 (N_28775,N_27831,N_27811);
xor U28776 (N_28776,N_27890,N_28002);
or U28777 (N_28777,N_28031,N_28095);
nor U28778 (N_28778,N_27949,N_27829);
nand U28779 (N_28779,N_27708,N_28106);
nor U28780 (N_28780,N_27985,N_27822);
nor U28781 (N_28781,N_28084,N_27635);
and U28782 (N_28782,N_27698,N_28003);
nand U28783 (N_28783,N_27945,N_27807);
xnor U28784 (N_28784,N_27993,N_27842);
nor U28785 (N_28785,N_27867,N_28164);
nand U28786 (N_28786,N_27626,N_27691);
or U28787 (N_28787,N_28022,N_27737);
nand U28788 (N_28788,N_27966,N_27950);
or U28789 (N_28789,N_28137,N_28141);
and U28790 (N_28790,N_27796,N_27865);
and U28791 (N_28791,N_28012,N_27960);
or U28792 (N_28792,N_27685,N_27871);
nor U28793 (N_28793,N_27844,N_28034);
and U28794 (N_28794,N_28134,N_28172);
or U28795 (N_28795,N_27998,N_27717);
and U28796 (N_28796,N_28107,N_27944);
nor U28797 (N_28797,N_28074,N_27904);
nand U28798 (N_28798,N_27648,N_27859);
nand U28799 (N_28799,N_28061,N_27747);
and U28800 (N_28800,N_28488,N_28487);
xnor U28801 (N_28801,N_28740,N_28261);
nor U28802 (N_28802,N_28599,N_28737);
nand U28803 (N_28803,N_28424,N_28337);
xor U28804 (N_28804,N_28315,N_28712);
nor U28805 (N_28805,N_28210,N_28279);
and U28806 (N_28806,N_28778,N_28223);
nand U28807 (N_28807,N_28573,N_28426);
and U28808 (N_28808,N_28471,N_28722);
and U28809 (N_28809,N_28705,N_28207);
nand U28810 (N_28810,N_28431,N_28638);
nand U28811 (N_28811,N_28280,N_28365);
nor U28812 (N_28812,N_28792,N_28617);
nand U28813 (N_28813,N_28597,N_28661);
or U28814 (N_28814,N_28414,N_28626);
nand U28815 (N_28815,N_28662,N_28641);
xnor U28816 (N_28816,N_28554,N_28256);
or U28817 (N_28817,N_28672,N_28578);
xor U28818 (N_28818,N_28743,N_28797);
xor U28819 (N_28819,N_28413,N_28265);
or U28820 (N_28820,N_28621,N_28741);
and U28821 (N_28821,N_28404,N_28252);
nand U28822 (N_28822,N_28347,N_28395);
nor U28823 (N_28823,N_28273,N_28614);
nor U28824 (N_28824,N_28334,N_28313);
or U28825 (N_28825,N_28720,N_28222);
nand U28826 (N_28826,N_28217,N_28714);
nand U28827 (N_28827,N_28655,N_28540);
and U28828 (N_28828,N_28787,N_28284);
nor U28829 (N_28829,N_28507,N_28303);
nand U28830 (N_28830,N_28477,N_28220);
nand U28831 (N_28831,N_28519,N_28522);
nor U28832 (N_28832,N_28286,N_28482);
xor U28833 (N_28833,N_28494,N_28676);
nor U28834 (N_28834,N_28379,N_28200);
or U28835 (N_28835,N_28491,N_28232);
or U28836 (N_28836,N_28465,N_28373);
xnor U28837 (N_28837,N_28250,N_28683);
or U28838 (N_28838,N_28734,N_28736);
and U28839 (N_28839,N_28325,N_28633);
xor U28840 (N_28840,N_28764,N_28237);
and U28841 (N_28841,N_28715,N_28526);
or U28842 (N_28842,N_28654,N_28269);
xnor U28843 (N_28843,N_28464,N_28370);
xnor U28844 (N_28844,N_28306,N_28480);
nor U28845 (N_28845,N_28652,N_28650);
nand U28846 (N_28846,N_28777,N_28615);
nand U28847 (N_28847,N_28755,N_28326);
xnor U28848 (N_28848,N_28535,N_28374);
nor U28849 (N_28849,N_28710,N_28344);
nand U28850 (N_28850,N_28233,N_28455);
xor U28851 (N_28851,N_28361,N_28765);
nand U28852 (N_28852,N_28645,N_28475);
nand U28853 (N_28853,N_28368,N_28731);
nor U28854 (N_28854,N_28706,N_28257);
nor U28855 (N_28855,N_28267,N_28761);
or U28856 (N_28856,N_28212,N_28735);
xor U28857 (N_28857,N_28634,N_28419);
xnor U28858 (N_28858,N_28432,N_28446);
and U28859 (N_28859,N_28644,N_28205);
nor U28860 (N_28860,N_28673,N_28203);
or U28861 (N_28861,N_28605,N_28649);
and U28862 (N_28862,N_28226,N_28292);
and U28863 (N_28863,N_28301,N_28758);
nor U28864 (N_28864,N_28732,N_28651);
nand U28865 (N_28865,N_28609,N_28786);
xor U28866 (N_28866,N_28266,N_28505);
and U28867 (N_28867,N_28208,N_28391);
and U28868 (N_28868,N_28246,N_28678);
nor U28869 (N_28869,N_28434,N_28698);
xor U28870 (N_28870,N_28251,N_28752);
and U28871 (N_28871,N_28445,N_28760);
nor U28872 (N_28872,N_28383,N_28713);
xor U28873 (N_28873,N_28328,N_28601);
or U28874 (N_28874,N_28497,N_28674);
nor U28875 (N_28875,N_28243,N_28581);
or U28876 (N_28876,N_28729,N_28509);
nor U28877 (N_28877,N_28503,N_28369);
and U28878 (N_28878,N_28263,N_28433);
nor U28879 (N_28879,N_28305,N_28258);
or U28880 (N_28880,N_28213,N_28454);
nor U28881 (N_28881,N_28687,N_28282);
nor U28882 (N_28882,N_28612,N_28759);
or U28883 (N_28883,N_28556,N_28523);
xnor U28884 (N_28884,N_28401,N_28399);
nor U28885 (N_28885,N_28646,N_28441);
nor U28886 (N_28886,N_28500,N_28584);
xor U28887 (N_28887,N_28703,N_28783);
nand U28888 (N_28888,N_28773,N_28580);
nor U28889 (N_28889,N_28772,N_28570);
xnor U28890 (N_28890,N_28481,N_28398);
xnor U28891 (N_28891,N_28219,N_28402);
or U28892 (N_28892,N_28575,N_28657);
and U28893 (N_28893,N_28671,N_28312);
xor U28894 (N_28894,N_28274,N_28354);
xor U28895 (N_28895,N_28586,N_28459);
xor U28896 (N_28896,N_28460,N_28766);
xnor U28897 (N_28897,N_28541,N_28642);
xor U28898 (N_28898,N_28211,N_28474);
and U28899 (N_28899,N_28763,N_28538);
or U28900 (N_28900,N_28342,N_28501);
and U28901 (N_28901,N_28717,N_28422);
and U28902 (N_28902,N_28593,N_28287);
xnor U28903 (N_28903,N_28542,N_28744);
or U28904 (N_28904,N_28511,N_28602);
or U28905 (N_28905,N_28780,N_28725);
xor U28906 (N_28906,N_28793,N_28591);
nand U28907 (N_28907,N_28314,N_28553);
nand U28908 (N_28908,N_28566,N_28299);
xnor U28909 (N_28909,N_28545,N_28429);
xor U28910 (N_28910,N_28510,N_28204);
xor U28911 (N_28911,N_28206,N_28295);
nand U28912 (N_28912,N_28619,N_28468);
nand U28913 (N_28913,N_28360,N_28548);
nand U28914 (N_28914,N_28514,N_28667);
nand U28915 (N_28915,N_28704,N_28366);
or U28916 (N_28916,N_28298,N_28456);
xnor U28917 (N_28917,N_28533,N_28727);
xnor U28918 (N_28918,N_28589,N_28750);
xor U28919 (N_28919,N_28255,N_28606);
xnor U28920 (N_28920,N_28508,N_28592);
and U28921 (N_28921,N_28253,N_28427);
nor U28922 (N_28922,N_28322,N_28350);
xor U28923 (N_28923,N_28516,N_28358);
and U28924 (N_28924,N_28234,N_28636);
xnor U28925 (N_28925,N_28216,N_28559);
and U28926 (N_28926,N_28603,N_28600);
or U28927 (N_28927,N_28338,N_28558);
nor U28928 (N_28928,N_28699,N_28668);
and U28929 (N_28929,N_28331,N_28451);
or U28930 (N_28930,N_28393,N_28564);
nand U28931 (N_28931,N_28469,N_28259);
and U28932 (N_28932,N_28275,N_28447);
nand U28933 (N_28933,N_28290,N_28440);
nand U28934 (N_28934,N_28406,N_28675);
or U28935 (N_28935,N_28518,N_28659);
and U28936 (N_28936,N_28483,N_28453);
and U28937 (N_28937,N_28225,N_28768);
nand U28938 (N_28938,N_28215,N_28416);
nand U28939 (N_28939,N_28608,N_28539);
xnor U28940 (N_28940,N_28632,N_28774);
nor U28941 (N_28941,N_28635,N_28435);
xnor U28942 (N_28942,N_28392,N_28707);
or U28943 (N_28943,N_28376,N_28549);
nor U28944 (N_28944,N_28604,N_28719);
or U28945 (N_28945,N_28443,N_28670);
and U28946 (N_28946,N_28798,N_28472);
xor U28947 (N_28947,N_28214,N_28679);
or U28948 (N_28948,N_28385,N_28262);
and U28949 (N_28949,N_28630,N_28389);
xnor U28950 (N_28950,N_28270,N_28622);
nand U28951 (N_28951,N_28779,N_28775);
nand U28952 (N_28952,N_28228,N_28436);
nor U28953 (N_28953,N_28264,N_28583);
xor U28954 (N_28954,N_28639,N_28364);
and U28955 (N_28955,N_28420,N_28478);
and U28956 (N_28956,N_28562,N_28247);
nand U28957 (N_28957,N_28378,N_28276);
or U28958 (N_28958,N_28356,N_28297);
xor U28959 (N_28959,N_28470,N_28355);
and U28960 (N_28960,N_28277,N_28682);
xnor U28961 (N_28961,N_28283,N_28784);
nor U28962 (N_28962,N_28590,N_28485);
and U28963 (N_28963,N_28218,N_28400);
or U28964 (N_28964,N_28458,N_28618);
xnor U28965 (N_28965,N_28403,N_28330);
and U28966 (N_28966,N_28227,N_28528);
and U28967 (N_28967,N_28620,N_28669);
and U28968 (N_28968,N_28421,N_28439);
and U28969 (N_28969,N_28349,N_28319);
or U28970 (N_28970,N_28377,N_28348);
nor U28971 (N_28971,N_28332,N_28762);
nor U28972 (N_28972,N_28381,N_28690);
and U28973 (N_28973,N_28663,N_28310);
nand U28974 (N_28974,N_28346,N_28484);
nor U28975 (N_28975,N_28423,N_28723);
and U28976 (N_28976,N_28693,N_28757);
or U28977 (N_28977,N_28771,N_28448);
and U28978 (N_28978,N_28409,N_28788);
xnor U28979 (N_28979,N_28579,N_28656);
and U28980 (N_28980,N_28230,N_28231);
and U28981 (N_28981,N_28323,N_28437);
nand U28982 (N_28982,N_28515,N_28594);
or U28983 (N_28983,N_28708,N_28329);
nand U28984 (N_28984,N_28794,N_28340);
xor U28985 (N_28985,N_28799,N_28607);
and U28986 (N_28986,N_28335,N_28236);
nor U28987 (N_28987,N_28351,N_28397);
nor U28988 (N_28988,N_28689,N_28380);
and U28989 (N_28989,N_28680,N_28567);
nand U28990 (N_28990,N_28384,N_28492);
nor U28991 (N_28991,N_28685,N_28746);
nor U28992 (N_28992,N_28595,N_28316);
xor U28993 (N_28993,N_28749,N_28320);
xor U28994 (N_28994,N_28209,N_28665);
xnor U28995 (N_28995,N_28701,N_28544);
or U28996 (N_28996,N_28343,N_28653);
or U28997 (N_28997,N_28688,N_28718);
nor U28998 (N_28998,N_28572,N_28696);
or U28999 (N_28999,N_28307,N_28462);
nand U29000 (N_29000,N_28527,N_28624);
nor U29001 (N_29001,N_28547,N_28643);
nand U29002 (N_29002,N_28613,N_28795);
nand U29003 (N_29003,N_28463,N_28739);
and U29004 (N_29004,N_28697,N_28577);
nor U29005 (N_29005,N_28691,N_28382);
xnor U29006 (N_29006,N_28260,N_28493);
xnor U29007 (N_29007,N_28336,N_28353);
nand U29008 (N_29008,N_28410,N_28552);
or U29009 (N_29009,N_28551,N_28271);
or U29010 (N_29010,N_28640,N_28625);
nand U29011 (N_29011,N_28543,N_28311);
xnor U29012 (N_29012,N_28702,N_28244);
nor U29013 (N_29013,N_28733,N_28461);
and U29014 (N_29014,N_28333,N_28405);
nand U29015 (N_29015,N_28585,N_28476);
or U29016 (N_29016,N_28628,N_28411);
and U29017 (N_29017,N_28496,N_28321);
nor U29018 (N_29018,N_28300,N_28238);
xnor U29019 (N_29019,N_28756,N_28498);
xor U29020 (N_29020,N_28202,N_28425);
and U29021 (N_29021,N_28466,N_28647);
or U29022 (N_29022,N_28695,N_28317);
or U29023 (N_29023,N_28318,N_28711);
or U29024 (N_29024,N_28293,N_28700);
nor U29025 (N_29025,N_28588,N_28367);
and U29026 (N_29026,N_28534,N_28686);
or U29027 (N_29027,N_28524,N_28388);
and U29028 (N_29028,N_28569,N_28596);
nand U29029 (N_29029,N_28561,N_28249);
xnor U29030 (N_29030,N_28289,N_28692);
and U29031 (N_29031,N_28296,N_28637);
nor U29032 (N_29032,N_28240,N_28684);
nor U29033 (N_29033,N_28531,N_28776);
or U29034 (N_29034,N_28574,N_28417);
nand U29035 (N_29035,N_28372,N_28341);
or U29036 (N_29036,N_28537,N_28489);
xnor U29037 (N_29037,N_28563,N_28576);
nor U29038 (N_29038,N_28648,N_28789);
nand U29039 (N_29039,N_28753,N_28241);
or U29040 (N_29040,N_28235,N_28560);
xor U29041 (N_29041,N_28442,N_28694);
xnor U29042 (N_29042,N_28291,N_28504);
xor U29043 (N_29043,N_28598,N_28473);
nor U29044 (N_29044,N_28610,N_28408);
nor U29045 (N_29045,N_28288,N_28302);
nor U29046 (N_29046,N_28502,N_28754);
and U29047 (N_29047,N_28728,N_28285);
or U29048 (N_29048,N_28221,N_28529);
nand U29049 (N_29049,N_28239,N_28677);
nand U29050 (N_29050,N_28742,N_28242);
and U29051 (N_29051,N_28345,N_28525);
xnor U29052 (N_29052,N_28546,N_28745);
or U29053 (N_29053,N_28412,N_28769);
xor U29054 (N_29054,N_28357,N_28664);
xnor U29055 (N_29055,N_28294,N_28438);
nand U29056 (N_29056,N_28430,N_28582);
xnor U29057 (N_29057,N_28730,N_28272);
xnor U29058 (N_29058,N_28520,N_28738);
nor U29059 (N_29059,N_28629,N_28536);
nor U29060 (N_29060,N_28268,N_28248);
or U29061 (N_29061,N_28428,N_28791);
xor U29062 (N_29062,N_28748,N_28362);
or U29063 (N_29063,N_28751,N_28394);
nand U29064 (N_29064,N_28517,N_28532);
or U29065 (N_29065,N_28201,N_28452);
nor U29066 (N_29066,N_28587,N_28390);
and U29067 (N_29067,N_28375,N_28339);
or U29068 (N_29068,N_28631,N_28681);
nand U29069 (N_29069,N_28709,N_28721);
and U29070 (N_29070,N_28716,N_28512);
nor U29071 (N_29071,N_28555,N_28506);
nor U29072 (N_29072,N_28568,N_28571);
xnor U29073 (N_29073,N_28324,N_28415);
and U29074 (N_29074,N_28363,N_28309);
nor U29075 (N_29075,N_28418,N_28490);
xor U29076 (N_29076,N_28495,N_28747);
nor U29077 (N_29077,N_28660,N_28499);
nor U29078 (N_29078,N_28450,N_28229);
or U29079 (N_29079,N_28449,N_28359);
nor U29080 (N_29080,N_28616,N_28224);
and U29081 (N_29081,N_28611,N_28386);
xor U29082 (N_29082,N_28726,N_28770);
nand U29083 (N_29083,N_28457,N_28782);
xor U29084 (N_29084,N_28781,N_28352);
nor U29085 (N_29085,N_28530,N_28565);
nand U29086 (N_29086,N_28557,N_28521);
and U29087 (N_29087,N_28623,N_28281);
and U29088 (N_29088,N_28790,N_28245);
nor U29089 (N_29089,N_28327,N_28396);
nor U29090 (N_29090,N_28785,N_28387);
nand U29091 (N_29091,N_28278,N_28796);
xnor U29092 (N_29092,N_28658,N_28467);
nor U29093 (N_29093,N_28254,N_28486);
and U29094 (N_29094,N_28513,N_28627);
nor U29095 (N_29095,N_28666,N_28444);
and U29096 (N_29096,N_28371,N_28304);
nand U29097 (N_29097,N_28724,N_28550);
and U29098 (N_29098,N_28479,N_28767);
xnor U29099 (N_29099,N_28308,N_28407);
nand U29100 (N_29100,N_28532,N_28456);
nor U29101 (N_29101,N_28347,N_28274);
xnor U29102 (N_29102,N_28739,N_28258);
nand U29103 (N_29103,N_28620,N_28663);
nand U29104 (N_29104,N_28232,N_28550);
or U29105 (N_29105,N_28599,N_28781);
nand U29106 (N_29106,N_28463,N_28573);
nand U29107 (N_29107,N_28567,N_28248);
nor U29108 (N_29108,N_28316,N_28322);
nand U29109 (N_29109,N_28584,N_28662);
nand U29110 (N_29110,N_28566,N_28370);
nand U29111 (N_29111,N_28694,N_28468);
nor U29112 (N_29112,N_28264,N_28537);
or U29113 (N_29113,N_28311,N_28377);
xnor U29114 (N_29114,N_28617,N_28471);
and U29115 (N_29115,N_28275,N_28238);
or U29116 (N_29116,N_28798,N_28274);
or U29117 (N_29117,N_28445,N_28378);
nand U29118 (N_29118,N_28785,N_28546);
or U29119 (N_29119,N_28450,N_28408);
nor U29120 (N_29120,N_28726,N_28203);
or U29121 (N_29121,N_28753,N_28215);
or U29122 (N_29122,N_28717,N_28386);
and U29123 (N_29123,N_28427,N_28655);
nand U29124 (N_29124,N_28444,N_28429);
or U29125 (N_29125,N_28458,N_28793);
nor U29126 (N_29126,N_28259,N_28296);
or U29127 (N_29127,N_28530,N_28254);
and U29128 (N_29128,N_28300,N_28558);
nand U29129 (N_29129,N_28465,N_28473);
nand U29130 (N_29130,N_28489,N_28510);
and U29131 (N_29131,N_28543,N_28723);
and U29132 (N_29132,N_28435,N_28754);
and U29133 (N_29133,N_28251,N_28755);
and U29134 (N_29134,N_28665,N_28502);
or U29135 (N_29135,N_28655,N_28625);
nand U29136 (N_29136,N_28528,N_28641);
xnor U29137 (N_29137,N_28676,N_28765);
and U29138 (N_29138,N_28343,N_28496);
xnor U29139 (N_29139,N_28449,N_28546);
xor U29140 (N_29140,N_28398,N_28724);
nor U29141 (N_29141,N_28268,N_28460);
nand U29142 (N_29142,N_28457,N_28203);
nand U29143 (N_29143,N_28734,N_28689);
and U29144 (N_29144,N_28651,N_28791);
and U29145 (N_29145,N_28695,N_28771);
xor U29146 (N_29146,N_28228,N_28255);
or U29147 (N_29147,N_28268,N_28528);
nand U29148 (N_29148,N_28369,N_28257);
xor U29149 (N_29149,N_28470,N_28740);
xnor U29150 (N_29150,N_28318,N_28452);
xnor U29151 (N_29151,N_28252,N_28769);
or U29152 (N_29152,N_28642,N_28206);
xor U29153 (N_29153,N_28373,N_28549);
nand U29154 (N_29154,N_28438,N_28293);
xnor U29155 (N_29155,N_28560,N_28251);
nand U29156 (N_29156,N_28744,N_28342);
or U29157 (N_29157,N_28554,N_28562);
nand U29158 (N_29158,N_28407,N_28641);
nand U29159 (N_29159,N_28781,N_28592);
nand U29160 (N_29160,N_28781,N_28261);
and U29161 (N_29161,N_28609,N_28455);
or U29162 (N_29162,N_28628,N_28490);
nand U29163 (N_29163,N_28734,N_28531);
and U29164 (N_29164,N_28441,N_28457);
nor U29165 (N_29165,N_28525,N_28758);
nand U29166 (N_29166,N_28684,N_28429);
nand U29167 (N_29167,N_28470,N_28315);
or U29168 (N_29168,N_28549,N_28305);
xor U29169 (N_29169,N_28621,N_28379);
xor U29170 (N_29170,N_28706,N_28475);
nor U29171 (N_29171,N_28328,N_28398);
nor U29172 (N_29172,N_28253,N_28718);
nand U29173 (N_29173,N_28667,N_28479);
or U29174 (N_29174,N_28483,N_28336);
nor U29175 (N_29175,N_28267,N_28759);
and U29176 (N_29176,N_28545,N_28550);
nor U29177 (N_29177,N_28399,N_28700);
and U29178 (N_29178,N_28687,N_28445);
nand U29179 (N_29179,N_28422,N_28678);
or U29180 (N_29180,N_28761,N_28608);
nand U29181 (N_29181,N_28232,N_28681);
xnor U29182 (N_29182,N_28415,N_28396);
and U29183 (N_29183,N_28707,N_28582);
or U29184 (N_29184,N_28323,N_28730);
nand U29185 (N_29185,N_28321,N_28459);
or U29186 (N_29186,N_28736,N_28683);
and U29187 (N_29187,N_28350,N_28415);
nor U29188 (N_29188,N_28508,N_28774);
or U29189 (N_29189,N_28256,N_28504);
nand U29190 (N_29190,N_28330,N_28373);
nand U29191 (N_29191,N_28343,N_28372);
xor U29192 (N_29192,N_28464,N_28706);
nor U29193 (N_29193,N_28754,N_28586);
and U29194 (N_29194,N_28695,N_28790);
and U29195 (N_29195,N_28460,N_28390);
or U29196 (N_29196,N_28512,N_28439);
nand U29197 (N_29197,N_28403,N_28617);
nand U29198 (N_29198,N_28603,N_28681);
or U29199 (N_29199,N_28513,N_28465);
and U29200 (N_29200,N_28499,N_28729);
xor U29201 (N_29201,N_28698,N_28242);
xnor U29202 (N_29202,N_28231,N_28491);
and U29203 (N_29203,N_28795,N_28735);
and U29204 (N_29204,N_28269,N_28704);
nor U29205 (N_29205,N_28783,N_28309);
xnor U29206 (N_29206,N_28333,N_28767);
xor U29207 (N_29207,N_28398,N_28508);
xnor U29208 (N_29208,N_28258,N_28566);
nor U29209 (N_29209,N_28410,N_28268);
xor U29210 (N_29210,N_28639,N_28347);
nand U29211 (N_29211,N_28344,N_28283);
nand U29212 (N_29212,N_28668,N_28277);
nand U29213 (N_29213,N_28232,N_28362);
xor U29214 (N_29214,N_28585,N_28204);
or U29215 (N_29215,N_28395,N_28294);
or U29216 (N_29216,N_28779,N_28409);
or U29217 (N_29217,N_28547,N_28478);
nand U29218 (N_29218,N_28498,N_28345);
or U29219 (N_29219,N_28661,N_28269);
or U29220 (N_29220,N_28397,N_28331);
or U29221 (N_29221,N_28234,N_28618);
and U29222 (N_29222,N_28567,N_28433);
or U29223 (N_29223,N_28268,N_28352);
xor U29224 (N_29224,N_28636,N_28653);
and U29225 (N_29225,N_28256,N_28321);
or U29226 (N_29226,N_28453,N_28223);
or U29227 (N_29227,N_28245,N_28682);
nor U29228 (N_29228,N_28738,N_28321);
or U29229 (N_29229,N_28293,N_28569);
xor U29230 (N_29230,N_28607,N_28349);
xnor U29231 (N_29231,N_28303,N_28361);
xor U29232 (N_29232,N_28778,N_28251);
or U29233 (N_29233,N_28541,N_28746);
or U29234 (N_29234,N_28722,N_28448);
and U29235 (N_29235,N_28484,N_28403);
nand U29236 (N_29236,N_28464,N_28248);
and U29237 (N_29237,N_28612,N_28408);
xnor U29238 (N_29238,N_28463,N_28506);
and U29239 (N_29239,N_28505,N_28584);
xor U29240 (N_29240,N_28706,N_28329);
nand U29241 (N_29241,N_28214,N_28497);
or U29242 (N_29242,N_28248,N_28398);
xnor U29243 (N_29243,N_28787,N_28653);
xnor U29244 (N_29244,N_28296,N_28613);
or U29245 (N_29245,N_28610,N_28529);
or U29246 (N_29246,N_28706,N_28388);
nand U29247 (N_29247,N_28429,N_28287);
nand U29248 (N_29248,N_28743,N_28236);
and U29249 (N_29249,N_28772,N_28579);
or U29250 (N_29250,N_28746,N_28394);
or U29251 (N_29251,N_28353,N_28708);
xnor U29252 (N_29252,N_28507,N_28786);
or U29253 (N_29253,N_28537,N_28743);
and U29254 (N_29254,N_28214,N_28237);
or U29255 (N_29255,N_28232,N_28332);
xnor U29256 (N_29256,N_28313,N_28294);
nand U29257 (N_29257,N_28721,N_28647);
and U29258 (N_29258,N_28217,N_28708);
nand U29259 (N_29259,N_28660,N_28567);
nor U29260 (N_29260,N_28743,N_28302);
nor U29261 (N_29261,N_28586,N_28404);
xor U29262 (N_29262,N_28506,N_28348);
and U29263 (N_29263,N_28226,N_28332);
or U29264 (N_29264,N_28384,N_28559);
xor U29265 (N_29265,N_28711,N_28570);
or U29266 (N_29266,N_28263,N_28342);
or U29267 (N_29267,N_28200,N_28734);
nor U29268 (N_29268,N_28348,N_28399);
and U29269 (N_29269,N_28344,N_28382);
or U29270 (N_29270,N_28515,N_28236);
nand U29271 (N_29271,N_28708,N_28300);
nor U29272 (N_29272,N_28688,N_28454);
nand U29273 (N_29273,N_28461,N_28225);
xor U29274 (N_29274,N_28774,N_28717);
or U29275 (N_29275,N_28251,N_28703);
xnor U29276 (N_29276,N_28365,N_28665);
nand U29277 (N_29277,N_28795,N_28299);
or U29278 (N_29278,N_28415,N_28708);
or U29279 (N_29279,N_28291,N_28481);
nand U29280 (N_29280,N_28654,N_28246);
nand U29281 (N_29281,N_28710,N_28392);
nor U29282 (N_29282,N_28357,N_28442);
or U29283 (N_29283,N_28626,N_28778);
nand U29284 (N_29284,N_28537,N_28650);
nand U29285 (N_29285,N_28371,N_28357);
and U29286 (N_29286,N_28730,N_28213);
and U29287 (N_29287,N_28638,N_28282);
xor U29288 (N_29288,N_28593,N_28292);
or U29289 (N_29289,N_28542,N_28601);
or U29290 (N_29290,N_28402,N_28561);
nor U29291 (N_29291,N_28533,N_28514);
nand U29292 (N_29292,N_28529,N_28469);
and U29293 (N_29293,N_28735,N_28433);
xor U29294 (N_29294,N_28783,N_28272);
nand U29295 (N_29295,N_28522,N_28257);
and U29296 (N_29296,N_28714,N_28378);
nor U29297 (N_29297,N_28306,N_28254);
nor U29298 (N_29298,N_28591,N_28293);
nor U29299 (N_29299,N_28417,N_28241);
or U29300 (N_29300,N_28471,N_28774);
or U29301 (N_29301,N_28756,N_28240);
xor U29302 (N_29302,N_28645,N_28419);
xnor U29303 (N_29303,N_28668,N_28565);
xor U29304 (N_29304,N_28248,N_28560);
and U29305 (N_29305,N_28527,N_28744);
xnor U29306 (N_29306,N_28436,N_28759);
or U29307 (N_29307,N_28638,N_28777);
xnor U29308 (N_29308,N_28542,N_28694);
or U29309 (N_29309,N_28673,N_28380);
or U29310 (N_29310,N_28402,N_28232);
or U29311 (N_29311,N_28467,N_28519);
nor U29312 (N_29312,N_28289,N_28673);
xor U29313 (N_29313,N_28648,N_28300);
xor U29314 (N_29314,N_28779,N_28232);
and U29315 (N_29315,N_28524,N_28576);
and U29316 (N_29316,N_28397,N_28733);
nand U29317 (N_29317,N_28777,N_28244);
nor U29318 (N_29318,N_28294,N_28222);
xor U29319 (N_29319,N_28221,N_28719);
nand U29320 (N_29320,N_28228,N_28262);
nor U29321 (N_29321,N_28227,N_28761);
nor U29322 (N_29322,N_28347,N_28773);
or U29323 (N_29323,N_28463,N_28732);
or U29324 (N_29324,N_28432,N_28319);
or U29325 (N_29325,N_28547,N_28493);
and U29326 (N_29326,N_28723,N_28530);
and U29327 (N_29327,N_28784,N_28289);
and U29328 (N_29328,N_28720,N_28674);
and U29329 (N_29329,N_28416,N_28783);
nand U29330 (N_29330,N_28384,N_28529);
nor U29331 (N_29331,N_28424,N_28726);
nor U29332 (N_29332,N_28561,N_28538);
and U29333 (N_29333,N_28286,N_28640);
xnor U29334 (N_29334,N_28481,N_28634);
nand U29335 (N_29335,N_28481,N_28477);
xor U29336 (N_29336,N_28696,N_28255);
xnor U29337 (N_29337,N_28360,N_28525);
nor U29338 (N_29338,N_28523,N_28504);
nor U29339 (N_29339,N_28326,N_28588);
and U29340 (N_29340,N_28524,N_28789);
and U29341 (N_29341,N_28585,N_28716);
nand U29342 (N_29342,N_28351,N_28587);
or U29343 (N_29343,N_28208,N_28370);
xnor U29344 (N_29344,N_28513,N_28466);
nor U29345 (N_29345,N_28364,N_28501);
and U29346 (N_29346,N_28724,N_28596);
and U29347 (N_29347,N_28589,N_28707);
xor U29348 (N_29348,N_28411,N_28226);
or U29349 (N_29349,N_28509,N_28470);
xnor U29350 (N_29350,N_28759,N_28456);
and U29351 (N_29351,N_28608,N_28468);
xor U29352 (N_29352,N_28488,N_28474);
nor U29353 (N_29353,N_28343,N_28237);
xor U29354 (N_29354,N_28659,N_28232);
or U29355 (N_29355,N_28726,N_28783);
or U29356 (N_29356,N_28321,N_28397);
and U29357 (N_29357,N_28403,N_28236);
nand U29358 (N_29358,N_28759,N_28535);
nor U29359 (N_29359,N_28451,N_28637);
xor U29360 (N_29360,N_28578,N_28444);
nand U29361 (N_29361,N_28397,N_28572);
nor U29362 (N_29362,N_28393,N_28260);
xnor U29363 (N_29363,N_28415,N_28494);
xnor U29364 (N_29364,N_28649,N_28563);
xor U29365 (N_29365,N_28630,N_28601);
nand U29366 (N_29366,N_28465,N_28580);
nand U29367 (N_29367,N_28288,N_28201);
and U29368 (N_29368,N_28793,N_28688);
or U29369 (N_29369,N_28525,N_28208);
xnor U29370 (N_29370,N_28509,N_28382);
nand U29371 (N_29371,N_28543,N_28481);
nor U29372 (N_29372,N_28621,N_28243);
or U29373 (N_29373,N_28718,N_28290);
xor U29374 (N_29374,N_28630,N_28576);
and U29375 (N_29375,N_28371,N_28595);
or U29376 (N_29376,N_28694,N_28383);
or U29377 (N_29377,N_28312,N_28771);
nand U29378 (N_29378,N_28621,N_28668);
nor U29379 (N_29379,N_28592,N_28505);
xnor U29380 (N_29380,N_28258,N_28699);
and U29381 (N_29381,N_28334,N_28225);
nand U29382 (N_29382,N_28758,N_28732);
xor U29383 (N_29383,N_28672,N_28250);
and U29384 (N_29384,N_28210,N_28703);
and U29385 (N_29385,N_28203,N_28661);
nand U29386 (N_29386,N_28773,N_28324);
and U29387 (N_29387,N_28670,N_28404);
and U29388 (N_29388,N_28748,N_28406);
xor U29389 (N_29389,N_28585,N_28250);
and U29390 (N_29390,N_28338,N_28219);
nor U29391 (N_29391,N_28451,N_28381);
or U29392 (N_29392,N_28500,N_28275);
nor U29393 (N_29393,N_28487,N_28332);
nand U29394 (N_29394,N_28686,N_28309);
and U29395 (N_29395,N_28540,N_28788);
and U29396 (N_29396,N_28596,N_28497);
or U29397 (N_29397,N_28251,N_28632);
nor U29398 (N_29398,N_28706,N_28339);
nor U29399 (N_29399,N_28494,N_28506);
nand U29400 (N_29400,N_29266,N_28938);
xnor U29401 (N_29401,N_28986,N_29190);
and U29402 (N_29402,N_28931,N_29146);
xnor U29403 (N_29403,N_29366,N_29149);
nor U29404 (N_29404,N_29013,N_29303);
and U29405 (N_29405,N_29377,N_28858);
xnor U29406 (N_29406,N_29359,N_29219);
nand U29407 (N_29407,N_29070,N_28823);
xor U29408 (N_29408,N_29282,N_29069);
xnor U29409 (N_29409,N_29179,N_28946);
or U29410 (N_29410,N_29301,N_29187);
and U29411 (N_29411,N_29031,N_29376);
nor U29412 (N_29412,N_28884,N_28876);
xnor U29413 (N_29413,N_29135,N_29308);
or U29414 (N_29414,N_28817,N_28837);
nor U29415 (N_29415,N_29141,N_28965);
xnor U29416 (N_29416,N_29169,N_28933);
nand U29417 (N_29417,N_29261,N_28936);
nand U29418 (N_29418,N_28802,N_29383);
xnor U29419 (N_29419,N_29089,N_29192);
and U29420 (N_29420,N_28958,N_29307);
or U29421 (N_29421,N_29157,N_29051);
and U29422 (N_29422,N_29207,N_29355);
or U29423 (N_29423,N_29127,N_29033);
and U29424 (N_29424,N_29218,N_29072);
xnor U29425 (N_29425,N_29114,N_29351);
and U29426 (N_29426,N_29185,N_28840);
nand U29427 (N_29427,N_29058,N_29107);
or U29428 (N_29428,N_29319,N_28810);
or U29429 (N_29429,N_29059,N_29382);
nand U29430 (N_29430,N_29224,N_28914);
nand U29431 (N_29431,N_29186,N_28964);
nand U29432 (N_29432,N_28897,N_28870);
nand U29433 (N_29433,N_28902,N_29133);
and U29434 (N_29434,N_29361,N_29164);
xnor U29435 (N_29435,N_28970,N_29317);
nor U29436 (N_29436,N_28832,N_28932);
and U29437 (N_29437,N_29309,N_29021);
or U29438 (N_29438,N_28906,N_28918);
xnor U29439 (N_29439,N_29145,N_29083);
nand U29440 (N_29440,N_29387,N_28903);
or U29441 (N_29441,N_29291,N_29123);
and U29442 (N_29442,N_28998,N_29062);
nor U29443 (N_29443,N_29230,N_28819);
nor U29444 (N_29444,N_29060,N_29269);
nor U29445 (N_29445,N_28816,N_29106);
nand U29446 (N_29446,N_29209,N_29128);
xor U29447 (N_29447,N_29144,N_28989);
nand U29448 (N_29448,N_29158,N_28907);
xnor U29449 (N_29449,N_29053,N_29182);
or U29450 (N_29450,N_29028,N_28800);
and U29451 (N_29451,N_28934,N_29034);
nand U29452 (N_29452,N_28821,N_29203);
xor U29453 (N_29453,N_29322,N_29332);
or U29454 (N_29454,N_29241,N_29094);
nand U29455 (N_29455,N_29140,N_29205);
nor U29456 (N_29456,N_29167,N_29172);
xnor U29457 (N_29457,N_28867,N_29109);
nand U29458 (N_29458,N_29280,N_28888);
nor U29459 (N_29459,N_29002,N_28893);
or U29460 (N_29460,N_29281,N_28868);
nand U29461 (N_29461,N_29392,N_29258);
nand U29462 (N_29462,N_29288,N_29386);
xor U29463 (N_29463,N_28953,N_29314);
or U29464 (N_29464,N_29056,N_28959);
and U29465 (N_29465,N_28904,N_29330);
or U29466 (N_29466,N_29357,N_28997);
xnor U29467 (N_29467,N_29247,N_29170);
nand U29468 (N_29468,N_29206,N_29321);
and U29469 (N_29469,N_29349,N_29183);
nor U29470 (N_29470,N_29102,N_29029);
nand U29471 (N_29471,N_28864,N_29112);
xnor U29472 (N_29472,N_28987,N_29333);
nor U29473 (N_29473,N_29380,N_29155);
and U29474 (N_29474,N_29043,N_29381);
and U29475 (N_29475,N_29299,N_28916);
nand U29476 (N_29476,N_28886,N_29120);
nand U29477 (N_29477,N_29345,N_28852);
or U29478 (N_29478,N_28833,N_29016);
and U29479 (N_29479,N_29079,N_29339);
nor U29480 (N_29480,N_28982,N_29335);
nor U29481 (N_29481,N_29118,N_29091);
or U29482 (N_29482,N_28996,N_28841);
or U29483 (N_29483,N_29006,N_28882);
nor U29484 (N_29484,N_29037,N_28863);
nand U29485 (N_29485,N_28928,N_29389);
xnor U29486 (N_29486,N_29244,N_28815);
nor U29487 (N_29487,N_28818,N_28873);
nor U29488 (N_29488,N_29151,N_28855);
or U29489 (N_29489,N_29344,N_29156);
and U29490 (N_29490,N_28900,N_28935);
or U29491 (N_29491,N_28875,N_29154);
nor U29492 (N_29492,N_28944,N_29071);
or U29493 (N_29493,N_29347,N_28920);
or U29494 (N_29494,N_29255,N_28968);
nand U29495 (N_29495,N_29180,N_28973);
nand U29496 (N_29496,N_28957,N_28985);
xnor U29497 (N_29497,N_29320,N_29152);
nand U29498 (N_29498,N_29289,N_29220);
nand U29499 (N_29499,N_29372,N_28850);
and U29500 (N_29500,N_29023,N_29108);
or U29501 (N_29501,N_29295,N_29188);
or U29502 (N_29502,N_29136,N_29310);
and U29503 (N_29503,N_29325,N_29286);
or U29504 (N_29504,N_29081,N_28809);
nand U29505 (N_29505,N_29005,N_28811);
nand U29506 (N_29506,N_29117,N_29181);
xnor U29507 (N_29507,N_29017,N_28942);
or U29508 (N_29508,N_28895,N_29040);
and U29509 (N_29509,N_28877,N_29233);
or U29510 (N_29510,N_29101,N_28801);
nor U29511 (N_29511,N_29012,N_29022);
nand U29512 (N_29512,N_29270,N_28930);
and U29513 (N_29513,N_28859,N_29068);
and U29514 (N_29514,N_28862,N_29126);
xnor U29515 (N_29515,N_29027,N_29358);
or U29516 (N_29516,N_29175,N_28826);
or U29517 (N_29517,N_29313,N_29393);
nor U29518 (N_29518,N_29371,N_29103);
nor U29519 (N_29519,N_29098,N_28993);
or U29520 (N_29520,N_29009,N_29085);
and U29521 (N_29521,N_29257,N_29001);
nand U29522 (N_29522,N_29353,N_28937);
nor U29523 (N_29523,N_29049,N_29113);
nand U29524 (N_29524,N_29138,N_29163);
xnor U29525 (N_29525,N_29297,N_28827);
nor U29526 (N_29526,N_29331,N_28943);
and U29527 (N_29527,N_28979,N_29150);
nand U29528 (N_29528,N_29214,N_29131);
or U29529 (N_29529,N_29076,N_29337);
nor U29530 (N_29530,N_29395,N_28908);
or U29531 (N_29531,N_28890,N_29160);
nand U29532 (N_29532,N_29242,N_29227);
nand U29533 (N_29533,N_29394,N_28865);
nor U29534 (N_29534,N_29055,N_28950);
nor U29535 (N_29535,N_29115,N_29239);
xnor U29536 (N_29536,N_29318,N_28869);
xnor U29537 (N_29537,N_29035,N_29228);
nor U29538 (N_29538,N_28971,N_29057);
nor U29539 (N_29539,N_29153,N_29193);
nand U29540 (N_29540,N_28824,N_29204);
and U29541 (N_29541,N_29132,N_29080);
or U29542 (N_29542,N_29119,N_28912);
xnor U29543 (N_29543,N_28836,N_29396);
nand U29544 (N_29544,N_29334,N_29041);
or U29545 (N_29545,N_28854,N_28975);
nor U29546 (N_29546,N_28804,N_29277);
nor U29547 (N_29547,N_29147,N_29312);
xnor U29548 (N_29548,N_29077,N_29348);
and U29549 (N_29549,N_29054,N_29370);
nor U29550 (N_29550,N_28992,N_28844);
xnor U29551 (N_29551,N_28891,N_29061);
nand U29552 (N_29552,N_28919,N_28806);
or U29553 (N_29553,N_28961,N_29238);
nand U29554 (N_29554,N_29384,N_29173);
nand U29555 (N_29555,N_29178,N_29200);
nand U29556 (N_29556,N_28954,N_29326);
xnor U29557 (N_29557,N_29195,N_29003);
nand U29558 (N_29558,N_28874,N_29336);
and U29559 (N_29559,N_28846,N_28960);
xor U29560 (N_29560,N_29290,N_29196);
nor U29561 (N_29561,N_28813,N_29036);
nand U29562 (N_29562,N_29082,N_28842);
and U29563 (N_29563,N_29311,N_29391);
nand U29564 (N_29564,N_28917,N_29217);
xor U29565 (N_29565,N_29298,N_29011);
nand U29566 (N_29566,N_29018,N_28939);
and U29567 (N_29567,N_29231,N_29341);
nor U29568 (N_29568,N_29189,N_29398);
nand U29569 (N_29569,N_28962,N_29092);
xor U29570 (N_29570,N_28983,N_28981);
xnor U29571 (N_29571,N_28848,N_29329);
nand U29572 (N_29572,N_29294,N_29168);
nor U29573 (N_29573,N_28845,N_28927);
xnor U29574 (N_29574,N_29385,N_28856);
nor U29575 (N_29575,N_29137,N_28872);
nand U29576 (N_29576,N_29240,N_28892);
and U29577 (N_29577,N_29216,N_28999);
xor U29578 (N_29578,N_29095,N_29225);
xor U29579 (N_29579,N_29259,N_28948);
nand U29580 (N_29580,N_28807,N_28911);
or U29581 (N_29581,N_29143,N_29315);
and U29582 (N_29582,N_29256,N_29350);
nor U29583 (N_29583,N_29300,N_28988);
or U29584 (N_29584,N_29197,N_28835);
xor U29585 (N_29585,N_29399,N_29226);
and U29586 (N_29586,N_29379,N_28820);
nor U29587 (N_29587,N_29279,N_29050);
xnor U29588 (N_29588,N_28922,N_29161);
nand U29589 (N_29589,N_29296,N_29222);
or U29590 (N_29590,N_28866,N_29162);
xnor U29591 (N_29591,N_28838,N_29174);
nor U29592 (N_29592,N_29073,N_29020);
or U29593 (N_29593,N_28966,N_29210);
xnor U29594 (N_29594,N_29248,N_28969);
and U29595 (N_29595,N_29087,N_29356);
or U29596 (N_29596,N_28945,N_29262);
nor U29597 (N_29597,N_29229,N_29304);
or U29598 (N_29598,N_28977,N_28913);
or U29599 (N_29599,N_29202,N_29323);
and U29600 (N_29600,N_29124,N_29265);
nor U29601 (N_29601,N_28926,N_29007);
nand U29602 (N_29602,N_29096,N_29032);
nand U29603 (N_29603,N_29075,N_29283);
nand U29604 (N_29604,N_29369,N_28896);
xor U29605 (N_29605,N_28881,N_29139);
nor U29606 (N_29606,N_29268,N_29374);
or U29607 (N_29607,N_28857,N_29285);
xor U29608 (N_29608,N_28830,N_29198);
nor U29609 (N_29609,N_29078,N_28929);
nand U29610 (N_29610,N_28851,N_29234);
and U29611 (N_29611,N_29273,N_29275);
xnor U29612 (N_29612,N_28828,N_29360);
and U29613 (N_29613,N_29246,N_29191);
or U29614 (N_29614,N_28825,N_29252);
and U29615 (N_29615,N_28905,N_28853);
nand U29616 (N_29616,N_28990,N_28843);
nand U29617 (N_29617,N_29039,N_29024);
nand U29618 (N_29618,N_28974,N_28963);
xor U29619 (N_29619,N_29338,N_29166);
xnor U29620 (N_29620,N_28839,N_28861);
nand U29621 (N_29621,N_29368,N_29271);
nor U29622 (N_29622,N_29327,N_29272);
nand U29623 (N_29623,N_29110,N_29223);
xnor U29624 (N_29624,N_29159,N_29354);
or U29625 (N_29625,N_29088,N_28940);
nand U29626 (N_29626,N_29121,N_28814);
nand U29627 (N_29627,N_29194,N_29042);
nand U29628 (N_29628,N_29184,N_28822);
and U29629 (N_29629,N_29276,N_29074);
and U29630 (N_29630,N_29253,N_29293);
or U29631 (N_29631,N_28967,N_29104);
or U29632 (N_29632,N_29008,N_29397);
or U29633 (N_29633,N_29045,N_29364);
or U29634 (N_29634,N_28994,N_29343);
and U29635 (N_29635,N_29235,N_29105);
nor U29636 (N_29636,N_29260,N_29044);
and U29637 (N_29637,N_29199,N_28951);
or U29638 (N_29638,N_28991,N_29000);
xnor U29639 (N_29639,N_28923,N_28978);
nor U29640 (N_29640,N_29211,N_29052);
or U29641 (N_29641,N_29065,N_28910);
nand U29642 (N_29642,N_29264,N_29236);
or U29643 (N_29643,N_29324,N_29030);
nand U29644 (N_29644,N_29362,N_29086);
and U29645 (N_29645,N_28878,N_28956);
nand U29646 (N_29646,N_29090,N_29352);
and U29647 (N_29647,N_29004,N_29026);
nand U29648 (N_29648,N_28955,N_29249);
nand U29649 (N_29649,N_28921,N_28909);
xor U29650 (N_29650,N_28901,N_29063);
and U29651 (N_29651,N_29038,N_29373);
nor U29652 (N_29652,N_29213,N_29284);
nand U29653 (N_29653,N_28829,N_29340);
or U29654 (N_29654,N_29134,N_29306);
nor U29655 (N_29655,N_29305,N_29015);
nor U29656 (N_29656,N_28898,N_29237);
xnor U29657 (N_29657,N_29171,N_29243);
and U29658 (N_29658,N_29099,N_29025);
nand U29659 (N_29659,N_29215,N_29367);
nand U29660 (N_29660,N_28947,N_29142);
nor U29661 (N_29661,N_29251,N_29208);
or U29662 (N_29662,N_29375,N_28803);
nand U29663 (N_29663,N_29212,N_28984);
nor U29664 (N_29664,N_28860,N_29254);
xnor U29665 (N_29665,N_29093,N_29125);
and U29666 (N_29666,N_28831,N_28941);
nor U29667 (N_29667,N_29263,N_29267);
or U29668 (N_29668,N_29316,N_28972);
nor U29669 (N_29669,N_29292,N_29176);
and U29670 (N_29670,N_29067,N_29287);
nor U29671 (N_29671,N_29302,N_29048);
nand U29672 (N_29672,N_29097,N_29047);
or U29673 (N_29673,N_28894,N_28949);
xnor U29674 (N_29674,N_29019,N_29221);
xor U29675 (N_29675,N_28889,N_28885);
nand U29676 (N_29676,N_28925,N_29130);
xnor U29677 (N_29677,N_29129,N_29363);
or U29678 (N_29678,N_28808,N_29084);
nand U29679 (N_29679,N_29232,N_28924);
or U29680 (N_29680,N_29274,N_29346);
xor U29681 (N_29681,N_29378,N_28879);
xnor U29682 (N_29682,N_29014,N_29165);
nor U29683 (N_29683,N_28980,N_29046);
nor U29684 (N_29684,N_29390,N_29388);
xnor U29685 (N_29685,N_29328,N_29342);
or U29686 (N_29686,N_28952,N_28880);
nand U29687 (N_29687,N_29100,N_28887);
nand U29688 (N_29688,N_28995,N_29116);
nor U29689 (N_29689,N_28976,N_28805);
or U29690 (N_29690,N_29111,N_28834);
and U29691 (N_29691,N_29278,N_29365);
nor U29692 (N_29692,N_29250,N_28899);
or U29693 (N_29693,N_29201,N_29122);
or U29694 (N_29694,N_28883,N_29177);
nand U29695 (N_29695,N_29148,N_29066);
nor U29696 (N_29696,N_28812,N_29010);
or U29697 (N_29697,N_29064,N_29245);
and U29698 (N_29698,N_28847,N_28871);
nor U29699 (N_29699,N_28849,N_28915);
nand U29700 (N_29700,N_28952,N_28891);
nor U29701 (N_29701,N_28831,N_28975);
nand U29702 (N_29702,N_29000,N_29002);
nand U29703 (N_29703,N_29194,N_28881);
xor U29704 (N_29704,N_29274,N_28987);
nand U29705 (N_29705,N_29317,N_29111);
and U29706 (N_29706,N_29050,N_29107);
or U29707 (N_29707,N_28851,N_29071);
nand U29708 (N_29708,N_29019,N_28884);
or U29709 (N_29709,N_28978,N_29201);
nand U29710 (N_29710,N_28804,N_29389);
xor U29711 (N_29711,N_29062,N_28821);
nand U29712 (N_29712,N_29030,N_29326);
or U29713 (N_29713,N_28839,N_29121);
nand U29714 (N_29714,N_29061,N_29298);
or U29715 (N_29715,N_29023,N_29044);
xor U29716 (N_29716,N_28885,N_29000);
xor U29717 (N_29717,N_28914,N_29025);
xor U29718 (N_29718,N_28984,N_29348);
and U29719 (N_29719,N_29130,N_29328);
nand U29720 (N_29720,N_28857,N_28903);
nor U29721 (N_29721,N_29151,N_28864);
and U29722 (N_29722,N_29016,N_29307);
xnor U29723 (N_29723,N_29021,N_28945);
or U29724 (N_29724,N_29171,N_29224);
nor U29725 (N_29725,N_29381,N_28924);
nand U29726 (N_29726,N_29177,N_29308);
nand U29727 (N_29727,N_29345,N_29121);
nand U29728 (N_29728,N_28906,N_29334);
xnor U29729 (N_29729,N_28902,N_29393);
and U29730 (N_29730,N_29124,N_29308);
nor U29731 (N_29731,N_28962,N_29057);
and U29732 (N_29732,N_29091,N_29240);
xnor U29733 (N_29733,N_28835,N_28866);
nor U29734 (N_29734,N_29342,N_29103);
nand U29735 (N_29735,N_29315,N_29390);
or U29736 (N_29736,N_29231,N_28922);
nor U29737 (N_29737,N_29301,N_28924);
and U29738 (N_29738,N_29279,N_29277);
or U29739 (N_29739,N_29358,N_29229);
and U29740 (N_29740,N_28915,N_29164);
nor U29741 (N_29741,N_28988,N_29143);
xnor U29742 (N_29742,N_28899,N_28972);
or U29743 (N_29743,N_28823,N_29109);
nor U29744 (N_29744,N_28929,N_28847);
xnor U29745 (N_29745,N_28842,N_29057);
xnor U29746 (N_29746,N_29361,N_29282);
or U29747 (N_29747,N_29391,N_28882);
or U29748 (N_29748,N_28943,N_28820);
nor U29749 (N_29749,N_28998,N_29007);
or U29750 (N_29750,N_28827,N_29308);
xnor U29751 (N_29751,N_29315,N_28934);
nor U29752 (N_29752,N_28826,N_28923);
and U29753 (N_29753,N_29204,N_29233);
nand U29754 (N_29754,N_28882,N_28816);
or U29755 (N_29755,N_29117,N_28942);
xnor U29756 (N_29756,N_29209,N_29340);
nor U29757 (N_29757,N_29369,N_29135);
nand U29758 (N_29758,N_29112,N_29255);
xor U29759 (N_29759,N_29318,N_29319);
and U29760 (N_29760,N_29176,N_28821);
or U29761 (N_29761,N_29165,N_29222);
and U29762 (N_29762,N_29013,N_29219);
and U29763 (N_29763,N_29385,N_29200);
and U29764 (N_29764,N_29124,N_29116);
nor U29765 (N_29765,N_28889,N_28977);
nand U29766 (N_29766,N_28922,N_28948);
and U29767 (N_29767,N_28849,N_29215);
xor U29768 (N_29768,N_28927,N_29018);
nor U29769 (N_29769,N_29033,N_28998);
or U29770 (N_29770,N_28807,N_29267);
nand U29771 (N_29771,N_29084,N_29292);
and U29772 (N_29772,N_29067,N_29017);
nor U29773 (N_29773,N_29042,N_29035);
nand U29774 (N_29774,N_29342,N_29027);
or U29775 (N_29775,N_29142,N_29247);
xor U29776 (N_29776,N_29228,N_29123);
nor U29777 (N_29777,N_29192,N_29343);
xnor U29778 (N_29778,N_29058,N_28832);
and U29779 (N_29779,N_29158,N_29280);
and U29780 (N_29780,N_28954,N_28881);
xor U29781 (N_29781,N_29106,N_29208);
xor U29782 (N_29782,N_29300,N_29030);
nor U29783 (N_29783,N_29167,N_29002);
nand U29784 (N_29784,N_28891,N_28801);
and U29785 (N_29785,N_29285,N_29135);
nor U29786 (N_29786,N_29019,N_28899);
nand U29787 (N_29787,N_29033,N_28931);
nor U29788 (N_29788,N_29368,N_28889);
or U29789 (N_29789,N_29291,N_29371);
xnor U29790 (N_29790,N_29140,N_29310);
and U29791 (N_29791,N_29305,N_29340);
or U29792 (N_29792,N_28833,N_29276);
nand U29793 (N_29793,N_29142,N_28882);
nand U29794 (N_29794,N_29200,N_29290);
nand U29795 (N_29795,N_29177,N_29108);
and U29796 (N_29796,N_28901,N_29113);
nand U29797 (N_29797,N_29179,N_28969);
xnor U29798 (N_29798,N_29176,N_29095);
nor U29799 (N_29799,N_28840,N_29169);
or U29800 (N_29800,N_29148,N_29307);
or U29801 (N_29801,N_28913,N_29146);
xnor U29802 (N_29802,N_29376,N_29059);
and U29803 (N_29803,N_29134,N_29103);
and U29804 (N_29804,N_29242,N_28945);
nor U29805 (N_29805,N_28938,N_29251);
and U29806 (N_29806,N_28920,N_29378);
xor U29807 (N_29807,N_29271,N_29339);
nand U29808 (N_29808,N_29009,N_29104);
and U29809 (N_29809,N_29139,N_29317);
and U29810 (N_29810,N_29333,N_29002);
and U29811 (N_29811,N_28823,N_29353);
nand U29812 (N_29812,N_29276,N_29145);
and U29813 (N_29813,N_29017,N_29263);
xnor U29814 (N_29814,N_29207,N_28829);
and U29815 (N_29815,N_29286,N_28862);
xnor U29816 (N_29816,N_29011,N_29207);
nor U29817 (N_29817,N_29308,N_29017);
nor U29818 (N_29818,N_29206,N_29396);
nand U29819 (N_29819,N_28881,N_29230);
nor U29820 (N_29820,N_28983,N_29299);
nand U29821 (N_29821,N_29131,N_28818);
and U29822 (N_29822,N_29228,N_28825);
and U29823 (N_29823,N_28937,N_28814);
and U29824 (N_29824,N_29167,N_28801);
nor U29825 (N_29825,N_29101,N_29261);
or U29826 (N_29826,N_29361,N_28934);
and U29827 (N_29827,N_29088,N_29246);
nand U29828 (N_29828,N_29269,N_29384);
nor U29829 (N_29829,N_29363,N_29276);
or U29830 (N_29830,N_28944,N_29087);
xnor U29831 (N_29831,N_28866,N_29284);
and U29832 (N_29832,N_29160,N_28851);
or U29833 (N_29833,N_29289,N_29151);
nor U29834 (N_29834,N_29100,N_29253);
and U29835 (N_29835,N_29219,N_29398);
xor U29836 (N_29836,N_28828,N_29316);
xnor U29837 (N_29837,N_29070,N_29391);
nor U29838 (N_29838,N_29230,N_29041);
and U29839 (N_29839,N_29143,N_29327);
xnor U29840 (N_29840,N_28958,N_28968);
or U29841 (N_29841,N_29114,N_28925);
xor U29842 (N_29842,N_29233,N_28929);
nand U29843 (N_29843,N_29183,N_29101);
and U29844 (N_29844,N_28857,N_29187);
or U29845 (N_29845,N_29384,N_28960);
nor U29846 (N_29846,N_29204,N_29365);
and U29847 (N_29847,N_29305,N_29029);
nor U29848 (N_29848,N_29133,N_29268);
and U29849 (N_29849,N_29143,N_29231);
nor U29850 (N_29850,N_29109,N_29038);
or U29851 (N_29851,N_29304,N_29192);
nand U29852 (N_29852,N_29371,N_28851);
xor U29853 (N_29853,N_29308,N_29037);
and U29854 (N_29854,N_29114,N_28947);
nand U29855 (N_29855,N_28823,N_29232);
nand U29856 (N_29856,N_28908,N_29135);
nand U29857 (N_29857,N_29166,N_29156);
or U29858 (N_29858,N_28981,N_29072);
nor U29859 (N_29859,N_29230,N_29395);
nand U29860 (N_29860,N_29103,N_29101);
nor U29861 (N_29861,N_29057,N_29096);
xnor U29862 (N_29862,N_29027,N_28931);
nand U29863 (N_29863,N_28976,N_28852);
xor U29864 (N_29864,N_29170,N_28822);
nor U29865 (N_29865,N_28847,N_28950);
nand U29866 (N_29866,N_29315,N_28831);
or U29867 (N_29867,N_29393,N_29024);
xor U29868 (N_29868,N_29218,N_29379);
and U29869 (N_29869,N_28815,N_28829);
or U29870 (N_29870,N_29081,N_29039);
or U29871 (N_29871,N_28920,N_28869);
nand U29872 (N_29872,N_29146,N_29016);
or U29873 (N_29873,N_28849,N_29263);
or U29874 (N_29874,N_29281,N_29373);
or U29875 (N_29875,N_29089,N_29110);
xor U29876 (N_29876,N_28950,N_29045);
and U29877 (N_29877,N_28857,N_29028);
nor U29878 (N_29878,N_29253,N_29046);
xor U29879 (N_29879,N_29124,N_29042);
and U29880 (N_29880,N_29374,N_28938);
xor U29881 (N_29881,N_28835,N_28901);
or U29882 (N_29882,N_29389,N_28961);
nand U29883 (N_29883,N_28971,N_29292);
and U29884 (N_29884,N_29176,N_29354);
xnor U29885 (N_29885,N_28806,N_29067);
or U29886 (N_29886,N_29197,N_29135);
xor U29887 (N_29887,N_29071,N_29075);
xnor U29888 (N_29888,N_28930,N_29323);
nor U29889 (N_29889,N_29067,N_29187);
and U29890 (N_29890,N_29272,N_29082);
xor U29891 (N_29891,N_28970,N_29077);
or U29892 (N_29892,N_29301,N_28853);
or U29893 (N_29893,N_28951,N_29298);
nor U29894 (N_29894,N_29387,N_29329);
or U29895 (N_29895,N_29384,N_28831);
nand U29896 (N_29896,N_29051,N_29334);
and U29897 (N_29897,N_29384,N_29280);
nand U29898 (N_29898,N_29122,N_29359);
nand U29899 (N_29899,N_29056,N_28862);
xnor U29900 (N_29900,N_29165,N_29005);
or U29901 (N_29901,N_29262,N_29283);
xor U29902 (N_29902,N_28944,N_28824);
or U29903 (N_29903,N_28851,N_29356);
or U29904 (N_29904,N_29387,N_29013);
and U29905 (N_29905,N_29187,N_29224);
nor U29906 (N_29906,N_29212,N_29223);
nor U29907 (N_29907,N_29349,N_28872);
xnor U29908 (N_29908,N_29040,N_29285);
and U29909 (N_29909,N_29277,N_29060);
xnor U29910 (N_29910,N_28888,N_29302);
nor U29911 (N_29911,N_29350,N_29288);
xor U29912 (N_29912,N_29247,N_29383);
nand U29913 (N_29913,N_29340,N_29214);
and U29914 (N_29914,N_29219,N_29232);
and U29915 (N_29915,N_29146,N_28840);
nand U29916 (N_29916,N_28939,N_28856);
xor U29917 (N_29917,N_28921,N_29365);
and U29918 (N_29918,N_29107,N_28828);
nor U29919 (N_29919,N_29128,N_28805);
and U29920 (N_29920,N_28849,N_29351);
nand U29921 (N_29921,N_28814,N_29289);
or U29922 (N_29922,N_29309,N_29296);
nor U29923 (N_29923,N_29097,N_29062);
nand U29924 (N_29924,N_29355,N_29363);
nor U29925 (N_29925,N_29239,N_29121);
or U29926 (N_29926,N_28886,N_28922);
xor U29927 (N_29927,N_28934,N_29280);
nor U29928 (N_29928,N_28816,N_29280);
nor U29929 (N_29929,N_29015,N_28926);
nand U29930 (N_29930,N_28905,N_28805);
xnor U29931 (N_29931,N_29291,N_29127);
or U29932 (N_29932,N_29107,N_28970);
nand U29933 (N_29933,N_29380,N_29294);
xnor U29934 (N_29934,N_29226,N_28931);
or U29935 (N_29935,N_28898,N_28999);
nand U29936 (N_29936,N_29329,N_29166);
nand U29937 (N_29937,N_29378,N_29012);
or U29938 (N_29938,N_29337,N_28821);
and U29939 (N_29939,N_29366,N_29220);
xor U29940 (N_29940,N_28975,N_29353);
or U29941 (N_29941,N_29048,N_29098);
xor U29942 (N_29942,N_28982,N_29040);
nor U29943 (N_29943,N_29375,N_29230);
xor U29944 (N_29944,N_29247,N_29018);
or U29945 (N_29945,N_28877,N_28828);
and U29946 (N_29946,N_28819,N_28965);
nor U29947 (N_29947,N_29093,N_29164);
xnor U29948 (N_29948,N_28874,N_29290);
nor U29949 (N_29949,N_29125,N_29031);
and U29950 (N_29950,N_29178,N_28917);
nand U29951 (N_29951,N_29174,N_29096);
nor U29952 (N_29952,N_29232,N_29394);
nor U29953 (N_29953,N_28963,N_29344);
nor U29954 (N_29954,N_28824,N_28978);
xor U29955 (N_29955,N_28981,N_29210);
nand U29956 (N_29956,N_28847,N_29040);
xor U29957 (N_29957,N_29240,N_29050);
nand U29958 (N_29958,N_28962,N_29368);
and U29959 (N_29959,N_29346,N_28972);
xnor U29960 (N_29960,N_28963,N_28800);
and U29961 (N_29961,N_29223,N_29256);
xnor U29962 (N_29962,N_28876,N_28973);
xnor U29963 (N_29963,N_29025,N_28807);
and U29964 (N_29964,N_29082,N_29238);
nor U29965 (N_29965,N_29027,N_29297);
or U29966 (N_29966,N_28843,N_29333);
and U29967 (N_29967,N_28834,N_28910);
xnor U29968 (N_29968,N_29311,N_28833);
nor U29969 (N_29969,N_29123,N_28995);
or U29970 (N_29970,N_29022,N_28974);
or U29971 (N_29971,N_29175,N_29363);
and U29972 (N_29972,N_29014,N_28882);
or U29973 (N_29973,N_29140,N_29142);
xor U29974 (N_29974,N_29388,N_29152);
and U29975 (N_29975,N_29031,N_29015);
nand U29976 (N_29976,N_29176,N_28842);
nand U29977 (N_29977,N_28876,N_29061);
xnor U29978 (N_29978,N_29353,N_28822);
nor U29979 (N_29979,N_29157,N_28952);
nor U29980 (N_29980,N_28936,N_28920);
or U29981 (N_29981,N_29230,N_29162);
xor U29982 (N_29982,N_28940,N_29387);
or U29983 (N_29983,N_28850,N_29009);
nor U29984 (N_29984,N_28918,N_28981);
xor U29985 (N_29985,N_29218,N_29049);
xor U29986 (N_29986,N_28827,N_28885);
nand U29987 (N_29987,N_29192,N_29368);
nand U29988 (N_29988,N_29100,N_29283);
or U29989 (N_29989,N_29036,N_28868);
nor U29990 (N_29990,N_29004,N_29103);
xor U29991 (N_29991,N_29137,N_29035);
nor U29992 (N_29992,N_29027,N_28867);
or U29993 (N_29993,N_28863,N_28935);
or U29994 (N_29994,N_28841,N_29048);
and U29995 (N_29995,N_29204,N_28827);
xor U29996 (N_29996,N_29050,N_29074);
or U29997 (N_29997,N_29372,N_29143);
xor U29998 (N_29998,N_29277,N_29349);
or U29999 (N_29999,N_28991,N_29216);
xnor UO_0 (O_0,N_29844,N_29428);
or UO_1 (O_1,N_29523,N_29920);
or UO_2 (O_2,N_29611,N_29777);
and UO_3 (O_3,N_29785,N_29446);
nand UO_4 (O_4,N_29524,N_29616);
and UO_5 (O_5,N_29940,N_29765);
nand UO_6 (O_6,N_29612,N_29815);
nor UO_7 (O_7,N_29707,N_29697);
nor UO_8 (O_8,N_29591,N_29727);
xnor UO_9 (O_9,N_29571,N_29775);
or UO_10 (O_10,N_29967,N_29676);
nand UO_11 (O_11,N_29580,N_29534);
or UO_12 (O_12,N_29643,N_29772);
xnor UO_13 (O_13,N_29514,N_29980);
or UO_14 (O_14,N_29512,N_29749);
nor UO_15 (O_15,N_29813,N_29682);
or UO_16 (O_16,N_29829,N_29963);
nand UO_17 (O_17,N_29873,N_29850);
and UO_18 (O_18,N_29740,N_29584);
nor UO_19 (O_19,N_29566,N_29706);
or UO_20 (O_20,N_29672,N_29687);
and UO_21 (O_21,N_29631,N_29444);
xnor UO_22 (O_22,N_29503,N_29704);
xor UO_23 (O_23,N_29909,N_29652);
or UO_24 (O_24,N_29413,N_29932);
and UO_25 (O_25,N_29575,N_29482);
xor UO_26 (O_26,N_29739,N_29821);
nand UO_27 (O_27,N_29864,N_29721);
and UO_28 (O_28,N_29702,N_29748);
nand UO_29 (O_29,N_29817,N_29780);
nor UO_30 (O_30,N_29500,N_29890);
and UO_31 (O_31,N_29507,N_29870);
xor UO_32 (O_32,N_29766,N_29581);
xnor UO_33 (O_33,N_29404,N_29724);
and UO_34 (O_34,N_29690,N_29502);
nand UO_35 (O_35,N_29496,N_29730);
nor UO_36 (O_36,N_29915,N_29786);
xor UO_37 (O_37,N_29722,N_29541);
and UO_38 (O_38,N_29495,N_29912);
or UO_39 (O_39,N_29768,N_29550);
and UO_40 (O_40,N_29622,N_29568);
nor UO_41 (O_41,N_29686,N_29617);
xor UO_42 (O_42,N_29804,N_29484);
and UO_43 (O_43,N_29798,N_29480);
xnor UO_44 (O_44,N_29883,N_29421);
nor UO_45 (O_45,N_29475,N_29825);
or UO_46 (O_46,N_29752,N_29640);
or UO_47 (O_47,N_29924,N_29792);
or UO_48 (O_48,N_29645,N_29809);
nand UO_49 (O_49,N_29939,N_29756);
xor UO_50 (O_50,N_29443,N_29710);
or UO_51 (O_51,N_29543,N_29906);
and UO_52 (O_52,N_29695,N_29412);
or UO_53 (O_53,N_29982,N_29891);
nand UO_54 (O_54,N_29615,N_29888);
xnor UO_55 (O_55,N_29471,N_29726);
xnor UO_56 (O_56,N_29598,N_29958);
nand UO_57 (O_57,N_29790,N_29876);
nor UO_58 (O_58,N_29972,N_29983);
nor UO_59 (O_59,N_29538,N_29973);
nand UO_60 (O_60,N_29455,N_29565);
nand UO_61 (O_61,N_29981,N_29681);
or UO_62 (O_62,N_29636,N_29540);
xnor UO_63 (O_63,N_29411,N_29819);
xor UO_64 (O_64,N_29409,N_29713);
and UO_65 (O_65,N_29732,N_29468);
or UO_66 (O_66,N_29564,N_29606);
or UO_67 (O_67,N_29991,N_29644);
nand UO_68 (O_68,N_29782,N_29593);
nand UO_69 (O_69,N_29634,N_29814);
or UO_70 (O_70,N_29483,N_29789);
nor UO_71 (O_71,N_29557,N_29947);
xnor UO_72 (O_72,N_29429,N_29918);
xor UO_73 (O_73,N_29406,N_29755);
nand UO_74 (O_74,N_29859,N_29460);
and UO_75 (O_75,N_29402,N_29653);
or UO_76 (O_76,N_29922,N_29490);
nand UO_77 (O_77,N_29826,N_29989);
and UO_78 (O_78,N_29678,N_29492);
nand UO_79 (O_79,N_29951,N_29916);
xnor UO_80 (O_80,N_29843,N_29555);
xor UO_81 (O_81,N_29810,N_29868);
and UO_82 (O_82,N_29667,N_29688);
and UO_83 (O_83,N_29552,N_29491);
and UO_84 (O_84,N_29520,N_29419);
nor UO_85 (O_85,N_29486,N_29497);
nand UO_86 (O_86,N_29589,N_29453);
or UO_87 (O_87,N_29999,N_29791);
and UO_88 (O_88,N_29579,N_29563);
nand UO_89 (O_89,N_29527,N_29965);
or UO_90 (O_90,N_29624,N_29769);
and UO_91 (O_91,N_29669,N_29416);
and UO_92 (O_92,N_29554,N_29797);
and UO_93 (O_93,N_29609,N_29910);
and UO_94 (O_94,N_29731,N_29937);
nor UO_95 (O_95,N_29662,N_29424);
or UO_96 (O_96,N_29608,N_29641);
and UO_97 (O_97,N_29614,N_29974);
and UO_98 (O_98,N_29637,N_29470);
and UO_99 (O_99,N_29917,N_29767);
xnor UO_100 (O_100,N_29773,N_29998);
and UO_101 (O_101,N_29833,N_29699);
xor UO_102 (O_102,N_29417,N_29881);
nor UO_103 (O_103,N_29400,N_29546);
nor UO_104 (O_104,N_29418,N_29473);
nand UO_105 (O_105,N_29592,N_29405);
and UO_106 (O_106,N_29865,N_29807);
and UO_107 (O_107,N_29990,N_29816);
nand UO_108 (O_108,N_29458,N_29465);
xor UO_109 (O_109,N_29671,N_29898);
nor UO_110 (O_110,N_29479,N_29853);
and UO_111 (O_111,N_29505,N_29956);
and UO_112 (O_112,N_29832,N_29494);
and UO_113 (O_113,N_29855,N_29863);
nor UO_114 (O_114,N_29633,N_29802);
or UO_115 (O_115,N_29913,N_29733);
xor UO_116 (O_116,N_29587,N_29900);
and UO_117 (O_117,N_29680,N_29577);
or UO_118 (O_118,N_29753,N_29911);
xor UO_119 (O_119,N_29812,N_29747);
or UO_120 (O_120,N_29808,N_29574);
xnor UO_121 (O_121,N_29501,N_29811);
or UO_122 (O_122,N_29582,N_29858);
and UO_123 (O_123,N_29744,N_29685);
nor UO_124 (O_124,N_29978,N_29668);
and UO_125 (O_125,N_29403,N_29720);
and UO_126 (O_126,N_29759,N_29472);
or UO_127 (O_127,N_29701,N_29447);
and UO_128 (O_128,N_29683,N_29799);
nand UO_129 (O_129,N_29892,N_29877);
nor UO_130 (O_130,N_29728,N_29474);
or UO_131 (O_131,N_29996,N_29845);
and UO_132 (O_132,N_29547,N_29698);
nand UO_133 (O_133,N_29905,N_29950);
or UO_134 (O_134,N_29602,N_29570);
or UO_135 (O_135,N_29462,N_29800);
or UO_136 (O_136,N_29851,N_29549);
and UO_137 (O_137,N_29971,N_29806);
or UO_138 (O_138,N_29415,N_29757);
nor UO_139 (O_139,N_29871,N_29528);
and UO_140 (O_140,N_29992,N_29679);
nand UO_141 (O_141,N_29481,N_29935);
and UO_142 (O_142,N_29432,N_29793);
or UO_143 (O_143,N_29499,N_29774);
and UO_144 (O_144,N_29613,N_29839);
or UO_145 (O_145,N_29510,N_29831);
nor UO_146 (O_146,N_29887,N_29776);
nand UO_147 (O_147,N_29788,N_29542);
xor UO_148 (O_148,N_29944,N_29830);
or UO_149 (O_149,N_29860,N_29869);
nand UO_150 (O_150,N_29493,N_29504);
nand UO_151 (O_151,N_29738,N_29431);
xor UO_152 (O_152,N_29840,N_29573);
and UO_153 (O_153,N_29969,N_29452);
and UO_154 (O_154,N_29993,N_29854);
xnor UO_155 (O_155,N_29878,N_29626);
xor UO_156 (O_156,N_29664,N_29723);
or UO_157 (O_157,N_29457,N_29834);
xnor UO_158 (O_158,N_29977,N_29604);
or UO_159 (O_159,N_29955,N_29919);
xor UO_160 (O_160,N_29422,N_29796);
and UO_161 (O_161,N_29410,N_29879);
or UO_162 (O_162,N_29805,N_29658);
nor UO_163 (O_163,N_29841,N_29908);
xor UO_164 (O_164,N_29885,N_29477);
xnor UO_165 (O_165,N_29567,N_29530);
nand UO_166 (O_166,N_29619,N_29539);
or UO_167 (O_167,N_29561,N_29449);
nand UO_168 (O_168,N_29556,N_29929);
and UO_169 (O_169,N_29770,N_29838);
xor UO_170 (O_170,N_29938,N_29737);
xor UO_171 (O_171,N_29875,N_29795);
nand UO_172 (O_172,N_29642,N_29849);
or UO_173 (O_173,N_29880,N_29434);
nor UO_174 (O_174,N_29709,N_29425);
and UO_175 (O_175,N_29670,N_29866);
or UO_176 (O_176,N_29901,N_29933);
xnor UO_177 (O_177,N_29628,N_29848);
xor UO_178 (O_178,N_29674,N_29522);
or UO_179 (O_179,N_29435,N_29985);
and UO_180 (O_180,N_29525,N_29560);
nor UO_181 (O_181,N_29648,N_29954);
nor UO_182 (O_182,N_29407,N_29454);
or UO_183 (O_183,N_29605,N_29521);
nor UO_184 (O_184,N_29941,N_29837);
nor UO_185 (O_185,N_29735,N_29625);
nor UO_186 (O_186,N_29957,N_29758);
or UO_187 (O_187,N_29448,N_29513);
nor UO_188 (O_188,N_29894,N_29533);
nand UO_189 (O_189,N_29976,N_29907);
and UO_190 (O_190,N_29590,N_29746);
xnor UO_191 (O_191,N_29842,N_29548);
and UO_192 (O_192,N_29559,N_29536);
and UO_193 (O_193,N_29703,N_29714);
nor UO_194 (O_194,N_29466,N_29818);
and UO_195 (O_195,N_29856,N_29741);
nand UO_196 (O_196,N_29961,N_29923);
or UO_197 (O_197,N_29588,N_29517);
nand UO_198 (O_198,N_29902,N_29930);
nand UO_199 (O_199,N_29433,N_29437);
and UO_200 (O_200,N_29659,N_29635);
or UO_201 (O_201,N_29820,N_29595);
xnor UO_202 (O_202,N_29666,N_29899);
nor UO_203 (O_203,N_29884,N_29927);
nand UO_204 (O_204,N_29762,N_29600);
nor UO_205 (O_205,N_29716,N_29632);
and UO_206 (O_206,N_29948,N_29994);
and UO_207 (O_207,N_29784,N_29836);
nor UO_208 (O_208,N_29962,N_29966);
and UO_209 (O_209,N_29692,N_29651);
nor UO_210 (O_210,N_29787,N_29596);
xor UO_211 (O_211,N_29953,N_29456);
or UO_212 (O_212,N_29488,N_29427);
nand UO_213 (O_213,N_29846,N_29712);
or UO_214 (O_214,N_29464,N_29896);
nor UO_215 (O_215,N_29618,N_29903);
nor UO_216 (O_216,N_29675,N_29509);
nor UO_217 (O_217,N_29526,N_29979);
or UO_218 (O_218,N_29751,N_29964);
xnor UO_219 (O_219,N_29673,N_29544);
nor UO_220 (O_220,N_29997,N_29914);
nor UO_221 (O_221,N_29426,N_29694);
xnor UO_222 (O_222,N_29578,N_29943);
nand UO_223 (O_223,N_29511,N_29778);
and UO_224 (O_224,N_29754,N_29897);
nor UO_225 (O_225,N_29771,N_29705);
xnor UO_226 (O_226,N_29439,N_29931);
xnor UO_227 (O_227,N_29408,N_29764);
and UO_228 (O_228,N_29663,N_29857);
nand UO_229 (O_229,N_29506,N_29760);
and UO_230 (O_230,N_29599,N_29414);
nor UO_231 (O_231,N_29779,N_29742);
xor UO_232 (O_232,N_29441,N_29485);
nand UO_233 (O_233,N_29750,N_29401);
nor UO_234 (O_234,N_29691,N_29968);
xnor UO_235 (O_235,N_29803,N_29715);
xor UO_236 (O_236,N_29655,N_29597);
xor UO_237 (O_237,N_29459,N_29783);
and UO_238 (O_238,N_29970,N_29987);
and UO_239 (O_239,N_29586,N_29984);
nor UO_240 (O_240,N_29629,N_29835);
xor UO_241 (O_241,N_29508,N_29696);
nand UO_242 (O_242,N_29516,N_29423);
and UO_243 (O_243,N_29921,N_29646);
xor UO_244 (O_244,N_29558,N_29824);
nand UO_245 (O_245,N_29975,N_29576);
or UO_246 (O_246,N_29620,N_29562);
or UO_247 (O_247,N_29665,N_29736);
and UO_248 (O_248,N_29420,N_29700);
or UO_249 (O_249,N_29719,N_29654);
and UO_250 (O_250,N_29450,N_29445);
and UO_251 (O_251,N_29630,N_29545);
and UO_252 (O_252,N_29729,N_29861);
nor UO_253 (O_253,N_29828,N_29794);
and UO_254 (O_254,N_29693,N_29822);
and UO_255 (O_255,N_29489,N_29717);
or UO_256 (O_256,N_29551,N_29874);
nor UO_257 (O_257,N_29518,N_29601);
nor UO_258 (O_258,N_29451,N_29743);
and UO_259 (O_259,N_29478,N_29708);
nand UO_260 (O_260,N_29781,N_29761);
xor UO_261 (O_261,N_29904,N_29519);
xnor UO_262 (O_262,N_29827,N_29936);
nand UO_263 (O_263,N_29531,N_29585);
and UO_264 (O_264,N_29610,N_29893);
nor UO_265 (O_265,N_29438,N_29487);
nand UO_266 (O_266,N_29677,N_29461);
or UO_267 (O_267,N_29661,N_29718);
and UO_268 (O_268,N_29430,N_29532);
or UO_269 (O_269,N_29436,N_29607);
and UO_270 (O_270,N_29657,N_29476);
and UO_271 (O_271,N_29515,N_29537);
or UO_272 (O_272,N_29952,N_29734);
or UO_273 (O_273,N_29942,N_29960);
xor UO_274 (O_274,N_29725,N_29745);
nand UO_275 (O_275,N_29623,N_29603);
and UO_276 (O_276,N_29882,N_29862);
xor UO_277 (O_277,N_29959,N_29711);
nor UO_278 (O_278,N_29852,N_29529);
nor UO_279 (O_279,N_29801,N_29535);
nor UO_280 (O_280,N_29650,N_29945);
and UO_281 (O_281,N_29627,N_29660);
and UO_282 (O_282,N_29442,N_29689);
nor UO_283 (O_283,N_29934,N_29498);
or UO_284 (O_284,N_29867,N_29440);
and UO_285 (O_285,N_29572,N_29926);
and UO_286 (O_286,N_29889,N_29847);
nand UO_287 (O_287,N_29469,N_29895);
nor UO_288 (O_288,N_29684,N_29823);
and UO_289 (O_289,N_29986,N_29886);
nand UO_290 (O_290,N_29594,N_29946);
nand UO_291 (O_291,N_29553,N_29949);
xnor UO_292 (O_292,N_29569,N_29621);
nor UO_293 (O_293,N_29647,N_29649);
xnor UO_294 (O_294,N_29463,N_29638);
and UO_295 (O_295,N_29763,N_29639);
and UO_296 (O_296,N_29925,N_29995);
or UO_297 (O_297,N_29467,N_29928);
xnor UO_298 (O_298,N_29583,N_29872);
nand UO_299 (O_299,N_29656,N_29988);
xor UO_300 (O_300,N_29812,N_29651);
or UO_301 (O_301,N_29881,N_29964);
nand UO_302 (O_302,N_29834,N_29692);
nand UO_303 (O_303,N_29787,N_29662);
nand UO_304 (O_304,N_29641,N_29499);
or UO_305 (O_305,N_29518,N_29740);
or UO_306 (O_306,N_29876,N_29571);
xor UO_307 (O_307,N_29877,N_29511);
xnor UO_308 (O_308,N_29990,N_29846);
and UO_309 (O_309,N_29597,N_29472);
xnor UO_310 (O_310,N_29504,N_29748);
and UO_311 (O_311,N_29945,N_29432);
nand UO_312 (O_312,N_29507,N_29468);
nor UO_313 (O_313,N_29616,N_29622);
or UO_314 (O_314,N_29982,N_29417);
xnor UO_315 (O_315,N_29530,N_29891);
xnor UO_316 (O_316,N_29543,N_29781);
or UO_317 (O_317,N_29447,N_29543);
nand UO_318 (O_318,N_29470,N_29716);
or UO_319 (O_319,N_29930,N_29982);
or UO_320 (O_320,N_29564,N_29773);
and UO_321 (O_321,N_29456,N_29812);
xnor UO_322 (O_322,N_29602,N_29723);
or UO_323 (O_323,N_29905,N_29705);
nor UO_324 (O_324,N_29829,N_29491);
nand UO_325 (O_325,N_29833,N_29905);
nand UO_326 (O_326,N_29429,N_29420);
xnor UO_327 (O_327,N_29569,N_29588);
nand UO_328 (O_328,N_29909,N_29613);
or UO_329 (O_329,N_29517,N_29490);
or UO_330 (O_330,N_29721,N_29897);
or UO_331 (O_331,N_29471,N_29665);
or UO_332 (O_332,N_29665,N_29893);
nor UO_333 (O_333,N_29928,N_29631);
nand UO_334 (O_334,N_29451,N_29763);
or UO_335 (O_335,N_29972,N_29700);
nor UO_336 (O_336,N_29433,N_29417);
nand UO_337 (O_337,N_29958,N_29483);
or UO_338 (O_338,N_29657,N_29443);
xnor UO_339 (O_339,N_29679,N_29837);
xnor UO_340 (O_340,N_29411,N_29829);
xor UO_341 (O_341,N_29463,N_29525);
or UO_342 (O_342,N_29525,N_29610);
and UO_343 (O_343,N_29466,N_29554);
and UO_344 (O_344,N_29864,N_29553);
and UO_345 (O_345,N_29451,N_29813);
nor UO_346 (O_346,N_29672,N_29944);
nor UO_347 (O_347,N_29707,N_29603);
nand UO_348 (O_348,N_29819,N_29733);
or UO_349 (O_349,N_29566,N_29915);
xor UO_350 (O_350,N_29664,N_29663);
or UO_351 (O_351,N_29862,N_29953);
and UO_352 (O_352,N_29723,N_29550);
and UO_353 (O_353,N_29702,N_29444);
and UO_354 (O_354,N_29411,N_29966);
nand UO_355 (O_355,N_29923,N_29559);
nor UO_356 (O_356,N_29428,N_29584);
or UO_357 (O_357,N_29884,N_29955);
xnor UO_358 (O_358,N_29483,N_29996);
or UO_359 (O_359,N_29687,N_29849);
and UO_360 (O_360,N_29685,N_29463);
xnor UO_361 (O_361,N_29913,N_29657);
nor UO_362 (O_362,N_29948,N_29663);
and UO_363 (O_363,N_29753,N_29885);
and UO_364 (O_364,N_29694,N_29876);
nor UO_365 (O_365,N_29667,N_29839);
nor UO_366 (O_366,N_29891,N_29694);
nand UO_367 (O_367,N_29704,N_29999);
xor UO_368 (O_368,N_29790,N_29580);
nand UO_369 (O_369,N_29999,N_29552);
nand UO_370 (O_370,N_29835,N_29672);
xor UO_371 (O_371,N_29629,N_29764);
nor UO_372 (O_372,N_29780,N_29921);
and UO_373 (O_373,N_29507,N_29767);
nor UO_374 (O_374,N_29486,N_29570);
and UO_375 (O_375,N_29826,N_29646);
nand UO_376 (O_376,N_29879,N_29616);
or UO_377 (O_377,N_29778,N_29763);
nand UO_378 (O_378,N_29873,N_29502);
nor UO_379 (O_379,N_29710,N_29470);
nand UO_380 (O_380,N_29745,N_29889);
or UO_381 (O_381,N_29858,N_29615);
or UO_382 (O_382,N_29615,N_29672);
xnor UO_383 (O_383,N_29730,N_29888);
nand UO_384 (O_384,N_29951,N_29463);
or UO_385 (O_385,N_29465,N_29873);
nor UO_386 (O_386,N_29970,N_29404);
nor UO_387 (O_387,N_29669,N_29802);
xnor UO_388 (O_388,N_29978,N_29804);
nand UO_389 (O_389,N_29933,N_29413);
nand UO_390 (O_390,N_29576,N_29686);
and UO_391 (O_391,N_29889,N_29905);
xor UO_392 (O_392,N_29968,N_29743);
and UO_393 (O_393,N_29693,N_29700);
nor UO_394 (O_394,N_29664,N_29526);
nand UO_395 (O_395,N_29582,N_29789);
and UO_396 (O_396,N_29741,N_29617);
nand UO_397 (O_397,N_29629,N_29682);
xnor UO_398 (O_398,N_29854,N_29852);
xor UO_399 (O_399,N_29552,N_29864);
nor UO_400 (O_400,N_29951,N_29455);
nor UO_401 (O_401,N_29912,N_29946);
nand UO_402 (O_402,N_29690,N_29965);
and UO_403 (O_403,N_29795,N_29854);
and UO_404 (O_404,N_29994,N_29411);
nor UO_405 (O_405,N_29963,N_29786);
nor UO_406 (O_406,N_29653,N_29533);
xor UO_407 (O_407,N_29488,N_29538);
nor UO_408 (O_408,N_29649,N_29760);
and UO_409 (O_409,N_29808,N_29792);
nor UO_410 (O_410,N_29694,N_29818);
nor UO_411 (O_411,N_29567,N_29600);
and UO_412 (O_412,N_29699,N_29918);
and UO_413 (O_413,N_29845,N_29968);
or UO_414 (O_414,N_29975,N_29612);
or UO_415 (O_415,N_29431,N_29736);
nor UO_416 (O_416,N_29508,N_29700);
and UO_417 (O_417,N_29473,N_29731);
nand UO_418 (O_418,N_29881,N_29610);
or UO_419 (O_419,N_29948,N_29494);
nand UO_420 (O_420,N_29893,N_29604);
xnor UO_421 (O_421,N_29416,N_29650);
nor UO_422 (O_422,N_29970,N_29827);
xor UO_423 (O_423,N_29895,N_29602);
or UO_424 (O_424,N_29582,N_29958);
xnor UO_425 (O_425,N_29738,N_29479);
or UO_426 (O_426,N_29842,N_29451);
xnor UO_427 (O_427,N_29842,N_29690);
nor UO_428 (O_428,N_29921,N_29683);
xnor UO_429 (O_429,N_29683,N_29626);
xor UO_430 (O_430,N_29900,N_29872);
or UO_431 (O_431,N_29516,N_29503);
and UO_432 (O_432,N_29407,N_29825);
xor UO_433 (O_433,N_29520,N_29611);
or UO_434 (O_434,N_29900,N_29600);
or UO_435 (O_435,N_29677,N_29546);
xnor UO_436 (O_436,N_29661,N_29671);
and UO_437 (O_437,N_29703,N_29887);
nor UO_438 (O_438,N_29866,N_29516);
and UO_439 (O_439,N_29762,N_29407);
xor UO_440 (O_440,N_29512,N_29572);
nand UO_441 (O_441,N_29998,N_29713);
or UO_442 (O_442,N_29910,N_29468);
and UO_443 (O_443,N_29465,N_29803);
and UO_444 (O_444,N_29494,N_29784);
nor UO_445 (O_445,N_29826,N_29539);
and UO_446 (O_446,N_29660,N_29753);
nor UO_447 (O_447,N_29402,N_29920);
nor UO_448 (O_448,N_29684,N_29712);
and UO_449 (O_449,N_29981,N_29882);
nand UO_450 (O_450,N_29517,N_29445);
nand UO_451 (O_451,N_29644,N_29446);
and UO_452 (O_452,N_29415,N_29932);
xnor UO_453 (O_453,N_29782,N_29610);
and UO_454 (O_454,N_29787,N_29448);
or UO_455 (O_455,N_29720,N_29588);
or UO_456 (O_456,N_29699,N_29480);
or UO_457 (O_457,N_29661,N_29895);
or UO_458 (O_458,N_29547,N_29695);
nand UO_459 (O_459,N_29856,N_29505);
xnor UO_460 (O_460,N_29880,N_29966);
and UO_461 (O_461,N_29642,N_29885);
or UO_462 (O_462,N_29636,N_29879);
or UO_463 (O_463,N_29733,N_29569);
nand UO_464 (O_464,N_29779,N_29471);
nor UO_465 (O_465,N_29820,N_29508);
nand UO_466 (O_466,N_29787,N_29929);
xnor UO_467 (O_467,N_29816,N_29573);
nand UO_468 (O_468,N_29702,N_29845);
nor UO_469 (O_469,N_29513,N_29829);
or UO_470 (O_470,N_29666,N_29730);
nor UO_471 (O_471,N_29657,N_29740);
xor UO_472 (O_472,N_29772,N_29722);
nor UO_473 (O_473,N_29408,N_29478);
xor UO_474 (O_474,N_29986,N_29954);
nand UO_475 (O_475,N_29666,N_29464);
xnor UO_476 (O_476,N_29853,N_29459);
xnor UO_477 (O_477,N_29405,N_29951);
nor UO_478 (O_478,N_29953,N_29485);
and UO_479 (O_479,N_29586,N_29623);
nor UO_480 (O_480,N_29502,N_29849);
nor UO_481 (O_481,N_29418,N_29553);
nand UO_482 (O_482,N_29629,N_29872);
nand UO_483 (O_483,N_29674,N_29946);
xnor UO_484 (O_484,N_29641,N_29752);
or UO_485 (O_485,N_29862,N_29528);
and UO_486 (O_486,N_29485,N_29474);
or UO_487 (O_487,N_29694,N_29540);
nor UO_488 (O_488,N_29457,N_29771);
or UO_489 (O_489,N_29962,N_29973);
nor UO_490 (O_490,N_29650,N_29861);
xor UO_491 (O_491,N_29577,N_29424);
or UO_492 (O_492,N_29447,N_29912);
or UO_493 (O_493,N_29584,N_29562);
nand UO_494 (O_494,N_29545,N_29541);
xnor UO_495 (O_495,N_29614,N_29886);
nor UO_496 (O_496,N_29837,N_29993);
nor UO_497 (O_497,N_29970,N_29998);
nand UO_498 (O_498,N_29439,N_29757);
xor UO_499 (O_499,N_29785,N_29428);
or UO_500 (O_500,N_29946,N_29801);
nand UO_501 (O_501,N_29848,N_29414);
or UO_502 (O_502,N_29600,N_29666);
xnor UO_503 (O_503,N_29804,N_29902);
or UO_504 (O_504,N_29497,N_29922);
nand UO_505 (O_505,N_29800,N_29951);
and UO_506 (O_506,N_29858,N_29581);
xnor UO_507 (O_507,N_29525,N_29432);
nand UO_508 (O_508,N_29796,N_29735);
and UO_509 (O_509,N_29704,N_29875);
nor UO_510 (O_510,N_29423,N_29560);
nand UO_511 (O_511,N_29651,N_29492);
nand UO_512 (O_512,N_29454,N_29692);
nand UO_513 (O_513,N_29754,N_29478);
or UO_514 (O_514,N_29471,N_29423);
or UO_515 (O_515,N_29752,N_29569);
or UO_516 (O_516,N_29747,N_29620);
and UO_517 (O_517,N_29984,N_29495);
or UO_518 (O_518,N_29415,N_29849);
and UO_519 (O_519,N_29475,N_29888);
xnor UO_520 (O_520,N_29812,N_29654);
nand UO_521 (O_521,N_29905,N_29911);
or UO_522 (O_522,N_29833,N_29426);
or UO_523 (O_523,N_29499,N_29473);
or UO_524 (O_524,N_29478,N_29554);
and UO_525 (O_525,N_29567,N_29882);
xnor UO_526 (O_526,N_29788,N_29445);
nand UO_527 (O_527,N_29537,N_29630);
nor UO_528 (O_528,N_29524,N_29853);
xor UO_529 (O_529,N_29583,N_29841);
xnor UO_530 (O_530,N_29994,N_29509);
nor UO_531 (O_531,N_29436,N_29762);
or UO_532 (O_532,N_29716,N_29581);
or UO_533 (O_533,N_29599,N_29510);
nand UO_534 (O_534,N_29990,N_29944);
nand UO_535 (O_535,N_29532,N_29755);
and UO_536 (O_536,N_29421,N_29442);
or UO_537 (O_537,N_29400,N_29741);
or UO_538 (O_538,N_29930,N_29445);
nor UO_539 (O_539,N_29915,N_29461);
or UO_540 (O_540,N_29603,N_29804);
nor UO_541 (O_541,N_29989,N_29484);
xor UO_542 (O_542,N_29652,N_29956);
and UO_543 (O_543,N_29527,N_29748);
xor UO_544 (O_544,N_29682,N_29871);
nand UO_545 (O_545,N_29821,N_29507);
nor UO_546 (O_546,N_29812,N_29429);
xnor UO_547 (O_547,N_29696,N_29809);
nand UO_548 (O_548,N_29766,N_29460);
and UO_549 (O_549,N_29537,N_29933);
and UO_550 (O_550,N_29852,N_29737);
and UO_551 (O_551,N_29942,N_29623);
nor UO_552 (O_552,N_29913,N_29725);
nand UO_553 (O_553,N_29784,N_29587);
nor UO_554 (O_554,N_29788,N_29602);
nand UO_555 (O_555,N_29774,N_29440);
nand UO_556 (O_556,N_29983,N_29431);
nand UO_557 (O_557,N_29933,N_29929);
nor UO_558 (O_558,N_29752,N_29416);
xor UO_559 (O_559,N_29915,N_29927);
nor UO_560 (O_560,N_29486,N_29725);
nand UO_561 (O_561,N_29822,N_29852);
xor UO_562 (O_562,N_29501,N_29642);
and UO_563 (O_563,N_29900,N_29879);
nand UO_564 (O_564,N_29570,N_29477);
nor UO_565 (O_565,N_29591,N_29682);
nand UO_566 (O_566,N_29830,N_29906);
xor UO_567 (O_567,N_29551,N_29969);
and UO_568 (O_568,N_29593,N_29750);
nor UO_569 (O_569,N_29954,N_29915);
nor UO_570 (O_570,N_29722,N_29451);
xnor UO_571 (O_571,N_29538,N_29774);
or UO_572 (O_572,N_29679,N_29637);
nand UO_573 (O_573,N_29623,N_29778);
and UO_574 (O_574,N_29798,N_29689);
nor UO_575 (O_575,N_29730,N_29663);
or UO_576 (O_576,N_29855,N_29770);
nor UO_577 (O_577,N_29899,N_29501);
and UO_578 (O_578,N_29813,N_29977);
nor UO_579 (O_579,N_29976,N_29460);
nand UO_580 (O_580,N_29590,N_29942);
and UO_581 (O_581,N_29770,N_29422);
nand UO_582 (O_582,N_29600,N_29645);
or UO_583 (O_583,N_29493,N_29777);
nand UO_584 (O_584,N_29751,N_29866);
or UO_585 (O_585,N_29664,N_29759);
or UO_586 (O_586,N_29782,N_29909);
xnor UO_587 (O_587,N_29459,N_29851);
xor UO_588 (O_588,N_29904,N_29699);
or UO_589 (O_589,N_29471,N_29878);
and UO_590 (O_590,N_29630,N_29976);
and UO_591 (O_591,N_29914,N_29647);
or UO_592 (O_592,N_29506,N_29497);
or UO_593 (O_593,N_29644,N_29555);
nor UO_594 (O_594,N_29481,N_29417);
nor UO_595 (O_595,N_29970,N_29525);
and UO_596 (O_596,N_29666,N_29468);
and UO_597 (O_597,N_29491,N_29539);
nand UO_598 (O_598,N_29718,N_29580);
nand UO_599 (O_599,N_29570,N_29457);
nand UO_600 (O_600,N_29980,N_29755);
or UO_601 (O_601,N_29448,N_29490);
nand UO_602 (O_602,N_29982,N_29859);
xor UO_603 (O_603,N_29707,N_29592);
nor UO_604 (O_604,N_29538,N_29477);
nand UO_605 (O_605,N_29672,N_29888);
nor UO_606 (O_606,N_29969,N_29560);
nand UO_607 (O_607,N_29557,N_29598);
and UO_608 (O_608,N_29652,N_29889);
nor UO_609 (O_609,N_29529,N_29729);
nand UO_610 (O_610,N_29723,N_29496);
or UO_611 (O_611,N_29698,N_29559);
or UO_612 (O_612,N_29491,N_29610);
nand UO_613 (O_613,N_29960,N_29768);
or UO_614 (O_614,N_29594,N_29794);
nand UO_615 (O_615,N_29954,N_29944);
or UO_616 (O_616,N_29814,N_29699);
xor UO_617 (O_617,N_29460,N_29417);
nor UO_618 (O_618,N_29587,N_29845);
and UO_619 (O_619,N_29876,N_29463);
or UO_620 (O_620,N_29905,N_29716);
nor UO_621 (O_621,N_29492,N_29828);
nand UO_622 (O_622,N_29859,N_29819);
or UO_623 (O_623,N_29978,N_29583);
nor UO_624 (O_624,N_29547,N_29965);
and UO_625 (O_625,N_29829,N_29998);
and UO_626 (O_626,N_29719,N_29562);
nand UO_627 (O_627,N_29883,N_29938);
nand UO_628 (O_628,N_29929,N_29534);
xnor UO_629 (O_629,N_29883,N_29507);
or UO_630 (O_630,N_29432,N_29419);
or UO_631 (O_631,N_29584,N_29894);
xor UO_632 (O_632,N_29427,N_29594);
xor UO_633 (O_633,N_29882,N_29754);
xor UO_634 (O_634,N_29546,N_29607);
nand UO_635 (O_635,N_29444,N_29697);
and UO_636 (O_636,N_29541,N_29717);
and UO_637 (O_637,N_29877,N_29717);
xnor UO_638 (O_638,N_29717,N_29702);
nor UO_639 (O_639,N_29911,N_29681);
xor UO_640 (O_640,N_29992,N_29895);
nand UO_641 (O_641,N_29466,N_29509);
nand UO_642 (O_642,N_29927,N_29417);
or UO_643 (O_643,N_29653,N_29628);
nand UO_644 (O_644,N_29966,N_29922);
xnor UO_645 (O_645,N_29709,N_29934);
xnor UO_646 (O_646,N_29791,N_29519);
xor UO_647 (O_647,N_29432,N_29854);
and UO_648 (O_648,N_29852,N_29673);
nand UO_649 (O_649,N_29904,N_29508);
nor UO_650 (O_650,N_29939,N_29619);
nand UO_651 (O_651,N_29421,N_29503);
and UO_652 (O_652,N_29816,N_29539);
nand UO_653 (O_653,N_29787,N_29684);
xor UO_654 (O_654,N_29532,N_29913);
nor UO_655 (O_655,N_29495,N_29668);
or UO_656 (O_656,N_29559,N_29599);
nor UO_657 (O_657,N_29893,N_29761);
nor UO_658 (O_658,N_29885,N_29655);
and UO_659 (O_659,N_29704,N_29852);
and UO_660 (O_660,N_29737,N_29544);
and UO_661 (O_661,N_29656,N_29606);
or UO_662 (O_662,N_29675,N_29899);
and UO_663 (O_663,N_29790,N_29414);
xnor UO_664 (O_664,N_29721,N_29746);
or UO_665 (O_665,N_29941,N_29933);
or UO_666 (O_666,N_29887,N_29830);
or UO_667 (O_667,N_29819,N_29830);
nand UO_668 (O_668,N_29653,N_29549);
nor UO_669 (O_669,N_29822,N_29738);
xnor UO_670 (O_670,N_29553,N_29873);
and UO_671 (O_671,N_29417,N_29404);
xor UO_672 (O_672,N_29920,N_29961);
and UO_673 (O_673,N_29651,N_29780);
xnor UO_674 (O_674,N_29910,N_29802);
nand UO_675 (O_675,N_29778,N_29516);
nand UO_676 (O_676,N_29662,N_29676);
or UO_677 (O_677,N_29842,N_29957);
nor UO_678 (O_678,N_29922,N_29940);
or UO_679 (O_679,N_29476,N_29451);
and UO_680 (O_680,N_29591,N_29574);
or UO_681 (O_681,N_29810,N_29851);
nor UO_682 (O_682,N_29767,N_29681);
and UO_683 (O_683,N_29443,N_29738);
or UO_684 (O_684,N_29848,N_29769);
nand UO_685 (O_685,N_29548,N_29794);
nor UO_686 (O_686,N_29616,N_29907);
nor UO_687 (O_687,N_29637,N_29748);
nand UO_688 (O_688,N_29936,N_29938);
and UO_689 (O_689,N_29798,N_29479);
nand UO_690 (O_690,N_29753,N_29948);
nand UO_691 (O_691,N_29529,N_29915);
and UO_692 (O_692,N_29535,N_29807);
or UO_693 (O_693,N_29806,N_29657);
nand UO_694 (O_694,N_29881,N_29497);
nand UO_695 (O_695,N_29589,N_29648);
nor UO_696 (O_696,N_29446,N_29860);
xor UO_697 (O_697,N_29931,N_29996);
xor UO_698 (O_698,N_29481,N_29509);
or UO_699 (O_699,N_29656,N_29892);
nand UO_700 (O_700,N_29856,N_29821);
xor UO_701 (O_701,N_29833,N_29505);
nand UO_702 (O_702,N_29963,N_29620);
xor UO_703 (O_703,N_29603,N_29952);
nor UO_704 (O_704,N_29871,N_29526);
or UO_705 (O_705,N_29515,N_29803);
nor UO_706 (O_706,N_29842,N_29910);
xor UO_707 (O_707,N_29861,N_29888);
nor UO_708 (O_708,N_29921,N_29588);
xnor UO_709 (O_709,N_29628,N_29631);
or UO_710 (O_710,N_29655,N_29843);
nand UO_711 (O_711,N_29737,N_29680);
or UO_712 (O_712,N_29838,N_29798);
xor UO_713 (O_713,N_29637,N_29907);
or UO_714 (O_714,N_29799,N_29448);
nand UO_715 (O_715,N_29416,N_29979);
nor UO_716 (O_716,N_29680,N_29422);
and UO_717 (O_717,N_29431,N_29773);
and UO_718 (O_718,N_29832,N_29965);
xor UO_719 (O_719,N_29870,N_29920);
and UO_720 (O_720,N_29573,N_29574);
and UO_721 (O_721,N_29836,N_29463);
nor UO_722 (O_722,N_29783,N_29410);
and UO_723 (O_723,N_29467,N_29559);
nand UO_724 (O_724,N_29613,N_29850);
and UO_725 (O_725,N_29614,N_29928);
nor UO_726 (O_726,N_29411,N_29862);
xnor UO_727 (O_727,N_29807,N_29805);
nor UO_728 (O_728,N_29599,N_29616);
xor UO_729 (O_729,N_29629,N_29796);
nand UO_730 (O_730,N_29923,N_29527);
xnor UO_731 (O_731,N_29719,N_29914);
or UO_732 (O_732,N_29986,N_29887);
nand UO_733 (O_733,N_29418,N_29864);
or UO_734 (O_734,N_29864,N_29695);
and UO_735 (O_735,N_29965,N_29757);
nand UO_736 (O_736,N_29886,N_29546);
xnor UO_737 (O_737,N_29573,N_29675);
nand UO_738 (O_738,N_29981,N_29837);
xnor UO_739 (O_739,N_29927,N_29447);
or UO_740 (O_740,N_29837,N_29457);
or UO_741 (O_741,N_29956,N_29901);
or UO_742 (O_742,N_29893,N_29483);
or UO_743 (O_743,N_29723,N_29813);
or UO_744 (O_744,N_29429,N_29944);
nand UO_745 (O_745,N_29402,N_29950);
and UO_746 (O_746,N_29760,N_29799);
and UO_747 (O_747,N_29778,N_29966);
xnor UO_748 (O_748,N_29427,N_29838);
xnor UO_749 (O_749,N_29626,N_29817);
nor UO_750 (O_750,N_29433,N_29744);
nand UO_751 (O_751,N_29418,N_29985);
xor UO_752 (O_752,N_29472,N_29820);
or UO_753 (O_753,N_29873,N_29489);
and UO_754 (O_754,N_29785,N_29714);
nor UO_755 (O_755,N_29713,N_29419);
nor UO_756 (O_756,N_29435,N_29481);
nand UO_757 (O_757,N_29468,N_29867);
and UO_758 (O_758,N_29839,N_29738);
xor UO_759 (O_759,N_29802,N_29749);
nand UO_760 (O_760,N_29537,N_29514);
xnor UO_761 (O_761,N_29921,N_29609);
or UO_762 (O_762,N_29616,N_29999);
nor UO_763 (O_763,N_29833,N_29518);
nand UO_764 (O_764,N_29683,N_29833);
xor UO_765 (O_765,N_29493,N_29900);
xor UO_766 (O_766,N_29539,N_29964);
and UO_767 (O_767,N_29953,N_29531);
nand UO_768 (O_768,N_29779,N_29904);
nor UO_769 (O_769,N_29628,N_29552);
nor UO_770 (O_770,N_29538,N_29606);
or UO_771 (O_771,N_29402,N_29524);
nor UO_772 (O_772,N_29813,N_29907);
and UO_773 (O_773,N_29888,N_29889);
xor UO_774 (O_774,N_29513,N_29792);
nor UO_775 (O_775,N_29827,N_29894);
nand UO_776 (O_776,N_29654,N_29705);
xnor UO_777 (O_777,N_29527,N_29995);
and UO_778 (O_778,N_29852,N_29769);
xor UO_779 (O_779,N_29920,N_29714);
xor UO_780 (O_780,N_29709,N_29501);
nand UO_781 (O_781,N_29665,N_29756);
or UO_782 (O_782,N_29664,N_29469);
nor UO_783 (O_783,N_29831,N_29621);
nor UO_784 (O_784,N_29813,N_29559);
nand UO_785 (O_785,N_29580,N_29583);
and UO_786 (O_786,N_29622,N_29713);
or UO_787 (O_787,N_29430,N_29580);
nor UO_788 (O_788,N_29607,N_29624);
nor UO_789 (O_789,N_29470,N_29756);
xor UO_790 (O_790,N_29585,N_29553);
nand UO_791 (O_791,N_29664,N_29684);
nor UO_792 (O_792,N_29440,N_29974);
nand UO_793 (O_793,N_29579,N_29874);
nor UO_794 (O_794,N_29435,N_29938);
or UO_795 (O_795,N_29638,N_29968);
xor UO_796 (O_796,N_29408,N_29978);
xnor UO_797 (O_797,N_29465,N_29722);
xor UO_798 (O_798,N_29560,N_29861);
nor UO_799 (O_799,N_29752,N_29473);
and UO_800 (O_800,N_29595,N_29413);
nor UO_801 (O_801,N_29554,N_29842);
and UO_802 (O_802,N_29977,N_29529);
and UO_803 (O_803,N_29619,N_29541);
and UO_804 (O_804,N_29986,N_29847);
nor UO_805 (O_805,N_29828,N_29874);
or UO_806 (O_806,N_29635,N_29887);
nor UO_807 (O_807,N_29535,N_29676);
and UO_808 (O_808,N_29693,N_29437);
and UO_809 (O_809,N_29737,N_29669);
nand UO_810 (O_810,N_29468,N_29849);
nand UO_811 (O_811,N_29866,N_29737);
nor UO_812 (O_812,N_29928,N_29601);
nand UO_813 (O_813,N_29624,N_29474);
nor UO_814 (O_814,N_29819,N_29749);
and UO_815 (O_815,N_29661,N_29703);
and UO_816 (O_816,N_29444,N_29558);
or UO_817 (O_817,N_29456,N_29486);
and UO_818 (O_818,N_29762,N_29553);
or UO_819 (O_819,N_29583,N_29961);
nand UO_820 (O_820,N_29466,N_29804);
nand UO_821 (O_821,N_29936,N_29523);
xor UO_822 (O_822,N_29951,N_29586);
nand UO_823 (O_823,N_29754,N_29615);
and UO_824 (O_824,N_29421,N_29615);
nand UO_825 (O_825,N_29832,N_29496);
or UO_826 (O_826,N_29792,N_29509);
or UO_827 (O_827,N_29663,N_29600);
nand UO_828 (O_828,N_29602,N_29840);
and UO_829 (O_829,N_29592,N_29652);
nor UO_830 (O_830,N_29802,N_29518);
and UO_831 (O_831,N_29516,N_29781);
or UO_832 (O_832,N_29889,N_29801);
or UO_833 (O_833,N_29560,N_29803);
and UO_834 (O_834,N_29735,N_29970);
xor UO_835 (O_835,N_29931,N_29736);
nor UO_836 (O_836,N_29683,N_29788);
or UO_837 (O_837,N_29767,N_29873);
xor UO_838 (O_838,N_29922,N_29919);
and UO_839 (O_839,N_29623,N_29893);
and UO_840 (O_840,N_29570,N_29879);
nand UO_841 (O_841,N_29556,N_29456);
xnor UO_842 (O_842,N_29662,N_29778);
nor UO_843 (O_843,N_29777,N_29559);
and UO_844 (O_844,N_29530,N_29826);
or UO_845 (O_845,N_29812,N_29609);
and UO_846 (O_846,N_29651,N_29957);
and UO_847 (O_847,N_29547,N_29953);
nand UO_848 (O_848,N_29926,N_29814);
or UO_849 (O_849,N_29870,N_29431);
and UO_850 (O_850,N_29640,N_29498);
nor UO_851 (O_851,N_29772,N_29760);
or UO_852 (O_852,N_29775,N_29465);
nand UO_853 (O_853,N_29954,N_29406);
nand UO_854 (O_854,N_29717,N_29866);
nand UO_855 (O_855,N_29858,N_29941);
and UO_856 (O_856,N_29507,N_29463);
xor UO_857 (O_857,N_29969,N_29634);
nor UO_858 (O_858,N_29675,N_29456);
xor UO_859 (O_859,N_29456,N_29639);
nand UO_860 (O_860,N_29853,N_29750);
xor UO_861 (O_861,N_29685,N_29519);
or UO_862 (O_862,N_29454,N_29731);
or UO_863 (O_863,N_29875,N_29604);
xor UO_864 (O_864,N_29585,N_29704);
nor UO_865 (O_865,N_29575,N_29885);
nor UO_866 (O_866,N_29795,N_29966);
nor UO_867 (O_867,N_29910,N_29964);
xor UO_868 (O_868,N_29703,N_29979);
nand UO_869 (O_869,N_29995,N_29871);
xor UO_870 (O_870,N_29686,N_29820);
xor UO_871 (O_871,N_29764,N_29898);
nor UO_872 (O_872,N_29843,N_29967);
and UO_873 (O_873,N_29945,N_29737);
nand UO_874 (O_874,N_29900,N_29440);
and UO_875 (O_875,N_29722,N_29702);
nand UO_876 (O_876,N_29497,N_29629);
xnor UO_877 (O_877,N_29540,N_29684);
and UO_878 (O_878,N_29562,N_29418);
xor UO_879 (O_879,N_29876,N_29705);
nand UO_880 (O_880,N_29540,N_29556);
nand UO_881 (O_881,N_29443,N_29668);
xnor UO_882 (O_882,N_29906,N_29677);
nor UO_883 (O_883,N_29736,N_29587);
nand UO_884 (O_884,N_29732,N_29413);
or UO_885 (O_885,N_29410,N_29465);
and UO_886 (O_886,N_29510,N_29475);
nand UO_887 (O_887,N_29648,N_29498);
nand UO_888 (O_888,N_29783,N_29774);
nand UO_889 (O_889,N_29417,N_29488);
nor UO_890 (O_890,N_29694,N_29728);
xor UO_891 (O_891,N_29601,N_29822);
xor UO_892 (O_892,N_29846,N_29640);
nand UO_893 (O_893,N_29667,N_29629);
xor UO_894 (O_894,N_29492,N_29403);
and UO_895 (O_895,N_29689,N_29616);
xor UO_896 (O_896,N_29541,N_29503);
nor UO_897 (O_897,N_29443,N_29692);
nand UO_898 (O_898,N_29861,N_29962);
nor UO_899 (O_899,N_29571,N_29836);
nor UO_900 (O_900,N_29892,N_29416);
or UO_901 (O_901,N_29503,N_29654);
nand UO_902 (O_902,N_29881,N_29561);
and UO_903 (O_903,N_29541,N_29735);
nand UO_904 (O_904,N_29834,N_29967);
or UO_905 (O_905,N_29521,N_29618);
or UO_906 (O_906,N_29424,N_29994);
xor UO_907 (O_907,N_29561,N_29408);
nand UO_908 (O_908,N_29686,N_29621);
or UO_909 (O_909,N_29517,N_29605);
nor UO_910 (O_910,N_29563,N_29989);
nor UO_911 (O_911,N_29981,N_29824);
nand UO_912 (O_912,N_29672,N_29542);
nor UO_913 (O_913,N_29905,N_29506);
xor UO_914 (O_914,N_29754,N_29637);
nor UO_915 (O_915,N_29532,N_29920);
xor UO_916 (O_916,N_29498,N_29964);
nand UO_917 (O_917,N_29668,N_29422);
and UO_918 (O_918,N_29842,N_29983);
nor UO_919 (O_919,N_29913,N_29997);
or UO_920 (O_920,N_29571,N_29428);
nor UO_921 (O_921,N_29998,N_29418);
xnor UO_922 (O_922,N_29565,N_29615);
nor UO_923 (O_923,N_29565,N_29808);
nor UO_924 (O_924,N_29927,N_29987);
xor UO_925 (O_925,N_29954,N_29617);
xnor UO_926 (O_926,N_29717,N_29821);
and UO_927 (O_927,N_29457,N_29965);
nand UO_928 (O_928,N_29775,N_29891);
nor UO_929 (O_929,N_29839,N_29479);
nand UO_930 (O_930,N_29602,N_29695);
xnor UO_931 (O_931,N_29597,N_29537);
xnor UO_932 (O_932,N_29575,N_29517);
xnor UO_933 (O_933,N_29641,N_29600);
xor UO_934 (O_934,N_29581,N_29876);
nand UO_935 (O_935,N_29930,N_29788);
or UO_936 (O_936,N_29493,N_29926);
or UO_937 (O_937,N_29472,N_29760);
xnor UO_938 (O_938,N_29560,N_29406);
nor UO_939 (O_939,N_29740,N_29651);
nand UO_940 (O_940,N_29887,N_29452);
xor UO_941 (O_941,N_29988,N_29536);
nand UO_942 (O_942,N_29994,N_29747);
and UO_943 (O_943,N_29944,N_29765);
or UO_944 (O_944,N_29710,N_29999);
nand UO_945 (O_945,N_29945,N_29766);
or UO_946 (O_946,N_29902,N_29876);
or UO_947 (O_947,N_29498,N_29755);
and UO_948 (O_948,N_29522,N_29618);
nand UO_949 (O_949,N_29943,N_29882);
xor UO_950 (O_950,N_29665,N_29588);
nand UO_951 (O_951,N_29719,N_29530);
nand UO_952 (O_952,N_29426,N_29782);
or UO_953 (O_953,N_29625,N_29503);
or UO_954 (O_954,N_29628,N_29419);
nand UO_955 (O_955,N_29997,N_29583);
nand UO_956 (O_956,N_29755,N_29697);
and UO_957 (O_957,N_29785,N_29551);
and UO_958 (O_958,N_29533,N_29435);
nor UO_959 (O_959,N_29727,N_29512);
nor UO_960 (O_960,N_29638,N_29433);
nor UO_961 (O_961,N_29998,N_29883);
and UO_962 (O_962,N_29666,N_29409);
and UO_963 (O_963,N_29683,N_29641);
nand UO_964 (O_964,N_29420,N_29688);
nand UO_965 (O_965,N_29788,N_29421);
xor UO_966 (O_966,N_29601,N_29824);
xor UO_967 (O_967,N_29694,N_29417);
xor UO_968 (O_968,N_29983,N_29760);
and UO_969 (O_969,N_29470,N_29763);
or UO_970 (O_970,N_29643,N_29513);
or UO_971 (O_971,N_29632,N_29648);
xor UO_972 (O_972,N_29615,N_29961);
xor UO_973 (O_973,N_29869,N_29501);
and UO_974 (O_974,N_29902,N_29654);
nor UO_975 (O_975,N_29438,N_29755);
nor UO_976 (O_976,N_29732,N_29758);
nand UO_977 (O_977,N_29467,N_29516);
nand UO_978 (O_978,N_29460,N_29982);
nand UO_979 (O_979,N_29555,N_29528);
and UO_980 (O_980,N_29479,N_29409);
nand UO_981 (O_981,N_29627,N_29972);
xnor UO_982 (O_982,N_29417,N_29666);
nor UO_983 (O_983,N_29495,N_29561);
xor UO_984 (O_984,N_29796,N_29814);
and UO_985 (O_985,N_29732,N_29869);
and UO_986 (O_986,N_29680,N_29988);
or UO_987 (O_987,N_29653,N_29880);
xnor UO_988 (O_988,N_29896,N_29430);
nor UO_989 (O_989,N_29491,N_29616);
nor UO_990 (O_990,N_29741,N_29527);
nor UO_991 (O_991,N_29919,N_29667);
and UO_992 (O_992,N_29504,N_29861);
and UO_993 (O_993,N_29666,N_29807);
nand UO_994 (O_994,N_29676,N_29648);
xor UO_995 (O_995,N_29934,N_29928);
nor UO_996 (O_996,N_29736,N_29565);
and UO_997 (O_997,N_29739,N_29832);
nor UO_998 (O_998,N_29773,N_29463);
and UO_999 (O_999,N_29409,N_29638);
nand UO_1000 (O_1000,N_29501,N_29403);
and UO_1001 (O_1001,N_29572,N_29882);
or UO_1002 (O_1002,N_29531,N_29949);
nand UO_1003 (O_1003,N_29732,N_29568);
nor UO_1004 (O_1004,N_29520,N_29454);
and UO_1005 (O_1005,N_29430,N_29780);
xor UO_1006 (O_1006,N_29943,N_29552);
xnor UO_1007 (O_1007,N_29762,N_29855);
and UO_1008 (O_1008,N_29730,N_29613);
nor UO_1009 (O_1009,N_29534,N_29855);
xor UO_1010 (O_1010,N_29774,N_29651);
nor UO_1011 (O_1011,N_29459,N_29836);
xnor UO_1012 (O_1012,N_29783,N_29764);
nor UO_1013 (O_1013,N_29587,N_29565);
and UO_1014 (O_1014,N_29428,N_29420);
xnor UO_1015 (O_1015,N_29806,N_29401);
and UO_1016 (O_1016,N_29459,N_29569);
nand UO_1017 (O_1017,N_29673,N_29722);
nor UO_1018 (O_1018,N_29896,N_29989);
and UO_1019 (O_1019,N_29558,N_29408);
xnor UO_1020 (O_1020,N_29412,N_29595);
nand UO_1021 (O_1021,N_29555,N_29816);
xnor UO_1022 (O_1022,N_29430,N_29957);
or UO_1023 (O_1023,N_29920,N_29657);
or UO_1024 (O_1024,N_29440,N_29478);
nor UO_1025 (O_1025,N_29733,N_29518);
nand UO_1026 (O_1026,N_29701,N_29912);
or UO_1027 (O_1027,N_29967,N_29503);
nor UO_1028 (O_1028,N_29607,N_29413);
or UO_1029 (O_1029,N_29691,N_29972);
or UO_1030 (O_1030,N_29930,N_29897);
nand UO_1031 (O_1031,N_29943,N_29783);
xnor UO_1032 (O_1032,N_29781,N_29859);
nor UO_1033 (O_1033,N_29655,N_29851);
xor UO_1034 (O_1034,N_29902,N_29669);
and UO_1035 (O_1035,N_29945,N_29619);
and UO_1036 (O_1036,N_29934,N_29958);
and UO_1037 (O_1037,N_29565,N_29483);
nand UO_1038 (O_1038,N_29761,N_29556);
xnor UO_1039 (O_1039,N_29869,N_29635);
and UO_1040 (O_1040,N_29576,N_29506);
nand UO_1041 (O_1041,N_29932,N_29647);
or UO_1042 (O_1042,N_29721,N_29628);
or UO_1043 (O_1043,N_29930,N_29799);
and UO_1044 (O_1044,N_29611,N_29837);
nand UO_1045 (O_1045,N_29900,N_29569);
or UO_1046 (O_1046,N_29593,N_29959);
and UO_1047 (O_1047,N_29426,N_29939);
nand UO_1048 (O_1048,N_29475,N_29620);
xor UO_1049 (O_1049,N_29978,N_29842);
and UO_1050 (O_1050,N_29763,N_29753);
xor UO_1051 (O_1051,N_29777,N_29904);
nor UO_1052 (O_1052,N_29531,N_29843);
and UO_1053 (O_1053,N_29767,N_29545);
nand UO_1054 (O_1054,N_29886,N_29949);
or UO_1055 (O_1055,N_29863,N_29417);
and UO_1056 (O_1056,N_29605,N_29981);
xor UO_1057 (O_1057,N_29944,N_29919);
nand UO_1058 (O_1058,N_29459,N_29993);
or UO_1059 (O_1059,N_29630,N_29900);
and UO_1060 (O_1060,N_29848,N_29782);
nand UO_1061 (O_1061,N_29495,N_29505);
xnor UO_1062 (O_1062,N_29530,N_29961);
or UO_1063 (O_1063,N_29567,N_29698);
nand UO_1064 (O_1064,N_29958,N_29914);
nor UO_1065 (O_1065,N_29472,N_29593);
and UO_1066 (O_1066,N_29658,N_29786);
xnor UO_1067 (O_1067,N_29567,N_29520);
or UO_1068 (O_1068,N_29576,N_29815);
nor UO_1069 (O_1069,N_29937,N_29544);
nor UO_1070 (O_1070,N_29486,N_29902);
nor UO_1071 (O_1071,N_29905,N_29818);
nand UO_1072 (O_1072,N_29683,N_29484);
nor UO_1073 (O_1073,N_29434,N_29419);
nor UO_1074 (O_1074,N_29812,N_29585);
xor UO_1075 (O_1075,N_29431,N_29999);
and UO_1076 (O_1076,N_29428,N_29790);
nor UO_1077 (O_1077,N_29455,N_29752);
and UO_1078 (O_1078,N_29924,N_29491);
xnor UO_1079 (O_1079,N_29820,N_29446);
xor UO_1080 (O_1080,N_29951,N_29862);
nand UO_1081 (O_1081,N_29408,N_29993);
xor UO_1082 (O_1082,N_29502,N_29414);
xor UO_1083 (O_1083,N_29790,N_29837);
nor UO_1084 (O_1084,N_29735,N_29641);
nand UO_1085 (O_1085,N_29772,N_29991);
and UO_1086 (O_1086,N_29655,N_29635);
or UO_1087 (O_1087,N_29711,N_29527);
nand UO_1088 (O_1088,N_29962,N_29605);
and UO_1089 (O_1089,N_29977,N_29641);
and UO_1090 (O_1090,N_29822,N_29730);
nor UO_1091 (O_1091,N_29528,N_29901);
nand UO_1092 (O_1092,N_29526,N_29654);
nor UO_1093 (O_1093,N_29618,N_29979);
or UO_1094 (O_1094,N_29659,N_29472);
nand UO_1095 (O_1095,N_29971,N_29419);
xnor UO_1096 (O_1096,N_29488,N_29571);
nor UO_1097 (O_1097,N_29557,N_29544);
and UO_1098 (O_1098,N_29826,N_29788);
xnor UO_1099 (O_1099,N_29540,N_29928);
xor UO_1100 (O_1100,N_29962,N_29413);
or UO_1101 (O_1101,N_29657,N_29711);
xnor UO_1102 (O_1102,N_29548,N_29912);
and UO_1103 (O_1103,N_29836,N_29902);
nor UO_1104 (O_1104,N_29992,N_29898);
xor UO_1105 (O_1105,N_29627,N_29656);
xor UO_1106 (O_1106,N_29563,N_29713);
xnor UO_1107 (O_1107,N_29562,N_29855);
nor UO_1108 (O_1108,N_29925,N_29465);
nor UO_1109 (O_1109,N_29579,N_29983);
or UO_1110 (O_1110,N_29624,N_29701);
nand UO_1111 (O_1111,N_29766,N_29410);
nand UO_1112 (O_1112,N_29617,N_29696);
or UO_1113 (O_1113,N_29473,N_29996);
nand UO_1114 (O_1114,N_29993,N_29628);
and UO_1115 (O_1115,N_29749,N_29849);
or UO_1116 (O_1116,N_29445,N_29801);
or UO_1117 (O_1117,N_29723,N_29470);
or UO_1118 (O_1118,N_29938,N_29656);
xnor UO_1119 (O_1119,N_29527,N_29686);
or UO_1120 (O_1120,N_29806,N_29681);
and UO_1121 (O_1121,N_29883,N_29427);
nand UO_1122 (O_1122,N_29573,N_29741);
and UO_1123 (O_1123,N_29513,N_29633);
xnor UO_1124 (O_1124,N_29974,N_29512);
nand UO_1125 (O_1125,N_29407,N_29750);
or UO_1126 (O_1126,N_29792,N_29657);
xnor UO_1127 (O_1127,N_29900,N_29679);
nor UO_1128 (O_1128,N_29614,N_29986);
xor UO_1129 (O_1129,N_29531,N_29862);
xnor UO_1130 (O_1130,N_29523,N_29864);
and UO_1131 (O_1131,N_29689,N_29667);
nor UO_1132 (O_1132,N_29716,N_29669);
nor UO_1133 (O_1133,N_29721,N_29896);
or UO_1134 (O_1134,N_29892,N_29585);
and UO_1135 (O_1135,N_29529,N_29720);
or UO_1136 (O_1136,N_29918,N_29745);
nand UO_1137 (O_1137,N_29934,N_29887);
nand UO_1138 (O_1138,N_29993,N_29883);
or UO_1139 (O_1139,N_29923,N_29907);
and UO_1140 (O_1140,N_29489,N_29849);
and UO_1141 (O_1141,N_29920,N_29400);
nor UO_1142 (O_1142,N_29579,N_29832);
and UO_1143 (O_1143,N_29480,N_29711);
nand UO_1144 (O_1144,N_29406,N_29604);
or UO_1145 (O_1145,N_29671,N_29850);
or UO_1146 (O_1146,N_29712,N_29940);
xnor UO_1147 (O_1147,N_29857,N_29865);
or UO_1148 (O_1148,N_29948,N_29430);
or UO_1149 (O_1149,N_29523,N_29949);
nor UO_1150 (O_1150,N_29806,N_29921);
nor UO_1151 (O_1151,N_29477,N_29873);
xor UO_1152 (O_1152,N_29494,N_29807);
or UO_1153 (O_1153,N_29754,N_29532);
nor UO_1154 (O_1154,N_29420,N_29925);
nor UO_1155 (O_1155,N_29561,N_29627);
or UO_1156 (O_1156,N_29672,N_29818);
nand UO_1157 (O_1157,N_29720,N_29816);
nand UO_1158 (O_1158,N_29866,N_29618);
nand UO_1159 (O_1159,N_29929,N_29427);
xor UO_1160 (O_1160,N_29851,N_29471);
and UO_1161 (O_1161,N_29604,N_29796);
or UO_1162 (O_1162,N_29947,N_29678);
xnor UO_1163 (O_1163,N_29667,N_29441);
xnor UO_1164 (O_1164,N_29894,N_29745);
xnor UO_1165 (O_1165,N_29746,N_29671);
nor UO_1166 (O_1166,N_29844,N_29657);
nor UO_1167 (O_1167,N_29488,N_29742);
nor UO_1168 (O_1168,N_29782,N_29726);
nand UO_1169 (O_1169,N_29798,N_29897);
or UO_1170 (O_1170,N_29585,N_29803);
nor UO_1171 (O_1171,N_29759,N_29479);
or UO_1172 (O_1172,N_29706,N_29406);
xnor UO_1173 (O_1173,N_29881,N_29671);
nand UO_1174 (O_1174,N_29864,N_29551);
xor UO_1175 (O_1175,N_29450,N_29616);
nand UO_1176 (O_1176,N_29400,N_29528);
and UO_1177 (O_1177,N_29642,N_29939);
nand UO_1178 (O_1178,N_29850,N_29498);
or UO_1179 (O_1179,N_29496,N_29696);
nand UO_1180 (O_1180,N_29418,N_29518);
xnor UO_1181 (O_1181,N_29961,N_29601);
nor UO_1182 (O_1182,N_29833,N_29921);
or UO_1183 (O_1183,N_29680,N_29603);
and UO_1184 (O_1184,N_29570,N_29917);
xnor UO_1185 (O_1185,N_29684,N_29876);
nand UO_1186 (O_1186,N_29695,N_29829);
and UO_1187 (O_1187,N_29456,N_29475);
or UO_1188 (O_1188,N_29903,N_29621);
or UO_1189 (O_1189,N_29601,N_29548);
or UO_1190 (O_1190,N_29510,N_29646);
xor UO_1191 (O_1191,N_29904,N_29444);
nor UO_1192 (O_1192,N_29760,N_29801);
and UO_1193 (O_1193,N_29419,N_29672);
xor UO_1194 (O_1194,N_29900,N_29631);
xor UO_1195 (O_1195,N_29793,N_29510);
nor UO_1196 (O_1196,N_29583,N_29863);
nor UO_1197 (O_1197,N_29670,N_29920);
and UO_1198 (O_1198,N_29931,N_29452);
nor UO_1199 (O_1199,N_29925,N_29458);
nand UO_1200 (O_1200,N_29918,N_29822);
nor UO_1201 (O_1201,N_29750,N_29535);
or UO_1202 (O_1202,N_29852,N_29825);
nor UO_1203 (O_1203,N_29982,N_29958);
and UO_1204 (O_1204,N_29883,N_29932);
xor UO_1205 (O_1205,N_29864,N_29910);
and UO_1206 (O_1206,N_29713,N_29725);
nor UO_1207 (O_1207,N_29844,N_29559);
or UO_1208 (O_1208,N_29932,N_29896);
xor UO_1209 (O_1209,N_29486,N_29533);
nand UO_1210 (O_1210,N_29494,N_29818);
or UO_1211 (O_1211,N_29468,N_29655);
and UO_1212 (O_1212,N_29851,N_29880);
nand UO_1213 (O_1213,N_29459,N_29764);
nor UO_1214 (O_1214,N_29440,N_29514);
xor UO_1215 (O_1215,N_29656,N_29919);
or UO_1216 (O_1216,N_29446,N_29537);
and UO_1217 (O_1217,N_29463,N_29675);
and UO_1218 (O_1218,N_29777,N_29866);
and UO_1219 (O_1219,N_29534,N_29982);
or UO_1220 (O_1220,N_29916,N_29668);
or UO_1221 (O_1221,N_29899,N_29491);
xor UO_1222 (O_1222,N_29508,N_29663);
or UO_1223 (O_1223,N_29468,N_29525);
nand UO_1224 (O_1224,N_29965,N_29846);
xnor UO_1225 (O_1225,N_29478,N_29687);
and UO_1226 (O_1226,N_29418,N_29835);
nand UO_1227 (O_1227,N_29949,N_29481);
or UO_1228 (O_1228,N_29887,N_29454);
nor UO_1229 (O_1229,N_29762,N_29618);
or UO_1230 (O_1230,N_29854,N_29746);
nand UO_1231 (O_1231,N_29696,N_29753);
nor UO_1232 (O_1232,N_29921,N_29476);
nor UO_1233 (O_1233,N_29941,N_29822);
nor UO_1234 (O_1234,N_29541,N_29651);
and UO_1235 (O_1235,N_29951,N_29513);
nor UO_1236 (O_1236,N_29530,N_29914);
nor UO_1237 (O_1237,N_29923,N_29450);
xor UO_1238 (O_1238,N_29517,N_29953);
nand UO_1239 (O_1239,N_29654,N_29763);
or UO_1240 (O_1240,N_29884,N_29505);
nand UO_1241 (O_1241,N_29590,N_29705);
nand UO_1242 (O_1242,N_29641,N_29568);
and UO_1243 (O_1243,N_29948,N_29832);
nor UO_1244 (O_1244,N_29409,N_29576);
xor UO_1245 (O_1245,N_29425,N_29758);
or UO_1246 (O_1246,N_29582,N_29555);
xnor UO_1247 (O_1247,N_29565,N_29903);
xnor UO_1248 (O_1248,N_29733,N_29675);
nand UO_1249 (O_1249,N_29833,N_29892);
nor UO_1250 (O_1250,N_29539,N_29951);
or UO_1251 (O_1251,N_29728,N_29656);
nand UO_1252 (O_1252,N_29765,N_29472);
or UO_1253 (O_1253,N_29843,N_29863);
nor UO_1254 (O_1254,N_29622,N_29774);
xor UO_1255 (O_1255,N_29966,N_29680);
xor UO_1256 (O_1256,N_29767,N_29700);
nand UO_1257 (O_1257,N_29787,N_29603);
xor UO_1258 (O_1258,N_29555,N_29586);
and UO_1259 (O_1259,N_29566,N_29983);
nand UO_1260 (O_1260,N_29848,N_29886);
and UO_1261 (O_1261,N_29972,N_29522);
nor UO_1262 (O_1262,N_29830,N_29552);
or UO_1263 (O_1263,N_29802,N_29629);
and UO_1264 (O_1264,N_29478,N_29625);
nand UO_1265 (O_1265,N_29901,N_29426);
nor UO_1266 (O_1266,N_29450,N_29650);
or UO_1267 (O_1267,N_29858,N_29678);
and UO_1268 (O_1268,N_29423,N_29855);
xor UO_1269 (O_1269,N_29829,N_29781);
xnor UO_1270 (O_1270,N_29638,N_29541);
and UO_1271 (O_1271,N_29538,N_29808);
or UO_1272 (O_1272,N_29734,N_29776);
xnor UO_1273 (O_1273,N_29950,N_29975);
or UO_1274 (O_1274,N_29454,N_29756);
and UO_1275 (O_1275,N_29955,N_29538);
nand UO_1276 (O_1276,N_29586,N_29713);
nor UO_1277 (O_1277,N_29500,N_29608);
nand UO_1278 (O_1278,N_29433,N_29989);
and UO_1279 (O_1279,N_29576,N_29423);
nand UO_1280 (O_1280,N_29570,N_29838);
and UO_1281 (O_1281,N_29753,N_29793);
xnor UO_1282 (O_1282,N_29579,N_29934);
and UO_1283 (O_1283,N_29890,N_29753);
nor UO_1284 (O_1284,N_29521,N_29526);
or UO_1285 (O_1285,N_29795,N_29477);
and UO_1286 (O_1286,N_29686,N_29481);
and UO_1287 (O_1287,N_29806,N_29810);
xor UO_1288 (O_1288,N_29661,N_29443);
nand UO_1289 (O_1289,N_29731,N_29693);
nand UO_1290 (O_1290,N_29664,N_29864);
and UO_1291 (O_1291,N_29966,N_29639);
nor UO_1292 (O_1292,N_29906,N_29496);
nand UO_1293 (O_1293,N_29782,N_29906);
nor UO_1294 (O_1294,N_29682,N_29610);
nor UO_1295 (O_1295,N_29930,N_29821);
or UO_1296 (O_1296,N_29867,N_29493);
nor UO_1297 (O_1297,N_29529,N_29974);
and UO_1298 (O_1298,N_29723,N_29840);
or UO_1299 (O_1299,N_29607,N_29645);
nor UO_1300 (O_1300,N_29961,N_29780);
xor UO_1301 (O_1301,N_29586,N_29575);
and UO_1302 (O_1302,N_29417,N_29758);
nor UO_1303 (O_1303,N_29751,N_29626);
nor UO_1304 (O_1304,N_29825,N_29928);
xnor UO_1305 (O_1305,N_29707,N_29776);
nor UO_1306 (O_1306,N_29899,N_29678);
xor UO_1307 (O_1307,N_29953,N_29648);
or UO_1308 (O_1308,N_29445,N_29495);
or UO_1309 (O_1309,N_29771,N_29785);
or UO_1310 (O_1310,N_29448,N_29421);
or UO_1311 (O_1311,N_29518,N_29863);
and UO_1312 (O_1312,N_29726,N_29723);
xor UO_1313 (O_1313,N_29888,N_29854);
xnor UO_1314 (O_1314,N_29824,N_29771);
and UO_1315 (O_1315,N_29969,N_29731);
xnor UO_1316 (O_1316,N_29635,N_29800);
xor UO_1317 (O_1317,N_29753,N_29540);
and UO_1318 (O_1318,N_29573,N_29854);
xnor UO_1319 (O_1319,N_29884,N_29721);
or UO_1320 (O_1320,N_29435,N_29587);
or UO_1321 (O_1321,N_29787,N_29426);
and UO_1322 (O_1322,N_29853,N_29966);
nor UO_1323 (O_1323,N_29581,N_29597);
nand UO_1324 (O_1324,N_29590,N_29974);
nand UO_1325 (O_1325,N_29516,N_29479);
and UO_1326 (O_1326,N_29898,N_29427);
or UO_1327 (O_1327,N_29525,N_29711);
nor UO_1328 (O_1328,N_29557,N_29589);
nand UO_1329 (O_1329,N_29658,N_29777);
or UO_1330 (O_1330,N_29622,N_29452);
and UO_1331 (O_1331,N_29932,N_29776);
nand UO_1332 (O_1332,N_29835,N_29459);
and UO_1333 (O_1333,N_29629,N_29439);
and UO_1334 (O_1334,N_29431,N_29612);
or UO_1335 (O_1335,N_29691,N_29701);
nand UO_1336 (O_1336,N_29879,N_29597);
xnor UO_1337 (O_1337,N_29887,N_29808);
nand UO_1338 (O_1338,N_29662,N_29991);
and UO_1339 (O_1339,N_29809,N_29415);
xor UO_1340 (O_1340,N_29501,N_29975);
xor UO_1341 (O_1341,N_29462,N_29689);
or UO_1342 (O_1342,N_29971,N_29946);
or UO_1343 (O_1343,N_29650,N_29956);
and UO_1344 (O_1344,N_29792,N_29620);
nand UO_1345 (O_1345,N_29809,N_29834);
nor UO_1346 (O_1346,N_29481,N_29685);
or UO_1347 (O_1347,N_29481,N_29962);
nand UO_1348 (O_1348,N_29731,N_29644);
xnor UO_1349 (O_1349,N_29437,N_29937);
nor UO_1350 (O_1350,N_29702,N_29639);
or UO_1351 (O_1351,N_29881,N_29795);
nor UO_1352 (O_1352,N_29873,N_29808);
and UO_1353 (O_1353,N_29450,N_29439);
or UO_1354 (O_1354,N_29965,N_29565);
nor UO_1355 (O_1355,N_29576,N_29938);
and UO_1356 (O_1356,N_29995,N_29822);
and UO_1357 (O_1357,N_29730,N_29701);
nand UO_1358 (O_1358,N_29679,N_29922);
nand UO_1359 (O_1359,N_29420,N_29986);
nand UO_1360 (O_1360,N_29422,N_29759);
or UO_1361 (O_1361,N_29696,N_29538);
nor UO_1362 (O_1362,N_29651,N_29968);
or UO_1363 (O_1363,N_29486,N_29782);
xor UO_1364 (O_1364,N_29621,N_29504);
or UO_1365 (O_1365,N_29781,N_29896);
and UO_1366 (O_1366,N_29729,N_29985);
or UO_1367 (O_1367,N_29842,N_29609);
nor UO_1368 (O_1368,N_29516,N_29582);
or UO_1369 (O_1369,N_29705,N_29510);
and UO_1370 (O_1370,N_29495,N_29462);
and UO_1371 (O_1371,N_29949,N_29495);
or UO_1372 (O_1372,N_29429,N_29638);
nand UO_1373 (O_1373,N_29688,N_29884);
xor UO_1374 (O_1374,N_29624,N_29458);
xor UO_1375 (O_1375,N_29623,N_29962);
nand UO_1376 (O_1376,N_29835,N_29828);
or UO_1377 (O_1377,N_29839,N_29487);
xnor UO_1378 (O_1378,N_29435,N_29600);
nor UO_1379 (O_1379,N_29696,N_29527);
nand UO_1380 (O_1380,N_29500,N_29671);
nor UO_1381 (O_1381,N_29935,N_29854);
or UO_1382 (O_1382,N_29748,N_29571);
or UO_1383 (O_1383,N_29775,N_29941);
xnor UO_1384 (O_1384,N_29487,N_29845);
nand UO_1385 (O_1385,N_29402,N_29447);
nor UO_1386 (O_1386,N_29724,N_29596);
nor UO_1387 (O_1387,N_29451,N_29798);
nor UO_1388 (O_1388,N_29801,N_29728);
nand UO_1389 (O_1389,N_29852,N_29523);
nand UO_1390 (O_1390,N_29784,N_29705);
nand UO_1391 (O_1391,N_29655,N_29934);
or UO_1392 (O_1392,N_29860,N_29876);
and UO_1393 (O_1393,N_29820,N_29979);
xnor UO_1394 (O_1394,N_29927,N_29735);
or UO_1395 (O_1395,N_29481,N_29413);
nor UO_1396 (O_1396,N_29872,N_29518);
nand UO_1397 (O_1397,N_29941,N_29818);
and UO_1398 (O_1398,N_29981,N_29420);
nor UO_1399 (O_1399,N_29954,N_29407);
xor UO_1400 (O_1400,N_29617,N_29895);
xnor UO_1401 (O_1401,N_29506,N_29640);
nor UO_1402 (O_1402,N_29435,N_29791);
nor UO_1403 (O_1403,N_29444,N_29909);
nand UO_1404 (O_1404,N_29764,N_29465);
nor UO_1405 (O_1405,N_29567,N_29725);
and UO_1406 (O_1406,N_29993,N_29613);
nor UO_1407 (O_1407,N_29455,N_29804);
nor UO_1408 (O_1408,N_29576,N_29889);
nor UO_1409 (O_1409,N_29472,N_29877);
nor UO_1410 (O_1410,N_29454,N_29738);
and UO_1411 (O_1411,N_29563,N_29434);
nand UO_1412 (O_1412,N_29502,N_29671);
nor UO_1413 (O_1413,N_29489,N_29620);
xor UO_1414 (O_1414,N_29979,N_29450);
or UO_1415 (O_1415,N_29730,N_29987);
xor UO_1416 (O_1416,N_29408,N_29532);
or UO_1417 (O_1417,N_29861,N_29809);
xor UO_1418 (O_1418,N_29971,N_29736);
nor UO_1419 (O_1419,N_29523,N_29803);
nand UO_1420 (O_1420,N_29901,N_29563);
and UO_1421 (O_1421,N_29773,N_29571);
and UO_1422 (O_1422,N_29609,N_29884);
nand UO_1423 (O_1423,N_29969,N_29919);
and UO_1424 (O_1424,N_29400,N_29919);
nor UO_1425 (O_1425,N_29443,N_29971);
nor UO_1426 (O_1426,N_29483,N_29595);
or UO_1427 (O_1427,N_29542,N_29812);
xnor UO_1428 (O_1428,N_29783,N_29944);
or UO_1429 (O_1429,N_29693,N_29686);
and UO_1430 (O_1430,N_29838,N_29639);
or UO_1431 (O_1431,N_29697,N_29756);
or UO_1432 (O_1432,N_29629,N_29852);
or UO_1433 (O_1433,N_29622,N_29632);
and UO_1434 (O_1434,N_29694,N_29934);
or UO_1435 (O_1435,N_29659,N_29484);
or UO_1436 (O_1436,N_29912,N_29456);
xor UO_1437 (O_1437,N_29625,N_29529);
nor UO_1438 (O_1438,N_29551,N_29692);
nand UO_1439 (O_1439,N_29750,N_29723);
xor UO_1440 (O_1440,N_29623,N_29633);
xor UO_1441 (O_1441,N_29923,N_29502);
xor UO_1442 (O_1442,N_29914,N_29602);
nor UO_1443 (O_1443,N_29936,N_29597);
or UO_1444 (O_1444,N_29911,N_29687);
or UO_1445 (O_1445,N_29631,N_29484);
and UO_1446 (O_1446,N_29630,N_29853);
xor UO_1447 (O_1447,N_29656,N_29578);
nor UO_1448 (O_1448,N_29566,N_29602);
or UO_1449 (O_1449,N_29743,N_29819);
xor UO_1450 (O_1450,N_29400,N_29946);
nand UO_1451 (O_1451,N_29800,N_29806);
and UO_1452 (O_1452,N_29578,N_29707);
or UO_1453 (O_1453,N_29758,N_29400);
nor UO_1454 (O_1454,N_29526,N_29696);
nand UO_1455 (O_1455,N_29972,N_29784);
xnor UO_1456 (O_1456,N_29810,N_29666);
or UO_1457 (O_1457,N_29652,N_29475);
nand UO_1458 (O_1458,N_29529,N_29471);
xor UO_1459 (O_1459,N_29712,N_29937);
xor UO_1460 (O_1460,N_29571,N_29564);
or UO_1461 (O_1461,N_29845,N_29573);
xnor UO_1462 (O_1462,N_29717,N_29833);
nor UO_1463 (O_1463,N_29546,N_29498);
and UO_1464 (O_1464,N_29770,N_29969);
and UO_1465 (O_1465,N_29645,N_29598);
nor UO_1466 (O_1466,N_29624,N_29860);
xor UO_1467 (O_1467,N_29436,N_29748);
xor UO_1468 (O_1468,N_29910,N_29617);
or UO_1469 (O_1469,N_29961,N_29828);
nand UO_1470 (O_1470,N_29618,N_29421);
nand UO_1471 (O_1471,N_29456,N_29784);
nor UO_1472 (O_1472,N_29540,N_29462);
nor UO_1473 (O_1473,N_29943,N_29576);
xor UO_1474 (O_1474,N_29710,N_29581);
and UO_1475 (O_1475,N_29573,N_29655);
nand UO_1476 (O_1476,N_29632,N_29488);
and UO_1477 (O_1477,N_29907,N_29734);
and UO_1478 (O_1478,N_29550,N_29982);
xnor UO_1479 (O_1479,N_29922,N_29825);
nand UO_1480 (O_1480,N_29849,N_29827);
nor UO_1481 (O_1481,N_29814,N_29983);
and UO_1482 (O_1482,N_29701,N_29464);
nor UO_1483 (O_1483,N_29889,N_29623);
nand UO_1484 (O_1484,N_29547,N_29830);
or UO_1485 (O_1485,N_29521,N_29848);
xor UO_1486 (O_1486,N_29651,N_29755);
nor UO_1487 (O_1487,N_29788,N_29669);
and UO_1488 (O_1488,N_29885,N_29788);
or UO_1489 (O_1489,N_29522,N_29998);
or UO_1490 (O_1490,N_29872,N_29997);
and UO_1491 (O_1491,N_29881,N_29928);
nor UO_1492 (O_1492,N_29842,N_29471);
xnor UO_1493 (O_1493,N_29551,N_29437);
xnor UO_1494 (O_1494,N_29451,N_29742);
nand UO_1495 (O_1495,N_29412,N_29797);
or UO_1496 (O_1496,N_29761,N_29736);
xor UO_1497 (O_1497,N_29571,N_29708);
nand UO_1498 (O_1498,N_29855,N_29403);
or UO_1499 (O_1499,N_29766,N_29954);
xor UO_1500 (O_1500,N_29778,N_29957);
or UO_1501 (O_1501,N_29891,N_29847);
xor UO_1502 (O_1502,N_29943,N_29444);
or UO_1503 (O_1503,N_29693,N_29547);
or UO_1504 (O_1504,N_29758,N_29959);
nor UO_1505 (O_1505,N_29520,N_29614);
and UO_1506 (O_1506,N_29667,N_29516);
or UO_1507 (O_1507,N_29753,N_29940);
nor UO_1508 (O_1508,N_29664,N_29658);
and UO_1509 (O_1509,N_29509,N_29581);
or UO_1510 (O_1510,N_29563,N_29893);
nand UO_1511 (O_1511,N_29508,N_29758);
and UO_1512 (O_1512,N_29692,N_29655);
and UO_1513 (O_1513,N_29769,N_29606);
nor UO_1514 (O_1514,N_29729,N_29617);
or UO_1515 (O_1515,N_29892,N_29775);
or UO_1516 (O_1516,N_29879,N_29808);
nand UO_1517 (O_1517,N_29889,N_29613);
and UO_1518 (O_1518,N_29484,N_29497);
nand UO_1519 (O_1519,N_29450,N_29491);
nand UO_1520 (O_1520,N_29799,N_29516);
or UO_1521 (O_1521,N_29797,N_29854);
xor UO_1522 (O_1522,N_29563,N_29749);
nand UO_1523 (O_1523,N_29629,N_29732);
nand UO_1524 (O_1524,N_29791,N_29610);
xnor UO_1525 (O_1525,N_29959,N_29454);
nand UO_1526 (O_1526,N_29905,N_29467);
and UO_1527 (O_1527,N_29870,N_29976);
and UO_1528 (O_1528,N_29546,N_29635);
xor UO_1529 (O_1529,N_29808,N_29914);
nand UO_1530 (O_1530,N_29605,N_29651);
and UO_1531 (O_1531,N_29703,N_29740);
or UO_1532 (O_1532,N_29499,N_29568);
nor UO_1533 (O_1533,N_29840,N_29836);
or UO_1534 (O_1534,N_29486,N_29824);
xnor UO_1535 (O_1535,N_29967,N_29456);
and UO_1536 (O_1536,N_29813,N_29594);
or UO_1537 (O_1537,N_29512,N_29503);
nand UO_1538 (O_1538,N_29612,N_29858);
xor UO_1539 (O_1539,N_29610,N_29654);
or UO_1540 (O_1540,N_29870,N_29737);
nand UO_1541 (O_1541,N_29876,N_29641);
or UO_1542 (O_1542,N_29973,N_29857);
nor UO_1543 (O_1543,N_29824,N_29712);
or UO_1544 (O_1544,N_29936,N_29926);
and UO_1545 (O_1545,N_29644,N_29886);
or UO_1546 (O_1546,N_29959,N_29644);
or UO_1547 (O_1547,N_29773,N_29578);
and UO_1548 (O_1548,N_29544,N_29407);
or UO_1549 (O_1549,N_29987,N_29716);
nand UO_1550 (O_1550,N_29895,N_29851);
xnor UO_1551 (O_1551,N_29651,N_29463);
nor UO_1552 (O_1552,N_29974,N_29908);
nand UO_1553 (O_1553,N_29526,N_29582);
and UO_1554 (O_1554,N_29765,N_29959);
or UO_1555 (O_1555,N_29943,N_29707);
xnor UO_1556 (O_1556,N_29854,N_29842);
or UO_1557 (O_1557,N_29981,N_29566);
xnor UO_1558 (O_1558,N_29448,N_29953);
or UO_1559 (O_1559,N_29722,N_29609);
nor UO_1560 (O_1560,N_29870,N_29532);
xnor UO_1561 (O_1561,N_29717,N_29506);
nand UO_1562 (O_1562,N_29787,N_29860);
and UO_1563 (O_1563,N_29419,N_29939);
and UO_1564 (O_1564,N_29819,N_29600);
and UO_1565 (O_1565,N_29885,N_29964);
nor UO_1566 (O_1566,N_29613,N_29946);
nor UO_1567 (O_1567,N_29854,N_29973);
and UO_1568 (O_1568,N_29775,N_29676);
xor UO_1569 (O_1569,N_29458,N_29674);
or UO_1570 (O_1570,N_29489,N_29407);
and UO_1571 (O_1571,N_29654,N_29977);
xor UO_1572 (O_1572,N_29889,N_29504);
xnor UO_1573 (O_1573,N_29541,N_29587);
and UO_1574 (O_1574,N_29913,N_29714);
nor UO_1575 (O_1575,N_29665,N_29525);
nand UO_1576 (O_1576,N_29612,N_29693);
nand UO_1577 (O_1577,N_29879,N_29489);
nor UO_1578 (O_1578,N_29456,N_29811);
nor UO_1579 (O_1579,N_29603,N_29402);
or UO_1580 (O_1580,N_29990,N_29475);
or UO_1581 (O_1581,N_29445,N_29481);
xor UO_1582 (O_1582,N_29556,N_29679);
xnor UO_1583 (O_1583,N_29868,N_29648);
nand UO_1584 (O_1584,N_29740,N_29734);
nand UO_1585 (O_1585,N_29793,N_29913);
nand UO_1586 (O_1586,N_29926,N_29684);
nor UO_1587 (O_1587,N_29769,N_29812);
nand UO_1588 (O_1588,N_29514,N_29867);
xnor UO_1589 (O_1589,N_29993,N_29423);
and UO_1590 (O_1590,N_29441,N_29588);
nor UO_1591 (O_1591,N_29439,N_29611);
nor UO_1592 (O_1592,N_29946,N_29872);
xor UO_1593 (O_1593,N_29773,N_29897);
nor UO_1594 (O_1594,N_29917,N_29539);
or UO_1595 (O_1595,N_29864,N_29979);
nor UO_1596 (O_1596,N_29673,N_29845);
xnor UO_1597 (O_1597,N_29533,N_29495);
or UO_1598 (O_1598,N_29481,N_29616);
or UO_1599 (O_1599,N_29707,N_29949);
or UO_1600 (O_1600,N_29582,N_29427);
xnor UO_1601 (O_1601,N_29574,N_29699);
xor UO_1602 (O_1602,N_29483,N_29931);
xor UO_1603 (O_1603,N_29666,N_29575);
nor UO_1604 (O_1604,N_29689,N_29565);
nor UO_1605 (O_1605,N_29555,N_29804);
nor UO_1606 (O_1606,N_29401,N_29496);
xor UO_1607 (O_1607,N_29976,N_29759);
xor UO_1608 (O_1608,N_29601,N_29633);
and UO_1609 (O_1609,N_29553,N_29655);
and UO_1610 (O_1610,N_29483,N_29991);
nor UO_1611 (O_1611,N_29409,N_29668);
nor UO_1612 (O_1612,N_29951,N_29901);
or UO_1613 (O_1613,N_29835,N_29856);
nand UO_1614 (O_1614,N_29968,N_29613);
nor UO_1615 (O_1615,N_29546,N_29643);
xor UO_1616 (O_1616,N_29594,N_29827);
nand UO_1617 (O_1617,N_29485,N_29823);
nand UO_1618 (O_1618,N_29413,N_29887);
nor UO_1619 (O_1619,N_29759,N_29409);
nor UO_1620 (O_1620,N_29469,N_29787);
xnor UO_1621 (O_1621,N_29509,N_29745);
nand UO_1622 (O_1622,N_29766,N_29438);
or UO_1623 (O_1623,N_29974,N_29539);
xnor UO_1624 (O_1624,N_29716,N_29770);
nand UO_1625 (O_1625,N_29497,N_29562);
xor UO_1626 (O_1626,N_29567,N_29587);
and UO_1627 (O_1627,N_29646,N_29647);
or UO_1628 (O_1628,N_29806,N_29718);
or UO_1629 (O_1629,N_29472,N_29782);
or UO_1630 (O_1630,N_29453,N_29997);
xor UO_1631 (O_1631,N_29928,N_29458);
nor UO_1632 (O_1632,N_29788,N_29658);
nand UO_1633 (O_1633,N_29602,N_29423);
and UO_1634 (O_1634,N_29579,N_29576);
and UO_1635 (O_1635,N_29481,N_29410);
nor UO_1636 (O_1636,N_29860,N_29952);
or UO_1637 (O_1637,N_29585,N_29935);
xnor UO_1638 (O_1638,N_29521,N_29495);
or UO_1639 (O_1639,N_29892,N_29802);
xnor UO_1640 (O_1640,N_29842,N_29443);
xor UO_1641 (O_1641,N_29911,N_29719);
nor UO_1642 (O_1642,N_29954,N_29468);
or UO_1643 (O_1643,N_29965,N_29722);
and UO_1644 (O_1644,N_29691,N_29682);
and UO_1645 (O_1645,N_29849,N_29485);
xnor UO_1646 (O_1646,N_29708,N_29432);
or UO_1647 (O_1647,N_29509,N_29506);
nand UO_1648 (O_1648,N_29707,N_29950);
nor UO_1649 (O_1649,N_29889,N_29622);
nand UO_1650 (O_1650,N_29521,N_29884);
nor UO_1651 (O_1651,N_29472,N_29750);
and UO_1652 (O_1652,N_29520,N_29694);
xnor UO_1653 (O_1653,N_29957,N_29879);
and UO_1654 (O_1654,N_29901,N_29681);
nand UO_1655 (O_1655,N_29432,N_29970);
and UO_1656 (O_1656,N_29881,N_29554);
nand UO_1657 (O_1657,N_29578,N_29923);
nand UO_1658 (O_1658,N_29756,N_29469);
nor UO_1659 (O_1659,N_29879,N_29826);
nand UO_1660 (O_1660,N_29954,N_29859);
or UO_1661 (O_1661,N_29592,N_29617);
or UO_1662 (O_1662,N_29517,N_29813);
and UO_1663 (O_1663,N_29913,N_29454);
nand UO_1664 (O_1664,N_29413,N_29843);
nand UO_1665 (O_1665,N_29411,N_29595);
xor UO_1666 (O_1666,N_29536,N_29727);
xor UO_1667 (O_1667,N_29595,N_29928);
or UO_1668 (O_1668,N_29671,N_29889);
nand UO_1669 (O_1669,N_29458,N_29537);
and UO_1670 (O_1670,N_29503,N_29862);
nand UO_1671 (O_1671,N_29463,N_29797);
nor UO_1672 (O_1672,N_29813,N_29754);
nor UO_1673 (O_1673,N_29909,N_29680);
or UO_1674 (O_1674,N_29980,N_29650);
nor UO_1675 (O_1675,N_29818,N_29536);
xnor UO_1676 (O_1676,N_29928,N_29471);
or UO_1677 (O_1677,N_29875,N_29930);
nor UO_1678 (O_1678,N_29610,N_29816);
or UO_1679 (O_1679,N_29507,N_29466);
nor UO_1680 (O_1680,N_29971,N_29854);
xor UO_1681 (O_1681,N_29531,N_29639);
and UO_1682 (O_1682,N_29686,N_29498);
and UO_1683 (O_1683,N_29855,N_29923);
nand UO_1684 (O_1684,N_29862,N_29494);
nor UO_1685 (O_1685,N_29622,N_29526);
or UO_1686 (O_1686,N_29941,N_29907);
nor UO_1687 (O_1687,N_29862,N_29468);
or UO_1688 (O_1688,N_29824,N_29986);
xor UO_1689 (O_1689,N_29471,N_29468);
xnor UO_1690 (O_1690,N_29697,N_29803);
xor UO_1691 (O_1691,N_29917,N_29953);
nand UO_1692 (O_1692,N_29903,N_29940);
xnor UO_1693 (O_1693,N_29776,N_29720);
or UO_1694 (O_1694,N_29898,N_29655);
xnor UO_1695 (O_1695,N_29990,N_29532);
or UO_1696 (O_1696,N_29450,N_29882);
nor UO_1697 (O_1697,N_29993,N_29692);
or UO_1698 (O_1698,N_29763,N_29716);
and UO_1699 (O_1699,N_29781,N_29897);
nand UO_1700 (O_1700,N_29615,N_29696);
nand UO_1701 (O_1701,N_29421,N_29936);
nand UO_1702 (O_1702,N_29901,N_29465);
or UO_1703 (O_1703,N_29801,N_29455);
and UO_1704 (O_1704,N_29876,N_29637);
and UO_1705 (O_1705,N_29514,N_29818);
or UO_1706 (O_1706,N_29664,N_29981);
nand UO_1707 (O_1707,N_29780,N_29840);
nor UO_1708 (O_1708,N_29917,N_29754);
xor UO_1709 (O_1709,N_29989,N_29684);
nand UO_1710 (O_1710,N_29426,N_29822);
xor UO_1711 (O_1711,N_29930,N_29611);
nor UO_1712 (O_1712,N_29681,N_29663);
nor UO_1713 (O_1713,N_29838,N_29449);
nor UO_1714 (O_1714,N_29973,N_29813);
nand UO_1715 (O_1715,N_29476,N_29528);
xor UO_1716 (O_1716,N_29807,N_29957);
nor UO_1717 (O_1717,N_29409,N_29606);
and UO_1718 (O_1718,N_29834,N_29772);
and UO_1719 (O_1719,N_29861,N_29746);
xor UO_1720 (O_1720,N_29847,N_29692);
and UO_1721 (O_1721,N_29634,N_29688);
or UO_1722 (O_1722,N_29490,N_29806);
and UO_1723 (O_1723,N_29678,N_29747);
and UO_1724 (O_1724,N_29693,N_29649);
xor UO_1725 (O_1725,N_29805,N_29637);
xnor UO_1726 (O_1726,N_29561,N_29968);
nand UO_1727 (O_1727,N_29459,N_29945);
or UO_1728 (O_1728,N_29697,N_29591);
and UO_1729 (O_1729,N_29438,N_29510);
nor UO_1730 (O_1730,N_29911,N_29980);
nand UO_1731 (O_1731,N_29966,N_29819);
nand UO_1732 (O_1732,N_29940,N_29533);
or UO_1733 (O_1733,N_29558,N_29653);
or UO_1734 (O_1734,N_29400,N_29974);
or UO_1735 (O_1735,N_29805,N_29961);
or UO_1736 (O_1736,N_29854,N_29711);
nand UO_1737 (O_1737,N_29800,N_29501);
or UO_1738 (O_1738,N_29435,N_29680);
nor UO_1739 (O_1739,N_29979,N_29749);
and UO_1740 (O_1740,N_29864,N_29706);
and UO_1741 (O_1741,N_29903,N_29547);
nor UO_1742 (O_1742,N_29870,N_29491);
xor UO_1743 (O_1743,N_29722,N_29978);
and UO_1744 (O_1744,N_29448,N_29404);
nand UO_1745 (O_1745,N_29577,N_29797);
nor UO_1746 (O_1746,N_29659,N_29863);
nand UO_1747 (O_1747,N_29486,N_29630);
or UO_1748 (O_1748,N_29810,N_29554);
nand UO_1749 (O_1749,N_29450,N_29821);
and UO_1750 (O_1750,N_29448,N_29944);
or UO_1751 (O_1751,N_29518,N_29612);
xor UO_1752 (O_1752,N_29607,N_29926);
and UO_1753 (O_1753,N_29880,N_29789);
xor UO_1754 (O_1754,N_29851,N_29454);
or UO_1755 (O_1755,N_29441,N_29821);
xor UO_1756 (O_1756,N_29786,N_29660);
xor UO_1757 (O_1757,N_29581,N_29939);
and UO_1758 (O_1758,N_29532,N_29734);
nor UO_1759 (O_1759,N_29441,N_29636);
nor UO_1760 (O_1760,N_29785,N_29596);
and UO_1761 (O_1761,N_29991,N_29621);
nand UO_1762 (O_1762,N_29613,N_29915);
xnor UO_1763 (O_1763,N_29765,N_29630);
nand UO_1764 (O_1764,N_29513,N_29728);
nor UO_1765 (O_1765,N_29645,N_29430);
and UO_1766 (O_1766,N_29993,N_29543);
nand UO_1767 (O_1767,N_29666,N_29608);
and UO_1768 (O_1768,N_29816,N_29566);
nand UO_1769 (O_1769,N_29651,N_29799);
nor UO_1770 (O_1770,N_29726,N_29714);
nand UO_1771 (O_1771,N_29694,N_29627);
xor UO_1772 (O_1772,N_29433,N_29464);
nand UO_1773 (O_1773,N_29452,N_29741);
and UO_1774 (O_1774,N_29511,N_29671);
and UO_1775 (O_1775,N_29515,N_29437);
nand UO_1776 (O_1776,N_29462,N_29466);
and UO_1777 (O_1777,N_29951,N_29762);
or UO_1778 (O_1778,N_29406,N_29516);
and UO_1779 (O_1779,N_29483,N_29772);
xnor UO_1780 (O_1780,N_29610,N_29493);
or UO_1781 (O_1781,N_29756,N_29945);
xor UO_1782 (O_1782,N_29480,N_29704);
or UO_1783 (O_1783,N_29500,N_29567);
and UO_1784 (O_1784,N_29806,N_29489);
and UO_1785 (O_1785,N_29987,N_29988);
or UO_1786 (O_1786,N_29642,N_29944);
nand UO_1787 (O_1787,N_29488,N_29675);
xor UO_1788 (O_1788,N_29887,N_29943);
xnor UO_1789 (O_1789,N_29725,N_29811);
nor UO_1790 (O_1790,N_29571,N_29904);
and UO_1791 (O_1791,N_29506,N_29885);
xor UO_1792 (O_1792,N_29469,N_29778);
and UO_1793 (O_1793,N_29766,N_29655);
xnor UO_1794 (O_1794,N_29464,N_29432);
or UO_1795 (O_1795,N_29439,N_29835);
nand UO_1796 (O_1796,N_29916,N_29710);
nand UO_1797 (O_1797,N_29985,N_29816);
nand UO_1798 (O_1798,N_29596,N_29892);
or UO_1799 (O_1799,N_29803,N_29591);
nor UO_1800 (O_1800,N_29921,N_29650);
or UO_1801 (O_1801,N_29877,N_29526);
or UO_1802 (O_1802,N_29741,N_29534);
and UO_1803 (O_1803,N_29452,N_29759);
xnor UO_1804 (O_1804,N_29816,N_29653);
and UO_1805 (O_1805,N_29487,N_29910);
xnor UO_1806 (O_1806,N_29664,N_29956);
nor UO_1807 (O_1807,N_29864,N_29856);
and UO_1808 (O_1808,N_29505,N_29453);
or UO_1809 (O_1809,N_29795,N_29525);
nor UO_1810 (O_1810,N_29600,N_29612);
and UO_1811 (O_1811,N_29729,N_29515);
and UO_1812 (O_1812,N_29606,N_29406);
nor UO_1813 (O_1813,N_29968,N_29582);
nand UO_1814 (O_1814,N_29952,N_29858);
and UO_1815 (O_1815,N_29622,N_29957);
xnor UO_1816 (O_1816,N_29501,N_29704);
or UO_1817 (O_1817,N_29747,N_29404);
xor UO_1818 (O_1818,N_29421,N_29585);
nand UO_1819 (O_1819,N_29774,N_29608);
and UO_1820 (O_1820,N_29608,N_29689);
nand UO_1821 (O_1821,N_29790,N_29804);
or UO_1822 (O_1822,N_29563,N_29789);
and UO_1823 (O_1823,N_29877,N_29554);
nand UO_1824 (O_1824,N_29676,N_29590);
nand UO_1825 (O_1825,N_29846,N_29614);
xor UO_1826 (O_1826,N_29562,N_29445);
nor UO_1827 (O_1827,N_29960,N_29499);
nor UO_1828 (O_1828,N_29490,N_29697);
xor UO_1829 (O_1829,N_29499,N_29489);
nor UO_1830 (O_1830,N_29923,N_29803);
nand UO_1831 (O_1831,N_29613,N_29950);
and UO_1832 (O_1832,N_29924,N_29445);
nand UO_1833 (O_1833,N_29950,N_29551);
nor UO_1834 (O_1834,N_29412,N_29553);
or UO_1835 (O_1835,N_29462,N_29812);
and UO_1836 (O_1836,N_29909,N_29668);
or UO_1837 (O_1837,N_29807,N_29896);
nor UO_1838 (O_1838,N_29940,N_29610);
and UO_1839 (O_1839,N_29829,N_29848);
or UO_1840 (O_1840,N_29538,N_29784);
or UO_1841 (O_1841,N_29744,N_29985);
nor UO_1842 (O_1842,N_29500,N_29967);
nand UO_1843 (O_1843,N_29487,N_29642);
nor UO_1844 (O_1844,N_29750,N_29518);
nor UO_1845 (O_1845,N_29834,N_29730);
and UO_1846 (O_1846,N_29914,N_29449);
or UO_1847 (O_1847,N_29997,N_29485);
and UO_1848 (O_1848,N_29894,N_29821);
xnor UO_1849 (O_1849,N_29754,N_29844);
xor UO_1850 (O_1850,N_29448,N_29812);
nand UO_1851 (O_1851,N_29596,N_29938);
xnor UO_1852 (O_1852,N_29775,N_29577);
and UO_1853 (O_1853,N_29607,N_29720);
nor UO_1854 (O_1854,N_29743,N_29891);
or UO_1855 (O_1855,N_29896,N_29569);
nor UO_1856 (O_1856,N_29666,N_29853);
and UO_1857 (O_1857,N_29756,N_29421);
nor UO_1858 (O_1858,N_29409,N_29500);
xnor UO_1859 (O_1859,N_29912,N_29550);
xor UO_1860 (O_1860,N_29705,N_29552);
and UO_1861 (O_1861,N_29937,N_29702);
or UO_1862 (O_1862,N_29858,N_29991);
xor UO_1863 (O_1863,N_29788,N_29740);
nor UO_1864 (O_1864,N_29670,N_29793);
xor UO_1865 (O_1865,N_29797,N_29409);
and UO_1866 (O_1866,N_29893,N_29469);
nand UO_1867 (O_1867,N_29412,N_29581);
nor UO_1868 (O_1868,N_29840,N_29963);
nor UO_1869 (O_1869,N_29757,N_29705);
and UO_1870 (O_1870,N_29584,N_29566);
and UO_1871 (O_1871,N_29602,N_29448);
nand UO_1872 (O_1872,N_29786,N_29669);
nand UO_1873 (O_1873,N_29612,N_29898);
or UO_1874 (O_1874,N_29537,N_29524);
or UO_1875 (O_1875,N_29598,N_29874);
and UO_1876 (O_1876,N_29951,N_29857);
and UO_1877 (O_1877,N_29648,N_29738);
or UO_1878 (O_1878,N_29724,N_29673);
and UO_1879 (O_1879,N_29735,N_29536);
nand UO_1880 (O_1880,N_29477,N_29741);
or UO_1881 (O_1881,N_29605,N_29558);
or UO_1882 (O_1882,N_29659,N_29993);
nand UO_1883 (O_1883,N_29674,N_29418);
nand UO_1884 (O_1884,N_29667,N_29970);
and UO_1885 (O_1885,N_29750,N_29739);
xor UO_1886 (O_1886,N_29859,N_29595);
or UO_1887 (O_1887,N_29464,N_29610);
xnor UO_1888 (O_1888,N_29554,N_29984);
or UO_1889 (O_1889,N_29439,N_29969);
and UO_1890 (O_1890,N_29820,N_29894);
xnor UO_1891 (O_1891,N_29640,N_29553);
nand UO_1892 (O_1892,N_29930,N_29437);
or UO_1893 (O_1893,N_29783,N_29733);
nor UO_1894 (O_1894,N_29468,N_29529);
nand UO_1895 (O_1895,N_29547,N_29796);
nor UO_1896 (O_1896,N_29659,N_29683);
xor UO_1897 (O_1897,N_29686,N_29891);
nor UO_1898 (O_1898,N_29674,N_29851);
xor UO_1899 (O_1899,N_29529,N_29962);
xor UO_1900 (O_1900,N_29930,N_29912);
nor UO_1901 (O_1901,N_29726,N_29931);
xnor UO_1902 (O_1902,N_29443,N_29917);
nand UO_1903 (O_1903,N_29777,N_29653);
nand UO_1904 (O_1904,N_29756,N_29845);
xnor UO_1905 (O_1905,N_29842,N_29637);
xnor UO_1906 (O_1906,N_29523,N_29584);
nor UO_1907 (O_1907,N_29471,N_29874);
or UO_1908 (O_1908,N_29918,N_29668);
or UO_1909 (O_1909,N_29625,N_29839);
and UO_1910 (O_1910,N_29556,N_29508);
or UO_1911 (O_1911,N_29649,N_29764);
or UO_1912 (O_1912,N_29542,N_29894);
and UO_1913 (O_1913,N_29595,N_29999);
nand UO_1914 (O_1914,N_29875,N_29606);
nor UO_1915 (O_1915,N_29473,N_29511);
and UO_1916 (O_1916,N_29581,N_29810);
nor UO_1917 (O_1917,N_29486,N_29966);
nand UO_1918 (O_1918,N_29792,N_29596);
nor UO_1919 (O_1919,N_29731,N_29907);
and UO_1920 (O_1920,N_29537,N_29885);
nand UO_1921 (O_1921,N_29468,N_29786);
xor UO_1922 (O_1922,N_29996,N_29588);
and UO_1923 (O_1923,N_29668,N_29599);
xnor UO_1924 (O_1924,N_29577,N_29972);
nor UO_1925 (O_1925,N_29824,N_29780);
and UO_1926 (O_1926,N_29903,N_29576);
or UO_1927 (O_1927,N_29443,N_29926);
or UO_1928 (O_1928,N_29880,N_29463);
xor UO_1929 (O_1929,N_29661,N_29833);
or UO_1930 (O_1930,N_29929,N_29846);
nand UO_1931 (O_1931,N_29996,N_29593);
xor UO_1932 (O_1932,N_29711,N_29874);
nand UO_1933 (O_1933,N_29990,N_29521);
nor UO_1934 (O_1934,N_29488,N_29621);
nor UO_1935 (O_1935,N_29692,N_29648);
and UO_1936 (O_1936,N_29804,N_29916);
and UO_1937 (O_1937,N_29784,N_29638);
or UO_1938 (O_1938,N_29641,N_29487);
and UO_1939 (O_1939,N_29893,N_29735);
or UO_1940 (O_1940,N_29557,N_29467);
and UO_1941 (O_1941,N_29648,N_29911);
nor UO_1942 (O_1942,N_29687,N_29554);
or UO_1943 (O_1943,N_29433,N_29480);
or UO_1944 (O_1944,N_29976,N_29790);
xnor UO_1945 (O_1945,N_29912,N_29680);
nor UO_1946 (O_1946,N_29760,N_29830);
nor UO_1947 (O_1947,N_29495,N_29995);
and UO_1948 (O_1948,N_29684,N_29954);
or UO_1949 (O_1949,N_29816,N_29540);
xnor UO_1950 (O_1950,N_29735,N_29859);
or UO_1951 (O_1951,N_29886,N_29829);
and UO_1952 (O_1952,N_29892,N_29651);
nor UO_1953 (O_1953,N_29716,N_29811);
nand UO_1954 (O_1954,N_29623,N_29991);
xor UO_1955 (O_1955,N_29508,N_29977);
nand UO_1956 (O_1956,N_29547,N_29517);
xnor UO_1957 (O_1957,N_29787,N_29493);
and UO_1958 (O_1958,N_29675,N_29993);
nor UO_1959 (O_1959,N_29459,N_29573);
and UO_1960 (O_1960,N_29932,N_29544);
nor UO_1961 (O_1961,N_29875,N_29557);
and UO_1962 (O_1962,N_29836,N_29922);
nand UO_1963 (O_1963,N_29430,N_29748);
nand UO_1964 (O_1964,N_29505,N_29426);
or UO_1965 (O_1965,N_29820,N_29680);
nand UO_1966 (O_1966,N_29425,N_29741);
nand UO_1967 (O_1967,N_29761,N_29676);
nor UO_1968 (O_1968,N_29765,N_29728);
nor UO_1969 (O_1969,N_29520,N_29477);
nand UO_1970 (O_1970,N_29448,N_29479);
nand UO_1971 (O_1971,N_29453,N_29751);
nand UO_1972 (O_1972,N_29449,N_29586);
xnor UO_1973 (O_1973,N_29517,N_29572);
nand UO_1974 (O_1974,N_29752,N_29618);
xnor UO_1975 (O_1975,N_29669,N_29659);
nand UO_1976 (O_1976,N_29770,N_29528);
or UO_1977 (O_1977,N_29801,N_29567);
or UO_1978 (O_1978,N_29481,N_29905);
and UO_1979 (O_1979,N_29422,N_29571);
nor UO_1980 (O_1980,N_29778,N_29718);
nor UO_1981 (O_1981,N_29988,N_29452);
or UO_1982 (O_1982,N_29548,N_29578);
nor UO_1983 (O_1983,N_29734,N_29908);
nand UO_1984 (O_1984,N_29476,N_29726);
and UO_1985 (O_1985,N_29848,N_29477);
and UO_1986 (O_1986,N_29713,N_29607);
or UO_1987 (O_1987,N_29680,N_29536);
or UO_1988 (O_1988,N_29662,N_29468);
nand UO_1989 (O_1989,N_29678,N_29422);
and UO_1990 (O_1990,N_29787,N_29726);
xnor UO_1991 (O_1991,N_29512,N_29676);
and UO_1992 (O_1992,N_29683,N_29637);
nor UO_1993 (O_1993,N_29698,N_29494);
nand UO_1994 (O_1994,N_29771,N_29598);
nor UO_1995 (O_1995,N_29492,N_29500);
xor UO_1996 (O_1996,N_29557,N_29698);
nor UO_1997 (O_1997,N_29953,N_29463);
nor UO_1998 (O_1998,N_29455,N_29579);
or UO_1999 (O_1999,N_29737,N_29806);
and UO_2000 (O_2000,N_29930,N_29404);
and UO_2001 (O_2001,N_29625,N_29410);
and UO_2002 (O_2002,N_29652,N_29649);
and UO_2003 (O_2003,N_29649,N_29473);
nand UO_2004 (O_2004,N_29466,N_29969);
and UO_2005 (O_2005,N_29703,N_29978);
nor UO_2006 (O_2006,N_29828,N_29908);
xnor UO_2007 (O_2007,N_29909,N_29935);
xnor UO_2008 (O_2008,N_29640,N_29884);
xnor UO_2009 (O_2009,N_29732,N_29674);
nor UO_2010 (O_2010,N_29867,N_29761);
nand UO_2011 (O_2011,N_29754,N_29963);
and UO_2012 (O_2012,N_29627,N_29634);
nand UO_2013 (O_2013,N_29445,N_29872);
or UO_2014 (O_2014,N_29837,N_29576);
xor UO_2015 (O_2015,N_29471,N_29621);
nor UO_2016 (O_2016,N_29494,N_29664);
nor UO_2017 (O_2017,N_29621,N_29468);
and UO_2018 (O_2018,N_29701,N_29630);
xnor UO_2019 (O_2019,N_29879,N_29999);
and UO_2020 (O_2020,N_29608,N_29938);
or UO_2021 (O_2021,N_29867,N_29985);
xor UO_2022 (O_2022,N_29682,N_29465);
and UO_2023 (O_2023,N_29701,N_29705);
or UO_2024 (O_2024,N_29895,N_29886);
and UO_2025 (O_2025,N_29810,N_29493);
or UO_2026 (O_2026,N_29424,N_29705);
xor UO_2027 (O_2027,N_29719,N_29858);
and UO_2028 (O_2028,N_29837,N_29707);
nor UO_2029 (O_2029,N_29621,N_29645);
or UO_2030 (O_2030,N_29671,N_29440);
nand UO_2031 (O_2031,N_29982,N_29646);
and UO_2032 (O_2032,N_29455,N_29838);
nor UO_2033 (O_2033,N_29543,N_29903);
nor UO_2034 (O_2034,N_29560,N_29403);
or UO_2035 (O_2035,N_29551,N_29523);
nor UO_2036 (O_2036,N_29690,N_29474);
xor UO_2037 (O_2037,N_29514,N_29776);
and UO_2038 (O_2038,N_29465,N_29539);
xnor UO_2039 (O_2039,N_29432,N_29707);
nor UO_2040 (O_2040,N_29955,N_29781);
nor UO_2041 (O_2041,N_29730,N_29661);
xnor UO_2042 (O_2042,N_29534,N_29655);
nor UO_2043 (O_2043,N_29890,N_29663);
nand UO_2044 (O_2044,N_29766,N_29865);
xor UO_2045 (O_2045,N_29429,N_29546);
nor UO_2046 (O_2046,N_29886,N_29431);
nand UO_2047 (O_2047,N_29754,N_29907);
nor UO_2048 (O_2048,N_29589,N_29994);
xor UO_2049 (O_2049,N_29828,N_29550);
or UO_2050 (O_2050,N_29474,N_29852);
nand UO_2051 (O_2051,N_29665,N_29570);
or UO_2052 (O_2052,N_29411,N_29578);
nand UO_2053 (O_2053,N_29502,N_29729);
or UO_2054 (O_2054,N_29993,N_29571);
or UO_2055 (O_2055,N_29407,N_29602);
and UO_2056 (O_2056,N_29716,N_29681);
and UO_2057 (O_2057,N_29608,N_29843);
xor UO_2058 (O_2058,N_29824,N_29700);
nand UO_2059 (O_2059,N_29528,N_29535);
nand UO_2060 (O_2060,N_29726,N_29659);
or UO_2061 (O_2061,N_29761,N_29844);
nor UO_2062 (O_2062,N_29975,N_29465);
nand UO_2063 (O_2063,N_29768,N_29552);
or UO_2064 (O_2064,N_29704,N_29788);
nor UO_2065 (O_2065,N_29479,N_29651);
nand UO_2066 (O_2066,N_29542,N_29904);
and UO_2067 (O_2067,N_29434,N_29473);
or UO_2068 (O_2068,N_29419,N_29968);
nand UO_2069 (O_2069,N_29856,N_29448);
nand UO_2070 (O_2070,N_29752,N_29418);
nand UO_2071 (O_2071,N_29581,N_29456);
nand UO_2072 (O_2072,N_29841,N_29610);
and UO_2073 (O_2073,N_29746,N_29729);
and UO_2074 (O_2074,N_29594,N_29895);
nand UO_2075 (O_2075,N_29459,N_29805);
nand UO_2076 (O_2076,N_29604,N_29520);
nor UO_2077 (O_2077,N_29641,N_29966);
nor UO_2078 (O_2078,N_29832,N_29624);
or UO_2079 (O_2079,N_29940,N_29559);
nor UO_2080 (O_2080,N_29948,N_29674);
nand UO_2081 (O_2081,N_29534,N_29675);
xor UO_2082 (O_2082,N_29478,N_29905);
and UO_2083 (O_2083,N_29466,N_29766);
and UO_2084 (O_2084,N_29863,N_29403);
nand UO_2085 (O_2085,N_29631,N_29468);
or UO_2086 (O_2086,N_29838,N_29628);
or UO_2087 (O_2087,N_29797,N_29987);
xnor UO_2088 (O_2088,N_29963,N_29463);
and UO_2089 (O_2089,N_29725,N_29514);
xor UO_2090 (O_2090,N_29457,N_29791);
nor UO_2091 (O_2091,N_29764,N_29665);
or UO_2092 (O_2092,N_29865,N_29658);
xor UO_2093 (O_2093,N_29451,N_29655);
nand UO_2094 (O_2094,N_29407,N_29657);
or UO_2095 (O_2095,N_29618,N_29469);
and UO_2096 (O_2096,N_29631,N_29932);
nor UO_2097 (O_2097,N_29572,N_29529);
xnor UO_2098 (O_2098,N_29804,N_29958);
and UO_2099 (O_2099,N_29401,N_29976);
nor UO_2100 (O_2100,N_29896,N_29750);
and UO_2101 (O_2101,N_29537,N_29936);
or UO_2102 (O_2102,N_29972,N_29803);
or UO_2103 (O_2103,N_29859,N_29594);
nand UO_2104 (O_2104,N_29837,N_29509);
and UO_2105 (O_2105,N_29403,N_29801);
xor UO_2106 (O_2106,N_29427,N_29954);
or UO_2107 (O_2107,N_29553,N_29960);
nor UO_2108 (O_2108,N_29803,N_29516);
or UO_2109 (O_2109,N_29429,N_29450);
nand UO_2110 (O_2110,N_29591,N_29548);
and UO_2111 (O_2111,N_29943,N_29646);
or UO_2112 (O_2112,N_29585,N_29918);
xnor UO_2113 (O_2113,N_29999,N_29881);
nand UO_2114 (O_2114,N_29496,N_29853);
nor UO_2115 (O_2115,N_29449,N_29992);
xor UO_2116 (O_2116,N_29442,N_29469);
or UO_2117 (O_2117,N_29406,N_29800);
xnor UO_2118 (O_2118,N_29402,N_29553);
xnor UO_2119 (O_2119,N_29487,N_29891);
xor UO_2120 (O_2120,N_29963,N_29432);
xnor UO_2121 (O_2121,N_29840,N_29489);
or UO_2122 (O_2122,N_29639,N_29441);
or UO_2123 (O_2123,N_29843,N_29779);
and UO_2124 (O_2124,N_29662,N_29881);
nor UO_2125 (O_2125,N_29993,N_29657);
or UO_2126 (O_2126,N_29733,N_29525);
or UO_2127 (O_2127,N_29474,N_29687);
xnor UO_2128 (O_2128,N_29841,N_29916);
xor UO_2129 (O_2129,N_29449,N_29745);
xor UO_2130 (O_2130,N_29725,N_29630);
nand UO_2131 (O_2131,N_29619,N_29681);
and UO_2132 (O_2132,N_29670,N_29829);
xnor UO_2133 (O_2133,N_29511,N_29740);
and UO_2134 (O_2134,N_29488,N_29520);
nand UO_2135 (O_2135,N_29410,N_29663);
or UO_2136 (O_2136,N_29955,N_29485);
nor UO_2137 (O_2137,N_29840,N_29514);
nand UO_2138 (O_2138,N_29764,N_29406);
and UO_2139 (O_2139,N_29807,N_29866);
nor UO_2140 (O_2140,N_29577,N_29955);
or UO_2141 (O_2141,N_29897,N_29636);
xnor UO_2142 (O_2142,N_29680,N_29755);
or UO_2143 (O_2143,N_29792,N_29870);
or UO_2144 (O_2144,N_29999,N_29744);
nand UO_2145 (O_2145,N_29893,N_29743);
and UO_2146 (O_2146,N_29616,N_29545);
nand UO_2147 (O_2147,N_29659,N_29580);
nor UO_2148 (O_2148,N_29586,N_29401);
and UO_2149 (O_2149,N_29970,N_29510);
nor UO_2150 (O_2150,N_29993,N_29793);
nor UO_2151 (O_2151,N_29602,N_29473);
nor UO_2152 (O_2152,N_29579,N_29559);
xor UO_2153 (O_2153,N_29503,N_29717);
nor UO_2154 (O_2154,N_29548,N_29682);
and UO_2155 (O_2155,N_29661,N_29825);
xnor UO_2156 (O_2156,N_29626,N_29813);
xor UO_2157 (O_2157,N_29493,N_29487);
nand UO_2158 (O_2158,N_29764,N_29729);
nor UO_2159 (O_2159,N_29995,N_29569);
nand UO_2160 (O_2160,N_29460,N_29736);
xnor UO_2161 (O_2161,N_29854,N_29987);
or UO_2162 (O_2162,N_29831,N_29634);
xnor UO_2163 (O_2163,N_29403,N_29624);
and UO_2164 (O_2164,N_29778,N_29595);
xor UO_2165 (O_2165,N_29453,N_29936);
nor UO_2166 (O_2166,N_29435,N_29990);
xor UO_2167 (O_2167,N_29892,N_29450);
nand UO_2168 (O_2168,N_29692,N_29733);
and UO_2169 (O_2169,N_29788,N_29528);
xnor UO_2170 (O_2170,N_29571,N_29717);
nor UO_2171 (O_2171,N_29616,N_29615);
nor UO_2172 (O_2172,N_29549,N_29849);
and UO_2173 (O_2173,N_29986,N_29838);
and UO_2174 (O_2174,N_29460,N_29911);
nor UO_2175 (O_2175,N_29550,N_29613);
xor UO_2176 (O_2176,N_29515,N_29935);
or UO_2177 (O_2177,N_29667,N_29549);
and UO_2178 (O_2178,N_29480,N_29758);
or UO_2179 (O_2179,N_29435,N_29936);
and UO_2180 (O_2180,N_29784,N_29418);
or UO_2181 (O_2181,N_29437,N_29966);
nand UO_2182 (O_2182,N_29437,N_29556);
or UO_2183 (O_2183,N_29427,N_29530);
nand UO_2184 (O_2184,N_29550,N_29594);
nand UO_2185 (O_2185,N_29629,N_29903);
nor UO_2186 (O_2186,N_29715,N_29524);
nor UO_2187 (O_2187,N_29939,N_29902);
nand UO_2188 (O_2188,N_29665,N_29595);
or UO_2189 (O_2189,N_29849,N_29953);
xnor UO_2190 (O_2190,N_29957,N_29978);
nor UO_2191 (O_2191,N_29686,N_29532);
and UO_2192 (O_2192,N_29986,N_29424);
nor UO_2193 (O_2193,N_29428,N_29485);
and UO_2194 (O_2194,N_29632,N_29474);
and UO_2195 (O_2195,N_29812,N_29831);
xnor UO_2196 (O_2196,N_29675,N_29804);
or UO_2197 (O_2197,N_29617,N_29432);
xor UO_2198 (O_2198,N_29988,N_29880);
xnor UO_2199 (O_2199,N_29881,N_29816);
nor UO_2200 (O_2200,N_29821,N_29676);
and UO_2201 (O_2201,N_29930,N_29710);
or UO_2202 (O_2202,N_29720,N_29745);
xnor UO_2203 (O_2203,N_29495,N_29400);
and UO_2204 (O_2204,N_29964,N_29888);
xnor UO_2205 (O_2205,N_29824,N_29935);
xnor UO_2206 (O_2206,N_29957,N_29634);
or UO_2207 (O_2207,N_29607,N_29752);
nor UO_2208 (O_2208,N_29706,N_29958);
nor UO_2209 (O_2209,N_29586,N_29745);
nand UO_2210 (O_2210,N_29993,N_29911);
nand UO_2211 (O_2211,N_29960,N_29703);
and UO_2212 (O_2212,N_29668,N_29583);
nor UO_2213 (O_2213,N_29839,N_29518);
xor UO_2214 (O_2214,N_29942,N_29706);
or UO_2215 (O_2215,N_29711,N_29617);
and UO_2216 (O_2216,N_29664,N_29846);
and UO_2217 (O_2217,N_29804,N_29976);
xor UO_2218 (O_2218,N_29560,N_29768);
and UO_2219 (O_2219,N_29580,N_29813);
and UO_2220 (O_2220,N_29795,N_29617);
nor UO_2221 (O_2221,N_29674,N_29749);
or UO_2222 (O_2222,N_29478,N_29657);
xor UO_2223 (O_2223,N_29907,N_29870);
or UO_2224 (O_2224,N_29936,N_29853);
xor UO_2225 (O_2225,N_29794,N_29585);
xor UO_2226 (O_2226,N_29792,N_29425);
xor UO_2227 (O_2227,N_29952,N_29551);
nor UO_2228 (O_2228,N_29534,N_29463);
or UO_2229 (O_2229,N_29451,N_29693);
nor UO_2230 (O_2230,N_29901,N_29427);
nor UO_2231 (O_2231,N_29931,N_29819);
nand UO_2232 (O_2232,N_29877,N_29988);
or UO_2233 (O_2233,N_29661,N_29734);
xor UO_2234 (O_2234,N_29732,N_29546);
or UO_2235 (O_2235,N_29706,N_29861);
nor UO_2236 (O_2236,N_29895,N_29447);
xnor UO_2237 (O_2237,N_29473,N_29984);
and UO_2238 (O_2238,N_29578,N_29607);
or UO_2239 (O_2239,N_29990,N_29654);
or UO_2240 (O_2240,N_29500,N_29648);
xnor UO_2241 (O_2241,N_29947,N_29617);
nand UO_2242 (O_2242,N_29462,N_29686);
nor UO_2243 (O_2243,N_29859,N_29416);
nand UO_2244 (O_2244,N_29700,N_29855);
and UO_2245 (O_2245,N_29834,N_29602);
nor UO_2246 (O_2246,N_29889,N_29841);
or UO_2247 (O_2247,N_29962,N_29616);
xnor UO_2248 (O_2248,N_29472,N_29634);
nor UO_2249 (O_2249,N_29949,N_29907);
xnor UO_2250 (O_2250,N_29977,N_29627);
xor UO_2251 (O_2251,N_29693,N_29948);
nor UO_2252 (O_2252,N_29477,N_29864);
or UO_2253 (O_2253,N_29755,N_29817);
or UO_2254 (O_2254,N_29430,N_29921);
or UO_2255 (O_2255,N_29746,N_29713);
nand UO_2256 (O_2256,N_29598,N_29538);
and UO_2257 (O_2257,N_29498,N_29739);
nor UO_2258 (O_2258,N_29874,N_29484);
xor UO_2259 (O_2259,N_29565,N_29478);
nor UO_2260 (O_2260,N_29834,N_29996);
and UO_2261 (O_2261,N_29423,N_29873);
or UO_2262 (O_2262,N_29411,N_29478);
or UO_2263 (O_2263,N_29867,N_29642);
nand UO_2264 (O_2264,N_29447,N_29724);
xor UO_2265 (O_2265,N_29414,N_29874);
nand UO_2266 (O_2266,N_29468,N_29544);
xnor UO_2267 (O_2267,N_29691,N_29463);
nand UO_2268 (O_2268,N_29562,N_29624);
or UO_2269 (O_2269,N_29512,N_29821);
nand UO_2270 (O_2270,N_29597,N_29996);
nand UO_2271 (O_2271,N_29787,N_29892);
xor UO_2272 (O_2272,N_29526,N_29967);
nor UO_2273 (O_2273,N_29558,N_29805);
or UO_2274 (O_2274,N_29765,N_29619);
nor UO_2275 (O_2275,N_29687,N_29948);
and UO_2276 (O_2276,N_29604,N_29576);
nand UO_2277 (O_2277,N_29461,N_29851);
nor UO_2278 (O_2278,N_29562,N_29568);
or UO_2279 (O_2279,N_29823,N_29724);
or UO_2280 (O_2280,N_29966,N_29841);
nor UO_2281 (O_2281,N_29557,N_29667);
or UO_2282 (O_2282,N_29885,N_29874);
xor UO_2283 (O_2283,N_29773,N_29913);
and UO_2284 (O_2284,N_29774,N_29752);
and UO_2285 (O_2285,N_29635,N_29470);
or UO_2286 (O_2286,N_29550,N_29448);
or UO_2287 (O_2287,N_29924,N_29937);
nand UO_2288 (O_2288,N_29460,N_29531);
nor UO_2289 (O_2289,N_29543,N_29824);
nor UO_2290 (O_2290,N_29855,N_29799);
nand UO_2291 (O_2291,N_29663,N_29965);
nand UO_2292 (O_2292,N_29731,N_29955);
or UO_2293 (O_2293,N_29585,N_29680);
or UO_2294 (O_2294,N_29807,N_29568);
nand UO_2295 (O_2295,N_29976,N_29717);
nand UO_2296 (O_2296,N_29653,N_29532);
xor UO_2297 (O_2297,N_29631,N_29528);
or UO_2298 (O_2298,N_29823,N_29756);
and UO_2299 (O_2299,N_29979,N_29740);
xor UO_2300 (O_2300,N_29569,N_29532);
nor UO_2301 (O_2301,N_29576,N_29630);
nand UO_2302 (O_2302,N_29609,N_29883);
xnor UO_2303 (O_2303,N_29806,N_29499);
and UO_2304 (O_2304,N_29598,N_29840);
and UO_2305 (O_2305,N_29747,N_29929);
nand UO_2306 (O_2306,N_29488,N_29884);
or UO_2307 (O_2307,N_29525,N_29487);
nor UO_2308 (O_2308,N_29749,N_29938);
nand UO_2309 (O_2309,N_29698,N_29718);
nand UO_2310 (O_2310,N_29780,N_29602);
and UO_2311 (O_2311,N_29846,N_29488);
or UO_2312 (O_2312,N_29433,N_29755);
and UO_2313 (O_2313,N_29810,N_29490);
and UO_2314 (O_2314,N_29866,N_29426);
and UO_2315 (O_2315,N_29457,N_29678);
or UO_2316 (O_2316,N_29433,N_29976);
xor UO_2317 (O_2317,N_29919,N_29805);
nand UO_2318 (O_2318,N_29793,N_29948);
xnor UO_2319 (O_2319,N_29762,N_29433);
nand UO_2320 (O_2320,N_29739,N_29614);
or UO_2321 (O_2321,N_29508,N_29723);
nor UO_2322 (O_2322,N_29860,N_29464);
nor UO_2323 (O_2323,N_29979,N_29807);
or UO_2324 (O_2324,N_29922,N_29999);
nor UO_2325 (O_2325,N_29982,N_29501);
or UO_2326 (O_2326,N_29449,N_29709);
xnor UO_2327 (O_2327,N_29551,N_29972);
and UO_2328 (O_2328,N_29707,N_29841);
xor UO_2329 (O_2329,N_29441,N_29891);
and UO_2330 (O_2330,N_29459,N_29973);
nand UO_2331 (O_2331,N_29599,N_29591);
xor UO_2332 (O_2332,N_29729,N_29791);
or UO_2333 (O_2333,N_29712,N_29930);
or UO_2334 (O_2334,N_29914,N_29532);
nand UO_2335 (O_2335,N_29578,N_29443);
or UO_2336 (O_2336,N_29741,N_29655);
nand UO_2337 (O_2337,N_29467,N_29668);
xor UO_2338 (O_2338,N_29589,N_29918);
xor UO_2339 (O_2339,N_29869,N_29980);
or UO_2340 (O_2340,N_29818,N_29602);
or UO_2341 (O_2341,N_29691,N_29688);
and UO_2342 (O_2342,N_29752,N_29860);
xnor UO_2343 (O_2343,N_29927,N_29543);
nand UO_2344 (O_2344,N_29716,N_29684);
xor UO_2345 (O_2345,N_29569,N_29667);
and UO_2346 (O_2346,N_29812,N_29878);
nand UO_2347 (O_2347,N_29448,N_29660);
nand UO_2348 (O_2348,N_29703,N_29583);
xor UO_2349 (O_2349,N_29931,N_29559);
and UO_2350 (O_2350,N_29684,N_29983);
and UO_2351 (O_2351,N_29978,N_29986);
nor UO_2352 (O_2352,N_29867,N_29789);
and UO_2353 (O_2353,N_29856,N_29510);
xor UO_2354 (O_2354,N_29573,N_29862);
or UO_2355 (O_2355,N_29823,N_29584);
xnor UO_2356 (O_2356,N_29943,N_29830);
and UO_2357 (O_2357,N_29785,N_29731);
and UO_2358 (O_2358,N_29520,N_29683);
and UO_2359 (O_2359,N_29926,N_29416);
and UO_2360 (O_2360,N_29904,N_29452);
or UO_2361 (O_2361,N_29573,N_29804);
and UO_2362 (O_2362,N_29958,N_29692);
nor UO_2363 (O_2363,N_29526,N_29872);
nand UO_2364 (O_2364,N_29905,N_29970);
and UO_2365 (O_2365,N_29418,N_29912);
nor UO_2366 (O_2366,N_29496,N_29984);
or UO_2367 (O_2367,N_29822,N_29969);
or UO_2368 (O_2368,N_29495,N_29588);
and UO_2369 (O_2369,N_29654,N_29431);
and UO_2370 (O_2370,N_29694,N_29996);
nor UO_2371 (O_2371,N_29705,N_29496);
nand UO_2372 (O_2372,N_29798,N_29627);
xor UO_2373 (O_2373,N_29731,N_29853);
xor UO_2374 (O_2374,N_29422,N_29771);
nor UO_2375 (O_2375,N_29893,N_29500);
and UO_2376 (O_2376,N_29745,N_29445);
and UO_2377 (O_2377,N_29443,N_29689);
xor UO_2378 (O_2378,N_29954,N_29829);
and UO_2379 (O_2379,N_29950,N_29526);
or UO_2380 (O_2380,N_29969,N_29490);
xor UO_2381 (O_2381,N_29881,N_29886);
or UO_2382 (O_2382,N_29600,N_29785);
and UO_2383 (O_2383,N_29996,N_29799);
or UO_2384 (O_2384,N_29662,N_29810);
nor UO_2385 (O_2385,N_29734,N_29563);
nor UO_2386 (O_2386,N_29859,N_29617);
xnor UO_2387 (O_2387,N_29440,N_29451);
or UO_2388 (O_2388,N_29639,N_29931);
nand UO_2389 (O_2389,N_29502,N_29755);
nand UO_2390 (O_2390,N_29712,N_29474);
or UO_2391 (O_2391,N_29783,N_29548);
nand UO_2392 (O_2392,N_29668,N_29999);
xnor UO_2393 (O_2393,N_29964,N_29673);
nor UO_2394 (O_2394,N_29528,N_29404);
and UO_2395 (O_2395,N_29658,N_29969);
xor UO_2396 (O_2396,N_29873,N_29988);
and UO_2397 (O_2397,N_29687,N_29628);
xor UO_2398 (O_2398,N_29556,N_29406);
and UO_2399 (O_2399,N_29946,N_29554);
nor UO_2400 (O_2400,N_29832,N_29859);
nor UO_2401 (O_2401,N_29641,N_29644);
or UO_2402 (O_2402,N_29638,N_29957);
nor UO_2403 (O_2403,N_29603,N_29498);
nand UO_2404 (O_2404,N_29507,N_29923);
and UO_2405 (O_2405,N_29665,N_29897);
or UO_2406 (O_2406,N_29423,N_29937);
nand UO_2407 (O_2407,N_29877,N_29550);
or UO_2408 (O_2408,N_29812,N_29997);
or UO_2409 (O_2409,N_29988,N_29994);
nor UO_2410 (O_2410,N_29874,N_29780);
nand UO_2411 (O_2411,N_29928,N_29853);
or UO_2412 (O_2412,N_29946,N_29896);
xor UO_2413 (O_2413,N_29785,N_29975);
or UO_2414 (O_2414,N_29462,N_29502);
nand UO_2415 (O_2415,N_29748,N_29624);
nand UO_2416 (O_2416,N_29922,N_29579);
and UO_2417 (O_2417,N_29452,N_29559);
and UO_2418 (O_2418,N_29405,N_29859);
or UO_2419 (O_2419,N_29538,N_29462);
xnor UO_2420 (O_2420,N_29922,N_29964);
or UO_2421 (O_2421,N_29986,N_29453);
or UO_2422 (O_2422,N_29920,N_29665);
nor UO_2423 (O_2423,N_29666,N_29876);
nand UO_2424 (O_2424,N_29605,N_29591);
and UO_2425 (O_2425,N_29451,N_29599);
nor UO_2426 (O_2426,N_29592,N_29529);
xnor UO_2427 (O_2427,N_29585,N_29592);
xnor UO_2428 (O_2428,N_29426,N_29614);
or UO_2429 (O_2429,N_29768,N_29439);
nand UO_2430 (O_2430,N_29909,N_29861);
nor UO_2431 (O_2431,N_29559,N_29440);
nand UO_2432 (O_2432,N_29586,N_29647);
xor UO_2433 (O_2433,N_29910,N_29629);
xor UO_2434 (O_2434,N_29579,N_29575);
xor UO_2435 (O_2435,N_29475,N_29931);
and UO_2436 (O_2436,N_29574,N_29869);
xnor UO_2437 (O_2437,N_29965,N_29622);
xor UO_2438 (O_2438,N_29753,N_29959);
and UO_2439 (O_2439,N_29761,N_29679);
and UO_2440 (O_2440,N_29864,N_29890);
xor UO_2441 (O_2441,N_29684,N_29824);
nor UO_2442 (O_2442,N_29823,N_29588);
xor UO_2443 (O_2443,N_29937,N_29631);
nand UO_2444 (O_2444,N_29706,N_29962);
nor UO_2445 (O_2445,N_29679,N_29671);
nor UO_2446 (O_2446,N_29858,N_29555);
or UO_2447 (O_2447,N_29842,N_29570);
xnor UO_2448 (O_2448,N_29751,N_29686);
nand UO_2449 (O_2449,N_29706,N_29731);
and UO_2450 (O_2450,N_29484,N_29905);
nand UO_2451 (O_2451,N_29975,N_29461);
nand UO_2452 (O_2452,N_29618,N_29746);
and UO_2453 (O_2453,N_29786,N_29442);
nor UO_2454 (O_2454,N_29832,N_29737);
nand UO_2455 (O_2455,N_29686,N_29926);
nor UO_2456 (O_2456,N_29439,N_29461);
nand UO_2457 (O_2457,N_29473,N_29489);
nor UO_2458 (O_2458,N_29610,N_29742);
or UO_2459 (O_2459,N_29860,N_29872);
xor UO_2460 (O_2460,N_29631,N_29737);
nor UO_2461 (O_2461,N_29444,N_29980);
or UO_2462 (O_2462,N_29719,N_29954);
xnor UO_2463 (O_2463,N_29407,N_29477);
and UO_2464 (O_2464,N_29804,N_29543);
xnor UO_2465 (O_2465,N_29527,N_29659);
or UO_2466 (O_2466,N_29934,N_29691);
or UO_2467 (O_2467,N_29737,N_29712);
nor UO_2468 (O_2468,N_29983,N_29561);
and UO_2469 (O_2469,N_29426,N_29674);
xnor UO_2470 (O_2470,N_29400,N_29805);
and UO_2471 (O_2471,N_29604,N_29476);
nand UO_2472 (O_2472,N_29516,N_29878);
nor UO_2473 (O_2473,N_29772,N_29852);
and UO_2474 (O_2474,N_29706,N_29825);
and UO_2475 (O_2475,N_29950,N_29833);
nand UO_2476 (O_2476,N_29509,N_29510);
nor UO_2477 (O_2477,N_29685,N_29710);
and UO_2478 (O_2478,N_29733,N_29670);
or UO_2479 (O_2479,N_29953,N_29449);
or UO_2480 (O_2480,N_29885,N_29998);
xor UO_2481 (O_2481,N_29617,N_29897);
nor UO_2482 (O_2482,N_29683,N_29616);
and UO_2483 (O_2483,N_29476,N_29962);
xor UO_2484 (O_2484,N_29538,N_29767);
and UO_2485 (O_2485,N_29444,N_29669);
xor UO_2486 (O_2486,N_29564,N_29454);
or UO_2487 (O_2487,N_29845,N_29750);
nand UO_2488 (O_2488,N_29548,N_29733);
nand UO_2489 (O_2489,N_29416,N_29794);
and UO_2490 (O_2490,N_29716,N_29870);
or UO_2491 (O_2491,N_29680,N_29989);
and UO_2492 (O_2492,N_29961,N_29420);
or UO_2493 (O_2493,N_29871,N_29446);
nand UO_2494 (O_2494,N_29512,N_29771);
xor UO_2495 (O_2495,N_29936,N_29811);
nor UO_2496 (O_2496,N_29443,N_29965);
and UO_2497 (O_2497,N_29632,N_29694);
and UO_2498 (O_2498,N_29458,N_29942);
and UO_2499 (O_2499,N_29459,N_29602);
and UO_2500 (O_2500,N_29494,N_29749);
nand UO_2501 (O_2501,N_29572,N_29459);
or UO_2502 (O_2502,N_29685,N_29553);
nor UO_2503 (O_2503,N_29992,N_29707);
and UO_2504 (O_2504,N_29668,N_29867);
nand UO_2505 (O_2505,N_29720,N_29823);
nor UO_2506 (O_2506,N_29703,N_29807);
nor UO_2507 (O_2507,N_29631,N_29551);
or UO_2508 (O_2508,N_29732,N_29553);
xor UO_2509 (O_2509,N_29606,N_29831);
or UO_2510 (O_2510,N_29590,N_29679);
nand UO_2511 (O_2511,N_29587,N_29473);
or UO_2512 (O_2512,N_29803,N_29832);
or UO_2513 (O_2513,N_29587,N_29582);
nand UO_2514 (O_2514,N_29775,N_29723);
nand UO_2515 (O_2515,N_29413,N_29570);
nor UO_2516 (O_2516,N_29591,N_29772);
nor UO_2517 (O_2517,N_29691,N_29981);
nor UO_2518 (O_2518,N_29711,N_29792);
nand UO_2519 (O_2519,N_29824,N_29666);
and UO_2520 (O_2520,N_29783,N_29792);
nor UO_2521 (O_2521,N_29769,N_29919);
and UO_2522 (O_2522,N_29703,N_29805);
nand UO_2523 (O_2523,N_29993,N_29709);
nand UO_2524 (O_2524,N_29534,N_29475);
and UO_2525 (O_2525,N_29787,N_29834);
nand UO_2526 (O_2526,N_29664,N_29787);
nand UO_2527 (O_2527,N_29915,N_29947);
nor UO_2528 (O_2528,N_29953,N_29659);
and UO_2529 (O_2529,N_29882,N_29631);
nand UO_2530 (O_2530,N_29435,N_29812);
and UO_2531 (O_2531,N_29870,N_29544);
or UO_2532 (O_2532,N_29635,N_29734);
and UO_2533 (O_2533,N_29885,N_29878);
nor UO_2534 (O_2534,N_29966,N_29565);
nand UO_2535 (O_2535,N_29426,N_29552);
nand UO_2536 (O_2536,N_29510,N_29908);
nor UO_2537 (O_2537,N_29868,N_29741);
or UO_2538 (O_2538,N_29985,N_29807);
or UO_2539 (O_2539,N_29710,N_29557);
or UO_2540 (O_2540,N_29523,N_29946);
xor UO_2541 (O_2541,N_29788,N_29616);
xor UO_2542 (O_2542,N_29456,N_29641);
xnor UO_2543 (O_2543,N_29606,N_29702);
nand UO_2544 (O_2544,N_29612,N_29646);
nor UO_2545 (O_2545,N_29861,N_29423);
and UO_2546 (O_2546,N_29933,N_29538);
or UO_2547 (O_2547,N_29809,N_29733);
xnor UO_2548 (O_2548,N_29487,N_29812);
xnor UO_2549 (O_2549,N_29698,N_29936);
nor UO_2550 (O_2550,N_29865,N_29494);
or UO_2551 (O_2551,N_29818,N_29788);
nor UO_2552 (O_2552,N_29457,N_29691);
nor UO_2553 (O_2553,N_29942,N_29527);
and UO_2554 (O_2554,N_29707,N_29965);
and UO_2555 (O_2555,N_29665,N_29630);
nand UO_2556 (O_2556,N_29829,N_29589);
and UO_2557 (O_2557,N_29980,N_29981);
nor UO_2558 (O_2558,N_29744,N_29827);
and UO_2559 (O_2559,N_29891,N_29616);
nor UO_2560 (O_2560,N_29765,N_29430);
or UO_2561 (O_2561,N_29610,N_29771);
and UO_2562 (O_2562,N_29657,N_29518);
xnor UO_2563 (O_2563,N_29413,N_29862);
nor UO_2564 (O_2564,N_29852,N_29975);
xnor UO_2565 (O_2565,N_29968,N_29823);
or UO_2566 (O_2566,N_29794,N_29815);
nor UO_2567 (O_2567,N_29825,N_29749);
and UO_2568 (O_2568,N_29921,N_29952);
xor UO_2569 (O_2569,N_29601,N_29428);
and UO_2570 (O_2570,N_29513,N_29843);
or UO_2571 (O_2571,N_29720,N_29936);
xnor UO_2572 (O_2572,N_29938,N_29457);
and UO_2573 (O_2573,N_29764,N_29832);
nor UO_2574 (O_2574,N_29595,N_29964);
and UO_2575 (O_2575,N_29760,N_29673);
nor UO_2576 (O_2576,N_29858,N_29661);
nor UO_2577 (O_2577,N_29699,N_29464);
and UO_2578 (O_2578,N_29620,N_29925);
or UO_2579 (O_2579,N_29427,N_29914);
and UO_2580 (O_2580,N_29469,N_29423);
nor UO_2581 (O_2581,N_29706,N_29828);
or UO_2582 (O_2582,N_29972,N_29903);
nand UO_2583 (O_2583,N_29413,N_29741);
and UO_2584 (O_2584,N_29836,N_29829);
nor UO_2585 (O_2585,N_29415,N_29566);
and UO_2586 (O_2586,N_29815,N_29860);
nand UO_2587 (O_2587,N_29508,N_29634);
and UO_2588 (O_2588,N_29980,N_29551);
nor UO_2589 (O_2589,N_29895,N_29834);
xor UO_2590 (O_2590,N_29434,N_29821);
nor UO_2591 (O_2591,N_29624,N_29742);
or UO_2592 (O_2592,N_29709,N_29937);
xnor UO_2593 (O_2593,N_29707,N_29625);
or UO_2594 (O_2594,N_29544,N_29961);
xnor UO_2595 (O_2595,N_29750,N_29570);
nor UO_2596 (O_2596,N_29681,N_29700);
or UO_2597 (O_2597,N_29988,N_29746);
nor UO_2598 (O_2598,N_29726,N_29882);
xnor UO_2599 (O_2599,N_29552,N_29758);
and UO_2600 (O_2600,N_29891,N_29625);
nand UO_2601 (O_2601,N_29505,N_29886);
xor UO_2602 (O_2602,N_29692,N_29418);
xor UO_2603 (O_2603,N_29844,N_29507);
and UO_2604 (O_2604,N_29803,N_29575);
xnor UO_2605 (O_2605,N_29646,N_29502);
nor UO_2606 (O_2606,N_29728,N_29593);
xor UO_2607 (O_2607,N_29844,N_29593);
nand UO_2608 (O_2608,N_29976,N_29470);
or UO_2609 (O_2609,N_29624,N_29905);
xor UO_2610 (O_2610,N_29848,N_29768);
nor UO_2611 (O_2611,N_29800,N_29980);
nand UO_2612 (O_2612,N_29856,N_29923);
nor UO_2613 (O_2613,N_29710,N_29844);
nand UO_2614 (O_2614,N_29622,N_29547);
or UO_2615 (O_2615,N_29552,N_29515);
and UO_2616 (O_2616,N_29823,N_29625);
or UO_2617 (O_2617,N_29754,N_29491);
or UO_2618 (O_2618,N_29889,N_29713);
nand UO_2619 (O_2619,N_29647,N_29673);
xor UO_2620 (O_2620,N_29764,N_29615);
nor UO_2621 (O_2621,N_29670,N_29930);
nor UO_2622 (O_2622,N_29603,N_29838);
nand UO_2623 (O_2623,N_29560,N_29452);
and UO_2624 (O_2624,N_29887,N_29991);
and UO_2625 (O_2625,N_29419,N_29890);
and UO_2626 (O_2626,N_29597,N_29808);
nor UO_2627 (O_2627,N_29767,N_29971);
nand UO_2628 (O_2628,N_29799,N_29835);
and UO_2629 (O_2629,N_29620,N_29523);
xnor UO_2630 (O_2630,N_29966,N_29791);
or UO_2631 (O_2631,N_29982,N_29887);
nor UO_2632 (O_2632,N_29853,N_29466);
or UO_2633 (O_2633,N_29879,N_29451);
nand UO_2634 (O_2634,N_29719,N_29501);
xnor UO_2635 (O_2635,N_29839,N_29687);
nand UO_2636 (O_2636,N_29444,N_29844);
nand UO_2637 (O_2637,N_29551,N_29944);
nor UO_2638 (O_2638,N_29852,N_29797);
or UO_2639 (O_2639,N_29431,N_29661);
nor UO_2640 (O_2640,N_29441,N_29973);
nor UO_2641 (O_2641,N_29761,N_29428);
nor UO_2642 (O_2642,N_29728,N_29827);
or UO_2643 (O_2643,N_29449,N_29929);
nor UO_2644 (O_2644,N_29741,N_29782);
nor UO_2645 (O_2645,N_29709,N_29561);
and UO_2646 (O_2646,N_29724,N_29622);
nor UO_2647 (O_2647,N_29976,N_29887);
xnor UO_2648 (O_2648,N_29831,N_29594);
or UO_2649 (O_2649,N_29720,N_29625);
nor UO_2650 (O_2650,N_29638,N_29467);
xnor UO_2651 (O_2651,N_29553,N_29565);
nand UO_2652 (O_2652,N_29687,N_29445);
nand UO_2653 (O_2653,N_29816,N_29520);
xor UO_2654 (O_2654,N_29500,N_29840);
or UO_2655 (O_2655,N_29987,N_29763);
or UO_2656 (O_2656,N_29841,N_29899);
nand UO_2657 (O_2657,N_29949,N_29728);
or UO_2658 (O_2658,N_29669,N_29997);
xor UO_2659 (O_2659,N_29766,N_29804);
or UO_2660 (O_2660,N_29487,N_29923);
nor UO_2661 (O_2661,N_29915,N_29571);
nor UO_2662 (O_2662,N_29842,N_29949);
and UO_2663 (O_2663,N_29495,N_29751);
nor UO_2664 (O_2664,N_29828,N_29705);
nor UO_2665 (O_2665,N_29706,N_29886);
xnor UO_2666 (O_2666,N_29405,N_29829);
or UO_2667 (O_2667,N_29492,N_29955);
and UO_2668 (O_2668,N_29875,N_29849);
and UO_2669 (O_2669,N_29659,N_29787);
or UO_2670 (O_2670,N_29899,N_29892);
nand UO_2671 (O_2671,N_29687,N_29414);
or UO_2672 (O_2672,N_29765,N_29674);
nand UO_2673 (O_2673,N_29707,N_29567);
or UO_2674 (O_2674,N_29441,N_29774);
xor UO_2675 (O_2675,N_29895,N_29732);
xnor UO_2676 (O_2676,N_29938,N_29716);
nor UO_2677 (O_2677,N_29861,N_29785);
xor UO_2678 (O_2678,N_29852,N_29656);
nor UO_2679 (O_2679,N_29410,N_29818);
or UO_2680 (O_2680,N_29637,N_29636);
nor UO_2681 (O_2681,N_29956,N_29804);
or UO_2682 (O_2682,N_29465,N_29435);
or UO_2683 (O_2683,N_29448,N_29691);
nor UO_2684 (O_2684,N_29866,N_29403);
and UO_2685 (O_2685,N_29445,N_29853);
nor UO_2686 (O_2686,N_29539,N_29442);
and UO_2687 (O_2687,N_29828,N_29834);
and UO_2688 (O_2688,N_29887,N_29831);
nand UO_2689 (O_2689,N_29952,N_29798);
nor UO_2690 (O_2690,N_29967,N_29519);
xor UO_2691 (O_2691,N_29655,N_29576);
nand UO_2692 (O_2692,N_29551,N_29726);
xor UO_2693 (O_2693,N_29504,N_29968);
xor UO_2694 (O_2694,N_29930,N_29637);
nand UO_2695 (O_2695,N_29633,N_29966);
xor UO_2696 (O_2696,N_29672,N_29400);
or UO_2697 (O_2697,N_29664,N_29980);
nand UO_2698 (O_2698,N_29684,N_29742);
nor UO_2699 (O_2699,N_29406,N_29593);
xnor UO_2700 (O_2700,N_29410,N_29513);
or UO_2701 (O_2701,N_29965,N_29640);
nor UO_2702 (O_2702,N_29623,N_29616);
or UO_2703 (O_2703,N_29476,N_29929);
and UO_2704 (O_2704,N_29624,N_29851);
nand UO_2705 (O_2705,N_29425,N_29677);
and UO_2706 (O_2706,N_29786,N_29821);
xor UO_2707 (O_2707,N_29999,N_29988);
nor UO_2708 (O_2708,N_29610,N_29476);
and UO_2709 (O_2709,N_29451,N_29562);
and UO_2710 (O_2710,N_29442,N_29707);
and UO_2711 (O_2711,N_29513,N_29827);
nand UO_2712 (O_2712,N_29903,N_29760);
and UO_2713 (O_2713,N_29683,N_29552);
or UO_2714 (O_2714,N_29979,N_29929);
nor UO_2715 (O_2715,N_29757,N_29563);
and UO_2716 (O_2716,N_29708,N_29730);
or UO_2717 (O_2717,N_29694,N_29454);
nand UO_2718 (O_2718,N_29542,N_29937);
xnor UO_2719 (O_2719,N_29656,N_29537);
and UO_2720 (O_2720,N_29499,N_29625);
xnor UO_2721 (O_2721,N_29677,N_29746);
and UO_2722 (O_2722,N_29954,N_29977);
xor UO_2723 (O_2723,N_29505,N_29568);
and UO_2724 (O_2724,N_29689,N_29888);
and UO_2725 (O_2725,N_29511,N_29411);
nand UO_2726 (O_2726,N_29728,N_29840);
or UO_2727 (O_2727,N_29696,N_29866);
or UO_2728 (O_2728,N_29723,N_29512);
or UO_2729 (O_2729,N_29488,N_29653);
nor UO_2730 (O_2730,N_29498,N_29843);
nor UO_2731 (O_2731,N_29476,N_29424);
or UO_2732 (O_2732,N_29445,N_29534);
and UO_2733 (O_2733,N_29654,N_29414);
nor UO_2734 (O_2734,N_29898,N_29678);
nor UO_2735 (O_2735,N_29862,N_29589);
xor UO_2736 (O_2736,N_29573,N_29952);
nand UO_2737 (O_2737,N_29952,N_29792);
nand UO_2738 (O_2738,N_29792,N_29728);
xnor UO_2739 (O_2739,N_29860,N_29511);
or UO_2740 (O_2740,N_29451,N_29439);
nor UO_2741 (O_2741,N_29943,N_29626);
xnor UO_2742 (O_2742,N_29753,N_29561);
and UO_2743 (O_2743,N_29674,N_29578);
or UO_2744 (O_2744,N_29745,N_29405);
nand UO_2745 (O_2745,N_29773,N_29933);
nand UO_2746 (O_2746,N_29697,N_29915);
and UO_2747 (O_2747,N_29932,N_29867);
xor UO_2748 (O_2748,N_29415,N_29498);
nor UO_2749 (O_2749,N_29417,N_29984);
xnor UO_2750 (O_2750,N_29472,N_29650);
xnor UO_2751 (O_2751,N_29577,N_29925);
nand UO_2752 (O_2752,N_29484,N_29465);
nand UO_2753 (O_2753,N_29673,N_29723);
and UO_2754 (O_2754,N_29723,N_29610);
xnor UO_2755 (O_2755,N_29973,N_29644);
and UO_2756 (O_2756,N_29904,N_29413);
or UO_2757 (O_2757,N_29767,N_29949);
nand UO_2758 (O_2758,N_29940,N_29698);
nand UO_2759 (O_2759,N_29935,N_29880);
and UO_2760 (O_2760,N_29573,N_29622);
and UO_2761 (O_2761,N_29712,N_29729);
nand UO_2762 (O_2762,N_29646,N_29678);
and UO_2763 (O_2763,N_29911,N_29895);
xnor UO_2764 (O_2764,N_29553,N_29980);
nand UO_2765 (O_2765,N_29948,N_29458);
nand UO_2766 (O_2766,N_29782,N_29483);
or UO_2767 (O_2767,N_29900,N_29939);
xor UO_2768 (O_2768,N_29455,N_29821);
nor UO_2769 (O_2769,N_29562,N_29874);
nand UO_2770 (O_2770,N_29945,N_29510);
and UO_2771 (O_2771,N_29631,N_29815);
xnor UO_2772 (O_2772,N_29906,N_29518);
nand UO_2773 (O_2773,N_29570,N_29576);
xor UO_2774 (O_2774,N_29768,N_29546);
nor UO_2775 (O_2775,N_29914,N_29888);
xnor UO_2776 (O_2776,N_29851,N_29434);
nand UO_2777 (O_2777,N_29581,N_29439);
and UO_2778 (O_2778,N_29490,N_29518);
or UO_2779 (O_2779,N_29966,N_29433);
xor UO_2780 (O_2780,N_29816,N_29548);
xor UO_2781 (O_2781,N_29977,N_29432);
xor UO_2782 (O_2782,N_29906,N_29946);
or UO_2783 (O_2783,N_29688,N_29969);
xnor UO_2784 (O_2784,N_29501,N_29566);
xor UO_2785 (O_2785,N_29495,N_29815);
and UO_2786 (O_2786,N_29719,N_29581);
xnor UO_2787 (O_2787,N_29686,N_29485);
nand UO_2788 (O_2788,N_29953,N_29626);
nand UO_2789 (O_2789,N_29815,N_29436);
xnor UO_2790 (O_2790,N_29956,N_29613);
xor UO_2791 (O_2791,N_29467,N_29878);
nor UO_2792 (O_2792,N_29643,N_29832);
and UO_2793 (O_2793,N_29515,N_29426);
or UO_2794 (O_2794,N_29408,N_29848);
and UO_2795 (O_2795,N_29533,N_29561);
nor UO_2796 (O_2796,N_29990,N_29660);
xor UO_2797 (O_2797,N_29691,N_29455);
xor UO_2798 (O_2798,N_29984,N_29957);
or UO_2799 (O_2799,N_29834,N_29521);
and UO_2800 (O_2800,N_29710,N_29551);
nand UO_2801 (O_2801,N_29860,N_29507);
or UO_2802 (O_2802,N_29515,N_29517);
nand UO_2803 (O_2803,N_29500,N_29738);
xnor UO_2804 (O_2804,N_29608,N_29927);
and UO_2805 (O_2805,N_29913,N_29617);
nand UO_2806 (O_2806,N_29997,N_29929);
xor UO_2807 (O_2807,N_29783,N_29712);
nor UO_2808 (O_2808,N_29593,N_29820);
xor UO_2809 (O_2809,N_29631,N_29674);
or UO_2810 (O_2810,N_29685,N_29994);
xnor UO_2811 (O_2811,N_29712,N_29899);
nand UO_2812 (O_2812,N_29935,N_29710);
nor UO_2813 (O_2813,N_29516,N_29762);
nor UO_2814 (O_2814,N_29524,N_29470);
nor UO_2815 (O_2815,N_29996,N_29600);
and UO_2816 (O_2816,N_29948,N_29956);
nor UO_2817 (O_2817,N_29743,N_29471);
nor UO_2818 (O_2818,N_29995,N_29948);
xnor UO_2819 (O_2819,N_29817,N_29440);
and UO_2820 (O_2820,N_29971,N_29428);
nor UO_2821 (O_2821,N_29486,N_29741);
or UO_2822 (O_2822,N_29463,N_29521);
and UO_2823 (O_2823,N_29537,N_29760);
nand UO_2824 (O_2824,N_29631,N_29491);
nor UO_2825 (O_2825,N_29559,N_29411);
and UO_2826 (O_2826,N_29762,N_29710);
and UO_2827 (O_2827,N_29499,N_29965);
nand UO_2828 (O_2828,N_29922,N_29492);
and UO_2829 (O_2829,N_29462,N_29444);
nor UO_2830 (O_2830,N_29433,N_29777);
nand UO_2831 (O_2831,N_29602,N_29729);
or UO_2832 (O_2832,N_29542,N_29637);
xnor UO_2833 (O_2833,N_29732,N_29882);
nand UO_2834 (O_2834,N_29654,N_29869);
nor UO_2835 (O_2835,N_29876,N_29440);
or UO_2836 (O_2836,N_29771,N_29519);
xor UO_2837 (O_2837,N_29643,N_29549);
and UO_2838 (O_2838,N_29496,N_29944);
xor UO_2839 (O_2839,N_29651,N_29886);
nand UO_2840 (O_2840,N_29689,N_29761);
nor UO_2841 (O_2841,N_29982,N_29599);
nand UO_2842 (O_2842,N_29762,N_29958);
nor UO_2843 (O_2843,N_29536,N_29449);
nand UO_2844 (O_2844,N_29691,N_29584);
nand UO_2845 (O_2845,N_29893,N_29582);
xor UO_2846 (O_2846,N_29579,N_29868);
xor UO_2847 (O_2847,N_29710,N_29782);
and UO_2848 (O_2848,N_29491,N_29605);
or UO_2849 (O_2849,N_29940,N_29485);
and UO_2850 (O_2850,N_29540,N_29682);
nand UO_2851 (O_2851,N_29862,N_29677);
nand UO_2852 (O_2852,N_29989,N_29971);
nand UO_2853 (O_2853,N_29826,N_29468);
nand UO_2854 (O_2854,N_29480,N_29898);
and UO_2855 (O_2855,N_29979,N_29937);
nor UO_2856 (O_2856,N_29847,N_29432);
xnor UO_2857 (O_2857,N_29846,N_29984);
nand UO_2858 (O_2858,N_29828,N_29888);
nand UO_2859 (O_2859,N_29919,N_29724);
and UO_2860 (O_2860,N_29466,N_29875);
xnor UO_2861 (O_2861,N_29664,N_29885);
xor UO_2862 (O_2862,N_29960,N_29676);
nor UO_2863 (O_2863,N_29782,N_29620);
nand UO_2864 (O_2864,N_29745,N_29729);
nor UO_2865 (O_2865,N_29949,N_29843);
nand UO_2866 (O_2866,N_29965,N_29405);
xor UO_2867 (O_2867,N_29928,N_29919);
nor UO_2868 (O_2868,N_29466,N_29511);
and UO_2869 (O_2869,N_29437,N_29773);
and UO_2870 (O_2870,N_29543,N_29451);
and UO_2871 (O_2871,N_29518,N_29475);
xor UO_2872 (O_2872,N_29604,N_29566);
xor UO_2873 (O_2873,N_29807,N_29545);
and UO_2874 (O_2874,N_29857,N_29793);
or UO_2875 (O_2875,N_29863,N_29492);
and UO_2876 (O_2876,N_29686,N_29704);
nand UO_2877 (O_2877,N_29422,N_29716);
nor UO_2878 (O_2878,N_29936,N_29621);
xnor UO_2879 (O_2879,N_29564,N_29897);
xor UO_2880 (O_2880,N_29939,N_29854);
nor UO_2881 (O_2881,N_29854,N_29610);
and UO_2882 (O_2882,N_29460,N_29667);
or UO_2883 (O_2883,N_29958,N_29658);
nand UO_2884 (O_2884,N_29493,N_29618);
nor UO_2885 (O_2885,N_29796,N_29925);
and UO_2886 (O_2886,N_29423,N_29463);
nor UO_2887 (O_2887,N_29858,N_29771);
or UO_2888 (O_2888,N_29531,N_29699);
or UO_2889 (O_2889,N_29612,N_29743);
and UO_2890 (O_2890,N_29723,N_29810);
or UO_2891 (O_2891,N_29940,N_29976);
xor UO_2892 (O_2892,N_29685,N_29485);
or UO_2893 (O_2893,N_29478,N_29836);
nor UO_2894 (O_2894,N_29794,N_29409);
or UO_2895 (O_2895,N_29678,N_29435);
xnor UO_2896 (O_2896,N_29624,N_29469);
and UO_2897 (O_2897,N_29865,N_29440);
and UO_2898 (O_2898,N_29810,N_29646);
or UO_2899 (O_2899,N_29832,N_29901);
or UO_2900 (O_2900,N_29781,N_29744);
xor UO_2901 (O_2901,N_29820,N_29675);
or UO_2902 (O_2902,N_29440,N_29830);
or UO_2903 (O_2903,N_29739,N_29428);
nand UO_2904 (O_2904,N_29690,N_29774);
xnor UO_2905 (O_2905,N_29470,N_29720);
xor UO_2906 (O_2906,N_29407,N_29417);
xnor UO_2907 (O_2907,N_29560,N_29866);
nor UO_2908 (O_2908,N_29832,N_29630);
nand UO_2909 (O_2909,N_29809,N_29957);
xor UO_2910 (O_2910,N_29852,N_29877);
nand UO_2911 (O_2911,N_29781,N_29789);
nand UO_2912 (O_2912,N_29494,N_29915);
xor UO_2913 (O_2913,N_29574,N_29551);
xnor UO_2914 (O_2914,N_29635,N_29577);
or UO_2915 (O_2915,N_29545,N_29564);
nand UO_2916 (O_2916,N_29945,N_29805);
xnor UO_2917 (O_2917,N_29546,N_29919);
nand UO_2918 (O_2918,N_29858,N_29475);
and UO_2919 (O_2919,N_29964,N_29645);
nand UO_2920 (O_2920,N_29521,N_29552);
nand UO_2921 (O_2921,N_29646,N_29861);
nor UO_2922 (O_2922,N_29724,N_29485);
nand UO_2923 (O_2923,N_29516,N_29571);
nand UO_2924 (O_2924,N_29579,N_29675);
xor UO_2925 (O_2925,N_29939,N_29473);
xnor UO_2926 (O_2926,N_29612,N_29770);
xor UO_2927 (O_2927,N_29787,N_29840);
nand UO_2928 (O_2928,N_29474,N_29661);
xnor UO_2929 (O_2929,N_29473,N_29529);
nand UO_2930 (O_2930,N_29544,N_29952);
and UO_2931 (O_2931,N_29987,N_29752);
nor UO_2932 (O_2932,N_29407,N_29968);
xnor UO_2933 (O_2933,N_29492,N_29546);
and UO_2934 (O_2934,N_29713,N_29621);
nor UO_2935 (O_2935,N_29480,N_29513);
nand UO_2936 (O_2936,N_29773,N_29675);
and UO_2937 (O_2937,N_29893,N_29959);
or UO_2938 (O_2938,N_29939,N_29872);
and UO_2939 (O_2939,N_29757,N_29632);
or UO_2940 (O_2940,N_29677,N_29865);
nor UO_2941 (O_2941,N_29535,N_29923);
xnor UO_2942 (O_2942,N_29682,N_29421);
or UO_2943 (O_2943,N_29872,N_29859);
nor UO_2944 (O_2944,N_29844,N_29679);
and UO_2945 (O_2945,N_29583,N_29686);
xor UO_2946 (O_2946,N_29860,N_29796);
or UO_2947 (O_2947,N_29654,N_29974);
nand UO_2948 (O_2948,N_29652,N_29989);
or UO_2949 (O_2949,N_29495,N_29596);
xnor UO_2950 (O_2950,N_29946,N_29992);
nor UO_2951 (O_2951,N_29707,N_29542);
or UO_2952 (O_2952,N_29838,N_29565);
and UO_2953 (O_2953,N_29895,N_29481);
nand UO_2954 (O_2954,N_29593,N_29516);
nor UO_2955 (O_2955,N_29537,N_29869);
nor UO_2956 (O_2956,N_29566,N_29645);
nor UO_2957 (O_2957,N_29730,N_29905);
xor UO_2958 (O_2958,N_29760,N_29675);
nor UO_2959 (O_2959,N_29422,N_29682);
xnor UO_2960 (O_2960,N_29625,N_29494);
or UO_2961 (O_2961,N_29887,N_29439);
nor UO_2962 (O_2962,N_29670,N_29761);
xnor UO_2963 (O_2963,N_29536,N_29637);
xnor UO_2964 (O_2964,N_29894,N_29705);
xnor UO_2965 (O_2965,N_29688,N_29459);
and UO_2966 (O_2966,N_29788,N_29442);
and UO_2967 (O_2967,N_29820,N_29585);
nor UO_2968 (O_2968,N_29868,N_29724);
xor UO_2969 (O_2969,N_29875,N_29984);
nor UO_2970 (O_2970,N_29725,N_29937);
nor UO_2971 (O_2971,N_29612,N_29912);
or UO_2972 (O_2972,N_29589,N_29819);
and UO_2973 (O_2973,N_29859,N_29791);
nand UO_2974 (O_2974,N_29444,N_29435);
xor UO_2975 (O_2975,N_29666,N_29598);
or UO_2976 (O_2976,N_29581,N_29424);
nor UO_2977 (O_2977,N_29894,N_29704);
nand UO_2978 (O_2978,N_29960,N_29705);
nor UO_2979 (O_2979,N_29860,N_29647);
nor UO_2980 (O_2980,N_29638,N_29603);
nand UO_2981 (O_2981,N_29477,N_29439);
nor UO_2982 (O_2982,N_29428,N_29792);
nand UO_2983 (O_2983,N_29543,N_29587);
nand UO_2984 (O_2984,N_29646,N_29696);
xor UO_2985 (O_2985,N_29461,N_29504);
nand UO_2986 (O_2986,N_29984,N_29660);
xor UO_2987 (O_2987,N_29626,N_29671);
and UO_2988 (O_2988,N_29451,N_29428);
and UO_2989 (O_2989,N_29688,N_29445);
and UO_2990 (O_2990,N_29442,N_29589);
nand UO_2991 (O_2991,N_29972,N_29782);
or UO_2992 (O_2992,N_29510,N_29997);
nand UO_2993 (O_2993,N_29868,N_29899);
xor UO_2994 (O_2994,N_29517,N_29621);
xnor UO_2995 (O_2995,N_29564,N_29633);
xor UO_2996 (O_2996,N_29996,N_29934);
nand UO_2997 (O_2997,N_29954,N_29577);
and UO_2998 (O_2998,N_29763,N_29745);
or UO_2999 (O_2999,N_29910,N_29463);
and UO_3000 (O_3000,N_29402,N_29438);
and UO_3001 (O_3001,N_29910,N_29871);
nor UO_3002 (O_3002,N_29679,N_29944);
xor UO_3003 (O_3003,N_29872,N_29837);
nor UO_3004 (O_3004,N_29688,N_29942);
and UO_3005 (O_3005,N_29960,N_29958);
or UO_3006 (O_3006,N_29499,N_29918);
nand UO_3007 (O_3007,N_29483,N_29430);
xor UO_3008 (O_3008,N_29443,N_29930);
nor UO_3009 (O_3009,N_29890,N_29781);
xnor UO_3010 (O_3010,N_29417,N_29727);
or UO_3011 (O_3011,N_29461,N_29875);
and UO_3012 (O_3012,N_29576,N_29773);
nor UO_3013 (O_3013,N_29490,N_29640);
xor UO_3014 (O_3014,N_29621,N_29703);
xnor UO_3015 (O_3015,N_29416,N_29899);
nand UO_3016 (O_3016,N_29502,N_29977);
nand UO_3017 (O_3017,N_29474,N_29876);
or UO_3018 (O_3018,N_29595,N_29718);
nand UO_3019 (O_3019,N_29462,N_29839);
xnor UO_3020 (O_3020,N_29593,N_29719);
nand UO_3021 (O_3021,N_29530,N_29803);
nor UO_3022 (O_3022,N_29981,N_29688);
xnor UO_3023 (O_3023,N_29993,N_29458);
nor UO_3024 (O_3024,N_29913,N_29885);
nand UO_3025 (O_3025,N_29491,N_29465);
xnor UO_3026 (O_3026,N_29958,N_29620);
nor UO_3027 (O_3027,N_29697,N_29979);
and UO_3028 (O_3028,N_29466,N_29513);
nand UO_3029 (O_3029,N_29715,N_29539);
or UO_3030 (O_3030,N_29619,N_29740);
nand UO_3031 (O_3031,N_29820,N_29967);
and UO_3032 (O_3032,N_29941,N_29407);
nand UO_3033 (O_3033,N_29409,N_29783);
nand UO_3034 (O_3034,N_29944,N_29710);
nor UO_3035 (O_3035,N_29420,N_29409);
xnor UO_3036 (O_3036,N_29904,N_29626);
nor UO_3037 (O_3037,N_29962,N_29417);
nor UO_3038 (O_3038,N_29466,N_29479);
and UO_3039 (O_3039,N_29846,N_29449);
nor UO_3040 (O_3040,N_29879,N_29672);
or UO_3041 (O_3041,N_29567,N_29471);
and UO_3042 (O_3042,N_29945,N_29899);
and UO_3043 (O_3043,N_29951,N_29537);
and UO_3044 (O_3044,N_29810,N_29800);
and UO_3045 (O_3045,N_29568,N_29645);
nor UO_3046 (O_3046,N_29537,N_29499);
nor UO_3047 (O_3047,N_29876,N_29913);
xnor UO_3048 (O_3048,N_29923,N_29750);
xor UO_3049 (O_3049,N_29867,N_29638);
xor UO_3050 (O_3050,N_29838,N_29769);
xor UO_3051 (O_3051,N_29826,N_29902);
nor UO_3052 (O_3052,N_29598,N_29900);
nor UO_3053 (O_3053,N_29580,N_29767);
or UO_3054 (O_3054,N_29406,N_29848);
or UO_3055 (O_3055,N_29548,N_29535);
xor UO_3056 (O_3056,N_29770,N_29654);
and UO_3057 (O_3057,N_29842,N_29726);
nor UO_3058 (O_3058,N_29572,N_29874);
or UO_3059 (O_3059,N_29641,N_29637);
or UO_3060 (O_3060,N_29803,N_29645);
nor UO_3061 (O_3061,N_29519,N_29943);
nor UO_3062 (O_3062,N_29954,N_29686);
xnor UO_3063 (O_3063,N_29477,N_29955);
nor UO_3064 (O_3064,N_29615,N_29688);
or UO_3065 (O_3065,N_29709,N_29577);
nand UO_3066 (O_3066,N_29989,N_29615);
and UO_3067 (O_3067,N_29556,N_29808);
nand UO_3068 (O_3068,N_29406,N_29751);
nor UO_3069 (O_3069,N_29552,N_29447);
xor UO_3070 (O_3070,N_29798,N_29837);
or UO_3071 (O_3071,N_29569,N_29921);
or UO_3072 (O_3072,N_29452,N_29737);
nor UO_3073 (O_3073,N_29936,N_29768);
and UO_3074 (O_3074,N_29521,N_29889);
nand UO_3075 (O_3075,N_29929,N_29861);
xor UO_3076 (O_3076,N_29916,N_29601);
xor UO_3077 (O_3077,N_29864,N_29463);
nor UO_3078 (O_3078,N_29734,N_29500);
nand UO_3079 (O_3079,N_29467,N_29533);
xor UO_3080 (O_3080,N_29658,N_29927);
or UO_3081 (O_3081,N_29939,N_29493);
or UO_3082 (O_3082,N_29793,N_29487);
and UO_3083 (O_3083,N_29670,N_29442);
or UO_3084 (O_3084,N_29938,N_29746);
nand UO_3085 (O_3085,N_29947,N_29624);
nand UO_3086 (O_3086,N_29625,N_29875);
and UO_3087 (O_3087,N_29759,N_29880);
nand UO_3088 (O_3088,N_29465,N_29698);
and UO_3089 (O_3089,N_29653,N_29633);
or UO_3090 (O_3090,N_29964,N_29793);
nand UO_3091 (O_3091,N_29865,N_29402);
nor UO_3092 (O_3092,N_29471,N_29927);
nor UO_3093 (O_3093,N_29593,N_29729);
and UO_3094 (O_3094,N_29752,N_29749);
and UO_3095 (O_3095,N_29861,N_29567);
and UO_3096 (O_3096,N_29788,N_29772);
and UO_3097 (O_3097,N_29970,N_29943);
and UO_3098 (O_3098,N_29776,N_29676);
or UO_3099 (O_3099,N_29814,N_29902);
xor UO_3100 (O_3100,N_29437,N_29557);
xor UO_3101 (O_3101,N_29496,N_29407);
nand UO_3102 (O_3102,N_29497,N_29871);
or UO_3103 (O_3103,N_29442,N_29527);
nor UO_3104 (O_3104,N_29713,N_29910);
nand UO_3105 (O_3105,N_29879,N_29840);
or UO_3106 (O_3106,N_29781,N_29513);
or UO_3107 (O_3107,N_29954,N_29872);
nand UO_3108 (O_3108,N_29995,N_29511);
xor UO_3109 (O_3109,N_29737,N_29661);
nor UO_3110 (O_3110,N_29606,N_29674);
and UO_3111 (O_3111,N_29630,N_29685);
or UO_3112 (O_3112,N_29695,N_29776);
or UO_3113 (O_3113,N_29716,N_29507);
nor UO_3114 (O_3114,N_29608,N_29821);
xor UO_3115 (O_3115,N_29438,N_29645);
nor UO_3116 (O_3116,N_29405,N_29540);
nand UO_3117 (O_3117,N_29961,N_29779);
nor UO_3118 (O_3118,N_29917,N_29971);
xnor UO_3119 (O_3119,N_29654,N_29555);
nand UO_3120 (O_3120,N_29731,N_29479);
or UO_3121 (O_3121,N_29560,N_29578);
nor UO_3122 (O_3122,N_29982,N_29544);
nand UO_3123 (O_3123,N_29688,N_29799);
nand UO_3124 (O_3124,N_29572,N_29744);
nor UO_3125 (O_3125,N_29813,N_29769);
or UO_3126 (O_3126,N_29914,N_29652);
or UO_3127 (O_3127,N_29415,N_29666);
xor UO_3128 (O_3128,N_29756,N_29834);
and UO_3129 (O_3129,N_29835,N_29727);
nor UO_3130 (O_3130,N_29595,N_29940);
nand UO_3131 (O_3131,N_29559,N_29684);
xor UO_3132 (O_3132,N_29977,N_29853);
or UO_3133 (O_3133,N_29741,N_29568);
xnor UO_3134 (O_3134,N_29405,N_29644);
xor UO_3135 (O_3135,N_29962,N_29575);
or UO_3136 (O_3136,N_29899,N_29464);
nor UO_3137 (O_3137,N_29504,N_29835);
and UO_3138 (O_3138,N_29514,N_29811);
or UO_3139 (O_3139,N_29909,N_29404);
nand UO_3140 (O_3140,N_29841,N_29958);
and UO_3141 (O_3141,N_29688,N_29784);
xor UO_3142 (O_3142,N_29613,N_29826);
nor UO_3143 (O_3143,N_29464,N_29806);
nor UO_3144 (O_3144,N_29938,N_29919);
nand UO_3145 (O_3145,N_29896,N_29471);
xor UO_3146 (O_3146,N_29810,N_29464);
nor UO_3147 (O_3147,N_29484,N_29805);
nand UO_3148 (O_3148,N_29505,N_29938);
and UO_3149 (O_3149,N_29498,N_29494);
or UO_3150 (O_3150,N_29714,N_29844);
or UO_3151 (O_3151,N_29605,N_29739);
or UO_3152 (O_3152,N_29510,N_29927);
or UO_3153 (O_3153,N_29554,N_29651);
nand UO_3154 (O_3154,N_29601,N_29501);
nand UO_3155 (O_3155,N_29543,N_29673);
xor UO_3156 (O_3156,N_29830,N_29986);
and UO_3157 (O_3157,N_29879,N_29497);
xnor UO_3158 (O_3158,N_29466,N_29478);
and UO_3159 (O_3159,N_29692,N_29407);
nor UO_3160 (O_3160,N_29485,N_29699);
nand UO_3161 (O_3161,N_29984,N_29891);
and UO_3162 (O_3162,N_29961,N_29928);
xor UO_3163 (O_3163,N_29603,N_29499);
nor UO_3164 (O_3164,N_29829,N_29830);
nor UO_3165 (O_3165,N_29611,N_29995);
nand UO_3166 (O_3166,N_29584,N_29552);
nor UO_3167 (O_3167,N_29540,N_29654);
nand UO_3168 (O_3168,N_29929,N_29613);
nand UO_3169 (O_3169,N_29698,N_29684);
and UO_3170 (O_3170,N_29753,N_29762);
nand UO_3171 (O_3171,N_29529,N_29810);
nor UO_3172 (O_3172,N_29915,N_29893);
and UO_3173 (O_3173,N_29425,N_29589);
nand UO_3174 (O_3174,N_29779,N_29997);
and UO_3175 (O_3175,N_29871,N_29539);
and UO_3176 (O_3176,N_29722,N_29798);
xor UO_3177 (O_3177,N_29541,N_29650);
or UO_3178 (O_3178,N_29996,N_29621);
or UO_3179 (O_3179,N_29619,N_29600);
or UO_3180 (O_3180,N_29833,N_29911);
or UO_3181 (O_3181,N_29904,N_29680);
xnor UO_3182 (O_3182,N_29485,N_29952);
and UO_3183 (O_3183,N_29915,N_29934);
nand UO_3184 (O_3184,N_29913,N_29620);
or UO_3185 (O_3185,N_29639,N_29920);
and UO_3186 (O_3186,N_29694,N_29766);
or UO_3187 (O_3187,N_29952,N_29890);
xor UO_3188 (O_3188,N_29820,N_29703);
nand UO_3189 (O_3189,N_29554,N_29580);
and UO_3190 (O_3190,N_29965,N_29839);
or UO_3191 (O_3191,N_29671,N_29678);
xor UO_3192 (O_3192,N_29778,N_29403);
or UO_3193 (O_3193,N_29743,N_29701);
xnor UO_3194 (O_3194,N_29888,N_29511);
and UO_3195 (O_3195,N_29973,N_29561);
and UO_3196 (O_3196,N_29525,N_29896);
and UO_3197 (O_3197,N_29909,N_29850);
and UO_3198 (O_3198,N_29658,N_29829);
nor UO_3199 (O_3199,N_29497,N_29690);
nor UO_3200 (O_3200,N_29534,N_29919);
xor UO_3201 (O_3201,N_29854,N_29601);
nor UO_3202 (O_3202,N_29736,N_29867);
and UO_3203 (O_3203,N_29404,N_29950);
and UO_3204 (O_3204,N_29718,N_29786);
nand UO_3205 (O_3205,N_29886,N_29454);
nor UO_3206 (O_3206,N_29988,N_29710);
nand UO_3207 (O_3207,N_29932,N_29760);
or UO_3208 (O_3208,N_29489,N_29476);
and UO_3209 (O_3209,N_29962,N_29794);
and UO_3210 (O_3210,N_29879,N_29953);
xor UO_3211 (O_3211,N_29778,N_29865);
and UO_3212 (O_3212,N_29565,N_29654);
nor UO_3213 (O_3213,N_29811,N_29549);
and UO_3214 (O_3214,N_29827,N_29605);
and UO_3215 (O_3215,N_29800,N_29519);
nand UO_3216 (O_3216,N_29897,N_29661);
and UO_3217 (O_3217,N_29585,N_29946);
and UO_3218 (O_3218,N_29624,N_29498);
or UO_3219 (O_3219,N_29815,N_29648);
nor UO_3220 (O_3220,N_29417,N_29484);
and UO_3221 (O_3221,N_29586,N_29434);
and UO_3222 (O_3222,N_29958,N_29991);
or UO_3223 (O_3223,N_29780,N_29987);
or UO_3224 (O_3224,N_29655,N_29786);
or UO_3225 (O_3225,N_29497,N_29846);
nand UO_3226 (O_3226,N_29545,N_29561);
nor UO_3227 (O_3227,N_29679,N_29930);
xnor UO_3228 (O_3228,N_29773,N_29523);
nor UO_3229 (O_3229,N_29429,N_29999);
and UO_3230 (O_3230,N_29872,N_29752);
and UO_3231 (O_3231,N_29745,N_29574);
and UO_3232 (O_3232,N_29931,N_29865);
nor UO_3233 (O_3233,N_29879,N_29797);
or UO_3234 (O_3234,N_29865,N_29988);
and UO_3235 (O_3235,N_29815,N_29427);
nand UO_3236 (O_3236,N_29467,N_29646);
xnor UO_3237 (O_3237,N_29451,N_29797);
nand UO_3238 (O_3238,N_29837,N_29448);
or UO_3239 (O_3239,N_29509,N_29925);
or UO_3240 (O_3240,N_29762,N_29671);
and UO_3241 (O_3241,N_29604,N_29790);
and UO_3242 (O_3242,N_29686,N_29859);
nor UO_3243 (O_3243,N_29904,N_29692);
nand UO_3244 (O_3244,N_29832,N_29440);
xor UO_3245 (O_3245,N_29969,N_29403);
nand UO_3246 (O_3246,N_29779,N_29862);
nand UO_3247 (O_3247,N_29936,N_29504);
xor UO_3248 (O_3248,N_29828,N_29944);
nand UO_3249 (O_3249,N_29988,N_29607);
and UO_3250 (O_3250,N_29870,N_29856);
nand UO_3251 (O_3251,N_29849,N_29867);
and UO_3252 (O_3252,N_29808,N_29790);
nand UO_3253 (O_3253,N_29540,N_29606);
or UO_3254 (O_3254,N_29815,N_29431);
or UO_3255 (O_3255,N_29401,N_29530);
nor UO_3256 (O_3256,N_29893,N_29756);
xnor UO_3257 (O_3257,N_29932,N_29835);
nor UO_3258 (O_3258,N_29912,N_29944);
and UO_3259 (O_3259,N_29582,N_29437);
xor UO_3260 (O_3260,N_29585,N_29728);
and UO_3261 (O_3261,N_29868,N_29433);
nand UO_3262 (O_3262,N_29465,N_29652);
and UO_3263 (O_3263,N_29833,N_29804);
nor UO_3264 (O_3264,N_29424,N_29993);
xnor UO_3265 (O_3265,N_29489,N_29978);
xnor UO_3266 (O_3266,N_29893,N_29906);
nor UO_3267 (O_3267,N_29446,N_29697);
or UO_3268 (O_3268,N_29563,N_29625);
and UO_3269 (O_3269,N_29814,N_29836);
nor UO_3270 (O_3270,N_29575,N_29905);
nand UO_3271 (O_3271,N_29928,N_29670);
and UO_3272 (O_3272,N_29676,N_29616);
xnor UO_3273 (O_3273,N_29417,N_29931);
or UO_3274 (O_3274,N_29999,N_29502);
or UO_3275 (O_3275,N_29719,N_29614);
or UO_3276 (O_3276,N_29705,N_29683);
or UO_3277 (O_3277,N_29491,N_29596);
nor UO_3278 (O_3278,N_29664,N_29757);
nand UO_3279 (O_3279,N_29836,N_29962);
nor UO_3280 (O_3280,N_29526,N_29466);
xnor UO_3281 (O_3281,N_29924,N_29780);
nor UO_3282 (O_3282,N_29771,N_29585);
or UO_3283 (O_3283,N_29955,N_29607);
nand UO_3284 (O_3284,N_29884,N_29845);
nor UO_3285 (O_3285,N_29840,N_29730);
xor UO_3286 (O_3286,N_29594,N_29839);
nand UO_3287 (O_3287,N_29525,N_29441);
nor UO_3288 (O_3288,N_29729,N_29629);
nand UO_3289 (O_3289,N_29629,N_29544);
xor UO_3290 (O_3290,N_29763,N_29591);
nand UO_3291 (O_3291,N_29941,N_29805);
and UO_3292 (O_3292,N_29469,N_29461);
nand UO_3293 (O_3293,N_29876,N_29457);
and UO_3294 (O_3294,N_29446,N_29861);
and UO_3295 (O_3295,N_29520,N_29506);
xor UO_3296 (O_3296,N_29666,N_29805);
or UO_3297 (O_3297,N_29631,N_29713);
nand UO_3298 (O_3298,N_29476,N_29504);
or UO_3299 (O_3299,N_29516,N_29811);
xor UO_3300 (O_3300,N_29459,N_29804);
and UO_3301 (O_3301,N_29934,N_29687);
and UO_3302 (O_3302,N_29934,N_29748);
and UO_3303 (O_3303,N_29787,N_29975);
xor UO_3304 (O_3304,N_29558,N_29847);
or UO_3305 (O_3305,N_29662,N_29691);
xnor UO_3306 (O_3306,N_29918,N_29413);
xor UO_3307 (O_3307,N_29889,N_29768);
xor UO_3308 (O_3308,N_29813,N_29424);
xor UO_3309 (O_3309,N_29988,N_29534);
xor UO_3310 (O_3310,N_29664,N_29531);
nand UO_3311 (O_3311,N_29815,N_29996);
or UO_3312 (O_3312,N_29481,N_29488);
or UO_3313 (O_3313,N_29588,N_29815);
and UO_3314 (O_3314,N_29671,N_29788);
nor UO_3315 (O_3315,N_29741,N_29767);
or UO_3316 (O_3316,N_29430,N_29835);
and UO_3317 (O_3317,N_29951,N_29623);
nor UO_3318 (O_3318,N_29988,N_29598);
and UO_3319 (O_3319,N_29489,N_29704);
nor UO_3320 (O_3320,N_29834,N_29791);
and UO_3321 (O_3321,N_29974,N_29446);
and UO_3322 (O_3322,N_29556,N_29400);
and UO_3323 (O_3323,N_29665,N_29437);
nor UO_3324 (O_3324,N_29910,N_29429);
nor UO_3325 (O_3325,N_29974,N_29583);
and UO_3326 (O_3326,N_29660,N_29512);
nor UO_3327 (O_3327,N_29865,N_29589);
and UO_3328 (O_3328,N_29650,N_29554);
nor UO_3329 (O_3329,N_29679,N_29757);
or UO_3330 (O_3330,N_29490,N_29456);
nor UO_3331 (O_3331,N_29662,N_29858);
or UO_3332 (O_3332,N_29883,N_29748);
xnor UO_3333 (O_3333,N_29691,N_29935);
nand UO_3334 (O_3334,N_29657,N_29708);
and UO_3335 (O_3335,N_29703,N_29701);
and UO_3336 (O_3336,N_29843,N_29625);
xor UO_3337 (O_3337,N_29463,N_29612);
xor UO_3338 (O_3338,N_29565,N_29756);
nor UO_3339 (O_3339,N_29902,N_29692);
nand UO_3340 (O_3340,N_29537,N_29490);
nand UO_3341 (O_3341,N_29669,N_29765);
nand UO_3342 (O_3342,N_29852,N_29565);
xor UO_3343 (O_3343,N_29907,N_29523);
and UO_3344 (O_3344,N_29787,N_29653);
xnor UO_3345 (O_3345,N_29557,N_29997);
nand UO_3346 (O_3346,N_29475,N_29784);
and UO_3347 (O_3347,N_29652,N_29709);
nor UO_3348 (O_3348,N_29766,N_29608);
xnor UO_3349 (O_3349,N_29585,N_29577);
and UO_3350 (O_3350,N_29697,N_29568);
nor UO_3351 (O_3351,N_29741,N_29504);
nand UO_3352 (O_3352,N_29933,N_29532);
xnor UO_3353 (O_3353,N_29923,N_29938);
or UO_3354 (O_3354,N_29992,N_29532);
xnor UO_3355 (O_3355,N_29640,N_29632);
nor UO_3356 (O_3356,N_29776,N_29638);
nor UO_3357 (O_3357,N_29980,N_29748);
and UO_3358 (O_3358,N_29445,N_29435);
or UO_3359 (O_3359,N_29712,N_29873);
xnor UO_3360 (O_3360,N_29789,N_29804);
nor UO_3361 (O_3361,N_29555,N_29595);
nand UO_3362 (O_3362,N_29769,N_29469);
and UO_3363 (O_3363,N_29651,N_29802);
nor UO_3364 (O_3364,N_29639,N_29642);
nand UO_3365 (O_3365,N_29944,N_29610);
nand UO_3366 (O_3366,N_29890,N_29561);
and UO_3367 (O_3367,N_29570,N_29488);
and UO_3368 (O_3368,N_29813,N_29500);
xnor UO_3369 (O_3369,N_29617,N_29514);
nor UO_3370 (O_3370,N_29624,N_29888);
xor UO_3371 (O_3371,N_29747,N_29655);
nand UO_3372 (O_3372,N_29716,N_29477);
nor UO_3373 (O_3373,N_29559,N_29895);
and UO_3374 (O_3374,N_29563,N_29692);
nor UO_3375 (O_3375,N_29497,N_29577);
or UO_3376 (O_3376,N_29901,N_29452);
xor UO_3377 (O_3377,N_29960,N_29455);
xor UO_3378 (O_3378,N_29983,N_29806);
nor UO_3379 (O_3379,N_29997,N_29946);
nand UO_3380 (O_3380,N_29811,N_29682);
xor UO_3381 (O_3381,N_29943,N_29480);
xnor UO_3382 (O_3382,N_29765,N_29492);
or UO_3383 (O_3383,N_29816,N_29624);
and UO_3384 (O_3384,N_29985,N_29950);
and UO_3385 (O_3385,N_29427,N_29961);
or UO_3386 (O_3386,N_29847,N_29662);
nand UO_3387 (O_3387,N_29433,N_29955);
nand UO_3388 (O_3388,N_29609,N_29692);
or UO_3389 (O_3389,N_29898,N_29709);
and UO_3390 (O_3390,N_29593,N_29500);
and UO_3391 (O_3391,N_29603,N_29561);
nor UO_3392 (O_3392,N_29496,N_29550);
and UO_3393 (O_3393,N_29760,N_29835);
and UO_3394 (O_3394,N_29492,N_29571);
nand UO_3395 (O_3395,N_29466,N_29831);
nand UO_3396 (O_3396,N_29445,N_29523);
xnor UO_3397 (O_3397,N_29980,N_29402);
nor UO_3398 (O_3398,N_29590,N_29588);
xnor UO_3399 (O_3399,N_29805,N_29806);
or UO_3400 (O_3400,N_29540,N_29908);
xnor UO_3401 (O_3401,N_29437,N_29973);
nand UO_3402 (O_3402,N_29448,N_29828);
and UO_3403 (O_3403,N_29939,N_29432);
xnor UO_3404 (O_3404,N_29400,N_29596);
nand UO_3405 (O_3405,N_29745,N_29527);
xor UO_3406 (O_3406,N_29795,N_29835);
and UO_3407 (O_3407,N_29525,N_29509);
nand UO_3408 (O_3408,N_29986,N_29591);
or UO_3409 (O_3409,N_29726,N_29873);
nand UO_3410 (O_3410,N_29681,N_29869);
and UO_3411 (O_3411,N_29631,N_29960);
and UO_3412 (O_3412,N_29815,N_29789);
xor UO_3413 (O_3413,N_29966,N_29412);
or UO_3414 (O_3414,N_29856,N_29515);
xor UO_3415 (O_3415,N_29821,N_29662);
nand UO_3416 (O_3416,N_29449,N_29615);
and UO_3417 (O_3417,N_29956,N_29523);
and UO_3418 (O_3418,N_29858,N_29683);
nand UO_3419 (O_3419,N_29476,N_29445);
nor UO_3420 (O_3420,N_29610,N_29500);
or UO_3421 (O_3421,N_29930,N_29772);
xor UO_3422 (O_3422,N_29599,N_29888);
nor UO_3423 (O_3423,N_29681,N_29576);
or UO_3424 (O_3424,N_29798,N_29669);
or UO_3425 (O_3425,N_29699,N_29888);
nor UO_3426 (O_3426,N_29726,N_29564);
nor UO_3427 (O_3427,N_29411,N_29621);
or UO_3428 (O_3428,N_29552,N_29800);
nand UO_3429 (O_3429,N_29771,N_29569);
nand UO_3430 (O_3430,N_29789,N_29639);
or UO_3431 (O_3431,N_29669,N_29809);
xor UO_3432 (O_3432,N_29688,N_29458);
xnor UO_3433 (O_3433,N_29837,N_29891);
nand UO_3434 (O_3434,N_29972,N_29850);
nor UO_3435 (O_3435,N_29796,N_29718);
xor UO_3436 (O_3436,N_29924,N_29493);
xnor UO_3437 (O_3437,N_29799,N_29738);
xnor UO_3438 (O_3438,N_29661,N_29874);
xnor UO_3439 (O_3439,N_29743,N_29726);
and UO_3440 (O_3440,N_29689,N_29434);
or UO_3441 (O_3441,N_29676,N_29586);
or UO_3442 (O_3442,N_29729,N_29926);
nand UO_3443 (O_3443,N_29560,N_29878);
nor UO_3444 (O_3444,N_29848,N_29732);
xnor UO_3445 (O_3445,N_29586,N_29618);
and UO_3446 (O_3446,N_29613,N_29690);
and UO_3447 (O_3447,N_29629,N_29598);
xnor UO_3448 (O_3448,N_29475,N_29721);
xor UO_3449 (O_3449,N_29534,N_29799);
or UO_3450 (O_3450,N_29763,N_29868);
nor UO_3451 (O_3451,N_29876,N_29516);
xor UO_3452 (O_3452,N_29807,N_29632);
nor UO_3453 (O_3453,N_29868,N_29465);
or UO_3454 (O_3454,N_29830,N_29507);
xnor UO_3455 (O_3455,N_29891,N_29885);
and UO_3456 (O_3456,N_29586,N_29514);
and UO_3457 (O_3457,N_29628,N_29783);
nor UO_3458 (O_3458,N_29914,N_29536);
xor UO_3459 (O_3459,N_29977,N_29655);
xor UO_3460 (O_3460,N_29653,N_29401);
nor UO_3461 (O_3461,N_29496,N_29948);
xnor UO_3462 (O_3462,N_29775,N_29800);
and UO_3463 (O_3463,N_29871,N_29864);
nand UO_3464 (O_3464,N_29564,N_29653);
nand UO_3465 (O_3465,N_29611,N_29533);
xnor UO_3466 (O_3466,N_29492,N_29709);
nand UO_3467 (O_3467,N_29477,N_29785);
and UO_3468 (O_3468,N_29871,N_29585);
nor UO_3469 (O_3469,N_29834,N_29735);
and UO_3470 (O_3470,N_29947,N_29800);
nor UO_3471 (O_3471,N_29534,N_29477);
xnor UO_3472 (O_3472,N_29583,N_29680);
and UO_3473 (O_3473,N_29657,N_29448);
nand UO_3474 (O_3474,N_29978,N_29861);
and UO_3475 (O_3475,N_29780,N_29614);
nor UO_3476 (O_3476,N_29668,N_29491);
xor UO_3477 (O_3477,N_29617,N_29917);
nor UO_3478 (O_3478,N_29418,N_29757);
nor UO_3479 (O_3479,N_29465,N_29691);
nor UO_3480 (O_3480,N_29550,N_29644);
or UO_3481 (O_3481,N_29582,N_29954);
nor UO_3482 (O_3482,N_29872,N_29527);
and UO_3483 (O_3483,N_29400,N_29818);
and UO_3484 (O_3484,N_29873,N_29648);
xor UO_3485 (O_3485,N_29698,N_29896);
or UO_3486 (O_3486,N_29603,N_29407);
xor UO_3487 (O_3487,N_29506,N_29894);
or UO_3488 (O_3488,N_29512,N_29458);
and UO_3489 (O_3489,N_29839,N_29921);
and UO_3490 (O_3490,N_29442,N_29840);
or UO_3491 (O_3491,N_29688,N_29881);
or UO_3492 (O_3492,N_29628,N_29702);
or UO_3493 (O_3493,N_29512,N_29505);
and UO_3494 (O_3494,N_29901,N_29991);
nand UO_3495 (O_3495,N_29549,N_29648);
or UO_3496 (O_3496,N_29836,N_29917);
xor UO_3497 (O_3497,N_29577,N_29664);
xnor UO_3498 (O_3498,N_29810,N_29428);
or UO_3499 (O_3499,N_29825,N_29454);
endmodule