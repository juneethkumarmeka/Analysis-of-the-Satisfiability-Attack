module basic_2000_20000_2500_25_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1004,In_270);
and U1 (N_1,In_1431,In_1732);
nand U2 (N_2,In_566,In_1779);
nand U3 (N_3,In_1644,In_570);
nor U4 (N_4,In_137,In_1029);
xnor U5 (N_5,In_609,In_1462);
nand U6 (N_6,In_1047,In_1436);
or U7 (N_7,In_719,In_1618);
and U8 (N_8,In_970,In_1061);
xnor U9 (N_9,In_1355,In_41);
nor U10 (N_10,In_728,In_1719);
or U11 (N_11,In_1095,In_356);
xor U12 (N_12,In_573,In_938);
and U13 (N_13,In_937,In_1681);
and U14 (N_14,In_1789,In_1999);
xor U15 (N_15,In_439,In_1115);
nand U16 (N_16,In_939,In_209);
or U17 (N_17,In_662,In_1149);
nor U18 (N_18,In_1476,In_1870);
or U19 (N_19,In_1888,In_614);
nand U20 (N_20,In_697,In_1545);
xor U21 (N_21,In_1552,In_1235);
or U22 (N_22,In_948,In_433);
and U23 (N_23,In_362,In_1464);
nand U24 (N_24,In_220,In_695);
or U25 (N_25,In_159,In_1030);
nand U26 (N_26,In_546,In_116);
nor U27 (N_27,In_920,In_1072);
or U28 (N_28,In_388,In_1676);
nor U29 (N_29,In_1786,In_1829);
xor U30 (N_30,In_815,In_967);
nand U31 (N_31,In_1527,In_124);
and U32 (N_32,In_1494,In_637);
nor U33 (N_33,In_480,In_1682);
xnor U34 (N_34,In_1725,In_419);
xnor U35 (N_35,In_1271,In_361);
nor U36 (N_36,In_1643,In_942);
nor U37 (N_37,In_1289,In_468);
nand U38 (N_38,In_1019,In_1743);
nor U39 (N_39,In_454,In_1435);
and U40 (N_40,In_77,In_1112);
nand U41 (N_41,In_1420,In_1210);
or U42 (N_42,In_615,In_422);
xnor U43 (N_43,In_1784,In_758);
nand U44 (N_44,In_1157,In_10);
and U45 (N_45,In_223,In_24);
xor U46 (N_46,In_997,In_12);
or U47 (N_47,In_1066,In_909);
or U48 (N_48,In_1317,In_1724);
nand U49 (N_49,In_814,In_1071);
and U50 (N_50,In_371,In_1553);
and U51 (N_51,In_389,In_868);
or U52 (N_52,In_1814,In_1300);
xor U53 (N_53,In_1600,In_976);
and U54 (N_54,In_803,In_1524);
nor U55 (N_55,In_230,In_1642);
nand U56 (N_56,In_1109,In_1002);
nor U57 (N_57,In_1148,In_1150);
and U58 (N_58,In_1983,In_996);
nand U59 (N_59,In_375,In_1986);
or U60 (N_60,In_114,In_1329);
nand U61 (N_61,In_1890,In_737);
or U62 (N_62,In_1469,In_1201);
nand U63 (N_63,In_105,In_608);
nand U64 (N_64,In_430,In_1224);
xnor U65 (N_65,In_1914,In_743);
nand U66 (N_66,In_723,In_485);
or U67 (N_67,In_1141,In_1144);
xor U68 (N_68,In_1471,In_515);
or U69 (N_69,In_1873,In_1186);
and U70 (N_70,In_139,In_1176);
xnor U71 (N_71,In_1972,In_765);
nand U72 (N_72,In_108,In_1933);
and U73 (N_73,In_796,In_1470);
nand U74 (N_74,In_953,In_67);
nor U75 (N_75,In_613,In_1799);
or U76 (N_76,In_1065,In_530);
or U77 (N_77,In_1133,In_880);
nor U78 (N_78,In_23,In_1119);
nand U79 (N_79,In_238,In_1415);
nor U80 (N_80,In_1497,In_1231);
and U81 (N_81,In_1008,In_556);
nor U82 (N_82,In_1191,In_1465);
xnor U83 (N_83,In_150,In_1882);
nor U84 (N_84,In_951,In_256);
nand U85 (N_85,In_869,In_1493);
and U86 (N_86,In_1121,In_1569);
and U87 (N_87,In_1969,In_376);
or U88 (N_88,In_331,In_1542);
or U89 (N_89,In_828,In_1632);
xor U90 (N_90,In_604,In_1174);
and U91 (N_91,In_755,In_1843);
and U92 (N_92,In_821,In_208);
and U93 (N_93,In_1484,In_456);
or U94 (N_94,In_1684,In_1889);
nand U95 (N_95,In_1874,In_739);
nor U96 (N_96,In_1306,In_500);
xor U97 (N_97,In_1871,In_1366);
nor U98 (N_98,In_807,In_1404);
nor U99 (N_99,In_450,In_1909);
nor U100 (N_100,In_287,In_146);
nand U101 (N_101,In_777,In_1380);
nand U102 (N_102,In_1111,In_1661);
or U103 (N_103,In_427,In_1279);
xnor U104 (N_104,In_104,In_340);
and U105 (N_105,In_28,In_25);
nand U106 (N_106,In_269,In_1816);
xnor U107 (N_107,In_1190,In_1383);
nand U108 (N_108,In_1165,In_1568);
or U109 (N_109,In_1713,In_1537);
xnor U110 (N_110,In_883,In_636);
nor U111 (N_111,In_1802,In_1158);
xnor U112 (N_112,In_235,In_464);
or U113 (N_113,In_959,In_1244);
nand U114 (N_114,In_543,In_1063);
or U115 (N_115,In_369,In_1598);
or U116 (N_116,In_972,In_113);
nand U117 (N_117,In_517,In_1624);
xnor U118 (N_118,In_15,In_1260);
nor U119 (N_119,In_1280,In_1045);
nand U120 (N_120,In_1345,In_1987);
and U121 (N_121,In_1297,In_1594);
or U122 (N_122,In_62,In_804);
or U123 (N_123,In_1502,In_1204);
and U124 (N_124,In_479,In_156);
xor U125 (N_125,In_1920,In_866);
and U126 (N_126,In_277,In_179);
or U127 (N_127,In_386,In_467);
xor U128 (N_128,In_483,In_761);
nor U129 (N_129,In_887,In_335);
nand U130 (N_130,In_1589,In_805);
xnor U131 (N_131,In_1532,In_696);
and U132 (N_132,In_1267,In_1769);
or U133 (N_133,In_710,In_94);
nand U134 (N_134,In_3,In_347);
xor U135 (N_135,In_452,In_503);
nand U136 (N_136,In_720,In_1685);
nand U137 (N_137,In_1400,In_73);
nor U138 (N_138,In_1183,In_1722);
and U139 (N_139,In_1671,In_1391);
and U140 (N_140,In_1554,In_1012);
xnor U141 (N_141,In_961,In_1284);
nor U142 (N_142,In_1927,In_32);
and U143 (N_143,In_1822,In_22);
or U144 (N_144,In_1641,In_1525);
nand U145 (N_145,In_1790,In_603);
nor U146 (N_146,In_158,In_1707);
nor U147 (N_147,In_586,In_706);
nand U148 (N_148,In_445,In_245);
and U149 (N_149,In_1311,In_1766);
xor U150 (N_150,In_1339,In_1556);
xnor U151 (N_151,In_1935,In_1302);
xnor U152 (N_152,In_559,In_523);
and U153 (N_153,In_487,In_436);
and U154 (N_154,In_1526,In_472);
or U155 (N_155,In_244,In_1372);
and U156 (N_156,In_1529,In_1978);
nand U157 (N_157,In_342,In_1474);
or U158 (N_158,In_1023,In_1377);
nor U159 (N_159,In_992,In_749);
nor U160 (N_160,In_329,In_325);
nand U161 (N_161,In_1084,In_820);
or U162 (N_162,In_308,In_687);
xor U163 (N_163,In_492,In_63);
nand U164 (N_164,In_1196,In_1636);
or U165 (N_165,In_644,In_1450);
and U166 (N_166,In_1958,In_1916);
nor U167 (N_167,In_1374,In_628);
xor U168 (N_168,In_750,In_1197);
and U169 (N_169,In_1562,In_1699);
or U170 (N_170,In_1437,In_1804);
nor U171 (N_171,In_53,In_1336);
xnor U172 (N_172,In_395,In_178);
nand U173 (N_173,In_1155,In_1495);
nor U174 (N_174,In_1659,In_1467);
xor U175 (N_175,In_1513,In_567);
and U176 (N_176,In_213,In_120);
xor U177 (N_177,In_1223,In_1102);
nor U178 (N_178,In_518,In_1209);
xor U179 (N_179,In_1396,In_438);
and U180 (N_180,In_634,In_0);
nor U181 (N_181,In_1670,In_411);
nand U182 (N_182,In_1832,In_396);
nand U183 (N_183,In_971,In_571);
and U184 (N_184,In_501,In_656);
xor U185 (N_185,In_840,In_1511);
and U186 (N_186,In_1950,In_1473);
nor U187 (N_187,In_966,In_1550);
and U188 (N_188,In_1449,In_1098);
xnor U189 (N_189,In_228,In_536);
xnor U190 (N_190,In_425,In_877);
xnor U191 (N_191,In_237,In_551);
or U192 (N_192,In_92,In_1427);
or U193 (N_193,In_1205,In_198);
nor U194 (N_194,In_888,In_1357);
xor U195 (N_195,In_694,In_384);
nand U196 (N_196,In_254,In_1451);
nand U197 (N_197,In_1973,In_381);
xor U198 (N_198,In_1519,In_1033);
and U199 (N_199,In_1240,In_393);
nor U200 (N_200,In_1479,In_58);
xnor U201 (N_201,In_314,In_688);
nand U202 (N_202,In_1964,In_257);
or U203 (N_203,In_838,In_1337);
nand U204 (N_204,In_713,In_304);
nand U205 (N_205,In_1386,In_1831);
nand U206 (N_206,In_1412,In_236);
nand U207 (N_207,In_1359,In_811);
or U208 (N_208,In_1487,In_177);
and U209 (N_209,In_1960,In_185);
and U210 (N_210,In_1514,In_444);
xor U211 (N_211,In_1957,In_36);
xnor U212 (N_212,In_1664,In_1665);
xnor U213 (N_213,In_1937,In_404);
or U214 (N_214,In_572,In_1988);
and U215 (N_215,In_635,In_933);
and U216 (N_216,In_339,In_372);
or U217 (N_217,In_654,In_852);
nor U218 (N_218,In_1602,In_1215);
and U219 (N_219,In_1152,In_1965);
and U220 (N_220,In_884,In_311);
or U221 (N_221,In_537,In_1915);
nor U222 (N_222,In_771,In_75);
and U223 (N_223,In_207,In_1801);
xnor U224 (N_224,In_272,In_1567);
or U225 (N_225,In_1895,In_1696);
and U226 (N_226,In_1859,In_798);
xnor U227 (N_227,In_562,In_1884);
or U228 (N_228,In_1839,In_867);
xnor U229 (N_229,In_786,In_526);
nor U230 (N_230,In_629,In_157);
and U231 (N_231,In_923,In_831);
xnor U232 (N_232,In_1857,In_215);
and U233 (N_233,In_169,In_56);
nor U234 (N_234,In_851,In_931);
or U235 (N_235,In_1040,In_239);
nor U236 (N_236,In_957,In_847);
and U237 (N_237,In_509,In_962);
nand U238 (N_238,In_736,In_1765);
and U239 (N_239,In_1118,In_1264);
and U240 (N_240,In_1154,In_789);
nand U241 (N_241,In_1227,In_1947);
or U242 (N_242,In_1213,In_1130);
and U243 (N_243,In_1961,In_1295);
or U244 (N_244,In_1747,In_206);
nor U245 (N_245,In_310,In_529);
and U246 (N_246,In_494,In_908);
and U247 (N_247,In_46,In_872);
or U248 (N_248,In_398,In_1352);
or U249 (N_249,In_733,In_544);
xor U250 (N_250,In_1423,In_281);
xor U251 (N_251,In_471,In_1089);
nand U252 (N_252,In_31,In_1499);
and U253 (N_253,In_1277,In_320);
and U254 (N_254,In_300,In_1202);
nor U255 (N_255,In_1036,In_845);
nor U256 (N_256,In_752,In_1614);
nor U257 (N_257,In_1031,In_1597);
xnor U258 (N_258,In_1698,In_447);
or U259 (N_259,In_585,In_597);
or U260 (N_260,In_1419,In_886);
xor U261 (N_261,In_1561,In_940);
xnor U262 (N_262,In_1875,In_193);
and U263 (N_263,In_1037,In_252);
nor U264 (N_264,In_1523,In_4);
and U265 (N_265,In_1193,In_240);
nand U266 (N_266,In_476,In_1966);
xor U267 (N_267,In_1485,In_1821);
and U268 (N_268,In_1516,In_1251);
nor U269 (N_269,In_850,In_1243);
xor U270 (N_270,In_1869,In_1207);
and U271 (N_271,In_588,In_1924);
xor U272 (N_272,In_1100,In_258);
nor U273 (N_273,In_598,In_1269);
nor U274 (N_274,In_1990,In_1222);
or U275 (N_275,In_1335,In_1912);
nand U276 (N_276,In_683,In_377);
xor U277 (N_277,In_892,In_1997);
xnor U278 (N_278,In_283,In_186);
nand U279 (N_279,In_1541,In_1265);
and U280 (N_280,In_741,In_627);
xnor U281 (N_281,In_459,In_1233);
and U282 (N_282,In_1456,In_1563);
or U283 (N_283,In_1667,In_1880);
or U284 (N_284,In_623,In_893);
xor U285 (N_285,In_165,In_735);
or U286 (N_286,In_865,In_85);
xor U287 (N_287,In_881,In_1482);
and U288 (N_288,In_1077,In_904);
nor U289 (N_289,In_1086,In_776);
nand U290 (N_290,In_1078,In_1605);
and U291 (N_291,In_1830,In_547);
nor U292 (N_292,In_1778,In_1395);
nand U293 (N_293,In_1225,In_147);
xor U294 (N_294,In_11,In_166);
and U295 (N_295,In_1901,In_1448);
xnor U296 (N_296,In_751,In_763);
or U297 (N_297,In_412,In_936);
or U298 (N_298,In_44,In_344);
and U299 (N_299,In_1310,In_1211);
nor U300 (N_300,In_1576,In_790);
xor U301 (N_301,In_461,In_793);
and U302 (N_302,In_68,In_1468);
and U303 (N_303,In_1261,In_373);
and U304 (N_304,In_1020,In_1087);
xnor U305 (N_305,In_138,In_652);
nand U306 (N_306,In_1459,In_1447);
nand U307 (N_307,In_1740,In_1807);
or U308 (N_308,In_301,In_1143);
or U309 (N_309,In_407,In_856);
xor U310 (N_310,In_168,In_1728);
xnor U311 (N_311,In_1976,In_1793);
nand U312 (N_312,In_1985,In_1863);
and U313 (N_313,In_397,In_69);
nand U314 (N_314,In_592,In_1236);
nand U315 (N_315,In_918,In_343);
and U316 (N_316,In_975,In_899);
nor U317 (N_317,In_1268,In_246);
or U318 (N_318,In_1263,In_1745);
nor U319 (N_319,In_1534,In_675);
or U320 (N_320,In_1586,In_1628);
and U321 (N_321,In_1139,In_729);
or U322 (N_322,In_1738,In_705);
nor U323 (N_323,In_1539,In_1134);
and U324 (N_324,In_271,In_650);
nand U325 (N_325,In_33,In_410);
nor U326 (N_326,In_400,In_1281);
nor U327 (N_327,In_1005,In_1257);
nand U328 (N_328,In_401,In_1906);
or U329 (N_329,In_91,In_646);
or U330 (N_330,In_112,In_1866);
nor U331 (N_331,In_968,In_1616);
and U332 (N_332,In_276,In_101);
nand U333 (N_333,In_7,In_1585);
and U334 (N_334,In_357,In_1818);
nor U335 (N_335,In_191,In_1619);
and U336 (N_336,In_837,In_941);
and U337 (N_337,In_1989,In_764);
nor U338 (N_338,In_553,In_292);
and U339 (N_339,In_717,In_382);
xnor U340 (N_340,In_14,In_1107);
nand U341 (N_341,In_16,In_1848);
nand U342 (N_342,In_1823,In_1825);
xor U343 (N_343,In_93,In_1457);
nor U344 (N_344,In_1810,In_1188);
nand U345 (N_345,In_135,In_1504);
nand U346 (N_346,In_1051,In_1373);
nand U347 (N_347,In_1893,In_1852);
xnor U348 (N_348,In_234,In_374);
nor U349 (N_349,In_895,In_1056);
xor U350 (N_350,In_921,In_879);
or U351 (N_351,In_1575,In_1027);
xnor U352 (N_352,In_714,In_1613);
or U353 (N_353,In_1518,In_1757);
xor U354 (N_354,In_988,In_1646);
nand U355 (N_355,In_1153,In_651);
and U356 (N_356,In_72,In_1623);
nor U357 (N_357,In_99,In_1455);
nor U358 (N_358,In_1414,In_721);
nor U359 (N_359,In_784,In_582);
or U360 (N_360,In_708,In_666);
or U361 (N_361,In_1840,In_296);
and U362 (N_362,In_816,In_1371);
nand U363 (N_363,In_1416,In_1198);
xnor U364 (N_364,In_225,In_660);
nor U365 (N_365,In_1291,In_1606);
or U366 (N_366,In_825,In_192);
or U367 (N_367,In_1797,In_1967);
xor U368 (N_368,In_1746,In_1813);
or U369 (N_369,In_1774,In_1543);
nor U370 (N_370,In_986,In_1445);
and U371 (N_371,In_1409,In_1126);
nand U372 (N_372,In_348,In_1160);
and U373 (N_373,In_605,In_218);
nand U374 (N_374,In_385,In_744);
nand U375 (N_375,In_291,In_1424);
or U376 (N_376,In_1686,In_745);
nand U377 (N_377,In_1853,In_183);
nor U378 (N_378,In_1753,In_1060);
or U379 (N_379,In_889,In_611);
or U380 (N_380,In_1483,In_201);
and U381 (N_381,In_409,In_1142);
or U382 (N_382,In_143,In_1610);
nor U383 (N_383,In_1577,In_943);
and U384 (N_384,In_1252,In_1410);
or U385 (N_385,In_111,In_1919);
nand U386 (N_386,In_1105,In_1708);
or U387 (N_387,In_1730,In_282);
and U388 (N_388,In_863,In_1953);
nor U389 (N_389,In_699,In_435);
nand U390 (N_390,In_328,In_1551);
nand U391 (N_391,In_1764,In_1718);
xor U392 (N_392,In_1253,In_315);
xnor U393 (N_393,In_919,In_1016);
nor U394 (N_394,In_1255,In_1320);
nor U395 (N_395,In_1171,In_1695);
and U396 (N_396,In_742,In_993);
nand U397 (N_397,In_359,In_658);
nand U398 (N_398,In_1385,In_1248);
nor U399 (N_399,In_30,In_698);
xnor U400 (N_400,In_1305,In_273);
xnor U401 (N_401,In_580,In_560);
and U402 (N_402,In_1220,In_1630);
nor U403 (N_403,In_875,In_1940);
and U404 (N_404,In_229,In_999);
or U405 (N_405,In_1481,In_224);
and U406 (N_406,In_1206,In_1792);
or U407 (N_407,In_730,In_1101);
and U408 (N_408,In_496,In_1566);
nor U409 (N_409,In_189,In_1785);
nand U410 (N_410,In_643,In_1422);
nand U411 (N_411,In_337,In_1540);
and U412 (N_412,In_17,In_754);
and U413 (N_413,In_153,In_5);
nand U414 (N_414,In_414,In_1170);
nand U415 (N_415,In_1748,In_122);
nand U416 (N_416,In_274,In_915);
and U417 (N_417,In_1073,In_358);
and U418 (N_418,In_154,In_1921);
nand U419 (N_419,In_475,In_1454);
xnor U420 (N_420,In_1315,In_647);
or U421 (N_421,In_497,In_1234);
nor U422 (N_422,In_279,In_1900);
and U423 (N_423,In_606,In_1788);
nor U424 (N_424,In_1313,In_669);
nand U425 (N_425,In_1181,In_136);
nor U426 (N_426,In_1783,In_295);
nor U427 (N_427,In_1717,In_1894);
nand U428 (N_428,In_724,In_498);
and U429 (N_429,In_1138,In_760);
nor U430 (N_430,In_405,In_1634);
nand U431 (N_431,In_1998,In_87);
nor U432 (N_432,In_1035,In_1951);
nand U433 (N_433,In_955,In_649);
nor U434 (N_434,In_1808,In_341);
nor U435 (N_435,In_286,In_1057);
nand U436 (N_436,In_1677,In_221);
nand U437 (N_437,In_704,In_74);
or U438 (N_438,In_1607,In_896);
and U439 (N_439,In_925,In_1530);
and U440 (N_440,In_693,In_554);
nand U441 (N_441,In_1262,In_1573);
and U442 (N_442,In_248,In_1603);
nor U443 (N_443,In_1342,In_1944);
or U444 (N_444,In_1876,In_1275);
and U445 (N_445,In_510,In_312);
nand U446 (N_446,In_575,In_934);
or U447 (N_447,In_1425,In_190);
xor U448 (N_448,In_1058,In_668);
or U449 (N_449,In_781,In_859);
and U450 (N_450,In_545,In_1819);
nand U451 (N_451,In_1347,In_1461);
or U452 (N_452,In_8,In_211);
or U453 (N_453,In_259,In_1564);
or U454 (N_454,In_794,In_1129);
nand U455 (N_455,In_928,In_1941);
nor U456 (N_456,In_1963,In_1434);
or U457 (N_457,In_1403,In_505);
nor U458 (N_458,In_672,In_1907);
or U459 (N_459,In_1712,In_1164);
and U460 (N_460,In_806,In_1382);
nor U461 (N_461,In_1715,In_1147);
or U462 (N_462,In_1096,In_1929);
xnor U463 (N_463,In_1787,In_1544);
xnor U464 (N_464,In_149,In_770);
and U465 (N_465,In_443,In_1506);
and U466 (N_466,In_200,In_1136);
or U467 (N_467,In_474,In_1421);
or U468 (N_468,In_772,In_490);
and U469 (N_469,In_1446,In_214);
or U470 (N_470,In_565,In_19);
or U471 (N_471,In_1582,In_1307);
and U472 (N_472,In_1599,In_1656);
or U473 (N_473,In_365,In_1418);
xor U474 (N_474,In_963,In_679);
nand U475 (N_475,In_1392,In_1943);
and U476 (N_476,In_57,In_125);
xor U477 (N_477,In_1872,In_834);
nor U478 (N_478,In_413,In_1923);
and U479 (N_479,In_1156,In_6);
nand U480 (N_480,In_1453,In_929);
xor U481 (N_481,In_685,In_801);
nor U482 (N_482,In_979,In_1555);
xnor U483 (N_483,In_1500,In_1322);
or U484 (N_484,In_1074,In_460);
and U485 (N_485,In_368,In_1817);
or U486 (N_486,In_1104,In_1756);
nand U487 (N_487,In_164,In_1120);
xnor U488 (N_488,In_1510,In_489);
and U489 (N_489,In_1127,In_118);
or U490 (N_490,In_620,In_1675);
xor U491 (N_491,In_659,In_973);
nor U492 (N_492,In_1521,In_533);
or U493 (N_493,In_1678,In_351);
nand U494 (N_494,In_1496,In_1574);
nand U495 (N_495,In_1179,In_1388);
nand U496 (N_496,In_1674,In_1159);
xnor U497 (N_497,In_1535,In_148);
nor U498 (N_498,In_521,In_493);
and U499 (N_499,In_550,In_21);
nor U500 (N_500,In_1680,In_1798);
or U501 (N_501,In_1203,In_528);
nand U502 (N_502,In_1938,In_232);
and U503 (N_503,In_579,In_1498);
nor U504 (N_504,In_1655,In_355);
and U505 (N_505,In_352,In_1861);
nand U506 (N_506,In_601,In_1137);
or U507 (N_507,In_525,In_981);
nand U508 (N_508,In_52,In_1595);
and U509 (N_509,In_552,In_76);
or U510 (N_510,In_1440,In_1601);
xnor U511 (N_511,In_568,In_1749);
nor U512 (N_512,In_1184,In_703);
and U513 (N_513,In_1172,In_1741);
nor U514 (N_514,In_326,In_60);
nor U515 (N_515,In_1701,In_1917);
and U516 (N_516,In_1736,In_1579);
and U517 (N_517,In_1549,In_1835);
nand U518 (N_518,In_162,In_1316);
or U519 (N_519,In_1367,In_690);
xnor U520 (N_520,In_383,In_1490);
nor U521 (N_521,In_416,In_1565);
xor U522 (N_522,In_1114,In_1982);
xor U523 (N_523,In_455,In_1581);
xnor U524 (N_524,In_624,In_511);
or U525 (N_525,In_1508,In_902);
nor U526 (N_526,In_226,In_1097);
nor U527 (N_527,In_1851,In_1343);
nor U528 (N_528,In_1113,In_563);
xnor U529 (N_529,In_1276,In_1411);
nor U530 (N_530,In_1522,In_79);
nand U531 (N_531,In_1013,In_944);
xnor U532 (N_532,In_1723,In_1024);
xor U533 (N_533,In_1520,In_266);
and U534 (N_534,In_1956,In_1480);
and U535 (N_535,In_299,In_1228);
or U536 (N_536,In_1489,In_1079);
or U537 (N_537,In_394,In_1389);
or U538 (N_538,In_1885,In_1854);
and U539 (N_539,In_621,In_1195);
nand U540 (N_540,In_431,In_1844);
and U541 (N_541,In_830,In_59);
or U542 (N_542,In_670,In_1402);
or U543 (N_543,In_633,In_1083);
nor U544 (N_544,In_788,In_1583);
xor U545 (N_545,In_524,In_227);
and U546 (N_546,In_1216,In_663);
or U547 (N_547,In_709,In_1332);
and U548 (N_548,In_391,In_268);
nor U549 (N_549,In_1358,In_469);
nand U550 (N_550,In_462,In_906);
nand U551 (N_551,In_898,In_1596);
and U552 (N_552,In_964,In_1363);
nand U553 (N_553,In_421,In_50);
or U554 (N_554,In_1076,In_332);
xnor U555 (N_555,In_1841,In_330);
and U556 (N_556,In_914,In_140);
xor U557 (N_557,In_1131,In_160);
and U558 (N_558,In_1794,In_451);
and U559 (N_559,In_1401,In_989);
nor U560 (N_560,In_1587,In_618);
xnor U561 (N_561,In_1633,In_1175);
xnor U562 (N_562,In_1046,In_819);
and U563 (N_563,In_453,In_1980);
nand U564 (N_564,In_1826,In_426);
nor U565 (N_565,In_345,In_1761);
or U566 (N_566,In_558,In_1417);
nor U567 (N_567,In_594,In_826);
and U568 (N_568,In_130,In_774);
or U569 (N_569,In_861,In_1731);
nand U570 (N_570,In_791,In_54);
or U571 (N_571,In_1286,In_1936);
nor U572 (N_572,In_1501,In_1334);
nor U573 (N_573,In_222,In_1673);
or U574 (N_574,In_1365,In_1845);
nor U575 (N_575,In_1959,In_121);
xor U576 (N_576,In_506,In_1653);
and U577 (N_577,In_1691,In_862);
nor U578 (N_578,In_1772,In_1879);
nand U579 (N_579,In_1803,In_1727);
nand U580 (N_580,In_1700,In_1625);
or U581 (N_581,In_1654,In_141);
xnor U582 (N_582,In_1742,In_1250);
nand U583 (N_583,In_1330,In_602);
nor U584 (N_584,In_366,In_96);
or U585 (N_585,In_1608,In_1621);
or U586 (N_586,In_1189,In_477);
xor U587 (N_587,In_1928,In_734);
nand U588 (N_588,In_18,In_34);
and U589 (N_589,In_1883,In_639);
and U590 (N_590,In_134,In_202);
or U591 (N_591,In_243,In_1229);
xor U592 (N_592,In_1631,In_495);
nor U593 (N_593,In_950,In_673);
nand U594 (N_594,In_638,In_870);
nand U595 (N_595,In_1278,In_1734);
and U596 (N_596,In_738,In_876);
and U597 (N_597,In_231,In_1232);
and U598 (N_598,In_1390,In_1546);
xnor U599 (N_599,In_1393,In_1571);
nand U600 (N_600,In_849,In_1617);
and U601 (N_601,In_309,In_930);
xnor U602 (N_602,In_903,In_625);
nor U603 (N_603,In_1351,In_499);
nor U604 (N_604,In_1081,In_1706);
nor U605 (N_605,In_370,In_747);
and U606 (N_606,In_1026,In_289);
xnor U607 (N_607,In_1992,In_1006);
xnor U608 (N_608,In_641,In_1770);
nor U609 (N_609,In_1294,In_466);
and U610 (N_610,In_255,In_1809);
nor U611 (N_611,In_1834,In_1626);
nand U612 (N_612,In_1399,In_718);
or U613 (N_613,In_1572,In_1259);
or U614 (N_614,In_1751,In_127);
nand U615 (N_615,In_616,In_1782);
or U616 (N_616,In_1000,In_1239);
xnor U617 (N_617,In_64,In_1820);
and U618 (N_618,In_110,In_1292);
or U619 (N_619,In_1217,In_653);
or U620 (N_620,In_319,In_1948);
and U621 (N_621,In_133,In_418);
nor U622 (N_622,In_1258,In_1931);
xnor U623 (N_623,In_1318,In_1735);
nand U624 (N_624,In_132,In_894);
nand U625 (N_625,In_655,In_917);
nand U626 (N_626,In_1693,In_701);
xnor U627 (N_627,In_549,In_767);
xnor U628 (N_628,In_583,In_491);
nor U629 (N_629,In_293,In_1652);
nand U630 (N_630,In_1771,In_911);
nand U631 (N_631,In_775,In_175);
xnor U632 (N_632,In_1043,In_415);
and U633 (N_633,In_1348,In_144);
or U634 (N_634,In_722,In_657);
xor U635 (N_635,In_954,In_1075);
nand U636 (N_636,In_61,In_288);
or U637 (N_637,In_667,In_1034);
nand U638 (N_638,In_1760,In_916);
xor U639 (N_639,In_1168,In_457);
xnor U640 (N_640,In_1777,In_1580);
nand U641 (N_641,In_1689,In_682);
and U642 (N_642,In_890,In_1962);
and U643 (N_643,In_1800,In_664);
nor U644 (N_644,In_1650,In_757);
nand U645 (N_645,In_1702,In_1088);
and U646 (N_646,In_188,In_678);
or U647 (N_647,In_1117,In_622);
and U648 (N_648,In_242,In_661);
and U649 (N_649,In_1714,In_645);
nand U650 (N_650,In_1282,In_1902);
nor U651 (N_651,In_103,In_1426);
and U652 (N_652,In_1812,In_1230);
nor U653 (N_653,In_607,In_1321);
or U654 (N_654,In_2,In_1773);
and U655 (N_655,In_1824,In_1862);
xnor U656 (N_656,In_145,In_97);
nor U657 (N_657,In_1977,In_924);
xor U658 (N_658,In_1327,In_1221);
nor U659 (N_659,In_810,In_1846);
and U660 (N_660,In_1662,In_782);
or U661 (N_661,In_1309,In_205);
nand U662 (N_662,In_1910,In_1169);
nor U663 (N_663,In_1219,In_1177);
nor U664 (N_664,In_284,In_576);
or U665 (N_665,In_969,In_83);
nor U666 (N_666,In_336,In_1952);
nand U667 (N_667,In_1886,In_1995);
or U668 (N_668,In_965,In_569);
xnor U669 (N_669,In_1049,In_913);
and U670 (N_670,In_65,In_1180);
xor U671 (N_671,In_129,In_187);
and U672 (N_672,In_596,In_945);
or U673 (N_673,In_1570,In_1704);
xor U674 (N_674,In_958,In_1903);
nand U675 (N_675,In_648,In_1091);
nand U676 (N_676,In_106,In_49);
xor U677 (N_677,In_1161,In_278);
or U678 (N_678,In_522,In_1319);
nor U679 (N_679,In_151,In_538);
nor U680 (N_680,In_1478,In_167);
and U681 (N_681,In_1199,In_1767);
nor U682 (N_682,In_680,In_182);
xnor U683 (N_683,In_321,In_978);
and U684 (N_684,In_305,In_1442);
and U685 (N_685,In_1984,In_1052);
and U686 (N_686,In_1443,In_1021);
and U687 (N_687,In_985,In_1303);
nand U688 (N_688,In_1241,In_1298);
or U689 (N_689,In_691,In_1833);
nand U690 (N_690,In_1949,In_1697);
nand U691 (N_691,In_204,In_1639);
nor U692 (N_692,In_1106,In_783);
xnor U693 (N_693,In_117,In_354);
and U694 (N_694,In_746,In_322);
or U695 (N_695,In_1609,In_808);
nand U696 (N_696,In_564,In_1067);
nor U697 (N_697,In_1942,In_1128);
nor U698 (N_698,In_465,In_333);
and U699 (N_699,In_1324,In_1911);
and U700 (N_700,In_90,In_1979);
and U701 (N_701,In_261,In_1647);
xor U702 (N_702,In_843,In_1022);
or U703 (N_703,In_1925,In_203);
and U704 (N_704,In_1328,In_265);
and U705 (N_705,In_561,In_172);
nand U706 (N_706,In_885,In_1679);
nor U707 (N_707,In_1093,In_626);
xnor U708 (N_708,In_619,In_1492);
nand U709 (N_709,In_1407,In_1452);
nand U710 (N_710,In_1273,In_399);
nor U711 (N_711,In_88,In_47);
and U712 (N_712,In_488,In_593);
and U713 (N_713,In_778,In_1406);
nor U714 (N_714,In_548,In_1397);
nor U715 (N_715,In_1369,In_1430);
xor U716 (N_716,In_264,In_260);
or U717 (N_717,In_126,In_1429);
and U718 (N_718,In_665,In_1173);
and U719 (N_719,In_1877,In_417);
and U720 (N_720,In_1640,In_1710);
nor U721 (N_721,In_1971,In_82);
xnor U722 (N_722,In_1975,In_595);
nand U723 (N_723,In_89,In_1053);
xnor U724 (N_724,In_1018,In_1360);
and U725 (N_725,In_346,In_390);
xnor U726 (N_726,In_712,In_1378);
nand U727 (N_727,In_1379,In_519);
nand U728 (N_728,In_196,In_1945);
xor U729 (N_729,In_578,In_1750);
nand U730 (N_730,In_1475,In_35);
xor U731 (N_731,In_1364,In_779);
and U732 (N_732,In_905,In_408);
or U733 (N_733,In_990,In_1064);
or U734 (N_734,In_1590,In_247);
and U735 (N_735,In_1226,In_473);
nand U736 (N_736,In_1353,In_1505);
and U737 (N_737,In_1285,In_527);
and U738 (N_738,In_512,In_1865);
xor U739 (N_739,In_1578,In_324);
xor U740 (N_740,In_882,In_66);
or U741 (N_741,In_1913,In_1145);
or U742 (N_742,In_1729,In_1370);
or U743 (N_743,In_267,In_1991);
xnor U744 (N_744,In_306,In_1968);
nor U745 (N_745,In_753,In_1955);
or U746 (N_746,In_403,In_353);
xnor U747 (N_747,In_900,In_442);
xnor U748 (N_748,In_350,In_1867);
and U749 (N_749,In_71,In_98);
nor U750 (N_750,In_1283,In_1588);
and U751 (N_751,In_128,In_1663);
nor U752 (N_752,In_960,In_759);
xnor U753 (N_753,In_285,In_773);
nor U754 (N_754,In_1759,In_181);
xnor U755 (N_755,In_212,In_631);
and U756 (N_756,In_115,In_1038);
nor U757 (N_757,In_313,In_1356);
nor U758 (N_758,In_949,In_1042);
or U759 (N_759,In_360,In_1296);
nor U760 (N_760,In_1003,In_20);
and U761 (N_761,In_1110,In_907);
nor U762 (N_762,In_1559,In_1891);
nor U763 (N_763,In_1488,In_428);
or U764 (N_764,In_1458,In_1146);
nor U765 (N_765,In_1349,In_612);
or U766 (N_766,In_632,In_1238);
nor U767 (N_767,In_1604,In_1811);
nand U768 (N_768,In_956,In_1908);
xnor U769 (N_769,In_910,In_1692);
or U770 (N_770,In_171,In_367);
nor U771 (N_771,In_617,In_1762);
nand U772 (N_772,In_1433,In_45);
nand U773 (N_773,In_446,In_1394);
or U774 (N_774,In_163,In_1413);
and U775 (N_775,In_1711,In_1694);
nor U776 (N_776,In_1806,In_1200);
nor U777 (N_777,In_250,In_1247);
nor U778 (N_778,In_640,In_1637);
or U779 (N_779,In_557,In_1344);
xor U780 (N_780,In_1108,In_827);
or U781 (N_781,In_809,In_1287);
nand U782 (N_782,In_795,In_1721);
nand U783 (N_783,In_392,In_197);
nand U784 (N_784,In_1896,In_1);
xnor U785 (N_785,In_871,In_1512);
or U786 (N_786,In_1858,In_78);
nor U787 (N_787,In_1726,In_1847);
or U788 (N_788,In_13,In_123);
and U789 (N_789,In_1558,In_1151);
nor U790 (N_790,In_387,In_1354);
and U791 (N_791,In_1716,In_520);
nor U792 (N_792,In_1192,In_1791);
nor U793 (N_793,In_1658,In_542);
xnor U794 (N_794,In_822,In_935);
nand U795 (N_795,In_334,In_402);
or U796 (N_796,In_994,In_1123);
and U797 (N_797,In_1752,In_1466);
and U798 (N_798,In_1242,In_1266);
xor U799 (N_799,In_406,In_1635);
xnor U800 (N_800,In_1361,N_157);
or U801 (N_801,N_503,N_321);
nand U802 (N_802,N_129,N_758);
xnor U803 (N_803,In_681,In_726);
or U804 (N_804,N_92,N_381);
nand U805 (N_805,N_665,N_423);
and U806 (N_806,In_420,N_782);
and U807 (N_807,N_340,N_633);
or U808 (N_808,In_677,In_170);
and U809 (N_809,N_374,In_1515);
or U810 (N_810,N_577,N_424);
or U811 (N_811,N_163,In_437);
nand U812 (N_812,N_465,N_105);
xor U813 (N_813,N_48,N_375);
and U814 (N_814,N_567,N_448);
nand U815 (N_815,N_371,N_662);
nand U816 (N_816,N_263,N_692);
nor U817 (N_817,N_439,In_1082);
and U818 (N_818,N_139,N_628);
nand U819 (N_819,N_500,N_365);
nand U820 (N_820,In_1398,N_142);
xnor U821 (N_821,N_42,In_39);
or U822 (N_822,N_660,N_774);
nor U823 (N_823,N_15,In_874);
or U824 (N_824,N_416,In_1405);
xnor U825 (N_825,N_85,N_21);
and U826 (N_826,In_195,In_1070);
nand U827 (N_827,N_703,N_579);
or U828 (N_828,N_286,In_364);
xor U829 (N_829,N_71,N_655);
and U830 (N_830,In_318,N_175);
xnor U831 (N_831,N_214,N_311);
and U832 (N_832,In_48,In_470);
xnor U833 (N_833,N_495,In_1930);
xnor U834 (N_834,In_1926,N_553);
xnor U835 (N_835,In_684,In_1842);
nor U836 (N_836,N_138,In_1669);
and U837 (N_837,N_132,In_858);
xor U838 (N_838,N_741,N_41);
xnor U839 (N_839,In_799,N_191);
nand U840 (N_840,N_686,N_319);
and U841 (N_841,N_56,N_638);
nor U842 (N_842,N_629,In_1094);
nor U843 (N_843,In_1062,N_775);
xor U844 (N_844,N_17,In_599);
xor U845 (N_845,N_685,In_873);
nand U846 (N_846,In_1754,In_901);
and U847 (N_847,N_677,N_199);
nand U848 (N_848,In_1509,N_196);
xnor U849 (N_849,In_307,N_390);
and U850 (N_850,N_277,In_584);
and U851 (N_851,N_536,N_480);
nor U852 (N_852,N_338,N_152);
nand U853 (N_853,N_46,N_149);
nor U854 (N_854,In_1720,N_168);
nand U855 (N_855,N_258,In_1124);
and U856 (N_856,N_678,In_184);
nand U857 (N_857,In_833,N_278);
or U858 (N_858,N_507,In_1304);
or U859 (N_859,N_642,In_513);
nand U860 (N_860,N_476,In_1994);
nor U861 (N_861,N_187,N_491);
and U862 (N_862,In_1218,In_86);
nand U863 (N_863,N_569,In_1254);
nand U864 (N_864,In_600,In_676);
or U865 (N_865,N_380,In_1878);
and U866 (N_866,In_1092,N_1);
nor U867 (N_867,N_275,N_88);
nand U868 (N_868,In_1187,N_329);
xor U869 (N_869,N_438,N_674);
and U870 (N_870,N_298,In_674);
and U871 (N_871,N_490,N_563);
or U872 (N_872,N_304,N_538);
nor U873 (N_873,N_370,N_493);
and U874 (N_874,N_483,N_724);
and U875 (N_875,N_458,N_444);
and U876 (N_876,In_423,N_714);
nor U877 (N_877,N_583,N_641);
and U878 (N_878,In_100,In_107);
and U879 (N_879,N_45,N_442);
nor U880 (N_880,In_484,In_1887);
and U881 (N_881,N_206,In_432);
or U882 (N_882,N_357,N_723);
or U883 (N_883,N_292,N_82);
and U884 (N_884,In_303,N_449);
nand U885 (N_885,In_1010,In_532);
nor U886 (N_886,N_300,N_302);
xor U887 (N_887,N_26,N_450);
xor U888 (N_888,N_100,N_167);
nor U889 (N_889,N_61,N_443);
or U890 (N_890,N_344,N_757);
xnor U891 (N_891,N_466,In_1651);
nor U892 (N_892,N_565,N_713);
and U893 (N_893,N_515,N_314);
or U894 (N_894,N_350,N_705);
or U895 (N_895,In_152,In_878);
and U896 (N_896,N_188,N_634);
and U897 (N_897,N_462,N_143);
xor U898 (N_898,N_798,N_429);
nor U899 (N_899,N_578,In_1103);
nand U900 (N_900,N_24,N_243);
and U901 (N_901,In_1325,N_355);
nor U902 (N_902,In_1996,N_180);
nor U903 (N_903,In_797,N_236);
or U904 (N_904,N_607,In_448);
and U905 (N_905,N_254,N_654);
nor U906 (N_906,N_64,N_178);
or U907 (N_907,N_29,N_60);
nand U908 (N_908,N_760,N_763);
or U909 (N_909,N_352,In_686);
nor U910 (N_910,In_926,N_54);
or U911 (N_911,N_575,N_737);
nor U912 (N_912,N_229,In_516);
xor U913 (N_913,In_1970,In_363);
xnor U914 (N_914,N_485,N_524);
or U915 (N_915,N_245,N_4);
xnor U916 (N_916,In_860,N_91);
nor U917 (N_917,N_605,In_1080);
and U918 (N_918,N_222,N_151);
or U919 (N_919,N_389,N_769);
nand U920 (N_920,N_637,In_338);
and U921 (N_921,N_299,N_532);
nor U922 (N_922,In_1892,N_512);
xor U923 (N_923,N_791,In_1245);
and U924 (N_924,N_727,N_430);
or U925 (N_925,N_657,N_471);
and U926 (N_926,N_744,N_6);
and U927 (N_927,N_122,N_447);
xor U928 (N_928,N_467,N_559);
nor U929 (N_929,N_732,In_1432);
nor U930 (N_930,N_750,N_514);
nor U931 (N_931,N_145,N_494);
xnor U932 (N_932,N_320,In_581);
and U933 (N_933,In_38,N_382);
nor U934 (N_934,In_1776,N_764);
nand U935 (N_935,N_508,In_1472);
nor U936 (N_936,In_1627,N_534);
xor U937 (N_937,N_602,N_110);
and U938 (N_938,In_95,In_1905);
or U939 (N_939,N_581,In_702);
xor U940 (N_940,N_79,N_341);
xor U941 (N_941,N_210,N_377);
nand U942 (N_942,N_257,N_646);
nor U943 (N_943,N_411,In_55);
nand U944 (N_944,In_1069,In_180);
nand U945 (N_945,N_781,In_1132);
xor U946 (N_946,N_250,In_1340);
and U947 (N_947,In_539,In_590);
and U948 (N_948,N_604,In_1932);
or U949 (N_949,N_373,N_67);
nor U950 (N_950,In_1557,N_83);
and U951 (N_951,N_36,N_787);
nor U952 (N_952,N_197,N_256);
and U953 (N_953,N_274,N_618);
nand U954 (N_954,N_179,N_74);
and U955 (N_955,N_378,N_486);
xor U956 (N_956,N_0,In_768);
or U957 (N_957,In_424,N_401);
and U958 (N_958,In_1167,In_1125);
nor U959 (N_959,N_13,N_386);
and U960 (N_960,N_496,In_1346);
or U961 (N_961,In_1376,N_5);
and U962 (N_962,N_742,N_574);
xor U963 (N_963,N_738,N_648);
nand U964 (N_964,N_632,In_1122);
xnor U965 (N_965,N_599,N_606);
or U966 (N_966,N_409,N_325);
nor U967 (N_967,N_523,N_455);
or U968 (N_968,In_839,In_1838);
and U969 (N_969,N_47,N_270);
or U970 (N_970,N_339,In_731);
nor U971 (N_971,N_399,N_269);
or U972 (N_972,N_192,N_630);
nor U973 (N_973,N_533,N_473);
and U974 (N_974,In_977,N_747);
nor U975 (N_975,N_531,N_676);
nand U976 (N_976,N_394,N_363);
or U977 (N_977,N_582,N_573);
xnor U978 (N_978,N_722,In_317);
xor U979 (N_979,N_227,In_1898);
or U980 (N_980,N_474,N_130);
nor U981 (N_981,N_470,N_543);
nor U982 (N_982,In_440,N_52);
nor U983 (N_983,N_498,N_420);
xnor U984 (N_984,N_115,N_786);
nand U985 (N_985,In_441,N_680);
nor U986 (N_986,N_649,In_27);
nand U987 (N_987,N_309,N_253);
xnor U988 (N_988,N_104,In_689);
xnor U989 (N_989,In_1428,N_631);
or U990 (N_990,N_545,In_1660);
or U991 (N_991,N_405,N_619);
xor U992 (N_992,In_1212,N_322);
xnor U993 (N_993,In_1528,N_224);
nor U994 (N_994,N_87,In_1055);
or U995 (N_995,In_1703,N_108);
or U996 (N_996,In_540,N_398);
nand U997 (N_997,N_376,N_489);
nand U998 (N_998,N_735,In_1763);
and U999 (N_999,N_10,N_711);
or U1000 (N_1000,N_177,N_431);
nor U1001 (N_1001,N_65,N_580);
and U1002 (N_1002,In_380,N_281);
and U1003 (N_1003,N_667,N_343);
and U1004 (N_1004,N_356,In_854);
and U1005 (N_1005,N_318,N_217);
nor U1006 (N_1006,N_133,N_402);
or U1007 (N_1007,N_772,N_159);
nor U1008 (N_1008,N_162,N_223);
and U1009 (N_1009,N_689,N_481);
nor U1010 (N_1010,N_57,N_622);
nor U1011 (N_1011,In_482,In_756);
and U1012 (N_1012,In_1611,In_1758);
xor U1013 (N_1013,N_384,N_135);
nand U1014 (N_1014,In_535,N_564);
or U1015 (N_1015,In_857,In_37);
nand U1016 (N_1016,In_1796,N_427);
or U1017 (N_1017,N_457,N_521);
nand U1018 (N_1018,N_392,N_174);
nor U1019 (N_1019,In_1011,N_661);
nor U1020 (N_1020,N_793,In_1850);
nand U1021 (N_1021,In_1387,N_762);
xor U1022 (N_1022,N_164,N_591);
or U1023 (N_1023,N_90,In_349);
nor U1024 (N_1024,In_1733,In_1547);
nand U1025 (N_1025,N_20,In_280);
and U1026 (N_1026,In_1438,N_460);
and U1027 (N_1027,N_600,In_119);
and U1028 (N_1028,In_1017,N_610);
and U1029 (N_1029,N_235,In_298);
or U1030 (N_1030,In_316,N_93);
nand U1031 (N_1031,In_835,N_432);
nand U1032 (N_1032,N_330,N_522);
xnor U1033 (N_1033,N_289,N_789);
and U1034 (N_1034,N_25,N_700);
nand U1035 (N_1035,In_481,N_413);
and U1036 (N_1036,N_440,N_726);
and U1037 (N_1037,N_644,N_621);
or U1038 (N_1038,N_454,N_748);
nand U1039 (N_1039,N_123,N_702);
and U1040 (N_1040,N_97,In_922);
and U1041 (N_1041,In_1054,In_841);
or U1042 (N_1042,N_589,N_294);
xnor U1043 (N_1043,N_464,N_659);
or U1044 (N_1044,In_1993,N_172);
or U1045 (N_1045,In_241,In_800);
or U1046 (N_1046,In_1237,N_316);
xnor U1047 (N_1047,In_1116,In_1444);
xnor U1048 (N_1048,N_617,N_8);
nand U1049 (N_1049,In_1560,In_1904);
xnor U1050 (N_1050,N_557,In_29);
and U1051 (N_1051,In_932,N_699);
or U1052 (N_1052,In_813,N_81);
or U1053 (N_1053,N_623,In_844);
nand U1054 (N_1054,N_240,In_1705);
nand U1055 (N_1055,In_263,N_673);
nor U1056 (N_1056,N_34,N_283);
xor U1057 (N_1057,In_829,In_1312);
xor U1058 (N_1058,In_1536,N_280);
nor U1059 (N_1059,N_183,N_771);
nand U1060 (N_1060,N_9,N_767);
and U1061 (N_1061,In_1683,In_210);
nor U1062 (N_1062,N_73,N_75);
nor U1063 (N_1063,N_154,N_799);
nand U1064 (N_1064,N_753,N_354);
and U1065 (N_1065,N_379,N_367);
and U1066 (N_1066,In_812,In_577);
nand U1067 (N_1067,N_117,In_194);
or U1068 (N_1068,N_160,In_1441);
and U1069 (N_1069,N_120,N_182);
or U1070 (N_1070,In_1856,N_221);
nor U1071 (N_1071,N_246,N_19);
nand U1072 (N_1072,N_368,N_241);
nor U1073 (N_1073,N_746,N_282);
or U1074 (N_1074,N_548,N_488);
nor U1075 (N_1075,N_584,N_248);
xnor U1076 (N_1076,N_710,N_66);
or U1077 (N_1077,N_118,In_1849);
or U1078 (N_1078,N_358,N_194);
nand U1079 (N_1079,N_234,N_276);
nor U1080 (N_1080,N_482,In_302);
xnor U1081 (N_1081,N_131,N_406);
xor U1082 (N_1082,N_198,N_50);
or U1083 (N_1083,N_561,N_756);
or U1084 (N_1084,N_336,In_1533);
nor U1085 (N_1085,N_730,N_396);
nor U1086 (N_1086,N_716,In_43);
xnor U1087 (N_1087,In_1439,N_2);
nor U1088 (N_1088,In_587,N_696);
xor U1089 (N_1089,N_211,N_252);
xnor U1090 (N_1090,N_576,N_111);
xnor U1091 (N_1091,N_520,N_525);
nand U1092 (N_1092,N_261,In_1491);
xnor U1093 (N_1093,N_249,N_230);
nand U1094 (N_1094,N_588,N_428);
nand U1095 (N_1095,In_1090,N_213);
nand U1096 (N_1096,N_539,In_1827);
or U1097 (N_1097,In_1672,N_647);
xnor U1098 (N_1098,In_792,N_63);
nor U1099 (N_1099,In_1140,N_364);
or U1100 (N_1100,In_297,N_668);
nor U1101 (N_1101,N_671,In_42);
or U1102 (N_1102,N_301,N_134);
xnor U1103 (N_1103,N_158,N_719);
nor U1104 (N_1104,N_445,N_614);
or U1105 (N_1105,N_89,In_1014);
or U1106 (N_1106,In_1507,N_451);
nand U1107 (N_1107,N_505,N_785);
and U1108 (N_1108,N_310,N_656);
nand U1109 (N_1109,N_267,N_366);
nor U1110 (N_1110,N_652,N_101);
and U1111 (N_1111,In_1463,In_531);
nand U1112 (N_1112,N_627,In_1615);
xnor U1113 (N_1113,In_1333,N_94);
and U1114 (N_1114,In_1899,In_1214);
nand U1115 (N_1115,In_1477,N_541);
and U1116 (N_1116,In_987,In_630);
nand U1117 (N_1117,In_983,N_720);
nand U1118 (N_1118,N_777,N_492);
xor U1119 (N_1119,N_415,N_369);
and U1120 (N_1120,In_1897,In_1657);
nand U1121 (N_1121,N_783,N_190);
or U1122 (N_1122,N_506,N_780);
nand U1123 (N_1123,N_640,In_1837);
or U1124 (N_1124,N_40,N_663);
nand U1125 (N_1125,N_239,In_1341);
nand U1126 (N_1126,N_529,N_27);
xnor U1127 (N_1127,In_486,N_408);
or U1128 (N_1128,In_1548,N_126);
xnor U1129 (N_1129,N_562,In_982);
and U1130 (N_1130,N_106,N_620);
nor U1131 (N_1131,N_698,N_147);
nand U1132 (N_1132,N_736,N_315);
or U1133 (N_1133,In_1918,N_593);
nor U1134 (N_1134,N_436,N_546);
nor U1135 (N_1135,In_912,In_1274);
nor U1136 (N_1136,In_824,N_16);
nand U1137 (N_1137,N_80,In_1981);
nand U1138 (N_1138,N_479,In_9);
and U1139 (N_1139,N_414,N_12);
nand U1140 (N_1140,In_1059,N_247);
or U1141 (N_1141,N_765,N_306);
or U1142 (N_1142,In_1649,N_537);
nand U1143 (N_1143,In_275,In_504);
or U1144 (N_1144,In_1860,In_1272);
nand U1145 (N_1145,In_262,In_864);
nand U1146 (N_1146,N_30,In_1868);
nor U1147 (N_1147,N_570,In_217);
xor U1148 (N_1148,N_346,N_124);
or U1149 (N_1149,N_422,N_287);
or U1150 (N_1150,N_285,In_991);
and U1151 (N_1151,N_317,N_547);
nor U1152 (N_1152,N_342,N_77);
nand U1153 (N_1153,In_1068,In_161);
or U1154 (N_1154,N_335,N_226);
nor U1155 (N_1155,N_201,In_109);
and U1156 (N_1156,In_327,In_1163);
or U1157 (N_1157,N_136,N_70);
and U1158 (N_1158,N_76,In_1085);
or U1159 (N_1159,In_769,In_1362);
nor U1160 (N_1160,N_518,In_1178);
nor U1161 (N_1161,N_153,In_1384);
nand U1162 (N_1162,N_612,In_1299);
or U1163 (N_1163,In_1032,In_897);
nand U1164 (N_1164,N_3,N_259);
and U1165 (N_1165,N_527,N_717);
or U1166 (N_1166,N_468,N_33);
nand U1167 (N_1167,N_776,N_189);
and U1168 (N_1168,N_790,N_170);
and U1169 (N_1169,In_429,N_397);
nor U1170 (N_1170,N_425,N_708);
xnor U1171 (N_1171,In_541,In_534);
xor U1172 (N_1172,N_690,N_102);
xnor U1173 (N_1173,N_770,N_144);
nor U1174 (N_1174,N_146,N_303);
nor U1175 (N_1175,N_308,N_43);
xnor U1176 (N_1176,N_596,N_32);
nor U1177 (N_1177,In_51,N_232);
or U1178 (N_1178,In_1737,N_497);
xnor U1179 (N_1179,N_238,N_434);
and U1180 (N_1180,N_516,In_1486);
xnor U1181 (N_1181,N_361,In_155);
or U1182 (N_1182,In_26,N_193);
xor U1183 (N_1183,N_729,In_1629);
nor U1184 (N_1184,N_658,N_773);
nand U1185 (N_1185,N_566,N_233);
or U1186 (N_1186,In_927,N_613);
nand U1187 (N_1187,N_171,In_1308);
or U1188 (N_1188,In_766,In_1331);
nand U1189 (N_1189,In_1048,In_233);
and U1190 (N_1190,N_345,N_412);
nand U1191 (N_1191,In_1246,N_51);
nand U1192 (N_1192,N_597,N_718);
xor U1193 (N_1193,N_62,N_395);
or U1194 (N_1194,N_264,N_526);
or U1195 (N_1195,In_216,In_1041);
nor U1196 (N_1196,N_296,In_802);
and U1197 (N_1197,In_715,In_449);
nand U1198 (N_1198,In_1954,N_752);
xnor U1199 (N_1199,N_437,N_550);
xnor U1200 (N_1200,In_700,In_1503);
nor U1201 (N_1201,N_733,N_218);
nor U1202 (N_1202,N_446,In_748);
xnor U1203 (N_1203,In_998,N_441);
xor U1204 (N_1204,N_555,N_195);
nand U1205 (N_1205,N_544,In_253);
and U1206 (N_1206,In_1099,In_1350);
nor U1207 (N_1207,N_461,N_400);
xor U1208 (N_1208,N_166,N_348);
nor U1209 (N_1209,In_995,N_421);
and U1210 (N_1210,N_517,In_1620);
and U1211 (N_1211,In_1648,In_952);
or U1212 (N_1212,In_1668,N_39);
or U1213 (N_1213,N_484,In_1460);
and U1214 (N_1214,N_208,N_552);
nand U1215 (N_1215,N_291,N_324);
xnor U1216 (N_1216,N_704,N_202);
and U1217 (N_1217,In_199,N_215);
or U1218 (N_1218,N_797,In_832);
xnor U1219 (N_1219,N_307,N_609);
nor U1220 (N_1220,N_501,In_1864);
nand U1221 (N_1221,N_44,N_639);
or U1222 (N_1222,N_69,In_980);
and U1223 (N_1223,N_694,N_636);
nand U1224 (N_1224,N_140,In_478);
nor U1225 (N_1225,In_1768,In_1194);
xor U1226 (N_1226,N_419,N_107);
nand U1227 (N_1227,In_787,N_707);
nand U1228 (N_1228,In_1007,N_616);
xor U1229 (N_1229,N_86,In_1028);
nand U1230 (N_1230,In_1795,N_103);
and U1231 (N_1231,In_846,N_58);
xnor U1232 (N_1232,In_1775,In_323);
nand U1233 (N_1233,In_1688,N_433);
xor U1234 (N_1234,In_1256,In_891);
or U1235 (N_1235,N_615,N_558);
nand U1236 (N_1236,N_768,N_99);
nand U1237 (N_1237,In_1015,N_734);
nand U1238 (N_1238,N_653,N_255);
xnor U1239 (N_1239,N_754,N_387);
and U1240 (N_1240,N_568,N_205);
nor U1241 (N_1241,N_796,In_70);
and U1242 (N_1242,N_551,N_209);
nand U1243 (N_1243,N_792,In_1368);
xor U1244 (N_1244,N_200,In_294);
xnor U1245 (N_1245,N_595,In_1946);
nand U1246 (N_1246,N_161,N_7);
nand U1247 (N_1247,N_666,N_332);
or U1248 (N_1248,N_18,N_313);
nand U1249 (N_1249,N_554,N_403);
or U1250 (N_1250,In_692,N_169);
or U1251 (N_1251,N_351,N_284);
and U1252 (N_1252,N_794,In_249);
or U1253 (N_1253,N_333,In_725);
nor U1254 (N_1254,N_670,N_410);
and U1255 (N_1255,N_116,In_947);
or U1256 (N_1256,N_435,In_80);
and U1257 (N_1257,In_780,In_1828);
nor U1258 (N_1258,N_68,N_643);
xor U1259 (N_1259,In_1934,N_509);
or U1260 (N_1260,N_383,N_586);
or U1261 (N_1261,N_745,N_35);
or U1262 (N_1262,N_31,N_472);
xnor U1263 (N_1263,N_778,In_732);
nor U1264 (N_1264,N_137,In_1974);
nand U1265 (N_1265,N_549,N_279);
nand U1266 (N_1266,N_688,In_1517);
nor U1267 (N_1267,N_560,N_795);
nand U1268 (N_1268,N_404,N_216);
nand U1269 (N_1269,N_113,In_591);
nor U1270 (N_1270,In_848,N_603);
nor U1271 (N_1271,N_262,N_556);
xnor U1272 (N_1272,N_141,N_72);
xnor U1273 (N_1273,In_1538,N_186);
nand U1274 (N_1274,N_295,In_555);
xor U1275 (N_1275,In_836,N_212);
nor U1276 (N_1276,N_456,N_585);
xnor U1277 (N_1277,N_684,In_508);
xor U1278 (N_1278,N_38,In_1622);
or U1279 (N_1279,N_360,N_426);
nand U1280 (N_1280,N_594,N_272);
nand U1281 (N_1281,N_542,In_1050);
nor U1282 (N_1282,N_535,N_96);
and U1283 (N_1283,In_1922,In_817);
xnor U1284 (N_1284,In_40,N_78);
and U1285 (N_1285,In_131,N_260);
or U1286 (N_1286,In_1135,In_102);
nand U1287 (N_1287,N_695,In_727);
or U1288 (N_1288,N_788,N_127);
or U1289 (N_1289,In_1881,In_842);
and U1290 (N_1290,In_716,In_1162);
nor U1291 (N_1291,In_507,N_682);
and U1292 (N_1292,N_150,In_984);
or U1293 (N_1293,In_1025,In_434);
nand U1294 (N_1294,N_697,N_293);
and U1295 (N_1295,In_574,N_779);
xnor U1296 (N_1296,In_1638,N_693);
xnor U1297 (N_1297,N_511,In_610);
nor U1298 (N_1298,N_290,In_1009);
or U1299 (N_1299,N_478,In_711);
or U1300 (N_1300,N_650,In_1836);
and U1301 (N_1301,N_587,In_1780);
nor U1302 (N_1302,In_1805,In_1666);
nor U1303 (N_1303,N_125,N_181);
xor U1304 (N_1304,N_337,In_1531);
and U1305 (N_1305,In_219,In_853);
and U1306 (N_1306,In_1314,In_1690);
nor U1307 (N_1307,In_1855,N_721);
nand U1308 (N_1308,N_11,N_266);
xor U1309 (N_1309,In_1166,N_55);
and U1310 (N_1310,N_477,N_237);
nor U1311 (N_1311,In_1781,In_458);
xor U1312 (N_1312,N_592,N_119);
and U1313 (N_1313,N_362,In_946);
and U1314 (N_1314,N_23,N_469);
xnor U1315 (N_1315,N_203,In_1375);
nand U1316 (N_1316,N_759,In_1381);
nand U1317 (N_1317,In_785,N_625);
xnor U1318 (N_1318,In_1591,N_49);
nor U1319 (N_1319,N_530,N_326);
and U1320 (N_1320,N_459,In_173);
and U1321 (N_1321,N_590,N_645);
nand U1322 (N_1322,N_372,N_155);
xnor U1323 (N_1323,In_1408,In_1815);
nor U1324 (N_1324,N_624,N_385);
nand U1325 (N_1325,N_701,N_519);
nand U1326 (N_1326,N_418,In_707);
nor U1327 (N_1327,N_571,N_359);
or U1328 (N_1328,N_740,In_1939);
and U1329 (N_1329,N_706,N_453);
xnor U1330 (N_1330,In_1755,N_626);
xor U1331 (N_1331,N_761,N_651);
nand U1332 (N_1332,N_743,N_265);
nor U1333 (N_1333,N_323,N_725);
nor U1334 (N_1334,N_393,N_204);
nand U1335 (N_1335,In_1338,N_251);
or U1336 (N_1336,In_818,N_672);
xor U1337 (N_1337,N_513,N_452);
and U1338 (N_1338,N_784,In_174);
and U1339 (N_1339,N_14,In_1323);
nand U1340 (N_1340,In_1593,In_251);
or U1341 (N_1341,N_739,N_173);
or U1342 (N_1342,In_379,N_683);
nor U1343 (N_1343,N_608,N_305);
nor U1344 (N_1344,N_185,N_327);
or U1345 (N_1345,N_679,N_499);
nand U1346 (N_1346,N_601,N_219);
or U1347 (N_1347,N_504,In_1208);
and U1348 (N_1348,In_1270,N_675);
xor U1349 (N_1349,In_81,N_28);
nor U1350 (N_1350,In_176,N_687);
nand U1351 (N_1351,In_1687,In_1744);
nor U1352 (N_1352,N_475,N_664);
nor U1353 (N_1353,N_510,N_334);
xnor U1354 (N_1354,N_407,N_244);
or U1355 (N_1355,N_487,N_328);
and U1356 (N_1356,N_347,In_1645);
nor U1357 (N_1357,In_974,N_691);
nor U1358 (N_1358,N_388,N_95);
nor U1359 (N_1359,N_528,N_755);
nand U1360 (N_1360,N_165,In_1182);
or U1361 (N_1361,N_220,N_98);
or U1362 (N_1362,N_59,In_642);
or U1363 (N_1363,N_312,N_611);
nand U1364 (N_1364,In_142,N_598);
and U1365 (N_1365,N_572,N_121);
or U1366 (N_1366,N_176,N_681);
or U1367 (N_1367,In_740,In_1185);
xor U1368 (N_1368,In_762,In_589);
nand U1369 (N_1369,In_823,N_288);
nand U1370 (N_1370,N_148,N_349);
nor U1371 (N_1371,In_1326,N_273);
nand U1372 (N_1372,N_112,In_1290);
or U1373 (N_1373,N_242,N_84);
nand U1374 (N_1374,In_1709,In_378);
nor U1375 (N_1375,N_712,In_514);
and U1376 (N_1376,N_728,In_502);
nor U1377 (N_1377,N_156,N_540);
xor U1378 (N_1378,In_855,N_766);
xor U1379 (N_1379,In_1584,In_84);
nand U1380 (N_1380,N_502,N_207);
nand U1381 (N_1381,N_731,In_1739);
nand U1382 (N_1382,N_22,N_391);
nand U1383 (N_1383,In_1249,N_709);
nor U1384 (N_1384,N_37,N_271);
nor U1385 (N_1385,N_184,N_463);
nor U1386 (N_1386,N_268,In_1612);
xor U1387 (N_1387,In_1301,N_715);
and U1388 (N_1388,N_128,N_114);
xor U1389 (N_1389,N_225,In_671);
xnor U1390 (N_1390,N_751,In_1293);
xor U1391 (N_1391,In_1039,N_297);
and U1392 (N_1392,In_463,N_331);
nor U1393 (N_1393,N_353,In_1001);
nor U1394 (N_1394,In_1592,N_749);
nand U1395 (N_1395,N_635,N_53);
xor U1396 (N_1396,In_290,N_417);
and U1397 (N_1397,N_231,N_228);
xor U1398 (N_1398,In_1288,N_109);
and U1399 (N_1399,In_1044,N_669);
xnor U1400 (N_1400,In_1304,N_738);
or U1401 (N_1401,N_648,In_1099);
xor U1402 (N_1402,In_1612,N_673);
or U1403 (N_1403,N_188,N_311);
nand U1404 (N_1404,N_761,N_387);
or U1405 (N_1405,N_206,In_1687);
and U1406 (N_1406,N_394,N_498);
and U1407 (N_1407,N_132,In_947);
and U1408 (N_1408,N_74,N_613);
or U1409 (N_1409,N_681,N_362);
and U1410 (N_1410,N_741,N_715);
or U1411 (N_1411,In_210,N_13);
nand U1412 (N_1412,In_1350,In_974);
nand U1413 (N_1413,N_487,N_593);
nand U1414 (N_1414,In_263,N_114);
nand U1415 (N_1415,In_932,In_48);
nor U1416 (N_1416,N_564,N_793);
and U1417 (N_1417,In_715,N_249);
xor U1418 (N_1418,In_600,In_1934);
nor U1419 (N_1419,N_699,N_168);
xnor U1420 (N_1420,In_1068,N_149);
xor U1421 (N_1421,N_78,N_96);
and U1422 (N_1422,In_1405,In_1560);
xnor U1423 (N_1423,In_1612,N_157);
and U1424 (N_1424,In_37,N_178);
xor U1425 (N_1425,N_456,In_1028);
nand U1426 (N_1426,N_706,N_40);
xnor U1427 (N_1427,In_51,N_329);
xor U1428 (N_1428,N_59,N_683);
nand U1429 (N_1429,N_149,In_297);
and U1430 (N_1430,N_180,N_280);
nor U1431 (N_1431,N_47,N_715);
and U1432 (N_1432,N_680,N_82);
xor U1433 (N_1433,N_55,In_1099);
nand U1434 (N_1434,In_39,In_43);
xnor U1435 (N_1435,In_762,N_70);
nor U1436 (N_1436,N_615,N_636);
or U1437 (N_1437,N_413,N_177);
and U1438 (N_1438,In_858,N_602);
xor U1439 (N_1439,N_727,In_873);
nor U1440 (N_1440,N_773,N_163);
nand U1441 (N_1441,In_1182,N_481);
nor U1442 (N_1442,N_445,N_66);
xor U1443 (N_1443,N_44,N_517);
nor U1444 (N_1444,N_64,N_592);
nand U1445 (N_1445,N_381,N_79);
or U1446 (N_1446,N_424,In_199);
or U1447 (N_1447,N_623,In_1375);
nor U1448 (N_1448,N_422,In_842);
xor U1449 (N_1449,In_692,N_417);
nand U1450 (N_1450,N_244,N_29);
xor U1451 (N_1451,In_581,In_1135);
xor U1452 (N_1452,In_1533,In_1615);
and U1453 (N_1453,N_410,N_648);
nand U1454 (N_1454,N_367,N_476);
or U1455 (N_1455,N_51,In_1477);
or U1456 (N_1456,N_311,N_737);
nor U1457 (N_1457,N_726,In_1041);
or U1458 (N_1458,In_1080,In_1333);
xor U1459 (N_1459,In_1381,In_800);
nor U1460 (N_1460,N_40,In_1032);
xor U1461 (N_1461,N_97,In_912);
nor U1462 (N_1462,N_365,N_277);
nor U1463 (N_1463,N_382,N_189);
or U1464 (N_1464,N_233,N_532);
nor U1465 (N_1465,In_1688,In_253);
xnor U1466 (N_1466,N_489,In_262);
nor U1467 (N_1467,N_757,N_32);
nor U1468 (N_1468,N_712,N_773);
and U1469 (N_1469,N_150,N_611);
xor U1470 (N_1470,In_1050,N_793);
nand U1471 (N_1471,N_736,N_506);
nand U1472 (N_1472,N_105,N_434);
or U1473 (N_1473,N_94,N_583);
xor U1474 (N_1474,N_221,In_173);
xor U1475 (N_1475,N_62,N_593);
nand U1476 (N_1476,N_573,N_313);
nor U1477 (N_1477,N_205,In_253);
nor U1478 (N_1478,In_1849,In_180);
and U1479 (N_1479,N_763,N_265);
xor U1480 (N_1480,N_424,N_275);
and U1481 (N_1481,In_591,N_18);
nand U1482 (N_1482,In_1974,N_127);
nand U1483 (N_1483,N_661,N_426);
or U1484 (N_1484,In_1611,N_75);
and U1485 (N_1485,N_522,In_1649);
or U1486 (N_1486,In_674,In_740);
and U1487 (N_1487,N_431,In_1011);
xnor U1488 (N_1488,N_391,N_84);
and U1489 (N_1489,N_766,In_980);
nor U1490 (N_1490,N_150,N_414);
and U1491 (N_1491,In_952,In_1611);
and U1492 (N_1492,N_448,N_687);
and U1493 (N_1493,N_47,In_1044);
nand U1494 (N_1494,In_700,In_1981);
nand U1495 (N_1495,In_977,In_748);
or U1496 (N_1496,In_1299,N_371);
and U1497 (N_1497,N_360,N_251);
nand U1498 (N_1498,N_102,In_715);
or U1499 (N_1499,In_303,N_313);
or U1500 (N_1500,N_551,N_134);
and U1501 (N_1501,N_361,In_484);
and U1502 (N_1502,N_329,N_564);
nor U1503 (N_1503,N_248,In_131);
and U1504 (N_1504,N_201,In_195);
nand U1505 (N_1505,N_702,N_115);
nand U1506 (N_1506,N_89,In_349);
and U1507 (N_1507,N_89,N_186);
nand U1508 (N_1508,In_241,N_543);
and U1509 (N_1509,N_561,In_732);
xnor U1510 (N_1510,N_376,N_547);
and U1511 (N_1511,N_66,N_448);
nor U1512 (N_1512,N_116,N_241);
or U1513 (N_1513,In_1592,N_753);
xor U1514 (N_1514,N_566,N_494);
nand U1515 (N_1515,N_202,In_40);
xor U1516 (N_1516,In_380,N_62);
nor U1517 (N_1517,N_302,N_462);
nand U1518 (N_1518,N_627,N_67);
nand U1519 (N_1519,N_783,N_204);
nand U1520 (N_1520,N_293,In_513);
or U1521 (N_1521,N_287,In_984);
xnor U1522 (N_1522,N_402,N_415);
xnor U1523 (N_1523,N_428,In_787);
nor U1524 (N_1524,N_566,N_445);
xnor U1525 (N_1525,In_513,In_323);
or U1526 (N_1526,In_152,N_74);
nand U1527 (N_1527,N_21,In_841);
and U1528 (N_1528,In_531,In_1666);
xor U1529 (N_1529,N_169,N_710);
nand U1530 (N_1530,In_841,N_675);
and U1531 (N_1531,N_531,N_757);
or U1532 (N_1532,In_316,N_737);
xnor U1533 (N_1533,N_423,N_798);
xor U1534 (N_1534,N_251,N_108);
nand U1535 (N_1535,N_793,In_449);
nor U1536 (N_1536,In_102,In_1993);
xnor U1537 (N_1537,In_1341,N_625);
nand U1538 (N_1538,N_274,In_785);
and U1539 (N_1539,In_1428,N_530);
xor U1540 (N_1540,N_799,In_1208);
nand U1541 (N_1541,N_192,N_541);
or U1542 (N_1542,N_279,In_991);
or U1543 (N_1543,In_878,In_1864);
or U1544 (N_1544,N_363,N_793);
and U1545 (N_1545,N_508,N_646);
and U1546 (N_1546,In_766,N_290);
xor U1547 (N_1547,N_475,N_477);
xor U1548 (N_1548,N_686,In_478);
nand U1549 (N_1549,N_768,N_71);
and U1550 (N_1550,N_142,N_181);
nor U1551 (N_1551,N_727,In_1028);
or U1552 (N_1552,N_59,N_277);
nand U1553 (N_1553,N_295,N_611);
and U1554 (N_1554,In_1860,N_538);
xor U1555 (N_1555,In_829,N_343);
xnor U1556 (N_1556,N_700,N_602);
nor U1557 (N_1557,In_27,N_451);
and U1558 (N_1558,In_1376,In_1301);
xnor U1559 (N_1559,N_217,N_143);
and U1560 (N_1560,N_487,N_76);
xnor U1561 (N_1561,In_303,N_280);
nand U1562 (N_1562,N_780,In_1638);
nor U1563 (N_1563,N_312,In_1408);
or U1564 (N_1564,In_715,N_253);
xnor U1565 (N_1565,In_379,N_657);
or U1566 (N_1566,N_716,N_664);
xnor U1567 (N_1567,In_1828,N_390);
xnor U1568 (N_1568,N_173,In_1059);
nor U1569 (N_1569,In_253,N_365);
or U1570 (N_1570,In_176,N_79);
nor U1571 (N_1571,In_1905,N_161);
or U1572 (N_1572,N_559,In_732);
xor U1573 (N_1573,N_334,N_168);
nand U1574 (N_1574,N_340,N_224);
nor U1575 (N_1575,N_759,In_1758);
nor U1576 (N_1576,In_1054,N_312);
and U1577 (N_1577,In_1926,In_176);
and U1578 (N_1578,N_449,In_574);
and U1579 (N_1579,N_148,N_751);
xor U1580 (N_1580,In_1439,N_760);
and U1581 (N_1581,In_780,N_487);
xnor U1582 (N_1582,N_138,In_1531);
or U1583 (N_1583,N_299,N_50);
nor U1584 (N_1584,N_642,N_629);
nand U1585 (N_1585,In_1669,N_370);
nand U1586 (N_1586,N_118,N_594);
or U1587 (N_1587,N_317,N_320);
or U1588 (N_1588,N_760,N_71);
nor U1589 (N_1589,N_703,N_415);
xor U1590 (N_1590,N_102,In_470);
xnor U1591 (N_1591,In_1996,In_174);
nand U1592 (N_1592,N_656,N_541);
and U1593 (N_1593,N_103,N_739);
and U1594 (N_1594,In_824,In_1974);
or U1595 (N_1595,In_1946,N_475);
nor U1596 (N_1596,In_249,N_608);
or U1597 (N_1597,In_1162,N_774);
xnor U1598 (N_1598,N_295,In_1781);
nor U1599 (N_1599,N_683,N_761);
or U1600 (N_1600,N_812,N_1267);
or U1601 (N_1601,N_1076,N_1155);
nor U1602 (N_1602,N_1486,N_1350);
and U1603 (N_1603,N_864,N_1016);
and U1604 (N_1604,N_1571,N_1420);
xnor U1605 (N_1605,N_1331,N_1322);
nor U1606 (N_1606,N_1552,N_1159);
nand U1607 (N_1607,N_1090,N_875);
nand U1608 (N_1608,N_1590,N_1026);
xor U1609 (N_1609,N_1098,N_1270);
nand U1610 (N_1610,N_991,N_983);
nor U1611 (N_1611,N_1162,N_1091);
or U1612 (N_1612,N_1277,N_1115);
xor U1613 (N_1613,N_1490,N_960);
nor U1614 (N_1614,N_1087,N_1376);
nor U1615 (N_1615,N_866,N_907);
and U1616 (N_1616,N_1004,N_1374);
xor U1617 (N_1617,N_827,N_880);
nand U1618 (N_1618,N_1360,N_1167);
or U1619 (N_1619,N_1422,N_965);
or U1620 (N_1620,N_1089,N_1278);
nand U1621 (N_1621,N_850,N_1522);
nand U1622 (N_1622,N_1104,N_1453);
nor U1623 (N_1623,N_1592,N_952);
nand U1624 (N_1624,N_1367,N_846);
nand U1625 (N_1625,N_1263,N_1371);
and U1626 (N_1626,N_1046,N_1209);
xnor U1627 (N_1627,N_1314,N_912);
xor U1628 (N_1628,N_1538,N_914);
nor U1629 (N_1629,N_1218,N_1107);
nor U1630 (N_1630,N_1359,N_927);
and U1631 (N_1631,N_968,N_862);
and U1632 (N_1632,N_1388,N_1041);
or U1633 (N_1633,N_1212,N_1300);
nor U1634 (N_1634,N_1363,N_1495);
xnor U1635 (N_1635,N_1001,N_1430);
nor U1636 (N_1636,N_1311,N_985);
and U1637 (N_1637,N_1273,N_1321);
nor U1638 (N_1638,N_1346,N_1061);
and U1639 (N_1639,N_1465,N_1228);
nand U1640 (N_1640,N_853,N_877);
nand U1641 (N_1641,N_1492,N_1403);
xor U1642 (N_1642,N_1445,N_1187);
or U1643 (N_1643,N_919,N_1512);
nor U1644 (N_1644,N_845,N_1247);
and U1645 (N_1645,N_1597,N_1250);
nand U1646 (N_1646,N_1306,N_1148);
nor U1647 (N_1647,N_1121,N_891);
nand U1648 (N_1648,N_838,N_1096);
nand U1649 (N_1649,N_1020,N_1546);
or U1650 (N_1650,N_1160,N_1528);
xor U1651 (N_1651,N_1013,N_989);
and U1652 (N_1652,N_1578,N_1544);
xnor U1653 (N_1653,N_1223,N_1560);
nor U1654 (N_1654,N_1054,N_1058);
xnor U1655 (N_1655,N_1498,N_1535);
xnor U1656 (N_1656,N_1339,N_1274);
xnor U1657 (N_1657,N_1395,N_1040);
nor U1658 (N_1658,N_1432,N_1084);
xor U1659 (N_1659,N_1125,N_1410);
and U1660 (N_1660,N_1372,N_1165);
xor U1661 (N_1661,N_1017,N_1405);
and U1662 (N_1662,N_1200,N_1014);
xor U1663 (N_1663,N_837,N_1312);
or U1664 (N_1664,N_909,N_1503);
nand U1665 (N_1665,N_1586,N_1565);
xor U1666 (N_1666,N_964,N_1128);
or U1667 (N_1667,N_1369,N_1483);
and U1668 (N_1668,N_1100,N_994);
nand U1669 (N_1669,N_1464,N_888);
xor U1670 (N_1670,N_1358,N_1351);
and U1671 (N_1671,N_1497,N_1450);
xnor U1672 (N_1672,N_1508,N_1393);
or U1673 (N_1673,N_1563,N_1518);
or U1674 (N_1674,N_1392,N_1309);
nor U1675 (N_1675,N_955,N_982);
and U1676 (N_1676,N_1409,N_1334);
nor U1677 (N_1677,N_1295,N_1293);
nor U1678 (N_1678,N_937,N_953);
xor U1679 (N_1679,N_1303,N_958);
xor U1680 (N_1680,N_1182,N_1328);
nor U1681 (N_1681,N_1072,N_1177);
nand U1682 (N_1682,N_938,N_1166);
nor U1683 (N_1683,N_1556,N_1461);
or U1684 (N_1684,N_1336,N_993);
xor U1685 (N_1685,N_802,N_923);
nor U1686 (N_1686,N_957,N_1067);
xnor U1687 (N_1687,N_1285,N_1261);
xnor U1688 (N_1688,N_1063,N_1525);
nor U1689 (N_1689,N_1401,N_1010);
xnor U1690 (N_1690,N_1255,N_1158);
nor U1691 (N_1691,N_1554,N_1417);
xor U1692 (N_1692,N_1025,N_809);
nor U1693 (N_1693,N_1437,N_951);
xor U1694 (N_1694,N_1305,N_1480);
xor U1695 (N_1695,N_820,N_945);
and U1696 (N_1696,N_1039,N_1352);
and U1697 (N_1697,N_905,N_1326);
or U1698 (N_1698,N_1124,N_1254);
or U1699 (N_1699,N_984,N_899);
or U1700 (N_1700,N_906,N_1414);
nand U1701 (N_1701,N_1170,N_1353);
xnor U1702 (N_1702,N_1493,N_828);
xor U1703 (N_1703,N_1572,N_933);
xnor U1704 (N_1704,N_1206,N_895);
nor U1705 (N_1705,N_1226,N_1479);
and U1706 (N_1706,N_1559,N_915);
and U1707 (N_1707,N_997,N_1071);
or U1708 (N_1708,N_1361,N_829);
and U1709 (N_1709,N_1216,N_1217);
or U1710 (N_1710,N_1284,N_1438);
and U1711 (N_1711,N_1567,N_1561);
nand U1712 (N_1712,N_1418,N_1411);
nor U1713 (N_1713,N_885,N_857);
nand U1714 (N_1714,N_1362,N_813);
and U1715 (N_1715,N_939,N_1031);
or U1716 (N_1716,N_943,N_1118);
nand U1717 (N_1717,N_1564,N_1421);
or U1718 (N_1718,N_1557,N_1074);
xnor U1719 (N_1719,N_1068,N_1019);
xnor U1720 (N_1720,N_1536,N_852);
and U1721 (N_1721,N_1488,N_1034);
xor U1722 (N_1722,N_848,N_1385);
nor U1723 (N_1723,N_1221,N_807);
and U1724 (N_1724,N_1378,N_1570);
xor U1725 (N_1725,N_865,N_894);
nor U1726 (N_1726,N_1229,N_1070);
xnor U1727 (N_1727,N_1587,N_1407);
nor U1728 (N_1728,N_1269,N_918);
xor U1729 (N_1729,N_1215,N_1164);
or U1730 (N_1730,N_1175,N_1398);
and U1731 (N_1731,N_975,N_841);
nand U1732 (N_1732,N_1537,N_1122);
xnor U1733 (N_1733,N_913,N_1241);
nand U1734 (N_1734,N_1207,N_978);
nand U1735 (N_1735,N_1514,N_1198);
and U1736 (N_1736,N_1294,N_1595);
or U1737 (N_1737,N_1481,N_1332);
and U1738 (N_1738,N_931,N_1506);
nand U1739 (N_1739,N_1179,N_1341);
or U1740 (N_1740,N_815,N_969);
nand U1741 (N_1741,N_1348,N_1073);
nand U1742 (N_1742,N_1062,N_1235);
xnor U1743 (N_1743,N_1575,N_1012);
nand U1744 (N_1744,N_1455,N_1429);
xnor U1745 (N_1745,N_1545,N_1018);
and U1746 (N_1746,N_1236,N_934);
xnor U1747 (N_1747,N_1387,N_1373);
or U1748 (N_1748,N_910,N_1591);
or U1749 (N_1749,N_816,N_1349);
nor U1750 (N_1750,N_1279,N_823);
nand U1751 (N_1751,N_801,N_1153);
or U1752 (N_1752,N_1172,N_1021);
nor U1753 (N_1753,N_1583,N_908);
and U1754 (N_1754,N_962,N_1057);
xor U1755 (N_1755,N_971,N_1171);
nand U1756 (N_1756,N_879,N_1291);
xnor U1757 (N_1757,N_1059,N_1183);
and U1758 (N_1758,N_902,N_1534);
nor U1759 (N_1759,N_1547,N_1214);
xnor U1760 (N_1760,N_1402,N_1489);
or U1761 (N_1761,N_1368,N_1441);
or U1762 (N_1762,N_868,N_950);
nor U1763 (N_1763,N_1022,N_1130);
nor U1764 (N_1764,N_1242,N_1365);
and U1765 (N_1765,N_1213,N_1262);
and U1766 (N_1766,N_976,N_804);
or U1767 (N_1767,N_1327,N_1458);
nand U1768 (N_1768,N_1555,N_1467);
xor U1769 (N_1769,N_1335,N_1006);
and U1770 (N_1770,N_1095,N_884);
nand U1771 (N_1771,N_890,N_947);
nor U1772 (N_1772,N_1077,N_1008);
nor U1773 (N_1773,N_1268,N_1507);
and U1774 (N_1774,N_1195,N_1333);
xor U1775 (N_1775,N_1265,N_1501);
xnor U1776 (N_1776,N_917,N_1375);
or U1777 (N_1777,N_863,N_1007);
nand U1778 (N_1778,N_832,N_1028);
or U1779 (N_1779,N_1035,N_1259);
xor U1780 (N_1780,N_1169,N_1240);
nor U1781 (N_1781,N_1211,N_1382);
xor U1782 (N_1782,N_1151,N_1029);
xor U1783 (N_1783,N_1131,N_1454);
or U1784 (N_1784,N_1027,N_1282);
or U1785 (N_1785,N_1345,N_1502);
xnor U1786 (N_1786,N_1106,N_928);
nand U1787 (N_1787,N_1103,N_1548);
nand U1788 (N_1788,N_903,N_1542);
or U1789 (N_1789,N_940,N_1078);
nor U1790 (N_1790,N_1189,N_876);
xnor U1791 (N_1791,N_948,N_1243);
nand U1792 (N_1792,N_1473,N_1135);
nor U1793 (N_1793,N_1364,N_1504);
nor U1794 (N_1794,N_1092,N_1568);
nand U1795 (N_1795,N_1474,N_1251);
xor U1796 (N_1796,N_871,N_1500);
nor U1797 (N_1797,N_979,N_949);
and U1798 (N_1798,N_839,N_1289);
nor U1799 (N_1799,N_1584,N_1320);
and U1800 (N_1800,N_922,N_1114);
xor U1801 (N_1801,N_1319,N_1266);
xnor U1802 (N_1802,N_1413,N_1313);
nor U1803 (N_1803,N_1337,N_1456);
or U1804 (N_1804,N_1541,N_1325);
nor U1805 (N_1805,N_1354,N_898);
nand U1806 (N_1806,N_1094,N_1150);
nor U1807 (N_1807,N_1272,N_1252);
xor U1808 (N_1808,N_1412,N_1310);
xor U1809 (N_1809,N_1086,N_1400);
and U1810 (N_1810,N_1540,N_834);
and U1811 (N_1811,N_1000,N_1472);
or U1812 (N_1812,N_1064,N_1047);
or U1813 (N_1813,N_889,N_981);
xnor U1814 (N_1814,N_1470,N_1245);
nand U1815 (N_1815,N_1042,N_844);
and U1816 (N_1816,N_810,N_1475);
and U1817 (N_1817,N_1539,N_1119);
nor U1818 (N_1818,N_818,N_1318);
or U1819 (N_1819,N_1051,N_1576);
or U1820 (N_1820,N_1370,N_1126);
or U1821 (N_1821,N_1137,N_1386);
nand U1822 (N_1822,N_1009,N_1045);
nor U1823 (N_1823,N_967,N_1109);
or U1824 (N_1824,N_932,N_946);
nor U1825 (N_1825,N_836,N_1330);
nor U1826 (N_1826,N_1434,N_874);
and U1827 (N_1827,N_826,N_822);
nand U1828 (N_1828,N_1142,N_1173);
and U1829 (N_1829,N_1315,N_1210);
nand U1830 (N_1830,N_1239,N_1099);
nor U1831 (N_1831,N_1343,N_1123);
xor U1832 (N_1832,N_1196,N_1384);
nor U1833 (N_1833,N_1530,N_1427);
or U1834 (N_1834,N_1484,N_1543);
nor U1835 (N_1835,N_1129,N_1088);
xor U1836 (N_1836,N_1231,N_1280);
nand U1837 (N_1837,N_924,N_1329);
nand U1838 (N_1838,N_1290,N_1258);
nand U1839 (N_1839,N_1185,N_1145);
nor U1840 (N_1840,N_1338,N_1227);
nor U1841 (N_1841,N_1582,N_970);
nand U1842 (N_1842,N_980,N_1281);
nand U1843 (N_1843,N_1275,N_1520);
nor U1844 (N_1844,N_1562,N_929);
xor U1845 (N_1845,N_1527,N_1144);
or U1846 (N_1846,N_1276,N_861);
and U1847 (N_1847,N_1199,N_1132);
nand U1848 (N_1848,N_961,N_1193);
and U1849 (N_1849,N_1204,N_1596);
or U1850 (N_1850,N_870,N_1161);
nand U1851 (N_1851,N_1079,N_851);
nand U1852 (N_1852,N_963,N_1133);
nand U1853 (N_1853,N_1381,N_1439);
nor U1854 (N_1854,N_1428,N_1066);
and U1855 (N_1855,N_1053,N_1080);
or U1856 (N_1856,N_1015,N_1580);
nand U1857 (N_1857,N_1435,N_1260);
nor U1858 (N_1858,N_1397,N_973);
and U1859 (N_1859,N_1509,N_1287);
and U1860 (N_1860,N_1519,N_1442);
nand U1861 (N_1861,N_1113,N_1032);
nand U1862 (N_1862,N_1317,N_1324);
xnor U1863 (N_1863,N_1487,N_987);
nor U1864 (N_1864,N_1205,N_1594);
nand U1865 (N_1865,N_1444,N_900);
or U1866 (N_1866,N_1307,N_1120);
and U1867 (N_1867,N_944,N_996);
nor U1868 (N_1868,N_911,N_959);
nand U1869 (N_1869,N_1023,N_1203);
xor U1870 (N_1870,N_1466,N_1396);
and U1871 (N_1871,N_1573,N_1531);
or U1872 (N_1872,N_1005,N_1069);
nor U1873 (N_1873,N_1147,N_872);
and U1874 (N_1874,N_1468,N_1271);
nor U1875 (N_1875,N_1419,N_1220);
xnor U1876 (N_1876,N_1127,N_1425);
nor U1877 (N_1877,N_1377,N_1224);
nor U1878 (N_1878,N_1589,N_1448);
and U1879 (N_1879,N_1237,N_1105);
xor U1880 (N_1880,N_873,N_833);
xnor U1881 (N_1881,N_1060,N_1383);
xnor U1882 (N_1882,N_1399,N_1390);
and U1883 (N_1883,N_887,N_1286);
nor U1884 (N_1884,N_1083,N_1344);
nand U1885 (N_1885,N_1093,N_843);
nand U1886 (N_1886,N_1256,N_805);
nand U1887 (N_1887,N_1257,N_1477);
xnor U1888 (N_1888,N_998,N_1234);
nor U1889 (N_1889,N_1476,N_808);
nand U1890 (N_1890,N_1176,N_1297);
xnor U1891 (N_1891,N_1011,N_1340);
nand U1892 (N_1892,N_1238,N_1598);
nand U1893 (N_1893,N_1457,N_831);
xor U1894 (N_1894,N_920,N_1406);
nor U1895 (N_1895,N_1152,N_896);
and U1896 (N_1896,N_1511,N_1513);
or U1897 (N_1897,N_1154,N_1423);
nor U1898 (N_1898,N_1002,N_1163);
or U1899 (N_1899,N_1517,N_1283);
nand U1900 (N_1900,N_840,N_1168);
nand U1901 (N_1901,N_1415,N_842);
nor U1902 (N_1902,N_1117,N_1136);
nor U1903 (N_1903,N_855,N_1178);
nor U1904 (N_1904,N_1085,N_1550);
nand U1905 (N_1905,N_1288,N_1516);
and U1906 (N_1906,N_1233,N_1380);
nand U1907 (N_1907,N_1478,N_1192);
nor U1908 (N_1908,N_1036,N_1055);
and U1909 (N_1909,N_1459,N_1532);
and U1910 (N_1910,N_1181,N_1452);
nor U1911 (N_1911,N_1201,N_1191);
nor U1912 (N_1912,N_1485,N_1451);
nor U1913 (N_1913,N_803,N_1588);
or U1914 (N_1914,N_921,N_1574);
nand U1915 (N_1915,N_1138,N_1404);
nand U1916 (N_1916,N_860,N_1246);
and U1917 (N_1917,N_1050,N_847);
nor U1918 (N_1918,N_926,N_1558);
nor U1919 (N_1919,N_1304,N_1024);
nor U1920 (N_1920,N_1194,N_1056);
nor U1921 (N_1921,N_1116,N_966);
xor U1922 (N_1922,N_1440,N_1551);
and U1923 (N_1923,N_1515,N_1391);
and U1924 (N_1924,N_800,N_811);
xor U1925 (N_1925,N_1521,N_1553);
or U1926 (N_1926,N_1585,N_1219);
and U1927 (N_1927,N_935,N_925);
nand U1928 (N_1928,N_1524,N_1357);
and U1929 (N_1929,N_941,N_1248);
xor U1930 (N_1930,N_1149,N_1299);
nor U1931 (N_1931,N_1436,N_1253);
and U1932 (N_1932,N_1342,N_821);
or U1933 (N_1933,N_1225,N_1230);
xnor U1934 (N_1934,N_1529,N_942);
xor U1935 (N_1935,N_856,N_1446);
nor U1936 (N_1936,N_1146,N_1577);
and U1937 (N_1937,N_1426,N_858);
nand U1938 (N_1938,N_825,N_859);
nand U1939 (N_1939,N_835,N_1111);
xor U1940 (N_1940,N_1157,N_1443);
nand U1941 (N_1941,N_1244,N_1134);
and U1942 (N_1942,N_1156,N_1449);
or U1943 (N_1943,N_1003,N_1408);
xor U1944 (N_1944,N_1316,N_1048);
and U1945 (N_1945,N_1302,N_1389);
nand U1946 (N_1946,N_974,N_1308);
xnor U1947 (N_1947,N_869,N_881);
nor U1948 (N_1948,N_1579,N_1222);
xnor U1949 (N_1949,N_1249,N_1499);
or U1950 (N_1950,N_897,N_1469);
and U1951 (N_1951,N_883,N_1581);
nor U1952 (N_1952,N_1599,N_893);
nand U1953 (N_1953,N_1394,N_901);
xnor U1954 (N_1954,N_1549,N_1102);
xnor U1955 (N_1955,N_1075,N_1030);
xnor U1956 (N_1956,N_1482,N_1298);
and U1957 (N_1957,N_882,N_817);
and U1958 (N_1958,N_1044,N_1184);
nor U1959 (N_1959,N_1505,N_892);
xnor U1960 (N_1960,N_990,N_916);
and U1961 (N_1961,N_1232,N_1356);
and U1962 (N_1962,N_1566,N_1491);
nor U1963 (N_1963,N_986,N_1180);
or U1964 (N_1964,N_1296,N_999);
or U1965 (N_1965,N_1097,N_1494);
xor U1966 (N_1966,N_1431,N_1141);
nand U1967 (N_1967,N_1038,N_824);
xnor U1968 (N_1968,N_1569,N_1460);
and U1969 (N_1969,N_1143,N_854);
nand U1970 (N_1970,N_1033,N_1471);
or U1971 (N_1971,N_1202,N_1462);
nand U1972 (N_1972,N_814,N_1533);
and U1973 (N_1973,N_972,N_954);
xor U1974 (N_1974,N_1292,N_1424);
nand U1975 (N_1975,N_1081,N_977);
nor U1976 (N_1976,N_886,N_988);
and U1977 (N_1977,N_930,N_1416);
and U1978 (N_1978,N_1526,N_1523);
nand U1979 (N_1979,N_1208,N_806);
and U1980 (N_1980,N_956,N_1347);
or U1981 (N_1981,N_1037,N_1049);
nand U1982 (N_1982,N_1043,N_878);
nor U1983 (N_1983,N_995,N_1188);
xor U1984 (N_1984,N_1174,N_1052);
xor U1985 (N_1985,N_1082,N_1190);
or U1986 (N_1986,N_1139,N_936);
nor U1987 (N_1987,N_1496,N_1433);
nor U1988 (N_1988,N_1140,N_1366);
or U1989 (N_1989,N_1463,N_1301);
or U1990 (N_1990,N_849,N_1110);
xnor U1991 (N_1991,N_867,N_830);
and U1992 (N_1992,N_1447,N_1065);
or U1993 (N_1993,N_1197,N_904);
or U1994 (N_1994,N_1323,N_1112);
nor U1995 (N_1995,N_992,N_1355);
xor U1996 (N_1996,N_1186,N_1101);
and U1997 (N_1997,N_1593,N_1108);
xor U1998 (N_1998,N_1264,N_1510);
xnor U1999 (N_1999,N_819,N_1379);
nand U2000 (N_2000,N_1303,N_1132);
nor U2001 (N_2001,N_841,N_885);
and U2002 (N_2002,N_1530,N_1213);
and U2003 (N_2003,N_1356,N_1202);
or U2004 (N_2004,N_824,N_1542);
xnor U2005 (N_2005,N_998,N_863);
nand U2006 (N_2006,N_1116,N_1567);
nand U2007 (N_2007,N_1070,N_1208);
xor U2008 (N_2008,N_905,N_1024);
nor U2009 (N_2009,N_1490,N_811);
and U2010 (N_2010,N_1050,N_800);
xnor U2011 (N_2011,N_1204,N_1177);
nand U2012 (N_2012,N_1062,N_964);
nor U2013 (N_2013,N_1484,N_1479);
or U2014 (N_2014,N_1415,N_806);
xor U2015 (N_2015,N_1211,N_1410);
nor U2016 (N_2016,N_870,N_1399);
nor U2017 (N_2017,N_1433,N_1579);
nand U2018 (N_2018,N_1335,N_1572);
and U2019 (N_2019,N_1030,N_1026);
and U2020 (N_2020,N_948,N_1029);
nand U2021 (N_2021,N_1000,N_832);
xor U2022 (N_2022,N_969,N_1063);
or U2023 (N_2023,N_940,N_1038);
nand U2024 (N_2024,N_897,N_1220);
nor U2025 (N_2025,N_950,N_879);
nor U2026 (N_2026,N_1372,N_863);
nor U2027 (N_2027,N_1292,N_1562);
nand U2028 (N_2028,N_1079,N_827);
nand U2029 (N_2029,N_1296,N_1051);
nand U2030 (N_2030,N_817,N_1016);
nor U2031 (N_2031,N_1102,N_1324);
nor U2032 (N_2032,N_1180,N_898);
and U2033 (N_2033,N_1106,N_1222);
xor U2034 (N_2034,N_1200,N_1049);
nor U2035 (N_2035,N_1419,N_853);
xnor U2036 (N_2036,N_915,N_1593);
xor U2037 (N_2037,N_945,N_1371);
nor U2038 (N_2038,N_1059,N_1207);
xor U2039 (N_2039,N_1268,N_1502);
and U2040 (N_2040,N_1042,N_1184);
or U2041 (N_2041,N_1200,N_1587);
xor U2042 (N_2042,N_855,N_892);
and U2043 (N_2043,N_1479,N_1010);
xnor U2044 (N_2044,N_1514,N_882);
nand U2045 (N_2045,N_1237,N_1153);
xnor U2046 (N_2046,N_826,N_1440);
or U2047 (N_2047,N_1390,N_1336);
and U2048 (N_2048,N_1494,N_1454);
and U2049 (N_2049,N_1519,N_1345);
xor U2050 (N_2050,N_1583,N_889);
nor U2051 (N_2051,N_1020,N_1193);
nand U2052 (N_2052,N_1097,N_1188);
nand U2053 (N_2053,N_1295,N_1550);
or U2054 (N_2054,N_892,N_1173);
nor U2055 (N_2055,N_1264,N_870);
and U2056 (N_2056,N_1000,N_1154);
or U2057 (N_2057,N_1509,N_942);
xnor U2058 (N_2058,N_1284,N_1054);
nor U2059 (N_2059,N_1025,N_1365);
or U2060 (N_2060,N_1288,N_1376);
xor U2061 (N_2061,N_955,N_990);
xnor U2062 (N_2062,N_958,N_990);
or U2063 (N_2063,N_967,N_1090);
nor U2064 (N_2064,N_969,N_1529);
and U2065 (N_2065,N_1176,N_1562);
and U2066 (N_2066,N_1311,N_1042);
xnor U2067 (N_2067,N_890,N_1485);
or U2068 (N_2068,N_1475,N_836);
nand U2069 (N_2069,N_1338,N_1407);
nand U2070 (N_2070,N_806,N_1224);
nand U2071 (N_2071,N_850,N_1238);
nand U2072 (N_2072,N_1536,N_1459);
nand U2073 (N_2073,N_1001,N_935);
or U2074 (N_2074,N_1200,N_1462);
nand U2075 (N_2075,N_933,N_1326);
xor U2076 (N_2076,N_1263,N_845);
nand U2077 (N_2077,N_906,N_1055);
nor U2078 (N_2078,N_1116,N_1020);
or U2079 (N_2079,N_911,N_914);
or U2080 (N_2080,N_1006,N_949);
or U2081 (N_2081,N_899,N_933);
or U2082 (N_2082,N_860,N_1331);
or U2083 (N_2083,N_1402,N_1473);
and U2084 (N_2084,N_1474,N_1094);
nor U2085 (N_2085,N_1464,N_1098);
and U2086 (N_2086,N_1469,N_1505);
xnor U2087 (N_2087,N_1385,N_1577);
or U2088 (N_2088,N_1131,N_1335);
xor U2089 (N_2089,N_1464,N_1223);
and U2090 (N_2090,N_1511,N_1372);
nand U2091 (N_2091,N_861,N_1072);
and U2092 (N_2092,N_1449,N_1380);
nand U2093 (N_2093,N_1187,N_1154);
xnor U2094 (N_2094,N_1437,N_1232);
or U2095 (N_2095,N_1492,N_1228);
and U2096 (N_2096,N_1064,N_1332);
or U2097 (N_2097,N_1430,N_1592);
nand U2098 (N_2098,N_922,N_982);
nor U2099 (N_2099,N_854,N_1277);
xor U2100 (N_2100,N_1206,N_965);
nand U2101 (N_2101,N_1121,N_929);
or U2102 (N_2102,N_1186,N_965);
xnor U2103 (N_2103,N_1218,N_1554);
or U2104 (N_2104,N_1564,N_1447);
xnor U2105 (N_2105,N_1310,N_1460);
and U2106 (N_2106,N_1078,N_1441);
or U2107 (N_2107,N_848,N_1177);
and U2108 (N_2108,N_1268,N_1261);
or U2109 (N_2109,N_1216,N_944);
and U2110 (N_2110,N_1555,N_1354);
or U2111 (N_2111,N_834,N_1111);
nand U2112 (N_2112,N_1010,N_1534);
or U2113 (N_2113,N_1108,N_1368);
nand U2114 (N_2114,N_910,N_1410);
xor U2115 (N_2115,N_1575,N_1114);
or U2116 (N_2116,N_1089,N_1071);
nor U2117 (N_2117,N_943,N_1224);
nor U2118 (N_2118,N_1588,N_1090);
and U2119 (N_2119,N_1078,N_1420);
nand U2120 (N_2120,N_1022,N_925);
nor U2121 (N_2121,N_1427,N_1206);
nor U2122 (N_2122,N_1173,N_1377);
xnor U2123 (N_2123,N_858,N_1149);
nor U2124 (N_2124,N_836,N_950);
and U2125 (N_2125,N_1482,N_898);
nor U2126 (N_2126,N_1039,N_845);
nor U2127 (N_2127,N_1341,N_1360);
and U2128 (N_2128,N_1377,N_1312);
xnor U2129 (N_2129,N_1027,N_1242);
xnor U2130 (N_2130,N_1405,N_1577);
nor U2131 (N_2131,N_1395,N_875);
and U2132 (N_2132,N_1317,N_1334);
nand U2133 (N_2133,N_859,N_937);
or U2134 (N_2134,N_1468,N_1493);
and U2135 (N_2135,N_1486,N_1581);
xor U2136 (N_2136,N_831,N_1044);
or U2137 (N_2137,N_1372,N_1294);
xnor U2138 (N_2138,N_1103,N_1055);
nand U2139 (N_2139,N_1453,N_1464);
nor U2140 (N_2140,N_1371,N_1282);
nor U2141 (N_2141,N_1305,N_909);
xor U2142 (N_2142,N_1294,N_1553);
nand U2143 (N_2143,N_1011,N_1048);
nand U2144 (N_2144,N_908,N_1171);
nand U2145 (N_2145,N_919,N_806);
or U2146 (N_2146,N_1197,N_1285);
or U2147 (N_2147,N_1024,N_1335);
xnor U2148 (N_2148,N_1412,N_1026);
and U2149 (N_2149,N_1462,N_821);
or U2150 (N_2150,N_1305,N_809);
nor U2151 (N_2151,N_1402,N_1048);
nand U2152 (N_2152,N_1366,N_874);
nand U2153 (N_2153,N_876,N_1107);
and U2154 (N_2154,N_1105,N_1178);
nor U2155 (N_2155,N_1249,N_1362);
and U2156 (N_2156,N_1037,N_1549);
nor U2157 (N_2157,N_887,N_983);
xor U2158 (N_2158,N_1465,N_1380);
or U2159 (N_2159,N_1206,N_1265);
and U2160 (N_2160,N_1549,N_863);
xor U2161 (N_2161,N_1394,N_854);
nor U2162 (N_2162,N_1114,N_1577);
and U2163 (N_2163,N_1382,N_1327);
and U2164 (N_2164,N_1229,N_838);
and U2165 (N_2165,N_905,N_1003);
nor U2166 (N_2166,N_1088,N_1256);
nor U2167 (N_2167,N_1078,N_1132);
or U2168 (N_2168,N_1052,N_812);
xor U2169 (N_2169,N_1377,N_1248);
xnor U2170 (N_2170,N_1109,N_1494);
xor U2171 (N_2171,N_1076,N_930);
and U2172 (N_2172,N_1138,N_1140);
or U2173 (N_2173,N_1280,N_1437);
nand U2174 (N_2174,N_812,N_827);
xor U2175 (N_2175,N_1446,N_1469);
and U2176 (N_2176,N_1499,N_1279);
or U2177 (N_2177,N_903,N_1069);
and U2178 (N_2178,N_846,N_1547);
nor U2179 (N_2179,N_1099,N_855);
and U2180 (N_2180,N_1349,N_1193);
nor U2181 (N_2181,N_829,N_1489);
and U2182 (N_2182,N_1486,N_1345);
and U2183 (N_2183,N_819,N_1090);
nand U2184 (N_2184,N_1570,N_1008);
nand U2185 (N_2185,N_1277,N_983);
nand U2186 (N_2186,N_1567,N_849);
nor U2187 (N_2187,N_951,N_981);
and U2188 (N_2188,N_1423,N_1422);
and U2189 (N_2189,N_968,N_1319);
or U2190 (N_2190,N_868,N_1295);
and U2191 (N_2191,N_1308,N_1069);
and U2192 (N_2192,N_1591,N_869);
or U2193 (N_2193,N_922,N_947);
nand U2194 (N_2194,N_1548,N_1287);
nor U2195 (N_2195,N_869,N_1081);
or U2196 (N_2196,N_1223,N_1264);
or U2197 (N_2197,N_1326,N_976);
xnor U2198 (N_2198,N_1024,N_1127);
nor U2199 (N_2199,N_1353,N_1137);
nand U2200 (N_2200,N_1475,N_1545);
nor U2201 (N_2201,N_1265,N_1083);
nor U2202 (N_2202,N_1305,N_1549);
xnor U2203 (N_2203,N_1291,N_1176);
xor U2204 (N_2204,N_1564,N_1290);
or U2205 (N_2205,N_1464,N_943);
and U2206 (N_2206,N_1309,N_1076);
and U2207 (N_2207,N_1558,N_984);
and U2208 (N_2208,N_991,N_1456);
nand U2209 (N_2209,N_1342,N_1262);
or U2210 (N_2210,N_898,N_1540);
nor U2211 (N_2211,N_1339,N_1225);
nand U2212 (N_2212,N_1394,N_1480);
and U2213 (N_2213,N_914,N_816);
xnor U2214 (N_2214,N_1591,N_1367);
nor U2215 (N_2215,N_1511,N_972);
or U2216 (N_2216,N_905,N_1135);
or U2217 (N_2217,N_1542,N_1537);
nand U2218 (N_2218,N_1298,N_1407);
or U2219 (N_2219,N_920,N_1518);
or U2220 (N_2220,N_1414,N_1141);
xor U2221 (N_2221,N_1161,N_1352);
and U2222 (N_2222,N_1367,N_1480);
nor U2223 (N_2223,N_1376,N_832);
or U2224 (N_2224,N_1154,N_1554);
nand U2225 (N_2225,N_829,N_890);
xnor U2226 (N_2226,N_1458,N_932);
nor U2227 (N_2227,N_1063,N_1397);
and U2228 (N_2228,N_1478,N_1417);
or U2229 (N_2229,N_860,N_1356);
and U2230 (N_2230,N_930,N_1049);
nor U2231 (N_2231,N_1535,N_1357);
or U2232 (N_2232,N_814,N_1014);
or U2233 (N_2233,N_1188,N_1570);
or U2234 (N_2234,N_1266,N_1300);
xnor U2235 (N_2235,N_926,N_858);
nand U2236 (N_2236,N_1295,N_1194);
xnor U2237 (N_2237,N_1053,N_1398);
nand U2238 (N_2238,N_951,N_1315);
nand U2239 (N_2239,N_1353,N_1594);
xor U2240 (N_2240,N_1479,N_1232);
nand U2241 (N_2241,N_921,N_1128);
nor U2242 (N_2242,N_1373,N_827);
and U2243 (N_2243,N_853,N_1445);
and U2244 (N_2244,N_1109,N_1471);
xor U2245 (N_2245,N_1507,N_1313);
nand U2246 (N_2246,N_1178,N_1119);
xnor U2247 (N_2247,N_1086,N_1032);
and U2248 (N_2248,N_1109,N_1501);
or U2249 (N_2249,N_828,N_1277);
nor U2250 (N_2250,N_1586,N_1307);
nand U2251 (N_2251,N_1582,N_1410);
xnor U2252 (N_2252,N_1242,N_921);
or U2253 (N_2253,N_1591,N_1125);
nor U2254 (N_2254,N_1091,N_1026);
nor U2255 (N_2255,N_1098,N_1113);
xnor U2256 (N_2256,N_1553,N_1188);
or U2257 (N_2257,N_938,N_1039);
nand U2258 (N_2258,N_952,N_1172);
and U2259 (N_2259,N_1342,N_1001);
nor U2260 (N_2260,N_1425,N_1058);
xor U2261 (N_2261,N_1383,N_994);
nand U2262 (N_2262,N_1589,N_978);
or U2263 (N_2263,N_841,N_953);
nor U2264 (N_2264,N_1599,N_1066);
nor U2265 (N_2265,N_882,N_1342);
nand U2266 (N_2266,N_1041,N_1182);
or U2267 (N_2267,N_1304,N_1282);
nor U2268 (N_2268,N_1010,N_1291);
nor U2269 (N_2269,N_1446,N_1312);
nand U2270 (N_2270,N_1591,N_912);
nand U2271 (N_2271,N_1237,N_1191);
and U2272 (N_2272,N_1120,N_805);
and U2273 (N_2273,N_1164,N_898);
or U2274 (N_2274,N_1358,N_1162);
or U2275 (N_2275,N_1017,N_1021);
nand U2276 (N_2276,N_933,N_902);
and U2277 (N_2277,N_993,N_1092);
nand U2278 (N_2278,N_801,N_1513);
and U2279 (N_2279,N_1245,N_1354);
and U2280 (N_2280,N_1293,N_890);
nand U2281 (N_2281,N_1559,N_1367);
and U2282 (N_2282,N_1581,N_1518);
or U2283 (N_2283,N_884,N_959);
nor U2284 (N_2284,N_1479,N_837);
nor U2285 (N_2285,N_1014,N_831);
nand U2286 (N_2286,N_909,N_919);
or U2287 (N_2287,N_1148,N_1296);
nand U2288 (N_2288,N_1149,N_874);
nand U2289 (N_2289,N_1548,N_1335);
and U2290 (N_2290,N_1039,N_825);
xor U2291 (N_2291,N_1154,N_1589);
or U2292 (N_2292,N_1549,N_1565);
nor U2293 (N_2293,N_1253,N_1529);
or U2294 (N_2294,N_808,N_1593);
or U2295 (N_2295,N_948,N_1362);
and U2296 (N_2296,N_811,N_1320);
xor U2297 (N_2297,N_1499,N_1099);
or U2298 (N_2298,N_1326,N_1287);
nor U2299 (N_2299,N_1272,N_1108);
nand U2300 (N_2300,N_867,N_1411);
nor U2301 (N_2301,N_1470,N_1453);
or U2302 (N_2302,N_1562,N_1094);
xor U2303 (N_2303,N_1575,N_1152);
nor U2304 (N_2304,N_1267,N_1336);
nand U2305 (N_2305,N_1441,N_1374);
xor U2306 (N_2306,N_1220,N_1106);
nand U2307 (N_2307,N_893,N_1011);
and U2308 (N_2308,N_852,N_1587);
xor U2309 (N_2309,N_1131,N_1472);
xor U2310 (N_2310,N_1552,N_1214);
and U2311 (N_2311,N_1095,N_1437);
or U2312 (N_2312,N_1408,N_1121);
nor U2313 (N_2313,N_1359,N_985);
or U2314 (N_2314,N_1273,N_1058);
nor U2315 (N_2315,N_858,N_1485);
nand U2316 (N_2316,N_871,N_807);
nor U2317 (N_2317,N_1309,N_1218);
xnor U2318 (N_2318,N_1378,N_1549);
nand U2319 (N_2319,N_1035,N_1005);
and U2320 (N_2320,N_872,N_1166);
and U2321 (N_2321,N_1510,N_839);
nand U2322 (N_2322,N_984,N_1391);
nor U2323 (N_2323,N_1431,N_1343);
nor U2324 (N_2324,N_989,N_1437);
xor U2325 (N_2325,N_853,N_825);
nor U2326 (N_2326,N_867,N_1103);
nand U2327 (N_2327,N_1248,N_860);
and U2328 (N_2328,N_913,N_1552);
nand U2329 (N_2329,N_1492,N_1204);
and U2330 (N_2330,N_1378,N_1504);
and U2331 (N_2331,N_1498,N_1201);
nand U2332 (N_2332,N_1014,N_1397);
xor U2333 (N_2333,N_1245,N_1560);
nand U2334 (N_2334,N_1091,N_810);
nand U2335 (N_2335,N_994,N_822);
nand U2336 (N_2336,N_1197,N_1078);
and U2337 (N_2337,N_978,N_880);
nor U2338 (N_2338,N_1410,N_1079);
xor U2339 (N_2339,N_1491,N_1374);
and U2340 (N_2340,N_1098,N_918);
nand U2341 (N_2341,N_1123,N_965);
nand U2342 (N_2342,N_903,N_1212);
nor U2343 (N_2343,N_936,N_959);
xor U2344 (N_2344,N_1304,N_1485);
nand U2345 (N_2345,N_948,N_1229);
or U2346 (N_2346,N_1493,N_1573);
xor U2347 (N_2347,N_1124,N_1205);
and U2348 (N_2348,N_952,N_1358);
nor U2349 (N_2349,N_1315,N_1052);
nand U2350 (N_2350,N_1588,N_991);
xor U2351 (N_2351,N_1564,N_1584);
and U2352 (N_2352,N_1342,N_1530);
nand U2353 (N_2353,N_936,N_1515);
nand U2354 (N_2354,N_1314,N_1477);
xnor U2355 (N_2355,N_1142,N_1522);
or U2356 (N_2356,N_1097,N_1273);
nor U2357 (N_2357,N_1503,N_1183);
xnor U2358 (N_2358,N_1302,N_1471);
and U2359 (N_2359,N_1005,N_1518);
nand U2360 (N_2360,N_1500,N_812);
xor U2361 (N_2361,N_1150,N_1436);
nand U2362 (N_2362,N_1341,N_948);
nor U2363 (N_2363,N_1271,N_1160);
or U2364 (N_2364,N_1314,N_1502);
and U2365 (N_2365,N_1587,N_1107);
xnor U2366 (N_2366,N_1182,N_1195);
and U2367 (N_2367,N_888,N_1530);
xnor U2368 (N_2368,N_1326,N_1134);
nor U2369 (N_2369,N_1191,N_853);
nor U2370 (N_2370,N_801,N_1210);
or U2371 (N_2371,N_1208,N_1279);
or U2372 (N_2372,N_989,N_1509);
and U2373 (N_2373,N_1403,N_928);
nor U2374 (N_2374,N_1301,N_996);
or U2375 (N_2375,N_1422,N_1355);
nand U2376 (N_2376,N_1003,N_894);
or U2377 (N_2377,N_1329,N_1222);
and U2378 (N_2378,N_1103,N_1194);
xnor U2379 (N_2379,N_1071,N_1193);
xnor U2380 (N_2380,N_1266,N_1541);
nor U2381 (N_2381,N_1236,N_1207);
xnor U2382 (N_2382,N_1013,N_891);
nand U2383 (N_2383,N_1331,N_1014);
nand U2384 (N_2384,N_1344,N_1225);
nor U2385 (N_2385,N_1413,N_927);
and U2386 (N_2386,N_1435,N_858);
xor U2387 (N_2387,N_1104,N_919);
nor U2388 (N_2388,N_1272,N_1568);
nand U2389 (N_2389,N_978,N_896);
nand U2390 (N_2390,N_1119,N_803);
and U2391 (N_2391,N_1341,N_1027);
or U2392 (N_2392,N_1050,N_1243);
and U2393 (N_2393,N_1404,N_1456);
nor U2394 (N_2394,N_1011,N_1551);
nand U2395 (N_2395,N_1571,N_1533);
nor U2396 (N_2396,N_1032,N_1542);
nor U2397 (N_2397,N_915,N_1365);
nand U2398 (N_2398,N_1118,N_1405);
nand U2399 (N_2399,N_1329,N_1226);
or U2400 (N_2400,N_1874,N_1899);
and U2401 (N_2401,N_1889,N_1677);
or U2402 (N_2402,N_1991,N_2052);
xnor U2403 (N_2403,N_2225,N_1912);
and U2404 (N_2404,N_1931,N_2131);
or U2405 (N_2405,N_1668,N_1978);
and U2406 (N_2406,N_2371,N_1855);
and U2407 (N_2407,N_1800,N_1806);
or U2408 (N_2408,N_2203,N_1607);
nor U2409 (N_2409,N_2228,N_2329);
and U2410 (N_2410,N_2336,N_2251);
and U2411 (N_2411,N_1670,N_1919);
nand U2412 (N_2412,N_2390,N_2397);
nand U2413 (N_2413,N_2367,N_1826);
nor U2414 (N_2414,N_2373,N_2326);
xnor U2415 (N_2415,N_1913,N_1904);
and U2416 (N_2416,N_2039,N_2117);
and U2417 (N_2417,N_2244,N_1842);
or U2418 (N_2418,N_2388,N_1831);
xor U2419 (N_2419,N_2159,N_2285);
nand U2420 (N_2420,N_2176,N_1704);
nand U2421 (N_2421,N_1972,N_1807);
nand U2422 (N_2422,N_2002,N_1973);
nand U2423 (N_2423,N_1953,N_1795);
and U2424 (N_2424,N_2182,N_2348);
nand U2425 (N_2425,N_1679,N_2211);
nand U2426 (N_2426,N_1986,N_2316);
or U2427 (N_2427,N_1849,N_2339);
nor U2428 (N_2428,N_1819,N_1603);
and U2429 (N_2429,N_1737,N_1772);
or U2430 (N_2430,N_1753,N_1735);
nor U2431 (N_2431,N_1657,N_1738);
and U2432 (N_2432,N_1703,N_1685);
xnor U2433 (N_2433,N_1941,N_1936);
and U2434 (N_2434,N_1834,N_1769);
or U2435 (N_2435,N_1960,N_1959);
nor U2436 (N_2436,N_1851,N_1693);
or U2437 (N_2437,N_1902,N_1832);
xnor U2438 (N_2438,N_1688,N_2255);
or U2439 (N_2439,N_1722,N_2178);
or U2440 (N_2440,N_2195,N_1761);
nor U2441 (N_2441,N_2340,N_2139);
and U2442 (N_2442,N_2116,N_1768);
xnor U2443 (N_2443,N_1837,N_1635);
or U2444 (N_2444,N_2238,N_1751);
xor U2445 (N_2445,N_2273,N_1955);
and U2446 (N_2446,N_2222,N_1905);
xor U2447 (N_2447,N_1921,N_2017);
and U2448 (N_2448,N_2383,N_2240);
nor U2449 (N_2449,N_2158,N_2020);
xor U2450 (N_2450,N_1760,N_1847);
nor U2451 (N_2451,N_2208,N_2346);
and U2452 (N_2452,N_2266,N_2028);
or U2453 (N_2453,N_1667,N_1746);
nand U2454 (N_2454,N_1713,N_1662);
xor U2455 (N_2455,N_2379,N_2221);
nor U2456 (N_2456,N_1928,N_1700);
or U2457 (N_2457,N_1780,N_2207);
nor U2458 (N_2458,N_1716,N_2217);
xor U2459 (N_2459,N_2179,N_2047);
and U2460 (N_2460,N_1830,N_2369);
xnor U2461 (N_2461,N_2130,N_2156);
xor U2462 (N_2462,N_1818,N_2059);
xnor U2463 (N_2463,N_1698,N_1814);
nor U2464 (N_2464,N_1995,N_1796);
xnor U2465 (N_2465,N_2107,N_2289);
or U2466 (N_2466,N_2065,N_2091);
nor U2467 (N_2467,N_2286,N_2387);
and U2468 (N_2468,N_1671,N_2302);
and U2469 (N_2469,N_2263,N_1648);
xnor U2470 (N_2470,N_2009,N_1721);
nand U2471 (N_2471,N_2145,N_2165);
xor U2472 (N_2472,N_2127,N_1985);
nor U2473 (N_2473,N_1997,N_2315);
and U2474 (N_2474,N_1625,N_2168);
nor U2475 (N_2475,N_2032,N_2301);
nor U2476 (N_2476,N_1621,N_2230);
and U2477 (N_2477,N_1647,N_1971);
and U2478 (N_2478,N_2331,N_2357);
xnor U2479 (N_2479,N_1894,N_2258);
or U2480 (N_2480,N_1803,N_1754);
xnor U2481 (N_2481,N_1695,N_1608);
xor U2482 (N_2482,N_2269,N_2354);
and U2483 (N_2483,N_2027,N_1639);
xnor U2484 (N_2484,N_2098,N_2325);
or U2485 (N_2485,N_2190,N_1654);
and U2486 (N_2486,N_2040,N_1665);
nand U2487 (N_2487,N_1739,N_1730);
and U2488 (N_2488,N_2134,N_1734);
or U2489 (N_2489,N_1797,N_1615);
or U2490 (N_2490,N_2186,N_1756);
and U2491 (N_2491,N_2295,N_1794);
nand U2492 (N_2492,N_1707,N_1788);
nand U2493 (N_2493,N_1645,N_2380);
nor U2494 (N_2494,N_2282,N_2236);
and U2495 (N_2495,N_2215,N_1990);
nand U2496 (N_2496,N_2100,N_2010);
and U2497 (N_2497,N_1669,N_2096);
or U2498 (N_2498,N_2046,N_2202);
xor U2499 (N_2499,N_2193,N_2389);
nor U2500 (N_2500,N_1619,N_1618);
xor U2501 (N_2501,N_2293,N_2092);
or U2502 (N_2502,N_1745,N_1964);
xnor U2503 (N_2503,N_2082,N_2259);
xnor U2504 (N_2504,N_1736,N_2344);
nand U2505 (N_2505,N_2265,N_2245);
or U2506 (N_2506,N_2035,N_2359);
nand U2507 (N_2507,N_1952,N_1873);
nor U2508 (N_2508,N_2055,N_1804);
or U2509 (N_2509,N_2093,N_1812);
nor U2510 (N_2510,N_2300,N_1929);
and U2511 (N_2511,N_2305,N_1845);
or U2512 (N_2512,N_2287,N_1970);
or U2513 (N_2513,N_2030,N_2112);
nand U2514 (N_2514,N_1755,N_1741);
or U2515 (N_2515,N_1610,N_1927);
or U2516 (N_2516,N_1701,N_2223);
and U2517 (N_2517,N_1763,N_2366);
nand U2518 (N_2518,N_2151,N_2235);
nand U2519 (N_2519,N_2088,N_1766);
xor U2520 (N_2520,N_1628,N_1752);
or U2521 (N_2521,N_2361,N_2123);
nand U2522 (N_2522,N_2114,N_2037);
and U2523 (N_2523,N_2386,N_2375);
and U2524 (N_2524,N_1916,N_1623);
or U2525 (N_2525,N_2162,N_1856);
xor U2526 (N_2526,N_2322,N_2142);
or U2527 (N_2527,N_2144,N_2070);
nor U2528 (N_2528,N_2256,N_1998);
xnor U2529 (N_2529,N_1785,N_1815);
nor U2530 (N_2530,N_2188,N_1809);
xor U2531 (N_2531,N_1731,N_1839);
and U2532 (N_2532,N_2050,N_1882);
xor U2533 (N_2533,N_2277,N_1881);
nand U2534 (N_2534,N_2137,N_2342);
nor U2535 (N_2535,N_1923,N_1965);
and U2536 (N_2536,N_1870,N_2081);
nand U2537 (N_2537,N_1903,N_2313);
or U2538 (N_2538,N_1655,N_1969);
or U2539 (N_2539,N_1664,N_1822);
or U2540 (N_2540,N_2033,N_2219);
nor U2541 (N_2541,N_1890,N_2353);
nand U2542 (N_2542,N_2038,N_1932);
or U2543 (N_2543,N_2013,N_2118);
and U2544 (N_2544,N_2220,N_1634);
and U2545 (N_2545,N_2053,N_2254);
nor U2546 (N_2546,N_1980,N_2119);
and U2547 (N_2547,N_2105,N_1641);
xnor U2548 (N_2548,N_2072,N_1827);
or U2549 (N_2549,N_2060,N_2253);
xor U2550 (N_2550,N_2062,N_1775);
or U2551 (N_2551,N_2011,N_2226);
nand U2552 (N_2552,N_1717,N_1644);
nand U2553 (N_2553,N_1656,N_2360);
nor U2554 (N_2554,N_2355,N_1816);
or U2555 (N_2555,N_2192,N_2095);
nand U2556 (N_2556,N_2057,N_1650);
or U2557 (N_2557,N_1757,N_2232);
nand U2558 (N_2558,N_2041,N_1974);
nand U2559 (N_2559,N_1900,N_1724);
nor U2560 (N_2560,N_2054,N_2174);
xor U2561 (N_2561,N_1793,N_2024);
nor U2562 (N_2562,N_1674,N_2304);
nor U2563 (N_2563,N_2381,N_2270);
or U2564 (N_2564,N_1954,N_1626);
or U2565 (N_2565,N_2078,N_2294);
xnor U2566 (N_2566,N_2163,N_2345);
xor U2567 (N_2567,N_1813,N_1779);
or U2568 (N_2568,N_2271,N_2278);
nand U2569 (N_2569,N_2362,N_1614);
and U2570 (N_2570,N_2323,N_2312);
and U2571 (N_2571,N_1999,N_1887);
nand U2572 (N_2572,N_2394,N_1786);
nand U2573 (N_2573,N_1801,N_2018);
nor U2574 (N_2574,N_2205,N_2372);
and U2575 (N_2575,N_2321,N_1629);
and U2576 (N_2576,N_2067,N_2272);
nor U2577 (N_2577,N_2043,N_1663);
nor U2578 (N_2578,N_2338,N_1767);
and U2579 (N_2579,N_1726,N_1939);
and U2580 (N_2580,N_2172,N_1778);
nand U2581 (N_2581,N_2309,N_1976);
xnor U2582 (N_2582,N_2352,N_2268);
nor U2583 (N_2583,N_1697,N_2169);
xnor U2584 (N_2584,N_1898,N_2104);
xor U2585 (N_2585,N_2187,N_1926);
xor U2586 (N_2586,N_1908,N_2370);
or U2587 (N_2587,N_2276,N_2080);
nand U2588 (N_2588,N_1861,N_1885);
and U2589 (N_2589,N_2141,N_1967);
xor U2590 (N_2590,N_1636,N_2297);
xnor U2591 (N_2591,N_2307,N_1850);
nor U2592 (N_2592,N_2153,N_1649);
nand U2593 (N_2593,N_1924,N_2110);
or U2594 (N_2594,N_2079,N_2022);
nand U2595 (N_2595,N_2173,N_2122);
or U2596 (N_2596,N_1732,N_1705);
xnor U2597 (N_2597,N_1702,N_1740);
nor U2598 (N_2598,N_2200,N_2003);
nand U2599 (N_2599,N_2347,N_2349);
nand U2600 (N_2600,N_1838,N_2196);
nand U2601 (N_2601,N_1787,N_2180);
or U2602 (N_2602,N_2183,N_2031);
nand U2603 (N_2603,N_1946,N_1863);
nor U2604 (N_2604,N_1875,N_1606);
or U2605 (N_2605,N_2281,N_1676);
or U2606 (N_2606,N_2292,N_1743);
nor U2607 (N_2607,N_1659,N_1854);
or U2608 (N_2608,N_2320,N_1872);
xnor U2609 (N_2609,N_2227,N_1930);
nand U2610 (N_2610,N_1948,N_1642);
nor U2611 (N_2611,N_2393,N_2029);
nor U2612 (N_2612,N_2101,N_2332);
and U2613 (N_2613,N_1977,N_1950);
and U2614 (N_2614,N_2194,N_2000);
and U2615 (N_2615,N_1661,N_1933);
nand U2616 (N_2616,N_2337,N_1880);
and U2617 (N_2617,N_1891,N_2016);
or U2618 (N_2618,N_1951,N_1984);
or U2619 (N_2619,N_2216,N_1867);
or U2620 (N_2620,N_2125,N_1947);
nand U2621 (N_2621,N_2121,N_1833);
or U2622 (N_2622,N_1683,N_1943);
nand U2623 (N_2623,N_2120,N_2191);
nor U2624 (N_2624,N_1949,N_1748);
xnor U2625 (N_2625,N_1802,N_2138);
xnor U2626 (N_2626,N_1937,N_2233);
nor U2627 (N_2627,N_2247,N_2181);
or U2628 (N_2628,N_1604,N_2314);
and U2629 (N_2629,N_1632,N_1859);
nand U2630 (N_2630,N_2036,N_2058);
or U2631 (N_2631,N_1733,N_2333);
and U2632 (N_2632,N_2257,N_1987);
nand U2633 (N_2633,N_2395,N_2385);
nand U2634 (N_2634,N_1600,N_1686);
xnor U2635 (N_2635,N_2275,N_1992);
xnor U2636 (N_2636,N_1725,N_1817);
xor U2637 (N_2637,N_1896,N_2056);
xnor U2638 (N_2638,N_1848,N_2102);
or U2639 (N_2639,N_2008,N_2076);
xor U2640 (N_2640,N_2063,N_1714);
and U2641 (N_2641,N_2262,N_1935);
nor U2642 (N_2642,N_1759,N_2274);
nand U2643 (N_2643,N_1956,N_1616);
and U2644 (N_2644,N_1765,N_1852);
and U2645 (N_2645,N_1824,N_2324);
and U2646 (N_2646,N_2264,N_2260);
or U2647 (N_2647,N_2214,N_1910);
or U2648 (N_2648,N_1934,N_2048);
and U2649 (N_2649,N_1771,N_2368);
xor U2650 (N_2650,N_2363,N_1602);
xor U2651 (N_2651,N_2239,N_1712);
xor U2652 (N_2652,N_1627,N_1694);
nand U2653 (N_2653,N_1773,N_1651);
nor U2654 (N_2654,N_1988,N_1710);
and U2655 (N_2655,N_2283,N_2006);
xor U2656 (N_2656,N_2068,N_1966);
xor U2657 (N_2657,N_2384,N_2136);
and U2658 (N_2658,N_1857,N_1811);
and U2659 (N_2659,N_1681,N_2106);
and U2660 (N_2660,N_1708,N_1605);
xor U2661 (N_2661,N_2087,N_2135);
nand U2662 (N_2662,N_1720,N_2201);
nand U2663 (N_2663,N_2288,N_2224);
nor U2664 (N_2664,N_1729,N_2124);
nand U2665 (N_2665,N_1790,N_1666);
xnor U2666 (N_2666,N_2001,N_1942);
or U2667 (N_2667,N_1633,N_2166);
nand U2668 (N_2668,N_2157,N_1911);
xor U2669 (N_2669,N_1958,N_2298);
or U2670 (N_2670,N_1624,N_2044);
nor U2671 (N_2671,N_1750,N_1783);
nand U2672 (N_2672,N_2167,N_1691);
xor U2673 (N_2673,N_1808,N_2356);
nand U2674 (N_2674,N_2376,N_2126);
and U2675 (N_2675,N_2132,N_1762);
or U2676 (N_2676,N_2160,N_2184);
and U2677 (N_2677,N_2197,N_2023);
nand U2678 (N_2678,N_1829,N_1853);
nor U2679 (N_2679,N_2382,N_2396);
nand U2680 (N_2680,N_1652,N_1637);
or U2681 (N_2681,N_2310,N_1920);
or U2682 (N_2682,N_2364,N_2358);
nor U2683 (N_2683,N_1915,N_2066);
or U2684 (N_2684,N_2249,N_1865);
or U2685 (N_2685,N_1728,N_2241);
or U2686 (N_2686,N_2077,N_1684);
or U2687 (N_2687,N_1825,N_1914);
or U2688 (N_2688,N_2242,N_2154);
or U2689 (N_2689,N_2164,N_2198);
or U2690 (N_2690,N_1617,N_2267);
nand U2691 (N_2691,N_1944,N_1901);
nand U2692 (N_2692,N_1836,N_2155);
nor U2693 (N_2693,N_1747,N_2374);
nor U2694 (N_2694,N_2299,N_2377);
or U2695 (N_2695,N_1820,N_1866);
nor U2696 (N_2696,N_2341,N_2319);
or U2697 (N_2697,N_2152,N_2243);
and U2698 (N_2698,N_2075,N_2365);
xnor U2699 (N_2699,N_2206,N_2335);
nand U2700 (N_2700,N_2170,N_1938);
or U2701 (N_2701,N_2034,N_1687);
xnor U2702 (N_2702,N_1613,N_1770);
xnor U2703 (N_2703,N_2073,N_1975);
nand U2704 (N_2704,N_2012,N_2334);
xnor U2705 (N_2705,N_2097,N_2071);
nand U2706 (N_2706,N_1799,N_2150);
xnor U2707 (N_2707,N_1696,N_2177);
and U2708 (N_2708,N_2290,N_1840);
or U2709 (N_2709,N_1884,N_2248);
nand U2710 (N_2710,N_1643,N_2280);
nand U2711 (N_2711,N_1996,N_1690);
nor U2712 (N_2712,N_1843,N_1611);
nor U2713 (N_2713,N_2115,N_2252);
and U2714 (N_2714,N_1620,N_2094);
nor U2715 (N_2715,N_2019,N_2140);
nor U2716 (N_2716,N_2025,N_1646);
or U2717 (N_2717,N_2045,N_1709);
nand U2718 (N_2718,N_2086,N_2084);
or U2719 (N_2719,N_1888,N_1860);
or U2720 (N_2720,N_1871,N_2231);
xnor U2721 (N_2721,N_2212,N_1989);
nor U2722 (N_2722,N_2199,N_2147);
nor U2723 (N_2723,N_2351,N_1835);
nor U2724 (N_2724,N_1886,N_2303);
and U2725 (N_2725,N_2343,N_1876);
xor U2726 (N_2726,N_2014,N_2099);
and U2727 (N_2727,N_1715,N_1622);
xor U2728 (N_2728,N_2210,N_1828);
xnor U2729 (N_2729,N_2111,N_1841);
nand U2730 (N_2730,N_1718,N_1660);
xor U2731 (N_2731,N_1981,N_2284);
xnor U2732 (N_2732,N_2318,N_1774);
or U2733 (N_2733,N_1719,N_2149);
nor U2734 (N_2734,N_2209,N_1961);
and U2735 (N_2735,N_1925,N_2399);
and U2736 (N_2736,N_1868,N_1893);
or U2737 (N_2737,N_2005,N_1630);
nand U2738 (N_2738,N_2229,N_2069);
nor U2739 (N_2739,N_2083,N_2085);
nor U2740 (N_2740,N_2051,N_1862);
nand U2741 (N_2741,N_2350,N_2327);
and U2742 (N_2742,N_1821,N_2213);
nor U2743 (N_2743,N_1675,N_1791);
xnor U2744 (N_2744,N_1673,N_1858);
nor U2745 (N_2745,N_1692,N_1957);
or U2746 (N_2746,N_1706,N_2103);
nand U2747 (N_2747,N_2074,N_2306);
xor U2748 (N_2748,N_1711,N_2328);
and U2749 (N_2749,N_1723,N_1883);
and U2750 (N_2750,N_2128,N_2234);
or U2751 (N_2751,N_1962,N_1922);
nor U2752 (N_2752,N_1940,N_1744);
nor U2753 (N_2753,N_1792,N_1640);
nor U2754 (N_2754,N_1777,N_2089);
or U2755 (N_2755,N_1638,N_2090);
nor U2756 (N_2756,N_1601,N_2015);
or U2757 (N_2757,N_2392,N_2398);
nor U2758 (N_2758,N_1879,N_1963);
xor U2759 (N_2759,N_2261,N_1699);
and U2760 (N_2760,N_1784,N_1994);
xnor U2761 (N_2761,N_1609,N_2317);
or U2762 (N_2762,N_2129,N_1658);
or U2763 (N_2763,N_2391,N_1612);
xor U2764 (N_2764,N_1897,N_1945);
and U2765 (N_2765,N_1918,N_2161);
nor U2766 (N_2766,N_2189,N_2026);
xnor U2767 (N_2767,N_1917,N_2146);
or U2768 (N_2768,N_2049,N_2218);
xor U2769 (N_2769,N_2143,N_1789);
or U2770 (N_2770,N_1869,N_1781);
or U2771 (N_2771,N_2296,N_2308);
nor U2772 (N_2772,N_1993,N_1846);
xor U2773 (N_2773,N_2246,N_1672);
and U2774 (N_2774,N_1864,N_1782);
or U2775 (N_2775,N_2175,N_1907);
nand U2776 (N_2776,N_1631,N_1689);
nand U2777 (N_2777,N_2237,N_2042);
or U2778 (N_2778,N_1653,N_2109);
and U2779 (N_2779,N_1909,N_2004);
xnor U2780 (N_2780,N_2007,N_1983);
xor U2781 (N_2781,N_2148,N_1810);
xnor U2782 (N_2782,N_1776,N_1878);
nor U2783 (N_2783,N_1892,N_2279);
and U2784 (N_2784,N_2061,N_2330);
and U2785 (N_2785,N_2171,N_2311);
and U2786 (N_2786,N_1678,N_1727);
nand U2787 (N_2787,N_2108,N_1906);
nand U2788 (N_2788,N_1877,N_2064);
and U2789 (N_2789,N_1982,N_1749);
and U2790 (N_2790,N_1844,N_1798);
nand U2791 (N_2791,N_1680,N_1758);
and U2792 (N_2792,N_1805,N_2133);
nor U2793 (N_2793,N_1823,N_2113);
or U2794 (N_2794,N_1968,N_2378);
nor U2795 (N_2795,N_1742,N_2291);
nand U2796 (N_2796,N_2250,N_1682);
xnor U2797 (N_2797,N_1895,N_1764);
and U2798 (N_2798,N_1979,N_2021);
nand U2799 (N_2799,N_2185,N_2204);
nor U2800 (N_2800,N_1688,N_2305);
or U2801 (N_2801,N_2302,N_1716);
nand U2802 (N_2802,N_1851,N_1815);
xnor U2803 (N_2803,N_2116,N_1782);
nor U2804 (N_2804,N_1707,N_2330);
and U2805 (N_2805,N_2326,N_1946);
nand U2806 (N_2806,N_1782,N_1619);
or U2807 (N_2807,N_2166,N_2352);
nand U2808 (N_2808,N_1774,N_1697);
nand U2809 (N_2809,N_2145,N_1722);
nor U2810 (N_2810,N_2203,N_2170);
or U2811 (N_2811,N_1749,N_2317);
or U2812 (N_2812,N_1898,N_1952);
nor U2813 (N_2813,N_1834,N_2254);
xor U2814 (N_2814,N_1979,N_2107);
nor U2815 (N_2815,N_1817,N_2081);
nand U2816 (N_2816,N_1971,N_1645);
and U2817 (N_2817,N_2319,N_2295);
nand U2818 (N_2818,N_1620,N_2380);
or U2819 (N_2819,N_1846,N_1787);
xnor U2820 (N_2820,N_2340,N_1850);
and U2821 (N_2821,N_1902,N_2088);
or U2822 (N_2822,N_2333,N_1874);
or U2823 (N_2823,N_1762,N_1949);
nor U2824 (N_2824,N_1710,N_2254);
nand U2825 (N_2825,N_2328,N_1648);
nor U2826 (N_2826,N_2364,N_2391);
nor U2827 (N_2827,N_1645,N_1947);
xor U2828 (N_2828,N_1693,N_1670);
and U2829 (N_2829,N_1954,N_1776);
nand U2830 (N_2830,N_2290,N_2165);
nand U2831 (N_2831,N_1845,N_2216);
nor U2832 (N_2832,N_1817,N_1626);
or U2833 (N_2833,N_1637,N_2309);
xnor U2834 (N_2834,N_2177,N_1991);
xor U2835 (N_2835,N_1757,N_2367);
nand U2836 (N_2836,N_2213,N_2248);
or U2837 (N_2837,N_1833,N_2285);
xnor U2838 (N_2838,N_2006,N_2177);
nor U2839 (N_2839,N_1852,N_1924);
or U2840 (N_2840,N_2301,N_1897);
and U2841 (N_2841,N_1720,N_2383);
nor U2842 (N_2842,N_2316,N_1720);
and U2843 (N_2843,N_1989,N_2121);
and U2844 (N_2844,N_2043,N_1811);
xor U2845 (N_2845,N_2166,N_2016);
and U2846 (N_2846,N_2369,N_1734);
and U2847 (N_2847,N_2270,N_1695);
nand U2848 (N_2848,N_1664,N_1844);
nor U2849 (N_2849,N_1933,N_1699);
xor U2850 (N_2850,N_1632,N_2147);
and U2851 (N_2851,N_1817,N_1925);
and U2852 (N_2852,N_2154,N_1653);
and U2853 (N_2853,N_1667,N_1794);
and U2854 (N_2854,N_2073,N_2175);
nor U2855 (N_2855,N_1935,N_1736);
and U2856 (N_2856,N_1783,N_2209);
or U2857 (N_2857,N_2137,N_2233);
and U2858 (N_2858,N_1975,N_1977);
or U2859 (N_2859,N_1980,N_1643);
xnor U2860 (N_2860,N_1739,N_1633);
nor U2861 (N_2861,N_1653,N_2059);
or U2862 (N_2862,N_2206,N_2281);
nor U2863 (N_2863,N_2001,N_1700);
nand U2864 (N_2864,N_2250,N_1686);
and U2865 (N_2865,N_1979,N_1838);
xnor U2866 (N_2866,N_1821,N_1761);
nand U2867 (N_2867,N_2121,N_1602);
or U2868 (N_2868,N_1996,N_1969);
nor U2869 (N_2869,N_2023,N_1960);
nor U2870 (N_2870,N_1971,N_1782);
or U2871 (N_2871,N_2210,N_2392);
nand U2872 (N_2872,N_2145,N_2090);
nor U2873 (N_2873,N_2287,N_1988);
xor U2874 (N_2874,N_1759,N_1942);
or U2875 (N_2875,N_1846,N_1612);
nand U2876 (N_2876,N_2295,N_1854);
nand U2877 (N_2877,N_1836,N_1705);
xnor U2878 (N_2878,N_1761,N_1980);
or U2879 (N_2879,N_2152,N_2139);
xor U2880 (N_2880,N_1716,N_2341);
or U2881 (N_2881,N_2333,N_1613);
xor U2882 (N_2882,N_1960,N_1666);
nand U2883 (N_2883,N_2248,N_1704);
nor U2884 (N_2884,N_1870,N_2291);
xnor U2885 (N_2885,N_1811,N_2033);
and U2886 (N_2886,N_2306,N_2259);
nor U2887 (N_2887,N_1919,N_1602);
nand U2888 (N_2888,N_1603,N_1693);
or U2889 (N_2889,N_2188,N_1759);
nand U2890 (N_2890,N_1663,N_2009);
xnor U2891 (N_2891,N_1690,N_1751);
nand U2892 (N_2892,N_2099,N_1714);
nor U2893 (N_2893,N_2371,N_2297);
and U2894 (N_2894,N_2353,N_2053);
nand U2895 (N_2895,N_2076,N_2104);
or U2896 (N_2896,N_1988,N_1859);
nor U2897 (N_2897,N_1938,N_1772);
nor U2898 (N_2898,N_2238,N_1624);
nand U2899 (N_2899,N_2297,N_2254);
or U2900 (N_2900,N_1966,N_1989);
nand U2901 (N_2901,N_1692,N_1983);
xor U2902 (N_2902,N_1653,N_1806);
or U2903 (N_2903,N_1707,N_2136);
nand U2904 (N_2904,N_2040,N_1888);
and U2905 (N_2905,N_1881,N_2266);
nor U2906 (N_2906,N_1834,N_1662);
nor U2907 (N_2907,N_1927,N_1658);
or U2908 (N_2908,N_1756,N_2131);
xnor U2909 (N_2909,N_2349,N_1744);
and U2910 (N_2910,N_1748,N_2223);
nand U2911 (N_2911,N_1827,N_2103);
nand U2912 (N_2912,N_1793,N_1761);
and U2913 (N_2913,N_1872,N_1713);
nor U2914 (N_2914,N_1973,N_2157);
nor U2915 (N_2915,N_1640,N_1752);
xnor U2916 (N_2916,N_1967,N_2040);
nor U2917 (N_2917,N_1998,N_2258);
nor U2918 (N_2918,N_2040,N_1815);
or U2919 (N_2919,N_1996,N_2087);
xnor U2920 (N_2920,N_2233,N_1663);
and U2921 (N_2921,N_2295,N_2225);
and U2922 (N_2922,N_2242,N_1699);
or U2923 (N_2923,N_1968,N_1952);
nor U2924 (N_2924,N_2247,N_2177);
nand U2925 (N_2925,N_1718,N_1981);
and U2926 (N_2926,N_1902,N_1908);
and U2927 (N_2927,N_2328,N_1754);
nor U2928 (N_2928,N_2009,N_1637);
nand U2929 (N_2929,N_1866,N_1792);
nor U2930 (N_2930,N_2322,N_1800);
nor U2931 (N_2931,N_1849,N_1688);
or U2932 (N_2932,N_2056,N_1619);
and U2933 (N_2933,N_1821,N_1709);
nand U2934 (N_2934,N_1716,N_2079);
or U2935 (N_2935,N_1885,N_1911);
nor U2936 (N_2936,N_1876,N_2264);
nor U2937 (N_2937,N_2082,N_2076);
and U2938 (N_2938,N_1980,N_2254);
or U2939 (N_2939,N_1765,N_2015);
or U2940 (N_2940,N_1985,N_1699);
nand U2941 (N_2941,N_2324,N_2093);
and U2942 (N_2942,N_1628,N_2244);
nor U2943 (N_2943,N_1938,N_1875);
nand U2944 (N_2944,N_1874,N_2215);
and U2945 (N_2945,N_1925,N_2157);
or U2946 (N_2946,N_1672,N_2235);
nor U2947 (N_2947,N_1864,N_1679);
or U2948 (N_2948,N_2337,N_2211);
or U2949 (N_2949,N_1790,N_1685);
and U2950 (N_2950,N_2372,N_1793);
and U2951 (N_2951,N_2178,N_2311);
nand U2952 (N_2952,N_1825,N_2074);
nand U2953 (N_2953,N_2198,N_2387);
or U2954 (N_2954,N_1864,N_1861);
and U2955 (N_2955,N_1801,N_2102);
xnor U2956 (N_2956,N_2278,N_2330);
nand U2957 (N_2957,N_1926,N_2363);
xor U2958 (N_2958,N_1774,N_1735);
xnor U2959 (N_2959,N_2108,N_1950);
nor U2960 (N_2960,N_2205,N_2147);
and U2961 (N_2961,N_1600,N_1943);
nand U2962 (N_2962,N_1968,N_2106);
xnor U2963 (N_2963,N_2100,N_2032);
and U2964 (N_2964,N_1684,N_2300);
and U2965 (N_2965,N_2139,N_1775);
nor U2966 (N_2966,N_2093,N_2298);
and U2967 (N_2967,N_1630,N_1793);
nor U2968 (N_2968,N_1632,N_2233);
nor U2969 (N_2969,N_2324,N_1693);
or U2970 (N_2970,N_1814,N_2373);
nand U2971 (N_2971,N_2302,N_2268);
and U2972 (N_2972,N_1959,N_2301);
nand U2973 (N_2973,N_2294,N_1864);
nand U2974 (N_2974,N_1637,N_1771);
nor U2975 (N_2975,N_1914,N_2101);
nor U2976 (N_2976,N_2256,N_1971);
or U2977 (N_2977,N_1608,N_2196);
xnor U2978 (N_2978,N_1970,N_2098);
nor U2979 (N_2979,N_2131,N_1972);
or U2980 (N_2980,N_2278,N_1901);
nand U2981 (N_2981,N_1928,N_2206);
nand U2982 (N_2982,N_2011,N_2066);
and U2983 (N_2983,N_2387,N_1732);
nor U2984 (N_2984,N_2215,N_2267);
and U2985 (N_2985,N_2228,N_2114);
and U2986 (N_2986,N_2165,N_1894);
nand U2987 (N_2987,N_2214,N_2121);
or U2988 (N_2988,N_1762,N_1872);
nor U2989 (N_2989,N_2353,N_1719);
and U2990 (N_2990,N_2121,N_2205);
and U2991 (N_2991,N_2390,N_1642);
nor U2992 (N_2992,N_1625,N_1656);
and U2993 (N_2993,N_2375,N_2311);
nor U2994 (N_2994,N_2191,N_2068);
or U2995 (N_2995,N_1990,N_2353);
xnor U2996 (N_2996,N_1662,N_1883);
nor U2997 (N_2997,N_1948,N_2067);
nand U2998 (N_2998,N_2096,N_1899);
nor U2999 (N_2999,N_1622,N_1794);
and U3000 (N_3000,N_2009,N_2068);
nor U3001 (N_3001,N_1892,N_1760);
xor U3002 (N_3002,N_1970,N_2177);
or U3003 (N_3003,N_1933,N_2382);
nor U3004 (N_3004,N_1877,N_1667);
or U3005 (N_3005,N_2008,N_2302);
and U3006 (N_3006,N_1933,N_2082);
or U3007 (N_3007,N_2158,N_1841);
nand U3008 (N_3008,N_2338,N_2184);
and U3009 (N_3009,N_1961,N_1973);
nor U3010 (N_3010,N_1676,N_2014);
xor U3011 (N_3011,N_2256,N_2090);
xor U3012 (N_3012,N_1946,N_2338);
or U3013 (N_3013,N_1981,N_1700);
nand U3014 (N_3014,N_2287,N_1999);
and U3015 (N_3015,N_2362,N_2284);
xnor U3016 (N_3016,N_2255,N_1740);
nand U3017 (N_3017,N_2026,N_1881);
nor U3018 (N_3018,N_1798,N_1977);
nor U3019 (N_3019,N_1967,N_2298);
xnor U3020 (N_3020,N_1920,N_1695);
xnor U3021 (N_3021,N_1811,N_1764);
or U3022 (N_3022,N_2127,N_2245);
or U3023 (N_3023,N_2241,N_2159);
and U3024 (N_3024,N_1753,N_1775);
or U3025 (N_3025,N_1960,N_2306);
and U3026 (N_3026,N_1734,N_2080);
and U3027 (N_3027,N_2299,N_2292);
xnor U3028 (N_3028,N_2040,N_2236);
nand U3029 (N_3029,N_2105,N_1681);
and U3030 (N_3030,N_1631,N_2371);
nand U3031 (N_3031,N_2083,N_2239);
nor U3032 (N_3032,N_1833,N_1758);
and U3033 (N_3033,N_2083,N_1743);
and U3034 (N_3034,N_1723,N_1858);
nor U3035 (N_3035,N_2372,N_2385);
nor U3036 (N_3036,N_2219,N_2124);
or U3037 (N_3037,N_1744,N_1615);
or U3038 (N_3038,N_2154,N_2025);
or U3039 (N_3039,N_2287,N_1692);
xor U3040 (N_3040,N_1728,N_1650);
nand U3041 (N_3041,N_2272,N_2137);
or U3042 (N_3042,N_1982,N_1860);
nor U3043 (N_3043,N_2351,N_2232);
and U3044 (N_3044,N_2158,N_2334);
xnor U3045 (N_3045,N_2069,N_2113);
nand U3046 (N_3046,N_2318,N_1933);
or U3047 (N_3047,N_1904,N_2303);
nand U3048 (N_3048,N_2197,N_1784);
or U3049 (N_3049,N_1825,N_2105);
nand U3050 (N_3050,N_2115,N_2309);
or U3051 (N_3051,N_2186,N_2323);
or U3052 (N_3052,N_1825,N_1788);
or U3053 (N_3053,N_2162,N_2381);
and U3054 (N_3054,N_1634,N_1966);
or U3055 (N_3055,N_2293,N_2339);
xnor U3056 (N_3056,N_1611,N_2259);
nor U3057 (N_3057,N_1652,N_2232);
or U3058 (N_3058,N_1766,N_2209);
and U3059 (N_3059,N_1608,N_1742);
and U3060 (N_3060,N_2236,N_2051);
or U3061 (N_3061,N_2033,N_1827);
nor U3062 (N_3062,N_1802,N_2243);
nand U3063 (N_3063,N_2023,N_2059);
xnor U3064 (N_3064,N_2299,N_2182);
and U3065 (N_3065,N_1831,N_2362);
nand U3066 (N_3066,N_1680,N_2154);
and U3067 (N_3067,N_2237,N_2160);
or U3068 (N_3068,N_1713,N_1976);
nor U3069 (N_3069,N_2019,N_2284);
nor U3070 (N_3070,N_2393,N_2001);
xor U3071 (N_3071,N_2340,N_1616);
nand U3072 (N_3072,N_2259,N_2137);
and U3073 (N_3073,N_1665,N_2302);
nor U3074 (N_3074,N_2357,N_2168);
nand U3075 (N_3075,N_2339,N_1927);
and U3076 (N_3076,N_2366,N_1751);
nand U3077 (N_3077,N_2271,N_2184);
and U3078 (N_3078,N_2127,N_2250);
or U3079 (N_3079,N_1786,N_1608);
and U3080 (N_3080,N_1970,N_1731);
and U3081 (N_3081,N_2095,N_1727);
xnor U3082 (N_3082,N_1845,N_1966);
nand U3083 (N_3083,N_2332,N_2335);
nor U3084 (N_3084,N_1791,N_1703);
nand U3085 (N_3085,N_1672,N_1976);
xor U3086 (N_3086,N_2342,N_2246);
nand U3087 (N_3087,N_1829,N_2023);
or U3088 (N_3088,N_2312,N_1651);
nand U3089 (N_3089,N_1822,N_1791);
or U3090 (N_3090,N_1990,N_2122);
or U3091 (N_3091,N_1809,N_1992);
or U3092 (N_3092,N_1664,N_2170);
nor U3093 (N_3093,N_2194,N_1620);
nand U3094 (N_3094,N_2356,N_2295);
and U3095 (N_3095,N_2076,N_1785);
nor U3096 (N_3096,N_1848,N_1955);
xor U3097 (N_3097,N_2284,N_2077);
and U3098 (N_3098,N_1652,N_1714);
xnor U3099 (N_3099,N_2137,N_1605);
nand U3100 (N_3100,N_2330,N_2313);
and U3101 (N_3101,N_1782,N_2165);
or U3102 (N_3102,N_2024,N_2198);
xor U3103 (N_3103,N_2018,N_2245);
and U3104 (N_3104,N_1846,N_2018);
nand U3105 (N_3105,N_1823,N_1697);
xnor U3106 (N_3106,N_2033,N_2080);
and U3107 (N_3107,N_1813,N_2120);
nor U3108 (N_3108,N_2245,N_1876);
nor U3109 (N_3109,N_2294,N_2241);
nand U3110 (N_3110,N_2032,N_1660);
nand U3111 (N_3111,N_2143,N_2219);
or U3112 (N_3112,N_1681,N_1886);
nor U3113 (N_3113,N_1786,N_2354);
nand U3114 (N_3114,N_1700,N_2322);
or U3115 (N_3115,N_1929,N_2050);
xnor U3116 (N_3116,N_2350,N_2287);
nand U3117 (N_3117,N_2121,N_1747);
and U3118 (N_3118,N_2251,N_2198);
and U3119 (N_3119,N_2251,N_1688);
and U3120 (N_3120,N_1970,N_2218);
nand U3121 (N_3121,N_1924,N_2387);
xor U3122 (N_3122,N_1762,N_1780);
or U3123 (N_3123,N_2130,N_2304);
xnor U3124 (N_3124,N_1893,N_1894);
nand U3125 (N_3125,N_2294,N_1915);
and U3126 (N_3126,N_1952,N_2216);
and U3127 (N_3127,N_1992,N_1610);
nand U3128 (N_3128,N_1614,N_2146);
or U3129 (N_3129,N_2138,N_2301);
nand U3130 (N_3130,N_2278,N_2083);
nor U3131 (N_3131,N_1963,N_1768);
and U3132 (N_3132,N_1883,N_1748);
xnor U3133 (N_3133,N_2248,N_1639);
or U3134 (N_3134,N_1823,N_1943);
or U3135 (N_3135,N_1688,N_1840);
nor U3136 (N_3136,N_1811,N_2115);
and U3137 (N_3137,N_2313,N_2179);
nor U3138 (N_3138,N_2077,N_1930);
or U3139 (N_3139,N_1775,N_1642);
nor U3140 (N_3140,N_1808,N_1769);
nor U3141 (N_3141,N_1651,N_2042);
nor U3142 (N_3142,N_2169,N_1659);
and U3143 (N_3143,N_1742,N_2126);
xnor U3144 (N_3144,N_2315,N_2117);
nor U3145 (N_3145,N_1637,N_1947);
xor U3146 (N_3146,N_2052,N_2034);
nand U3147 (N_3147,N_1919,N_2120);
xnor U3148 (N_3148,N_2081,N_2205);
nor U3149 (N_3149,N_1774,N_2395);
nand U3150 (N_3150,N_1751,N_2389);
nand U3151 (N_3151,N_2083,N_1833);
nand U3152 (N_3152,N_1892,N_2303);
and U3153 (N_3153,N_1868,N_1604);
or U3154 (N_3154,N_2361,N_1827);
and U3155 (N_3155,N_1755,N_1730);
xnor U3156 (N_3156,N_1656,N_2021);
nor U3157 (N_3157,N_2352,N_2384);
nor U3158 (N_3158,N_2015,N_1681);
nand U3159 (N_3159,N_2213,N_2156);
nor U3160 (N_3160,N_1844,N_1675);
or U3161 (N_3161,N_2027,N_1907);
or U3162 (N_3162,N_1882,N_1715);
or U3163 (N_3163,N_1911,N_1716);
and U3164 (N_3164,N_2026,N_1705);
nor U3165 (N_3165,N_1712,N_1756);
and U3166 (N_3166,N_1785,N_1690);
xnor U3167 (N_3167,N_2029,N_1802);
and U3168 (N_3168,N_1755,N_1681);
nor U3169 (N_3169,N_1703,N_1755);
nand U3170 (N_3170,N_1786,N_2015);
nor U3171 (N_3171,N_2263,N_1695);
and U3172 (N_3172,N_2021,N_1708);
xnor U3173 (N_3173,N_1927,N_1714);
nand U3174 (N_3174,N_1965,N_1611);
and U3175 (N_3175,N_2336,N_1717);
xnor U3176 (N_3176,N_1898,N_1691);
or U3177 (N_3177,N_1885,N_1638);
nand U3178 (N_3178,N_1693,N_2313);
nor U3179 (N_3179,N_1692,N_1607);
nor U3180 (N_3180,N_1726,N_1866);
nand U3181 (N_3181,N_2168,N_2291);
nor U3182 (N_3182,N_1776,N_1705);
nand U3183 (N_3183,N_1806,N_2322);
nor U3184 (N_3184,N_1625,N_2236);
and U3185 (N_3185,N_2111,N_1980);
xor U3186 (N_3186,N_2286,N_2252);
xnor U3187 (N_3187,N_1999,N_2340);
or U3188 (N_3188,N_2339,N_1605);
nor U3189 (N_3189,N_1784,N_1799);
xor U3190 (N_3190,N_2204,N_1995);
or U3191 (N_3191,N_2386,N_2141);
nand U3192 (N_3192,N_1844,N_2186);
and U3193 (N_3193,N_2243,N_1764);
and U3194 (N_3194,N_1901,N_2232);
xor U3195 (N_3195,N_1947,N_1821);
nor U3196 (N_3196,N_2089,N_1760);
and U3197 (N_3197,N_2219,N_1787);
nor U3198 (N_3198,N_1644,N_2286);
xnor U3199 (N_3199,N_2076,N_2157);
nor U3200 (N_3200,N_3038,N_2941);
and U3201 (N_3201,N_3006,N_2903);
nand U3202 (N_3202,N_2747,N_3167);
xor U3203 (N_3203,N_3021,N_3134);
nand U3204 (N_3204,N_2987,N_2957);
and U3205 (N_3205,N_2897,N_2539);
and U3206 (N_3206,N_3194,N_2924);
and U3207 (N_3207,N_2898,N_2517);
nor U3208 (N_3208,N_3061,N_2908);
and U3209 (N_3209,N_3102,N_2852);
nor U3210 (N_3210,N_2600,N_2454);
or U3211 (N_3211,N_3059,N_3029);
nand U3212 (N_3212,N_2889,N_2739);
xor U3213 (N_3213,N_2563,N_2905);
and U3214 (N_3214,N_3013,N_2726);
nand U3215 (N_3215,N_2416,N_2942);
nand U3216 (N_3216,N_3025,N_3090);
nand U3217 (N_3217,N_2583,N_3123);
nor U3218 (N_3218,N_2459,N_3072);
xor U3219 (N_3219,N_2945,N_3108);
nand U3220 (N_3220,N_2627,N_2564);
nor U3221 (N_3221,N_2493,N_2749);
xnor U3222 (N_3222,N_2460,N_2642);
nand U3223 (N_3223,N_3015,N_2954);
and U3224 (N_3224,N_2814,N_2592);
nor U3225 (N_3225,N_2746,N_2877);
nor U3226 (N_3226,N_2405,N_3149);
nor U3227 (N_3227,N_2951,N_2891);
and U3228 (N_3228,N_2571,N_2439);
or U3229 (N_3229,N_2588,N_3164);
nand U3230 (N_3230,N_2499,N_2964);
or U3231 (N_3231,N_3126,N_3054);
nor U3232 (N_3232,N_2411,N_2615);
and U3233 (N_3233,N_2607,N_2773);
xnor U3234 (N_3234,N_2569,N_2855);
nand U3235 (N_3235,N_2829,N_2846);
or U3236 (N_3236,N_2516,N_2966);
nand U3237 (N_3237,N_2890,N_2839);
and U3238 (N_3238,N_2755,N_2408);
or U3239 (N_3239,N_2512,N_2502);
nor U3240 (N_3240,N_2614,N_3027);
nor U3241 (N_3241,N_2520,N_2778);
xnor U3242 (N_3242,N_3098,N_2689);
and U3243 (N_3243,N_3182,N_2929);
nor U3244 (N_3244,N_2596,N_2425);
or U3245 (N_3245,N_2716,N_2663);
nor U3246 (N_3246,N_3136,N_2494);
nor U3247 (N_3247,N_2878,N_2617);
xor U3248 (N_3248,N_2863,N_2522);
xor U3249 (N_3249,N_2496,N_2559);
or U3250 (N_3250,N_2692,N_2697);
or U3251 (N_3251,N_3100,N_3103);
nor U3252 (N_3252,N_2787,N_2529);
xnor U3253 (N_3253,N_2651,N_2955);
nor U3254 (N_3254,N_2703,N_2501);
and U3255 (N_3255,N_3160,N_3191);
and U3256 (N_3256,N_2680,N_2526);
or U3257 (N_3257,N_2906,N_2751);
and U3258 (N_3258,N_3095,N_2476);
xnor U3259 (N_3259,N_2543,N_3002);
and U3260 (N_3260,N_3060,N_2561);
nor U3261 (N_3261,N_2469,N_2487);
and U3262 (N_3262,N_2448,N_2506);
nor U3263 (N_3263,N_2622,N_2928);
nor U3264 (N_3264,N_2546,N_3141);
nor U3265 (N_3265,N_3030,N_2871);
or U3266 (N_3266,N_2545,N_2734);
nor U3267 (N_3267,N_2780,N_2503);
and U3268 (N_3268,N_2407,N_2925);
nor U3269 (N_3269,N_2451,N_2758);
or U3270 (N_3270,N_3009,N_2597);
or U3271 (N_3271,N_2582,N_2834);
nor U3272 (N_3272,N_2444,N_2712);
xor U3273 (N_3273,N_2748,N_3058);
nand U3274 (N_3274,N_2631,N_2585);
nand U3275 (N_3275,N_2532,N_2720);
xor U3276 (N_3276,N_2616,N_2800);
nor U3277 (N_3277,N_2518,N_3169);
xnor U3278 (N_3278,N_2899,N_2489);
nand U3279 (N_3279,N_2468,N_2847);
nor U3280 (N_3280,N_2511,N_2844);
and U3281 (N_3281,N_2472,N_2687);
nor U3282 (N_3282,N_2798,N_2817);
or U3283 (N_3283,N_2523,N_2541);
and U3284 (N_3284,N_2816,N_2785);
or U3285 (N_3285,N_2854,N_3173);
and U3286 (N_3286,N_2648,N_2760);
nor U3287 (N_3287,N_2686,N_2804);
or U3288 (N_3288,N_2790,N_2887);
and U3289 (N_3289,N_2827,N_2638);
or U3290 (N_3290,N_2447,N_2477);
or U3291 (N_3291,N_3017,N_3119);
and U3292 (N_3292,N_3028,N_3171);
and U3293 (N_3293,N_3089,N_2603);
and U3294 (N_3294,N_2473,N_2996);
xor U3295 (N_3295,N_2811,N_2693);
xnor U3296 (N_3296,N_2431,N_2741);
nor U3297 (N_3297,N_2437,N_2728);
nor U3298 (N_3298,N_2786,N_2880);
nand U3299 (N_3299,N_2730,N_2450);
xor U3300 (N_3300,N_2762,N_3032);
and U3301 (N_3301,N_2885,N_2842);
and U3302 (N_3302,N_2462,N_2576);
nor U3303 (N_3303,N_2930,N_2590);
nor U3304 (N_3304,N_2649,N_2401);
and U3305 (N_3305,N_2536,N_2981);
nand U3306 (N_3306,N_2990,N_3178);
xor U3307 (N_3307,N_2409,N_3037);
or U3308 (N_3308,N_3196,N_3165);
or U3309 (N_3309,N_2774,N_2997);
nor U3310 (N_3310,N_2655,N_2574);
xor U3311 (N_3311,N_3082,N_2659);
or U3312 (N_3312,N_2573,N_2643);
xnor U3313 (N_3313,N_3073,N_3185);
nand U3314 (N_3314,N_2848,N_3065);
nor U3315 (N_3315,N_2915,N_2534);
xor U3316 (N_3316,N_3024,N_2613);
or U3317 (N_3317,N_2736,N_3135);
nor U3318 (N_3318,N_2772,N_2538);
xnor U3319 (N_3319,N_2552,N_2791);
or U3320 (N_3320,N_2436,N_3106);
or U3321 (N_3321,N_2861,N_2510);
nor U3322 (N_3322,N_2952,N_2604);
xnor U3323 (N_3323,N_2420,N_2808);
or U3324 (N_3324,N_3138,N_3057);
nor U3325 (N_3325,N_3071,N_2701);
and U3326 (N_3326,N_2630,N_2490);
or U3327 (N_3327,N_2806,N_2868);
and U3328 (N_3328,N_3117,N_2652);
xor U3329 (N_3329,N_2531,N_2828);
nor U3330 (N_3330,N_2919,N_3174);
nand U3331 (N_3331,N_2535,N_2418);
nand U3332 (N_3332,N_3133,N_2892);
nand U3333 (N_3333,N_2667,N_2986);
and U3334 (N_3334,N_2644,N_2833);
nor U3335 (N_3335,N_2479,N_2722);
nand U3336 (N_3336,N_2896,N_2429);
or U3337 (N_3337,N_2938,N_2883);
or U3338 (N_3338,N_2738,N_3018);
and U3339 (N_3339,N_2637,N_2918);
xnor U3340 (N_3340,N_2632,N_2611);
nor U3341 (N_3341,N_3120,N_2936);
xor U3342 (N_3342,N_3070,N_2881);
xor U3343 (N_3343,N_2442,N_2540);
or U3344 (N_3344,N_2795,N_2403);
nand U3345 (N_3345,N_3150,N_2624);
nor U3346 (N_3346,N_2402,N_2700);
xor U3347 (N_3347,N_2732,N_3074);
or U3348 (N_3348,N_2645,N_2524);
and U3349 (N_3349,N_3139,N_2481);
nand U3350 (N_3350,N_3033,N_2963);
and U3351 (N_3351,N_2708,N_2423);
nor U3352 (N_3352,N_3069,N_2620);
or U3353 (N_3353,N_2554,N_2713);
or U3354 (N_3354,N_2756,N_2681);
nor U3355 (N_3355,N_2587,N_2544);
or U3356 (N_3356,N_2969,N_3016);
or U3357 (N_3357,N_2933,N_3066);
nand U3358 (N_3358,N_3091,N_2830);
xor U3359 (N_3359,N_2799,N_2464);
or U3360 (N_3360,N_2625,N_2836);
and U3361 (N_3361,N_2610,N_2654);
and U3362 (N_3362,N_2685,N_3068);
or U3363 (N_3363,N_2984,N_3156);
xor U3364 (N_3364,N_2873,N_2949);
nor U3365 (N_3365,N_2907,N_3044);
nand U3366 (N_3366,N_2639,N_2400);
or U3367 (N_3367,N_2406,N_2466);
xnor U3368 (N_3368,N_2428,N_2609);
nand U3369 (N_3369,N_3170,N_3081);
nor U3370 (N_3370,N_2542,N_2968);
nand U3371 (N_3371,N_2983,N_2792);
and U3372 (N_3372,N_2943,N_2788);
nor U3373 (N_3373,N_2683,N_3092);
nor U3374 (N_3374,N_2505,N_2482);
xnor U3375 (N_3375,N_2882,N_2452);
nand U3376 (N_3376,N_2463,N_2671);
xnor U3377 (N_3377,N_3148,N_2684);
nor U3378 (N_3378,N_2467,N_3198);
xor U3379 (N_3379,N_2940,N_2864);
nor U3380 (N_3380,N_2677,N_2803);
or U3381 (N_3381,N_2674,N_2551);
xnor U3382 (N_3382,N_2641,N_2724);
nor U3383 (N_3383,N_2434,N_2740);
nand U3384 (N_3384,N_2455,N_2975);
or U3385 (N_3385,N_2737,N_3043);
xor U3386 (N_3386,N_2706,N_2618);
or U3387 (N_3387,N_2521,N_2950);
nand U3388 (N_3388,N_2553,N_3007);
nor U3389 (N_3389,N_2427,N_2558);
and U3390 (N_3390,N_2865,N_2488);
nand U3391 (N_3391,N_2783,N_3166);
nand U3392 (N_3392,N_2937,N_2805);
xor U3393 (N_3393,N_2676,N_2960);
xnor U3394 (N_3394,N_2858,N_2438);
or U3395 (N_3395,N_2498,N_2628);
nor U3396 (N_3396,N_3062,N_2660);
and U3397 (N_3397,N_2824,N_2843);
and U3398 (N_3398,N_2530,N_3175);
nand U3399 (N_3399,N_2812,N_2884);
xnor U3400 (N_3400,N_2784,N_3010);
nor U3401 (N_3401,N_2599,N_2761);
nand U3402 (N_3402,N_2766,N_3187);
xor U3403 (N_3403,N_2764,N_2876);
nand U3404 (N_3404,N_3104,N_3154);
xor U3405 (N_3405,N_2931,N_3051);
nand U3406 (N_3406,N_2417,N_3112);
or U3407 (N_3407,N_2446,N_2965);
or U3408 (N_3408,N_2633,N_2958);
and U3409 (N_3409,N_2533,N_2980);
or U3410 (N_3410,N_2895,N_3083);
and U3411 (N_3411,N_2959,N_2572);
xnor U3412 (N_3412,N_2935,N_2888);
and U3413 (N_3413,N_3161,N_2822);
xnor U3414 (N_3414,N_2796,N_2557);
and U3415 (N_3415,N_3000,N_2714);
xnor U3416 (N_3416,N_2991,N_2840);
and U3417 (N_3417,N_2695,N_3153);
and U3418 (N_3418,N_3195,N_3008);
and U3419 (N_3419,N_2721,N_3183);
nor U3420 (N_3420,N_2995,N_2579);
or U3421 (N_3421,N_3144,N_2461);
nand U3422 (N_3422,N_3003,N_3023);
or U3423 (N_3423,N_2497,N_2456);
nand U3424 (N_3424,N_3087,N_3036);
or U3425 (N_3425,N_3050,N_2668);
or U3426 (N_3426,N_3053,N_3022);
xnor U3427 (N_3427,N_3049,N_2771);
or U3428 (N_3428,N_2912,N_2675);
and U3429 (N_3429,N_3125,N_3132);
nand U3430 (N_3430,N_2527,N_2879);
nor U3431 (N_3431,N_2753,N_2850);
nand U3432 (N_3432,N_2670,N_2775);
nand U3433 (N_3433,N_3181,N_2484);
nor U3434 (N_3434,N_2718,N_3162);
xor U3435 (N_3435,N_2470,N_2849);
or U3436 (N_3436,N_2989,N_2626);
nor U3437 (N_3437,N_2691,N_2415);
or U3438 (N_3438,N_3158,N_3197);
xor U3439 (N_3439,N_3146,N_2922);
nand U3440 (N_3440,N_2742,N_2927);
xnor U3441 (N_3441,N_2653,N_2458);
nor U3442 (N_3442,N_2856,N_2443);
nand U3443 (N_3443,N_2977,N_3085);
xnor U3444 (N_3444,N_2513,N_2900);
and U3445 (N_3445,N_2673,N_3177);
or U3446 (N_3446,N_3041,N_2913);
and U3447 (N_3447,N_2821,N_2519);
or U3448 (N_3448,N_2661,N_2646);
and U3449 (N_3449,N_2413,N_2802);
and U3450 (N_3450,N_2664,N_2979);
and U3451 (N_3451,N_2733,N_2514);
nor U3452 (N_3452,N_2507,N_2421);
nor U3453 (N_3453,N_3113,N_3193);
nand U3454 (N_3454,N_3101,N_2723);
or U3455 (N_3455,N_2548,N_2910);
and U3456 (N_3456,N_3151,N_3042);
and U3457 (N_3457,N_2710,N_2662);
nand U3458 (N_3458,N_3048,N_2682);
nand U3459 (N_3459,N_3142,N_3145);
nor U3460 (N_3460,N_2635,N_2765);
xor U3461 (N_3461,N_2727,N_2962);
nor U3462 (N_3462,N_2605,N_2602);
nor U3463 (N_3463,N_2801,N_3111);
and U3464 (N_3464,N_2867,N_2698);
nor U3465 (N_3465,N_2433,N_2743);
nand U3466 (N_3466,N_3047,N_2825);
or U3467 (N_3467,N_2449,N_2819);
or U3468 (N_3468,N_2593,N_2650);
or U3469 (N_3469,N_2715,N_3067);
xor U3470 (N_3470,N_3011,N_2426);
and U3471 (N_3471,N_2870,N_2575);
or U3472 (N_3472,N_2595,N_2601);
nand U3473 (N_3473,N_2580,N_3046);
or U3474 (N_3474,N_2537,N_2767);
nand U3475 (N_3475,N_2647,N_2636);
xnor U3476 (N_3476,N_2789,N_2939);
and U3477 (N_3477,N_3004,N_2424);
and U3478 (N_3478,N_2699,N_2901);
nand U3479 (N_3479,N_2750,N_2862);
xor U3480 (N_3480,N_2577,N_3115);
xor U3481 (N_3481,N_2591,N_2992);
nand U3482 (N_3482,N_2744,N_2948);
nor U3483 (N_3483,N_2550,N_2809);
and U3484 (N_3484,N_2731,N_2866);
or U3485 (N_3485,N_3076,N_2893);
xor U3486 (N_3486,N_3129,N_2956);
nor U3487 (N_3487,N_2475,N_2944);
and U3488 (N_3488,N_3118,N_2665);
or U3489 (N_3489,N_3105,N_2904);
or U3490 (N_3490,N_2404,N_3168);
and U3491 (N_3491,N_3099,N_2886);
and U3492 (N_3492,N_2999,N_2634);
or U3493 (N_3493,N_2859,N_3163);
nor U3494 (N_3494,N_2457,N_2953);
or U3495 (N_3495,N_2770,N_2422);
or U3496 (N_3496,N_2471,N_3020);
or U3497 (N_3497,N_2666,N_3189);
nor U3498 (N_3498,N_2619,N_2832);
and U3499 (N_3499,N_3188,N_2797);
and U3500 (N_3500,N_3130,N_2973);
xor U3501 (N_3501,N_2946,N_3140);
xnor U3502 (N_3502,N_3184,N_2920);
nor U3503 (N_3503,N_2810,N_2669);
xnor U3504 (N_3504,N_2492,N_2894);
or U3505 (N_3505,N_2976,N_2853);
nor U3506 (N_3506,N_3116,N_2932);
or U3507 (N_3507,N_2719,N_3172);
nand U3508 (N_3508,N_2947,N_3186);
nand U3509 (N_3509,N_2911,N_2508);
and U3510 (N_3510,N_2412,N_2562);
xor U3511 (N_3511,N_2807,N_2782);
and U3512 (N_3512,N_3026,N_2581);
nor U3513 (N_3513,N_2820,N_2629);
nor U3514 (N_3514,N_3155,N_2851);
or U3515 (N_3515,N_2690,N_2769);
and U3516 (N_3516,N_2586,N_2921);
or U3517 (N_3517,N_2656,N_3107);
nor U3518 (N_3518,N_2725,N_2515);
nand U3519 (N_3519,N_3179,N_2860);
and U3520 (N_3520,N_2917,N_2974);
xnor U3521 (N_3521,N_3121,N_2967);
xor U3522 (N_3522,N_2566,N_2547);
nor U3523 (N_3523,N_3056,N_3143);
nand U3524 (N_3524,N_2757,N_2776);
or U3525 (N_3525,N_2465,N_2621);
or U3526 (N_3526,N_3124,N_2478);
nand U3527 (N_3527,N_3110,N_3128);
nand U3528 (N_3528,N_3080,N_2598);
or U3529 (N_3529,N_3034,N_2768);
nor U3530 (N_3530,N_2994,N_2556);
nor U3531 (N_3531,N_3094,N_2694);
or U3532 (N_3532,N_2831,N_2500);
or U3533 (N_3533,N_2432,N_2754);
or U3534 (N_3534,N_3176,N_2678);
nand U3535 (N_3535,N_2838,N_2752);
or U3536 (N_3536,N_2779,N_3147);
nor U3537 (N_3537,N_2875,N_2971);
nand U3538 (N_3538,N_3109,N_2679);
nand U3539 (N_3539,N_3199,N_2504);
nor U3540 (N_3540,N_2549,N_2410);
and U3541 (N_3541,N_3159,N_3031);
or U3542 (N_3542,N_3064,N_3093);
nor U3543 (N_3543,N_2658,N_2440);
nand U3544 (N_3544,N_2435,N_3097);
nor U3545 (N_3545,N_2528,N_2525);
or U3546 (N_3546,N_2486,N_2709);
nand U3547 (N_3547,N_2837,N_3052);
nand U3548 (N_3548,N_2640,N_2688);
and U3549 (N_3549,N_2578,N_2777);
xor U3550 (N_3550,N_3019,N_2480);
and U3551 (N_3551,N_2793,N_3001);
and U3552 (N_3552,N_2606,N_3035);
or U3553 (N_3553,N_2491,N_2560);
nand U3554 (N_3554,N_2453,N_3014);
nand U3555 (N_3555,N_2985,N_2993);
or U3556 (N_3556,N_3063,N_2735);
xor U3557 (N_3557,N_2509,N_2794);
nand U3558 (N_3558,N_3137,N_2608);
nor U3559 (N_3559,N_2841,N_2555);
nand U3560 (N_3560,N_3086,N_2565);
nand U3561 (N_3561,N_2570,N_2926);
nor U3562 (N_3562,N_3045,N_3114);
xnor U3563 (N_3563,N_2916,N_2414);
nor U3564 (N_3564,N_2845,N_3096);
nand U3565 (N_3565,N_2445,N_2909);
or U3566 (N_3566,N_2902,N_2568);
and U3567 (N_3567,N_2872,N_2923);
or U3568 (N_3568,N_2914,N_2982);
nor U3569 (N_3569,N_2826,N_2474);
and U3570 (N_3570,N_2934,N_2623);
nor U3571 (N_3571,N_2869,N_2781);
and U3572 (N_3572,N_3078,N_2857);
or U3573 (N_3573,N_3122,N_2978);
and U3574 (N_3574,N_3075,N_3180);
or U3575 (N_3575,N_2589,N_2813);
xnor U3576 (N_3576,N_3190,N_3039);
and U3577 (N_3577,N_2729,N_2961);
xnor U3578 (N_3578,N_2419,N_2823);
xor U3579 (N_3579,N_3077,N_3152);
nor U3580 (N_3580,N_2988,N_2696);
xnor U3581 (N_3581,N_2998,N_2485);
nand U3582 (N_3582,N_2835,N_3005);
or U3583 (N_3583,N_2430,N_2705);
nand U3584 (N_3584,N_2970,N_2717);
or U3585 (N_3585,N_3040,N_2759);
or U3586 (N_3586,N_3088,N_3055);
nor U3587 (N_3587,N_2483,N_2704);
nand U3588 (N_3588,N_2815,N_2672);
nor U3589 (N_3589,N_2745,N_3192);
nor U3590 (N_3590,N_2495,N_3127);
or U3591 (N_3591,N_2818,N_2972);
nor U3592 (N_3592,N_2657,N_3084);
nand U3593 (N_3593,N_2567,N_3157);
or U3594 (N_3594,N_2584,N_2711);
xor U3595 (N_3595,N_2441,N_2707);
and U3596 (N_3596,N_3079,N_2702);
xor U3597 (N_3597,N_2874,N_2594);
xor U3598 (N_3598,N_2612,N_2763);
and U3599 (N_3599,N_3012,N_3131);
and U3600 (N_3600,N_2897,N_3138);
or U3601 (N_3601,N_2592,N_2635);
xnor U3602 (N_3602,N_2984,N_2967);
and U3603 (N_3603,N_3065,N_2688);
nor U3604 (N_3604,N_2634,N_2621);
nor U3605 (N_3605,N_2402,N_2505);
nand U3606 (N_3606,N_2648,N_3078);
or U3607 (N_3607,N_2573,N_2786);
nor U3608 (N_3608,N_2508,N_3004);
xor U3609 (N_3609,N_2430,N_2483);
xor U3610 (N_3610,N_2937,N_2492);
and U3611 (N_3611,N_2495,N_2552);
xor U3612 (N_3612,N_3088,N_2524);
or U3613 (N_3613,N_2545,N_2696);
or U3614 (N_3614,N_2896,N_2643);
nor U3615 (N_3615,N_2520,N_2449);
and U3616 (N_3616,N_3135,N_2834);
nand U3617 (N_3617,N_2861,N_3102);
and U3618 (N_3618,N_2492,N_2778);
xor U3619 (N_3619,N_2914,N_3029);
nand U3620 (N_3620,N_3196,N_3008);
or U3621 (N_3621,N_2615,N_2744);
xnor U3622 (N_3622,N_2863,N_3121);
nand U3623 (N_3623,N_2849,N_2630);
xor U3624 (N_3624,N_2582,N_3180);
or U3625 (N_3625,N_2745,N_2880);
or U3626 (N_3626,N_2775,N_3144);
nor U3627 (N_3627,N_2448,N_3000);
xnor U3628 (N_3628,N_2852,N_2580);
xnor U3629 (N_3629,N_3073,N_3099);
and U3630 (N_3630,N_2553,N_2998);
xor U3631 (N_3631,N_2706,N_2467);
xor U3632 (N_3632,N_2457,N_3170);
nand U3633 (N_3633,N_2874,N_2743);
or U3634 (N_3634,N_2734,N_2416);
or U3635 (N_3635,N_2894,N_2639);
nand U3636 (N_3636,N_3023,N_2879);
xor U3637 (N_3637,N_2507,N_3047);
nand U3638 (N_3638,N_3091,N_3055);
nor U3639 (N_3639,N_2410,N_2879);
nand U3640 (N_3640,N_2793,N_3185);
and U3641 (N_3641,N_2853,N_2753);
nand U3642 (N_3642,N_2747,N_2719);
and U3643 (N_3643,N_2906,N_3066);
and U3644 (N_3644,N_2680,N_2624);
and U3645 (N_3645,N_2409,N_2934);
xnor U3646 (N_3646,N_3114,N_3095);
or U3647 (N_3647,N_2530,N_3038);
xor U3648 (N_3648,N_2414,N_2586);
xnor U3649 (N_3649,N_2472,N_2673);
nor U3650 (N_3650,N_2780,N_3109);
nor U3651 (N_3651,N_2708,N_2642);
nor U3652 (N_3652,N_3092,N_2771);
nor U3653 (N_3653,N_3108,N_2832);
xnor U3654 (N_3654,N_2428,N_2722);
nor U3655 (N_3655,N_2905,N_2478);
nand U3656 (N_3656,N_2754,N_2791);
xor U3657 (N_3657,N_2954,N_2868);
and U3658 (N_3658,N_2534,N_2586);
xor U3659 (N_3659,N_2683,N_3180);
nand U3660 (N_3660,N_2615,N_3020);
xnor U3661 (N_3661,N_2628,N_2751);
or U3662 (N_3662,N_2841,N_2478);
and U3663 (N_3663,N_3027,N_2514);
and U3664 (N_3664,N_2421,N_2731);
nor U3665 (N_3665,N_2607,N_2524);
nor U3666 (N_3666,N_2955,N_2705);
nor U3667 (N_3667,N_2565,N_2645);
and U3668 (N_3668,N_3053,N_2704);
nor U3669 (N_3669,N_2657,N_2996);
nand U3670 (N_3670,N_2997,N_2508);
and U3671 (N_3671,N_2633,N_2409);
nand U3672 (N_3672,N_2510,N_2555);
xor U3673 (N_3673,N_3172,N_2921);
and U3674 (N_3674,N_2777,N_2749);
nand U3675 (N_3675,N_2804,N_3089);
nand U3676 (N_3676,N_2610,N_2899);
xnor U3677 (N_3677,N_2657,N_2753);
nand U3678 (N_3678,N_2898,N_2797);
or U3679 (N_3679,N_2430,N_2520);
and U3680 (N_3680,N_2724,N_2751);
xnor U3681 (N_3681,N_2506,N_2802);
xor U3682 (N_3682,N_2906,N_2464);
xor U3683 (N_3683,N_3121,N_3015);
nand U3684 (N_3684,N_3031,N_2541);
or U3685 (N_3685,N_2767,N_3037);
and U3686 (N_3686,N_2425,N_2443);
or U3687 (N_3687,N_2894,N_2948);
and U3688 (N_3688,N_2877,N_3098);
nand U3689 (N_3689,N_2621,N_3110);
or U3690 (N_3690,N_3072,N_2892);
xnor U3691 (N_3691,N_2671,N_2750);
or U3692 (N_3692,N_2969,N_2673);
or U3693 (N_3693,N_2710,N_3165);
nor U3694 (N_3694,N_2632,N_2844);
nand U3695 (N_3695,N_2548,N_2885);
xor U3696 (N_3696,N_2507,N_2494);
nand U3697 (N_3697,N_2452,N_2990);
and U3698 (N_3698,N_2740,N_2634);
and U3699 (N_3699,N_3188,N_3033);
and U3700 (N_3700,N_3096,N_3092);
and U3701 (N_3701,N_3155,N_2770);
nand U3702 (N_3702,N_2741,N_2480);
nand U3703 (N_3703,N_2437,N_3110);
nand U3704 (N_3704,N_2995,N_3106);
xor U3705 (N_3705,N_2674,N_3021);
nor U3706 (N_3706,N_3087,N_3022);
xor U3707 (N_3707,N_2441,N_2805);
nor U3708 (N_3708,N_2621,N_2832);
xnor U3709 (N_3709,N_2575,N_2840);
xnor U3710 (N_3710,N_2926,N_2795);
and U3711 (N_3711,N_3178,N_2866);
nand U3712 (N_3712,N_3075,N_2510);
nor U3713 (N_3713,N_3112,N_3021);
xor U3714 (N_3714,N_2485,N_2559);
nor U3715 (N_3715,N_2525,N_3199);
nand U3716 (N_3716,N_2633,N_2477);
nor U3717 (N_3717,N_2577,N_2816);
xor U3718 (N_3718,N_2832,N_2578);
and U3719 (N_3719,N_2527,N_3034);
xor U3720 (N_3720,N_2517,N_2490);
nor U3721 (N_3721,N_2628,N_2806);
nor U3722 (N_3722,N_2446,N_2402);
and U3723 (N_3723,N_2762,N_2831);
or U3724 (N_3724,N_2778,N_3163);
and U3725 (N_3725,N_3107,N_2606);
nor U3726 (N_3726,N_2567,N_2482);
xor U3727 (N_3727,N_2902,N_2599);
nor U3728 (N_3728,N_2894,N_3157);
or U3729 (N_3729,N_2466,N_2892);
nor U3730 (N_3730,N_2606,N_2795);
and U3731 (N_3731,N_2879,N_3009);
and U3732 (N_3732,N_2975,N_2765);
nand U3733 (N_3733,N_2942,N_2787);
xnor U3734 (N_3734,N_2550,N_3120);
xor U3735 (N_3735,N_2867,N_2646);
nand U3736 (N_3736,N_2560,N_2837);
or U3737 (N_3737,N_2740,N_2478);
nor U3738 (N_3738,N_2515,N_3177);
or U3739 (N_3739,N_2504,N_2859);
or U3740 (N_3740,N_3116,N_3186);
or U3741 (N_3741,N_2606,N_2514);
and U3742 (N_3742,N_3108,N_2861);
and U3743 (N_3743,N_2724,N_2849);
or U3744 (N_3744,N_2538,N_2475);
or U3745 (N_3745,N_2916,N_2457);
nor U3746 (N_3746,N_2930,N_2597);
xor U3747 (N_3747,N_3013,N_2812);
nand U3748 (N_3748,N_3136,N_2436);
or U3749 (N_3749,N_2576,N_2657);
or U3750 (N_3750,N_2945,N_3071);
and U3751 (N_3751,N_2834,N_2496);
and U3752 (N_3752,N_3128,N_2567);
xor U3753 (N_3753,N_3024,N_2952);
nand U3754 (N_3754,N_2868,N_2982);
xor U3755 (N_3755,N_2575,N_3154);
nor U3756 (N_3756,N_2463,N_2789);
nand U3757 (N_3757,N_2569,N_2705);
and U3758 (N_3758,N_2840,N_3024);
and U3759 (N_3759,N_3146,N_2916);
nor U3760 (N_3760,N_2991,N_2855);
xor U3761 (N_3761,N_3052,N_2475);
and U3762 (N_3762,N_2850,N_2811);
or U3763 (N_3763,N_2424,N_3056);
xnor U3764 (N_3764,N_2563,N_2593);
or U3765 (N_3765,N_2552,N_3000);
xor U3766 (N_3766,N_2672,N_2936);
or U3767 (N_3767,N_2471,N_3105);
or U3768 (N_3768,N_2676,N_2436);
or U3769 (N_3769,N_2800,N_2860);
and U3770 (N_3770,N_3183,N_2479);
nor U3771 (N_3771,N_2723,N_2891);
xor U3772 (N_3772,N_3060,N_2487);
xnor U3773 (N_3773,N_2805,N_2627);
xor U3774 (N_3774,N_2956,N_2771);
nand U3775 (N_3775,N_2614,N_2490);
nand U3776 (N_3776,N_2584,N_2590);
and U3777 (N_3777,N_2442,N_3191);
and U3778 (N_3778,N_3199,N_2918);
nor U3779 (N_3779,N_3125,N_2894);
nor U3780 (N_3780,N_2450,N_2922);
or U3781 (N_3781,N_2776,N_3073);
and U3782 (N_3782,N_2469,N_2968);
xor U3783 (N_3783,N_2994,N_2783);
xor U3784 (N_3784,N_2595,N_2514);
xor U3785 (N_3785,N_2967,N_2875);
xor U3786 (N_3786,N_2496,N_3088);
nand U3787 (N_3787,N_3148,N_2977);
nand U3788 (N_3788,N_2981,N_3051);
xnor U3789 (N_3789,N_2413,N_2570);
nand U3790 (N_3790,N_2641,N_2979);
nor U3791 (N_3791,N_2873,N_2721);
nor U3792 (N_3792,N_2711,N_2463);
or U3793 (N_3793,N_3009,N_2747);
and U3794 (N_3794,N_2958,N_2663);
and U3795 (N_3795,N_3044,N_3169);
and U3796 (N_3796,N_2636,N_2761);
nand U3797 (N_3797,N_3085,N_3099);
nor U3798 (N_3798,N_2727,N_2504);
xnor U3799 (N_3799,N_2852,N_3127);
or U3800 (N_3800,N_2747,N_2715);
and U3801 (N_3801,N_2952,N_2711);
nand U3802 (N_3802,N_2924,N_3185);
nor U3803 (N_3803,N_3198,N_2583);
nor U3804 (N_3804,N_2920,N_2668);
nor U3805 (N_3805,N_3130,N_3041);
nor U3806 (N_3806,N_2971,N_2665);
and U3807 (N_3807,N_2932,N_3028);
nand U3808 (N_3808,N_2880,N_3006);
or U3809 (N_3809,N_2993,N_2964);
nor U3810 (N_3810,N_2697,N_3077);
xor U3811 (N_3811,N_2688,N_3136);
and U3812 (N_3812,N_3023,N_2597);
or U3813 (N_3813,N_3133,N_2447);
nor U3814 (N_3814,N_2696,N_2882);
and U3815 (N_3815,N_2646,N_2464);
xnor U3816 (N_3816,N_2689,N_2474);
xor U3817 (N_3817,N_2705,N_2693);
xnor U3818 (N_3818,N_3153,N_2473);
and U3819 (N_3819,N_2659,N_2708);
xnor U3820 (N_3820,N_3044,N_2496);
nand U3821 (N_3821,N_2623,N_3137);
and U3822 (N_3822,N_2932,N_3100);
and U3823 (N_3823,N_3010,N_2818);
nor U3824 (N_3824,N_2937,N_2430);
or U3825 (N_3825,N_3090,N_3181);
nand U3826 (N_3826,N_2793,N_2675);
xnor U3827 (N_3827,N_3197,N_2945);
nand U3828 (N_3828,N_2919,N_2570);
nor U3829 (N_3829,N_2902,N_2470);
and U3830 (N_3830,N_3111,N_3046);
and U3831 (N_3831,N_2460,N_3181);
or U3832 (N_3832,N_2810,N_3027);
xor U3833 (N_3833,N_3189,N_3023);
or U3834 (N_3834,N_2753,N_2924);
or U3835 (N_3835,N_2599,N_3053);
xnor U3836 (N_3836,N_2404,N_3156);
nand U3837 (N_3837,N_3189,N_2664);
and U3838 (N_3838,N_2856,N_3167);
and U3839 (N_3839,N_2455,N_2743);
nand U3840 (N_3840,N_2949,N_2966);
nor U3841 (N_3841,N_2646,N_2607);
or U3842 (N_3842,N_2757,N_2611);
xnor U3843 (N_3843,N_3062,N_2705);
nor U3844 (N_3844,N_2544,N_2903);
nor U3845 (N_3845,N_2971,N_2535);
xor U3846 (N_3846,N_2933,N_2453);
or U3847 (N_3847,N_3106,N_3081);
and U3848 (N_3848,N_2888,N_3190);
nand U3849 (N_3849,N_2945,N_3026);
nor U3850 (N_3850,N_2833,N_2733);
nor U3851 (N_3851,N_2408,N_2852);
and U3852 (N_3852,N_2514,N_2860);
nand U3853 (N_3853,N_2485,N_2521);
or U3854 (N_3854,N_3012,N_3122);
xor U3855 (N_3855,N_2668,N_2661);
xor U3856 (N_3856,N_2854,N_3137);
xor U3857 (N_3857,N_2982,N_2841);
or U3858 (N_3858,N_2734,N_2761);
nor U3859 (N_3859,N_3067,N_2797);
or U3860 (N_3860,N_2963,N_2880);
nor U3861 (N_3861,N_2974,N_2517);
nor U3862 (N_3862,N_3126,N_2615);
and U3863 (N_3863,N_2969,N_2746);
and U3864 (N_3864,N_2758,N_2853);
xnor U3865 (N_3865,N_2554,N_2960);
or U3866 (N_3866,N_2592,N_2999);
or U3867 (N_3867,N_3032,N_2735);
nor U3868 (N_3868,N_2487,N_3029);
and U3869 (N_3869,N_3095,N_2930);
or U3870 (N_3870,N_2480,N_2808);
nor U3871 (N_3871,N_2930,N_2894);
nand U3872 (N_3872,N_3149,N_2948);
or U3873 (N_3873,N_2982,N_2636);
and U3874 (N_3874,N_2650,N_2514);
or U3875 (N_3875,N_2421,N_3131);
or U3876 (N_3876,N_3157,N_2591);
xnor U3877 (N_3877,N_3172,N_2586);
and U3878 (N_3878,N_2750,N_2476);
and U3879 (N_3879,N_2610,N_2443);
xnor U3880 (N_3880,N_3009,N_2608);
nor U3881 (N_3881,N_2614,N_3005);
nor U3882 (N_3882,N_2406,N_2969);
xor U3883 (N_3883,N_3132,N_2679);
nand U3884 (N_3884,N_2572,N_2993);
xor U3885 (N_3885,N_3087,N_3027);
xor U3886 (N_3886,N_3069,N_2746);
or U3887 (N_3887,N_2445,N_3149);
nor U3888 (N_3888,N_3014,N_2617);
nand U3889 (N_3889,N_2916,N_2472);
xnor U3890 (N_3890,N_2578,N_2839);
xor U3891 (N_3891,N_2806,N_2877);
and U3892 (N_3892,N_2405,N_2579);
nand U3893 (N_3893,N_2842,N_3077);
xnor U3894 (N_3894,N_2626,N_3025);
and U3895 (N_3895,N_2833,N_2808);
or U3896 (N_3896,N_2727,N_2620);
nand U3897 (N_3897,N_2488,N_2911);
xnor U3898 (N_3898,N_2770,N_3167);
or U3899 (N_3899,N_2854,N_2596);
xor U3900 (N_3900,N_3125,N_2720);
nor U3901 (N_3901,N_3168,N_2446);
xnor U3902 (N_3902,N_2803,N_2476);
nor U3903 (N_3903,N_2551,N_2566);
xor U3904 (N_3904,N_2433,N_3099);
nand U3905 (N_3905,N_3090,N_3052);
xnor U3906 (N_3906,N_2707,N_3015);
nor U3907 (N_3907,N_2748,N_3134);
and U3908 (N_3908,N_2670,N_2522);
nor U3909 (N_3909,N_2706,N_2809);
or U3910 (N_3910,N_3134,N_2853);
nand U3911 (N_3911,N_2814,N_2490);
nand U3912 (N_3912,N_2463,N_2656);
nor U3913 (N_3913,N_2755,N_3003);
nor U3914 (N_3914,N_3048,N_2714);
and U3915 (N_3915,N_2636,N_2450);
nor U3916 (N_3916,N_2967,N_2428);
xor U3917 (N_3917,N_3049,N_2673);
nor U3918 (N_3918,N_2579,N_2852);
nor U3919 (N_3919,N_3041,N_3134);
nor U3920 (N_3920,N_3006,N_3005);
and U3921 (N_3921,N_2518,N_3123);
xor U3922 (N_3922,N_2640,N_3176);
xnor U3923 (N_3923,N_2775,N_2506);
nor U3924 (N_3924,N_2996,N_3189);
xor U3925 (N_3925,N_2505,N_3023);
or U3926 (N_3926,N_2918,N_2418);
and U3927 (N_3927,N_2823,N_3173);
or U3928 (N_3928,N_2449,N_2689);
or U3929 (N_3929,N_3145,N_2591);
nor U3930 (N_3930,N_2814,N_2515);
and U3931 (N_3931,N_3166,N_2488);
nand U3932 (N_3932,N_2750,N_2967);
or U3933 (N_3933,N_3089,N_2710);
nor U3934 (N_3934,N_2936,N_2545);
xnor U3935 (N_3935,N_2436,N_3162);
nor U3936 (N_3936,N_3097,N_2650);
and U3937 (N_3937,N_2619,N_2502);
nand U3938 (N_3938,N_2984,N_2760);
and U3939 (N_3939,N_3015,N_2611);
and U3940 (N_3940,N_3129,N_2519);
nor U3941 (N_3941,N_3026,N_2910);
and U3942 (N_3942,N_2742,N_2587);
nand U3943 (N_3943,N_2517,N_2686);
nand U3944 (N_3944,N_3030,N_2918);
xnor U3945 (N_3945,N_2658,N_3025);
nor U3946 (N_3946,N_2768,N_2548);
nor U3947 (N_3947,N_2804,N_2970);
xor U3948 (N_3948,N_3162,N_2406);
or U3949 (N_3949,N_2501,N_2832);
nand U3950 (N_3950,N_2432,N_2743);
and U3951 (N_3951,N_2522,N_2923);
nand U3952 (N_3952,N_2630,N_2869);
nand U3953 (N_3953,N_3160,N_3067);
and U3954 (N_3954,N_2846,N_3170);
xor U3955 (N_3955,N_2897,N_2871);
or U3956 (N_3956,N_3057,N_2716);
or U3957 (N_3957,N_2879,N_3116);
or U3958 (N_3958,N_2806,N_2673);
or U3959 (N_3959,N_2974,N_2703);
and U3960 (N_3960,N_2725,N_2709);
or U3961 (N_3961,N_2565,N_3122);
nor U3962 (N_3962,N_2894,N_2664);
and U3963 (N_3963,N_2889,N_2937);
and U3964 (N_3964,N_2869,N_2739);
and U3965 (N_3965,N_2819,N_2570);
nand U3966 (N_3966,N_2968,N_2870);
xnor U3967 (N_3967,N_2576,N_2701);
or U3968 (N_3968,N_2462,N_3079);
xor U3969 (N_3969,N_3180,N_2728);
and U3970 (N_3970,N_2607,N_2538);
and U3971 (N_3971,N_2661,N_2513);
and U3972 (N_3972,N_2580,N_2883);
xnor U3973 (N_3973,N_2811,N_2914);
nand U3974 (N_3974,N_2613,N_3111);
nor U3975 (N_3975,N_3104,N_2835);
xnor U3976 (N_3976,N_2720,N_2644);
nand U3977 (N_3977,N_3031,N_3151);
nand U3978 (N_3978,N_2947,N_3078);
xnor U3979 (N_3979,N_2805,N_2938);
and U3980 (N_3980,N_2482,N_2884);
nor U3981 (N_3981,N_2871,N_3144);
or U3982 (N_3982,N_3079,N_2650);
nand U3983 (N_3983,N_2554,N_2693);
or U3984 (N_3984,N_3132,N_3189);
xor U3985 (N_3985,N_2956,N_2973);
xnor U3986 (N_3986,N_3059,N_2700);
nor U3987 (N_3987,N_2864,N_2526);
and U3988 (N_3988,N_2470,N_2839);
nor U3989 (N_3989,N_2660,N_2852);
nand U3990 (N_3990,N_2747,N_3112);
nor U3991 (N_3991,N_2596,N_2957);
or U3992 (N_3992,N_3057,N_2524);
nor U3993 (N_3993,N_3038,N_2638);
and U3994 (N_3994,N_2830,N_2408);
and U3995 (N_3995,N_2881,N_2694);
nor U3996 (N_3996,N_2851,N_2866);
xor U3997 (N_3997,N_2973,N_2968);
and U3998 (N_3998,N_3078,N_2771);
nand U3999 (N_3999,N_2557,N_2899);
or U4000 (N_4000,N_3827,N_3466);
nor U4001 (N_4001,N_3345,N_3458);
and U4002 (N_4002,N_3501,N_3294);
xor U4003 (N_4003,N_3956,N_3262);
and U4004 (N_4004,N_3611,N_3768);
or U4005 (N_4005,N_3227,N_3223);
and U4006 (N_4006,N_3797,N_3798);
and U4007 (N_4007,N_3918,N_3464);
or U4008 (N_4008,N_3642,N_3689);
xor U4009 (N_4009,N_3468,N_3832);
nand U4010 (N_4010,N_3384,N_3792);
or U4011 (N_4011,N_3625,N_3891);
and U4012 (N_4012,N_3505,N_3606);
or U4013 (N_4013,N_3692,N_3705);
nor U4014 (N_4014,N_3872,N_3762);
or U4015 (N_4015,N_3856,N_3779);
nand U4016 (N_4016,N_3440,N_3946);
and U4017 (N_4017,N_3914,N_3803);
xnor U4018 (N_4018,N_3397,N_3900);
and U4019 (N_4019,N_3698,N_3351);
and U4020 (N_4020,N_3386,N_3691);
xnor U4021 (N_4021,N_3737,N_3251);
or U4022 (N_4022,N_3860,N_3765);
and U4023 (N_4023,N_3631,N_3562);
nor U4024 (N_4024,N_3534,N_3998);
nor U4025 (N_4025,N_3229,N_3320);
nand U4026 (N_4026,N_3919,N_3876);
nor U4027 (N_4027,N_3819,N_3252);
or U4028 (N_4028,N_3361,N_3371);
nand U4029 (N_4029,N_3927,N_3713);
and U4030 (N_4030,N_3341,N_3271);
nand U4031 (N_4031,N_3484,N_3554);
nand U4032 (N_4032,N_3994,N_3428);
and U4033 (N_4033,N_3436,N_3590);
or U4034 (N_4034,N_3742,N_3548);
or U4035 (N_4035,N_3204,N_3382);
nor U4036 (N_4036,N_3766,N_3981);
and U4037 (N_4037,N_3416,N_3888);
or U4038 (N_4038,N_3308,N_3461);
and U4039 (N_4039,N_3411,N_3884);
and U4040 (N_4040,N_3771,N_3926);
nor U4041 (N_4041,N_3365,N_3896);
nand U4042 (N_4042,N_3745,N_3527);
or U4043 (N_4043,N_3561,N_3995);
nand U4044 (N_4044,N_3323,N_3623);
nor U4045 (N_4045,N_3530,N_3759);
xor U4046 (N_4046,N_3254,N_3493);
nor U4047 (N_4047,N_3859,N_3373);
xnor U4048 (N_4048,N_3736,N_3201);
and U4049 (N_4049,N_3756,N_3697);
nand U4050 (N_4050,N_3482,N_3208);
or U4051 (N_4051,N_3282,N_3321);
and U4052 (N_4052,N_3454,N_3857);
nand U4053 (N_4053,N_3935,N_3302);
xnor U4054 (N_4054,N_3268,N_3734);
xor U4055 (N_4055,N_3376,N_3673);
xnor U4056 (N_4056,N_3659,N_3979);
or U4057 (N_4057,N_3586,N_3209);
nand U4058 (N_4058,N_3239,N_3634);
nand U4059 (N_4059,N_3350,N_3487);
nor U4060 (N_4060,N_3526,N_3267);
or U4061 (N_4061,N_3471,N_3406);
and U4062 (N_4062,N_3494,N_3894);
xnor U4063 (N_4063,N_3377,N_3917);
nand U4064 (N_4064,N_3322,N_3353);
and U4065 (N_4065,N_3617,N_3300);
or U4066 (N_4066,N_3887,N_3824);
or U4067 (N_4067,N_3543,N_3870);
or U4068 (N_4068,N_3687,N_3773);
or U4069 (N_4069,N_3746,N_3336);
and U4070 (N_4070,N_3408,N_3712);
or U4071 (N_4071,N_3751,N_3863);
and U4072 (N_4072,N_3304,N_3843);
and U4073 (N_4073,N_3709,N_3491);
or U4074 (N_4074,N_3865,N_3715);
and U4075 (N_4075,N_3629,N_3791);
or U4076 (N_4076,N_3654,N_3975);
xor U4077 (N_4077,N_3473,N_3265);
nor U4078 (N_4078,N_3389,N_3758);
and U4079 (N_4079,N_3477,N_3582);
xnor U4080 (N_4080,N_3702,N_3503);
xnor U4081 (N_4081,N_3546,N_3690);
nand U4082 (N_4082,N_3840,N_3982);
nand U4083 (N_4083,N_3842,N_3839);
and U4084 (N_4084,N_3815,N_3885);
xnor U4085 (N_4085,N_3895,N_3807);
or U4086 (N_4086,N_3696,N_3783);
nand U4087 (N_4087,N_3986,N_3708);
and U4088 (N_4088,N_3788,N_3646);
and U4089 (N_4089,N_3513,N_3287);
nor U4090 (N_4090,N_3816,N_3362);
nor U4091 (N_4091,N_3537,N_3882);
and U4092 (N_4092,N_3948,N_3971);
xnor U4093 (N_4093,N_3937,N_3347);
and U4094 (N_4094,N_3786,N_3695);
nor U4095 (N_4095,N_3729,N_3288);
nand U4096 (N_4096,N_3584,N_3851);
nor U4097 (N_4097,N_3793,N_3977);
or U4098 (N_4098,N_3460,N_3913);
and U4099 (N_4099,N_3557,N_3412);
nor U4100 (N_4100,N_3380,N_3396);
nor U4101 (N_4101,N_3923,N_3280);
or U4102 (N_4102,N_3472,N_3245);
or U4103 (N_4103,N_3735,N_3740);
and U4104 (N_4104,N_3565,N_3243);
nor U4105 (N_4105,N_3938,N_3366);
or U4106 (N_4106,N_3718,N_3647);
nand U4107 (N_4107,N_3355,N_3307);
nor U4108 (N_4108,N_3492,N_3834);
or U4109 (N_4109,N_3790,N_3645);
and U4110 (N_4110,N_3772,N_3508);
nand U4111 (N_4111,N_3587,N_3656);
xor U4112 (N_4112,N_3478,N_3244);
nand U4113 (N_4113,N_3560,N_3372);
and U4114 (N_4114,N_3680,N_3298);
and U4115 (N_4115,N_3855,N_3489);
or U4116 (N_4116,N_3480,N_3422);
or U4117 (N_4117,N_3669,N_3206);
or U4118 (N_4118,N_3306,N_3655);
or U4119 (N_4119,N_3983,N_3607);
or U4120 (N_4120,N_3214,N_3342);
nand U4121 (N_4121,N_3374,N_3359);
xor U4122 (N_4122,N_3533,N_3886);
nand U4123 (N_4123,N_3782,N_3674);
xnor U4124 (N_4124,N_3952,N_3398);
and U4125 (N_4125,N_3423,N_3552);
and U4126 (N_4126,N_3922,N_3542);
xnor U4127 (N_4127,N_3732,N_3987);
or U4128 (N_4128,N_3583,N_3499);
and U4129 (N_4129,N_3445,N_3749);
or U4130 (N_4130,N_3344,N_3720);
nand U4131 (N_4131,N_3609,N_3310);
and U4132 (N_4132,N_3662,N_3441);
xnor U4133 (N_4133,N_3540,N_3539);
nand U4134 (N_4134,N_3414,N_3932);
xor U4135 (N_4135,N_3760,N_3898);
nand U4136 (N_4136,N_3281,N_3675);
nand U4137 (N_4137,N_3593,N_3610);
or U4138 (N_4138,N_3504,N_3388);
or U4139 (N_4139,N_3812,N_3984);
xor U4140 (N_4140,N_3684,N_3597);
nand U4141 (N_4141,N_3621,N_3580);
and U4142 (N_4142,N_3969,N_3936);
nand U4143 (N_4143,N_3326,N_3405);
or U4144 (N_4144,N_3523,N_3248);
nor U4145 (N_4145,N_3947,N_3438);
and U4146 (N_4146,N_3949,N_3910);
and U4147 (N_4147,N_3272,N_3972);
nand U4148 (N_4148,N_3536,N_3589);
xor U4149 (N_4149,N_3991,N_3875);
or U4150 (N_4150,N_3448,N_3879);
nand U4151 (N_4151,N_3598,N_3453);
or U4152 (N_4152,N_3930,N_3837);
nand U4153 (N_4153,N_3763,N_3403);
and U4154 (N_4154,N_3550,N_3908);
or U4155 (N_4155,N_3578,N_3253);
or U4156 (N_4156,N_3595,N_3638);
and U4157 (N_4157,N_3385,N_3568);
or U4158 (N_4158,N_3592,N_3963);
xnor U4159 (N_4159,N_3943,N_3528);
xor U4160 (N_4160,N_3479,N_3219);
and U4161 (N_4161,N_3430,N_3228);
and U4162 (N_4162,N_3240,N_3420);
nand U4163 (N_4163,N_3614,N_3340);
nor U4164 (N_4164,N_3278,N_3805);
and U4165 (N_4165,N_3305,N_3725);
and U4166 (N_4166,N_3509,N_3928);
or U4167 (N_4167,N_3301,N_3439);
or U4168 (N_4168,N_3512,N_3230);
or U4169 (N_4169,N_3719,N_3902);
nor U4170 (N_4170,N_3474,N_3957);
and U4171 (N_4171,N_3613,N_3459);
or U4172 (N_4172,N_3821,N_3657);
nand U4173 (N_4173,N_3835,N_3814);
or U4174 (N_4174,N_3563,N_3225);
and U4175 (N_4175,N_3789,N_3427);
nand U4176 (N_4176,N_3699,N_3990);
or U4177 (N_4177,N_3360,N_3663);
nand U4178 (N_4178,N_3831,N_3434);
or U4179 (N_4179,N_3878,N_3522);
or U4180 (N_4180,N_3500,N_3337);
xor U4181 (N_4181,N_3847,N_3212);
nor U4182 (N_4182,N_3999,N_3324);
xnor U4183 (N_4183,N_3313,N_3246);
xor U4184 (N_4184,N_3848,N_3871);
nor U4185 (N_4185,N_3688,N_3640);
nand U4186 (N_4186,N_3748,N_3604);
and U4187 (N_4187,N_3330,N_3616);
nor U4188 (N_4188,N_3289,N_3600);
and U4189 (N_4189,N_3541,N_3869);
xnor U4190 (N_4190,N_3588,N_3311);
xnor U4191 (N_4191,N_3241,N_3258);
and U4192 (N_4192,N_3841,N_3232);
nand U4193 (N_4193,N_3899,N_3802);
nand U4194 (N_4194,N_3387,N_3905);
and U4195 (N_4195,N_3775,N_3576);
xor U4196 (N_4196,N_3309,N_3711);
nand U4197 (N_4197,N_3318,N_3612);
or U4198 (N_4198,N_3476,N_3391);
and U4199 (N_4199,N_3700,N_3714);
nor U4200 (N_4200,N_3635,N_3224);
and U4201 (N_4201,N_3497,N_3770);
nor U4202 (N_4202,N_3238,N_3432);
xor U4203 (N_4203,N_3222,N_3721);
nand U4204 (N_4204,N_3658,N_3897);
xor U4205 (N_4205,N_3653,N_3573);
or U4206 (N_4206,N_3437,N_3545);
nor U4207 (N_4207,N_3925,N_3596);
and U4208 (N_4208,N_3261,N_3681);
nor U4209 (N_4209,N_3602,N_3706);
nand U4210 (N_4210,N_3942,N_3202);
xor U4211 (N_4211,N_3383,N_3475);
or U4212 (N_4212,N_3652,N_3951);
or U4213 (N_4213,N_3495,N_3955);
nand U4214 (N_4214,N_3339,N_3915);
or U4215 (N_4215,N_3933,N_3348);
and U4216 (N_4216,N_3643,N_3375);
and U4217 (N_4217,N_3467,N_3808);
nand U4218 (N_4218,N_3618,N_3874);
nor U4219 (N_4219,N_3784,N_3757);
nand U4220 (N_4220,N_3764,N_3717);
xnor U4221 (N_4221,N_3993,N_3524);
nor U4222 (N_4222,N_3970,N_3818);
and U4223 (N_4223,N_3683,N_3394);
and U4224 (N_4224,N_3838,N_3510);
nand U4225 (N_4225,N_3585,N_3579);
or U4226 (N_4226,N_3833,N_3250);
nor U4227 (N_4227,N_3393,N_3907);
and U4228 (N_4228,N_3854,N_3744);
xnor U4229 (N_4229,N_3670,N_3236);
and U4230 (N_4230,N_3633,N_3378);
xnor U4231 (N_4231,N_3973,N_3517);
or U4232 (N_4232,N_3518,N_3769);
nand U4233 (N_4233,N_3447,N_3531);
and U4234 (N_4234,N_3911,N_3996);
xnor U4235 (N_4235,N_3456,N_3794);
nand U4236 (N_4236,N_3331,N_3678);
nand U4237 (N_4237,N_3877,N_3215);
and U4238 (N_4238,N_3893,N_3682);
and U4239 (N_4239,N_3203,N_3415);
xnor U4240 (N_4240,N_3485,N_3810);
nor U4241 (N_4241,N_3507,N_3776);
nor U4242 (N_4242,N_3486,N_3354);
xor U4243 (N_4243,N_3502,N_3242);
nand U4244 (N_4244,N_3599,N_3303);
xnor U4245 (N_4245,N_3968,N_3953);
nor U4246 (N_4246,N_3433,N_3753);
nor U4247 (N_4247,N_3519,N_3426);
nor U4248 (N_4248,N_3247,N_3574);
or U4249 (N_4249,N_3273,N_3358);
and U4250 (N_4250,N_3845,N_3672);
and U4251 (N_4251,N_3916,N_3904);
nand U4252 (N_4252,N_3231,N_3334);
and U4253 (N_4253,N_3980,N_3864);
nand U4254 (N_4254,N_3319,N_3551);
and U4255 (N_4255,N_3958,N_3525);
or U4256 (N_4256,N_3813,N_3777);
nand U4257 (N_4257,N_3210,N_3664);
nand U4258 (N_4258,N_3727,N_3627);
nand U4259 (N_4259,N_3892,N_3452);
nand U4260 (N_4260,N_3409,N_3685);
and U4261 (N_4261,N_3266,N_3976);
or U4262 (N_4262,N_3290,N_3463);
xnor U4263 (N_4263,N_3924,N_3569);
or U4264 (N_4264,N_3636,N_3451);
or U4265 (N_4265,N_3873,N_3315);
xor U4266 (N_4266,N_3858,N_3285);
and U4267 (N_4267,N_3823,N_3328);
nor U4268 (N_4268,N_3880,N_3444);
or U4269 (N_4269,N_3407,N_3667);
and U4270 (N_4270,N_3279,N_3395);
xnor U4271 (N_4271,N_3752,N_3716);
nor U4272 (N_4272,N_3269,N_3628);
nand U4273 (N_4273,N_3686,N_3293);
and U4274 (N_4274,N_3828,N_3449);
and U4275 (N_4275,N_3920,N_3939);
xnor U4276 (N_4276,N_3811,N_3694);
xnor U4277 (N_4277,N_3964,N_3577);
nand U4278 (N_4278,N_3778,N_3967);
nand U4279 (N_4279,N_3723,N_3470);
or U4280 (N_4280,N_3966,N_3619);
and U4281 (N_4281,N_3277,N_3520);
xnor U4282 (N_4282,N_3226,N_3558);
xor U4283 (N_4283,N_3274,N_3553);
xnor U4284 (N_4284,N_3676,N_3338);
or U4285 (N_4285,N_3710,N_3668);
xnor U4286 (N_4286,N_3852,N_3974);
nor U4287 (N_4287,N_3650,N_3529);
nor U4288 (N_4288,N_3862,N_3417);
nor U4289 (N_4289,N_3940,N_3799);
xnor U4290 (N_4290,N_3761,N_3327);
nand U4291 (N_4291,N_3603,N_3259);
nand U4292 (N_4292,N_3216,N_3255);
xnor U4293 (N_4293,N_3462,N_3796);
nand U4294 (N_4294,N_3379,N_3237);
xor U4295 (N_4295,N_3853,N_3890);
nand U4296 (N_4296,N_3787,N_3591);
and U4297 (N_4297,N_3465,N_3883);
nor U4298 (N_4298,N_3624,N_3850);
xnor U4299 (N_4299,N_3822,N_3564);
and U4300 (N_4300,N_3774,N_3220);
or U4301 (N_4301,N_3989,N_3992);
nor U4302 (N_4302,N_3481,N_3570);
xor U4303 (N_4303,N_3800,N_3844);
or U4304 (N_4304,N_3649,N_3665);
or U4305 (N_4305,N_3903,N_3299);
or U4306 (N_4306,N_3249,N_3260);
nand U4307 (N_4307,N_3496,N_3724);
and U4308 (N_4308,N_3620,N_3200);
nand U4309 (N_4309,N_3648,N_3400);
nor U4310 (N_4310,N_3825,N_3795);
nand U4311 (N_4311,N_3312,N_3516);
xnor U4312 (N_4312,N_3264,N_3965);
or U4313 (N_4313,N_3419,N_3651);
nand U4314 (N_4314,N_3929,N_3424);
xnor U4315 (N_4315,N_3572,N_3429);
xnor U4316 (N_4316,N_3747,N_3867);
or U4317 (N_4317,N_3335,N_3521);
xor U4318 (N_4318,N_3402,N_3731);
and U4319 (N_4319,N_3661,N_3442);
nand U4320 (N_4320,N_3829,N_3605);
nor U4321 (N_4321,N_3641,N_3703);
nand U4322 (N_4322,N_3276,N_3934);
and U4323 (N_4323,N_3901,N_3671);
and U4324 (N_4324,N_3931,N_3701);
and U4325 (N_4325,N_3483,N_3404);
xor U4326 (N_4326,N_3944,N_3544);
or U4327 (N_4327,N_3535,N_3780);
nand U4328 (N_4328,N_3733,N_3233);
nand U4329 (N_4329,N_3959,N_3660);
nor U4330 (N_4330,N_3511,N_3555);
nor U4331 (N_4331,N_3785,N_3263);
and U4332 (N_4332,N_3549,N_3960);
xor U4333 (N_4333,N_3352,N_3704);
nand U4334 (N_4334,N_3889,N_3817);
and U4335 (N_4335,N_3314,N_3217);
xnor U4336 (N_4336,N_3368,N_3413);
and U4337 (N_4337,N_3978,N_3804);
or U4338 (N_4338,N_3211,N_3962);
and U4339 (N_4339,N_3622,N_3488);
or U4340 (N_4340,N_3912,N_3988);
and U4341 (N_4341,N_3270,N_3571);
xor U4342 (N_4342,N_3921,N_3909);
xnor U4343 (N_4343,N_3349,N_3626);
and U4344 (N_4344,N_3566,N_3325);
or U4345 (N_4345,N_3861,N_3256);
and U4346 (N_4346,N_3559,N_3291);
nor U4347 (N_4347,N_3961,N_3849);
or U4348 (N_4348,N_3601,N_3399);
and U4349 (N_4349,N_3317,N_3450);
or U4350 (N_4350,N_3235,N_3425);
nand U4351 (N_4351,N_3275,N_3755);
nand U4352 (N_4352,N_3431,N_3781);
xor U4353 (N_4353,N_3632,N_3205);
or U4354 (N_4354,N_3881,N_3741);
nor U4355 (N_4355,N_3329,N_3722);
or U4356 (N_4356,N_3950,N_3356);
or U4357 (N_4357,N_3469,N_3213);
nor U4358 (N_4358,N_3868,N_3644);
xor U4359 (N_4359,N_3435,N_3809);
nor U4360 (N_4360,N_3750,N_3346);
and U4361 (N_4361,N_3728,N_3381);
or U4362 (N_4362,N_3506,N_3666);
and U4363 (N_4363,N_3295,N_3221);
and U4364 (N_4364,N_3846,N_3594);
and U4365 (N_4365,N_3806,N_3954);
or U4366 (N_4366,N_3754,N_3446);
nand U4367 (N_4367,N_3457,N_3739);
nand U4368 (N_4368,N_3836,N_3421);
or U4369 (N_4369,N_3639,N_3801);
or U4370 (N_4370,N_3693,N_3390);
and U4371 (N_4371,N_3637,N_3532);
or U4372 (N_4372,N_3410,N_3498);
xor U4373 (N_4373,N_3581,N_3369);
xor U4374 (N_4374,N_3679,N_3367);
nor U4375 (N_4375,N_3234,N_3333);
and U4376 (N_4376,N_3443,N_3297);
or U4377 (N_4377,N_3866,N_3615);
and U4378 (N_4378,N_3370,N_3707);
and U4379 (N_4379,N_3567,N_3401);
nor U4380 (N_4380,N_3207,N_3677);
and U4381 (N_4381,N_3738,N_3726);
or U4382 (N_4382,N_3945,N_3997);
or U4383 (N_4383,N_3556,N_3257);
xnor U4384 (N_4384,N_3743,N_3490);
nor U4385 (N_4385,N_3316,N_3515);
nor U4386 (N_4386,N_3630,N_3296);
nor U4387 (N_4387,N_3941,N_3218);
nand U4388 (N_4388,N_3575,N_3547);
or U4389 (N_4389,N_3906,N_3985);
xnor U4390 (N_4390,N_3826,N_3514);
nor U4391 (N_4391,N_3608,N_3363);
and U4392 (N_4392,N_3357,N_3292);
or U4393 (N_4393,N_3538,N_3820);
or U4394 (N_4394,N_3730,N_3343);
xor U4395 (N_4395,N_3392,N_3286);
or U4396 (N_4396,N_3283,N_3284);
nor U4397 (N_4397,N_3332,N_3767);
or U4398 (N_4398,N_3830,N_3455);
and U4399 (N_4399,N_3418,N_3364);
nand U4400 (N_4400,N_3495,N_3223);
xnor U4401 (N_4401,N_3280,N_3593);
nor U4402 (N_4402,N_3927,N_3215);
or U4403 (N_4403,N_3422,N_3871);
or U4404 (N_4404,N_3679,N_3502);
nor U4405 (N_4405,N_3672,N_3242);
nor U4406 (N_4406,N_3898,N_3571);
xor U4407 (N_4407,N_3711,N_3435);
nor U4408 (N_4408,N_3916,N_3521);
and U4409 (N_4409,N_3789,N_3778);
and U4410 (N_4410,N_3915,N_3316);
xnor U4411 (N_4411,N_3379,N_3911);
xor U4412 (N_4412,N_3966,N_3757);
xnor U4413 (N_4413,N_3913,N_3276);
nand U4414 (N_4414,N_3987,N_3212);
or U4415 (N_4415,N_3590,N_3792);
and U4416 (N_4416,N_3431,N_3758);
xnor U4417 (N_4417,N_3526,N_3880);
nand U4418 (N_4418,N_3204,N_3378);
nand U4419 (N_4419,N_3642,N_3351);
xor U4420 (N_4420,N_3705,N_3863);
xnor U4421 (N_4421,N_3931,N_3577);
nand U4422 (N_4422,N_3932,N_3787);
and U4423 (N_4423,N_3806,N_3490);
xor U4424 (N_4424,N_3602,N_3887);
xnor U4425 (N_4425,N_3346,N_3239);
nor U4426 (N_4426,N_3569,N_3534);
nor U4427 (N_4427,N_3352,N_3422);
nor U4428 (N_4428,N_3941,N_3799);
and U4429 (N_4429,N_3588,N_3829);
xor U4430 (N_4430,N_3288,N_3403);
xnor U4431 (N_4431,N_3353,N_3603);
nand U4432 (N_4432,N_3323,N_3297);
nor U4433 (N_4433,N_3835,N_3917);
nand U4434 (N_4434,N_3969,N_3702);
xor U4435 (N_4435,N_3368,N_3824);
nor U4436 (N_4436,N_3769,N_3990);
or U4437 (N_4437,N_3847,N_3255);
and U4438 (N_4438,N_3765,N_3314);
nor U4439 (N_4439,N_3717,N_3891);
or U4440 (N_4440,N_3208,N_3228);
or U4441 (N_4441,N_3813,N_3656);
xnor U4442 (N_4442,N_3330,N_3987);
and U4443 (N_4443,N_3769,N_3622);
xnor U4444 (N_4444,N_3840,N_3471);
xnor U4445 (N_4445,N_3434,N_3238);
or U4446 (N_4446,N_3901,N_3693);
xor U4447 (N_4447,N_3235,N_3565);
xor U4448 (N_4448,N_3458,N_3814);
nand U4449 (N_4449,N_3824,N_3631);
and U4450 (N_4450,N_3622,N_3730);
or U4451 (N_4451,N_3798,N_3344);
nor U4452 (N_4452,N_3811,N_3431);
nand U4453 (N_4453,N_3990,N_3265);
xnor U4454 (N_4454,N_3231,N_3757);
nor U4455 (N_4455,N_3533,N_3491);
or U4456 (N_4456,N_3467,N_3986);
and U4457 (N_4457,N_3524,N_3586);
nand U4458 (N_4458,N_3300,N_3243);
or U4459 (N_4459,N_3570,N_3421);
nand U4460 (N_4460,N_3340,N_3604);
and U4461 (N_4461,N_3849,N_3598);
nor U4462 (N_4462,N_3923,N_3255);
nor U4463 (N_4463,N_3773,N_3534);
nor U4464 (N_4464,N_3728,N_3655);
and U4465 (N_4465,N_3907,N_3564);
and U4466 (N_4466,N_3691,N_3918);
nor U4467 (N_4467,N_3894,N_3607);
nand U4468 (N_4468,N_3975,N_3464);
nand U4469 (N_4469,N_3873,N_3677);
and U4470 (N_4470,N_3716,N_3241);
nand U4471 (N_4471,N_3403,N_3669);
xor U4472 (N_4472,N_3365,N_3932);
nand U4473 (N_4473,N_3498,N_3940);
nand U4474 (N_4474,N_3968,N_3567);
nor U4475 (N_4475,N_3618,N_3238);
nand U4476 (N_4476,N_3910,N_3724);
nor U4477 (N_4477,N_3677,N_3374);
xor U4478 (N_4478,N_3867,N_3629);
nor U4479 (N_4479,N_3808,N_3679);
nor U4480 (N_4480,N_3975,N_3436);
and U4481 (N_4481,N_3820,N_3580);
or U4482 (N_4482,N_3277,N_3617);
nor U4483 (N_4483,N_3441,N_3621);
xnor U4484 (N_4484,N_3545,N_3504);
and U4485 (N_4485,N_3686,N_3947);
nor U4486 (N_4486,N_3580,N_3336);
nand U4487 (N_4487,N_3259,N_3598);
and U4488 (N_4488,N_3822,N_3972);
nor U4489 (N_4489,N_3975,N_3961);
xor U4490 (N_4490,N_3898,N_3470);
and U4491 (N_4491,N_3885,N_3842);
nand U4492 (N_4492,N_3280,N_3276);
and U4493 (N_4493,N_3745,N_3306);
nand U4494 (N_4494,N_3862,N_3665);
nand U4495 (N_4495,N_3819,N_3615);
xnor U4496 (N_4496,N_3922,N_3670);
or U4497 (N_4497,N_3858,N_3453);
nor U4498 (N_4498,N_3840,N_3990);
nand U4499 (N_4499,N_3336,N_3696);
xnor U4500 (N_4500,N_3686,N_3550);
xor U4501 (N_4501,N_3418,N_3261);
nor U4502 (N_4502,N_3327,N_3957);
or U4503 (N_4503,N_3882,N_3361);
nand U4504 (N_4504,N_3558,N_3259);
and U4505 (N_4505,N_3667,N_3294);
xor U4506 (N_4506,N_3536,N_3694);
and U4507 (N_4507,N_3662,N_3926);
or U4508 (N_4508,N_3729,N_3570);
and U4509 (N_4509,N_3992,N_3291);
nand U4510 (N_4510,N_3421,N_3687);
nand U4511 (N_4511,N_3635,N_3852);
xor U4512 (N_4512,N_3201,N_3473);
or U4513 (N_4513,N_3876,N_3859);
xor U4514 (N_4514,N_3856,N_3764);
nand U4515 (N_4515,N_3485,N_3565);
nor U4516 (N_4516,N_3470,N_3755);
and U4517 (N_4517,N_3261,N_3471);
xnor U4518 (N_4518,N_3651,N_3473);
nor U4519 (N_4519,N_3819,N_3918);
xnor U4520 (N_4520,N_3696,N_3921);
and U4521 (N_4521,N_3784,N_3947);
nor U4522 (N_4522,N_3668,N_3640);
and U4523 (N_4523,N_3469,N_3635);
nand U4524 (N_4524,N_3590,N_3448);
xnor U4525 (N_4525,N_3504,N_3814);
and U4526 (N_4526,N_3741,N_3387);
xnor U4527 (N_4527,N_3539,N_3427);
xor U4528 (N_4528,N_3204,N_3472);
nor U4529 (N_4529,N_3505,N_3514);
and U4530 (N_4530,N_3898,N_3244);
nand U4531 (N_4531,N_3666,N_3895);
and U4532 (N_4532,N_3324,N_3251);
or U4533 (N_4533,N_3617,N_3572);
nor U4534 (N_4534,N_3899,N_3792);
or U4535 (N_4535,N_3358,N_3625);
nor U4536 (N_4536,N_3501,N_3516);
or U4537 (N_4537,N_3395,N_3964);
or U4538 (N_4538,N_3528,N_3779);
and U4539 (N_4539,N_3748,N_3812);
nand U4540 (N_4540,N_3945,N_3547);
and U4541 (N_4541,N_3756,N_3890);
nand U4542 (N_4542,N_3560,N_3231);
xnor U4543 (N_4543,N_3337,N_3525);
nand U4544 (N_4544,N_3332,N_3620);
nand U4545 (N_4545,N_3336,N_3625);
or U4546 (N_4546,N_3414,N_3865);
or U4547 (N_4547,N_3779,N_3545);
nand U4548 (N_4548,N_3253,N_3407);
and U4549 (N_4549,N_3881,N_3434);
or U4550 (N_4550,N_3972,N_3428);
or U4551 (N_4551,N_3631,N_3625);
nand U4552 (N_4552,N_3780,N_3898);
nand U4553 (N_4553,N_3595,N_3456);
nand U4554 (N_4554,N_3344,N_3467);
and U4555 (N_4555,N_3405,N_3471);
or U4556 (N_4556,N_3584,N_3543);
nor U4557 (N_4557,N_3667,N_3349);
and U4558 (N_4558,N_3740,N_3485);
xor U4559 (N_4559,N_3958,N_3725);
nor U4560 (N_4560,N_3678,N_3216);
nand U4561 (N_4561,N_3763,N_3906);
nand U4562 (N_4562,N_3231,N_3268);
or U4563 (N_4563,N_3246,N_3318);
and U4564 (N_4564,N_3710,N_3974);
and U4565 (N_4565,N_3648,N_3451);
nand U4566 (N_4566,N_3285,N_3992);
nand U4567 (N_4567,N_3380,N_3924);
xnor U4568 (N_4568,N_3712,N_3896);
or U4569 (N_4569,N_3788,N_3740);
and U4570 (N_4570,N_3606,N_3725);
nand U4571 (N_4571,N_3983,N_3410);
nor U4572 (N_4572,N_3824,N_3810);
or U4573 (N_4573,N_3962,N_3400);
nor U4574 (N_4574,N_3211,N_3549);
nand U4575 (N_4575,N_3982,N_3868);
or U4576 (N_4576,N_3804,N_3604);
nand U4577 (N_4577,N_3308,N_3586);
nand U4578 (N_4578,N_3643,N_3252);
nor U4579 (N_4579,N_3593,N_3605);
and U4580 (N_4580,N_3432,N_3212);
xor U4581 (N_4581,N_3538,N_3473);
and U4582 (N_4582,N_3931,N_3562);
nand U4583 (N_4583,N_3861,N_3659);
or U4584 (N_4584,N_3651,N_3858);
or U4585 (N_4585,N_3316,N_3207);
and U4586 (N_4586,N_3712,N_3350);
and U4587 (N_4587,N_3658,N_3621);
and U4588 (N_4588,N_3887,N_3963);
nand U4589 (N_4589,N_3764,N_3438);
nand U4590 (N_4590,N_3277,N_3888);
and U4591 (N_4591,N_3825,N_3248);
nand U4592 (N_4592,N_3462,N_3777);
xnor U4593 (N_4593,N_3688,N_3610);
xnor U4594 (N_4594,N_3908,N_3684);
and U4595 (N_4595,N_3350,N_3721);
and U4596 (N_4596,N_3990,N_3827);
xnor U4597 (N_4597,N_3586,N_3786);
nand U4598 (N_4598,N_3680,N_3945);
and U4599 (N_4599,N_3953,N_3482);
nand U4600 (N_4600,N_3797,N_3355);
nor U4601 (N_4601,N_3615,N_3456);
xnor U4602 (N_4602,N_3965,N_3753);
xor U4603 (N_4603,N_3959,N_3688);
nand U4604 (N_4604,N_3737,N_3968);
xnor U4605 (N_4605,N_3549,N_3934);
xnor U4606 (N_4606,N_3389,N_3993);
xor U4607 (N_4607,N_3805,N_3396);
or U4608 (N_4608,N_3902,N_3686);
nand U4609 (N_4609,N_3680,N_3436);
nor U4610 (N_4610,N_3348,N_3582);
nor U4611 (N_4611,N_3368,N_3496);
nand U4612 (N_4612,N_3490,N_3549);
or U4613 (N_4613,N_3840,N_3651);
or U4614 (N_4614,N_3289,N_3516);
nand U4615 (N_4615,N_3271,N_3606);
or U4616 (N_4616,N_3492,N_3807);
or U4617 (N_4617,N_3908,N_3806);
or U4618 (N_4618,N_3382,N_3317);
nor U4619 (N_4619,N_3932,N_3847);
and U4620 (N_4620,N_3823,N_3401);
nand U4621 (N_4621,N_3667,N_3369);
nor U4622 (N_4622,N_3394,N_3722);
nand U4623 (N_4623,N_3742,N_3467);
or U4624 (N_4624,N_3272,N_3474);
xnor U4625 (N_4625,N_3634,N_3329);
nand U4626 (N_4626,N_3507,N_3805);
or U4627 (N_4627,N_3543,N_3900);
and U4628 (N_4628,N_3797,N_3529);
nor U4629 (N_4629,N_3583,N_3857);
nand U4630 (N_4630,N_3877,N_3995);
xor U4631 (N_4631,N_3807,N_3977);
and U4632 (N_4632,N_3236,N_3502);
nor U4633 (N_4633,N_3673,N_3337);
or U4634 (N_4634,N_3540,N_3714);
xor U4635 (N_4635,N_3782,N_3364);
nand U4636 (N_4636,N_3544,N_3606);
or U4637 (N_4637,N_3815,N_3660);
or U4638 (N_4638,N_3345,N_3469);
or U4639 (N_4639,N_3927,N_3414);
nand U4640 (N_4640,N_3563,N_3382);
or U4641 (N_4641,N_3700,N_3938);
nor U4642 (N_4642,N_3639,N_3297);
nor U4643 (N_4643,N_3890,N_3722);
or U4644 (N_4644,N_3512,N_3473);
nand U4645 (N_4645,N_3928,N_3967);
and U4646 (N_4646,N_3981,N_3216);
xnor U4647 (N_4647,N_3511,N_3819);
xor U4648 (N_4648,N_3949,N_3533);
nor U4649 (N_4649,N_3569,N_3446);
xnor U4650 (N_4650,N_3848,N_3923);
nor U4651 (N_4651,N_3480,N_3805);
nand U4652 (N_4652,N_3935,N_3562);
and U4653 (N_4653,N_3882,N_3459);
and U4654 (N_4654,N_3417,N_3523);
and U4655 (N_4655,N_3203,N_3783);
nand U4656 (N_4656,N_3736,N_3415);
and U4657 (N_4657,N_3990,N_3255);
nand U4658 (N_4658,N_3689,N_3398);
nand U4659 (N_4659,N_3341,N_3661);
xnor U4660 (N_4660,N_3775,N_3888);
nor U4661 (N_4661,N_3980,N_3236);
or U4662 (N_4662,N_3900,N_3554);
nand U4663 (N_4663,N_3757,N_3696);
and U4664 (N_4664,N_3871,N_3418);
nand U4665 (N_4665,N_3298,N_3352);
or U4666 (N_4666,N_3534,N_3301);
nor U4667 (N_4667,N_3642,N_3210);
or U4668 (N_4668,N_3307,N_3437);
nor U4669 (N_4669,N_3219,N_3211);
and U4670 (N_4670,N_3415,N_3222);
xor U4671 (N_4671,N_3324,N_3747);
nand U4672 (N_4672,N_3636,N_3535);
and U4673 (N_4673,N_3285,N_3938);
or U4674 (N_4674,N_3856,N_3278);
nand U4675 (N_4675,N_3401,N_3894);
nor U4676 (N_4676,N_3448,N_3872);
xnor U4677 (N_4677,N_3758,N_3289);
and U4678 (N_4678,N_3297,N_3894);
and U4679 (N_4679,N_3401,N_3659);
xnor U4680 (N_4680,N_3273,N_3648);
xnor U4681 (N_4681,N_3620,N_3428);
nor U4682 (N_4682,N_3374,N_3354);
nand U4683 (N_4683,N_3469,N_3686);
and U4684 (N_4684,N_3903,N_3545);
nand U4685 (N_4685,N_3876,N_3477);
xor U4686 (N_4686,N_3346,N_3218);
nand U4687 (N_4687,N_3239,N_3743);
or U4688 (N_4688,N_3616,N_3548);
or U4689 (N_4689,N_3565,N_3548);
nand U4690 (N_4690,N_3642,N_3743);
and U4691 (N_4691,N_3680,N_3902);
and U4692 (N_4692,N_3253,N_3972);
or U4693 (N_4693,N_3742,N_3249);
and U4694 (N_4694,N_3243,N_3806);
nand U4695 (N_4695,N_3561,N_3250);
and U4696 (N_4696,N_3975,N_3864);
nor U4697 (N_4697,N_3317,N_3285);
nor U4698 (N_4698,N_3559,N_3931);
and U4699 (N_4699,N_3491,N_3364);
or U4700 (N_4700,N_3295,N_3407);
and U4701 (N_4701,N_3321,N_3917);
xnor U4702 (N_4702,N_3589,N_3697);
xnor U4703 (N_4703,N_3896,N_3366);
nand U4704 (N_4704,N_3958,N_3765);
nor U4705 (N_4705,N_3636,N_3724);
nor U4706 (N_4706,N_3737,N_3351);
and U4707 (N_4707,N_3398,N_3604);
nor U4708 (N_4708,N_3270,N_3246);
nor U4709 (N_4709,N_3275,N_3304);
xnor U4710 (N_4710,N_3278,N_3925);
nand U4711 (N_4711,N_3946,N_3361);
nand U4712 (N_4712,N_3960,N_3477);
nor U4713 (N_4713,N_3491,N_3535);
and U4714 (N_4714,N_3405,N_3542);
nand U4715 (N_4715,N_3323,N_3711);
xor U4716 (N_4716,N_3424,N_3695);
nor U4717 (N_4717,N_3769,N_3980);
xnor U4718 (N_4718,N_3454,N_3337);
or U4719 (N_4719,N_3573,N_3465);
and U4720 (N_4720,N_3744,N_3701);
nor U4721 (N_4721,N_3868,N_3651);
nor U4722 (N_4722,N_3670,N_3310);
and U4723 (N_4723,N_3749,N_3223);
nor U4724 (N_4724,N_3405,N_3730);
or U4725 (N_4725,N_3749,N_3775);
nor U4726 (N_4726,N_3671,N_3274);
nand U4727 (N_4727,N_3407,N_3922);
or U4728 (N_4728,N_3229,N_3941);
nand U4729 (N_4729,N_3966,N_3342);
nor U4730 (N_4730,N_3546,N_3432);
nor U4731 (N_4731,N_3977,N_3969);
nor U4732 (N_4732,N_3602,N_3275);
xor U4733 (N_4733,N_3773,N_3665);
xnor U4734 (N_4734,N_3237,N_3992);
xor U4735 (N_4735,N_3229,N_3828);
nor U4736 (N_4736,N_3257,N_3280);
nand U4737 (N_4737,N_3928,N_3793);
xnor U4738 (N_4738,N_3616,N_3278);
and U4739 (N_4739,N_3327,N_3857);
and U4740 (N_4740,N_3475,N_3833);
or U4741 (N_4741,N_3316,N_3706);
and U4742 (N_4742,N_3476,N_3803);
nand U4743 (N_4743,N_3319,N_3931);
nor U4744 (N_4744,N_3914,N_3307);
nand U4745 (N_4745,N_3637,N_3577);
nor U4746 (N_4746,N_3838,N_3980);
and U4747 (N_4747,N_3639,N_3726);
nor U4748 (N_4748,N_3624,N_3992);
nor U4749 (N_4749,N_3379,N_3904);
and U4750 (N_4750,N_3544,N_3530);
or U4751 (N_4751,N_3859,N_3496);
nor U4752 (N_4752,N_3975,N_3278);
xor U4753 (N_4753,N_3720,N_3347);
and U4754 (N_4754,N_3744,N_3836);
or U4755 (N_4755,N_3856,N_3430);
nor U4756 (N_4756,N_3960,N_3826);
nor U4757 (N_4757,N_3743,N_3410);
or U4758 (N_4758,N_3926,N_3366);
xor U4759 (N_4759,N_3497,N_3350);
xor U4760 (N_4760,N_3882,N_3515);
and U4761 (N_4761,N_3429,N_3331);
nor U4762 (N_4762,N_3627,N_3730);
and U4763 (N_4763,N_3505,N_3610);
xor U4764 (N_4764,N_3706,N_3378);
xor U4765 (N_4765,N_3591,N_3398);
and U4766 (N_4766,N_3375,N_3768);
xnor U4767 (N_4767,N_3463,N_3706);
or U4768 (N_4768,N_3532,N_3819);
and U4769 (N_4769,N_3792,N_3424);
nand U4770 (N_4770,N_3953,N_3772);
and U4771 (N_4771,N_3809,N_3733);
and U4772 (N_4772,N_3344,N_3459);
or U4773 (N_4773,N_3826,N_3622);
nand U4774 (N_4774,N_3696,N_3890);
nand U4775 (N_4775,N_3758,N_3812);
or U4776 (N_4776,N_3251,N_3204);
nor U4777 (N_4777,N_3651,N_3326);
and U4778 (N_4778,N_3415,N_3847);
or U4779 (N_4779,N_3559,N_3926);
or U4780 (N_4780,N_3615,N_3264);
or U4781 (N_4781,N_3878,N_3843);
xnor U4782 (N_4782,N_3343,N_3572);
xnor U4783 (N_4783,N_3684,N_3471);
nand U4784 (N_4784,N_3335,N_3563);
xor U4785 (N_4785,N_3619,N_3995);
nand U4786 (N_4786,N_3285,N_3346);
and U4787 (N_4787,N_3820,N_3305);
or U4788 (N_4788,N_3829,N_3700);
or U4789 (N_4789,N_3689,N_3819);
xor U4790 (N_4790,N_3591,N_3725);
or U4791 (N_4791,N_3564,N_3898);
or U4792 (N_4792,N_3797,N_3393);
nor U4793 (N_4793,N_3571,N_3519);
xor U4794 (N_4794,N_3608,N_3470);
xor U4795 (N_4795,N_3982,N_3651);
or U4796 (N_4796,N_3949,N_3701);
or U4797 (N_4797,N_3752,N_3575);
nand U4798 (N_4798,N_3721,N_3634);
xnor U4799 (N_4799,N_3852,N_3213);
xor U4800 (N_4800,N_4706,N_4235);
nor U4801 (N_4801,N_4175,N_4022);
nand U4802 (N_4802,N_4359,N_4250);
and U4803 (N_4803,N_4561,N_4459);
and U4804 (N_4804,N_4742,N_4762);
and U4805 (N_4805,N_4255,N_4358);
and U4806 (N_4806,N_4215,N_4229);
xor U4807 (N_4807,N_4698,N_4398);
xnor U4808 (N_4808,N_4282,N_4313);
nor U4809 (N_4809,N_4604,N_4444);
nor U4810 (N_4810,N_4648,N_4288);
nor U4811 (N_4811,N_4478,N_4070);
xnor U4812 (N_4812,N_4009,N_4180);
nor U4813 (N_4813,N_4258,N_4060);
and U4814 (N_4814,N_4150,N_4073);
nor U4815 (N_4815,N_4120,N_4512);
nand U4816 (N_4816,N_4211,N_4731);
and U4817 (N_4817,N_4470,N_4681);
nor U4818 (N_4818,N_4671,N_4349);
nor U4819 (N_4819,N_4422,N_4787);
or U4820 (N_4820,N_4686,N_4602);
xor U4821 (N_4821,N_4216,N_4106);
and U4822 (N_4822,N_4270,N_4362);
xnor U4823 (N_4823,N_4179,N_4003);
nor U4824 (N_4824,N_4074,N_4432);
nor U4825 (N_4825,N_4791,N_4528);
xor U4826 (N_4826,N_4333,N_4661);
nand U4827 (N_4827,N_4663,N_4218);
nand U4828 (N_4828,N_4565,N_4506);
nand U4829 (N_4829,N_4361,N_4247);
xor U4830 (N_4830,N_4775,N_4522);
or U4831 (N_4831,N_4597,N_4057);
and U4832 (N_4832,N_4352,N_4161);
xor U4833 (N_4833,N_4507,N_4689);
nor U4834 (N_4834,N_4547,N_4222);
nor U4835 (N_4835,N_4371,N_4690);
and U4836 (N_4836,N_4101,N_4283);
nand U4837 (N_4837,N_4440,N_4578);
xnor U4838 (N_4838,N_4025,N_4510);
nor U4839 (N_4839,N_4027,N_4311);
nor U4840 (N_4840,N_4325,N_4401);
or U4841 (N_4841,N_4389,N_4103);
xor U4842 (N_4842,N_4607,N_4285);
nor U4843 (N_4843,N_4675,N_4557);
or U4844 (N_4844,N_4031,N_4276);
nor U4845 (N_4845,N_4062,N_4356);
xnor U4846 (N_4846,N_4296,N_4092);
xnor U4847 (N_4847,N_4188,N_4453);
nor U4848 (N_4848,N_4608,N_4201);
nor U4849 (N_4849,N_4720,N_4754);
nand U4850 (N_4850,N_4335,N_4368);
xor U4851 (N_4851,N_4600,N_4446);
nor U4852 (N_4852,N_4451,N_4035);
xor U4853 (N_4853,N_4643,N_4577);
nand U4854 (N_4854,N_4511,N_4743);
xnor U4855 (N_4855,N_4054,N_4007);
or U4856 (N_4856,N_4476,N_4580);
nand U4857 (N_4857,N_4078,N_4606);
nand U4858 (N_4858,N_4532,N_4550);
nand U4859 (N_4859,N_4526,N_4190);
and U4860 (N_4860,N_4384,N_4341);
or U4861 (N_4861,N_4403,N_4075);
nand U4862 (N_4862,N_4323,N_4688);
or U4863 (N_4863,N_4234,N_4677);
nor U4864 (N_4864,N_4518,N_4297);
and U4865 (N_4865,N_4122,N_4289);
and U4866 (N_4866,N_4579,N_4337);
nor U4867 (N_4867,N_4725,N_4394);
or U4868 (N_4868,N_4491,N_4248);
xnor U4869 (N_4869,N_4269,N_4588);
nand U4870 (N_4870,N_4280,N_4628);
and U4871 (N_4871,N_4146,N_4411);
nor U4872 (N_4872,N_4202,N_4082);
and U4873 (N_4873,N_4737,N_4366);
nand U4874 (N_4874,N_4438,N_4271);
and U4875 (N_4875,N_4264,N_4257);
xnor U4876 (N_4876,N_4065,N_4044);
nor U4877 (N_4877,N_4238,N_4474);
or U4878 (N_4878,N_4553,N_4773);
nor U4879 (N_4879,N_4590,N_4030);
or U4880 (N_4880,N_4575,N_4627);
or U4881 (N_4881,N_4166,N_4170);
or U4882 (N_4882,N_4709,N_4443);
xor U4883 (N_4883,N_4548,N_4716);
and U4884 (N_4884,N_4515,N_4680);
xnor U4885 (N_4885,N_4479,N_4441);
or U4886 (N_4886,N_4342,N_4149);
or U4887 (N_4887,N_4733,N_4041);
and U4888 (N_4888,N_4767,N_4763);
nor U4889 (N_4889,N_4402,N_4516);
and U4890 (N_4890,N_4480,N_4535);
nand U4891 (N_4891,N_4204,N_4284);
nand U4892 (N_4892,N_4562,N_4423);
xnor U4893 (N_4893,N_4094,N_4464);
xnor U4894 (N_4894,N_4231,N_4324);
nand U4895 (N_4895,N_4736,N_4496);
or U4896 (N_4896,N_4481,N_4447);
or U4897 (N_4897,N_4042,N_4712);
nand U4898 (N_4898,N_4461,N_4002);
nand U4899 (N_4899,N_4719,N_4387);
nand U4900 (N_4900,N_4372,N_4240);
xnor U4901 (N_4901,N_4585,N_4397);
xor U4902 (N_4902,N_4353,N_4412);
and U4903 (N_4903,N_4764,N_4158);
or U4904 (N_4904,N_4084,N_4263);
nor U4905 (N_4905,N_4710,N_4097);
or U4906 (N_4906,N_4584,N_4460);
nand U4907 (N_4907,N_4046,N_4458);
nor U4908 (N_4908,N_4406,N_4772);
and U4909 (N_4909,N_4336,N_4254);
or U4910 (N_4910,N_4208,N_4610);
xnor U4911 (N_4911,N_4052,N_4489);
nand U4912 (N_4912,N_4455,N_4755);
nand U4913 (N_4913,N_4430,N_4727);
or U4914 (N_4914,N_4020,N_4795);
nand U4915 (N_4915,N_4750,N_4252);
nand U4916 (N_4916,N_4650,N_4645);
xnor U4917 (N_4917,N_4644,N_4500);
nor U4918 (N_4918,N_4711,N_4129);
and U4919 (N_4919,N_4472,N_4262);
or U4920 (N_4920,N_4355,N_4088);
or U4921 (N_4921,N_4291,N_4753);
xnor U4922 (N_4922,N_4242,N_4135);
xor U4923 (N_4923,N_4564,N_4539);
and U4924 (N_4924,N_4182,N_4026);
or U4925 (N_4925,N_4312,N_4574);
nor U4926 (N_4926,N_4439,N_4452);
and U4927 (N_4927,N_4334,N_4164);
and U4928 (N_4928,N_4339,N_4345);
and U4929 (N_4929,N_4782,N_4249);
nor U4930 (N_4930,N_4195,N_4200);
or U4931 (N_4931,N_4601,N_4674);
nor U4932 (N_4932,N_4399,N_4653);
nand U4933 (N_4933,N_4793,N_4792);
nand U4934 (N_4934,N_4682,N_4300);
and U4935 (N_4935,N_4672,N_4523);
xor U4936 (N_4936,N_4064,N_4540);
nor U4937 (N_4937,N_4319,N_4000);
nand U4938 (N_4938,N_4330,N_4102);
nor U4939 (N_4939,N_4011,N_4147);
xnor U4940 (N_4940,N_4244,N_4327);
xor U4941 (N_4941,N_4437,N_4697);
and U4942 (N_4942,N_4056,N_4377);
or U4943 (N_4943,N_4373,N_4199);
and U4944 (N_4944,N_4008,N_4419);
nor U4945 (N_4945,N_4637,N_4486);
and U4946 (N_4946,N_4301,N_4369);
nor U4947 (N_4947,N_4294,N_4615);
and U4948 (N_4948,N_4251,N_4220);
or U4949 (N_4949,N_4531,N_4529);
nor U4950 (N_4950,N_4560,N_4729);
nand U4951 (N_4951,N_4622,N_4429);
nor U4952 (N_4952,N_4457,N_4237);
nor U4953 (N_4953,N_4721,N_4286);
nor U4954 (N_4954,N_4351,N_4173);
nand U4955 (N_4955,N_4141,N_4517);
nand U4956 (N_4956,N_4405,N_4108);
nor U4957 (N_4957,N_4114,N_4365);
xnor U4958 (N_4958,N_4281,N_4274);
nor U4959 (N_4959,N_4445,N_4024);
or U4960 (N_4960,N_4752,N_4587);
nor U4961 (N_4961,N_4794,N_4105);
or U4962 (N_4962,N_4685,N_4664);
nand U4963 (N_4963,N_4077,N_4219);
nor U4964 (N_4964,N_4536,N_4665);
nand U4965 (N_4965,N_4213,N_4107);
nand U4966 (N_4966,N_4467,N_4293);
nand U4967 (N_4967,N_4646,N_4181);
nor U4968 (N_4968,N_4408,N_4425);
or U4969 (N_4969,N_4555,N_4551);
and U4970 (N_4970,N_4509,N_4226);
or U4971 (N_4971,N_4570,N_4156);
xor U4972 (N_4972,N_4673,N_4477);
or U4973 (N_4973,N_4169,N_4694);
xnor U4974 (N_4974,N_4299,N_4050);
nand U4975 (N_4975,N_4519,N_4061);
nand U4976 (N_4976,N_4593,N_4450);
nor U4977 (N_4977,N_4413,N_4099);
nand U4978 (N_4978,N_4468,N_4045);
nand U4979 (N_4979,N_4168,N_4370);
and U4980 (N_4980,N_4314,N_4253);
xnor U4981 (N_4981,N_4131,N_4781);
xor U4982 (N_4982,N_4513,N_4048);
nor U4983 (N_4983,N_4189,N_4005);
nand U4984 (N_4984,N_4692,N_4683);
nand U4985 (N_4985,N_4656,N_4434);
and U4986 (N_4986,N_4144,N_4130);
xnor U4987 (N_4987,N_4163,N_4040);
nand U4988 (N_4988,N_4758,N_4265);
xor U4989 (N_4989,N_4599,N_4592);
and U4990 (N_4990,N_4124,N_4055);
nand U4991 (N_4991,N_4326,N_4051);
and U4992 (N_4992,N_4081,N_4514);
and U4993 (N_4993,N_4797,N_4657);
and U4994 (N_4994,N_4196,N_4594);
or U4995 (N_4995,N_4748,N_4230);
xnor U4996 (N_4996,N_4115,N_4520);
nor U4997 (N_4997,N_4649,N_4449);
nor U4998 (N_4998,N_4780,N_4212);
xnor U4999 (N_4999,N_4171,N_4724);
nor U5000 (N_5000,N_4471,N_4713);
nand U5001 (N_5001,N_4768,N_4110);
nand U5002 (N_5002,N_4634,N_4306);
nand U5003 (N_5003,N_4788,N_4347);
and U5004 (N_5004,N_4176,N_4383);
xnor U5005 (N_5005,N_4160,N_4310);
xnor U5006 (N_5006,N_4277,N_4396);
and U5007 (N_5007,N_4591,N_4693);
nor U5008 (N_5008,N_4400,N_4331);
or U5009 (N_5009,N_4209,N_4123);
nor U5010 (N_5010,N_4172,N_4783);
and U5011 (N_5011,N_4490,N_4089);
nor U5012 (N_5012,N_4162,N_4036);
and U5013 (N_5013,N_4165,N_4620);
xnor U5014 (N_5014,N_4224,N_4275);
nor U5015 (N_5015,N_4696,N_4542);
xnor U5016 (N_5016,N_4076,N_4626);
and U5017 (N_5017,N_4318,N_4796);
xnor U5018 (N_5018,N_4316,N_4143);
nor U5019 (N_5019,N_4360,N_4418);
nor U5020 (N_5020,N_4544,N_4687);
and U5021 (N_5021,N_4572,N_4223);
nor U5022 (N_5022,N_4053,N_4734);
nor U5023 (N_5023,N_4667,N_4521);
and U5024 (N_5024,N_4625,N_4098);
xor U5025 (N_5025,N_4328,N_4639);
nand U5026 (N_5026,N_4139,N_4501);
and U5027 (N_5027,N_4658,N_4485);
xor U5028 (N_5028,N_4295,N_4707);
xnor U5029 (N_5029,N_4708,N_4197);
and U5030 (N_5030,N_4395,N_4239);
and U5031 (N_5031,N_4183,N_4256);
xor U5032 (N_5032,N_4701,N_4730);
nand U5033 (N_5033,N_4636,N_4431);
and U5034 (N_5034,N_4746,N_4738);
nand U5035 (N_5035,N_4338,N_4571);
nand U5036 (N_5036,N_4699,N_4225);
and U5037 (N_5037,N_4037,N_4576);
nor U5038 (N_5038,N_4340,N_4740);
nor U5039 (N_5039,N_4187,N_4380);
nor U5040 (N_5040,N_4145,N_4136);
xor U5041 (N_5041,N_4777,N_4668);
or U5042 (N_5042,N_4603,N_4006);
nand U5043 (N_5043,N_4148,N_4494);
xor U5044 (N_5044,N_4379,N_4504);
and U5045 (N_5045,N_4072,N_4589);
nor U5046 (N_5046,N_4385,N_4483);
nand U5047 (N_5047,N_4635,N_4442);
xor U5048 (N_5048,N_4482,N_4344);
or U5049 (N_5049,N_4343,N_4315);
nor U5050 (N_5050,N_4524,N_4032);
xnor U5051 (N_5051,N_4140,N_4421);
xnor U5052 (N_5052,N_4534,N_4317);
nand U5053 (N_5053,N_4178,N_4221);
and U5054 (N_5054,N_4121,N_4760);
or U5055 (N_5055,N_4613,N_4016);
nor U5056 (N_5056,N_4266,N_4132);
or U5057 (N_5057,N_4066,N_4417);
nand U5058 (N_5058,N_4079,N_4320);
nor U5059 (N_5059,N_4420,N_4279);
xnor U5060 (N_5060,N_4354,N_4582);
nor U5061 (N_5061,N_4495,N_4757);
or U5062 (N_5062,N_4090,N_4367);
nor U5063 (N_5063,N_4382,N_4784);
nand U5064 (N_5064,N_4659,N_4722);
nand U5065 (N_5065,N_4033,N_4741);
or U5066 (N_5066,N_4670,N_4109);
or U5067 (N_5067,N_4798,N_4013);
and U5068 (N_5068,N_4463,N_4745);
nand U5069 (N_5069,N_4039,N_4184);
nand U5070 (N_5070,N_4116,N_4492);
or U5071 (N_5071,N_4018,N_4268);
nand U5072 (N_5072,N_4508,N_4038);
and U5073 (N_5073,N_4227,N_4647);
and U5074 (N_5074,N_4497,N_4475);
nor U5075 (N_5075,N_4774,N_4554);
nor U5076 (N_5076,N_4678,N_4567);
and U5077 (N_5077,N_4126,N_4205);
nor U5078 (N_5078,N_4302,N_4739);
or U5079 (N_5079,N_4014,N_4117);
or U5080 (N_5080,N_4785,N_4357);
or U5081 (N_5081,N_4614,N_4435);
nand U5082 (N_5082,N_4558,N_4393);
nor U5083 (N_5083,N_4154,N_4735);
nand U5084 (N_5084,N_4138,N_4428);
nor U5085 (N_5085,N_4546,N_4630);
nand U5086 (N_5086,N_4573,N_4505);
and U5087 (N_5087,N_4134,N_4083);
nor U5088 (N_5088,N_4616,N_4095);
nor U5089 (N_5089,N_4309,N_4290);
or U5090 (N_5090,N_4723,N_4069);
nor U5091 (N_5091,N_4043,N_4364);
and U5092 (N_5092,N_4426,N_4407);
nand U5093 (N_5093,N_4137,N_4769);
nand U5094 (N_5094,N_4391,N_4596);
nor U5095 (N_5095,N_4236,N_4029);
and U5096 (N_5096,N_4568,N_4228);
xor U5097 (N_5097,N_4642,N_4104);
nor U5098 (N_5098,N_4049,N_4203);
xnor U5099 (N_5099,N_4416,N_4086);
and U5100 (N_5100,N_4305,N_4566);
nand U5101 (N_5101,N_4718,N_4465);
or U5102 (N_5102,N_4456,N_4346);
xnor U5103 (N_5103,N_4655,N_4023);
and U5104 (N_5104,N_4779,N_4261);
xnor U5105 (N_5105,N_4404,N_4598);
or U5106 (N_5106,N_4638,N_4091);
nand U5107 (N_5107,N_4304,N_4058);
or U5108 (N_5108,N_4611,N_4631);
and U5109 (N_5109,N_4128,N_4632);
or U5110 (N_5110,N_4715,N_4194);
nor U5111 (N_5111,N_4619,N_4010);
xnor U5112 (N_5112,N_4100,N_4307);
or U5113 (N_5113,N_4068,N_4605);
or U5114 (N_5114,N_4153,N_4298);
xnor U5115 (N_5115,N_4569,N_4586);
nand U5116 (N_5116,N_4308,N_4332);
or U5117 (N_5117,N_4651,N_4770);
and U5118 (N_5118,N_4329,N_4527);
nor U5119 (N_5119,N_4087,N_4386);
xnor U5120 (N_5120,N_4776,N_4766);
xor U5121 (N_5121,N_4473,N_4155);
nand U5122 (N_5122,N_4217,N_4717);
and U5123 (N_5123,N_4113,N_4322);
nor U5124 (N_5124,N_4778,N_4388);
nand U5125 (N_5125,N_4498,N_4034);
or U5126 (N_5126,N_4378,N_4624);
or U5127 (N_5127,N_4621,N_4157);
xnor U5128 (N_5128,N_4125,N_4629);
nor U5129 (N_5129,N_4771,N_4206);
or U5130 (N_5130,N_4067,N_4207);
or U5131 (N_5131,N_4503,N_4749);
nand U5132 (N_5132,N_4454,N_4728);
or U5133 (N_5133,N_4543,N_4415);
and U5134 (N_5134,N_4744,N_4303);
or U5135 (N_5135,N_4028,N_4537);
nand U5136 (N_5136,N_4466,N_4676);
nand U5137 (N_5137,N_4595,N_4704);
and U5138 (N_5138,N_4159,N_4287);
nor U5139 (N_5139,N_4133,N_4177);
or U5140 (N_5140,N_4001,N_4243);
nor U5141 (N_5141,N_4112,N_4502);
and U5142 (N_5142,N_4583,N_4652);
xnor U5143 (N_5143,N_4414,N_4063);
or U5144 (N_5144,N_4633,N_4186);
xor U5145 (N_5145,N_4499,N_4666);
xor U5146 (N_5146,N_4702,N_4786);
xnor U5147 (N_5147,N_4695,N_4071);
or U5148 (N_5148,N_4462,N_4559);
xnor U5149 (N_5149,N_4538,N_4799);
or U5150 (N_5150,N_4375,N_4545);
or U5151 (N_5151,N_4623,N_4080);
nor U5152 (N_5152,N_4151,N_4533);
and U5153 (N_5153,N_4214,N_4167);
xnor U5154 (N_5154,N_4376,N_4759);
and U5155 (N_5155,N_4700,N_4732);
xor U5156 (N_5156,N_4267,N_4119);
or U5157 (N_5157,N_4192,N_4085);
nor U5158 (N_5158,N_4705,N_4245);
nand U5159 (N_5159,N_4618,N_4127);
or U5160 (N_5160,N_4390,N_4789);
and U5161 (N_5161,N_4392,N_4556);
and U5162 (N_5162,N_4409,N_4684);
nand U5163 (N_5163,N_4374,N_4617);
nor U5164 (N_5164,N_4273,N_4118);
xnor U5165 (N_5165,N_4487,N_4691);
nand U5166 (N_5166,N_4152,N_4669);
nor U5167 (N_5167,N_4260,N_4093);
or U5168 (N_5168,N_4609,N_4679);
nor U5169 (N_5169,N_4191,N_4272);
and U5170 (N_5170,N_4259,N_4790);
xor U5171 (N_5171,N_4484,N_4012);
and U5172 (N_5172,N_4552,N_4232);
or U5173 (N_5173,N_4427,N_4198);
or U5174 (N_5174,N_4424,N_4433);
or U5175 (N_5175,N_4726,N_4549);
and U5176 (N_5176,N_4047,N_4493);
or U5177 (N_5177,N_4448,N_4019);
or U5178 (N_5178,N_4541,N_4640);
nand U5179 (N_5179,N_4751,N_4348);
and U5180 (N_5180,N_4469,N_4241);
nand U5181 (N_5181,N_4662,N_4747);
or U5182 (N_5182,N_4714,N_4612);
xor U5183 (N_5183,N_4581,N_4185);
or U5184 (N_5184,N_4641,N_4436);
or U5185 (N_5185,N_4563,N_4021);
nor U5186 (N_5186,N_4059,N_4210);
or U5187 (N_5187,N_4233,N_4525);
and U5188 (N_5188,N_4321,N_4660);
and U5189 (N_5189,N_4246,N_4410);
xor U5190 (N_5190,N_4142,N_4017);
or U5191 (N_5191,N_4654,N_4292);
nor U5192 (N_5192,N_4096,N_4350);
nand U5193 (N_5193,N_4004,N_4363);
xor U5194 (N_5194,N_4756,N_4015);
and U5195 (N_5195,N_4703,N_4278);
nor U5196 (N_5196,N_4111,N_4174);
xor U5197 (N_5197,N_4381,N_4193);
nand U5198 (N_5198,N_4530,N_4488);
and U5199 (N_5199,N_4765,N_4761);
or U5200 (N_5200,N_4518,N_4058);
and U5201 (N_5201,N_4465,N_4569);
nand U5202 (N_5202,N_4667,N_4643);
or U5203 (N_5203,N_4482,N_4363);
or U5204 (N_5204,N_4238,N_4544);
or U5205 (N_5205,N_4168,N_4448);
and U5206 (N_5206,N_4529,N_4620);
or U5207 (N_5207,N_4654,N_4581);
and U5208 (N_5208,N_4328,N_4794);
and U5209 (N_5209,N_4433,N_4722);
nand U5210 (N_5210,N_4243,N_4355);
xor U5211 (N_5211,N_4792,N_4327);
xnor U5212 (N_5212,N_4469,N_4269);
or U5213 (N_5213,N_4021,N_4131);
or U5214 (N_5214,N_4520,N_4643);
and U5215 (N_5215,N_4386,N_4504);
nor U5216 (N_5216,N_4086,N_4099);
nor U5217 (N_5217,N_4310,N_4379);
nand U5218 (N_5218,N_4015,N_4100);
or U5219 (N_5219,N_4589,N_4176);
xnor U5220 (N_5220,N_4385,N_4523);
or U5221 (N_5221,N_4353,N_4506);
and U5222 (N_5222,N_4581,N_4749);
or U5223 (N_5223,N_4419,N_4518);
and U5224 (N_5224,N_4703,N_4369);
xnor U5225 (N_5225,N_4788,N_4512);
and U5226 (N_5226,N_4247,N_4025);
nor U5227 (N_5227,N_4408,N_4510);
or U5228 (N_5228,N_4347,N_4603);
and U5229 (N_5229,N_4767,N_4556);
or U5230 (N_5230,N_4019,N_4107);
nand U5231 (N_5231,N_4372,N_4224);
nand U5232 (N_5232,N_4720,N_4060);
or U5233 (N_5233,N_4399,N_4203);
and U5234 (N_5234,N_4410,N_4679);
or U5235 (N_5235,N_4388,N_4094);
nand U5236 (N_5236,N_4171,N_4339);
and U5237 (N_5237,N_4789,N_4036);
and U5238 (N_5238,N_4575,N_4674);
xnor U5239 (N_5239,N_4703,N_4101);
and U5240 (N_5240,N_4543,N_4758);
xnor U5241 (N_5241,N_4788,N_4496);
and U5242 (N_5242,N_4287,N_4734);
nand U5243 (N_5243,N_4294,N_4536);
nand U5244 (N_5244,N_4507,N_4456);
and U5245 (N_5245,N_4421,N_4563);
or U5246 (N_5246,N_4042,N_4080);
and U5247 (N_5247,N_4261,N_4736);
nor U5248 (N_5248,N_4245,N_4558);
or U5249 (N_5249,N_4529,N_4337);
xnor U5250 (N_5250,N_4548,N_4274);
and U5251 (N_5251,N_4766,N_4382);
nand U5252 (N_5252,N_4515,N_4268);
or U5253 (N_5253,N_4676,N_4630);
nor U5254 (N_5254,N_4546,N_4368);
and U5255 (N_5255,N_4689,N_4551);
nor U5256 (N_5256,N_4531,N_4014);
and U5257 (N_5257,N_4750,N_4081);
xnor U5258 (N_5258,N_4208,N_4040);
and U5259 (N_5259,N_4123,N_4098);
or U5260 (N_5260,N_4337,N_4610);
or U5261 (N_5261,N_4287,N_4439);
xor U5262 (N_5262,N_4643,N_4579);
or U5263 (N_5263,N_4472,N_4462);
or U5264 (N_5264,N_4537,N_4235);
or U5265 (N_5265,N_4678,N_4717);
nor U5266 (N_5266,N_4371,N_4784);
nor U5267 (N_5267,N_4287,N_4150);
and U5268 (N_5268,N_4572,N_4033);
or U5269 (N_5269,N_4228,N_4697);
and U5270 (N_5270,N_4225,N_4617);
xnor U5271 (N_5271,N_4146,N_4359);
or U5272 (N_5272,N_4791,N_4339);
xor U5273 (N_5273,N_4234,N_4409);
nor U5274 (N_5274,N_4023,N_4182);
and U5275 (N_5275,N_4197,N_4417);
nand U5276 (N_5276,N_4229,N_4475);
and U5277 (N_5277,N_4796,N_4220);
nand U5278 (N_5278,N_4714,N_4445);
nor U5279 (N_5279,N_4327,N_4240);
and U5280 (N_5280,N_4729,N_4723);
or U5281 (N_5281,N_4046,N_4524);
and U5282 (N_5282,N_4361,N_4258);
nand U5283 (N_5283,N_4119,N_4445);
xor U5284 (N_5284,N_4228,N_4042);
nor U5285 (N_5285,N_4758,N_4485);
nand U5286 (N_5286,N_4217,N_4764);
xor U5287 (N_5287,N_4619,N_4684);
nand U5288 (N_5288,N_4048,N_4313);
xnor U5289 (N_5289,N_4696,N_4021);
nor U5290 (N_5290,N_4620,N_4214);
nor U5291 (N_5291,N_4556,N_4020);
nand U5292 (N_5292,N_4715,N_4655);
nor U5293 (N_5293,N_4247,N_4279);
xnor U5294 (N_5294,N_4736,N_4516);
nor U5295 (N_5295,N_4519,N_4232);
nand U5296 (N_5296,N_4476,N_4656);
nor U5297 (N_5297,N_4539,N_4144);
nor U5298 (N_5298,N_4308,N_4325);
nand U5299 (N_5299,N_4550,N_4788);
nor U5300 (N_5300,N_4065,N_4118);
or U5301 (N_5301,N_4409,N_4322);
nand U5302 (N_5302,N_4172,N_4114);
nor U5303 (N_5303,N_4687,N_4512);
and U5304 (N_5304,N_4776,N_4330);
nor U5305 (N_5305,N_4791,N_4026);
or U5306 (N_5306,N_4541,N_4424);
nand U5307 (N_5307,N_4449,N_4201);
and U5308 (N_5308,N_4572,N_4018);
nor U5309 (N_5309,N_4364,N_4734);
xor U5310 (N_5310,N_4196,N_4599);
or U5311 (N_5311,N_4143,N_4360);
nor U5312 (N_5312,N_4129,N_4462);
nand U5313 (N_5313,N_4402,N_4496);
nand U5314 (N_5314,N_4551,N_4397);
xnor U5315 (N_5315,N_4465,N_4087);
and U5316 (N_5316,N_4059,N_4406);
xnor U5317 (N_5317,N_4182,N_4316);
and U5318 (N_5318,N_4547,N_4209);
and U5319 (N_5319,N_4747,N_4087);
xor U5320 (N_5320,N_4430,N_4482);
and U5321 (N_5321,N_4228,N_4710);
nand U5322 (N_5322,N_4656,N_4740);
and U5323 (N_5323,N_4556,N_4765);
or U5324 (N_5324,N_4624,N_4499);
nor U5325 (N_5325,N_4145,N_4359);
nand U5326 (N_5326,N_4541,N_4540);
nand U5327 (N_5327,N_4672,N_4440);
and U5328 (N_5328,N_4675,N_4787);
nor U5329 (N_5329,N_4271,N_4695);
nor U5330 (N_5330,N_4292,N_4272);
and U5331 (N_5331,N_4448,N_4598);
nor U5332 (N_5332,N_4139,N_4574);
and U5333 (N_5333,N_4346,N_4698);
or U5334 (N_5334,N_4240,N_4098);
nor U5335 (N_5335,N_4151,N_4676);
nor U5336 (N_5336,N_4193,N_4496);
xor U5337 (N_5337,N_4758,N_4732);
or U5338 (N_5338,N_4009,N_4265);
or U5339 (N_5339,N_4342,N_4230);
and U5340 (N_5340,N_4540,N_4715);
nor U5341 (N_5341,N_4078,N_4306);
xnor U5342 (N_5342,N_4166,N_4243);
nand U5343 (N_5343,N_4362,N_4569);
nand U5344 (N_5344,N_4763,N_4697);
nor U5345 (N_5345,N_4127,N_4400);
nor U5346 (N_5346,N_4436,N_4039);
and U5347 (N_5347,N_4706,N_4797);
nand U5348 (N_5348,N_4209,N_4549);
nor U5349 (N_5349,N_4738,N_4003);
and U5350 (N_5350,N_4010,N_4312);
and U5351 (N_5351,N_4248,N_4076);
nor U5352 (N_5352,N_4314,N_4743);
nand U5353 (N_5353,N_4607,N_4725);
and U5354 (N_5354,N_4567,N_4538);
or U5355 (N_5355,N_4510,N_4538);
xnor U5356 (N_5356,N_4359,N_4604);
nor U5357 (N_5357,N_4419,N_4547);
or U5358 (N_5358,N_4018,N_4229);
nand U5359 (N_5359,N_4504,N_4047);
nor U5360 (N_5360,N_4504,N_4750);
nand U5361 (N_5361,N_4292,N_4315);
and U5362 (N_5362,N_4191,N_4160);
nand U5363 (N_5363,N_4189,N_4767);
xnor U5364 (N_5364,N_4475,N_4112);
or U5365 (N_5365,N_4237,N_4791);
and U5366 (N_5366,N_4075,N_4741);
xnor U5367 (N_5367,N_4276,N_4734);
xor U5368 (N_5368,N_4056,N_4634);
nor U5369 (N_5369,N_4084,N_4133);
and U5370 (N_5370,N_4116,N_4650);
or U5371 (N_5371,N_4052,N_4668);
xor U5372 (N_5372,N_4690,N_4261);
and U5373 (N_5373,N_4599,N_4200);
nand U5374 (N_5374,N_4645,N_4490);
xnor U5375 (N_5375,N_4495,N_4558);
nor U5376 (N_5376,N_4389,N_4214);
xnor U5377 (N_5377,N_4402,N_4314);
or U5378 (N_5378,N_4549,N_4773);
nand U5379 (N_5379,N_4541,N_4726);
or U5380 (N_5380,N_4222,N_4061);
and U5381 (N_5381,N_4225,N_4019);
nor U5382 (N_5382,N_4189,N_4333);
and U5383 (N_5383,N_4569,N_4731);
or U5384 (N_5384,N_4515,N_4066);
nand U5385 (N_5385,N_4528,N_4404);
nor U5386 (N_5386,N_4734,N_4356);
xor U5387 (N_5387,N_4751,N_4361);
xnor U5388 (N_5388,N_4382,N_4362);
nor U5389 (N_5389,N_4344,N_4458);
and U5390 (N_5390,N_4314,N_4129);
xor U5391 (N_5391,N_4748,N_4260);
nor U5392 (N_5392,N_4391,N_4281);
and U5393 (N_5393,N_4478,N_4238);
and U5394 (N_5394,N_4173,N_4164);
or U5395 (N_5395,N_4761,N_4316);
nor U5396 (N_5396,N_4693,N_4098);
or U5397 (N_5397,N_4336,N_4754);
and U5398 (N_5398,N_4130,N_4060);
and U5399 (N_5399,N_4102,N_4155);
and U5400 (N_5400,N_4157,N_4735);
nand U5401 (N_5401,N_4495,N_4487);
xor U5402 (N_5402,N_4133,N_4120);
and U5403 (N_5403,N_4376,N_4578);
or U5404 (N_5404,N_4390,N_4043);
nor U5405 (N_5405,N_4270,N_4701);
nor U5406 (N_5406,N_4274,N_4702);
nor U5407 (N_5407,N_4570,N_4294);
nand U5408 (N_5408,N_4503,N_4234);
nand U5409 (N_5409,N_4398,N_4632);
xnor U5410 (N_5410,N_4547,N_4195);
nor U5411 (N_5411,N_4360,N_4244);
and U5412 (N_5412,N_4332,N_4367);
xnor U5413 (N_5413,N_4573,N_4767);
or U5414 (N_5414,N_4653,N_4197);
and U5415 (N_5415,N_4403,N_4256);
xor U5416 (N_5416,N_4067,N_4402);
nor U5417 (N_5417,N_4586,N_4649);
and U5418 (N_5418,N_4249,N_4781);
nor U5419 (N_5419,N_4411,N_4284);
xnor U5420 (N_5420,N_4302,N_4170);
nand U5421 (N_5421,N_4214,N_4270);
and U5422 (N_5422,N_4058,N_4415);
nand U5423 (N_5423,N_4351,N_4655);
and U5424 (N_5424,N_4500,N_4545);
nor U5425 (N_5425,N_4025,N_4327);
nand U5426 (N_5426,N_4598,N_4624);
nor U5427 (N_5427,N_4576,N_4506);
or U5428 (N_5428,N_4189,N_4787);
or U5429 (N_5429,N_4397,N_4388);
or U5430 (N_5430,N_4584,N_4589);
nor U5431 (N_5431,N_4199,N_4475);
xnor U5432 (N_5432,N_4707,N_4121);
xnor U5433 (N_5433,N_4366,N_4092);
nor U5434 (N_5434,N_4699,N_4707);
xor U5435 (N_5435,N_4202,N_4274);
and U5436 (N_5436,N_4397,N_4079);
nor U5437 (N_5437,N_4688,N_4040);
xor U5438 (N_5438,N_4313,N_4194);
or U5439 (N_5439,N_4675,N_4043);
or U5440 (N_5440,N_4012,N_4396);
xor U5441 (N_5441,N_4710,N_4717);
or U5442 (N_5442,N_4402,N_4151);
nor U5443 (N_5443,N_4423,N_4663);
nand U5444 (N_5444,N_4155,N_4171);
nand U5445 (N_5445,N_4771,N_4613);
nand U5446 (N_5446,N_4529,N_4082);
and U5447 (N_5447,N_4311,N_4131);
and U5448 (N_5448,N_4380,N_4456);
xor U5449 (N_5449,N_4591,N_4734);
or U5450 (N_5450,N_4688,N_4326);
xnor U5451 (N_5451,N_4287,N_4142);
nand U5452 (N_5452,N_4434,N_4029);
or U5453 (N_5453,N_4430,N_4499);
and U5454 (N_5454,N_4315,N_4306);
xnor U5455 (N_5455,N_4661,N_4396);
xor U5456 (N_5456,N_4647,N_4481);
and U5457 (N_5457,N_4006,N_4280);
xor U5458 (N_5458,N_4259,N_4346);
and U5459 (N_5459,N_4442,N_4470);
or U5460 (N_5460,N_4454,N_4528);
nor U5461 (N_5461,N_4602,N_4698);
nor U5462 (N_5462,N_4149,N_4550);
nand U5463 (N_5463,N_4127,N_4129);
or U5464 (N_5464,N_4263,N_4566);
and U5465 (N_5465,N_4117,N_4169);
xor U5466 (N_5466,N_4788,N_4303);
nand U5467 (N_5467,N_4564,N_4568);
nor U5468 (N_5468,N_4312,N_4081);
and U5469 (N_5469,N_4534,N_4344);
and U5470 (N_5470,N_4790,N_4414);
and U5471 (N_5471,N_4140,N_4767);
or U5472 (N_5472,N_4165,N_4614);
xnor U5473 (N_5473,N_4606,N_4317);
nor U5474 (N_5474,N_4014,N_4347);
nand U5475 (N_5475,N_4714,N_4523);
xor U5476 (N_5476,N_4742,N_4445);
and U5477 (N_5477,N_4470,N_4608);
or U5478 (N_5478,N_4552,N_4725);
and U5479 (N_5479,N_4714,N_4399);
xor U5480 (N_5480,N_4194,N_4172);
nand U5481 (N_5481,N_4047,N_4063);
xnor U5482 (N_5482,N_4081,N_4093);
or U5483 (N_5483,N_4053,N_4373);
nor U5484 (N_5484,N_4653,N_4058);
nand U5485 (N_5485,N_4040,N_4442);
and U5486 (N_5486,N_4643,N_4763);
xor U5487 (N_5487,N_4066,N_4208);
nand U5488 (N_5488,N_4371,N_4428);
and U5489 (N_5489,N_4784,N_4286);
nand U5490 (N_5490,N_4709,N_4010);
nand U5491 (N_5491,N_4340,N_4593);
nand U5492 (N_5492,N_4421,N_4218);
and U5493 (N_5493,N_4614,N_4177);
nand U5494 (N_5494,N_4545,N_4415);
nand U5495 (N_5495,N_4194,N_4464);
nor U5496 (N_5496,N_4376,N_4299);
xnor U5497 (N_5497,N_4369,N_4379);
nand U5498 (N_5498,N_4170,N_4210);
or U5499 (N_5499,N_4023,N_4379);
or U5500 (N_5500,N_4540,N_4549);
nor U5501 (N_5501,N_4105,N_4754);
nand U5502 (N_5502,N_4010,N_4434);
and U5503 (N_5503,N_4290,N_4477);
nor U5504 (N_5504,N_4578,N_4043);
and U5505 (N_5505,N_4182,N_4603);
or U5506 (N_5506,N_4582,N_4419);
nand U5507 (N_5507,N_4128,N_4743);
or U5508 (N_5508,N_4266,N_4225);
nand U5509 (N_5509,N_4798,N_4185);
or U5510 (N_5510,N_4545,N_4094);
xor U5511 (N_5511,N_4289,N_4764);
and U5512 (N_5512,N_4489,N_4334);
or U5513 (N_5513,N_4529,N_4471);
or U5514 (N_5514,N_4233,N_4386);
nand U5515 (N_5515,N_4754,N_4109);
and U5516 (N_5516,N_4618,N_4192);
or U5517 (N_5517,N_4435,N_4034);
or U5518 (N_5518,N_4108,N_4663);
xor U5519 (N_5519,N_4207,N_4206);
or U5520 (N_5520,N_4532,N_4605);
and U5521 (N_5521,N_4129,N_4405);
or U5522 (N_5522,N_4030,N_4015);
nand U5523 (N_5523,N_4211,N_4503);
and U5524 (N_5524,N_4417,N_4201);
xnor U5525 (N_5525,N_4782,N_4033);
xor U5526 (N_5526,N_4503,N_4529);
xnor U5527 (N_5527,N_4303,N_4686);
or U5528 (N_5528,N_4045,N_4008);
nand U5529 (N_5529,N_4199,N_4732);
and U5530 (N_5530,N_4744,N_4025);
xnor U5531 (N_5531,N_4509,N_4389);
or U5532 (N_5532,N_4599,N_4544);
and U5533 (N_5533,N_4288,N_4061);
and U5534 (N_5534,N_4251,N_4106);
and U5535 (N_5535,N_4313,N_4758);
nor U5536 (N_5536,N_4379,N_4519);
and U5537 (N_5537,N_4161,N_4426);
xnor U5538 (N_5538,N_4324,N_4396);
or U5539 (N_5539,N_4184,N_4053);
nand U5540 (N_5540,N_4707,N_4155);
nand U5541 (N_5541,N_4063,N_4455);
or U5542 (N_5542,N_4248,N_4367);
nor U5543 (N_5543,N_4519,N_4321);
and U5544 (N_5544,N_4735,N_4708);
nand U5545 (N_5545,N_4437,N_4701);
or U5546 (N_5546,N_4720,N_4490);
nor U5547 (N_5547,N_4452,N_4108);
or U5548 (N_5548,N_4500,N_4400);
nor U5549 (N_5549,N_4750,N_4725);
xnor U5550 (N_5550,N_4796,N_4444);
and U5551 (N_5551,N_4171,N_4778);
xnor U5552 (N_5552,N_4595,N_4260);
nand U5553 (N_5553,N_4737,N_4643);
or U5554 (N_5554,N_4618,N_4767);
nor U5555 (N_5555,N_4004,N_4024);
nor U5556 (N_5556,N_4500,N_4409);
nor U5557 (N_5557,N_4442,N_4284);
and U5558 (N_5558,N_4526,N_4745);
nand U5559 (N_5559,N_4081,N_4229);
nand U5560 (N_5560,N_4759,N_4029);
or U5561 (N_5561,N_4541,N_4423);
or U5562 (N_5562,N_4056,N_4391);
or U5563 (N_5563,N_4020,N_4717);
xnor U5564 (N_5564,N_4234,N_4048);
or U5565 (N_5565,N_4754,N_4771);
xnor U5566 (N_5566,N_4470,N_4443);
or U5567 (N_5567,N_4322,N_4435);
xor U5568 (N_5568,N_4216,N_4493);
nor U5569 (N_5569,N_4284,N_4318);
or U5570 (N_5570,N_4341,N_4245);
xor U5571 (N_5571,N_4038,N_4502);
xor U5572 (N_5572,N_4130,N_4279);
xnor U5573 (N_5573,N_4105,N_4740);
nor U5574 (N_5574,N_4541,N_4769);
or U5575 (N_5575,N_4787,N_4371);
nand U5576 (N_5576,N_4595,N_4273);
and U5577 (N_5577,N_4224,N_4562);
nor U5578 (N_5578,N_4546,N_4355);
nor U5579 (N_5579,N_4216,N_4567);
and U5580 (N_5580,N_4079,N_4118);
xor U5581 (N_5581,N_4645,N_4733);
and U5582 (N_5582,N_4229,N_4679);
or U5583 (N_5583,N_4392,N_4488);
xnor U5584 (N_5584,N_4012,N_4665);
and U5585 (N_5585,N_4583,N_4772);
or U5586 (N_5586,N_4273,N_4675);
and U5587 (N_5587,N_4621,N_4487);
nand U5588 (N_5588,N_4220,N_4712);
and U5589 (N_5589,N_4192,N_4689);
nand U5590 (N_5590,N_4721,N_4024);
nand U5591 (N_5591,N_4759,N_4352);
xor U5592 (N_5592,N_4566,N_4548);
or U5593 (N_5593,N_4443,N_4392);
nor U5594 (N_5594,N_4302,N_4588);
nor U5595 (N_5595,N_4783,N_4175);
and U5596 (N_5596,N_4401,N_4793);
xnor U5597 (N_5597,N_4544,N_4173);
and U5598 (N_5598,N_4087,N_4304);
and U5599 (N_5599,N_4627,N_4377);
nand U5600 (N_5600,N_5297,N_5431);
or U5601 (N_5601,N_5099,N_5408);
or U5602 (N_5602,N_4804,N_5442);
xor U5603 (N_5603,N_5142,N_5109);
nand U5604 (N_5604,N_5256,N_5368);
xor U5605 (N_5605,N_5048,N_4876);
and U5606 (N_5606,N_4802,N_5140);
and U5607 (N_5607,N_5113,N_4921);
nand U5608 (N_5608,N_5001,N_5502);
nand U5609 (N_5609,N_5576,N_5088);
and U5610 (N_5610,N_5483,N_5588);
xor U5611 (N_5611,N_5147,N_5059);
nor U5612 (N_5612,N_5380,N_5374);
nor U5613 (N_5613,N_5568,N_5129);
nand U5614 (N_5614,N_5296,N_5375);
and U5615 (N_5615,N_5014,N_5314);
and U5616 (N_5616,N_5178,N_5053);
xor U5617 (N_5617,N_4912,N_5285);
nor U5618 (N_5618,N_5095,N_5172);
or U5619 (N_5619,N_5400,N_4978);
nor U5620 (N_5620,N_4894,N_5518);
nor U5621 (N_5621,N_5184,N_5016);
and U5622 (N_5622,N_5527,N_5039);
and U5623 (N_5623,N_5487,N_5533);
or U5624 (N_5624,N_4819,N_5355);
or U5625 (N_5625,N_4857,N_5191);
nand U5626 (N_5626,N_5254,N_4803);
or U5627 (N_5627,N_5412,N_5583);
nand U5628 (N_5628,N_5318,N_5156);
or U5629 (N_5629,N_4893,N_5501);
xor U5630 (N_5630,N_5248,N_4911);
nor U5631 (N_5631,N_5108,N_5343);
xnor U5632 (N_5632,N_4948,N_5584);
xor U5633 (N_5633,N_5271,N_5276);
nor U5634 (N_5634,N_5457,N_5510);
or U5635 (N_5635,N_4847,N_4868);
and U5636 (N_5636,N_4903,N_5460);
nand U5637 (N_5637,N_5553,N_5132);
nand U5638 (N_5638,N_5466,N_5174);
and U5639 (N_5639,N_5468,N_5305);
nand U5640 (N_5640,N_5078,N_5532);
or U5641 (N_5641,N_4913,N_5045);
or U5642 (N_5642,N_5133,N_5282);
xnor U5643 (N_5643,N_4964,N_5218);
and U5644 (N_5644,N_5371,N_5206);
nor U5645 (N_5645,N_5398,N_5511);
nand U5646 (N_5646,N_5308,N_4837);
or U5647 (N_5647,N_5428,N_5017);
or U5648 (N_5648,N_5278,N_5443);
xnor U5649 (N_5649,N_5395,N_5542);
xnor U5650 (N_5650,N_5420,N_5061);
or U5651 (N_5651,N_5433,N_5198);
nor U5652 (N_5652,N_4929,N_5090);
nor U5653 (N_5653,N_5111,N_4945);
and U5654 (N_5654,N_4997,N_5513);
or U5655 (N_5655,N_5138,N_4817);
nor U5656 (N_5656,N_5549,N_4914);
xor U5657 (N_5657,N_5484,N_5454);
xor U5658 (N_5658,N_5227,N_5223);
nand U5659 (N_5659,N_5042,N_4854);
xor U5660 (N_5660,N_5245,N_4952);
xor U5661 (N_5661,N_5103,N_5134);
and U5662 (N_5662,N_5348,N_4916);
or U5663 (N_5663,N_5264,N_5159);
or U5664 (N_5664,N_5357,N_5161);
nor U5665 (N_5665,N_5505,N_5382);
and U5666 (N_5666,N_4946,N_5535);
or U5667 (N_5667,N_4947,N_5360);
or U5668 (N_5668,N_5192,N_5366);
or U5669 (N_5669,N_5515,N_4985);
and U5670 (N_5670,N_5240,N_5224);
and U5671 (N_5671,N_5175,N_5266);
or U5672 (N_5672,N_4933,N_4966);
nor U5673 (N_5673,N_5087,N_4987);
or U5674 (N_5674,N_5350,N_5461);
nand U5675 (N_5675,N_5397,N_5038);
and U5676 (N_5676,N_5424,N_5509);
nand U5677 (N_5677,N_4930,N_5473);
xnor U5678 (N_5678,N_5300,N_5071);
nand U5679 (N_5679,N_5054,N_5169);
xnor U5680 (N_5680,N_5194,N_4951);
xor U5681 (N_5681,N_4905,N_4998);
nor U5682 (N_5682,N_5516,N_5196);
xnor U5683 (N_5683,N_5562,N_4994);
or U5684 (N_5684,N_5574,N_5345);
or U5685 (N_5685,N_5028,N_5330);
or U5686 (N_5686,N_5289,N_5149);
or U5687 (N_5687,N_5467,N_5389);
nor U5688 (N_5688,N_5047,N_4896);
nand U5689 (N_5689,N_5411,N_5586);
nor U5690 (N_5690,N_5521,N_5494);
or U5691 (N_5691,N_5367,N_5277);
or U5692 (N_5692,N_5065,N_5128);
or U5693 (N_5693,N_5274,N_5525);
or U5694 (N_5694,N_4969,N_5427);
xor U5695 (N_5695,N_5127,N_5321);
and U5696 (N_5696,N_5358,N_4836);
nor U5697 (N_5697,N_5066,N_5449);
xor U5698 (N_5698,N_5550,N_4939);
xor U5699 (N_5699,N_5244,N_5577);
or U5700 (N_5700,N_5101,N_5036);
nor U5701 (N_5701,N_4875,N_5592);
nand U5702 (N_5702,N_5417,N_5237);
or U5703 (N_5703,N_5440,N_4890);
nand U5704 (N_5704,N_5554,N_4897);
nor U5705 (N_5705,N_5552,N_5506);
and U5706 (N_5706,N_5165,N_5100);
nor U5707 (N_5707,N_5107,N_4928);
and U5708 (N_5708,N_5137,N_5205);
and U5709 (N_5709,N_4919,N_4891);
or U5710 (N_5710,N_4850,N_5004);
nand U5711 (N_5711,N_5148,N_4956);
xnor U5712 (N_5712,N_5136,N_5067);
or U5713 (N_5713,N_4965,N_4865);
and U5714 (N_5714,N_5311,N_5563);
and U5715 (N_5715,N_5476,N_5465);
nor U5716 (N_5716,N_5164,N_5176);
or U5717 (N_5717,N_5182,N_5011);
xnor U5718 (N_5718,N_5226,N_5037);
xnor U5719 (N_5719,N_5558,N_4927);
and U5720 (N_5720,N_5019,N_4887);
or U5721 (N_5721,N_5210,N_5519);
and U5722 (N_5722,N_5504,N_4967);
nand U5723 (N_5723,N_5364,N_5410);
or U5724 (N_5724,N_5421,N_5503);
xor U5725 (N_5725,N_5450,N_5064);
or U5726 (N_5726,N_5597,N_4990);
nor U5727 (N_5727,N_5183,N_5288);
or U5728 (N_5728,N_5415,N_5168);
or U5729 (N_5729,N_5233,N_5596);
nand U5730 (N_5730,N_5263,N_4885);
nand U5731 (N_5731,N_4839,N_5005);
and U5732 (N_5732,N_5195,N_5204);
xnor U5733 (N_5733,N_5073,N_4950);
or U5734 (N_5734,N_5270,N_4949);
nand U5735 (N_5735,N_5238,N_5582);
nor U5736 (N_5736,N_5560,N_5377);
nand U5737 (N_5737,N_5075,N_4938);
nand U5738 (N_5738,N_5426,N_5339);
nand U5739 (N_5739,N_5546,N_5040);
nor U5740 (N_5740,N_4832,N_5021);
and U5741 (N_5741,N_5219,N_5098);
nand U5742 (N_5742,N_4859,N_5524);
nand U5743 (N_5743,N_5072,N_4879);
xor U5744 (N_5744,N_4892,N_5215);
nand U5745 (N_5745,N_5225,N_5260);
xor U5746 (N_5746,N_5080,N_4811);
nand U5747 (N_5747,N_5081,N_4871);
nand U5748 (N_5748,N_4920,N_5403);
and U5749 (N_5749,N_5447,N_5301);
nor U5750 (N_5750,N_5097,N_5077);
and U5751 (N_5751,N_4909,N_4867);
nand U5752 (N_5752,N_5253,N_5069);
or U5753 (N_5753,N_5146,N_4861);
nor U5754 (N_5754,N_5230,N_5453);
or U5755 (N_5755,N_5200,N_5145);
and U5756 (N_5756,N_5153,N_4813);
or U5757 (N_5757,N_5268,N_5291);
nor U5758 (N_5758,N_5435,N_5203);
nor U5759 (N_5759,N_5482,N_5528);
nor U5760 (N_5760,N_5262,N_5572);
and U5761 (N_5761,N_5056,N_4915);
and U5762 (N_5762,N_5459,N_4808);
xor U5763 (N_5763,N_5273,N_4821);
and U5764 (N_5764,N_5376,N_4878);
xor U5765 (N_5765,N_4958,N_4801);
or U5766 (N_5766,N_5458,N_5394);
nand U5767 (N_5767,N_5413,N_5561);
nand U5768 (N_5768,N_5488,N_5327);
xnor U5769 (N_5769,N_4999,N_5386);
or U5770 (N_5770,N_5115,N_4848);
and U5771 (N_5771,N_5439,N_5236);
nor U5772 (N_5772,N_4959,N_5281);
nand U5773 (N_5773,N_5250,N_5315);
and U5774 (N_5774,N_4873,N_4849);
nor U5775 (N_5775,N_5547,N_5463);
nor U5776 (N_5776,N_4979,N_5030);
nand U5777 (N_5777,N_5393,N_4851);
and U5778 (N_5778,N_5312,N_4858);
or U5779 (N_5779,N_5143,N_5406);
or U5780 (N_5780,N_5177,N_5020);
or U5781 (N_5781,N_5006,N_5340);
xor U5782 (N_5782,N_5157,N_4902);
xnor U5783 (N_5783,N_5462,N_5418);
xor U5784 (N_5784,N_5022,N_4968);
xnor U5785 (N_5785,N_5373,N_5491);
nand U5786 (N_5786,N_5079,N_5571);
or U5787 (N_5787,N_4953,N_5261);
or U5788 (N_5788,N_5565,N_4828);
or U5789 (N_5789,N_4826,N_4976);
xnor U5790 (N_5790,N_4869,N_5013);
and U5791 (N_5791,N_5500,N_5163);
and U5792 (N_5792,N_5049,N_4842);
or U5793 (N_5793,N_4863,N_5493);
or U5794 (N_5794,N_5388,N_5379);
nand U5795 (N_5795,N_5593,N_4936);
xnor U5796 (N_5796,N_4844,N_5492);
xnor U5797 (N_5797,N_5529,N_5255);
xor U5798 (N_5798,N_5122,N_5384);
or U5799 (N_5799,N_4957,N_5117);
xnor U5800 (N_5800,N_5520,N_5573);
xnor U5801 (N_5801,N_5279,N_5259);
nand U5802 (N_5802,N_4922,N_4996);
nor U5803 (N_5803,N_4810,N_5402);
nand U5804 (N_5804,N_4941,N_5027);
or U5805 (N_5805,N_5396,N_5119);
xnor U5806 (N_5806,N_5243,N_4822);
nor U5807 (N_5807,N_4841,N_5414);
xnor U5808 (N_5808,N_5008,N_5540);
nor U5809 (N_5809,N_5180,N_4977);
and U5810 (N_5810,N_5474,N_5155);
or U5811 (N_5811,N_5302,N_5246);
nor U5812 (N_5812,N_4931,N_4809);
and U5813 (N_5813,N_5580,N_5187);
xnor U5814 (N_5814,N_5213,N_5385);
and U5815 (N_5815,N_4831,N_4983);
xor U5816 (N_5816,N_5057,N_5123);
and U5817 (N_5817,N_4899,N_5526);
xor U5818 (N_5818,N_5570,N_4824);
xor U5819 (N_5819,N_5190,N_5472);
or U5820 (N_5820,N_5082,N_5110);
or U5821 (N_5821,N_5283,N_5211);
nand U5822 (N_5822,N_5370,N_5106);
nor U5823 (N_5823,N_5171,N_5423);
nor U5824 (N_5824,N_5430,N_5247);
nor U5825 (N_5825,N_4989,N_5114);
and U5826 (N_5826,N_5104,N_4963);
nor U5827 (N_5827,N_5197,N_4888);
and U5828 (N_5828,N_5102,N_5383);
nand U5829 (N_5829,N_4818,N_5217);
and U5830 (N_5830,N_5130,N_5295);
nor U5831 (N_5831,N_5490,N_5112);
xnor U5832 (N_5832,N_5092,N_4815);
and U5833 (N_5833,N_4940,N_5307);
and U5834 (N_5834,N_5131,N_4935);
and U5835 (N_5835,N_4960,N_5257);
or U5836 (N_5836,N_4971,N_4838);
xnor U5837 (N_5837,N_5162,N_5337);
nand U5838 (N_5838,N_5335,N_5316);
nand U5839 (N_5839,N_4800,N_5452);
and U5840 (N_5840,N_5025,N_5076);
xor U5841 (N_5841,N_4970,N_5578);
nand U5842 (N_5842,N_4812,N_5507);
and U5843 (N_5843,N_5508,N_5514);
nor U5844 (N_5844,N_5352,N_5498);
and U5845 (N_5845,N_5585,N_5589);
xnor U5846 (N_5846,N_5293,N_5438);
nand U5847 (N_5847,N_4923,N_4955);
or U5848 (N_5848,N_5170,N_5336);
nor U5849 (N_5849,N_5361,N_5326);
or U5850 (N_5850,N_5555,N_4986);
nand U5851 (N_5851,N_5551,N_5479);
and U5852 (N_5852,N_4973,N_5416);
nor U5853 (N_5853,N_5369,N_5023);
xor U5854 (N_5854,N_4907,N_4827);
xor U5855 (N_5855,N_5405,N_5126);
xnor U5856 (N_5856,N_5407,N_4910);
xor U5857 (N_5857,N_5587,N_4884);
xnor U5858 (N_5858,N_5419,N_5325);
or U5859 (N_5859,N_4925,N_5029);
or U5860 (N_5860,N_5242,N_5046);
and U5861 (N_5861,N_5455,N_5135);
nand U5862 (N_5862,N_5160,N_4877);
and U5863 (N_5863,N_5425,N_5310);
xor U5864 (N_5864,N_4908,N_5002);
nor U5865 (N_5865,N_5286,N_5309);
and U5866 (N_5866,N_4883,N_5537);
nand U5867 (N_5867,N_5456,N_4856);
and U5868 (N_5868,N_5522,N_5322);
and U5869 (N_5869,N_5469,N_4870);
and U5870 (N_5870,N_4981,N_4843);
or U5871 (N_5871,N_5347,N_4834);
nand U5872 (N_5872,N_5342,N_5470);
xnor U5873 (N_5873,N_5530,N_5151);
nor U5874 (N_5874,N_5249,N_5432);
nor U5875 (N_5875,N_4805,N_4932);
xor U5876 (N_5876,N_4904,N_5185);
nand U5877 (N_5877,N_5313,N_5018);
nor U5878 (N_5878,N_4982,N_5298);
or U5879 (N_5879,N_5284,N_5207);
and U5880 (N_5880,N_4874,N_5003);
nor U5881 (N_5881,N_5141,N_5575);
nor U5882 (N_5882,N_5173,N_5269);
xnor U5883 (N_5883,N_5579,N_5331);
and U5884 (N_5884,N_5486,N_4974);
or U5885 (N_5885,N_5334,N_5139);
xnor U5886 (N_5886,N_5272,N_5085);
nor U5887 (N_5887,N_5362,N_5392);
nand U5888 (N_5888,N_5186,N_5303);
or U5889 (N_5889,N_4961,N_4825);
and U5890 (N_5890,N_5598,N_4901);
and U5891 (N_5891,N_4820,N_4823);
or U5892 (N_5892,N_5445,N_5328);
or U5893 (N_5893,N_5280,N_5323);
nand U5894 (N_5894,N_5105,N_5356);
or U5895 (N_5895,N_5485,N_5199);
and U5896 (N_5896,N_5566,N_5595);
and U5897 (N_5897,N_5089,N_5010);
or U5898 (N_5898,N_5338,N_5222);
xor U5899 (N_5899,N_5094,N_5294);
or U5900 (N_5900,N_5031,N_5209);
or U5901 (N_5901,N_5118,N_5399);
and U5902 (N_5902,N_4918,N_5446);
or U5903 (N_5903,N_5252,N_4840);
or U5904 (N_5904,N_5234,N_5034);
nor U5905 (N_5905,N_5074,N_5341);
or U5906 (N_5906,N_4917,N_5032);
nor U5907 (N_5907,N_4835,N_5409);
nand U5908 (N_5908,N_5543,N_5292);
nand U5909 (N_5909,N_4855,N_5556);
or U5910 (N_5910,N_4937,N_5068);
xnor U5911 (N_5911,N_5070,N_4906);
or U5912 (N_5912,N_4860,N_5480);
xnor U5913 (N_5913,N_5451,N_5523);
xnor U5914 (N_5914,N_5591,N_5363);
or U5915 (N_5915,N_5332,N_4814);
nand U5916 (N_5916,N_4880,N_5544);
or U5917 (N_5917,N_5471,N_5599);
or U5918 (N_5918,N_5567,N_4926);
or U5919 (N_5919,N_5035,N_4872);
xor U5920 (N_5920,N_5317,N_5306);
or U5921 (N_5921,N_5512,N_5232);
or U5922 (N_5922,N_5381,N_5120);
or U5923 (N_5923,N_5365,N_5091);
and U5924 (N_5924,N_5026,N_5181);
nand U5925 (N_5925,N_5541,N_5116);
nand U5926 (N_5926,N_5083,N_5378);
nor U5927 (N_5927,N_4829,N_4852);
nand U5928 (N_5928,N_5436,N_5346);
nand U5929 (N_5929,N_4830,N_4954);
and U5930 (N_5930,N_4984,N_5324);
xnor U5931 (N_5931,N_5050,N_5559);
and U5932 (N_5932,N_4807,N_5096);
xnor U5933 (N_5933,N_5290,N_5124);
or U5934 (N_5934,N_5214,N_4816);
nor U5935 (N_5935,N_5007,N_5349);
or U5936 (N_5936,N_5539,N_4862);
and U5937 (N_5937,N_5429,N_5201);
or U5938 (N_5938,N_5545,N_5287);
nand U5939 (N_5939,N_5202,N_4898);
and U5940 (N_5940,N_4895,N_5564);
nand U5941 (N_5941,N_5189,N_4943);
and U5942 (N_5942,N_5043,N_5499);
or U5943 (N_5943,N_5536,N_5216);
and U5944 (N_5944,N_5320,N_5058);
nand U5945 (N_5945,N_5265,N_5251);
nor U5946 (N_5946,N_5534,N_5354);
or U5947 (N_5947,N_5372,N_5000);
xor U5948 (N_5948,N_5275,N_5391);
nor U5949 (N_5949,N_4972,N_5212);
or U5950 (N_5950,N_5084,N_5193);
nor U5951 (N_5951,N_5179,N_5024);
or U5952 (N_5952,N_5319,N_4889);
nand U5953 (N_5953,N_5052,N_5569);
nand U5954 (N_5954,N_5051,N_5166);
xor U5955 (N_5955,N_5538,N_5229);
nor U5956 (N_5956,N_5033,N_5154);
nand U5957 (N_5957,N_5437,N_5329);
or U5958 (N_5958,N_5060,N_5144);
and U5959 (N_5959,N_5359,N_4980);
nor U5960 (N_5960,N_5581,N_5009);
or U5961 (N_5961,N_5041,N_5448);
and U5962 (N_5962,N_5220,N_4924);
and U5963 (N_5963,N_4853,N_4881);
or U5964 (N_5964,N_5012,N_5158);
or U5965 (N_5965,N_4934,N_5444);
and U5966 (N_5966,N_4833,N_5333);
and U5967 (N_5967,N_5167,N_4866);
nand U5968 (N_5968,N_5228,N_4991);
xor U5969 (N_5969,N_4846,N_5422);
xnor U5970 (N_5970,N_5344,N_5496);
nor U5971 (N_5971,N_4975,N_5478);
or U5972 (N_5972,N_5152,N_5188);
and U5973 (N_5973,N_4944,N_5304);
or U5974 (N_5974,N_5231,N_4806);
xor U5975 (N_5975,N_5125,N_5401);
or U5976 (N_5976,N_5351,N_5477);
or U5977 (N_5977,N_5548,N_5241);
nand U5978 (N_5978,N_4995,N_4864);
nand U5979 (N_5979,N_5235,N_5221);
or U5980 (N_5980,N_5062,N_5441);
nand U5981 (N_5981,N_5055,N_5489);
nor U5982 (N_5982,N_5208,N_4993);
xor U5983 (N_5983,N_5015,N_5475);
or U5984 (N_5984,N_5434,N_4992);
and U5985 (N_5985,N_4886,N_4845);
nand U5986 (N_5986,N_5390,N_5086);
and U5987 (N_5987,N_5239,N_5044);
nor U5988 (N_5988,N_5387,N_5093);
nor U5989 (N_5989,N_5517,N_5497);
nand U5990 (N_5990,N_5590,N_5495);
and U5991 (N_5991,N_5150,N_4988);
nor U5992 (N_5992,N_5404,N_4962);
nand U5993 (N_5993,N_5464,N_5063);
and U5994 (N_5994,N_4900,N_4882);
nand U5995 (N_5995,N_5258,N_5531);
nand U5996 (N_5996,N_5299,N_5481);
nand U5997 (N_5997,N_4942,N_5121);
xnor U5998 (N_5998,N_5557,N_5267);
nand U5999 (N_5999,N_5594,N_5353);
nand U6000 (N_6000,N_5542,N_5034);
nor U6001 (N_6001,N_5346,N_5000);
or U6002 (N_6002,N_5297,N_5461);
nor U6003 (N_6003,N_5504,N_5432);
and U6004 (N_6004,N_5111,N_5021);
nor U6005 (N_6005,N_5347,N_5462);
nand U6006 (N_6006,N_4864,N_5532);
and U6007 (N_6007,N_5414,N_5506);
xnor U6008 (N_6008,N_5458,N_5452);
nand U6009 (N_6009,N_5350,N_5082);
nor U6010 (N_6010,N_5445,N_5538);
xnor U6011 (N_6011,N_5589,N_5211);
and U6012 (N_6012,N_5205,N_5357);
xnor U6013 (N_6013,N_4909,N_5495);
or U6014 (N_6014,N_5224,N_5512);
nand U6015 (N_6015,N_4847,N_4844);
and U6016 (N_6016,N_4951,N_4970);
and U6017 (N_6017,N_5134,N_4999);
nor U6018 (N_6018,N_5565,N_5361);
and U6019 (N_6019,N_5386,N_5232);
xor U6020 (N_6020,N_4809,N_5276);
xnor U6021 (N_6021,N_4823,N_4846);
and U6022 (N_6022,N_5288,N_5588);
or U6023 (N_6023,N_4806,N_5109);
or U6024 (N_6024,N_5236,N_5419);
and U6025 (N_6025,N_4937,N_5432);
xor U6026 (N_6026,N_5009,N_5249);
nor U6027 (N_6027,N_5268,N_4826);
nor U6028 (N_6028,N_5097,N_4986);
nor U6029 (N_6029,N_4931,N_5123);
xnor U6030 (N_6030,N_5166,N_4843);
xor U6031 (N_6031,N_4871,N_4979);
xor U6032 (N_6032,N_4921,N_4952);
xnor U6033 (N_6033,N_5555,N_4922);
and U6034 (N_6034,N_5545,N_5350);
or U6035 (N_6035,N_4872,N_5388);
xnor U6036 (N_6036,N_5183,N_4988);
and U6037 (N_6037,N_5095,N_5467);
nor U6038 (N_6038,N_5335,N_5204);
or U6039 (N_6039,N_5133,N_5550);
nand U6040 (N_6040,N_4984,N_5297);
nand U6041 (N_6041,N_4868,N_5553);
nor U6042 (N_6042,N_5485,N_5111);
or U6043 (N_6043,N_4810,N_5283);
and U6044 (N_6044,N_5352,N_4970);
or U6045 (N_6045,N_5447,N_5302);
and U6046 (N_6046,N_5178,N_5005);
nand U6047 (N_6047,N_4977,N_5404);
nor U6048 (N_6048,N_4981,N_5411);
nand U6049 (N_6049,N_5265,N_5591);
nand U6050 (N_6050,N_5291,N_5167);
and U6051 (N_6051,N_4832,N_5552);
and U6052 (N_6052,N_5511,N_5074);
xnor U6053 (N_6053,N_5029,N_4920);
nor U6054 (N_6054,N_5549,N_5143);
and U6055 (N_6055,N_5353,N_5381);
xor U6056 (N_6056,N_5022,N_5142);
and U6057 (N_6057,N_5392,N_4828);
nand U6058 (N_6058,N_5598,N_4909);
or U6059 (N_6059,N_4968,N_5079);
nor U6060 (N_6060,N_5073,N_5213);
nand U6061 (N_6061,N_5165,N_5291);
xor U6062 (N_6062,N_5331,N_5090);
xor U6063 (N_6063,N_5020,N_5252);
and U6064 (N_6064,N_5195,N_4911);
nand U6065 (N_6065,N_5568,N_5217);
nor U6066 (N_6066,N_5335,N_5065);
nand U6067 (N_6067,N_5269,N_5389);
and U6068 (N_6068,N_5113,N_4836);
nor U6069 (N_6069,N_5548,N_4928);
nor U6070 (N_6070,N_5185,N_5558);
xnor U6071 (N_6071,N_5521,N_5560);
or U6072 (N_6072,N_5569,N_5574);
and U6073 (N_6073,N_5561,N_4937);
and U6074 (N_6074,N_5156,N_5464);
or U6075 (N_6075,N_5001,N_5386);
or U6076 (N_6076,N_5475,N_4858);
nor U6077 (N_6077,N_5159,N_5546);
xor U6078 (N_6078,N_4808,N_5417);
or U6079 (N_6079,N_5059,N_5142);
or U6080 (N_6080,N_4939,N_5523);
nand U6081 (N_6081,N_5236,N_5579);
nor U6082 (N_6082,N_5439,N_4932);
xor U6083 (N_6083,N_5285,N_5298);
nand U6084 (N_6084,N_5327,N_5405);
and U6085 (N_6085,N_5020,N_5142);
nand U6086 (N_6086,N_4966,N_5276);
nor U6087 (N_6087,N_4945,N_5316);
xor U6088 (N_6088,N_5592,N_5485);
nand U6089 (N_6089,N_4903,N_4817);
and U6090 (N_6090,N_5073,N_5520);
nor U6091 (N_6091,N_5333,N_5184);
and U6092 (N_6092,N_5259,N_4930);
xor U6093 (N_6093,N_4802,N_4826);
nor U6094 (N_6094,N_5542,N_4860);
xnor U6095 (N_6095,N_5020,N_5488);
nor U6096 (N_6096,N_4938,N_5592);
and U6097 (N_6097,N_5275,N_5363);
or U6098 (N_6098,N_5189,N_5019);
nand U6099 (N_6099,N_5441,N_4886);
nand U6100 (N_6100,N_4849,N_4857);
nor U6101 (N_6101,N_5013,N_4851);
and U6102 (N_6102,N_4860,N_5478);
xor U6103 (N_6103,N_5208,N_4833);
and U6104 (N_6104,N_4995,N_4971);
and U6105 (N_6105,N_5330,N_5250);
or U6106 (N_6106,N_5106,N_5534);
or U6107 (N_6107,N_5151,N_5294);
or U6108 (N_6108,N_5219,N_5124);
nor U6109 (N_6109,N_5302,N_5448);
nor U6110 (N_6110,N_5357,N_4909);
or U6111 (N_6111,N_5474,N_5087);
or U6112 (N_6112,N_4885,N_5052);
xnor U6113 (N_6113,N_5477,N_5445);
nand U6114 (N_6114,N_4906,N_4927);
nor U6115 (N_6115,N_4861,N_5216);
nor U6116 (N_6116,N_4848,N_5212);
nor U6117 (N_6117,N_4892,N_4979);
nand U6118 (N_6118,N_5422,N_5489);
nor U6119 (N_6119,N_5589,N_5060);
and U6120 (N_6120,N_5094,N_5384);
and U6121 (N_6121,N_5370,N_5277);
nor U6122 (N_6122,N_5199,N_4965);
nand U6123 (N_6123,N_5467,N_5149);
nand U6124 (N_6124,N_5500,N_5358);
nand U6125 (N_6125,N_5343,N_4922);
and U6126 (N_6126,N_4924,N_5393);
and U6127 (N_6127,N_5377,N_4946);
nor U6128 (N_6128,N_5099,N_5507);
or U6129 (N_6129,N_5298,N_5396);
xnor U6130 (N_6130,N_4910,N_4844);
xnor U6131 (N_6131,N_4869,N_5492);
nand U6132 (N_6132,N_5096,N_5449);
or U6133 (N_6133,N_5012,N_5515);
or U6134 (N_6134,N_5214,N_4960);
and U6135 (N_6135,N_5178,N_5513);
nor U6136 (N_6136,N_5326,N_5042);
nand U6137 (N_6137,N_5068,N_5537);
and U6138 (N_6138,N_4920,N_5022);
nand U6139 (N_6139,N_5065,N_4801);
nand U6140 (N_6140,N_4982,N_5384);
and U6141 (N_6141,N_5121,N_4845);
and U6142 (N_6142,N_5572,N_4962);
nand U6143 (N_6143,N_5267,N_4977);
and U6144 (N_6144,N_5374,N_5016);
and U6145 (N_6145,N_5229,N_5124);
and U6146 (N_6146,N_5152,N_5473);
and U6147 (N_6147,N_4834,N_4962);
and U6148 (N_6148,N_4891,N_5002);
and U6149 (N_6149,N_5115,N_5102);
xnor U6150 (N_6150,N_5432,N_5122);
xor U6151 (N_6151,N_5426,N_5414);
nor U6152 (N_6152,N_5304,N_5513);
or U6153 (N_6153,N_5295,N_4885);
or U6154 (N_6154,N_5421,N_5297);
nor U6155 (N_6155,N_4831,N_5236);
and U6156 (N_6156,N_4867,N_5442);
nor U6157 (N_6157,N_5058,N_5382);
and U6158 (N_6158,N_4997,N_5126);
nor U6159 (N_6159,N_5598,N_5471);
or U6160 (N_6160,N_5516,N_4939);
xor U6161 (N_6161,N_4929,N_5094);
nor U6162 (N_6162,N_4951,N_5514);
nor U6163 (N_6163,N_5574,N_5210);
nor U6164 (N_6164,N_5265,N_4837);
and U6165 (N_6165,N_5499,N_5310);
or U6166 (N_6166,N_5276,N_5456);
nand U6167 (N_6167,N_5351,N_5085);
and U6168 (N_6168,N_4897,N_5445);
or U6169 (N_6169,N_4954,N_5504);
and U6170 (N_6170,N_5150,N_5492);
nor U6171 (N_6171,N_5488,N_5338);
nor U6172 (N_6172,N_5214,N_4907);
and U6173 (N_6173,N_5016,N_5489);
and U6174 (N_6174,N_5020,N_4953);
nor U6175 (N_6175,N_4804,N_5387);
nor U6176 (N_6176,N_5204,N_4827);
xnor U6177 (N_6177,N_5101,N_4970);
and U6178 (N_6178,N_5538,N_4840);
nand U6179 (N_6179,N_5550,N_5555);
or U6180 (N_6180,N_5301,N_5531);
xor U6181 (N_6181,N_5595,N_5174);
nand U6182 (N_6182,N_4861,N_5189);
and U6183 (N_6183,N_5193,N_5443);
nor U6184 (N_6184,N_5411,N_4901);
nor U6185 (N_6185,N_5069,N_4934);
nor U6186 (N_6186,N_5031,N_4950);
and U6187 (N_6187,N_5121,N_5218);
xor U6188 (N_6188,N_4921,N_4806);
and U6189 (N_6189,N_5498,N_5487);
nand U6190 (N_6190,N_4865,N_5379);
and U6191 (N_6191,N_5551,N_5456);
or U6192 (N_6192,N_5173,N_5224);
xnor U6193 (N_6193,N_4925,N_5161);
nor U6194 (N_6194,N_5197,N_5380);
and U6195 (N_6195,N_4969,N_5019);
or U6196 (N_6196,N_5178,N_5426);
nand U6197 (N_6197,N_5358,N_5266);
xor U6198 (N_6198,N_5432,N_5586);
nand U6199 (N_6199,N_5219,N_5022);
nor U6200 (N_6200,N_5341,N_5060);
and U6201 (N_6201,N_5268,N_5366);
xor U6202 (N_6202,N_4898,N_4943);
xnor U6203 (N_6203,N_5089,N_5009);
or U6204 (N_6204,N_5252,N_5547);
and U6205 (N_6205,N_5451,N_5378);
nor U6206 (N_6206,N_4822,N_5153);
nand U6207 (N_6207,N_5259,N_5554);
nand U6208 (N_6208,N_5439,N_4996);
nor U6209 (N_6209,N_5250,N_4850);
nand U6210 (N_6210,N_4900,N_5030);
nor U6211 (N_6211,N_5306,N_5107);
xor U6212 (N_6212,N_5478,N_5084);
xnor U6213 (N_6213,N_5101,N_5044);
xnor U6214 (N_6214,N_5319,N_5499);
or U6215 (N_6215,N_5594,N_5167);
xnor U6216 (N_6216,N_5327,N_5430);
or U6217 (N_6217,N_5263,N_5285);
nor U6218 (N_6218,N_5073,N_5294);
xor U6219 (N_6219,N_4869,N_4848);
nor U6220 (N_6220,N_5461,N_5049);
xor U6221 (N_6221,N_4875,N_5327);
and U6222 (N_6222,N_4878,N_5579);
and U6223 (N_6223,N_5297,N_5468);
xnor U6224 (N_6224,N_5513,N_5172);
nand U6225 (N_6225,N_5455,N_4895);
xor U6226 (N_6226,N_5382,N_4958);
xor U6227 (N_6227,N_5489,N_5007);
nand U6228 (N_6228,N_5117,N_5423);
and U6229 (N_6229,N_5488,N_4924);
and U6230 (N_6230,N_5163,N_4826);
nor U6231 (N_6231,N_5248,N_5288);
nor U6232 (N_6232,N_4938,N_4941);
xor U6233 (N_6233,N_5517,N_5479);
nor U6234 (N_6234,N_5128,N_5429);
xor U6235 (N_6235,N_5281,N_4978);
xnor U6236 (N_6236,N_5022,N_5414);
nand U6237 (N_6237,N_5025,N_5540);
and U6238 (N_6238,N_5494,N_5389);
or U6239 (N_6239,N_4943,N_5412);
nand U6240 (N_6240,N_4982,N_4862);
or U6241 (N_6241,N_5533,N_4855);
and U6242 (N_6242,N_4964,N_5472);
or U6243 (N_6243,N_5338,N_5412);
xnor U6244 (N_6244,N_5401,N_5156);
nor U6245 (N_6245,N_5312,N_5363);
or U6246 (N_6246,N_5055,N_5135);
xor U6247 (N_6247,N_5247,N_5292);
nor U6248 (N_6248,N_5219,N_5388);
nand U6249 (N_6249,N_5222,N_4846);
and U6250 (N_6250,N_5062,N_4994);
or U6251 (N_6251,N_5082,N_4809);
xnor U6252 (N_6252,N_5381,N_5478);
nor U6253 (N_6253,N_5080,N_4964);
or U6254 (N_6254,N_5002,N_4923);
nor U6255 (N_6255,N_5467,N_5195);
nor U6256 (N_6256,N_5114,N_5131);
or U6257 (N_6257,N_5112,N_5147);
nor U6258 (N_6258,N_5546,N_5192);
nor U6259 (N_6259,N_4931,N_4949);
nor U6260 (N_6260,N_4804,N_4892);
nand U6261 (N_6261,N_5559,N_4897);
or U6262 (N_6262,N_5170,N_4852);
or U6263 (N_6263,N_5538,N_5330);
nand U6264 (N_6264,N_5004,N_5083);
xor U6265 (N_6265,N_5447,N_5487);
or U6266 (N_6266,N_4902,N_4917);
and U6267 (N_6267,N_4826,N_5028);
nand U6268 (N_6268,N_5450,N_5492);
or U6269 (N_6269,N_5301,N_5425);
nand U6270 (N_6270,N_5257,N_5272);
xnor U6271 (N_6271,N_5440,N_5011);
and U6272 (N_6272,N_5486,N_5264);
nor U6273 (N_6273,N_5159,N_5281);
and U6274 (N_6274,N_5139,N_4867);
nor U6275 (N_6275,N_5197,N_5325);
nor U6276 (N_6276,N_5147,N_5330);
xor U6277 (N_6277,N_5251,N_5582);
or U6278 (N_6278,N_5096,N_5532);
and U6279 (N_6279,N_5584,N_5502);
and U6280 (N_6280,N_5474,N_5544);
or U6281 (N_6281,N_4828,N_5083);
or U6282 (N_6282,N_4826,N_5495);
xor U6283 (N_6283,N_5017,N_4976);
xnor U6284 (N_6284,N_5370,N_5294);
nand U6285 (N_6285,N_5560,N_5440);
nand U6286 (N_6286,N_5107,N_5215);
xor U6287 (N_6287,N_5351,N_5280);
or U6288 (N_6288,N_5392,N_5485);
nor U6289 (N_6289,N_4955,N_5100);
nor U6290 (N_6290,N_5414,N_4948);
and U6291 (N_6291,N_5419,N_5074);
xor U6292 (N_6292,N_5405,N_5367);
xnor U6293 (N_6293,N_5457,N_5059);
or U6294 (N_6294,N_5337,N_5347);
and U6295 (N_6295,N_5508,N_5553);
and U6296 (N_6296,N_4956,N_4905);
or U6297 (N_6297,N_5262,N_5329);
or U6298 (N_6298,N_5383,N_4912);
and U6299 (N_6299,N_5378,N_4821);
nand U6300 (N_6300,N_5298,N_4816);
and U6301 (N_6301,N_5082,N_4865);
nor U6302 (N_6302,N_4902,N_5437);
or U6303 (N_6303,N_5468,N_5293);
xor U6304 (N_6304,N_5134,N_5127);
nor U6305 (N_6305,N_4885,N_5105);
nor U6306 (N_6306,N_5117,N_5314);
xnor U6307 (N_6307,N_5246,N_4854);
nand U6308 (N_6308,N_5072,N_5096);
xor U6309 (N_6309,N_5026,N_5216);
and U6310 (N_6310,N_5074,N_5131);
nand U6311 (N_6311,N_5305,N_5463);
xor U6312 (N_6312,N_5346,N_5591);
nor U6313 (N_6313,N_5117,N_5577);
and U6314 (N_6314,N_5302,N_4843);
nor U6315 (N_6315,N_5481,N_5058);
nand U6316 (N_6316,N_4889,N_4974);
nand U6317 (N_6317,N_4800,N_5053);
nor U6318 (N_6318,N_5247,N_5422);
or U6319 (N_6319,N_5450,N_5550);
and U6320 (N_6320,N_4850,N_4987);
nor U6321 (N_6321,N_5554,N_5401);
or U6322 (N_6322,N_5430,N_5065);
and U6323 (N_6323,N_5393,N_5426);
xnor U6324 (N_6324,N_5390,N_5092);
or U6325 (N_6325,N_5208,N_5550);
and U6326 (N_6326,N_4943,N_4945);
nor U6327 (N_6327,N_4853,N_5297);
or U6328 (N_6328,N_5593,N_5461);
and U6329 (N_6329,N_4906,N_5342);
or U6330 (N_6330,N_5507,N_4982);
nor U6331 (N_6331,N_5005,N_5116);
and U6332 (N_6332,N_5189,N_4821);
and U6333 (N_6333,N_5503,N_5003);
nor U6334 (N_6334,N_5478,N_4864);
xnor U6335 (N_6335,N_5066,N_5237);
and U6336 (N_6336,N_4976,N_5318);
and U6337 (N_6337,N_5258,N_4849);
nor U6338 (N_6338,N_5201,N_5329);
xor U6339 (N_6339,N_5127,N_5415);
and U6340 (N_6340,N_5386,N_5595);
and U6341 (N_6341,N_5575,N_4839);
xnor U6342 (N_6342,N_5506,N_4923);
and U6343 (N_6343,N_5030,N_5185);
and U6344 (N_6344,N_4927,N_5509);
nor U6345 (N_6345,N_5572,N_5010);
xnor U6346 (N_6346,N_5366,N_5533);
or U6347 (N_6347,N_4884,N_5288);
or U6348 (N_6348,N_5307,N_4803);
nand U6349 (N_6349,N_4918,N_5248);
or U6350 (N_6350,N_5046,N_4955);
and U6351 (N_6351,N_5114,N_5054);
and U6352 (N_6352,N_4960,N_5132);
or U6353 (N_6353,N_5323,N_5166);
nor U6354 (N_6354,N_5127,N_5135);
and U6355 (N_6355,N_5049,N_5156);
and U6356 (N_6356,N_4905,N_5225);
nand U6357 (N_6357,N_5197,N_5128);
or U6358 (N_6358,N_4893,N_5417);
and U6359 (N_6359,N_5094,N_5534);
and U6360 (N_6360,N_5073,N_4955);
xor U6361 (N_6361,N_5162,N_5036);
and U6362 (N_6362,N_5153,N_5375);
nand U6363 (N_6363,N_5367,N_5323);
or U6364 (N_6364,N_4800,N_5280);
nor U6365 (N_6365,N_5445,N_5422);
xnor U6366 (N_6366,N_5101,N_4924);
xnor U6367 (N_6367,N_4949,N_5144);
and U6368 (N_6368,N_5505,N_4958);
and U6369 (N_6369,N_4805,N_5352);
nand U6370 (N_6370,N_5059,N_5563);
or U6371 (N_6371,N_5243,N_4896);
nor U6372 (N_6372,N_5352,N_4892);
xor U6373 (N_6373,N_5183,N_5210);
or U6374 (N_6374,N_5523,N_5318);
and U6375 (N_6375,N_5362,N_5251);
and U6376 (N_6376,N_5051,N_5459);
nand U6377 (N_6377,N_5408,N_5002);
nand U6378 (N_6378,N_4804,N_5060);
xor U6379 (N_6379,N_5255,N_5597);
xnor U6380 (N_6380,N_5533,N_4973);
or U6381 (N_6381,N_5220,N_5450);
nand U6382 (N_6382,N_5325,N_4808);
nor U6383 (N_6383,N_5052,N_4819);
or U6384 (N_6384,N_5109,N_5003);
xor U6385 (N_6385,N_5580,N_4911);
xor U6386 (N_6386,N_5387,N_5373);
or U6387 (N_6387,N_5045,N_4807);
nand U6388 (N_6388,N_5412,N_5318);
nor U6389 (N_6389,N_5198,N_5594);
xor U6390 (N_6390,N_5319,N_4823);
nor U6391 (N_6391,N_5548,N_5521);
nor U6392 (N_6392,N_4977,N_4981);
nand U6393 (N_6393,N_5013,N_5523);
or U6394 (N_6394,N_5592,N_5065);
or U6395 (N_6395,N_5005,N_5100);
nand U6396 (N_6396,N_5595,N_4948);
xor U6397 (N_6397,N_5189,N_5373);
nor U6398 (N_6398,N_5523,N_4993);
and U6399 (N_6399,N_5550,N_5153);
nand U6400 (N_6400,N_6173,N_6337);
nand U6401 (N_6401,N_5713,N_6089);
or U6402 (N_6402,N_6288,N_5899);
xnor U6403 (N_6403,N_6348,N_5941);
nand U6404 (N_6404,N_5655,N_6042);
xnor U6405 (N_6405,N_6182,N_6266);
nand U6406 (N_6406,N_5919,N_5819);
nand U6407 (N_6407,N_6259,N_6188);
nand U6408 (N_6408,N_6244,N_6021);
or U6409 (N_6409,N_6119,N_6009);
nand U6410 (N_6410,N_5780,N_5690);
nand U6411 (N_6411,N_5891,N_5975);
and U6412 (N_6412,N_6026,N_5779);
and U6413 (N_6413,N_6085,N_6181);
nor U6414 (N_6414,N_6396,N_6335);
nor U6415 (N_6415,N_6378,N_6349);
nand U6416 (N_6416,N_5886,N_6150);
and U6417 (N_6417,N_6315,N_5726);
xor U6418 (N_6418,N_5757,N_6243);
and U6419 (N_6419,N_5695,N_6330);
and U6420 (N_6420,N_5679,N_5820);
nor U6421 (N_6421,N_5796,N_6199);
and U6422 (N_6422,N_6193,N_5752);
or U6423 (N_6423,N_6286,N_6164);
or U6424 (N_6424,N_5784,N_6290);
nand U6425 (N_6425,N_5644,N_5683);
xnor U6426 (N_6426,N_6324,N_5746);
and U6427 (N_6427,N_5646,N_5730);
and U6428 (N_6428,N_5716,N_6232);
or U6429 (N_6429,N_6251,N_6344);
and U6430 (N_6430,N_6018,N_5635);
or U6431 (N_6431,N_5952,N_6139);
nand U6432 (N_6432,N_5856,N_6358);
and U6433 (N_6433,N_5883,N_5900);
and U6434 (N_6434,N_6005,N_5632);
xor U6435 (N_6435,N_5824,N_5788);
and U6436 (N_6436,N_6273,N_6377);
xor U6437 (N_6437,N_5927,N_5618);
xor U6438 (N_6438,N_6045,N_5848);
nand U6439 (N_6439,N_6316,N_5648);
and U6440 (N_6440,N_5966,N_5855);
and U6441 (N_6441,N_6012,N_6227);
and U6442 (N_6442,N_6058,N_5860);
or U6443 (N_6443,N_6000,N_5974);
or U6444 (N_6444,N_5770,N_6262);
nor U6445 (N_6445,N_5893,N_5715);
or U6446 (N_6446,N_5773,N_6351);
xor U6447 (N_6447,N_5877,N_6299);
xnor U6448 (N_6448,N_5607,N_5669);
or U6449 (N_6449,N_6131,N_5653);
xnor U6450 (N_6450,N_5994,N_6271);
or U6451 (N_6451,N_6168,N_5834);
xnor U6452 (N_6452,N_5745,N_5892);
or U6453 (N_6453,N_6109,N_5708);
or U6454 (N_6454,N_6054,N_6385);
and U6455 (N_6455,N_5762,N_5987);
and U6456 (N_6456,N_6350,N_6307);
and U6457 (N_6457,N_5818,N_5611);
nor U6458 (N_6458,N_5782,N_5787);
nand U6459 (N_6459,N_6121,N_5768);
or U6460 (N_6460,N_6136,N_5793);
xnor U6461 (N_6461,N_6379,N_5969);
xor U6462 (N_6462,N_6187,N_5928);
or U6463 (N_6463,N_6105,N_6143);
and U6464 (N_6464,N_6254,N_5685);
nor U6465 (N_6465,N_5874,N_5907);
nand U6466 (N_6466,N_6333,N_5677);
or U6467 (N_6467,N_5970,N_5605);
nor U6468 (N_6468,N_6013,N_6095);
xnor U6469 (N_6469,N_5875,N_5718);
and U6470 (N_6470,N_5687,N_6353);
or U6471 (N_6471,N_6008,N_5761);
nor U6472 (N_6472,N_5852,N_6142);
or U6473 (N_6473,N_5961,N_5917);
or U6474 (N_6474,N_5795,N_5766);
xor U6475 (N_6475,N_5932,N_5783);
xnor U6476 (N_6476,N_5758,N_5665);
nor U6477 (N_6477,N_5697,N_5674);
nor U6478 (N_6478,N_5634,N_5826);
and U6479 (N_6479,N_6137,N_5957);
and U6480 (N_6480,N_6276,N_6183);
nor U6481 (N_6481,N_6148,N_5986);
xor U6482 (N_6482,N_6154,N_5876);
nand U6483 (N_6483,N_6050,N_5809);
nor U6484 (N_6484,N_6103,N_6261);
and U6485 (N_6485,N_6197,N_5837);
and U6486 (N_6486,N_5955,N_5923);
xor U6487 (N_6487,N_5672,N_6192);
nor U6488 (N_6488,N_5616,N_6064);
xor U6489 (N_6489,N_6284,N_6293);
xor U6490 (N_6490,N_5640,N_5921);
xnor U6491 (N_6491,N_6091,N_5624);
xor U6492 (N_6492,N_5650,N_6102);
nor U6493 (N_6493,N_5951,N_5976);
or U6494 (N_6494,N_5915,N_6117);
or U6495 (N_6495,N_5850,N_6175);
nor U6496 (N_6496,N_5642,N_6057);
xor U6497 (N_6497,N_6036,N_5682);
or U6498 (N_6498,N_5910,N_6308);
nand U6499 (N_6499,N_5636,N_5673);
or U6500 (N_6500,N_5841,N_5866);
or U6501 (N_6501,N_5844,N_5980);
and U6502 (N_6502,N_6310,N_5728);
or U6503 (N_6503,N_5924,N_5991);
and U6504 (N_6504,N_5637,N_5777);
xor U6505 (N_6505,N_5967,N_6205);
xor U6506 (N_6506,N_5948,N_5939);
xnor U6507 (N_6507,N_5663,N_6368);
or U6508 (N_6508,N_6072,N_6287);
and U6509 (N_6509,N_6106,N_6252);
and U6510 (N_6510,N_6237,N_5739);
and U6511 (N_6511,N_6198,N_5950);
nor U6512 (N_6512,N_6208,N_5680);
xor U6513 (N_6513,N_5714,N_6135);
or U6514 (N_6514,N_6234,N_6086);
xnor U6515 (N_6515,N_6108,N_6221);
xor U6516 (N_6516,N_6365,N_6046);
and U6517 (N_6517,N_5664,N_5827);
nor U6518 (N_6518,N_6043,N_6247);
nor U6519 (N_6519,N_5754,N_5702);
xnor U6520 (N_6520,N_6170,N_6074);
and U6521 (N_6521,N_6246,N_6025);
nor U6522 (N_6522,N_6149,N_5743);
nor U6523 (N_6523,N_5906,N_6063);
and U6524 (N_6524,N_5811,N_5843);
nand U6525 (N_6525,N_6264,N_5721);
or U6526 (N_6526,N_5944,N_6144);
nand U6527 (N_6527,N_5705,N_6165);
nand U6528 (N_6528,N_5785,N_5678);
xnor U6529 (N_6529,N_6029,N_6278);
or U6530 (N_6530,N_5704,N_6028);
and U6531 (N_6531,N_6129,N_6283);
or U6532 (N_6532,N_6245,N_5775);
nand U6533 (N_6533,N_6049,N_6156);
and U6534 (N_6534,N_5861,N_6190);
nand U6535 (N_6535,N_5606,N_6145);
or U6536 (N_6536,N_5904,N_5814);
nor U6537 (N_6537,N_6120,N_6210);
xnor U6538 (N_6538,N_5964,N_6125);
nand U6539 (N_6539,N_6006,N_6393);
or U6540 (N_6540,N_6040,N_5959);
or U6541 (N_6541,N_5920,N_6322);
xnor U6542 (N_6542,N_5865,N_5608);
and U6543 (N_6543,N_6023,N_5619);
nand U6544 (N_6544,N_6179,N_6048);
xnor U6545 (N_6545,N_6285,N_5813);
and U6546 (N_6546,N_5997,N_6381);
nor U6547 (N_6547,N_6127,N_5999);
and U6548 (N_6548,N_5688,N_6067);
or U6549 (N_6549,N_5645,N_6389);
xor U6550 (N_6550,N_6313,N_6253);
nor U6551 (N_6551,N_6163,N_5882);
and U6552 (N_6552,N_5706,N_5949);
xor U6553 (N_6553,N_6073,N_6217);
nand U6554 (N_6554,N_6203,N_5838);
nor U6555 (N_6555,N_5890,N_5701);
nand U6556 (N_6556,N_5894,N_6314);
nor U6557 (N_6557,N_5696,N_5651);
and U6558 (N_6558,N_6060,N_5734);
or U6559 (N_6559,N_5990,N_5840);
nand U6560 (N_6560,N_6394,N_5615);
and U6561 (N_6561,N_6134,N_6001);
nor U6562 (N_6562,N_6367,N_5984);
xnor U6563 (N_6563,N_5765,N_5625);
or U6564 (N_6564,N_5749,N_5903);
nor U6565 (N_6565,N_5601,N_6263);
and U6566 (N_6566,N_5965,N_5914);
nand U6567 (N_6567,N_6122,N_6141);
nand U6568 (N_6568,N_5981,N_6357);
or U6569 (N_6569,N_5712,N_6255);
and U6570 (N_6570,N_5929,N_6189);
nor U6571 (N_6571,N_5934,N_6031);
nand U6572 (N_6572,N_6390,N_6305);
xor U6573 (N_6573,N_6032,N_5628);
nand U6574 (N_6574,N_5772,N_5871);
nand U6575 (N_6575,N_5895,N_5845);
or U6576 (N_6576,N_6354,N_5764);
or U6577 (N_6577,N_6382,N_5698);
nand U6578 (N_6578,N_6114,N_5759);
and U6579 (N_6579,N_5786,N_5709);
or U6580 (N_6580,N_6319,N_6019);
nand U6581 (N_6581,N_5804,N_5660);
nand U6582 (N_6582,N_6265,N_6070);
and U6583 (N_6583,N_6004,N_6162);
or U6584 (N_6584,N_5731,N_6138);
xor U6585 (N_6585,N_5985,N_6184);
or U6586 (N_6586,N_5700,N_6177);
xnor U6587 (N_6587,N_6159,N_6155);
nand U6588 (N_6588,N_5971,N_6303);
nand U6589 (N_6589,N_5854,N_5609);
nor U6590 (N_6590,N_5610,N_5922);
nor U6591 (N_6591,N_5960,N_6200);
nor U6592 (N_6592,N_6080,N_5807);
nand U6593 (N_6593,N_6325,N_5954);
nand U6594 (N_6594,N_5707,N_5753);
or U6595 (N_6595,N_5799,N_6171);
and U6596 (N_6596,N_6140,N_5719);
xnor U6597 (N_6597,N_6016,N_6123);
and U6598 (N_6598,N_6037,N_5756);
or U6599 (N_6599,N_6110,N_5869);
or U6600 (N_6600,N_5661,N_6115);
or U6601 (N_6601,N_6185,N_5626);
or U6602 (N_6602,N_5670,N_6280);
xor U6603 (N_6603,N_5815,N_6399);
and U6604 (N_6604,N_5620,N_5736);
and U6605 (N_6605,N_6239,N_6279);
or U6606 (N_6606,N_6130,N_6268);
nor U6607 (N_6607,N_6090,N_5600);
or U6608 (N_6608,N_5668,N_6225);
xnor U6609 (N_6609,N_5729,N_5681);
nand U6610 (N_6610,N_5846,N_5689);
and U6611 (N_6611,N_5872,N_6274);
xor U6612 (N_6612,N_6218,N_6151);
or U6613 (N_6613,N_6124,N_6281);
xor U6614 (N_6614,N_5885,N_6010);
and U6615 (N_6615,N_6157,N_5781);
nand U6616 (N_6616,N_5889,N_5778);
xnor U6617 (N_6617,N_6034,N_5662);
nor U6618 (N_6618,N_5797,N_6346);
or U6619 (N_6619,N_5717,N_6223);
or U6620 (N_6620,N_5847,N_5992);
nand U6621 (N_6621,N_5973,N_5613);
nand U6622 (N_6622,N_6291,N_6269);
xnor U6623 (N_6623,N_5751,N_5833);
nand U6624 (N_6624,N_5776,N_6206);
nand U6625 (N_6625,N_6180,N_6334);
xnor U6626 (N_6626,N_5732,N_5901);
and U6627 (N_6627,N_6309,N_6235);
nor U6628 (N_6628,N_6161,N_6242);
and U6629 (N_6629,N_5849,N_5755);
xor U6630 (N_6630,N_5935,N_5888);
or U6631 (N_6631,N_6300,N_5909);
nor U6632 (N_6632,N_6250,N_6212);
and U6633 (N_6633,N_6317,N_6336);
xor U6634 (N_6634,N_5733,N_6374);
nand U6635 (N_6635,N_5667,N_5978);
nor U6636 (N_6636,N_6107,N_5870);
xor U6637 (N_6637,N_5958,N_6258);
xor U6638 (N_6638,N_6201,N_6318);
nand U6639 (N_6639,N_6065,N_6014);
nor U6640 (N_6640,N_5943,N_5604);
or U6641 (N_6641,N_6147,N_5617);
xor U6642 (N_6642,N_5771,N_6345);
or U6643 (N_6643,N_6191,N_6097);
and U6644 (N_6644,N_6167,N_6002);
nand U6645 (N_6645,N_6295,N_6071);
xnor U6646 (N_6646,N_6079,N_5864);
xor U6647 (N_6647,N_5684,N_5897);
nor U6648 (N_6648,N_5735,N_5828);
and U6649 (N_6649,N_6272,N_6297);
or U6650 (N_6650,N_6301,N_5808);
or U6651 (N_6651,N_6364,N_6209);
xnor U6652 (N_6652,N_5614,N_6372);
nand U6653 (N_6653,N_6388,N_6196);
nor U6654 (N_6654,N_6062,N_6395);
and U6655 (N_6655,N_5930,N_6338);
or U6656 (N_6656,N_5794,N_6224);
and U6657 (N_6657,N_6370,N_5887);
nor U6658 (N_6658,N_6238,N_6275);
nand U6659 (N_6659,N_5858,N_6215);
nor U6660 (N_6660,N_6320,N_5913);
and U6661 (N_6661,N_5654,N_6128);
nor U6662 (N_6662,N_5962,N_6146);
and U6663 (N_6663,N_6326,N_6094);
nor U6664 (N_6664,N_6195,N_6373);
and U6665 (N_6665,N_5630,N_5938);
and U6666 (N_6666,N_5982,N_5633);
and U6667 (N_6667,N_6022,N_5806);
xnor U6668 (N_6668,N_6220,N_5691);
xnor U6669 (N_6669,N_5659,N_6039);
and U6670 (N_6670,N_5803,N_6306);
xor U6671 (N_6671,N_6007,N_6024);
and U6672 (N_6672,N_5925,N_6298);
nor U6673 (N_6673,N_5989,N_5623);
nand U6674 (N_6674,N_5658,N_6116);
or U6675 (N_6675,N_6363,N_5801);
or U6676 (N_6676,N_5983,N_6292);
nand U6677 (N_6677,N_5767,N_6248);
nor U6678 (N_6678,N_5693,N_6213);
or U6679 (N_6679,N_5737,N_6100);
or U6680 (N_6680,N_5742,N_6166);
and U6681 (N_6681,N_5612,N_6133);
xnor U6682 (N_6682,N_6321,N_5789);
nor U6683 (N_6683,N_6059,N_6053);
and U6684 (N_6684,N_5652,N_5744);
or U6685 (N_6685,N_5649,N_5656);
nand U6686 (N_6686,N_6088,N_5802);
nor U6687 (N_6687,N_5926,N_5643);
xnor U6688 (N_6688,N_6256,N_6329);
nand U6689 (N_6689,N_6371,N_6211);
nand U6690 (N_6690,N_5908,N_6098);
xor U6691 (N_6691,N_6312,N_6076);
xor U6692 (N_6692,N_5988,N_5947);
or U6693 (N_6693,N_5879,N_6087);
nand U6694 (N_6694,N_5829,N_6236);
xor U6695 (N_6695,N_6101,N_5798);
nand U6696 (N_6696,N_5671,N_6392);
nand U6697 (N_6697,N_6081,N_5998);
nor U6698 (N_6698,N_6084,N_6304);
and U6699 (N_6699,N_5812,N_6347);
and U6700 (N_6700,N_5816,N_5720);
nor U6701 (N_6701,N_6003,N_5851);
and U6702 (N_6702,N_6038,N_5996);
nand U6703 (N_6703,N_6342,N_5995);
xnor U6704 (N_6704,N_6066,N_6230);
nor U6705 (N_6705,N_5747,N_6343);
xnor U6706 (N_6706,N_5694,N_6207);
nand U6707 (N_6707,N_5863,N_6380);
xnor U6708 (N_6708,N_5703,N_5911);
and U6709 (N_6709,N_6033,N_6068);
or U6710 (N_6710,N_5769,N_6331);
xor U6711 (N_6711,N_6112,N_6035);
and U6712 (N_6712,N_5627,N_6222);
xor U6713 (N_6713,N_5741,N_6075);
xor U6714 (N_6714,N_5622,N_5791);
or U6715 (N_6715,N_6041,N_5993);
nor U6716 (N_6716,N_5868,N_5725);
nand U6717 (N_6717,N_6356,N_5936);
and U6718 (N_6718,N_6214,N_5880);
nand U6719 (N_6719,N_6289,N_5898);
xor U6720 (N_6720,N_6077,N_5675);
nand U6721 (N_6721,N_6257,N_5835);
xnor U6722 (N_6722,N_6327,N_6152);
xnor U6723 (N_6723,N_5629,N_6339);
or U6724 (N_6724,N_5956,N_5738);
nand U6725 (N_6725,N_6233,N_5676);
and U6726 (N_6726,N_5657,N_6267);
nand U6727 (N_6727,N_5896,N_6277);
xnor U6728 (N_6728,N_6176,N_5937);
nand U6729 (N_6729,N_6132,N_5699);
and U6730 (N_6730,N_6093,N_6369);
or U6731 (N_6731,N_5884,N_5942);
or U6732 (N_6732,N_6056,N_6229);
and U6733 (N_6733,N_6294,N_6174);
xnor U6734 (N_6734,N_6359,N_6323);
nor U6735 (N_6735,N_6332,N_5853);
xor U6736 (N_6736,N_6386,N_6204);
or U6737 (N_6737,N_5881,N_5724);
nand U6738 (N_6738,N_6397,N_5748);
nand U6739 (N_6739,N_5867,N_5723);
xnor U6740 (N_6740,N_6160,N_5666);
nand U6741 (N_6741,N_5692,N_6219);
or U6742 (N_6742,N_6027,N_5822);
nor U6743 (N_6743,N_6083,N_5763);
and U6744 (N_6744,N_6118,N_6194);
and U6745 (N_6745,N_6328,N_5602);
or U6746 (N_6746,N_6202,N_6011);
xor U6747 (N_6747,N_6398,N_6375);
or U6748 (N_6748,N_5831,N_6111);
xor U6749 (N_6749,N_5905,N_5750);
xnor U6750 (N_6750,N_5790,N_5727);
nor U6751 (N_6751,N_6340,N_6241);
nand U6752 (N_6752,N_6030,N_5603);
and U6753 (N_6753,N_5710,N_5711);
nor U6754 (N_6754,N_6153,N_5639);
nand U6755 (N_6755,N_5878,N_6052);
nand U6756 (N_6756,N_5918,N_5902);
xnor U6757 (N_6757,N_5953,N_5912);
nor U6758 (N_6758,N_5830,N_5821);
nand U6759 (N_6759,N_5931,N_6282);
or U6760 (N_6760,N_6366,N_6384);
and U6761 (N_6761,N_6260,N_6044);
xnor U6762 (N_6762,N_5825,N_6360);
or U6763 (N_6763,N_6158,N_5800);
xor U6764 (N_6764,N_6078,N_6352);
nor U6765 (N_6765,N_5641,N_6020);
nor U6766 (N_6766,N_5979,N_5946);
nand U6767 (N_6767,N_5638,N_6082);
and U6768 (N_6768,N_5977,N_5722);
nor U6769 (N_6769,N_5740,N_6126);
nor U6770 (N_6770,N_6015,N_5857);
nor U6771 (N_6771,N_5933,N_6047);
nand U6772 (N_6772,N_5972,N_5963);
or U6773 (N_6773,N_5842,N_6361);
xor U6774 (N_6774,N_5859,N_5836);
xor U6775 (N_6775,N_6231,N_6240);
xor U6776 (N_6776,N_5968,N_6362);
nand U6777 (N_6777,N_5940,N_5823);
xor U6778 (N_6778,N_5817,N_6376);
nor U6779 (N_6779,N_6169,N_5862);
nand U6780 (N_6780,N_6186,N_5873);
and U6781 (N_6781,N_5621,N_6017);
nand U6782 (N_6782,N_6216,N_6104);
or U6783 (N_6783,N_5810,N_5647);
nand U6784 (N_6784,N_6061,N_6383);
and U6785 (N_6785,N_6341,N_6226);
nand U6786 (N_6786,N_5686,N_6228);
nand U6787 (N_6787,N_6296,N_6387);
or U6788 (N_6788,N_5916,N_6051);
or U6789 (N_6789,N_6270,N_6172);
xor U6790 (N_6790,N_5774,N_6096);
or U6791 (N_6791,N_6055,N_5839);
xnor U6792 (N_6792,N_5805,N_5760);
and U6793 (N_6793,N_6069,N_5945);
nand U6794 (N_6794,N_6113,N_6311);
and U6795 (N_6795,N_6302,N_6391);
xor U6796 (N_6796,N_6249,N_5792);
nor U6797 (N_6797,N_6178,N_6092);
nand U6798 (N_6798,N_5832,N_6355);
and U6799 (N_6799,N_6099,N_5631);
nand U6800 (N_6800,N_6344,N_5867);
xnor U6801 (N_6801,N_6155,N_5847);
nand U6802 (N_6802,N_6079,N_6317);
and U6803 (N_6803,N_5820,N_6029);
nand U6804 (N_6804,N_6264,N_5833);
and U6805 (N_6805,N_5894,N_5665);
or U6806 (N_6806,N_6345,N_5966);
nor U6807 (N_6807,N_6161,N_6024);
nor U6808 (N_6808,N_6319,N_6040);
xnor U6809 (N_6809,N_5806,N_6175);
nand U6810 (N_6810,N_5611,N_6273);
nand U6811 (N_6811,N_5641,N_5893);
or U6812 (N_6812,N_6277,N_5743);
xor U6813 (N_6813,N_5974,N_6202);
nand U6814 (N_6814,N_6270,N_6352);
or U6815 (N_6815,N_6351,N_5856);
xor U6816 (N_6816,N_5837,N_5877);
and U6817 (N_6817,N_5861,N_6066);
nand U6818 (N_6818,N_5686,N_6265);
xor U6819 (N_6819,N_5641,N_5706);
xnor U6820 (N_6820,N_5603,N_6145);
xor U6821 (N_6821,N_5990,N_5904);
nand U6822 (N_6822,N_5964,N_5989);
and U6823 (N_6823,N_5854,N_5728);
nand U6824 (N_6824,N_6107,N_5754);
and U6825 (N_6825,N_6333,N_5694);
nand U6826 (N_6826,N_6263,N_5747);
xnor U6827 (N_6827,N_6258,N_6114);
xnor U6828 (N_6828,N_6215,N_6384);
nor U6829 (N_6829,N_6005,N_6383);
nand U6830 (N_6830,N_6026,N_6293);
nand U6831 (N_6831,N_6296,N_5805);
nor U6832 (N_6832,N_6098,N_6157);
nor U6833 (N_6833,N_6201,N_6111);
xor U6834 (N_6834,N_6350,N_5821);
nand U6835 (N_6835,N_6000,N_6138);
and U6836 (N_6836,N_5769,N_5990);
xnor U6837 (N_6837,N_5931,N_5666);
or U6838 (N_6838,N_6276,N_5827);
nor U6839 (N_6839,N_5717,N_5994);
nor U6840 (N_6840,N_6260,N_6034);
nand U6841 (N_6841,N_5790,N_6340);
xor U6842 (N_6842,N_5758,N_5934);
or U6843 (N_6843,N_5728,N_6325);
or U6844 (N_6844,N_6255,N_5655);
and U6845 (N_6845,N_6327,N_5984);
or U6846 (N_6846,N_5736,N_5996);
nor U6847 (N_6847,N_5792,N_6029);
xor U6848 (N_6848,N_5711,N_6312);
or U6849 (N_6849,N_6239,N_5914);
and U6850 (N_6850,N_6180,N_6194);
xor U6851 (N_6851,N_5935,N_5916);
nand U6852 (N_6852,N_5978,N_5611);
nor U6853 (N_6853,N_5835,N_5666);
nand U6854 (N_6854,N_5711,N_5652);
nand U6855 (N_6855,N_5986,N_6110);
nand U6856 (N_6856,N_6396,N_6138);
nand U6857 (N_6857,N_6142,N_6064);
nand U6858 (N_6858,N_6191,N_5856);
nand U6859 (N_6859,N_5624,N_6270);
xnor U6860 (N_6860,N_6120,N_5879);
xor U6861 (N_6861,N_5886,N_6204);
xor U6862 (N_6862,N_5760,N_5823);
nor U6863 (N_6863,N_5875,N_5939);
or U6864 (N_6864,N_5912,N_6017);
or U6865 (N_6865,N_5656,N_5945);
xnor U6866 (N_6866,N_6375,N_5743);
xnor U6867 (N_6867,N_6258,N_6245);
nand U6868 (N_6868,N_6169,N_5662);
xnor U6869 (N_6869,N_6090,N_5978);
nand U6870 (N_6870,N_6080,N_5713);
and U6871 (N_6871,N_5610,N_5908);
nand U6872 (N_6872,N_5760,N_5900);
xnor U6873 (N_6873,N_6385,N_6338);
or U6874 (N_6874,N_5613,N_5952);
nand U6875 (N_6875,N_6191,N_6287);
nor U6876 (N_6876,N_5904,N_5879);
xnor U6877 (N_6877,N_6339,N_5740);
and U6878 (N_6878,N_5948,N_5912);
xor U6879 (N_6879,N_5974,N_6112);
nand U6880 (N_6880,N_5925,N_6172);
xor U6881 (N_6881,N_5874,N_5900);
nor U6882 (N_6882,N_5830,N_5709);
xnor U6883 (N_6883,N_6268,N_6330);
xnor U6884 (N_6884,N_6024,N_6336);
nand U6885 (N_6885,N_5999,N_6317);
xnor U6886 (N_6886,N_6055,N_5670);
nor U6887 (N_6887,N_6043,N_5601);
nor U6888 (N_6888,N_6142,N_5642);
and U6889 (N_6889,N_5990,N_6071);
and U6890 (N_6890,N_5884,N_6201);
nand U6891 (N_6891,N_6256,N_6354);
nand U6892 (N_6892,N_5784,N_6230);
nand U6893 (N_6893,N_5813,N_6104);
and U6894 (N_6894,N_6285,N_6043);
nor U6895 (N_6895,N_5841,N_5621);
nor U6896 (N_6896,N_6398,N_6083);
nand U6897 (N_6897,N_6171,N_6182);
xnor U6898 (N_6898,N_5610,N_6034);
or U6899 (N_6899,N_6389,N_5857);
nor U6900 (N_6900,N_6184,N_6299);
nor U6901 (N_6901,N_6129,N_5886);
xor U6902 (N_6902,N_5989,N_5700);
nor U6903 (N_6903,N_6305,N_5679);
and U6904 (N_6904,N_6024,N_5669);
and U6905 (N_6905,N_6146,N_5783);
or U6906 (N_6906,N_6321,N_6358);
nor U6907 (N_6907,N_6238,N_5787);
nor U6908 (N_6908,N_6367,N_5780);
and U6909 (N_6909,N_5735,N_5708);
xor U6910 (N_6910,N_5832,N_6143);
nand U6911 (N_6911,N_6281,N_5772);
and U6912 (N_6912,N_5896,N_6216);
and U6913 (N_6913,N_6115,N_5905);
or U6914 (N_6914,N_5663,N_5990);
nand U6915 (N_6915,N_5883,N_5824);
nor U6916 (N_6916,N_5747,N_5869);
nand U6917 (N_6917,N_6039,N_5759);
nor U6918 (N_6918,N_6231,N_5746);
nand U6919 (N_6919,N_5603,N_6074);
nor U6920 (N_6920,N_6384,N_6370);
xor U6921 (N_6921,N_5713,N_5923);
and U6922 (N_6922,N_5904,N_5874);
nor U6923 (N_6923,N_6104,N_5647);
nand U6924 (N_6924,N_5762,N_6328);
or U6925 (N_6925,N_5991,N_6122);
nand U6926 (N_6926,N_6039,N_5999);
xnor U6927 (N_6927,N_6046,N_5688);
xnor U6928 (N_6928,N_6174,N_6396);
xnor U6929 (N_6929,N_5810,N_5970);
or U6930 (N_6930,N_5676,N_6399);
or U6931 (N_6931,N_6382,N_6343);
nor U6932 (N_6932,N_6284,N_5748);
xor U6933 (N_6933,N_6260,N_6011);
nor U6934 (N_6934,N_5864,N_5619);
xor U6935 (N_6935,N_5887,N_6261);
or U6936 (N_6936,N_6141,N_6134);
xor U6937 (N_6937,N_6319,N_6007);
or U6938 (N_6938,N_5870,N_5998);
xnor U6939 (N_6939,N_6002,N_5656);
or U6940 (N_6940,N_6055,N_5929);
xor U6941 (N_6941,N_5864,N_6146);
or U6942 (N_6942,N_5982,N_5946);
and U6943 (N_6943,N_5769,N_6260);
and U6944 (N_6944,N_6167,N_6275);
xnor U6945 (N_6945,N_5791,N_6240);
and U6946 (N_6946,N_5990,N_5739);
and U6947 (N_6947,N_5745,N_5806);
nand U6948 (N_6948,N_6355,N_5873);
or U6949 (N_6949,N_6208,N_5916);
xnor U6950 (N_6950,N_6119,N_6231);
nand U6951 (N_6951,N_5734,N_6389);
or U6952 (N_6952,N_6280,N_5627);
nor U6953 (N_6953,N_6273,N_6168);
nor U6954 (N_6954,N_6101,N_5767);
or U6955 (N_6955,N_6163,N_6185);
or U6956 (N_6956,N_6301,N_6267);
xor U6957 (N_6957,N_5608,N_5834);
xnor U6958 (N_6958,N_6361,N_6390);
and U6959 (N_6959,N_5828,N_6186);
nor U6960 (N_6960,N_5618,N_5952);
nor U6961 (N_6961,N_5709,N_6197);
and U6962 (N_6962,N_6266,N_6169);
xnor U6963 (N_6963,N_5826,N_5671);
and U6964 (N_6964,N_6373,N_5607);
nor U6965 (N_6965,N_6367,N_5888);
nand U6966 (N_6966,N_5883,N_6217);
nor U6967 (N_6967,N_6101,N_6379);
nor U6968 (N_6968,N_6060,N_5830);
xnor U6969 (N_6969,N_5759,N_5648);
nor U6970 (N_6970,N_5602,N_5911);
nand U6971 (N_6971,N_6386,N_5962);
xor U6972 (N_6972,N_5852,N_5665);
nand U6973 (N_6973,N_5754,N_6393);
xnor U6974 (N_6974,N_6136,N_5706);
or U6975 (N_6975,N_6201,N_5900);
nand U6976 (N_6976,N_6300,N_5888);
nor U6977 (N_6977,N_5830,N_6263);
or U6978 (N_6978,N_6209,N_6272);
and U6979 (N_6979,N_6127,N_6304);
or U6980 (N_6980,N_6395,N_5925);
xnor U6981 (N_6981,N_6349,N_5863);
and U6982 (N_6982,N_5718,N_5758);
nor U6983 (N_6983,N_5801,N_6115);
nor U6984 (N_6984,N_6160,N_6037);
or U6985 (N_6985,N_6218,N_5941);
nor U6986 (N_6986,N_5678,N_5985);
xor U6987 (N_6987,N_5769,N_5644);
and U6988 (N_6988,N_6337,N_5796);
nand U6989 (N_6989,N_6255,N_6133);
nor U6990 (N_6990,N_6344,N_5796);
and U6991 (N_6991,N_6397,N_5951);
nor U6992 (N_6992,N_6356,N_5809);
xnor U6993 (N_6993,N_6141,N_5859);
xnor U6994 (N_6994,N_6088,N_6164);
nand U6995 (N_6995,N_5865,N_5774);
xnor U6996 (N_6996,N_6135,N_5858);
or U6997 (N_6997,N_5829,N_6362);
xnor U6998 (N_6998,N_6207,N_5651);
and U6999 (N_6999,N_6144,N_5624);
and U7000 (N_7000,N_6162,N_5963);
nor U7001 (N_7001,N_6085,N_5837);
nor U7002 (N_7002,N_5925,N_5956);
nand U7003 (N_7003,N_5770,N_6004);
nor U7004 (N_7004,N_5987,N_5723);
nand U7005 (N_7005,N_6133,N_6355);
nor U7006 (N_7006,N_5775,N_5718);
nand U7007 (N_7007,N_6290,N_6108);
nor U7008 (N_7008,N_6030,N_5694);
nand U7009 (N_7009,N_5888,N_5924);
or U7010 (N_7010,N_6376,N_6360);
xor U7011 (N_7011,N_6333,N_6259);
or U7012 (N_7012,N_6397,N_5787);
and U7013 (N_7013,N_6311,N_6397);
and U7014 (N_7014,N_5697,N_6161);
nor U7015 (N_7015,N_6312,N_6096);
and U7016 (N_7016,N_6082,N_6291);
xor U7017 (N_7017,N_6356,N_5808);
or U7018 (N_7018,N_6103,N_6147);
or U7019 (N_7019,N_5644,N_5703);
nor U7020 (N_7020,N_6216,N_6280);
nand U7021 (N_7021,N_6237,N_5865);
or U7022 (N_7022,N_5990,N_6140);
and U7023 (N_7023,N_5932,N_5717);
or U7024 (N_7024,N_5847,N_5731);
and U7025 (N_7025,N_6324,N_6053);
nand U7026 (N_7026,N_6295,N_6001);
and U7027 (N_7027,N_5712,N_5955);
or U7028 (N_7028,N_5677,N_6086);
nor U7029 (N_7029,N_5735,N_6268);
and U7030 (N_7030,N_6307,N_5780);
or U7031 (N_7031,N_5956,N_6031);
xor U7032 (N_7032,N_5994,N_5934);
and U7033 (N_7033,N_6076,N_6092);
xor U7034 (N_7034,N_6006,N_5711);
xor U7035 (N_7035,N_5859,N_5644);
and U7036 (N_7036,N_6272,N_5750);
xnor U7037 (N_7037,N_6287,N_5919);
nand U7038 (N_7038,N_5730,N_5983);
nor U7039 (N_7039,N_6185,N_6096);
or U7040 (N_7040,N_6294,N_5863);
nor U7041 (N_7041,N_5835,N_6097);
or U7042 (N_7042,N_5754,N_5986);
nand U7043 (N_7043,N_6070,N_6075);
nor U7044 (N_7044,N_5775,N_6276);
or U7045 (N_7045,N_5718,N_6083);
nor U7046 (N_7046,N_6185,N_6385);
nor U7047 (N_7047,N_6062,N_6266);
xnor U7048 (N_7048,N_6138,N_5884);
and U7049 (N_7049,N_6369,N_6169);
and U7050 (N_7050,N_5916,N_6156);
or U7051 (N_7051,N_5793,N_6147);
nor U7052 (N_7052,N_6336,N_6331);
nand U7053 (N_7053,N_5830,N_6038);
nor U7054 (N_7054,N_5675,N_5890);
xnor U7055 (N_7055,N_5603,N_5657);
xor U7056 (N_7056,N_5631,N_6073);
and U7057 (N_7057,N_6032,N_5722);
and U7058 (N_7058,N_5968,N_6385);
nand U7059 (N_7059,N_5910,N_6105);
nor U7060 (N_7060,N_6265,N_6057);
nand U7061 (N_7061,N_6289,N_5921);
and U7062 (N_7062,N_5696,N_6310);
or U7063 (N_7063,N_5716,N_5795);
or U7064 (N_7064,N_5794,N_5786);
or U7065 (N_7065,N_5867,N_6104);
nor U7066 (N_7066,N_6135,N_5926);
nand U7067 (N_7067,N_6156,N_5621);
xnor U7068 (N_7068,N_6251,N_6092);
nand U7069 (N_7069,N_6145,N_6108);
nand U7070 (N_7070,N_5819,N_6270);
nor U7071 (N_7071,N_5689,N_5921);
nand U7072 (N_7072,N_6365,N_6384);
and U7073 (N_7073,N_5825,N_5743);
and U7074 (N_7074,N_5753,N_6381);
nor U7075 (N_7075,N_6309,N_6008);
nor U7076 (N_7076,N_6179,N_6393);
xor U7077 (N_7077,N_5675,N_5601);
xnor U7078 (N_7078,N_6321,N_6143);
nand U7079 (N_7079,N_6321,N_6141);
xnor U7080 (N_7080,N_5811,N_5638);
or U7081 (N_7081,N_6015,N_5999);
nand U7082 (N_7082,N_6015,N_6299);
and U7083 (N_7083,N_5900,N_5726);
or U7084 (N_7084,N_5853,N_6341);
xnor U7085 (N_7085,N_6132,N_5841);
and U7086 (N_7086,N_6244,N_6363);
or U7087 (N_7087,N_5703,N_6237);
nor U7088 (N_7088,N_5726,N_5613);
or U7089 (N_7089,N_5793,N_6393);
or U7090 (N_7090,N_6302,N_6062);
and U7091 (N_7091,N_6325,N_6215);
nor U7092 (N_7092,N_6352,N_5647);
or U7093 (N_7093,N_5922,N_6134);
nor U7094 (N_7094,N_5775,N_6164);
nor U7095 (N_7095,N_5813,N_6150);
xnor U7096 (N_7096,N_5991,N_6192);
xor U7097 (N_7097,N_5682,N_6025);
or U7098 (N_7098,N_6159,N_6309);
and U7099 (N_7099,N_5662,N_6204);
nor U7100 (N_7100,N_6080,N_5738);
nor U7101 (N_7101,N_5731,N_5873);
or U7102 (N_7102,N_5662,N_6207);
xnor U7103 (N_7103,N_5629,N_6275);
nor U7104 (N_7104,N_6264,N_6020);
nor U7105 (N_7105,N_5718,N_5692);
nor U7106 (N_7106,N_6190,N_6010);
nor U7107 (N_7107,N_5708,N_5654);
nor U7108 (N_7108,N_5775,N_6198);
and U7109 (N_7109,N_5690,N_5995);
nand U7110 (N_7110,N_6104,N_5603);
and U7111 (N_7111,N_5853,N_6015);
nand U7112 (N_7112,N_6131,N_5690);
nor U7113 (N_7113,N_5914,N_5864);
and U7114 (N_7114,N_5861,N_5796);
nor U7115 (N_7115,N_6284,N_6159);
nand U7116 (N_7116,N_5938,N_6301);
or U7117 (N_7117,N_6366,N_5968);
xnor U7118 (N_7118,N_5615,N_6336);
nand U7119 (N_7119,N_5775,N_6087);
or U7120 (N_7120,N_5792,N_6084);
or U7121 (N_7121,N_6338,N_6356);
and U7122 (N_7122,N_6042,N_5975);
nor U7123 (N_7123,N_5623,N_5903);
nand U7124 (N_7124,N_6348,N_5846);
xnor U7125 (N_7125,N_6298,N_5976);
xnor U7126 (N_7126,N_6286,N_6098);
xnor U7127 (N_7127,N_5776,N_6147);
and U7128 (N_7128,N_6327,N_6361);
xnor U7129 (N_7129,N_6300,N_5630);
or U7130 (N_7130,N_5670,N_6135);
nor U7131 (N_7131,N_6362,N_6260);
xor U7132 (N_7132,N_5983,N_5748);
or U7133 (N_7133,N_5990,N_5671);
or U7134 (N_7134,N_6262,N_6198);
or U7135 (N_7135,N_6277,N_5836);
or U7136 (N_7136,N_5900,N_6062);
nand U7137 (N_7137,N_6127,N_5906);
or U7138 (N_7138,N_6107,N_5640);
and U7139 (N_7139,N_5833,N_5825);
and U7140 (N_7140,N_6006,N_6305);
or U7141 (N_7141,N_5863,N_5661);
nand U7142 (N_7142,N_5628,N_5909);
and U7143 (N_7143,N_5671,N_6166);
xor U7144 (N_7144,N_6089,N_6237);
and U7145 (N_7145,N_5803,N_6172);
xor U7146 (N_7146,N_5614,N_6266);
and U7147 (N_7147,N_6225,N_6284);
nor U7148 (N_7148,N_6274,N_6234);
nor U7149 (N_7149,N_6220,N_6035);
xor U7150 (N_7150,N_5869,N_5911);
nand U7151 (N_7151,N_6345,N_5632);
and U7152 (N_7152,N_5743,N_6343);
or U7153 (N_7153,N_5690,N_6240);
nor U7154 (N_7154,N_5681,N_5652);
or U7155 (N_7155,N_6163,N_6256);
nor U7156 (N_7156,N_6171,N_5887);
nor U7157 (N_7157,N_6089,N_6159);
xor U7158 (N_7158,N_5895,N_6275);
xor U7159 (N_7159,N_6037,N_5634);
and U7160 (N_7160,N_6039,N_6126);
or U7161 (N_7161,N_5712,N_5634);
and U7162 (N_7162,N_6082,N_5642);
or U7163 (N_7163,N_6349,N_6365);
or U7164 (N_7164,N_6339,N_6397);
and U7165 (N_7165,N_6173,N_6287);
nand U7166 (N_7166,N_6348,N_5764);
or U7167 (N_7167,N_6275,N_5691);
xnor U7168 (N_7168,N_6174,N_6259);
or U7169 (N_7169,N_6320,N_6081);
nor U7170 (N_7170,N_5838,N_5781);
and U7171 (N_7171,N_5937,N_5722);
nor U7172 (N_7172,N_6231,N_6169);
nor U7173 (N_7173,N_5763,N_5866);
nand U7174 (N_7174,N_5789,N_5898);
or U7175 (N_7175,N_5669,N_6296);
xor U7176 (N_7176,N_5962,N_6315);
or U7177 (N_7177,N_6174,N_6225);
or U7178 (N_7178,N_5760,N_6386);
and U7179 (N_7179,N_5828,N_5800);
and U7180 (N_7180,N_6102,N_6345);
nor U7181 (N_7181,N_5837,N_6039);
nor U7182 (N_7182,N_6213,N_5910);
nand U7183 (N_7183,N_5748,N_6164);
nor U7184 (N_7184,N_5856,N_5688);
nor U7185 (N_7185,N_6140,N_5830);
nand U7186 (N_7186,N_5619,N_6176);
or U7187 (N_7187,N_5764,N_5854);
or U7188 (N_7188,N_5751,N_6373);
or U7189 (N_7189,N_5876,N_5780);
xor U7190 (N_7190,N_5689,N_5927);
and U7191 (N_7191,N_5812,N_5773);
nor U7192 (N_7192,N_6328,N_5844);
nor U7193 (N_7193,N_6351,N_5661);
and U7194 (N_7194,N_6067,N_5899);
or U7195 (N_7195,N_5763,N_5600);
nor U7196 (N_7196,N_6032,N_6291);
and U7197 (N_7197,N_6150,N_5736);
xor U7198 (N_7198,N_6043,N_5975);
xor U7199 (N_7199,N_6016,N_5891);
nand U7200 (N_7200,N_6932,N_6557);
and U7201 (N_7201,N_6729,N_6969);
and U7202 (N_7202,N_6825,N_7020);
nand U7203 (N_7203,N_7133,N_6527);
or U7204 (N_7204,N_7116,N_6695);
xor U7205 (N_7205,N_6828,N_6912);
and U7206 (N_7206,N_6673,N_6631);
or U7207 (N_7207,N_6649,N_6995);
or U7208 (N_7208,N_6724,N_6730);
nor U7209 (N_7209,N_6606,N_6589);
and U7210 (N_7210,N_6402,N_7087);
nand U7211 (N_7211,N_7148,N_6526);
xnor U7212 (N_7212,N_6771,N_7139);
or U7213 (N_7213,N_6736,N_6652);
nand U7214 (N_7214,N_6563,N_6561);
and U7215 (N_7215,N_6778,N_6613);
and U7216 (N_7216,N_6927,N_6740);
xor U7217 (N_7217,N_6566,N_7153);
xor U7218 (N_7218,N_7049,N_6734);
or U7219 (N_7219,N_6731,N_7100);
nand U7220 (N_7220,N_7007,N_7104);
and U7221 (N_7221,N_6627,N_7054);
and U7222 (N_7222,N_7085,N_6752);
xnor U7223 (N_7223,N_6821,N_6493);
and U7224 (N_7224,N_6915,N_6438);
xnor U7225 (N_7225,N_6766,N_6772);
xnor U7226 (N_7226,N_6898,N_6586);
nand U7227 (N_7227,N_6474,N_7015);
or U7228 (N_7228,N_6776,N_6416);
or U7229 (N_7229,N_7137,N_6931);
and U7230 (N_7230,N_6419,N_7109);
or U7231 (N_7231,N_6491,N_6986);
xnor U7232 (N_7232,N_7154,N_6536);
and U7233 (N_7233,N_6788,N_6868);
or U7234 (N_7234,N_6988,N_6899);
nand U7235 (N_7235,N_6540,N_6494);
and U7236 (N_7236,N_7019,N_6668);
nand U7237 (N_7237,N_6404,N_6829);
and U7238 (N_7238,N_6853,N_6807);
and U7239 (N_7239,N_6692,N_6746);
or U7240 (N_7240,N_7121,N_6948);
nor U7241 (N_7241,N_6694,N_7122);
xnor U7242 (N_7242,N_6794,N_7163);
nor U7243 (N_7243,N_6897,N_6591);
nor U7244 (N_7244,N_6654,N_7075);
or U7245 (N_7245,N_6637,N_7021);
or U7246 (N_7246,N_6625,N_6926);
nor U7247 (N_7247,N_7026,N_6508);
or U7248 (N_7248,N_6959,N_6859);
xor U7249 (N_7249,N_6601,N_6733);
nand U7250 (N_7250,N_7061,N_6976);
or U7251 (N_7251,N_6789,N_6609);
and U7252 (N_7252,N_7056,N_7016);
nand U7253 (N_7253,N_7002,N_6640);
nor U7254 (N_7254,N_6528,N_6618);
and U7255 (N_7255,N_6529,N_6817);
and U7256 (N_7256,N_6780,N_6801);
xnor U7257 (N_7257,N_6887,N_6908);
nand U7258 (N_7258,N_7107,N_7086);
and U7259 (N_7259,N_6764,N_6784);
and U7260 (N_7260,N_6497,N_6935);
xor U7261 (N_7261,N_6579,N_6624);
xnor U7262 (N_7262,N_6571,N_6551);
xnor U7263 (N_7263,N_7017,N_7005);
nor U7264 (N_7264,N_6687,N_6997);
xor U7265 (N_7265,N_6418,N_6934);
nand U7266 (N_7266,N_6775,N_7164);
nor U7267 (N_7267,N_7068,N_7199);
xnor U7268 (N_7268,N_7156,N_6517);
or U7269 (N_7269,N_6822,N_7057);
xnor U7270 (N_7270,N_6857,N_6860);
nand U7271 (N_7271,N_6457,N_7146);
xor U7272 (N_7272,N_6647,N_6412);
nor U7273 (N_7273,N_7080,N_6824);
xnor U7274 (N_7274,N_6975,N_7125);
and U7275 (N_7275,N_6666,N_6515);
and U7276 (N_7276,N_7180,N_7065);
nor U7277 (N_7277,N_6901,N_6851);
or U7278 (N_7278,N_6500,N_7149);
and U7279 (N_7279,N_7012,N_7000);
xnor U7280 (N_7280,N_6442,N_7124);
xnor U7281 (N_7281,N_6599,N_7039);
and U7282 (N_7282,N_6994,N_6506);
or U7283 (N_7283,N_6521,N_6698);
xor U7284 (N_7284,N_6567,N_7053);
or U7285 (N_7285,N_6406,N_6998);
xor U7286 (N_7286,N_7078,N_6578);
nor U7287 (N_7287,N_6799,N_6779);
xor U7288 (N_7288,N_7011,N_6475);
nand U7289 (N_7289,N_6634,N_7120);
xnor U7290 (N_7290,N_6808,N_6786);
nand U7291 (N_7291,N_6811,N_6690);
nor U7292 (N_7292,N_7177,N_6896);
xnor U7293 (N_7293,N_6711,N_6743);
or U7294 (N_7294,N_6888,N_7063);
nor U7295 (N_7295,N_6840,N_6511);
xnor U7296 (N_7296,N_7037,N_6773);
or U7297 (N_7297,N_6476,N_7141);
nor U7298 (N_7298,N_6795,N_6452);
nor U7299 (N_7299,N_7081,N_7031);
and U7300 (N_7300,N_6723,N_7105);
xor U7301 (N_7301,N_6646,N_6530);
nand U7302 (N_7302,N_7188,N_6573);
and U7303 (N_7303,N_6538,N_6620);
nor U7304 (N_7304,N_6558,N_7169);
and U7305 (N_7305,N_6437,N_6481);
or U7306 (N_7306,N_6965,N_6610);
nand U7307 (N_7307,N_7157,N_6676);
nand U7308 (N_7308,N_6655,N_6644);
and U7309 (N_7309,N_6950,N_7167);
or U7310 (N_7310,N_7010,N_6739);
xnor U7311 (N_7311,N_6728,N_6877);
and U7312 (N_7312,N_6993,N_6958);
and U7313 (N_7313,N_7166,N_6804);
nand U7314 (N_7314,N_6914,N_6663);
or U7315 (N_7315,N_6744,N_6623);
nor U7316 (N_7316,N_7052,N_6505);
nor U7317 (N_7317,N_6542,N_6755);
nand U7318 (N_7318,N_7159,N_6922);
xnor U7319 (N_7319,N_6798,N_6876);
or U7320 (N_7320,N_6465,N_7117);
and U7321 (N_7321,N_6466,N_6533);
nand U7322 (N_7322,N_6943,N_6410);
xnor U7323 (N_7323,N_6677,N_6972);
and U7324 (N_7324,N_6405,N_6702);
or U7325 (N_7325,N_6715,N_6524);
and U7326 (N_7326,N_6674,N_6957);
or U7327 (N_7327,N_7115,N_6518);
nor U7328 (N_7328,N_6450,N_6765);
or U7329 (N_7329,N_7191,N_7092);
and U7330 (N_7330,N_6871,N_6832);
nand U7331 (N_7331,N_6544,N_6835);
or U7332 (N_7332,N_6499,N_6565);
nor U7333 (N_7333,N_6662,N_6441);
nor U7334 (N_7334,N_6675,N_7171);
xnor U7335 (N_7335,N_7069,N_7040);
or U7336 (N_7336,N_7082,N_6569);
nor U7337 (N_7337,N_6575,N_6597);
xnor U7338 (N_7338,N_6917,N_7190);
nor U7339 (N_7339,N_6717,N_7132);
and U7340 (N_7340,N_7024,N_6564);
and U7341 (N_7341,N_7138,N_7098);
or U7342 (N_7342,N_6847,N_7055);
nor U7343 (N_7343,N_6459,N_7106);
nor U7344 (N_7344,N_6796,N_6920);
and U7345 (N_7345,N_7030,N_6921);
nor U7346 (N_7346,N_6545,N_6532);
xor U7347 (N_7347,N_6767,N_6440);
nor U7348 (N_7348,N_6495,N_6411);
or U7349 (N_7349,N_6890,N_6882);
nor U7350 (N_7350,N_6971,N_6839);
nand U7351 (N_7351,N_6486,N_7060);
xor U7352 (N_7352,N_7158,N_6885);
xnor U7353 (N_7353,N_6595,N_7102);
and U7354 (N_7354,N_6858,N_6759);
xor U7355 (N_7355,N_6490,N_7168);
xnor U7356 (N_7356,N_7189,N_6903);
nand U7357 (N_7357,N_6464,N_6823);
xnor U7358 (N_7358,N_6705,N_6628);
nor U7359 (N_7359,N_7076,N_6906);
or U7360 (N_7360,N_7088,N_6911);
nor U7361 (N_7361,N_6570,N_6814);
nand U7362 (N_7362,N_6435,N_7046);
nor U7363 (N_7363,N_6797,N_6710);
nand U7364 (N_7364,N_6554,N_6562);
nand U7365 (N_7365,N_7152,N_7155);
or U7366 (N_7366,N_6865,N_6802);
and U7367 (N_7367,N_6461,N_7165);
nor U7368 (N_7368,N_6426,N_6688);
or U7369 (N_7369,N_6421,N_6485);
or U7370 (N_7370,N_6682,N_7091);
xor U7371 (N_7371,N_7062,N_7111);
nand U7372 (N_7372,N_6408,N_7186);
and U7373 (N_7373,N_6856,N_6460);
xnor U7374 (N_7374,N_6576,N_6448);
nor U7375 (N_7375,N_6434,N_6880);
or U7376 (N_7376,N_6718,N_6816);
nand U7377 (N_7377,N_6820,N_6635);
nor U7378 (N_7378,N_6970,N_7130);
and U7379 (N_7379,N_6883,N_6604);
nor U7380 (N_7380,N_6866,N_7084);
xor U7381 (N_7381,N_6552,N_6905);
xor U7382 (N_7382,N_6944,N_6747);
nand U7383 (N_7383,N_6665,N_6608);
xnor U7384 (N_7384,N_6593,N_6872);
or U7385 (N_7385,N_6787,N_6879);
or U7386 (N_7386,N_6633,N_6977);
and U7387 (N_7387,N_6407,N_7013);
nand U7388 (N_7388,N_6621,N_6661);
xor U7389 (N_7389,N_6458,N_6598);
and U7390 (N_7390,N_7140,N_6791);
or U7391 (N_7391,N_6479,N_6725);
or U7392 (N_7392,N_6657,N_7004);
or U7393 (N_7393,N_6732,N_7147);
xnor U7394 (N_7394,N_6722,N_7018);
and U7395 (N_7395,N_6769,N_6619);
xor U7396 (N_7396,N_7198,N_7066);
or U7397 (N_7397,N_6684,N_6987);
xor U7398 (N_7398,N_7033,N_6881);
xor U7399 (N_7399,N_6547,N_6472);
xor U7400 (N_7400,N_6584,N_6894);
nor U7401 (N_7401,N_7173,N_7058);
nor U7402 (N_7402,N_7006,N_6504);
xnor U7403 (N_7403,N_6838,N_6955);
and U7404 (N_7404,N_7027,N_6946);
xnor U7405 (N_7405,N_6819,N_7064);
and U7406 (N_7406,N_6826,N_6895);
xnor U7407 (N_7407,N_6594,N_6503);
nor U7408 (N_7408,N_7113,N_6742);
nand U7409 (N_7409,N_6423,N_7048);
or U7410 (N_7410,N_6471,N_7036);
nand U7411 (N_7411,N_6774,N_6468);
nand U7412 (N_7412,N_6942,N_6873);
or U7413 (N_7413,N_6793,N_7083);
nand U7414 (N_7414,N_6629,N_6548);
or U7415 (N_7415,N_6681,N_6444);
nand U7416 (N_7416,N_6549,N_6933);
nor U7417 (N_7417,N_6680,N_6781);
or U7418 (N_7418,N_7182,N_7129);
nand U7419 (N_7419,N_7150,N_6445);
xor U7420 (N_7420,N_6745,N_6964);
nand U7421 (N_7421,N_6630,N_6727);
or U7422 (N_7422,N_6583,N_6487);
and U7423 (N_7423,N_6522,N_6537);
nor U7424 (N_7424,N_7044,N_7176);
xor U7425 (N_7425,N_6884,N_6941);
nor U7426 (N_7426,N_6449,N_6510);
xor U7427 (N_7427,N_7143,N_7008);
nor U7428 (N_7428,N_6430,N_6439);
xnor U7429 (N_7429,N_6667,N_6845);
xnor U7430 (N_7430,N_7183,N_7151);
xor U7431 (N_7431,N_6979,N_6966);
nor U7432 (N_7432,N_7038,N_6842);
or U7433 (N_7433,N_6520,N_6930);
xnor U7434 (N_7434,N_7022,N_6480);
or U7435 (N_7435,N_7035,N_7134);
nand U7436 (N_7436,N_6612,N_7043);
nand U7437 (N_7437,N_6909,N_6470);
or U7438 (N_7438,N_6812,N_6645);
xor U7439 (N_7439,N_6611,N_6753);
or U7440 (N_7440,N_7095,N_6737);
and U7441 (N_7441,N_6716,N_6703);
and U7442 (N_7442,N_6422,N_6900);
nand U7443 (N_7443,N_6642,N_7029);
and U7444 (N_7444,N_6617,N_6514);
nor U7445 (N_7445,N_6854,N_6425);
and U7446 (N_7446,N_6632,N_6990);
nand U7447 (N_7447,N_7074,N_7123);
xnor U7448 (N_7448,N_6961,N_6818);
xor U7449 (N_7449,N_6451,N_6719);
or U7450 (N_7450,N_6862,N_7090);
and U7451 (N_7451,N_6815,N_6937);
nand U7452 (N_7452,N_6462,N_6656);
nor U7453 (N_7453,N_7050,N_6580);
nor U7454 (N_7454,N_6659,N_6726);
nand U7455 (N_7455,N_6953,N_6874);
nand U7456 (N_7456,N_6701,N_6837);
or U7457 (N_7457,N_6768,N_6800);
and U7458 (N_7458,N_6918,N_7023);
xnor U7459 (N_7459,N_6539,N_6588);
nor U7460 (N_7460,N_6803,N_6864);
nand U7461 (N_7461,N_6770,N_6525);
nor U7462 (N_7462,N_7195,N_6678);
or U7463 (N_7463,N_6913,N_6446);
or U7464 (N_7464,N_6670,N_7172);
nor U7465 (N_7465,N_7135,N_6429);
and U7466 (N_7466,N_6827,N_6456);
nor U7467 (N_7467,N_6830,N_6555);
nor U7468 (N_7468,N_6886,N_6919);
and U7469 (N_7469,N_6891,N_6844);
and U7470 (N_7470,N_6978,N_6685);
nor U7471 (N_7471,N_6581,N_6974);
nor U7472 (N_7472,N_6714,N_6869);
or U7473 (N_7473,N_6850,N_6409);
nand U7474 (N_7474,N_6641,N_6478);
nand U7475 (N_7475,N_6841,N_6484);
nor U7476 (N_7476,N_6910,N_7059);
and U7477 (N_7477,N_6720,N_6924);
and U7478 (N_7478,N_6424,N_6651);
nand U7479 (N_7479,N_6763,N_6916);
or U7480 (N_7480,N_7093,N_6704);
xor U7481 (N_7481,N_7034,N_6400);
or U7482 (N_7482,N_6488,N_6420);
nand U7483 (N_7483,N_6512,N_6693);
nor U7484 (N_7484,N_7014,N_6636);
and U7485 (N_7485,N_6738,N_6639);
or U7486 (N_7486,N_6754,N_6498);
xnor U7487 (N_7487,N_6980,N_6697);
xor U7488 (N_7488,N_7070,N_6574);
nand U7489 (N_7489,N_6721,N_7028);
nor U7490 (N_7490,N_6492,N_6983);
nand U7491 (N_7491,N_6653,N_6550);
nand U7492 (N_7492,N_6749,N_7073);
and U7493 (N_7493,N_6699,N_6432);
nand U7494 (N_7494,N_7131,N_6758);
and U7495 (N_7495,N_6572,N_6892);
or U7496 (N_7496,N_6928,N_6401);
or U7497 (N_7497,N_6756,N_6750);
or U7498 (N_7498,N_6785,N_7119);
nor U7499 (N_7499,N_7089,N_6945);
nor U7500 (N_7500,N_6939,N_6672);
nor U7501 (N_7501,N_7142,N_7009);
nand U7502 (N_7502,N_6686,N_7077);
or U7503 (N_7503,N_7160,N_7175);
and U7504 (N_7504,N_7194,N_6664);
or U7505 (N_7505,N_6556,N_6870);
nand U7506 (N_7506,N_7118,N_6483);
nand U7507 (N_7507,N_7185,N_6952);
nand U7508 (N_7508,N_6519,N_6951);
xnor U7509 (N_7509,N_6960,N_6985);
nand U7510 (N_7510,N_7025,N_7067);
and U7511 (N_7511,N_6454,N_6560);
and U7512 (N_7512,N_6473,N_6683);
xnor U7513 (N_7513,N_6638,N_6616);
xnor U7514 (N_7514,N_6805,N_6614);
xnor U7515 (N_7515,N_6605,N_7001);
nor U7516 (N_7516,N_7184,N_6954);
nor U7517 (N_7517,N_6989,N_7045);
nor U7518 (N_7518,N_6843,N_6534);
nor U7519 (N_7519,N_6467,N_6689);
and U7520 (N_7520,N_6417,N_7193);
nand U7521 (N_7521,N_7072,N_6741);
or U7522 (N_7522,N_6582,N_6502);
and U7523 (N_7523,N_6650,N_7197);
nor U7524 (N_7524,N_6809,N_6496);
xor U7525 (N_7525,N_6709,N_6777);
nor U7526 (N_7526,N_6938,N_6516);
and U7527 (N_7527,N_7110,N_6783);
xor U7528 (N_7528,N_6999,N_6708);
xnor U7529 (N_7529,N_6751,N_6696);
nor U7530 (N_7530,N_6996,N_7003);
and U7531 (N_7531,N_7178,N_6615);
nand U7532 (N_7532,N_7071,N_6902);
xor U7533 (N_7533,N_7181,N_6691);
and U7534 (N_7534,N_6669,N_7097);
xnor U7535 (N_7535,N_6836,N_6600);
xnor U7536 (N_7536,N_7103,N_6559);
and U7537 (N_7537,N_7099,N_6507);
nand U7538 (N_7538,N_6431,N_7170);
xnor U7539 (N_7539,N_7144,N_6603);
or U7540 (N_7540,N_6992,N_6907);
xnor U7541 (N_7541,N_6607,N_6867);
and U7542 (N_7542,N_6501,N_6443);
xnor U7543 (N_7543,N_6735,N_7162);
xor U7544 (N_7544,N_6553,N_6956);
and U7545 (N_7545,N_6535,N_7196);
nand U7546 (N_7546,N_6543,N_6968);
nand U7547 (N_7547,N_7161,N_6602);
or U7548 (N_7548,N_6587,N_6622);
or U7549 (N_7549,N_6413,N_6878);
nand U7550 (N_7550,N_6967,N_6577);
or U7551 (N_7551,N_6469,N_6427);
and U7552 (N_7552,N_6833,N_6523);
nor U7553 (N_7553,N_7051,N_6541);
xnor U7554 (N_7554,N_6660,N_6893);
xnor U7555 (N_7555,N_6671,N_7047);
nand U7556 (N_7556,N_7108,N_6707);
or U7557 (N_7557,N_6706,N_6596);
and U7558 (N_7558,N_6863,N_6648);
or U7559 (N_7559,N_6834,N_7096);
nor U7560 (N_7560,N_6904,N_6782);
or U7561 (N_7561,N_6590,N_6949);
nor U7562 (N_7562,N_6455,N_6806);
nand U7563 (N_7563,N_7192,N_6415);
or U7564 (N_7564,N_7032,N_6463);
xnor U7565 (N_7565,N_6585,N_6973);
xor U7566 (N_7566,N_6875,N_6509);
nand U7567 (N_7567,N_6991,N_6813);
xor U7568 (N_7568,N_6482,N_7174);
or U7569 (N_7569,N_6700,N_6852);
xor U7570 (N_7570,N_6940,N_6403);
and U7571 (N_7571,N_6433,N_6981);
nor U7572 (N_7572,N_6849,N_7145);
nor U7573 (N_7573,N_6489,N_6923);
or U7574 (N_7574,N_6658,N_7179);
xnor U7575 (N_7575,N_6453,N_7128);
and U7576 (N_7576,N_6984,N_7136);
nor U7577 (N_7577,N_6592,N_6846);
xor U7578 (N_7578,N_6929,N_6762);
nor U7579 (N_7579,N_6477,N_6761);
or U7580 (N_7580,N_7127,N_6889);
nor U7581 (N_7581,N_6936,N_6414);
or U7582 (N_7582,N_6855,N_6982);
xor U7583 (N_7583,N_6643,N_6790);
and U7584 (N_7584,N_6428,N_6531);
or U7585 (N_7585,N_6757,N_7041);
nand U7586 (N_7586,N_6792,N_6436);
or U7587 (N_7587,N_7126,N_6947);
nand U7588 (N_7588,N_7042,N_7101);
nor U7589 (N_7589,N_7187,N_6925);
xor U7590 (N_7590,N_6810,N_6713);
and U7591 (N_7591,N_7094,N_6760);
or U7592 (N_7592,N_6447,N_6568);
and U7593 (N_7593,N_6962,N_6546);
xor U7594 (N_7594,N_6831,N_6679);
nand U7595 (N_7595,N_6861,N_6626);
xor U7596 (N_7596,N_6748,N_7079);
or U7597 (N_7597,N_6848,N_6513);
xor U7598 (N_7598,N_6963,N_6712);
nor U7599 (N_7599,N_7114,N_7112);
nand U7600 (N_7600,N_6789,N_7190);
xnor U7601 (N_7601,N_6560,N_7115);
nor U7602 (N_7602,N_6995,N_6842);
and U7603 (N_7603,N_7046,N_6616);
nand U7604 (N_7604,N_6596,N_6925);
nand U7605 (N_7605,N_6580,N_7143);
or U7606 (N_7606,N_6629,N_6878);
nor U7607 (N_7607,N_6453,N_6415);
and U7608 (N_7608,N_6819,N_6765);
xnor U7609 (N_7609,N_6883,N_6983);
xor U7610 (N_7610,N_6675,N_6543);
xnor U7611 (N_7611,N_6752,N_6713);
and U7612 (N_7612,N_6559,N_6861);
nor U7613 (N_7613,N_6997,N_6607);
or U7614 (N_7614,N_7057,N_6778);
and U7615 (N_7615,N_6866,N_6832);
nand U7616 (N_7616,N_6933,N_6415);
nor U7617 (N_7617,N_6564,N_7081);
xnor U7618 (N_7618,N_6907,N_6851);
xnor U7619 (N_7619,N_6531,N_6732);
xnor U7620 (N_7620,N_6627,N_6751);
nor U7621 (N_7621,N_6830,N_6632);
or U7622 (N_7622,N_7095,N_6983);
nand U7623 (N_7623,N_6670,N_6522);
and U7624 (N_7624,N_7009,N_7139);
nor U7625 (N_7625,N_6745,N_7084);
and U7626 (N_7626,N_7138,N_6966);
nor U7627 (N_7627,N_6742,N_6451);
nor U7628 (N_7628,N_6592,N_7193);
and U7629 (N_7629,N_6742,N_7079);
nor U7630 (N_7630,N_7034,N_6808);
and U7631 (N_7631,N_6810,N_7038);
xnor U7632 (N_7632,N_6931,N_6588);
and U7633 (N_7633,N_7074,N_6660);
nand U7634 (N_7634,N_7161,N_6600);
nor U7635 (N_7635,N_6676,N_6817);
nand U7636 (N_7636,N_6845,N_6456);
nor U7637 (N_7637,N_6909,N_6799);
nand U7638 (N_7638,N_6740,N_6723);
and U7639 (N_7639,N_6754,N_6862);
or U7640 (N_7640,N_6604,N_7097);
or U7641 (N_7641,N_7031,N_7102);
xor U7642 (N_7642,N_7111,N_6798);
xnor U7643 (N_7643,N_6404,N_7174);
and U7644 (N_7644,N_6472,N_6785);
nor U7645 (N_7645,N_6444,N_7189);
nor U7646 (N_7646,N_6418,N_6501);
nor U7647 (N_7647,N_6547,N_7149);
or U7648 (N_7648,N_6955,N_6525);
or U7649 (N_7649,N_6887,N_7114);
xor U7650 (N_7650,N_6536,N_7042);
or U7651 (N_7651,N_6782,N_6872);
or U7652 (N_7652,N_7028,N_7123);
nor U7653 (N_7653,N_6595,N_7119);
nand U7654 (N_7654,N_6682,N_6868);
and U7655 (N_7655,N_6530,N_7026);
and U7656 (N_7656,N_6732,N_6647);
and U7657 (N_7657,N_7175,N_7100);
xnor U7658 (N_7658,N_6844,N_7085);
and U7659 (N_7659,N_6929,N_6939);
nor U7660 (N_7660,N_6487,N_6428);
nand U7661 (N_7661,N_7108,N_6924);
and U7662 (N_7662,N_6540,N_7160);
or U7663 (N_7663,N_6916,N_6886);
nand U7664 (N_7664,N_6864,N_7016);
xnor U7665 (N_7665,N_7060,N_6521);
or U7666 (N_7666,N_6956,N_6656);
and U7667 (N_7667,N_7016,N_7034);
and U7668 (N_7668,N_7067,N_6410);
nand U7669 (N_7669,N_7016,N_6957);
nor U7670 (N_7670,N_6682,N_6801);
or U7671 (N_7671,N_7195,N_6639);
or U7672 (N_7672,N_6473,N_6434);
nand U7673 (N_7673,N_6974,N_6731);
or U7674 (N_7674,N_7172,N_6574);
xnor U7675 (N_7675,N_6443,N_6759);
and U7676 (N_7676,N_6816,N_6782);
nor U7677 (N_7677,N_6482,N_6764);
and U7678 (N_7678,N_6551,N_6827);
xnor U7679 (N_7679,N_6933,N_6735);
and U7680 (N_7680,N_7128,N_6505);
xor U7681 (N_7681,N_7166,N_6945);
nor U7682 (N_7682,N_6501,N_6820);
nand U7683 (N_7683,N_6829,N_6828);
nand U7684 (N_7684,N_6432,N_6422);
or U7685 (N_7685,N_6696,N_6475);
xnor U7686 (N_7686,N_6499,N_6919);
xor U7687 (N_7687,N_6883,N_6700);
xor U7688 (N_7688,N_6560,N_7085);
nand U7689 (N_7689,N_7104,N_7003);
nor U7690 (N_7690,N_6784,N_6419);
nor U7691 (N_7691,N_6954,N_7092);
nand U7692 (N_7692,N_6996,N_6897);
xnor U7693 (N_7693,N_6426,N_6592);
or U7694 (N_7694,N_6417,N_7118);
or U7695 (N_7695,N_6617,N_6482);
xnor U7696 (N_7696,N_6739,N_6906);
nor U7697 (N_7697,N_6850,N_6400);
nand U7698 (N_7698,N_6802,N_6685);
and U7699 (N_7699,N_6486,N_6989);
nand U7700 (N_7700,N_6692,N_6487);
and U7701 (N_7701,N_6917,N_6747);
xnor U7702 (N_7702,N_6657,N_6733);
and U7703 (N_7703,N_6801,N_6843);
nand U7704 (N_7704,N_6484,N_7023);
nand U7705 (N_7705,N_7084,N_7104);
and U7706 (N_7706,N_6947,N_6748);
or U7707 (N_7707,N_6875,N_6587);
nand U7708 (N_7708,N_6484,N_6433);
and U7709 (N_7709,N_6854,N_7144);
nor U7710 (N_7710,N_7096,N_6935);
xor U7711 (N_7711,N_7149,N_7090);
nor U7712 (N_7712,N_7029,N_6767);
or U7713 (N_7713,N_6788,N_6505);
nand U7714 (N_7714,N_6590,N_6475);
or U7715 (N_7715,N_6595,N_6707);
or U7716 (N_7716,N_7121,N_6491);
nor U7717 (N_7717,N_6997,N_6975);
xor U7718 (N_7718,N_7004,N_7003);
nor U7719 (N_7719,N_6672,N_6826);
nand U7720 (N_7720,N_6787,N_7003);
nor U7721 (N_7721,N_6528,N_6489);
nand U7722 (N_7722,N_7139,N_6495);
nor U7723 (N_7723,N_6875,N_6578);
or U7724 (N_7724,N_7058,N_6894);
or U7725 (N_7725,N_7190,N_7170);
and U7726 (N_7726,N_6466,N_7126);
nand U7727 (N_7727,N_6516,N_6659);
or U7728 (N_7728,N_6898,N_6627);
or U7729 (N_7729,N_6719,N_6730);
nor U7730 (N_7730,N_6859,N_6743);
nor U7731 (N_7731,N_7074,N_7084);
nand U7732 (N_7732,N_6457,N_6756);
nor U7733 (N_7733,N_6931,N_6690);
nor U7734 (N_7734,N_6859,N_6535);
or U7735 (N_7735,N_6782,N_6900);
and U7736 (N_7736,N_6528,N_6594);
or U7737 (N_7737,N_6981,N_6595);
or U7738 (N_7738,N_6588,N_7143);
xnor U7739 (N_7739,N_7058,N_6721);
nor U7740 (N_7740,N_6594,N_6576);
xor U7741 (N_7741,N_6561,N_6949);
and U7742 (N_7742,N_6768,N_6738);
and U7743 (N_7743,N_7070,N_6622);
nor U7744 (N_7744,N_6525,N_6934);
nor U7745 (N_7745,N_7108,N_6840);
or U7746 (N_7746,N_6904,N_7055);
nor U7747 (N_7747,N_6545,N_6651);
or U7748 (N_7748,N_6574,N_7164);
or U7749 (N_7749,N_6774,N_6656);
and U7750 (N_7750,N_6557,N_6900);
or U7751 (N_7751,N_6661,N_7073);
or U7752 (N_7752,N_6409,N_6642);
nand U7753 (N_7753,N_6594,N_6443);
xor U7754 (N_7754,N_6516,N_6504);
and U7755 (N_7755,N_6939,N_7117);
and U7756 (N_7756,N_6964,N_6751);
xnor U7757 (N_7757,N_6826,N_6671);
nor U7758 (N_7758,N_7071,N_6738);
and U7759 (N_7759,N_6944,N_6672);
nand U7760 (N_7760,N_6813,N_6695);
xor U7761 (N_7761,N_7079,N_6970);
and U7762 (N_7762,N_6417,N_6530);
or U7763 (N_7763,N_6445,N_6767);
or U7764 (N_7764,N_6745,N_6653);
xor U7765 (N_7765,N_6631,N_6475);
and U7766 (N_7766,N_6404,N_7046);
or U7767 (N_7767,N_6415,N_6948);
or U7768 (N_7768,N_6979,N_7123);
nor U7769 (N_7769,N_7106,N_7126);
and U7770 (N_7770,N_6730,N_6673);
nand U7771 (N_7771,N_6831,N_7021);
nand U7772 (N_7772,N_6728,N_6846);
nand U7773 (N_7773,N_6660,N_7158);
or U7774 (N_7774,N_6907,N_6630);
nand U7775 (N_7775,N_6893,N_7158);
nand U7776 (N_7776,N_6961,N_6893);
nand U7777 (N_7777,N_6952,N_6602);
or U7778 (N_7778,N_7150,N_7060);
or U7779 (N_7779,N_6917,N_6927);
nand U7780 (N_7780,N_6598,N_6940);
nand U7781 (N_7781,N_6926,N_6716);
or U7782 (N_7782,N_6671,N_6631);
or U7783 (N_7783,N_7122,N_7044);
nor U7784 (N_7784,N_6601,N_6824);
and U7785 (N_7785,N_7117,N_6562);
and U7786 (N_7786,N_6975,N_6596);
nand U7787 (N_7787,N_7115,N_6708);
and U7788 (N_7788,N_6965,N_6872);
nor U7789 (N_7789,N_6574,N_7138);
or U7790 (N_7790,N_6771,N_6426);
or U7791 (N_7791,N_7017,N_7111);
or U7792 (N_7792,N_7158,N_6873);
and U7793 (N_7793,N_6630,N_6666);
and U7794 (N_7794,N_6497,N_7137);
nor U7795 (N_7795,N_6728,N_6559);
xor U7796 (N_7796,N_6872,N_6679);
and U7797 (N_7797,N_6822,N_6854);
or U7798 (N_7798,N_6874,N_6643);
xnor U7799 (N_7799,N_7114,N_6832);
or U7800 (N_7800,N_6637,N_6480);
xor U7801 (N_7801,N_6763,N_7054);
or U7802 (N_7802,N_6747,N_6595);
xnor U7803 (N_7803,N_6515,N_6424);
nand U7804 (N_7804,N_6693,N_6481);
xor U7805 (N_7805,N_6633,N_6483);
nor U7806 (N_7806,N_6955,N_7171);
and U7807 (N_7807,N_6415,N_6763);
xnor U7808 (N_7808,N_7155,N_7028);
and U7809 (N_7809,N_6844,N_6438);
nand U7810 (N_7810,N_6667,N_6490);
nor U7811 (N_7811,N_6632,N_6598);
nor U7812 (N_7812,N_6494,N_6437);
xnor U7813 (N_7813,N_6768,N_7095);
xor U7814 (N_7814,N_6595,N_6783);
nand U7815 (N_7815,N_6718,N_7178);
or U7816 (N_7816,N_7067,N_6945);
xor U7817 (N_7817,N_6571,N_6836);
xor U7818 (N_7818,N_6709,N_6976);
xor U7819 (N_7819,N_6762,N_6766);
and U7820 (N_7820,N_7191,N_6518);
and U7821 (N_7821,N_6745,N_6715);
or U7822 (N_7822,N_6559,N_7140);
or U7823 (N_7823,N_6994,N_6950);
xor U7824 (N_7824,N_6494,N_6481);
nor U7825 (N_7825,N_7132,N_6526);
and U7826 (N_7826,N_7019,N_6459);
or U7827 (N_7827,N_7099,N_6473);
nand U7828 (N_7828,N_6835,N_6596);
or U7829 (N_7829,N_6414,N_6475);
and U7830 (N_7830,N_6499,N_6816);
xnor U7831 (N_7831,N_7138,N_6720);
and U7832 (N_7832,N_6493,N_6794);
or U7833 (N_7833,N_7126,N_6989);
nand U7834 (N_7834,N_6695,N_6635);
or U7835 (N_7835,N_6537,N_6685);
and U7836 (N_7836,N_6869,N_6809);
xor U7837 (N_7837,N_6554,N_7078);
nor U7838 (N_7838,N_6577,N_6858);
and U7839 (N_7839,N_7141,N_6847);
nor U7840 (N_7840,N_6618,N_6787);
nor U7841 (N_7841,N_7089,N_6919);
xor U7842 (N_7842,N_7157,N_6709);
nand U7843 (N_7843,N_6480,N_6828);
and U7844 (N_7844,N_7097,N_6963);
and U7845 (N_7845,N_7133,N_6626);
and U7846 (N_7846,N_6692,N_7152);
nand U7847 (N_7847,N_6532,N_6741);
and U7848 (N_7848,N_6614,N_7109);
xnor U7849 (N_7849,N_6560,N_6670);
and U7850 (N_7850,N_6548,N_7037);
or U7851 (N_7851,N_7118,N_6906);
nand U7852 (N_7852,N_6844,N_6847);
and U7853 (N_7853,N_6539,N_6998);
and U7854 (N_7854,N_6560,N_6710);
nand U7855 (N_7855,N_7101,N_6594);
or U7856 (N_7856,N_6447,N_6717);
and U7857 (N_7857,N_6602,N_6415);
or U7858 (N_7858,N_6675,N_6900);
xnor U7859 (N_7859,N_7057,N_6432);
and U7860 (N_7860,N_6859,N_6421);
and U7861 (N_7861,N_6780,N_7096);
or U7862 (N_7862,N_7194,N_6818);
or U7863 (N_7863,N_6832,N_6707);
or U7864 (N_7864,N_7168,N_6619);
or U7865 (N_7865,N_7065,N_7056);
or U7866 (N_7866,N_7020,N_6798);
nand U7867 (N_7867,N_6498,N_6789);
xnor U7868 (N_7868,N_6658,N_7012);
xor U7869 (N_7869,N_6763,N_7125);
or U7870 (N_7870,N_7164,N_6806);
xor U7871 (N_7871,N_7153,N_7171);
and U7872 (N_7872,N_6878,N_6447);
nand U7873 (N_7873,N_6505,N_6799);
nor U7874 (N_7874,N_6458,N_6675);
xor U7875 (N_7875,N_7019,N_6774);
or U7876 (N_7876,N_6709,N_6497);
nor U7877 (N_7877,N_6974,N_6851);
or U7878 (N_7878,N_6757,N_6454);
xnor U7879 (N_7879,N_6637,N_6823);
nor U7880 (N_7880,N_6521,N_6486);
or U7881 (N_7881,N_6545,N_6827);
nor U7882 (N_7882,N_6658,N_6646);
nor U7883 (N_7883,N_6534,N_6997);
nand U7884 (N_7884,N_6639,N_6758);
and U7885 (N_7885,N_7063,N_6518);
nor U7886 (N_7886,N_6576,N_7032);
and U7887 (N_7887,N_6436,N_6935);
and U7888 (N_7888,N_7120,N_7164);
nor U7889 (N_7889,N_7059,N_6654);
or U7890 (N_7890,N_7101,N_6785);
nand U7891 (N_7891,N_6849,N_6739);
nor U7892 (N_7892,N_7196,N_7031);
xnor U7893 (N_7893,N_6920,N_6795);
or U7894 (N_7894,N_6494,N_7171);
nor U7895 (N_7895,N_7175,N_6888);
nand U7896 (N_7896,N_6891,N_6442);
xor U7897 (N_7897,N_6888,N_6897);
nor U7898 (N_7898,N_7173,N_6792);
xnor U7899 (N_7899,N_6699,N_6570);
or U7900 (N_7900,N_6843,N_6762);
and U7901 (N_7901,N_6824,N_7097);
and U7902 (N_7902,N_7130,N_6486);
or U7903 (N_7903,N_7132,N_7062);
nor U7904 (N_7904,N_6628,N_6816);
xnor U7905 (N_7905,N_6704,N_6524);
and U7906 (N_7906,N_6975,N_7181);
nor U7907 (N_7907,N_6839,N_6895);
xor U7908 (N_7908,N_6836,N_6749);
xor U7909 (N_7909,N_6401,N_6499);
xnor U7910 (N_7910,N_6687,N_6972);
or U7911 (N_7911,N_7155,N_6903);
nor U7912 (N_7912,N_7017,N_6515);
nand U7913 (N_7913,N_6813,N_7028);
nor U7914 (N_7914,N_6881,N_6970);
and U7915 (N_7915,N_7070,N_6894);
nor U7916 (N_7916,N_7066,N_6446);
nand U7917 (N_7917,N_6837,N_6504);
xnor U7918 (N_7918,N_7029,N_6758);
nor U7919 (N_7919,N_6896,N_6994);
nand U7920 (N_7920,N_7152,N_7087);
nand U7921 (N_7921,N_6899,N_6871);
nor U7922 (N_7922,N_7108,N_7008);
nand U7923 (N_7923,N_6700,N_6632);
or U7924 (N_7924,N_6710,N_6501);
nand U7925 (N_7925,N_6724,N_6964);
xor U7926 (N_7926,N_6811,N_6442);
nor U7927 (N_7927,N_7016,N_6850);
or U7928 (N_7928,N_6509,N_7180);
xor U7929 (N_7929,N_6453,N_7072);
nor U7930 (N_7930,N_6699,N_6654);
and U7931 (N_7931,N_6869,N_6721);
and U7932 (N_7932,N_7143,N_7088);
nor U7933 (N_7933,N_6744,N_6579);
nand U7934 (N_7934,N_6896,N_6586);
or U7935 (N_7935,N_6802,N_6972);
nor U7936 (N_7936,N_6485,N_7156);
or U7937 (N_7937,N_6715,N_7135);
and U7938 (N_7938,N_6628,N_6561);
nand U7939 (N_7939,N_7084,N_6748);
or U7940 (N_7940,N_6703,N_6569);
or U7941 (N_7941,N_6416,N_6716);
xnor U7942 (N_7942,N_6697,N_6678);
or U7943 (N_7943,N_6432,N_7170);
nor U7944 (N_7944,N_7123,N_6754);
and U7945 (N_7945,N_6953,N_6658);
or U7946 (N_7946,N_6745,N_7006);
and U7947 (N_7947,N_7051,N_6847);
or U7948 (N_7948,N_7195,N_6640);
or U7949 (N_7949,N_7105,N_7152);
nor U7950 (N_7950,N_6696,N_7150);
nor U7951 (N_7951,N_6438,N_6632);
nand U7952 (N_7952,N_6811,N_6467);
nand U7953 (N_7953,N_6725,N_6634);
nor U7954 (N_7954,N_6863,N_6907);
or U7955 (N_7955,N_6807,N_6529);
and U7956 (N_7956,N_7195,N_7164);
and U7957 (N_7957,N_7156,N_6421);
nor U7958 (N_7958,N_7094,N_6727);
nor U7959 (N_7959,N_6949,N_6855);
xor U7960 (N_7960,N_6946,N_6444);
and U7961 (N_7961,N_7110,N_6690);
and U7962 (N_7962,N_6415,N_6606);
xnor U7963 (N_7963,N_6781,N_7022);
xor U7964 (N_7964,N_6923,N_7009);
xor U7965 (N_7965,N_6683,N_6514);
nor U7966 (N_7966,N_6561,N_6651);
and U7967 (N_7967,N_6698,N_6500);
or U7968 (N_7968,N_6520,N_6858);
nand U7969 (N_7969,N_6921,N_6470);
nor U7970 (N_7970,N_7089,N_6916);
nand U7971 (N_7971,N_6687,N_6749);
or U7972 (N_7972,N_6990,N_6792);
nand U7973 (N_7973,N_6750,N_6597);
nor U7974 (N_7974,N_7038,N_6646);
nor U7975 (N_7975,N_7099,N_7196);
xor U7976 (N_7976,N_6823,N_6762);
nand U7977 (N_7977,N_6484,N_6753);
nand U7978 (N_7978,N_6505,N_6585);
or U7979 (N_7979,N_7032,N_6654);
or U7980 (N_7980,N_6904,N_6551);
or U7981 (N_7981,N_6588,N_6612);
or U7982 (N_7982,N_6457,N_7197);
xnor U7983 (N_7983,N_6745,N_6786);
or U7984 (N_7984,N_6809,N_6418);
xnor U7985 (N_7985,N_6961,N_7066);
nand U7986 (N_7986,N_6738,N_6487);
or U7987 (N_7987,N_6620,N_6918);
nor U7988 (N_7988,N_7001,N_6805);
and U7989 (N_7989,N_6503,N_6950);
nor U7990 (N_7990,N_6811,N_6614);
nand U7991 (N_7991,N_6770,N_6500);
and U7992 (N_7992,N_7043,N_6943);
or U7993 (N_7993,N_7141,N_6912);
and U7994 (N_7994,N_6616,N_6605);
and U7995 (N_7995,N_6695,N_7089);
nor U7996 (N_7996,N_6551,N_6957);
nand U7997 (N_7997,N_6409,N_6534);
or U7998 (N_7998,N_7122,N_6765);
nand U7999 (N_7999,N_6962,N_7014);
nor U8000 (N_8000,N_7570,N_7720);
or U8001 (N_8001,N_7567,N_7363);
and U8002 (N_8002,N_7263,N_7943);
nand U8003 (N_8003,N_7215,N_7712);
and U8004 (N_8004,N_7826,N_7994);
xor U8005 (N_8005,N_7805,N_7484);
or U8006 (N_8006,N_7476,N_7339);
and U8007 (N_8007,N_7629,N_7514);
and U8008 (N_8008,N_7691,N_7600);
or U8009 (N_8009,N_7392,N_7391);
xnor U8010 (N_8010,N_7859,N_7465);
nand U8011 (N_8011,N_7858,N_7912);
xnor U8012 (N_8012,N_7808,N_7979);
xnor U8013 (N_8013,N_7445,N_7644);
nor U8014 (N_8014,N_7539,N_7690);
xor U8015 (N_8015,N_7839,N_7245);
or U8016 (N_8016,N_7229,N_7309);
xor U8017 (N_8017,N_7848,N_7298);
or U8018 (N_8018,N_7780,N_7918);
and U8019 (N_8019,N_7710,N_7524);
nor U8020 (N_8020,N_7910,N_7823);
nand U8021 (N_8021,N_7872,N_7250);
nor U8022 (N_8022,N_7834,N_7645);
nor U8023 (N_8023,N_7835,N_7988);
nand U8024 (N_8024,N_7334,N_7380);
nand U8025 (N_8025,N_7275,N_7743);
and U8026 (N_8026,N_7452,N_7674);
nor U8027 (N_8027,N_7734,N_7421);
nand U8028 (N_8028,N_7490,N_7474);
nand U8029 (N_8029,N_7828,N_7443);
and U8030 (N_8030,N_7272,N_7804);
and U8031 (N_8031,N_7602,N_7781);
nand U8032 (N_8032,N_7766,N_7967);
or U8033 (N_8033,N_7756,N_7706);
nand U8034 (N_8034,N_7417,N_7509);
or U8035 (N_8035,N_7537,N_7891);
xnor U8036 (N_8036,N_7702,N_7547);
xor U8037 (N_8037,N_7248,N_7396);
nand U8038 (N_8038,N_7696,N_7323);
and U8039 (N_8039,N_7224,N_7341);
and U8040 (N_8040,N_7221,N_7719);
xnor U8041 (N_8041,N_7282,N_7990);
xnor U8042 (N_8042,N_7599,N_7900);
nand U8043 (N_8043,N_7862,N_7888);
or U8044 (N_8044,N_7981,N_7203);
and U8045 (N_8045,N_7538,N_7966);
nor U8046 (N_8046,N_7387,N_7803);
or U8047 (N_8047,N_7882,N_7761);
and U8048 (N_8048,N_7786,N_7467);
xor U8049 (N_8049,N_7436,N_7242);
and U8050 (N_8050,N_7253,N_7646);
and U8051 (N_8051,N_7856,N_7814);
and U8052 (N_8052,N_7578,N_7843);
nor U8053 (N_8053,N_7614,N_7752);
nor U8054 (N_8054,N_7950,N_7665);
nor U8055 (N_8055,N_7532,N_7420);
xor U8056 (N_8056,N_7873,N_7505);
nor U8057 (N_8057,N_7362,N_7206);
xnor U8058 (N_8058,N_7493,N_7638);
and U8059 (N_8059,N_7640,N_7573);
nor U8060 (N_8060,N_7300,N_7962);
and U8061 (N_8061,N_7672,N_7355);
and U8062 (N_8062,N_7760,N_7475);
xnor U8063 (N_8063,N_7940,N_7757);
or U8064 (N_8064,N_7968,N_7543);
and U8065 (N_8065,N_7358,N_7499);
nor U8066 (N_8066,N_7855,N_7575);
or U8067 (N_8067,N_7878,N_7703);
nand U8068 (N_8068,N_7213,N_7963);
or U8069 (N_8069,N_7864,N_7208);
or U8070 (N_8070,N_7549,N_7502);
and U8071 (N_8071,N_7222,N_7899);
and U8072 (N_8072,N_7486,N_7378);
nand U8073 (N_8073,N_7832,N_7607);
or U8074 (N_8074,N_7931,N_7916);
xnor U8075 (N_8075,N_7764,N_7303);
or U8076 (N_8076,N_7792,N_7442);
and U8077 (N_8077,N_7955,N_7753);
and U8078 (N_8078,N_7620,N_7960);
xnor U8079 (N_8079,N_7218,N_7866);
and U8080 (N_8080,N_7301,N_7431);
xnor U8081 (N_8081,N_7359,N_7525);
nor U8082 (N_8082,N_7483,N_7914);
xor U8083 (N_8083,N_7513,N_7410);
and U8084 (N_8084,N_7244,N_7553);
and U8085 (N_8085,N_7928,N_7830);
or U8086 (N_8086,N_7783,N_7446);
nor U8087 (N_8087,N_7850,N_7729);
and U8088 (N_8088,N_7572,N_7209);
xnor U8089 (N_8089,N_7657,N_7906);
nor U8090 (N_8090,N_7508,N_7863);
or U8091 (N_8091,N_7820,N_7360);
xor U8092 (N_8092,N_7975,N_7308);
xor U8093 (N_8093,N_7874,N_7790);
or U8094 (N_8094,N_7273,N_7438);
nand U8095 (N_8095,N_7728,N_7892);
nand U8096 (N_8096,N_7297,N_7205);
and U8097 (N_8097,N_7302,N_7586);
and U8098 (N_8098,N_7503,N_7875);
xnor U8099 (N_8099,N_7938,N_7982);
nor U8100 (N_8100,N_7930,N_7909);
nor U8101 (N_8101,N_7664,N_7535);
nand U8102 (N_8102,N_7615,N_7220);
xnor U8103 (N_8103,N_7274,N_7344);
and U8104 (N_8104,N_7214,N_7330);
xnor U8105 (N_8105,N_7207,N_7371);
or U8106 (N_8106,N_7526,N_7773);
nor U8107 (N_8107,N_7501,N_7447);
nand U8108 (N_8108,N_7470,N_7292);
or U8109 (N_8109,N_7342,N_7777);
or U8110 (N_8110,N_7400,N_7705);
nand U8111 (N_8111,N_7802,N_7590);
xor U8112 (N_8112,N_7239,N_7592);
xor U8113 (N_8113,N_7317,N_7627);
xnor U8114 (N_8114,N_7472,N_7851);
and U8115 (N_8115,N_7243,N_7867);
nand U8116 (N_8116,N_7240,N_7279);
nor U8117 (N_8117,N_7701,N_7451);
or U8118 (N_8118,N_7349,N_7887);
and U8119 (N_8119,N_7869,N_7755);
and U8120 (N_8120,N_7210,N_7681);
nand U8121 (N_8121,N_7903,N_7458);
and U8122 (N_8122,N_7427,N_7929);
nor U8123 (N_8123,N_7852,N_7669);
nor U8124 (N_8124,N_7958,N_7594);
and U8125 (N_8125,N_7405,N_7890);
and U8126 (N_8126,N_7973,N_7384);
xnor U8127 (N_8127,N_7609,N_7544);
and U8128 (N_8128,N_7601,N_7324);
or U8129 (N_8129,N_7817,N_7422);
and U8130 (N_8130,N_7404,N_7934);
nand U8131 (N_8131,N_7683,N_7949);
nor U8132 (N_8132,N_7985,N_7225);
and U8133 (N_8133,N_7256,N_7932);
and U8134 (N_8134,N_7348,N_7726);
and U8135 (N_8135,N_7551,N_7722);
or U8136 (N_8136,N_7688,N_7398);
or U8137 (N_8137,N_7978,N_7550);
nand U8138 (N_8138,N_7546,N_7795);
nand U8139 (N_8139,N_7260,N_7618);
nor U8140 (N_8140,N_7937,N_7321);
or U8141 (N_8141,N_7810,N_7738);
xnor U8142 (N_8142,N_7419,N_7401);
nor U8143 (N_8143,N_7639,N_7763);
and U8144 (N_8144,N_7905,N_7412);
or U8145 (N_8145,N_7876,N_7587);
nand U8146 (N_8146,N_7226,N_7388);
and U8147 (N_8147,N_7845,N_7316);
and U8148 (N_8148,N_7351,N_7495);
or U8149 (N_8149,N_7313,N_7336);
nand U8150 (N_8150,N_7374,N_7418);
and U8151 (N_8151,N_7232,N_7439);
xnor U8152 (N_8152,N_7255,N_7736);
xor U8153 (N_8153,N_7557,N_7343);
xnor U8154 (N_8154,N_7633,N_7758);
xnor U8155 (N_8155,N_7998,N_7361);
nor U8156 (N_8156,N_7796,N_7558);
xnor U8157 (N_8157,N_7379,N_7643);
xnor U8158 (N_8158,N_7516,N_7849);
xor U8159 (N_8159,N_7699,N_7816);
xnor U8160 (N_8160,N_7376,N_7481);
xor U8161 (N_8161,N_7831,N_7449);
xnor U8162 (N_8162,N_7861,N_7574);
xor U8163 (N_8163,N_7842,N_7434);
nand U8164 (N_8164,N_7327,N_7433);
nand U8165 (N_8165,N_7373,N_7312);
and U8166 (N_8166,N_7662,N_7364);
or U8167 (N_8167,N_7715,N_7995);
xnor U8168 (N_8168,N_7304,N_7671);
or U8169 (N_8169,N_7993,N_7367);
and U8170 (N_8170,N_7577,N_7881);
nand U8171 (N_8171,N_7735,N_7907);
nor U8172 (N_8172,N_7588,N_7389);
nand U8173 (N_8173,N_7377,N_7860);
xor U8174 (N_8174,N_7991,N_7320);
xnor U8175 (N_8175,N_7247,N_7844);
or U8176 (N_8176,N_7723,N_7926);
or U8177 (N_8177,N_7840,N_7237);
nand U8178 (N_8178,N_7879,N_7459);
xor U8179 (N_8179,N_7822,N_7576);
nor U8180 (N_8180,N_7653,N_7463);
nor U8181 (N_8181,N_7782,N_7714);
xnor U8182 (N_8182,N_7406,N_7612);
xnor U8183 (N_8183,N_7440,N_7295);
nand U8184 (N_8184,N_7216,N_7437);
and U8185 (N_8185,N_7285,N_7326);
or U8186 (N_8186,N_7785,N_7515);
xor U8187 (N_8187,N_7896,N_7281);
xnor U8188 (N_8188,N_7754,N_7700);
nand U8189 (N_8189,N_7821,N_7211);
xor U8190 (N_8190,N_7774,N_7315);
nand U8191 (N_8191,N_7969,N_7429);
or U8192 (N_8192,N_7893,N_7280);
nor U8193 (N_8193,N_7485,N_7689);
nor U8194 (N_8194,N_7885,N_7491);
and U8195 (N_8195,N_7732,N_7825);
or U8196 (N_8196,N_7976,N_7622);
nor U8197 (N_8197,N_7325,N_7291);
xor U8198 (N_8198,N_7267,N_7654);
xor U8199 (N_8199,N_7530,N_7913);
nor U8200 (N_8200,N_7236,N_7692);
nor U8201 (N_8201,N_7974,N_7686);
nor U8202 (N_8202,N_7789,N_7517);
xnor U8203 (N_8203,N_7667,N_7673);
nand U8204 (N_8204,N_7277,N_7799);
nand U8205 (N_8205,N_7895,N_7563);
and U8206 (N_8206,N_7897,N_7269);
xnor U8207 (N_8207,N_7270,N_7693);
nand U8208 (N_8208,N_7911,N_7556);
nor U8209 (N_8209,N_7959,N_7886);
or U8210 (N_8210,N_7961,N_7871);
nor U8211 (N_8211,N_7286,N_7504);
nand U8212 (N_8212,N_7923,N_7322);
nor U8213 (N_8213,N_7454,N_7806);
nand U8214 (N_8214,N_7682,N_7748);
nor U8215 (N_8215,N_7611,N_7775);
nand U8216 (N_8216,N_7964,N_7647);
nor U8217 (N_8217,N_7372,N_7679);
and U8218 (N_8218,N_7428,N_7857);
nor U8219 (N_8219,N_7770,N_7718);
or U8220 (N_8220,N_7477,N_7744);
nor U8221 (N_8221,N_7251,N_7917);
or U8222 (N_8222,N_7534,N_7684);
or U8223 (N_8223,N_7507,N_7984);
and U8224 (N_8224,N_7740,N_7791);
and U8225 (N_8225,N_7290,N_7571);
and U8226 (N_8226,N_7939,N_7957);
or U8227 (N_8227,N_7545,N_7725);
nand U8228 (N_8228,N_7582,N_7980);
nor U8229 (N_8229,N_7779,N_7731);
nor U8230 (N_8230,N_7531,N_7564);
nand U8231 (N_8231,N_7658,N_7709);
or U8232 (N_8232,N_7983,N_7500);
xnor U8233 (N_8233,N_7569,N_7271);
or U8234 (N_8234,N_7711,N_7390);
or U8235 (N_8235,N_7494,N_7407);
nand U8236 (N_8236,N_7807,N_7289);
nor U8237 (N_8237,N_7261,N_7276);
and U8238 (N_8238,N_7730,N_7347);
or U8239 (N_8239,N_7996,N_7769);
nor U8240 (N_8240,N_7987,N_7265);
nor U8241 (N_8241,N_7337,N_7695);
or U8242 (N_8242,N_7927,N_7596);
xor U8243 (N_8243,N_7765,N_7293);
and U8244 (N_8244,N_7908,N_7555);
nor U8245 (N_8245,N_7787,N_7812);
and U8246 (N_8246,N_7331,N_7241);
nor U8247 (N_8247,N_7299,N_7945);
or U8248 (N_8248,N_7552,N_7462);
and U8249 (N_8249,N_7656,N_7307);
and U8250 (N_8250,N_7217,N_7680);
or U8251 (N_8251,N_7922,N_7579);
or U8252 (N_8252,N_7212,N_7370);
nor U8253 (N_8253,N_7473,N_7837);
nor U8254 (N_8254,N_7489,N_7335);
nor U8255 (N_8255,N_7455,N_7416);
nor U8256 (N_8256,N_7668,N_7708);
xnor U8257 (N_8257,N_7933,N_7511);
nand U8258 (N_8258,N_7258,N_7262);
and U8259 (N_8259,N_7227,N_7395);
nand U8260 (N_8260,N_7641,N_7617);
and U8261 (N_8261,N_7512,N_7460);
or U8262 (N_8262,N_7562,N_7580);
and U8263 (N_8263,N_7448,N_7631);
xnor U8264 (N_8264,N_7951,N_7624);
nor U8265 (N_8265,N_7464,N_7287);
and U8266 (N_8266,N_7642,N_7368);
and U8267 (N_8267,N_7619,N_7952);
or U8268 (N_8268,N_7529,N_7478);
and U8269 (N_8269,N_7687,N_7915);
nand U8270 (N_8270,N_7737,N_7997);
nand U8271 (N_8271,N_7651,N_7589);
xnor U8272 (N_8272,N_7824,N_7383);
and U8273 (N_8273,N_7435,N_7784);
xnor U8274 (N_8274,N_7597,N_7751);
or U8275 (N_8275,N_7759,N_7884);
and U8276 (N_8276,N_7605,N_7266);
nand U8277 (N_8277,N_7898,N_7257);
nand U8278 (N_8278,N_7528,N_7847);
or U8279 (N_8279,N_7634,N_7698);
nand U8280 (N_8280,N_7880,N_7519);
xor U8281 (N_8281,N_7801,N_7479);
and U8282 (N_8282,N_7883,N_7408);
and U8283 (N_8283,N_7469,N_7548);
or U8284 (N_8284,N_7284,N_7739);
nor U8285 (N_8285,N_7946,N_7685);
xnor U8286 (N_8286,N_7632,N_7369);
and U8287 (N_8287,N_7527,N_7354);
or U8288 (N_8288,N_7352,N_7249);
nor U8289 (N_8289,N_7310,N_7800);
nor U8290 (N_8290,N_7231,N_7965);
xor U8291 (N_8291,N_7393,N_7319);
and U8292 (N_8292,N_7561,N_7670);
nor U8293 (N_8293,N_7935,N_7523);
and U8294 (N_8294,N_7818,N_7704);
and U8295 (N_8295,N_7595,N_7397);
xor U8296 (N_8296,N_7432,N_7724);
xnor U8297 (N_8297,N_7846,N_7584);
nor U8298 (N_8298,N_7877,N_7450);
nand U8299 (N_8299,N_7953,N_7676);
nand U8300 (N_8300,N_7403,N_7733);
nor U8301 (N_8301,N_7252,N_7510);
or U8302 (N_8302,N_7836,N_7468);
nand U8303 (N_8303,N_7471,N_7741);
nand U8304 (N_8304,N_7466,N_7697);
nor U8305 (N_8305,N_7901,N_7677);
xor U8306 (N_8306,N_7498,N_7956);
nor U8307 (N_8307,N_7585,N_7488);
or U8308 (N_8308,N_7659,N_7727);
and U8309 (N_8309,N_7296,N_7794);
nand U8310 (N_8310,N_7660,N_7970);
nand U8311 (N_8311,N_7655,N_7314);
or U8312 (N_8312,N_7793,N_7332);
and U8313 (N_8313,N_7542,N_7350);
xnor U8314 (N_8314,N_7920,N_7560);
or U8315 (N_8315,N_7235,N_7385);
xor U8316 (N_8316,N_7649,N_7536);
nor U8317 (N_8317,N_7202,N_7414);
or U8318 (N_8318,N_7999,N_7533);
xnor U8319 (N_8319,N_7598,N_7283);
nand U8320 (N_8320,N_7233,N_7487);
nand U8321 (N_8321,N_7441,N_7853);
xnor U8322 (N_8322,N_7278,N_7568);
nor U8323 (N_8323,N_7833,N_7566);
nor U8324 (N_8324,N_7716,N_7650);
nor U8325 (N_8325,N_7621,N_7746);
nand U8326 (N_8326,N_7254,N_7626);
or U8327 (N_8327,N_7411,N_7606);
and U8328 (N_8328,N_7306,N_7522);
or U8329 (N_8329,N_7925,N_7457);
or U8330 (N_8330,N_7986,N_7461);
or U8331 (N_8331,N_7838,N_7591);
or U8332 (N_8332,N_7675,N_7413);
or U8333 (N_8333,N_7815,N_7889);
xnor U8334 (N_8334,N_7456,N_7771);
nand U8335 (N_8335,N_7305,N_7201);
nand U8336 (N_8336,N_7430,N_7954);
nand U8337 (N_8337,N_7204,N_7246);
nor U8338 (N_8338,N_7409,N_7496);
and U8339 (N_8339,N_7294,N_7497);
and U8340 (N_8340,N_7772,N_7424);
nor U8341 (N_8341,N_7581,N_7423);
and U8342 (N_8342,N_7717,N_7394);
nor U8343 (N_8343,N_7989,N_7329);
nand U8344 (N_8344,N_7230,N_7750);
xor U8345 (N_8345,N_7798,N_7648);
xnor U8346 (N_8346,N_7921,N_7333);
xor U8347 (N_8347,N_7778,N_7623);
nor U8348 (N_8348,N_7540,N_7868);
and U8349 (N_8349,N_7238,N_7870);
xnor U8350 (N_8350,N_7415,N_7345);
nor U8351 (N_8351,N_7357,N_7661);
nand U8352 (N_8352,N_7768,N_7616);
nand U8353 (N_8353,N_7541,N_7865);
xor U8354 (N_8354,N_7608,N_7328);
nand U8355 (N_8355,N_7767,N_7259);
xor U8356 (N_8356,N_7375,N_7904);
nor U8357 (N_8357,N_7268,N_7318);
xnor U8358 (N_8358,N_7636,N_7813);
or U8359 (N_8359,N_7749,N_7338);
and U8360 (N_8360,N_7223,N_7554);
or U8361 (N_8361,N_7776,N_7353);
nand U8362 (N_8362,N_7694,N_7971);
or U8363 (N_8363,N_7811,N_7944);
or U8364 (N_8364,N_7809,N_7628);
or U8365 (N_8365,N_7604,N_7745);
nand U8366 (N_8366,N_7948,N_7399);
nand U8367 (N_8367,N_7506,N_7635);
or U8368 (N_8368,N_7829,N_7402);
and U8369 (N_8369,N_7707,N_7841);
nor U8370 (N_8370,N_7747,N_7482);
or U8371 (N_8371,N_7518,N_7365);
nor U8372 (N_8372,N_7678,N_7721);
and U8373 (N_8373,N_7492,N_7827);
nand U8374 (N_8374,N_7894,N_7713);
xor U8375 (N_8375,N_7788,N_7311);
and U8376 (N_8376,N_7666,N_7425);
or U8377 (N_8377,N_7386,N_7652);
and U8378 (N_8378,N_7453,N_7797);
or U8379 (N_8379,N_7854,N_7480);
or U8380 (N_8380,N_7381,N_7288);
or U8381 (N_8381,N_7992,N_7941);
nor U8382 (N_8382,N_7762,N_7625);
and U8383 (N_8383,N_7637,N_7234);
xnor U8384 (N_8384,N_7346,N_7593);
and U8385 (N_8385,N_7356,N_7924);
xnor U8386 (N_8386,N_7919,N_7613);
or U8387 (N_8387,N_7366,N_7630);
or U8388 (N_8388,N_7819,N_7977);
or U8389 (N_8389,N_7565,N_7228);
nor U8390 (N_8390,N_7583,N_7520);
nor U8391 (N_8391,N_7444,N_7340);
xor U8392 (N_8392,N_7610,N_7559);
xnor U8393 (N_8393,N_7947,N_7200);
nand U8394 (N_8394,N_7219,N_7972);
nor U8395 (N_8395,N_7264,N_7521);
or U8396 (N_8396,N_7742,N_7426);
nand U8397 (N_8397,N_7942,N_7603);
nand U8398 (N_8398,N_7663,N_7936);
nand U8399 (N_8399,N_7902,N_7382);
xnor U8400 (N_8400,N_7484,N_7999);
nor U8401 (N_8401,N_7334,N_7577);
xor U8402 (N_8402,N_7422,N_7421);
nor U8403 (N_8403,N_7551,N_7909);
nor U8404 (N_8404,N_7823,N_7507);
nor U8405 (N_8405,N_7876,N_7689);
and U8406 (N_8406,N_7854,N_7399);
or U8407 (N_8407,N_7792,N_7375);
nor U8408 (N_8408,N_7557,N_7526);
or U8409 (N_8409,N_7846,N_7645);
nand U8410 (N_8410,N_7342,N_7875);
nor U8411 (N_8411,N_7413,N_7537);
or U8412 (N_8412,N_7585,N_7471);
or U8413 (N_8413,N_7761,N_7933);
nand U8414 (N_8414,N_7823,N_7623);
nand U8415 (N_8415,N_7417,N_7450);
or U8416 (N_8416,N_7336,N_7510);
and U8417 (N_8417,N_7213,N_7749);
nand U8418 (N_8418,N_7415,N_7818);
nor U8419 (N_8419,N_7846,N_7997);
or U8420 (N_8420,N_7475,N_7541);
and U8421 (N_8421,N_7434,N_7444);
or U8422 (N_8422,N_7253,N_7794);
xor U8423 (N_8423,N_7878,N_7204);
and U8424 (N_8424,N_7932,N_7523);
or U8425 (N_8425,N_7661,N_7768);
and U8426 (N_8426,N_7520,N_7925);
xnor U8427 (N_8427,N_7971,N_7947);
or U8428 (N_8428,N_7730,N_7965);
or U8429 (N_8429,N_7258,N_7370);
xor U8430 (N_8430,N_7762,N_7824);
nor U8431 (N_8431,N_7458,N_7624);
and U8432 (N_8432,N_7773,N_7785);
nor U8433 (N_8433,N_7764,N_7578);
nand U8434 (N_8434,N_7278,N_7776);
xor U8435 (N_8435,N_7669,N_7862);
nor U8436 (N_8436,N_7667,N_7771);
or U8437 (N_8437,N_7853,N_7922);
or U8438 (N_8438,N_7291,N_7835);
or U8439 (N_8439,N_7963,N_7526);
and U8440 (N_8440,N_7525,N_7547);
xor U8441 (N_8441,N_7318,N_7258);
nor U8442 (N_8442,N_7586,N_7256);
and U8443 (N_8443,N_7878,N_7439);
and U8444 (N_8444,N_7322,N_7950);
and U8445 (N_8445,N_7395,N_7350);
nand U8446 (N_8446,N_7870,N_7277);
and U8447 (N_8447,N_7662,N_7621);
and U8448 (N_8448,N_7596,N_7542);
xnor U8449 (N_8449,N_7399,N_7630);
or U8450 (N_8450,N_7816,N_7877);
or U8451 (N_8451,N_7336,N_7923);
nand U8452 (N_8452,N_7426,N_7321);
xor U8453 (N_8453,N_7797,N_7878);
xor U8454 (N_8454,N_7746,N_7260);
nand U8455 (N_8455,N_7236,N_7667);
nand U8456 (N_8456,N_7383,N_7478);
nand U8457 (N_8457,N_7645,N_7252);
nor U8458 (N_8458,N_7338,N_7702);
xor U8459 (N_8459,N_7782,N_7654);
nor U8460 (N_8460,N_7298,N_7571);
and U8461 (N_8461,N_7962,N_7747);
xor U8462 (N_8462,N_7206,N_7541);
or U8463 (N_8463,N_7752,N_7297);
and U8464 (N_8464,N_7781,N_7679);
and U8465 (N_8465,N_7776,N_7753);
nor U8466 (N_8466,N_7263,N_7812);
xor U8467 (N_8467,N_7809,N_7693);
or U8468 (N_8468,N_7840,N_7204);
or U8469 (N_8469,N_7387,N_7832);
or U8470 (N_8470,N_7371,N_7681);
or U8471 (N_8471,N_7805,N_7488);
xnor U8472 (N_8472,N_7720,N_7499);
nand U8473 (N_8473,N_7324,N_7813);
xnor U8474 (N_8474,N_7396,N_7944);
or U8475 (N_8475,N_7434,N_7376);
or U8476 (N_8476,N_7570,N_7564);
xor U8477 (N_8477,N_7401,N_7470);
and U8478 (N_8478,N_7341,N_7861);
and U8479 (N_8479,N_7359,N_7267);
xor U8480 (N_8480,N_7624,N_7328);
or U8481 (N_8481,N_7435,N_7853);
nor U8482 (N_8482,N_7591,N_7819);
and U8483 (N_8483,N_7941,N_7689);
or U8484 (N_8484,N_7513,N_7577);
nand U8485 (N_8485,N_7809,N_7802);
or U8486 (N_8486,N_7242,N_7455);
or U8487 (N_8487,N_7278,N_7560);
nor U8488 (N_8488,N_7247,N_7407);
or U8489 (N_8489,N_7822,N_7996);
and U8490 (N_8490,N_7262,N_7788);
and U8491 (N_8491,N_7415,N_7949);
nand U8492 (N_8492,N_7689,N_7602);
or U8493 (N_8493,N_7980,N_7323);
or U8494 (N_8494,N_7397,N_7810);
and U8495 (N_8495,N_7782,N_7594);
and U8496 (N_8496,N_7239,N_7870);
nand U8497 (N_8497,N_7459,N_7391);
nor U8498 (N_8498,N_7919,N_7847);
and U8499 (N_8499,N_7254,N_7585);
and U8500 (N_8500,N_7600,N_7834);
or U8501 (N_8501,N_7608,N_7864);
nor U8502 (N_8502,N_7822,N_7224);
xnor U8503 (N_8503,N_7315,N_7288);
or U8504 (N_8504,N_7638,N_7318);
and U8505 (N_8505,N_7347,N_7999);
and U8506 (N_8506,N_7968,N_7402);
nor U8507 (N_8507,N_7398,N_7442);
nand U8508 (N_8508,N_7482,N_7276);
nand U8509 (N_8509,N_7237,N_7729);
xor U8510 (N_8510,N_7488,N_7407);
nand U8511 (N_8511,N_7947,N_7372);
nand U8512 (N_8512,N_7533,N_7919);
nand U8513 (N_8513,N_7258,N_7782);
xnor U8514 (N_8514,N_7360,N_7589);
nand U8515 (N_8515,N_7305,N_7420);
nor U8516 (N_8516,N_7659,N_7500);
nor U8517 (N_8517,N_7925,N_7663);
and U8518 (N_8518,N_7633,N_7620);
and U8519 (N_8519,N_7495,N_7901);
or U8520 (N_8520,N_7734,N_7486);
nor U8521 (N_8521,N_7338,N_7786);
xor U8522 (N_8522,N_7672,N_7334);
nor U8523 (N_8523,N_7892,N_7296);
or U8524 (N_8524,N_7488,N_7618);
xor U8525 (N_8525,N_7790,N_7905);
and U8526 (N_8526,N_7393,N_7487);
and U8527 (N_8527,N_7485,N_7824);
nor U8528 (N_8528,N_7326,N_7443);
nor U8529 (N_8529,N_7323,N_7569);
nor U8530 (N_8530,N_7931,N_7961);
and U8531 (N_8531,N_7871,N_7918);
nor U8532 (N_8532,N_7347,N_7444);
xnor U8533 (N_8533,N_7717,N_7656);
and U8534 (N_8534,N_7661,N_7809);
xnor U8535 (N_8535,N_7413,N_7436);
or U8536 (N_8536,N_7509,N_7747);
xnor U8537 (N_8537,N_7645,N_7474);
or U8538 (N_8538,N_7557,N_7614);
or U8539 (N_8539,N_7678,N_7272);
xnor U8540 (N_8540,N_7874,N_7791);
nor U8541 (N_8541,N_7638,N_7700);
or U8542 (N_8542,N_7622,N_7685);
or U8543 (N_8543,N_7562,N_7684);
nor U8544 (N_8544,N_7988,N_7924);
xor U8545 (N_8545,N_7484,N_7688);
xnor U8546 (N_8546,N_7588,N_7294);
and U8547 (N_8547,N_7222,N_7522);
and U8548 (N_8548,N_7431,N_7706);
nor U8549 (N_8549,N_7300,N_7443);
or U8550 (N_8550,N_7295,N_7442);
or U8551 (N_8551,N_7811,N_7545);
nand U8552 (N_8552,N_7726,N_7677);
and U8553 (N_8553,N_7282,N_7842);
nor U8554 (N_8554,N_7244,N_7750);
and U8555 (N_8555,N_7212,N_7699);
nand U8556 (N_8556,N_7950,N_7841);
and U8557 (N_8557,N_7224,N_7236);
nor U8558 (N_8558,N_7975,N_7553);
nand U8559 (N_8559,N_7999,N_7603);
nor U8560 (N_8560,N_7381,N_7733);
nand U8561 (N_8561,N_7395,N_7275);
or U8562 (N_8562,N_7819,N_7409);
xnor U8563 (N_8563,N_7256,N_7909);
or U8564 (N_8564,N_7335,N_7979);
or U8565 (N_8565,N_7263,N_7645);
xor U8566 (N_8566,N_7824,N_7618);
nor U8567 (N_8567,N_7928,N_7505);
xnor U8568 (N_8568,N_7343,N_7312);
nand U8569 (N_8569,N_7205,N_7308);
xnor U8570 (N_8570,N_7951,N_7730);
or U8571 (N_8571,N_7277,N_7639);
and U8572 (N_8572,N_7610,N_7393);
xor U8573 (N_8573,N_7553,N_7974);
nor U8574 (N_8574,N_7961,N_7805);
xnor U8575 (N_8575,N_7796,N_7763);
and U8576 (N_8576,N_7774,N_7484);
and U8577 (N_8577,N_7929,N_7566);
nand U8578 (N_8578,N_7290,N_7669);
or U8579 (N_8579,N_7584,N_7807);
or U8580 (N_8580,N_7364,N_7464);
xor U8581 (N_8581,N_7594,N_7428);
or U8582 (N_8582,N_7834,N_7819);
and U8583 (N_8583,N_7267,N_7329);
nand U8584 (N_8584,N_7201,N_7661);
or U8585 (N_8585,N_7541,N_7498);
nand U8586 (N_8586,N_7959,N_7666);
or U8587 (N_8587,N_7370,N_7596);
nor U8588 (N_8588,N_7739,N_7749);
nand U8589 (N_8589,N_7804,N_7795);
nor U8590 (N_8590,N_7670,N_7899);
xnor U8591 (N_8591,N_7427,N_7673);
xnor U8592 (N_8592,N_7538,N_7375);
and U8593 (N_8593,N_7270,N_7508);
xor U8594 (N_8594,N_7715,N_7860);
nor U8595 (N_8595,N_7256,N_7988);
and U8596 (N_8596,N_7498,N_7876);
nand U8597 (N_8597,N_7865,N_7248);
or U8598 (N_8598,N_7509,N_7916);
or U8599 (N_8599,N_7766,N_7650);
or U8600 (N_8600,N_7913,N_7897);
and U8601 (N_8601,N_7660,N_7828);
xnor U8602 (N_8602,N_7657,N_7805);
nor U8603 (N_8603,N_7424,N_7950);
and U8604 (N_8604,N_7359,N_7762);
xnor U8605 (N_8605,N_7478,N_7999);
nand U8606 (N_8606,N_7621,N_7219);
or U8607 (N_8607,N_7593,N_7700);
or U8608 (N_8608,N_7648,N_7838);
nand U8609 (N_8609,N_7705,N_7203);
nand U8610 (N_8610,N_7568,N_7458);
xnor U8611 (N_8611,N_7871,N_7499);
or U8612 (N_8612,N_7873,N_7513);
or U8613 (N_8613,N_7760,N_7426);
nand U8614 (N_8614,N_7583,N_7712);
and U8615 (N_8615,N_7257,N_7442);
xnor U8616 (N_8616,N_7823,N_7650);
xor U8617 (N_8617,N_7578,N_7888);
and U8618 (N_8618,N_7374,N_7561);
and U8619 (N_8619,N_7304,N_7201);
nor U8620 (N_8620,N_7730,N_7411);
xor U8621 (N_8621,N_7436,N_7679);
nand U8622 (N_8622,N_7771,N_7669);
or U8623 (N_8623,N_7840,N_7517);
and U8624 (N_8624,N_7468,N_7412);
xnor U8625 (N_8625,N_7904,N_7731);
or U8626 (N_8626,N_7925,N_7773);
and U8627 (N_8627,N_7268,N_7467);
and U8628 (N_8628,N_7242,N_7480);
or U8629 (N_8629,N_7837,N_7679);
or U8630 (N_8630,N_7390,N_7700);
and U8631 (N_8631,N_7903,N_7901);
xnor U8632 (N_8632,N_7261,N_7869);
xnor U8633 (N_8633,N_7603,N_7521);
or U8634 (N_8634,N_7725,N_7840);
nand U8635 (N_8635,N_7684,N_7817);
and U8636 (N_8636,N_7706,N_7337);
xor U8637 (N_8637,N_7800,N_7608);
and U8638 (N_8638,N_7758,N_7587);
xnor U8639 (N_8639,N_7873,N_7472);
xor U8640 (N_8640,N_7797,N_7957);
xnor U8641 (N_8641,N_7214,N_7780);
nand U8642 (N_8642,N_7838,N_7317);
nor U8643 (N_8643,N_7657,N_7871);
xor U8644 (N_8644,N_7328,N_7905);
or U8645 (N_8645,N_7890,N_7256);
xnor U8646 (N_8646,N_7221,N_7277);
and U8647 (N_8647,N_7245,N_7541);
or U8648 (N_8648,N_7647,N_7398);
and U8649 (N_8649,N_7590,N_7584);
and U8650 (N_8650,N_7834,N_7991);
nor U8651 (N_8651,N_7868,N_7428);
nand U8652 (N_8652,N_7227,N_7493);
nor U8653 (N_8653,N_7260,N_7602);
nand U8654 (N_8654,N_7420,N_7951);
nand U8655 (N_8655,N_7493,N_7721);
nor U8656 (N_8656,N_7627,N_7475);
and U8657 (N_8657,N_7977,N_7466);
nor U8658 (N_8658,N_7885,N_7825);
xnor U8659 (N_8659,N_7902,N_7633);
or U8660 (N_8660,N_7702,N_7307);
nor U8661 (N_8661,N_7891,N_7814);
or U8662 (N_8662,N_7352,N_7319);
or U8663 (N_8663,N_7640,N_7444);
and U8664 (N_8664,N_7417,N_7277);
and U8665 (N_8665,N_7988,N_7625);
or U8666 (N_8666,N_7606,N_7583);
and U8667 (N_8667,N_7280,N_7674);
and U8668 (N_8668,N_7472,N_7374);
or U8669 (N_8669,N_7961,N_7783);
nand U8670 (N_8670,N_7496,N_7226);
nor U8671 (N_8671,N_7522,N_7483);
xnor U8672 (N_8672,N_7634,N_7958);
xnor U8673 (N_8673,N_7301,N_7753);
xor U8674 (N_8674,N_7921,N_7345);
xnor U8675 (N_8675,N_7416,N_7807);
xor U8676 (N_8676,N_7905,N_7919);
xor U8677 (N_8677,N_7710,N_7511);
or U8678 (N_8678,N_7965,N_7606);
nand U8679 (N_8679,N_7572,N_7897);
nand U8680 (N_8680,N_7573,N_7201);
xnor U8681 (N_8681,N_7936,N_7277);
nor U8682 (N_8682,N_7351,N_7784);
xnor U8683 (N_8683,N_7419,N_7478);
nand U8684 (N_8684,N_7781,N_7556);
and U8685 (N_8685,N_7363,N_7239);
and U8686 (N_8686,N_7398,N_7808);
nor U8687 (N_8687,N_7670,N_7646);
xor U8688 (N_8688,N_7454,N_7396);
nor U8689 (N_8689,N_7966,N_7843);
nand U8690 (N_8690,N_7359,N_7625);
nand U8691 (N_8691,N_7710,N_7316);
and U8692 (N_8692,N_7331,N_7599);
xnor U8693 (N_8693,N_7647,N_7417);
and U8694 (N_8694,N_7982,N_7637);
or U8695 (N_8695,N_7537,N_7288);
xor U8696 (N_8696,N_7382,N_7591);
and U8697 (N_8697,N_7816,N_7567);
and U8698 (N_8698,N_7678,N_7477);
nor U8699 (N_8699,N_7754,N_7655);
or U8700 (N_8700,N_7295,N_7711);
xnor U8701 (N_8701,N_7826,N_7546);
and U8702 (N_8702,N_7844,N_7269);
or U8703 (N_8703,N_7366,N_7567);
nand U8704 (N_8704,N_7665,N_7885);
nor U8705 (N_8705,N_7255,N_7597);
nand U8706 (N_8706,N_7635,N_7913);
or U8707 (N_8707,N_7217,N_7779);
and U8708 (N_8708,N_7517,N_7954);
or U8709 (N_8709,N_7671,N_7628);
nand U8710 (N_8710,N_7948,N_7734);
xor U8711 (N_8711,N_7528,N_7766);
and U8712 (N_8712,N_7817,N_7869);
and U8713 (N_8713,N_7218,N_7917);
nor U8714 (N_8714,N_7635,N_7647);
or U8715 (N_8715,N_7518,N_7805);
xnor U8716 (N_8716,N_7257,N_7532);
or U8717 (N_8717,N_7527,N_7981);
nor U8718 (N_8718,N_7556,N_7376);
nor U8719 (N_8719,N_7993,N_7790);
nor U8720 (N_8720,N_7544,N_7223);
or U8721 (N_8721,N_7708,N_7728);
nand U8722 (N_8722,N_7515,N_7500);
nor U8723 (N_8723,N_7529,N_7455);
nand U8724 (N_8724,N_7880,N_7984);
and U8725 (N_8725,N_7844,N_7481);
or U8726 (N_8726,N_7703,N_7830);
and U8727 (N_8727,N_7902,N_7524);
and U8728 (N_8728,N_7777,N_7352);
nand U8729 (N_8729,N_7431,N_7229);
xnor U8730 (N_8730,N_7411,N_7965);
xnor U8731 (N_8731,N_7658,N_7922);
nand U8732 (N_8732,N_7542,N_7499);
or U8733 (N_8733,N_7252,N_7709);
nor U8734 (N_8734,N_7326,N_7537);
and U8735 (N_8735,N_7983,N_7435);
nor U8736 (N_8736,N_7622,N_7802);
nand U8737 (N_8737,N_7295,N_7604);
xnor U8738 (N_8738,N_7600,N_7959);
and U8739 (N_8739,N_7808,N_7547);
or U8740 (N_8740,N_7792,N_7464);
nor U8741 (N_8741,N_7826,N_7272);
and U8742 (N_8742,N_7437,N_7822);
nand U8743 (N_8743,N_7244,N_7721);
and U8744 (N_8744,N_7315,N_7668);
nand U8745 (N_8745,N_7408,N_7599);
nor U8746 (N_8746,N_7431,N_7436);
xnor U8747 (N_8747,N_7525,N_7201);
nand U8748 (N_8748,N_7971,N_7584);
nand U8749 (N_8749,N_7242,N_7973);
nand U8750 (N_8750,N_7412,N_7728);
and U8751 (N_8751,N_7507,N_7229);
xnor U8752 (N_8752,N_7781,N_7512);
xor U8753 (N_8753,N_7715,N_7250);
and U8754 (N_8754,N_7681,N_7386);
or U8755 (N_8755,N_7549,N_7924);
nand U8756 (N_8756,N_7438,N_7676);
or U8757 (N_8757,N_7678,N_7329);
or U8758 (N_8758,N_7402,N_7622);
xor U8759 (N_8759,N_7404,N_7528);
or U8760 (N_8760,N_7556,N_7245);
and U8761 (N_8761,N_7417,N_7359);
nand U8762 (N_8762,N_7485,N_7272);
and U8763 (N_8763,N_7593,N_7551);
nand U8764 (N_8764,N_7515,N_7725);
xor U8765 (N_8765,N_7628,N_7892);
and U8766 (N_8766,N_7298,N_7348);
nand U8767 (N_8767,N_7462,N_7641);
or U8768 (N_8768,N_7891,N_7999);
xor U8769 (N_8769,N_7529,N_7341);
nor U8770 (N_8770,N_7886,N_7208);
or U8771 (N_8771,N_7278,N_7364);
and U8772 (N_8772,N_7267,N_7347);
xnor U8773 (N_8773,N_7555,N_7711);
or U8774 (N_8774,N_7572,N_7543);
nand U8775 (N_8775,N_7737,N_7642);
xnor U8776 (N_8776,N_7745,N_7712);
or U8777 (N_8777,N_7585,N_7451);
nor U8778 (N_8778,N_7551,N_7790);
and U8779 (N_8779,N_7990,N_7798);
nor U8780 (N_8780,N_7967,N_7444);
or U8781 (N_8781,N_7731,N_7845);
nand U8782 (N_8782,N_7348,N_7225);
or U8783 (N_8783,N_7688,N_7968);
and U8784 (N_8784,N_7595,N_7279);
and U8785 (N_8785,N_7881,N_7727);
or U8786 (N_8786,N_7737,N_7454);
xnor U8787 (N_8787,N_7918,N_7223);
nor U8788 (N_8788,N_7212,N_7235);
xnor U8789 (N_8789,N_7352,N_7628);
or U8790 (N_8790,N_7260,N_7378);
or U8791 (N_8791,N_7410,N_7634);
nand U8792 (N_8792,N_7251,N_7714);
or U8793 (N_8793,N_7907,N_7856);
nor U8794 (N_8794,N_7672,N_7453);
xnor U8795 (N_8795,N_7335,N_7256);
xor U8796 (N_8796,N_7535,N_7379);
nand U8797 (N_8797,N_7334,N_7737);
nand U8798 (N_8798,N_7702,N_7740);
nand U8799 (N_8799,N_7965,N_7490);
and U8800 (N_8800,N_8585,N_8507);
nor U8801 (N_8801,N_8782,N_8593);
or U8802 (N_8802,N_8510,N_8088);
nand U8803 (N_8803,N_8099,N_8634);
or U8804 (N_8804,N_8172,N_8660);
and U8805 (N_8805,N_8423,N_8098);
or U8806 (N_8806,N_8315,N_8466);
nand U8807 (N_8807,N_8054,N_8517);
nand U8808 (N_8808,N_8670,N_8582);
or U8809 (N_8809,N_8415,N_8633);
and U8810 (N_8810,N_8121,N_8064);
xnor U8811 (N_8811,N_8364,N_8650);
nand U8812 (N_8812,N_8482,N_8612);
nand U8813 (N_8813,N_8127,N_8003);
or U8814 (N_8814,N_8201,N_8200);
xor U8815 (N_8815,N_8046,N_8503);
nand U8816 (N_8816,N_8304,N_8717);
and U8817 (N_8817,N_8535,N_8268);
and U8818 (N_8818,N_8070,N_8218);
nand U8819 (N_8819,N_8011,N_8234);
xnor U8820 (N_8820,N_8117,N_8104);
xor U8821 (N_8821,N_8748,N_8513);
xor U8822 (N_8822,N_8402,N_8590);
nor U8823 (N_8823,N_8502,N_8225);
nand U8824 (N_8824,N_8547,N_8756);
xor U8825 (N_8825,N_8635,N_8375);
and U8826 (N_8826,N_8454,N_8282);
nand U8827 (N_8827,N_8223,N_8735);
nor U8828 (N_8828,N_8422,N_8641);
xnor U8829 (N_8829,N_8749,N_8712);
and U8830 (N_8830,N_8493,N_8654);
or U8831 (N_8831,N_8530,N_8055);
and U8832 (N_8832,N_8791,N_8559);
nand U8833 (N_8833,N_8414,N_8467);
xor U8834 (N_8834,N_8214,N_8430);
and U8835 (N_8835,N_8762,N_8529);
or U8836 (N_8836,N_8330,N_8427);
nand U8837 (N_8837,N_8368,N_8401);
and U8838 (N_8838,N_8344,N_8032);
nor U8839 (N_8839,N_8532,N_8085);
and U8840 (N_8840,N_8069,N_8229);
and U8841 (N_8841,N_8653,N_8014);
and U8842 (N_8842,N_8312,N_8391);
and U8843 (N_8843,N_8473,N_8403);
xor U8844 (N_8844,N_8307,N_8698);
or U8845 (N_8845,N_8061,N_8322);
nor U8846 (N_8846,N_8224,N_8656);
nor U8847 (N_8847,N_8460,N_8608);
nor U8848 (N_8848,N_8568,N_8640);
and U8849 (N_8849,N_8595,N_8526);
xor U8850 (N_8850,N_8638,N_8300);
or U8851 (N_8851,N_8065,N_8360);
xnor U8852 (N_8852,N_8584,N_8715);
nand U8853 (N_8853,N_8020,N_8620);
xnor U8854 (N_8854,N_8324,N_8133);
xnor U8855 (N_8855,N_8376,N_8270);
nand U8856 (N_8856,N_8233,N_8692);
xor U8857 (N_8857,N_8116,N_8159);
nor U8858 (N_8858,N_8586,N_8626);
and U8859 (N_8859,N_8577,N_8720);
nor U8860 (N_8860,N_8461,N_8275);
or U8861 (N_8861,N_8523,N_8188);
and U8862 (N_8862,N_8210,N_8134);
nand U8863 (N_8863,N_8674,N_8207);
or U8864 (N_8864,N_8760,N_8484);
nand U8865 (N_8865,N_8082,N_8063);
nand U8866 (N_8866,N_8228,N_8008);
and U8867 (N_8867,N_8028,N_8555);
and U8868 (N_8868,N_8095,N_8714);
nor U8869 (N_8869,N_8034,N_8739);
nor U8870 (N_8870,N_8351,N_8258);
xnor U8871 (N_8871,N_8354,N_8000);
nor U8872 (N_8872,N_8152,N_8107);
nand U8873 (N_8873,N_8349,N_8667);
xor U8874 (N_8874,N_8558,N_8248);
nand U8875 (N_8875,N_8074,N_8156);
or U8876 (N_8876,N_8279,N_8716);
xnor U8877 (N_8877,N_8102,N_8508);
or U8878 (N_8878,N_8338,N_8472);
and U8879 (N_8879,N_8652,N_8792);
nor U8880 (N_8880,N_8266,N_8109);
and U8881 (N_8881,N_8619,N_8398);
and U8882 (N_8882,N_8067,N_8009);
or U8883 (N_8883,N_8628,N_8496);
and U8884 (N_8884,N_8732,N_8179);
nor U8885 (N_8885,N_8004,N_8697);
and U8886 (N_8886,N_8786,N_8591);
xnor U8887 (N_8887,N_8168,N_8309);
xor U8888 (N_8888,N_8500,N_8292);
nor U8889 (N_8889,N_8409,N_8216);
or U8890 (N_8890,N_8777,N_8294);
and U8891 (N_8891,N_8780,N_8658);
and U8892 (N_8892,N_8078,N_8329);
nor U8893 (N_8893,N_8303,N_8580);
nor U8894 (N_8894,N_8611,N_8757);
xnor U8895 (N_8895,N_8736,N_8182);
xor U8896 (N_8896,N_8262,N_8793);
or U8897 (N_8897,N_8221,N_8217);
and U8898 (N_8898,N_8053,N_8776);
and U8899 (N_8899,N_8447,N_8036);
or U8900 (N_8900,N_8389,N_8724);
xor U8901 (N_8901,N_8564,N_8112);
and U8902 (N_8902,N_8546,N_8521);
nor U8903 (N_8903,N_8220,N_8336);
nor U8904 (N_8904,N_8106,N_8280);
nand U8905 (N_8905,N_8655,N_8537);
xnor U8906 (N_8906,N_8105,N_8710);
xor U8907 (N_8907,N_8783,N_8722);
or U8908 (N_8908,N_8689,N_8411);
or U8909 (N_8909,N_8672,N_8741);
nand U8910 (N_8910,N_8742,N_8313);
nand U8911 (N_8911,N_8442,N_8515);
or U8912 (N_8912,N_8249,N_8569);
nor U8913 (N_8913,N_8799,N_8153);
xnor U8914 (N_8914,N_8485,N_8348);
or U8915 (N_8915,N_8150,N_8663);
or U8916 (N_8916,N_8101,N_8281);
nor U8917 (N_8917,N_8708,N_8625);
or U8918 (N_8918,N_8245,N_8729);
nand U8919 (N_8919,N_8754,N_8400);
nand U8920 (N_8920,N_8060,N_8276);
and U8921 (N_8921,N_8199,N_8341);
or U8922 (N_8922,N_8075,N_8788);
and U8923 (N_8923,N_8155,N_8378);
and U8924 (N_8924,N_8058,N_8539);
xnor U8925 (N_8925,N_8534,N_8158);
and U8926 (N_8926,N_8334,N_8594);
nor U8927 (N_8927,N_8267,N_8583);
nand U8928 (N_8928,N_8678,N_8764);
and U8929 (N_8929,N_8092,N_8100);
xor U8930 (N_8930,N_8022,N_8601);
xnor U8931 (N_8931,N_8426,N_8671);
nor U8932 (N_8932,N_8311,N_8452);
and U8933 (N_8933,N_8318,N_8796);
or U8934 (N_8934,N_8683,N_8392);
and U8935 (N_8935,N_8596,N_8607);
nor U8936 (N_8936,N_8433,N_8388);
and U8937 (N_8937,N_8090,N_8421);
xnor U8938 (N_8938,N_8797,N_8752);
and U8939 (N_8939,N_8556,N_8614);
nand U8940 (N_8940,N_8242,N_8328);
and U8941 (N_8941,N_8277,N_8187);
or U8942 (N_8942,N_8299,N_8365);
nor U8943 (N_8943,N_8763,N_8027);
or U8944 (N_8944,N_8616,N_8615);
nand U8945 (N_8945,N_8072,N_8774);
xnor U8946 (N_8946,N_8097,N_8371);
xor U8947 (N_8947,N_8232,N_8361);
nor U8948 (N_8948,N_8527,N_8772);
nand U8949 (N_8949,N_8471,N_8450);
nand U8950 (N_8950,N_8056,N_8035);
or U8951 (N_8951,N_8213,N_8314);
nor U8952 (N_8952,N_8132,N_8769);
xnor U8953 (N_8953,N_8687,N_8044);
and U8954 (N_8954,N_8165,N_8709);
or U8955 (N_8955,N_8321,N_8481);
or U8956 (N_8956,N_8381,N_8491);
or U8957 (N_8957,N_8141,N_8428);
and U8958 (N_8958,N_8093,N_8413);
xnor U8959 (N_8959,N_8033,N_8498);
nand U8960 (N_8960,N_8059,N_8621);
nand U8961 (N_8961,N_8186,N_8347);
and U8962 (N_8962,N_8087,N_8528);
nor U8963 (N_8963,N_8298,N_8146);
xnor U8964 (N_8964,N_8123,N_8045);
xnor U8965 (N_8965,N_8637,N_8778);
and U8966 (N_8966,N_8648,N_8029);
or U8967 (N_8967,N_8369,N_8429);
or U8968 (N_8968,N_8190,N_8699);
and U8969 (N_8969,N_8030,N_8253);
nor U8970 (N_8970,N_8734,N_8352);
nand U8971 (N_8971,N_8366,N_8694);
and U8972 (N_8972,N_8598,N_8779);
and U8973 (N_8973,N_8682,N_8707);
and U8974 (N_8974,N_8103,N_8514);
nor U8975 (N_8975,N_8139,N_8259);
xnor U8976 (N_8976,N_8657,N_8789);
nor U8977 (N_8977,N_8509,N_8420);
xnor U8978 (N_8978,N_8175,N_8629);
xor U8979 (N_8979,N_8219,N_8451);
or U8980 (N_8980,N_8691,N_8609);
and U8981 (N_8981,N_8162,N_8163);
or U8982 (N_8982,N_8557,N_8323);
xor U8983 (N_8983,N_8355,N_8701);
xnor U8984 (N_8984,N_8377,N_8387);
and U8985 (N_8985,N_8549,N_8489);
nand U8986 (N_8986,N_8543,N_8721);
or U8987 (N_8987,N_8140,N_8393);
or U8988 (N_8988,N_8725,N_8448);
nand U8989 (N_8989,N_8096,N_8662);
or U8990 (N_8990,N_8272,N_8646);
and U8991 (N_8991,N_8702,N_8538);
nand U8992 (N_8992,N_8115,N_8531);
nand U8993 (N_8993,N_8181,N_8192);
nor U8994 (N_8994,N_8613,N_8206);
or U8995 (N_8995,N_8755,N_8195);
xor U8996 (N_8996,N_8787,N_8252);
nor U8997 (N_8997,N_8630,N_8157);
xor U8998 (N_8998,N_8129,N_8290);
nand U8999 (N_8999,N_8284,N_8073);
nand U9000 (N_9000,N_8302,N_8773);
nor U9001 (N_9001,N_8205,N_8295);
nor U9002 (N_9002,N_8264,N_8533);
nand U9003 (N_9003,N_8131,N_8340);
xnor U9004 (N_9004,N_8695,N_8790);
nor U9005 (N_9005,N_8647,N_8039);
and U9006 (N_9006,N_8643,N_8463);
and U9007 (N_9007,N_8688,N_8396);
nor U9008 (N_9008,N_8194,N_8296);
nand U9009 (N_9009,N_8669,N_8191);
xor U9010 (N_9010,N_8470,N_8645);
nand U9011 (N_9011,N_8571,N_8048);
nand U9012 (N_9012,N_8209,N_8015);
xnor U9013 (N_9013,N_8052,N_8077);
or U9014 (N_9014,N_8465,N_8287);
nor U9015 (N_9015,N_8337,N_8487);
or U9016 (N_9016,N_8226,N_8359);
and U9017 (N_9017,N_8166,N_8288);
nor U9018 (N_9018,N_8173,N_8738);
and U9019 (N_9019,N_8047,N_8419);
nor U9020 (N_9020,N_8444,N_8468);
and U9021 (N_9021,N_8622,N_8273);
nand U9022 (N_9022,N_8649,N_8703);
or U9023 (N_9023,N_8770,N_8383);
xor U9024 (N_9024,N_8042,N_8222);
and U9025 (N_9025,N_8142,N_8237);
nand U9026 (N_9026,N_8665,N_8386);
nand U9027 (N_9027,N_8407,N_8145);
nand U9028 (N_9028,N_8490,N_8488);
and U9029 (N_9029,N_8746,N_8696);
nand U9030 (N_9030,N_8581,N_8627);
xor U9031 (N_9031,N_8548,N_8504);
nor U9032 (N_9032,N_8236,N_8367);
xor U9033 (N_9033,N_8494,N_8327);
nand U9034 (N_9034,N_8208,N_8379);
nand U9035 (N_9035,N_8164,N_8128);
xor U9036 (N_9036,N_8243,N_8016);
and U9037 (N_9037,N_8363,N_8544);
xor U9038 (N_9038,N_8231,N_8642);
and U9039 (N_9039,N_8565,N_8552);
or U9040 (N_9040,N_8730,N_8184);
xor U9041 (N_9041,N_8317,N_8068);
and U9042 (N_9042,N_8346,N_8540);
and U9043 (N_9043,N_8587,N_8143);
or U9044 (N_9044,N_8562,N_8686);
xnor U9045 (N_9045,N_8438,N_8798);
and U9046 (N_9046,N_8435,N_8519);
and U9047 (N_9047,N_8639,N_8373);
and U9048 (N_9048,N_8137,N_8263);
and U9049 (N_9049,N_8291,N_8301);
nand U9050 (N_9050,N_8592,N_8416);
nor U9051 (N_9051,N_8700,N_8574);
nor U9052 (N_9052,N_8094,N_8525);
xor U9053 (N_9053,N_8486,N_8765);
nand U9054 (N_9054,N_8449,N_8554);
nand U9055 (N_9055,N_8589,N_8561);
xor U9056 (N_9056,N_8006,N_8728);
nand U9057 (N_9057,N_8512,N_8553);
nor U9058 (N_9058,N_8462,N_8197);
xor U9059 (N_9059,N_8439,N_8572);
nor U9060 (N_9060,N_8256,N_8254);
nand U9061 (N_9061,N_8325,N_8759);
and U9062 (N_9062,N_8459,N_8326);
nor U9063 (N_9063,N_8310,N_8124);
nand U9064 (N_9064,N_8305,N_8358);
nor U9065 (N_9065,N_8345,N_8332);
nand U9066 (N_9066,N_8436,N_8605);
or U9067 (N_9067,N_8050,N_8737);
nor U9068 (N_9068,N_8147,N_8417);
nor U9069 (N_9069,N_8474,N_8357);
nor U9070 (N_9070,N_8241,N_8676);
nor U9071 (N_9071,N_8342,N_8478);
nand U9072 (N_9072,N_8251,N_8469);
or U9073 (N_9073,N_8394,N_8684);
or U9074 (N_9074,N_8524,N_8624);
nor U9075 (N_9075,N_8130,N_8110);
and U9076 (N_9076,N_8434,N_8602);
or U9077 (N_9077,N_8768,N_8149);
xnor U9078 (N_9078,N_8545,N_8599);
nor U9079 (N_9079,N_8215,N_8606);
and U9080 (N_9080,N_8541,N_8551);
xnor U9081 (N_9081,N_8505,N_8244);
and U9082 (N_9082,N_8445,N_8084);
or U9083 (N_9083,N_8308,N_8726);
or U9084 (N_9084,N_8536,N_8603);
or U9085 (N_9085,N_8483,N_8285);
xnor U9086 (N_9086,N_8316,N_8271);
nand U9087 (N_9087,N_8125,N_8002);
and U9088 (N_9088,N_8227,N_8293);
and U9089 (N_9089,N_8010,N_8170);
nor U9090 (N_9090,N_8588,N_8644);
and U9091 (N_9091,N_8169,N_8511);
and U9092 (N_9092,N_8183,N_8677);
or U9093 (N_9093,N_8431,N_8176);
nor U9094 (N_9094,N_8516,N_8057);
nand U9095 (N_9095,N_8260,N_8240);
xnor U9096 (N_9096,N_8784,N_8475);
nor U9097 (N_9097,N_8560,N_8563);
nand U9098 (N_9098,N_8743,N_8193);
xor U9099 (N_9099,N_8731,N_8198);
nor U9100 (N_9100,N_8661,N_8753);
xor U9101 (N_9101,N_8230,N_8017);
nand U9102 (N_9102,N_8372,N_8021);
xnor U9103 (N_9103,N_8235,N_8353);
nand U9104 (N_9104,N_8212,N_8119);
nor U9105 (N_9105,N_8719,N_8501);
nand U9106 (N_9106,N_8713,N_8440);
nor U9107 (N_9107,N_8744,N_8204);
nand U9108 (N_9108,N_8480,N_8151);
or U9109 (N_9109,N_8666,N_8781);
and U9110 (N_9110,N_8066,N_8404);
xnor U9111 (N_9111,N_8012,N_8673);
and U9112 (N_9112,N_8664,N_8189);
xnor U9113 (N_9113,N_8455,N_8306);
or U9114 (N_9114,N_8111,N_8617);
nor U9115 (N_9115,N_8005,N_8331);
and U9116 (N_9116,N_8718,N_8750);
and U9117 (N_9117,N_8246,N_8406);
nand U9118 (N_9118,N_8499,N_8446);
and U9119 (N_9119,N_8081,N_8343);
nor U9120 (N_9120,N_8319,N_8086);
xnor U9121 (N_9121,N_8041,N_8618);
or U9122 (N_9122,N_8570,N_8289);
or U9123 (N_9123,N_8453,N_8390);
and U9124 (N_9124,N_8167,N_8136);
nor U9125 (N_9125,N_8610,N_8040);
nor U9126 (N_9126,N_8203,N_8408);
nor U9127 (N_9127,N_8680,N_8771);
nor U9128 (N_9128,N_8578,N_8135);
or U9129 (N_9129,N_8374,N_8178);
xnor U9130 (N_9130,N_8384,N_8575);
nor U9131 (N_9131,N_8395,N_8091);
nand U9132 (N_9132,N_8399,N_8542);
nand U9133 (N_9133,N_8255,N_8250);
nor U9134 (N_9134,N_8679,N_8007);
nand U9135 (N_9135,N_8566,N_8380);
and U9136 (N_9136,N_8118,N_8711);
xnor U9137 (N_9137,N_8579,N_8573);
nor U9138 (N_9138,N_8238,N_8747);
nor U9139 (N_9139,N_8775,N_8693);
or U9140 (N_9140,N_8350,N_8154);
and U9141 (N_9141,N_8794,N_8758);
and U9142 (N_9142,N_8457,N_8623);
or U9143 (N_9143,N_8138,N_8043);
nor U9144 (N_9144,N_8705,N_8604);
nor U9145 (N_9145,N_8297,N_8018);
nor U9146 (N_9146,N_8745,N_8600);
xor U9147 (N_9147,N_8443,N_8382);
nor U9148 (N_9148,N_8479,N_8202);
and U9149 (N_9149,N_8522,N_8019);
nand U9150 (N_9150,N_8492,N_8761);
nand U9151 (N_9151,N_8651,N_8767);
xor U9152 (N_9152,N_8706,N_8432);
and U9153 (N_9153,N_8339,N_8632);
and U9154 (N_9154,N_8013,N_8247);
or U9155 (N_9155,N_8083,N_8257);
or U9156 (N_9156,N_8668,N_8506);
xnor U9157 (N_9157,N_8476,N_8425);
or U9158 (N_9158,N_8286,N_8795);
xnor U9159 (N_9159,N_8122,N_8001);
and U9160 (N_9160,N_8464,N_8727);
nor U9161 (N_9161,N_8196,N_8397);
or U9162 (N_9162,N_8274,N_8024);
xnor U9163 (N_9163,N_8740,N_8089);
xor U9164 (N_9164,N_8320,N_8636);
xnor U9165 (N_9165,N_8239,N_8283);
nand U9166 (N_9166,N_8261,N_8458);
xor U9167 (N_9167,N_8071,N_8180);
or U9168 (N_9168,N_8418,N_8211);
nand U9169 (N_9169,N_8031,N_8265);
or U9170 (N_9170,N_8126,N_8410);
or U9171 (N_9171,N_8079,N_8370);
nand U9172 (N_9172,N_8362,N_8704);
nand U9173 (N_9173,N_8733,N_8076);
nor U9174 (N_9174,N_8062,N_8023);
and U9175 (N_9175,N_8456,N_8690);
nor U9176 (N_9176,N_8025,N_8766);
and U9177 (N_9177,N_8675,N_8497);
nand U9178 (N_9178,N_8038,N_8148);
and U9179 (N_9179,N_8518,N_8049);
xnor U9180 (N_9180,N_8751,N_8477);
or U9181 (N_9181,N_8495,N_8051);
nand U9182 (N_9182,N_8567,N_8185);
nand U9183 (N_9183,N_8171,N_8659);
or U9184 (N_9184,N_8437,N_8597);
and U9185 (N_9185,N_8174,N_8441);
nor U9186 (N_9186,N_8681,N_8405);
or U9187 (N_9187,N_8333,N_8520);
nor U9188 (N_9188,N_8723,N_8080);
nor U9189 (N_9189,N_8269,N_8161);
nor U9190 (N_9190,N_8412,N_8144);
nor U9191 (N_9191,N_8685,N_8631);
and U9192 (N_9192,N_8785,N_8113);
and U9193 (N_9193,N_8177,N_8120);
or U9194 (N_9194,N_8278,N_8037);
xor U9195 (N_9195,N_8108,N_8576);
nand U9196 (N_9196,N_8026,N_8550);
xor U9197 (N_9197,N_8335,N_8424);
xnor U9198 (N_9198,N_8160,N_8385);
nor U9199 (N_9199,N_8114,N_8356);
xnor U9200 (N_9200,N_8059,N_8370);
nand U9201 (N_9201,N_8669,N_8104);
and U9202 (N_9202,N_8087,N_8035);
xnor U9203 (N_9203,N_8735,N_8129);
and U9204 (N_9204,N_8216,N_8020);
xnor U9205 (N_9205,N_8729,N_8044);
and U9206 (N_9206,N_8552,N_8660);
and U9207 (N_9207,N_8312,N_8621);
and U9208 (N_9208,N_8491,N_8757);
or U9209 (N_9209,N_8775,N_8143);
and U9210 (N_9210,N_8064,N_8003);
and U9211 (N_9211,N_8681,N_8049);
xor U9212 (N_9212,N_8553,N_8283);
nand U9213 (N_9213,N_8557,N_8766);
nand U9214 (N_9214,N_8536,N_8729);
or U9215 (N_9215,N_8157,N_8697);
and U9216 (N_9216,N_8791,N_8029);
xnor U9217 (N_9217,N_8257,N_8421);
or U9218 (N_9218,N_8496,N_8230);
xnor U9219 (N_9219,N_8655,N_8153);
and U9220 (N_9220,N_8595,N_8048);
nand U9221 (N_9221,N_8325,N_8714);
nor U9222 (N_9222,N_8563,N_8785);
nor U9223 (N_9223,N_8150,N_8337);
nand U9224 (N_9224,N_8012,N_8406);
nor U9225 (N_9225,N_8030,N_8231);
and U9226 (N_9226,N_8595,N_8777);
and U9227 (N_9227,N_8268,N_8418);
or U9228 (N_9228,N_8004,N_8713);
nand U9229 (N_9229,N_8174,N_8493);
xor U9230 (N_9230,N_8000,N_8165);
nand U9231 (N_9231,N_8282,N_8554);
xnor U9232 (N_9232,N_8425,N_8614);
or U9233 (N_9233,N_8430,N_8024);
nand U9234 (N_9234,N_8063,N_8021);
and U9235 (N_9235,N_8023,N_8076);
nor U9236 (N_9236,N_8300,N_8756);
or U9237 (N_9237,N_8594,N_8672);
xor U9238 (N_9238,N_8372,N_8499);
nor U9239 (N_9239,N_8252,N_8025);
and U9240 (N_9240,N_8774,N_8277);
nor U9241 (N_9241,N_8508,N_8234);
xor U9242 (N_9242,N_8768,N_8232);
nor U9243 (N_9243,N_8726,N_8457);
xnor U9244 (N_9244,N_8358,N_8720);
or U9245 (N_9245,N_8470,N_8514);
nor U9246 (N_9246,N_8083,N_8423);
xnor U9247 (N_9247,N_8057,N_8654);
or U9248 (N_9248,N_8641,N_8775);
nor U9249 (N_9249,N_8207,N_8574);
xnor U9250 (N_9250,N_8745,N_8474);
and U9251 (N_9251,N_8626,N_8301);
and U9252 (N_9252,N_8000,N_8460);
and U9253 (N_9253,N_8602,N_8498);
and U9254 (N_9254,N_8590,N_8592);
nand U9255 (N_9255,N_8287,N_8293);
nor U9256 (N_9256,N_8067,N_8611);
and U9257 (N_9257,N_8260,N_8058);
nor U9258 (N_9258,N_8225,N_8388);
nor U9259 (N_9259,N_8694,N_8126);
or U9260 (N_9260,N_8212,N_8189);
xnor U9261 (N_9261,N_8032,N_8695);
nand U9262 (N_9262,N_8618,N_8250);
and U9263 (N_9263,N_8421,N_8193);
and U9264 (N_9264,N_8723,N_8107);
or U9265 (N_9265,N_8267,N_8286);
nand U9266 (N_9266,N_8019,N_8301);
nand U9267 (N_9267,N_8402,N_8510);
nand U9268 (N_9268,N_8758,N_8628);
xnor U9269 (N_9269,N_8139,N_8571);
xor U9270 (N_9270,N_8778,N_8414);
nand U9271 (N_9271,N_8345,N_8787);
nor U9272 (N_9272,N_8595,N_8384);
xnor U9273 (N_9273,N_8629,N_8222);
nor U9274 (N_9274,N_8147,N_8656);
or U9275 (N_9275,N_8385,N_8202);
nand U9276 (N_9276,N_8106,N_8161);
and U9277 (N_9277,N_8394,N_8636);
and U9278 (N_9278,N_8386,N_8709);
nor U9279 (N_9279,N_8261,N_8009);
or U9280 (N_9280,N_8590,N_8770);
nor U9281 (N_9281,N_8521,N_8645);
nor U9282 (N_9282,N_8348,N_8730);
nand U9283 (N_9283,N_8420,N_8584);
or U9284 (N_9284,N_8479,N_8779);
nand U9285 (N_9285,N_8481,N_8437);
xnor U9286 (N_9286,N_8119,N_8572);
nor U9287 (N_9287,N_8173,N_8186);
and U9288 (N_9288,N_8660,N_8726);
nor U9289 (N_9289,N_8588,N_8245);
and U9290 (N_9290,N_8452,N_8013);
and U9291 (N_9291,N_8093,N_8403);
and U9292 (N_9292,N_8201,N_8467);
xnor U9293 (N_9293,N_8445,N_8576);
nand U9294 (N_9294,N_8593,N_8019);
nand U9295 (N_9295,N_8679,N_8048);
xor U9296 (N_9296,N_8620,N_8666);
nor U9297 (N_9297,N_8785,N_8200);
nor U9298 (N_9298,N_8245,N_8404);
nand U9299 (N_9299,N_8196,N_8136);
and U9300 (N_9300,N_8010,N_8230);
or U9301 (N_9301,N_8127,N_8408);
or U9302 (N_9302,N_8390,N_8582);
or U9303 (N_9303,N_8038,N_8537);
nor U9304 (N_9304,N_8368,N_8298);
and U9305 (N_9305,N_8206,N_8211);
nand U9306 (N_9306,N_8622,N_8781);
nand U9307 (N_9307,N_8461,N_8459);
or U9308 (N_9308,N_8652,N_8155);
xor U9309 (N_9309,N_8405,N_8673);
nand U9310 (N_9310,N_8317,N_8666);
xnor U9311 (N_9311,N_8167,N_8581);
nand U9312 (N_9312,N_8575,N_8686);
nand U9313 (N_9313,N_8740,N_8252);
xnor U9314 (N_9314,N_8305,N_8457);
xnor U9315 (N_9315,N_8646,N_8209);
and U9316 (N_9316,N_8054,N_8698);
nor U9317 (N_9317,N_8321,N_8365);
xor U9318 (N_9318,N_8145,N_8731);
nand U9319 (N_9319,N_8198,N_8469);
and U9320 (N_9320,N_8309,N_8055);
nand U9321 (N_9321,N_8278,N_8606);
and U9322 (N_9322,N_8156,N_8216);
or U9323 (N_9323,N_8773,N_8473);
and U9324 (N_9324,N_8126,N_8365);
and U9325 (N_9325,N_8417,N_8547);
and U9326 (N_9326,N_8517,N_8327);
nand U9327 (N_9327,N_8208,N_8083);
and U9328 (N_9328,N_8382,N_8148);
nand U9329 (N_9329,N_8602,N_8422);
nand U9330 (N_9330,N_8764,N_8372);
nor U9331 (N_9331,N_8019,N_8531);
nand U9332 (N_9332,N_8336,N_8754);
nor U9333 (N_9333,N_8542,N_8675);
nor U9334 (N_9334,N_8423,N_8353);
xor U9335 (N_9335,N_8383,N_8681);
nand U9336 (N_9336,N_8111,N_8258);
or U9337 (N_9337,N_8414,N_8574);
nor U9338 (N_9338,N_8547,N_8257);
or U9339 (N_9339,N_8465,N_8299);
or U9340 (N_9340,N_8024,N_8231);
and U9341 (N_9341,N_8316,N_8092);
or U9342 (N_9342,N_8433,N_8412);
nor U9343 (N_9343,N_8694,N_8704);
xor U9344 (N_9344,N_8497,N_8053);
nor U9345 (N_9345,N_8478,N_8452);
xor U9346 (N_9346,N_8779,N_8421);
or U9347 (N_9347,N_8786,N_8404);
nand U9348 (N_9348,N_8647,N_8165);
and U9349 (N_9349,N_8018,N_8270);
nor U9350 (N_9350,N_8004,N_8693);
nor U9351 (N_9351,N_8651,N_8395);
or U9352 (N_9352,N_8591,N_8516);
and U9353 (N_9353,N_8744,N_8259);
xor U9354 (N_9354,N_8687,N_8616);
nand U9355 (N_9355,N_8760,N_8359);
nand U9356 (N_9356,N_8029,N_8058);
nand U9357 (N_9357,N_8707,N_8708);
nor U9358 (N_9358,N_8746,N_8047);
nor U9359 (N_9359,N_8104,N_8022);
nand U9360 (N_9360,N_8517,N_8246);
and U9361 (N_9361,N_8375,N_8452);
nand U9362 (N_9362,N_8289,N_8789);
nand U9363 (N_9363,N_8104,N_8215);
xor U9364 (N_9364,N_8770,N_8496);
or U9365 (N_9365,N_8419,N_8220);
and U9366 (N_9366,N_8494,N_8059);
xor U9367 (N_9367,N_8050,N_8608);
xnor U9368 (N_9368,N_8214,N_8600);
nor U9369 (N_9369,N_8157,N_8256);
nor U9370 (N_9370,N_8458,N_8294);
nand U9371 (N_9371,N_8007,N_8402);
nand U9372 (N_9372,N_8321,N_8327);
nand U9373 (N_9373,N_8336,N_8743);
and U9374 (N_9374,N_8791,N_8108);
and U9375 (N_9375,N_8308,N_8162);
nor U9376 (N_9376,N_8687,N_8701);
nand U9377 (N_9377,N_8174,N_8795);
nand U9378 (N_9378,N_8669,N_8612);
nor U9379 (N_9379,N_8608,N_8451);
or U9380 (N_9380,N_8183,N_8195);
xnor U9381 (N_9381,N_8066,N_8014);
and U9382 (N_9382,N_8680,N_8377);
or U9383 (N_9383,N_8543,N_8481);
or U9384 (N_9384,N_8382,N_8129);
and U9385 (N_9385,N_8113,N_8604);
nor U9386 (N_9386,N_8772,N_8337);
nor U9387 (N_9387,N_8600,N_8554);
nor U9388 (N_9388,N_8369,N_8395);
or U9389 (N_9389,N_8034,N_8620);
nand U9390 (N_9390,N_8556,N_8164);
and U9391 (N_9391,N_8764,N_8748);
nand U9392 (N_9392,N_8142,N_8565);
xor U9393 (N_9393,N_8514,N_8291);
or U9394 (N_9394,N_8029,N_8418);
or U9395 (N_9395,N_8544,N_8219);
nor U9396 (N_9396,N_8581,N_8704);
and U9397 (N_9397,N_8476,N_8566);
nor U9398 (N_9398,N_8201,N_8237);
nor U9399 (N_9399,N_8352,N_8631);
nor U9400 (N_9400,N_8253,N_8447);
xor U9401 (N_9401,N_8359,N_8049);
or U9402 (N_9402,N_8117,N_8387);
xnor U9403 (N_9403,N_8552,N_8070);
xnor U9404 (N_9404,N_8501,N_8208);
nand U9405 (N_9405,N_8256,N_8165);
and U9406 (N_9406,N_8236,N_8287);
nand U9407 (N_9407,N_8340,N_8699);
nor U9408 (N_9408,N_8170,N_8738);
and U9409 (N_9409,N_8311,N_8693);
nor U9410 (N_9410,N_8422,N_8128);
nor U9411 (N_9411,N_8773,N_8576);
xnor U9412 (N_9412,N_8174,N_8747);
nand U9413 (N_9413,N_8681,N_8342);
or U9414 (N_9414,N_8422,N_8785);
nand U9415 (N_9415,N_8361,N_8707);
and U9416 (N_9416,N_8124,N_8204);
or U9417 (N_9417,N_8568,N_8253);
and U9418 (N_9418,N_8247,N_8597);
xnor U9419 (N_9419,N_8347,N_8266);
or U9420 (N_9420,N_8475,N_8777);
nand U9421 (N_9421,N_8019,N_8608);
nand U9422 (N_9422,N_8521,N_8722);
nand U9423 (N_9423,N_8257,N_8033);
and U9424 (N_9424,N_8178,N_8639);
xor U9425 (N_9425,N_8505,N_8253);
nand U9426 (N_9426,N_8676,N_8026);
or U9427 (N_9427,N_8290,N_8234);
xnor U9428 (N_9428,N_8769,N_8586);
or U9429 (N_9429,N_8780,N_8194);
nand U9430 (N_9430,N_8195,N_8303);
nand U9431 (N_9431,N_8407,N_8678);
nor U9432 (N_9432,N_8000,N_8593);
and U9433 (N_9433,N_8132,N_8420);
nor U9434 (N_9434,N_8581,N_8607);
xnor U9435 (N_9435,N_8016,N_8100);
or U9436 (N_9436,N_8524,N_8478);
and U9437 (N_9437,N_8607,N_8413);
xor U9438 (N_9438,N_8665,N_8035);
nor U9439 (N_9439,N_8019,N_8099);
or U9440 (N_9440,N_8604,N_8655);
nor U9441 (N_9441,N_8080,N_8048);
nand U9442 (N_9442,N_8536,N_8202);
and U9443 (N_9443,N_8166,N_8131);
nor U9444 (N_9444,N_8430,N_8317);
and U9445 (N_9445,N_8436,N_8364);
xnor U9446 (N_9446,N_8341,N_8690);
nor U9447 (N_9447,N_8789,N_8522);
nand U9448 (N_9448,N_8287,N_8172);
and U9449 (N_9449,N_8100,N_8020);
or U9450 (N_9450,N_8535,N_8719);
and U9451 (N_9451,N_8494,N_8484);
nand U9452 (N_9452,N_8190,N_8562);
and U9453 (N_9453,N_8398,N_8780);
and U9454 (N_9454,N_8028,N_8474);
xnor U9455 (N_9455,N_8143,N_8638);
or U9456 (N_9456,N_8002,N_8471);
nor U9457 (N_9457,N_8363,N_8133);
nand U9458 (N_9458,N_8408,N_8574);
and U9459 (N_9459,N_8070,N_8392);
or U9460 (N_9460,N_8218,N_8334);
and U9461 (N_9461,N_8012,N_8317);
xor U9462 (N_9462,N_8732,N_8245);
xnor U9463 (N_9463,N_8747,N_8786);
or U9464 (N_9464,N_8151,N_8484);
and U9465 (N_9465,N_8504,N_8556);
xnor U9466 (N_9466,N_8499,N_8198);
nor U9467 (N_9467,N_8076,N_8355);
and U9468 (N_9468,N_8554,N_8481);
nand U9469 (N_9469,N_8067,N_8046);
or U9470 (N_9470,N_8560,N_8098);
nand U9471 (N_9471,N_8404,N_8340);
xor U9472 (N_9472,N_8793,N_8026);
nor U9473 (N_9473,N_8701,N_8390);
or U9474 (N_9474,N_8478,N_8143);
xor U9475 (N_9475,N_8597,N_8256);
or U9476 (N_9476,N_8074,N_8080);
or U9477 (N_9477,N_8336,N_8320);
xor U9478 (N_9478,N_8733,N_8067);
nand U9479 (N_9479,N_8411,N_8105);
and U9480 (N_9480,N_8370,N_8651);
nand U9481 (N_9481,N_8332,N_8112);
nor U9482 (N_9482,N_8681,N_8221);
and U9483 (N_9483,N_8427,N_8498);
and U9484 (N_9484,N_8118,N_8511);
or U9485 (N_9485,N_8626,N_8370);
and U9486 (N_9486,N_8504,N_8435);
or U9487 (N_9487,N_8696,N_8642);
xor U9488 (N_9488,N_8424,N_8519);
or U9489 (N_9489,N_8140,N_8024);
and U9490 (N_9490,N_8199,N_8644);
xor U9491 (N_9491,N_8030,N_8478);
nor U9492 (N_9492,N_8446,N_8343);
or U9493 (N_9493,N_8662,N_8634);
or U9494 (N_9494,N_8044,N_8561);
and U9495 (N_9495,N_8495,N_8031);
and U9496 (N_9496,N_8369,N_8269);
and U9497 (N_9497,N_8148,N_8693);
or U9498 (N_9498,N_8327,N_8416);
nor U9499 (N_9499,N_8498,N_8609);
or U9500 (N_9500,N_8592,N_8700);
nand U9501 (N_9501,N_8612,N_8666);
nand U9502 (N_9502,N_8353,N_8762);
and U9503 (N_9503,N_8146,N_8281);
nor U9504 (N_9504,N_8419,N_8119);
nand U9505 (N_9505,N_8731,N_8220);
nor U9506 (N_9506,N_8624,N_8160);
and U9507 (N_9507,N_8682,N_8083);
xor U9508 (N_9508,N_8375,N_8368);
or U9509 (N_9509,N_8549,N_8053);
or U9510 (N_9510,N_8068,N_8608);
and U9511 (N_9511,N_8688,N_8674);
nand U9512 (N_9512,N_8335,N_8439);
xnor U9513 (N_9513,N_8178,N_8794);
or U9514 (N_9514,N_8448,N_8219);
and U9515 (N_9515,N_8155,N_8451);
nor U9516 (N_9516,N_8145,N_8216);
or U9517 (N_9517,N_8481,N_8120);
or U9518 (N_9518,N_8161,N_8250);
nand U9519 (N_9519,N_8483,N_8269);
or U9520 (N_9520,N_8156,N_8637);
nand U9521 (N_9521,N_8650,N_8617);
xor U9522 (N_9522,N_8387,N_8291);
or U9523 (N_9523,N_8049,N_8692);
or U9524 (N_9524,N_8145,N_8590);
nand U9525 (N_9525,N_8568,N_8216);
nor U9526 (N_9526,N_8142,N_8784);
xnor U9527 (N_9527,N_8274,N_8169);
and U9528 (N_9528,N_8308,N_8715);
or U9529 (N_9529,N_8154,N_8644);
nand U9530 (N_9530,N_8174,N_8692);
and U9531 (N_9531,N_8058,N_8449);
or U9532 (N_9532,N_8208,N_8443);
nand U9533 (N_9533,N_8422,N_8038);
xnor U9534 (N_9534,N_8482,N_8213);
and U9535 (N_9535,N_8236,N_8154);
and U9536 (N_9536,N_8629,N_8150);
and U9537 (N_9537,N_8223,N_8714);
xnor U9538 (N_9538,N_8712,N_8719);
xor U9539 (N_9539,N_8123,N_8634);
xor U9540 (N_9540,N_8394,N_8663);
xor U9541 (N_9541,N_8783,N_8069);
and U9542 (N_9542,N_8365,N_8095);
nand U9543 (N_9543,N_8289,N_8033);
nor U9544 (N_9544,N_8132,N_8346);
nand U9545 (N_9545,N_8103,N_8204);
and U9546 (N_9546,N_8735,N_8435);
nand U9547 (N_9547,N_8094,N_8699);
or U9548 (N_9548,N_8616,N_8296);
or U9549 (N_9549,N_8316,N_8134);
nand U9550 (N_9550,N_8051,N_8130);
or U9551 (N_9551,N_8243,N_8445);
xnor U9552 (N_9552,N_8492,N_8042);
nor U9553 (N_9553,N_8378,N_8706);
nor U9554 (N_9554,N_8763,N_8395);
nand U9555 (N_9555,N_8616,N_8667);
or U9556 (N_9556,N_8236,N_8477);
or U9557 (N_9557,N_8592,N_8394);
nor U9558 (N_9558,N_8359,N_8755);
xnor U9559 (N_9559,N_8079,N_8421);
nand U9560 (N_9560,N_8424,N_8585);
nand U9561 (N_9561,N_8385,N_8390);
nor U9562 (N_9562,N_8349,N_8460);
nor U9563 (N_9563,N_8504,N_8394);
xnor U9564 (N_9564,N_8622,N_8013);
nand U9565 (N_9565,N_8795,N_8512);
nand U9566 (N_9566,N_8728,N_8202);
nor U9567 (N_9567,N_8289,N_8505);
nor U9568 (N_9568,N_8640,N_8520);
xor U9569 (N_9569,N_8321,N_8550);
nor U9570 (N_9570,N_8743,N_8210);
nor U9571 (N_9571,N_8678,N_8424);
xor U9572 (N_9572,N_8075,N_8280);
nor U9573 (N_9573,N_8069,N_8431);
or U9574 (N_9574,N_8340,N_8643);
xnor U9575 (N_9575,N_8334,N_8027);
nand U9576 (N_9576,N_8052,N_8164);
nor U9577 (N_9577,N_8746,N_8650);
or U9578 (N_9578,N_8775,N_8597);
xor U9579 (N_9579,N_8500,N_8485);
xnor U9580 (N_9580,N_8552,N_8393);
nand U9581 (N_9581,N_8278,N_8573);
xor U9582 (N_9582,N_8599,N_8308);
nand U9583 (N_9583,N_8266,N_8753);
nor U9584 (N_9584,N_8656,N_8717);
and U9585 (N_9585,N_8777,N_8289);
nand U9586 (N_9586,N_8084,N_8224);
nand U9587 (N_9587,N_8675,N_8369);
xor U9588 (N_9588,N_8218,N_8074);
xor U9589 (N_9589,N_8149,N_8331);
and U9590 (N_9590,N_8304,N_8619);
xnor U9591 (N_9591,N_8075,N_8431);
and U9592 (N_9592,N_8605,N_8334);
or U9593 (N_9593,N_8448,N_8034);
and U9594 (N_9594,N_8362,N_8543);
or U9595 (N_9595,N_8426,N_8381);
and U9596 (N_9596,N_8676,N_8590);
nor U9597 (N_9597,N_8111,N_8047);
nor U9598 (N_9598,N_8550,N_8035);
xor U9599 (N_9599,N_8581,N_8646);
or U9600 (N_9600,N_9475,N_9117);
and U9601 (N_9601,N_9197,N_9295);
or U9602 (N_9602,N_9551,N_9587);
xnor U9603 (N_9603,N_8885,N_9177);
or U9604 (N_9604,N_9502,N_8833);
xor U9605 (N_9605,N_9353,N_9289);
nand U9606 (N_9606,N_9188,N_9150);
or U9607 (N_9607,N_9156,N_8804);
and U9608 (N_9608,N_9566,N_9416);
nand U9609 (N_9609,N_8802,N_9064);
xor U9610 (N_9610,N_9506,N_8835);
nand U9611 (N_9611,N_9179,N_8925);
nand U9612 (N_9612,N_8811,N_8810);
nand U9613 (N_9613,N_9075,N_9272);
or U9614 (N_9614,N_9074,N_8886);
and U9615 (N_9615,N_9067,N_9335);
or U9616 (N_9616,N_9020,N_8901);
nand U9617 (N_9617,N_9255,N_9414);
and U9618 (N_9618,N_8836,N_9286);
and U9619 (N_9619,N_9223,N_8911);
and U9620 (N_9620,N_9128,N_8954);
or U9621 (N_9621,N_9509,N_8859);
and U9622 (N_9622,N_9523,N_9080);
and U9623 (N_9623,N_9470,N_8867);
or U9624 (N_9624,N_8921,N_9142);
nor U9625 (N_9625,N_9168,N_9578);
xnor U9626 (N_9626,N_9112,N_9015);
xnor U9627 (N_9627,N_9077,N_8861);
and U9628 (N_9628,N_9119,N_8838);
nor U9629 (N_9629,N_9013,N_9448);
or U9630 (N_9630,N_9061,N_9530);
xor U9631 (N_9631,N_8904,N_9468);
or U9632 (N_9632,N_8840,N_9497);
and U9633 (N_9633,N_8971,N_9565);
nand U9634 (N_9634,N_9171,N_9224);
xor U9635 (N_9635,N_8842,N_8941);
xnor U9636 (N_9636,N_8984,N_8860);
nor U9637 (N_9637,N_9437,N_8889);
nor U9638 (N_9638,N_8931,N_9323);
or U9639 (N_9639,N_8878,N_9352);
or U9640 (N_9640,N_9256,N_9594);
and U9641 (N_9641,N_8905,N_8936);
or U9642 (N_9642,N_9111,N_9181);
nor U9643 (N_9643,N_9248,N_9203);
xnor U9644 (N_9644,N_8942,N_9398);
nand U9645 (N_9645,N_9133,N_9554);
nor U9646 (N_9646,N_9297,N_9182);
nand U9647 (N_9647,N_9520,N_9158);
nor U9648 (N_9648,N_9311,N_9556);
and U9649 (N_9649,N_8816,N_9490);
xnor U9650 (N_9650,N_9407,N_9134);
nand U9651 (N_9651,N_9474,N_9400);
or U9652 (N_9652,N_8837,N_9366);
nand U9653 (N_9653,N_9595,N_9447);
nor U9654 (N_9654,N_9382,N_8934);
nor U9655 (N_9655,N_8903,N_9079);
and U9656 (N_9656,N_9550,N_9324);
nand U9657 (N_9657,N_9145,N_9419);
nor U9658 (N_9658,N_9331,N_9193);
and U9659 (N_9659,N_9371,N_9599);
nand U9660 (N_9660,N_9545,N_9521);
nand U9661 (N_9661,N_8820,N_9264);
nand U9662 (N_9662,N_9425,N_9147);
nor U9663 (N_9663,N_9000,N_9001);
and U9664 (N_9664,N_9367,N_9065);
xor U9665 (N_9665,N_8800,N_9327);
nor U9666 (N_9666,N_9279,N_9163);
xnor U9667 (N_9667,N_9436,N_9040);
xnor U9668 (N_9668,N_9380,N_8868);
nor U9669 (N_9669,N_9183,N_9273);
or U9670 (N_9670,N_9066,N_9069);
xnor U9671 (N_9671,N_8956,N_9581);
or U9672 (N_9672,N_9118,N_9591);
and U9673 (N_9673,N_9276,N_9009);
xor U9674 (N_9674,N_9317,N_9413);
or U9675 (N_9675,N_8897,N_9008);
and U9676 (N_9676,N_9121,N_8808);
and U9677 (N_9677,N_9073,N_9477);
and U9678 (N_9678,N_8947,N_8992);
nand U9679 (N_9679,N_9549,N_9430);
and U9680 (N_9680,N_9541,N_9123);
nor U9681 (N_9681,N_9356,N_9589);
or U9682 (N_9682,N_9495,N_8955);
nand U9683 (N_9683,N_9592,N_9051);
xor U9684 (N_9684,N_9338,N_9101);
or U9685 (N_9685,N_9078,N_9479);
or U9686 (N_9686,N_9499,N_9472);
and U9687 (N_9687,N_9035,N_9127);
and U9688 (N_9688,N_9387,N_9303);
nand U9689 (N_9689,N_9391,N_9573);
or U9690 (N_9690,N_9138,N_9143);
nor U9691 (N_9691,N_9024,N_9396);
or U9692 (N_9692,N_9226,N_8969);
nor U9693 (N_9693,N_9236,N_9410);
nor U9694 (N_9694,N_9007,N_9357);
nand U9695 (N_9695,N_8985,N_8929);
xnor U9696 (N_9696,N_8855,N_9308);
nor U9697 (N_9697,N_9374,N_9494);
or U9698 (N_9698,N_9508,N_8932);
or U9699 (N_9699,N_9211,N_9486);
nor U9700 (N_9700,N_9593,N_9381);
or U9701 (N_9701,N_9271,N_9547);
xor U9702 (N_9702,N_8953,N_8866);
and U9703 (N_9703,N_8862,N_9116);
and U9704 (N_9704,N_9326,N_9318);
or U9705 (N_9705,N_8926,N_9084);
xor U9706 (N_9706,N_9500,N_9044);
xor U9707 (N_9707,N_9011,N_8832);
nor U9708 (N_9708,N_9423,N_9483);
xor U9709 (N_9709,N_9584,N_9053);
xnor U9710 (N_9710,N_9103,N_9379);
nand U9711 (N_9711,N_9048,N_9131);
nor U9712 (N_9712,N_9515,N_8875);
nand U9713 (N_9713,N_9165,N_8857);
or U9714 (N_9714,N_9401,N_8966);
xnor U9715 (N_9715,N_9316,N_9322);
and U9716 (N_9716,N_9070,N_8960);
xnor U9717 (N_9717,N_9346,N_9350);
nand U9718 (N_9718,N_9347,N_8891);
xor U9719 (N_9719,N_9055,N_8809);
nand U9720 (N_9720,N_8963,N_9014);
and U9721 (N_9721,N_9451,N_9473);
nor U9722 (N_9722,N_9538,N_8846);
nor U9723 (N_9723,N_9298,N_9384);
or U9724 (N_9724,N_9296,N_8848);
nor U9725 (N_9725,N_9590,N_9212);
or U9726 (N_9726,N_9245,N_9415);
nand U9727 (N_9727,N_9375,N_9480);
xnor U9728 (N_9728,N_9247,N_9220);
nand U9729 (N_9729,N_9567,N_9453);
and U9730 (N_9730,N_8807,N_9540);
nand U9731 (N_9731,N_9446,N_8928);
nand U9732 (N_9732,N_9113,N_8962);
xnor U9733 (N_9733,N_8959,N_9155);
nand U9734 (N_9734,N_8937,N_9516);
nand U9735 (N_9735,N_9114,N_9358);
nor U9736 (N_9736,N_9083,N_9229);
nor U9737 (N_9737,N_9086,N_9124);
xnor U9738 (N_9738,N_9093,N_8986);
nand U9739 (N_9739,N_9032,N_9263);
xor U9740 (N_9740,N_9343,N_8918);
nand U9741 (N_9741,N_9246,N_9485);
nand U9742 (N_9742,N_9028,N_8923);
xnor U9743 (N_9743,N_9033,N_9056);
or U9744 (N_9744,N_8914,N_9433);
xor U9745 (N_9745,N_8823,N_9225);
xor U9746 (N_9746,N_8999,N_9240);
xnor U9747 (N_9747,N_8844,N_8972);
nand U9748 (N_9748,N_9186,N_9207);
or U9749 (N_9749,N_9478,N_9402);
or U9750 (N_9750,N_8913,N_9238);
and U9751 (N_9751,N_9090,N_8919);
nor U9752 (N_9752,N_9409,N_9002);
nand U9753 (N_9753,N_9404,N_9522);
and U9754 (N_9754,N_9458,N_9052);
nor U9755 (N_9755,N_8948,N_9455);
nor U9756 (N_9756,N_8871,N_9561);
nor U9757 (N_9757,N_9062,N_9144);
xor U9758 (N_9758,N_9089,N_9196);
nand U9759 (N_9759,N_8806,N_8949);
xor U9760 (N_9760,N_8829,N_9059);
and U9761 (N_9761,N_9249,N_9022);
or U9762 (N_9762,N_9135,N_9016);
and U9763 (N_9763,N_9095,N_9426);
or U9764 (N_9764,N_9385,N_9088);
xnor U9765 (N_9765,N_9208,N_9046);
xor U9766 (N_9766,N_9464,N_9319);
nand U9767 (N_9767,N_8847,N_9369);
or U9768 (N_9768,N_9287,N_9087);
xor U9769 (N_9769,N_8916,N_9222);
and U9770 (N_9770,N_9363,N_9463);
or U9771 (N_9771,N_9017,N_9570);
and U9772 (N_9772,N_8815,N_9159);
and U9773 (N_9773,N_8817,N_9325);
nor U9774 (N_9774,N_9452,N_9460);
nor U9775 (N_9775,N_8998,N_8909);
nand U9776 (N_9776,N_9031,N_9206);
or U9777 (N_9777,N_9493,N_8858);
and U9778 (N_9778,N_8907,N_9459);
or U9779 (N_9779,N_9050,N_9261);
and U9780 (N_9780,N_9543,N_9192);
nor U9781 (N_9781,N_9529,N_8818);
and U9782 (N_9782,N_9341,N_9300);
or U9783 (N_9783,N_9553,N_9106);
nand U9784 (N_9784,N_8912,N_8958);
xnor U9785 (N_9785,N_9390,N_9166);
or U9786 (N_9786,N_9408,N_9443);
nand U9787 (N_9787,N_9337,N_8803);
nand U9788 (N_9788,N_9422,N_8964);
and U9789 (N_9789,N_8924,N_9176);
or U9790 (N_9790,N_9244,N_8852);
xor U9791 (N_9791,N_9492,N_8906);
nand U9792 (N_9792,N_9585,N_9498);
nand U9793 (N_9793,N_9354,N_8888);
or U9794 (N_9794,N_9030,N_9057);
or U9795 (N_9795,N_9394,N_8967);
xor U9796 (N_9796,N_9038,N_9189);
or U9797 (N_9797,N_9162,N_9397);
nand U9798 (N_9798,N_9228,N_9466);
xnor U9799 (N_9799,N_9250,N_9227);
or U9800 (N_9800,N_9429,N_9568);
xor U9801 (N_9801,N_8910,N_9098);
or U9802 (N_9802,N_8896,N_9577);
xor U9803 (N_9803,N_8883,N_9469);
nand U9804 (N_9804,N_9488,N_9569);
or U9805 (N_9805,N_9536,N_9097);
or U9806 (N_9806,N_9370,N_9491);
nor U9807 (N_9807,N_9524,N_9285);
or U9808 (N_9808,N_9198,N_8977);
nor U9809 (N_9809,N_9525,N_8996);
nor U9810 (N_9810,N_9457,N_8987);
nand U9811 (N_9811,N_8973,N_9081);
xnor U9812 (N_9812,N_9294,N_9281);
nand U9813 (N_9813,N_9213,N_9005);
nand U9814 (N_9814,N_9544,N_9006);
and U9815 (N_9815,N_9094,N_9428);
or U9816 (N_9816,N_9068,N_9299);
nor U9817 (N_9817,N_9372,N_9424);
nand U9818 (N_9818,N_8821,N_9180);
and U9819 (N_9819,N_9596,N_8841);
xnor U9820 (N_9820,N_9539,N_9243);
nor U9821 (N_9821,N_9257,N_9377);
xnor U9822 (N_9822,N_9432,N_9489);
xnor U9823 (N_9823,N_9531,N_8944);
or U9824 (N_9824,N_9364,N_9102);
and U9825 (N_9825,N_8850,N_8880);
and U9826 (N_9826,N_8863,N_9586);
or U9827 (N_9827,N_8899,N_9125);
and U9828 (N_9828,N_9563,N_9167);
nand U9829 (N_9829,N_9290,N_8873);
nand U9830 (N_9830,N_8814,N_8957);
nor U9831 (N_9831,N_9512,N_9267);
or U9832 (N_9832,N_9321,N_9235);
nand U9833 (N_9833,N_9418,N_9292);
and U9834 (N_9834,N_9392,N_9012);
nand U9835 (N_9835,N_8943,N_9412);
xor U9836 (N_9836,N_9063,N_9164);
xor U9837 (N_9837,N_9120,N_9152);
xnor U9838 (N_9838,N_9018,N_9535);
nor U9839 (N_9839,N_8872,N_9200);
or U9840 (N_9840,N_9362,N_9293);
and U9841 (N_9841,N_9388,N_8991);
nor U9842 (N_9842,N_9395,N_9376);
nor U9843 (N_9843,N_9058,N_8945);
nand U9844 (N_9844,N_8952,N_9170);
xnor U9845 (N_9845,N_9484,N_9571);
nand U9846 (N_9846,N_9010,N_9234);
nor U9847 (N_9847,N_9481,N_9221);
nand U9848 (N_9848,N_8870,N_9190);
nand U9849 (N_9849,N_9204,N_9329);
nor U9850 (N_9850,N_9252,N_8865);
xnor U9851 (N_9851,N_9233,N_8995);
nand U9852 (N_9852,N_9450,N_9588);
and U9853 (N_9853,N_8882,N_8893);
nand U9854 (N_9854,N_9487,N_9438);
nor U9855 (N_9855,N_9383,N_8939);
nor U9856 (N_9856,N_9314,N_9187);
nor U9857 (N_9857,N_9173,N_9503);
nand U9858 (N_9858,N_9306,N_8849);
xnor U9859 (N_9859,N_8851,N_8974);
nand U9860 (N_9860,N_9456,N_9332);
nand U9861 (N_9861,N_9291,N_9036);
nand U9862 (N_9862,N_9185,N_8978);
and U9863 (N_9863,N_9154,N_9361);
and U9864 (N_9864,N_9442,N_9108);
xor U9865 (N_9865,N_8898,N_9260);
and U9866 (N_9866,N_8938,N_9403);
nor U9867 (N_9867,N_8895,N_8994);
xor U9868 (N_9868,N_9071,N_9060);
nor U9869 (N_9869,N_9148,N_8813);
and U9870 (N_9870,N_9519,N_9580);
or U9871 (N_9871,N_9386,N_8831);
and U9872 (N_9872,N_8902,N_8864);
xor U9873 (N_9873,N_9399,N_9471);
nand U9874 (N_9874,N_8981,N_8968);
or U9875 (N_9875,N_9340,N_8982);
nand U9876 (N_9876,N_9462,N_9355);
and U9877 (N_9877,N_8819,N_8980);
nor U9878 (N_9878,N_9411,N_8997);
nand U9879 (N_9879,N_9039,N_9439);
nand U9880 (N_9880,N_9461,N_9099);
nand U9881 (N_9881,N_8917,N_9542);
xor U9882 (N_9882,N_9169,N_8827);
and U9883 (N_9883,N_9305,N_8881);
and U9884 (N_9884,N_9269,N_9534);
nor U9885 (N_9885,N_9026,N_9107);
nor U9886 (N_9886,N_9199,N_9476);
and U9887 (N_9887,N_9546,N_8908);
or U9888 (N_9888,N_8884,N_8874);
and U9889 (N_9889,N_9122,N_9251);
and U9890 (N_9890,N_9184,N_8983);
nand U9891 (N_9891,N_8900,N_8839);
nor U9892 (N_9892,N_9049,N_9096);
xor U9893 (N_9893,N_9021,N_9130);
nand U9894 (N_9894,N_9427,N_9351);
nand U9895 (N_9895,N_9559,N_9526);
or U9896 (N_9896,N_9435,N_8979);
xnor U9897 (N_9897,N_9076,N_9149);
or U9898 (N_9898,N_9172,N_8856);
nor U9899 (N_9899,N_9085,N_9420);
xnor U9900 (N_9900,N_9239,N_9598);
nand U9901 (N_9901,N_9178,N_9518);
or U9902 (N_9902,N_9034,N_8843);
xnor U9903 (N_9903,N_9365,N_9575);
nand U9904 (N_9904,N_9449,N_9205);
or U9905 (N_9905,N_9348,N_9342);
xnor U9906 (N_9906,N_9309,N_9231);
or U9907 (N_9907,N_9557,N_8933);
nand U9908 (N_9908,N_9023,N_9140);
nand U9909 (N_9909,N_9537,N_8890);
xor U9910 (N_9910,N_9282,N_9045);
nor U9911 (N_9911,N_8812,N_9266);
xor U9912 (N_9912,N_9393,N_9548);
nor U9913 (N_9913,N_9174,N_9440);
nor U9914 (N_9914,N_8920,N_9219);
and U9915 (N_9915,N_8927,N_9389);
and U9916 (N_9916,N_8834,N_8965);
nand U9917 (N_9917,N_8975,N_9270);
nand U9918 (N_9918,N_9560,N_9302);
or U9919 (N_9919,N_9027,N_9501);
and U9920 (N_9920,N_8951,N_9445);
nor U9921 (N_9921,N_9334,N_9025);
and U9922 (N_9922,N_8869,N_8830);
and U9923 (N_9923,N_9406,N_8922);
xnor U9924 (N_9924,N_9232,N_9041);
xnor U9925 (N_9925,N_9517,N_9315);
and U9926 (N_9926,N_9265,N_9194);
nand U9927 (N_9927,N_8828,N_9161);
nand U9928 (N_9928,N_8877,N_9202);
xnor U9929 (N_9929,N_9216,N_8915);
or U9930 (N_9930,N_9209,N_8988);
or U9931 (N_9931,N_9558,N_9528);
nor U9932 (N_9932,N_9339,N_9141);
nor U9933 (N_9933,N_9359,N_9328);
and U9934 (N_9934,N_9082,N_9333);
and U9935 (N_9935,N_9230,N_9237);
or U9936 (N_9936,N_9310,N_9431);
nand U9937 (N_9937,N_8824,N_8822);
xor U9938 (N_9938,N_8854,N_8940);
or U9939 (N_9939,N_9283,N_9307);
or U9940 (N_9940,N_9160,N_8930);
and U9941 (N_9941,N_9268,N_9597);
xor U9942 (N_9942,N_9003,N_9054);
nand U9943 (N_9943,N_9241,N_9504);
xor U9944 (N_9944,N_9109,N_8805);
nand U9945 (N_9945,N_9210,N_9368);
or U9946 (N_9946,N_9320,N_9583);
nand U9947 (N_9947,N_8935,N_9242);
nand U9948 (N_9948,N_9574,N_9507);
xnor U9949 (N_9949,N_9579,N_9373);
nand U9950 (N_9950,N_9072,N_9254);
nor U9951 (N_9951,N_9218,N_9284);
or U9952 (N_9952,N_9511,N_9129);
or U9953 (N_9953,N_9100,N_9091);
xnor U9954 (N_9954,N_9288,N_9146);
or U9955 (N_9955,N_8976,N_8970);
nor U9956 (N_9956,N_8887,N_9110);
nand U9957 (N_9957,N_9482,N_9454);
nor U9958 (N_9958,N_9572,N_9465);
nand U9959 (N_9959,N_9301,N_9037);
nor U9960 (N_9960,N_8961,N_9582);
nor U9961 (N_9961,N_9304,N_9275);
nor U9962 (N_9962,N_9496,N_9153);
or U9963 (N_9963,N_8989,N_9157);
nor U9964 (N_9964,N_9405,N_9029);
xor U9965 (N_9965,N_9104,N_9562);
or U9966 (N_9966,N_9533,N_9042);
nand U9967 (N_9967,N_8801,N_8879);
and U9968 (N_9968,N_9552,N_9201);
and U9969 (N_9969,N_9278,N_8853);
nor U9970 (N_9970,N_9043,N_9345);
xnor U9971 (N_9971,N_9312,N_9564);
and U9972 (N_9972,N_9258,N_9195);
and U9973 (N_9973,N_9259,N_8876);
and U9974 (N_9974,N_9092,N_9467);
xnor U9975 (N_9975,N_9274,N_9417);
nor U9976 (N_9976,N_9262,N_8993);
nor U9977 (N_9977,N_8894,N_9105);
nor U9978 (N_9978,N_9019,N_8950);
xnor U9979 (N_9979,N_9510,N_9151);
nor U9980 (N_9980,N_9137,N_9513);
or U9981 (N_9981,N_8825,N_9555);
nand U9982 (N_9982,N_9215,N_9505);
and U9983 (N_9983,N_8845,N_9421);
xor U9984 (N_9984,N_9360,N_9336);
and U9985 (N_9985,N_9378,N_9175);
and U9986 (N_9986,N_9434,N_9527);
nor U9987 (N_9987,N_9514,N_9277);
or U9988 (N_9988,N_8892,N_9313);
and U9989 (N_9989,N_9441,N_9136);
xnor U9990 (N_9990,N_8946,N_9132);
and U9991 (N_9991,N_9004,N_9047);
nor U9992 (N_9992,N_9344,N_8990);
nand U9993 (N_9993,N_9126,N_9191);
or U9994 (N_9994,N_8826,N_9217);
xnor U9995 (N_9995,N_9115,N_9139);
nor U9996 (N_9996,N_9280,N_9532);
nor U9997 (N_9997,N_9253,N_9349);
xnor U9998 (N_9998,N_9444,N_9576);
or U9999 (N_9999,N_9330,N_9214);
nor U10000 (N_10000,N_8821,N_9027);
and U10001 (N_10001,N_8930,N_9350);
nor U10002 (N_10002,N_9226,N_8875);
xnor U10003 (N_10003,N_9419,N_9118);
nand U10004 (N_10004,N_9020,N_8827);
xnor U10005 (N_10005,N_9532,N_9144);
nand U10006 (N_10006,N_8906,N_8856);
nand U10007 (N_10007,N_9598,N_9254);
or U10008 (N_10008,N_8880,N_8966);
xnor U10009 (N_10009,N_9427,N_8935);
xor U10010 (N_10010,N_9068,N_8956);
nor U10011 (N_10011,N_9352,N_9545);
nor U10012 (N_10012,N_8885,N_8974);
nor U10013 (N_10013,N_8834,N_9322);
or U10014 (N_10014,N_9504,N_9102);
xor U10015 (N_10015,N_9372,N_9558);
nand U10016 (N_10016,N_9041,N_9102);
and U10017 (N_10017,N_9566,N_8912);
xnor U10018 (N_10018,N_8803,N_9384);
xnor U10019 (N_10019,N_8938,N_9518);
and U10020 (N_10020,N_9061,N_8923);
nand U10021 (N_10021,N_8882,N_8974);
xor U10022 (N_10022,N_9389,N_9212);
xnor U10023 (N_10023,N_9298,N_9019);
nand U10024 (N_10024,N_9066,N_9386);
xor U10025 (N_10025,N_9576,N_8814);
nand U10026 (N_10026,N_9350,N_9402);
nor U10027 (N_10027,N_8818,N_9249);
or U10028 (N_10028,N_9388,N_8825);
and U10029 (N_10029,N_8974,N_9574);
and U10030 (N_10030,N_9448,N_9237);
and U10031 (N_10031,N_8850,N_8993);
nor U10032 (N_10032,N_9512,N_8800);
nor U10033 (N_10033,N_9596,N_8959);
xnor U10034 (N_10034,N_9212,N_8891);
or U10035 (N_10035,N_9299,N_8995);
and U10036 (N_10036,N_9291,N_9235);
nor U10037 (N_10037,N_8819,N_9382);
xor U10038 (N_10038,N_9167,N_8914);
nand U10039 (N_10039,N_8864,N_8818);
nor U10040 (N_10040,N_9388,N_9091);
nor U10041 (N_10041,N_9230,N_9260);
and U10042 (N_10042,N_9258,N_9465);
xnor U10043 (N_10043,N_9082,N_9266);
nand U10044 (N_10044,N_9407,N_9191);
or U10045 (N_10045,N_9060,N_9184);
and U10046 (N_10046,N_9394,N_9311);
nand U10047 (N_10047,N_9232,N_9142);
nor U10048 (N_10048,N_8897,N_8941);
or U10049 (N_10049,N_9055,N_9372);
or U10050 (N_10050,N_8815,N_8937);
or U10051 (N_10051,N_9071,N_9339);
nor U10052 (N_10052,N_9438,N_9499);
and U10053 (N_10053,N_9058,N_9549);
or U10054 (N_10054,N_9288,N_9309);
and U10055 (N_10055,N_9361,N_8993);
xor U10056 (N_10056,N_9024,N_8905);
nand U10057 (N_10057,N_9454,N_9367);
and U10058 (N_10058,N_9363,N_8852);
or U10059 (N_10059,N_9152,N_9430);
xnor U10060 (N_10060,N_9286,N_9411);
nor U10061 (N_10061,N_9130,N_9276);
xor U10062 (N_10062,N_8822,N_8806);
nand U10063 (N_10063,N_8814,N_8901);
nand U10064 (N_10064,N_9281,N_9118);
and U10065 (N_10065,N_9471,N_8978);
nor U10066 (N_10066,N_9480,N_9542);
nor U10067 (N_10067,N_8803,N_9327);
nor U10068 (N_10068,N_9422,N_9181);
nand U10069 (N_10069,N_8936,N_9171);
and U10070 (N_10070,N_9046,N_9188);
or U10071 (N_10071,N_9084,N_9162);
or U10072 (N_10072,N_9209,N_9114);
xnor U10073 (N_10073,N_9326,N_9085);
nand U10074 (N_10074,N_9039,N_9100);
or U10075 (N_10075,N_9569,N_8921);
or U10076 (N_10076,N_9547,N_9451);
nor U10077 (N_10077,N_9404,N_9240);
nand U10078 (N_10078,N_9387,N_9032);
or U10079 (N_10079,N_9168,N_9191);
nand U10080 (N_10080,N_9085,N_8883);
nand U10081 (N_10081,N_9482,N_9545);
and U10082 (N_10082,N_8897,N_9285);
nor U10083 (N_10083,N_9146,N_8870);
and U10084 (N_10084,N_9262,N_9003);
nand U10085 (N_10085,N_8981,N_8850);
or U10086 (N_10086,N_9474,N_9193);
xor U10087 (N_10087,N_9308,N_9205);
and U10088 (N_10088,N_9221,N_9374);
nand U10089 (N_10089,N_8911,N_8993);
and U10090 (N_10090,N_9554,N_9536);
and U10091 (N_10091,N_9217,N_9160);
or U10092 (N_10092,N_9393,N_8825);
nand U10093 (N_10093,N_8884,N_9430);
nand U10094 (N_10094,N_9262,N_9548);
and U10095 (N_10095,N_9158,N_9078);
and U10096 (N_10096,N_9143,N_9348);
xnor U10097 (N_10097,N_8905,N_9526);
or U10098 (N_10098,N_8918,N_9404);
xnor U10099 (N_10099,N_9506,N_9212);
xor U10100 (N_10100,N_9290,N_9222);
nand U10101 (N_10101,N_8895,N_9296);
xor U10102 (N_10102,N_9315,N_9541);
nor U10103 (N_10103,N_9073,N_8887);
xor U10104 (N_10104,N_9058,N_9102);
and U10105 (N_10105,N_9568,N_9360);
and U10106 (N_10106,N_9304,N_8832);
xor U10107 (N_10107,N_9204,N_8820);
or U10108 (N_10108,N_8919,N_9232);
xor U10109 (N_10109,N_9077,N_8925);
nor U10110 (N_10110,N_9072,N_9599);
and U10111 (N_10111,N_9422,N_9482);
and U10112 (N_10112,N_9495,N_9453);
xnor U10113 (N_10113,N_9104,N_9037);
nand U10114 (N_10114,N_9445,N_9161);
xor U10115 (N_10115,N_9422,N_9087);
nor U10116 (N_10116,N_8994,N_9540);
nor U10117 (N_10117,N_9540,N_9594);
or U10118 (N_10118,N_8823,N_9279);
or U10119 (N_10119,N_9291,N_9261);
xor U10120 (N_10120,N_9298,N_9213);
or U10121 (N_10121,N_9063,N_9348);
or U10122 (N_10122,N_8996,N_9388);
or U10123 (N_10123,N_9400,N_9079);
and U10124 (N_10124,N_9591,N_9572);
and U10125 (N_10125,N_9251,N_9546);
xnor U10126 (N_10126,N_8945,N_8873);
nor U10127 (N_10127,N_9134,N_9307);
nor U10128 (N_10128,N_8875,N_9334);
nor U10129 (N_10129,N_9128,N_9020);
or U10130 (N_10130,N_9518,N_9484);
nand U10131 (N_10131,N_9267,N_9496);
nor U10132 (N_10132,N_9202,N_8907);
xnor U10133 (N_10133,N_8811,N_9565);
nand U10134 (N_10134,N_8860,N_9510);
or U10135 (N_10135,N_9510,N_9252);
xnor U10136 (N_10136,N_8987,N_9591);
and U10137 (N_10137,N_9124,N_9210);
xor U10138 (N_10138,N_9457,N_9138);
or U10139 (N_10139,N_9190,N_9163);
and U10140 (N_10140,N_9210,N_8864);
xnor U10141 (N_10141,N_9473,N_8810);
xnor U10142 (N_10142,N_9166,N_9452);
xor U10143 (N_10143,N_9103,N_8871);
nor U10144 (N_10144,N_8999,N_9442);
nand U10145 (N_10145,N_8940,N_8815);
nor U10146 (N_10146,N_9589,N_8907);
nand U10147 (N_10147,N_8928,N_8877);
or U10148 (N_10148,N_9262,N_9545);
nand U10149 (N_10149,N_9078,N_8800);
and U10150 (N_10150,N_9238,N_9378);
or U10151 (N_10151,N_9059,N_9292);
and U10152 (N_10152,N_9487,N_9044);
or U10153 (N_10153,N_9403,N_8869);
or U10154 (N_10154,N_9245,N_8842);
nand U10155 (N_10155,N_9498,N_8950);
or U10156 (N_10156,N_9229,N_8869);
xor U10157 (N_10157,N_9134,N_9492);
xor U10158 (N_10158,N_9303,N_8813);
nor U10159 (N_10159,N_9494,N_9090);
or U10160 (N_10160,N_8970,N_9243);
nor U10161 (N_10161,N_9154,N_8923);
nor U10162 (N_10162,N_8941,N_8930);
xnor U10163 (N_10163,N_9585,N_8899);
xnor U10164 (N_10164,N_9090,N_8904);
xnor U10165 (N_10165,N_8964,N_8824);
xor U10166 (N_10166,N_8877,N_9496);
nand U10167 (N_10167,N_8969,N_9313);
or U10168 (N_10168,N_9386,N_9510);
and U10169 (N_10169,N_9192,N_9577);
xor U10170 (N_10170,N_9179,N_9122);
nor U10171 (N_10171,N_9004,N_9048);
or U10172 (N_10172,N_9218,N_8914);
nand U10173 (N_10173,N_9299,N_9483);
and U10174 (N_10174,N_9109,N_8824);
xnor U10175 (N_10175,N_9423,N_9592);
xor U10176 (N_10176,N_9049,N_9156);
xnor U10177 (N_10177,N_8821,N_9000);
or U10178 (N_10178,N_9243,N_9279);
nor U10179 (N_10179,N_9539,N_9187);
nand U10180 (N_10180,N_8978,N_8943);
nand U10181 (N_10181,N_9291,N_9000);
xor U10182 (N_10182,N_9504,N_9599);
xor U10183 (N_10183,N_9409,N_9267);
or U10184 (N_10184,N_8954,N_9052);
or U10185 (N_10185,N_9310,N_8855);
nand U10186 (N_10186,N_9043,N_9516);
and U10187 (N_10187,N_9286,N_9299);
xor U10188 (N_10188,N_8969,N_9289);
or U10189 (N_10189,N_9502,N_9028);
xor U10190 (N_10190,N_9274,N_9438);
or U10191 (N_10191,N_9051,N_9520);
xnor U10192 (N_10192,N_9344,N_9051);
nor U10193 (N_10193,N_9279,N_8901);
and U10194 (N_10194,N_9398,N_9133);
nor U10195 (N_10195,N_8815,N_9041);
and U10196 (N_10196,N_8867,N_9180);
and U10197 (N_10197,N_8813,N_9532);
xor U10198 (N_10198,N_8876,N_9286);
nor U10199 (N_10199,N_9297,N_8863);
and U10200 (N_10200,N_9566,N_9032);
xor U10201 (N_10201,N_8864,N_9264);
nor U10202 (N_10202,N_9367,N_9373);
nor U10203 (N_10203,N_9295,N_9047);
nand U10204 (N_10204,N_9240,N_8930);
nand U10205 (N_10205,N_9599,N_8915);
and U10206 (N_10206,N_9368,N_9325);
nand U10207 (N_10207,N_8979,N_9213);
nor U10208 (N_10208,N_9074,N_9005);
or U10209 (N_10209,N_9298,N_9415);
or U10210 (N_10210,N_9037,N_9005);
or U10211 (N_10211,N_8803,N_9219);
or U10212 (N_10212,N_8833,N_8856);
nand U10213 (N_10213,N_9200,N_9036);
and U10214 (N_10214,N_9591,N_9410);
and U10215 (N_10215,N_8879,N_9425);
or U10216 (N_10216,N_8859,N_9510);
nor U10217 (N_10217,N_9269,N_8986);
or U10218 (N_10218,N_9434,N_9215);
and U10219 (N_10219,N_9274,N_8831);
xnor U10220 (N_10220,N_9218,N_9097);
and U10221 (N_10221,N_9107,N_9051);
nor U10222 (N_10222,N_8981,N_8992);
xnor U10223 (N_10223,N_8911,N_9087);
or U10224 (N_10224,N_9162,N_9359);
nand U10225 (N_10225,N_9132,N_8910);
or U10226 (N_10226,N_8859,N_9182);
xnor U10227 (N_10227,N_9221,N_9331);
nand U10228 (N_10228,N_9451,N_8933);
or U10229 (N_10229,N_9403,N_9155);
nor U10230 (N_10230,N_8920,N_9351);
xnor U10231 (N_10231,N_9315,N_8854);
nand U10232 (N_10232,N_8970,N_9252);
nor U10233 (N_10233,N_9371,N_9056);
nor U10234 (N_10234,N_8940,N_8990);
nand U10235 (N_10235,N_9344,N_8915);
and U10236 (N_10236,N_8844,N_9390);
nor U10237 (N_10237,N_9193,N_9156);
or U10238 (N_10238,N_9078,N_9502);
xor U10239 (N_10239,N_9559,N_9505);
nand U10240 (N_10240,N_8937,N_8922);
and U10241 (N_10241,N_9517,N_9004);
xor U10242 (N_10242,N_9006,N_9056);
nor U10243 (N_10243,N_9011,N_8994);
and U10244 (N_10244,N_9319,N_9599);
or U10245 (N_10245,N_9354,N_9448);
nor U10246 (N_10246,N_8812,N_9122);
xnor U10247 (N_10247,N_8869,N_9166);
and U10248 (N_10248,N_8889,N_9338);
nand U10249 (N_10249,N_8885,N_9283);
nand U10250 (N_10250,N_9127,N_9247);
xor U10251 (N_10251,N_8888,N_9417);
nand U10252 (N_10252,N_9366,N_9238);
and U10253 (N_10253,N_9090,N_9197);
or U10254 (N_10254,N_9349,N_9365);
and U10255 (N_10255,N_9386,N_9126);
xor U10256 (N_10256,N_9128,N_8966);
or U10257 (N_10257,N_9199,N_9146);
and U10258 (N_10258,N_9186,N_9263);
or U10259 (N_10259,N_9029,N_9195);
nor U10260 (N_10260,N_9435,N_9595);
and U10261 (N_10261,N_9197,N_9298);
and U10262 (N_10262,N_8893,N_9162);
nor U10263 (N_10263,N_8829,N_9468);
or U10264 (N_10264,N_9079,N_9179);
or U10265 (N_10265,N_9007,N_9552);
nand U10266 (N_10266,N_9448,N_9238);
nand U10267 (N_10267,N_9390,N_9551);
or U10268 (N_10268,N_9245,N_8965);
or U10269 (N_10269,N_8979,N_9335);
and U10270 (N_10270,N_9066,N_8920);
and U10271 (N_10271,N_8998,N_9462);
xnor U10272 (N_10272,N_8997,N_8867);
and U10273 (N_10273,N_9292,N_9062);
xor U10274 (N_10274,N_9391,N_8933);
xnor U10275 (N_10275,N_9400,N_9394);
xor U10276 (N_10276,N_9266,N_9120);
nor U10277 (N_10277,N_9433,N_9015);
and U10278 (N_10278,N_9258,N_8869);
nand U10279 (N_10279,N_8935,N_8987);
and U10280 (N_10280,N_9192,N_8893);
nor U10281 (N_10281,N_9068,N_9085);
and U10282 (N_10282,N_9057,N_8900);
nand U10283 (N_10283,N_9234,N_8992);
nor U10284 (N_10284,N_8912,N_9099);
and U10285 (N_10285,N_9198,N_9343);
nor U10286 (N_10286,N_9431,N_8866);
or U10287 (N_10287,N_9071,N_9208);
nand U10288 (N_10288,N_9508,N_9282);
or U10289 (N_10289,N_9181,N_8970);
or U10290 (N_10290,N_9513,N_9073);
nand U10291 (N_10291,N_9517,N_9152);
xnor U10292 (N_10292,N_8809,N_9140);
xnor U10293 (N_10293,N_9485,N_9322);
nor U10294 (N_10294,N_9572,N_8814);
and U10295 (N_10295,N_9578,N_9204);
nand U10296 (N_10296,N_9535,N_8868);
nor U10297 (N_10297,N_9252,N_9009);
nor U10298 (N_10298,N_8952,N_9165);
and U10299 (N_10299,N_9213,N_9366);
nor U10300 (N_10300,N_9534,N_8881);
xnor U10301 (N_10301,N_8985,N_9533);
xor U10302 (N_10302,N_9573,N_8802);
and U10303 (N_10303,N_9560,N_9536);
nand U10304 (N_10304,N_9455,N_9109);
nor U10305 (N_10305,N_9039,N_9170);
nand U10306 (N_10306,N_9178,N_9097);
or U10307 (N_10307,N_8982,N_9188);
xnor U10308 (N_10308,N_9088,N_9337);
nand U10309 (N_10309,N_9403,N_9458);
or U10310 (N_10310,N_9434,N_9008);
and U10311 (N_10311,N_9326,N_9417);
nand U10312 (N_10312,N_9231,N_9114);
xnor U10313 (N_10313,N_8945,N_8822);
nand U10314 (N_10314,N_9342,N_8994);
and U10315 (N_10315,N_9120,N_9153);
and U10316 (N_10316,N_8961,N_8973);
or U10317 (N_10317,N_9409,N_8890);
nor U10318 (N_10318,N_9172,N_9585);
nand U10319 (N_10319,N_9151,N_9324);
xnor U10320 (N_10320,N_8998,N_8888);
and U10321 (N_10321,N_9169,N_9166);
nand U10322 (N_10322,N_8857,N_9293);
nor U10323 (N_10323,N_9290,N_9029);
xor U10324 (N_10324,N_8982,N_8921);
xor U10325 (N_10325,N_9275,N_9153);
xor U10326 (N_10326,N_9466,N_9527);
and U10327 (N_10327,N_9507,N_8824);
or U10328 (N_10328,N_9051,N_9390);
nor U10329 (N_10329,N_9403,N_8823);
and U10330 (N_10330,N_9299,N_8827);
nand U10331 (N_10331,N_8826,N_9052);
nor U10332 (N_10332,N_9503,N_9486);
nor U10333 (N_10333,N_9303,N_9514);
or U10334 (N_10334,N_8894,N_9529);
xnor U10335 (N_10335,N_9373,N_9042);
xor U10336 (N_10336,N_9599,N_9004);
and U10337 (N_10337,N_9536,N_9474);
nor U10338 (N_10338,N_9407,N_9186);
or U10339 (N_10339,N_9136,N_8883);
xnor U10340 (N_10340,N_9532,N_8810);
nand U10341 (N_10341,N_8940,N_9264);
or U10342 (N_10342,N_9223,N_8921);
nand U10343 (N_10343,N_8906,N_9514);
and U10344 (N_10344,N_9339,N_8996);
or U10345 (N_10345,N_9195,N_8898);
or U10346 (N_10346,N_9507,N_9067);
and U10347 (N_10347,N_9317,N_9055);
or U10348 (N_10348,N_9461,N_9310);
or U10349 (N_10349,N_8802,N_9312);
nand U10350 (N_10350,N_9254,N_9321);
and U10351 (N_10351,N_9273,N_9027);
or U10352 (N_10352,N_9288,N_9484);
nor U10353 (N_10353,N_9486,N_9005);
nand U10354 (N_10354,N_9394,N_9263);
and U10355 (N_10355,N_9318,N_9245);
and U10356 (N_10356,N_8944,N_9420);
and U10357 (N_10357,N_9532,N_8937);
or U10358 (N_10358,N_9206,N_9202);
or U10359 (N_10359,N_9061,N_9592);
xnor U10360 (N_10360,N_9116,N_9341);
nor U10361 (N_10361,N_9500,N_9226);
or U10362 (N_10362,N_9369,N_8859);
xor U10363 (N_10363,N_8858,N_9491);
xor U10364 (N_10364,N_9458,N_8970);
or U10365 (N_10365,N_9523,N_8950);
xor U10366 (N_10366,N_9330,N_8919);
or U10367 (N_10367,N_8912,N_9320);
nand U10368 (N_10368,N_8951,N_9242);
and U10369 (N_10369,N_9426,N_9518);
nand U10370 (N_10370,N_9498,N_9218);
or U10371 (N_10371,N_9276,N_9238);
nand U10372 (N_10372,N_9248,N_9360);
nand U10373 (N_10373,N_9198,N_9258);
nor U10374 (N_10374,N_9573,N_8832);
or U10375 (N_10375,N_9333,N_8931);
nand U10376 (N_10376,N_9393,N_8918);
or U10377 (N_10377,N_9548,N_8839);
nand U10378 (N_10378,N_9247,N_9175);
or U10379 (N_10379,N_9069,N_9130);
xor U10380 (N_10380,N_9279,N_9094);
or U10381 (N_10381,N_9318,N_9482);
xor U10382 (N_10382,N_8980,N_9398);
nor U10383 (N_10383,N_9017,N_9326);
or U10384 (N_10384,N_9318,N_9323);
or U10385 (N_10385,N_9263,N_8908);
or U10386 (N_10386,N_9125,N_9329);
nand U10387 (N_10387,N_9095,N_9211);
xor U10388 (N_10388,N_9236,N_9495);
xnor U10389 (N_10389,N_9386,N_9325);
and U10390 (N_10390,N_9172,N_9096);
xor U10391 (N_10391,N_9299,N_9287);
or U10392 (N_10392,N_9312,N_9138);
xnor U10393 (N_10393,N_9337,N_9448);
nor U10394 (N_10394,N_9487,N_9007);
nor U10395 (N_10395,N_9047,N_8963);
nand U10396 (N_10396,N_9129,N_9030);
and U10397 (N_10397,N_9051,N_8918);
nor U10398 (N_10398,N_9076,N_9121);
and U10399 (N_10399,N_8985,N_9182);
nand U10400 (N_10400,N_10125,N_10139);
nand U10401 (N_10401,N_9818,N_9715);
and U10402 (N_10402,N_10208,N_9705);
or U10403 (N_10403,N_10345,N_9634);
and U10404 (N_10404,N_9768,N_9970);
xor U10405 (N_10405,N_9743,N_9793);
xor U10406 (N_10406,N_9624,N_10335);
nand U10407 (N_10407,N_9933,N_9686);
and U10408 (N_10408,N_9968,N_10079);
xnor U10409 (N_10409,N_9943,N_10106);
or U10410 (N_10410,N_9709,N_9742);
nor U10411 (N_10411,N_10020,N_10098);
xor U10412 (N_10412,N_10096,N_9910);
and U10413 (N_10413,N_9826,N_9744);
xnor U10414 (N_10414,N_10391,N_10319);
nand U10415 (N_10415,N_10305,N_9936);
or U10416 (N_10416,N_10193,N_9628);
and U10417 (N_10417,N_9856,N_10119);
xnor U10418 (N_10418,N_9736,N_10276);
and U10419 (N_10419,N_9913,N_10390);
nand U10420 (N_10420,N_9948,N_9771);
xor U10421 (N_10421,N_10171,N_10097);
and U10422 (N_10422,N_10282,N_10051);
xor U10423 (N_10423,N_9923,N_10281);
nand U10424 (N_10424,N_9710,N_9642);
or U10425 (N_10425,N_10374,N_9956);
or U10426 (N_10426,N_9617,N_9753);
nor U10427 (N_10427,N_10185,N_9799);
xor U10428 (N_10428,N_10304,N_10315);
or U10429 (N_10429,N_10126,N_10052);
nand U10430 (N_10430,N_10389,N_10267);
nand U10431 (N_10431,N_9606,N_10303);
or U10432 (N_10432,N_9700,N_10346);
nor U10433 (N_10433,N_10060,N_9684);
nand U10434 (N_10434,N_10279,N_9932);
or U10435 (N_10435,N_9635,N_9747);
nor U10436 (N_10436,N_10366,N_9735);
nand U10437 (N_10437,N_9612,N_9695);
nand U10438 (N_10438,N_9891,N_10294);
xnor U10439 (N_10439,N_10198,N_9730);
nand U10440 (N_10440,N_9934,N_10061);
or U10441 (N_10441,N_9692,N_10036);
xor U10442 (N_10442,N_10118,N_9655);
xnor U10443 (N_10443,N_10383,N_10209);
nor U10444 (N_10444,N_9912,N_10155);
or U10445 (N_10445,N_9806,N_10067);
xor U10446 (N_10446,N_9690,N_10316);
or U10447 (N_10447,N_10013,N_10202);
or U10448 (N_10448,N_10095,N_10221);
xor U10449 (N_10449,N_10252,N_9832);
xnor U10450 (N_10450,N_10322,N_10260);
and U10451 (N_10451,N_10004,N_10270);
or U10452 (N_10452,N_9696,N_9754);
and U10453 (N_10453,N_9904,N_10189);
xnor U10454 (N_10454,N_9967,N_10249);
nor U10455 (N_10455,N_10138,N_9972);
and U10456 (N_10456,N_10076,N_10320);
nor U10457 (N_10457,N_10378,N_9999);
or U10458 (N_10458,N_9966,N_10114);
nand U10459 (N_10459,N_9610,N_10234);
nor U10460 (N_10460,N_9662,N_10168);
or U10461 (N_10461,N_9924,N_9600);
xor U10462 (N_10462,N_10088,N_10222);
nand U10463 (N_10463,N_10159,N_9830);
xnor U10464 (N_10464,N_9660,N_10170);
nand U10465 (N_10465,N_9725,N_9882);
or U10466 (N_10466,N_9755,N_10003);
nor U10467 (N_10467,N_9955,N_10367);
nor U10468 (N_10468,N_9960,N_10115);
xor U10469 (N_10469,N_9845,N_9998);
and U10470 (N_10470,N_9841,N_10082);
or U10471 (N_10471,N_10018,N_10008);
nand U10472 (N_10472,N_9925,N_10100);
or U10473 (N_10473,N_9985,N_9680);
nand U10474 (N_10474,N_10215,N_10257);
and U10475 (N_10475,N_10205,N_10056);
nand U10476 (N_10476,N_10362,N_9727);
nand U10477 (N_10477,N_9773,N_10317);
nor U10478 (N_10478,N_10207,N_9720);
nand U10479 (N_10479,N_10031,N_10373);
nand U10480 (N_10480,N_9976,N_10089);
xnor U10481 (N_10481,N_10151,N_10360);
and U10482 (N_10482,N_9828,N_9822);
nand U10483 (N_10483,N_10358,N_9693);
and U10484 (N_10484,N_9641,N_9993);
xor U10485 (N_10485,N_10246,N_9905);
nor U10486 (N_10486,N_10102,N_9670);
xor U10487 (N_10487,N_10025,N_9643);
or U10488 (N_10488,N_10191,N_10262);
xor U10489 (N_10489,N_10005,N_10081);
nor U10490 (N_10490,N_10295,N_10214);
nand U10491 (N_10491,N_9875,N_9937);
or U10492 (N_10492,N_10230,N_10296);
nor U10493 (N_10493,N_9638,N_10277);
or U10494 (N_10494,N_9876,N_10064);
xor U10495 (N_10495,N_9677,N_9848);
nor U10496 (N_10496,N_9810,N_10349);
nor U10497 (N_10497,N_10261,N_9951);
nor U10498 (N_10498,N_10359,N_10328);
nor U10499 (N_10499,N_10121,N_9605);
nor U10500 (N_10500,N_10128,N_9780);
xnor U10501 (N_10501,N_9863,N_10188);
xnor U10502 (N_10502,N_9833,N_10053);
and U10503 (N_10503,N_9859,N_9911);
nor U10504 (N_10504,N_10110,N_10393);
xor U10505 (N_10505,N_9865,N_9774);
and U10506 (N_10506,N_9654,N_10132);
nand U10507 (N_10507,N_10045,N_9988);
nor U10508 (N_10508,N_9920,N_9615);
nand U10509 (N_10509,N_10156,N_9982);
and U10510 (N_10510,N_10157,N_9853);
nand U10511 (N_10511,N_10376,N_10101);
and U10512 (N_10512,N_9931,N_9922);
nor U10513 (N_10513,N_10306,N_10321);
xor U10514 (N_10514,N_10072,N_10184);
or U10515 (N_10515,N_9842,N_9778);
xor U10516 (N_10516,N_9792,N_9881);
and U10517 (N_10517,N_9728,N_10268);
xnor U10518 (N_10518,N_9941,N_10135);
and U10519 (N_10519,N_9873,N_9813);
nor U10520 (N_10520,N_10247,N_9629);
or U10521 (N_10521,N_10255,N_9867);
and U10522 (N_10522,N_9883,N_9978);
and U10523 (N_10523,N_10200,N_9779);
nand U10524 (N_10524,N_9839,N_9691);
nand U10525 (N_10525,N_10112,N_9829);
and U10526 (N_10526,N_9711,N_10023);
xnor U10527 (N_10527,N_10394,N_9917);
xnor U10528 (N_10528,N_10326,N_9887);
nor U10529 (N_10529,N_9639,N_9992);
nand U10530 (N_10530,N_10329,N_9994);
nor U10531 (N_10531,N_9620,N_10049);
and U10532 (N_10532,N_10299,N_10007);
xor U10533 (N_10533,N_10154,N_9697);
and U10534 (N_10534,N_10382,N_9740);
xnor U10535 (N_10535,N_10127,N_10340);
nor U10536 (N_10536,N_10371,N_9947);
nor U10537 (N_10537,N_9989,N_10080);
nand U10538 (N_10538,N_10289,N_10104);
nor U10539 (N_10539,N_9834,N_10074);
xor U10540 (N_10540,N_10334,N_9869);
xnor U10541 (N_10541,N_10010,N_10284);
nor U10542 (N_10542,N_9731,N_9894);
or U10543 (N_10543,N_10369,N_9798);
nor U10544 (N_10544,N_10269,N_10077);
xnor U10545 (N_10545,N_9987,N_9666);
or U10546 (N_10546,N_10350,N_9827);
nand U10547 (N_10547,N_10197,N_10105);
xnor U10548 (N_10548,N_10271,N_10111);
xnor U10549 (N_10549,N_10054,N_9878);
or U10550 (N_10550,N_10177,N_10314);
and U10551 (N_10551,N_10001,N_9930);
xnor U10552 (N_10552,N_9678,N_10062);
nor U10553 (N_10553,N_9738,N_10122);
and U10554 (N_10554,N_9946,N_9651);
and U10555 (N_10555,N_9734,N_9864);
nor U10556 (N_10556,N_10203,N_9892);
nand U10557 (N_10557,N_10307,N_9979);
or U10558 (N_10558,N_10273,N_9761);
or U10559 (N_10559,N_10002,N_9926);
nor U10560 (N_10560,N_9657,N_9969);
or U10561 (N_10561,N_10172,N_9723);
and U10562 (N_10562,N_10363,N_10368);
and U10563 (N_10563,N_9851,N_10057);
nand U10564 (N_10564,N_9961,N_10011);
or U10565 (N_10565,N_10140,N_10204);
nand U10566 (N_10566,N_10009,N_10375);
and U10567 (N_10567,N_10278,N_10050);
xor U10568 (N_10568,N_9921,N_10264);
nor U10569 (N_10569,N_9759,N_10006);
xnor U10570 (N_10570,N_9840,N_9850);
nor U10571 (N_10571,N_10353,N_10137);
nand U10572 (N_10572,N_9766,N_9732);
or U10573 (N_10573,N_10292,N_10186);
nand U10574 (N_10574,N_9667,N_9811);
nor U10575 (N_10575,N_10165,N_10083);
nand U10576 (N_10576,N_10206,N_10163);
or U10577 (N_10577,N_10336,N_9675);
and U10578 (N_10578,N_10381,N_9957);
nor U10579 (N_10579,N_10372,N_9718);
xnor U10580 (N_10580,N_9614,N_9964);
or U10581 (N_10581,N_10136,N_10038);
nand U10582 (N_10582,N_9739,N_10178);
nand U10583 (N_10583,N_10377,N_10392);
or U10584 (N_10584,N_9746,N_10028);
nand U10585 (N_10585,N_9627,N_10245);
xnor U10586 (N_10586,N_9789,N_10235);
and U10587 (N_10587,N_9602,N_10047);
nor U10588 (N_10588,N_9689,N_9914);
and U10589 (N_10589,N_9682,N_9698);
and U10590 (N_10590,N_9819,N_10216);
nor U10591 (N_10591,N_9973,N_9794);
or U10592 (N_10592,N_9939,N_9986);
nand U10593 (N_10593,N_10103,N_10091);
and U10594 (N_10594,N_9611,N_9650);
and U10595 (N_10595,N_9748,N_10039);
nand U10596 (N_10596,N_9616,N_10248);
nor U10597 (N_10597,N_10030,N_9907);
nand U10598 (N_10598,N_10070,N_9984);
nor U10599 (N_10599,N_9704,N_9645);
or U10600 (N_10600,N_10174,N_9805);
or U10601 (N_10601,N_9906,N_9980);
nand U10602 (N_10602,N_9676,N_10229);
nor U10603 (N_10603,N_9659,N_9637);
and U10604 (N_10604,N_9749,N_10032);
and U10605 (N_10605,N_9880,N_9706);
nand U10606 (N_10606,N_10120,N_9656);
xor U10607 (N_10607,N_10312,N_10055);
nand U10608 (N_10608,N_10133,N_10352);
nor U10609 (N_10609,N_10141,N_9847);
nor U10610 (N_10610,N_10256,N_10272);
nand U10611 (N_10611,N_9928,N_9765);
or U10612 (N_10612,N_10169,N_9940);
or U10613 (N_10613,N_9633,N_9714);
xnor U10614 (N_10614,N_10148,N_9983);
or U10615 (N_10615,N_9658,N_9702);
xnor U10616 (N_10616,N_9608,N_9750);
nor U10617 (N_10617,N_9942,N_9935);
and U10618 (N_10618,N_9663,N_9609);
and U10619 (N_10619,N_10339,N_9688);
nand U10620 (N_10620,N_9803,N_9716);
xor U10621 (N_10621,N_10073,N_9717);
nand U10622 (N_10622,N_9699,N_10090);
or U10623 (N_10623,N_10014,N_10201);
or U10624 (N_10624,N_10078,N_9665);
or U10625 (N_10625,N_9944,N_9896);
nor U10626 (N_10626,N_9997,N_9927);
or U10627 (N_10627,N_9713,N_10265);
nor U10628 (N_10628,N_10325,N_9855);
or U10629 (N_10629,N_10068,N_10243);
or U10630 (N_10630,N_9787,N_9919);
nor U10631 (N_10631,N_10293,N_10129);
and U10632 (N_10632,N_10254,N_10324);
nand U10633 (N_10633,N_10274,N_9604);
xor U10634 (N_10634,N_10175,N_10343);
nand U10635 (N_10635,N_9965,N_10259);
nand U10636 (N_10636,N_10370,N_9722);
and U10637 (N_10637,N_10354,N_10242);
or U10638 (N_10638,N_10232,N_10179);
nand U10639 (N_10639,N_10173,N_9632);
nor U10640 (N_10640,N_9795,N_10237);
xor U10641 (N_10641,N_10046,N_9900);
nand U10642 (N_10642,N_10117,N_9764);
xor U10643 (N_10643,N_10026,N_9797);
nand U10644 (N_10644,N_10220,N_9648);
xor U10645 (N_10645,N_10355,N_10071);
nor U10646 (N_10646,N_9949,N_9756);
nor U10647 (N_10647,N_9679,N_10286);
and U10648 (N_10648,N_10338,N_9915);
nor U10649 (N_10649,N_9975,N_9995);
or U10650 (N_10650,N_9758,N_10399);
nand U10651 (N_10651,N_10379,N_10227);
nand U10652 (N_10652,N_9953,N_10164);
nand U10653 (N_10653,N_10143,N_9785);
and U10654 (N_10654,N_10094,N_10093);
nand U10655 (N_10655,N_9821,N_9647);
xnor U10656 (N_10656,N_10251,N_9607);
xnor U10657 (N_10657,N_10182,N_10160);
nand U10658 (N_10658,N_9777,N_10063);
xor U10659 (N_10659,N_9962,N_10145);
and U10660 (N_10660,N_10142,N_9825);
nor U10661 (N_10661,N_10302,N_10059);
nand U10662 (N_10662,N_10194,N_10134);
or U10663 (N_10663,N_9959,N_10146);
and U10664 (N_10664,N_9603,N_10042);
xnor U10665 (N_10665,N_10395,N_9719);
nand U10666 (N_10666,N_9752,N_10034);
nor U10667 (N_10667,N_10219,N_9877);
nor U10668 (N_10668,N_10266,N_9858);
xnor U10669 (N_10669,N_10183,N_9636);
xnor U10670 (N_10670,N_10043,N_10092);
and U10671 (N_10671,N_9938,N_9644);
xnor U10672 (N_10672,N_9971,N_9741);
nor U10673 (N_10673,N_10087,N_9762);
nor U10674 (N_10674,N_9886,N_10385);
xor U10675 (N_10675,N_10301,N_9884);
and U10676 (N_10676,N_10396,N_10015);
and U10677 (N_10677,N_10361,N_9668);
nor U10678 (N_10678,N_9804,N_9945);
or U10679 (N_10679,N_9673,N_10029);
nand U10680 (N_10680,N_10075,N_10233);
or U10681 (N_10681,N_9823,N_10113);
xor U10682 (N_10682,N_10176,N_10019);
xnor U10683 (N_10683,N_10309,N_9909);
and U10684 (N_10684,N_9885,N_10150);
nand U10685 (N_10685,N_9929,N_9849);
nor U10686 (N_10686,N_10228,N_10158);
xor U10687 (N_10687,N_10297,N_10351);
nand U10688 (N_10688,N_10180,N_9661);
nor U10689 (N_10689,N_9775,N_10040);
nand U10690 (N_10690,N_9852,N_10287);
xor U10691 (N_10691,N_9838,N_10365);
or U10692 (N_10692,N_10199,N_9619);
and U10693 (N_10693,N_9950,N_9640);
xnor U10694 (N_10694,N_10226,N_10224);
or U10695 (N_10695,N_9649,N_9807);
nor U10696 (N_10696,N_9981,N_9908);
nor U10697 (N_10697,N_10211,N_9862);
and U10698 (N_10698,N_9890,N_9788);
nor U10699 (N_10699,N_9770,N_9767);
nor U10700 (N_10700,N_9703,N_9801);
and U10701 (N_10701,N_9796,N_9854);
nor U10702 (N_10702,N_9958,N_9751);
nor U10703 (N_10703,N_10217,N_9835);
xor U10704 (N_10704,N_10181,N_9815);
or U10705 (N_10705,N_9701,N_9729);
xor U10706 (N_10706,N_10167,N_9843);
and U10707 (N_10707,N_9860,N_9707);
and U10708 (N_10708,N_10311,N_9721);
nor U10709 (N_10709,N_10263,N_10318);
or U10710 (N_10710,N_10241,N_9664);
nand U10711 (N_10711,N_10323,N_9622);
xnor U10712 (N_10712,N_10161,N_9808);
and U10713 (N_10713,N_10069,N_9836);
and U10714 (N_10714,N_10313,N_10238);
nand U10715 (N_10715,N_9776,N_10310);
nand U10716 (N_10716,N_10398,N_9824);
xnor U10717 (N_10717,N_9990,N_9745);
nor U10718 (N_10718,N_10342,N_9674);
or U10719 (N_10719,N_10290,N_10331);
nor U10720 (N_10720,N_10024,N_10231);
or U10721 (N_10721,N_9772,N_10192);
or U10722 (N_10722,N_9652,N_10308);
xor U10723 (N_10723,N_9814,N_10327);
or U10724 (N_10724,N_9618,N_9952);
xor U10725 (N_10725,N_10131,N_9800);
or U10726 (N_10726,N_9871,N_10275);
or U10727 (N_10727,N_9724,N_10330);
xnor U10728 (N_10728,N_9837,N_9630);
nand U10729 (N_10729,N_9898,N_9726);
xnor U10730 (N_10730,N_10347,N_10384);
and U10731 (N_10731,N_9737,N_9763);
or U10732 (N_10732,N_10344,N_9977);
nand U10733 (N_10733,N_10190,N_9902);
xnor U10734 (N_10734,N_9760,N_9790);
xnor U10735 (N_10735,N_9916,N_10058);
and U10736 (N_10736,N_9782,N_10107);
nand U10737 (N_10737,N_9672,N_9954);
and U10738 (N_10738,N_9872,N_10213);
xor U10739 (N_10739,N_10223,N_10152);
nor U10740 (N_10740,N_9897,N_10041);
xor U10741 (N_10741,N_9626,N_9996);
nand U10742 (N_10742,N_9903,N_9861);
nand U10743 (N_10743,N_10017,N_10357);
or U10744 (N_10744,N_10035,N_10124);
or U10745 (N_10745,N_10250,N_10291);
and U10746 (N_10746,N_10337,N_9646);
or U10747 (N_10747,N_9653,N_9809);
and U10748 (N_10748,N_10196,N_10244);
xnor U10749 (N_10749,N_10225,N_9757);
or U10750 (N_10750,N_9781,N_9817);
xor U10751 (N_10751,N_10283,N_9991);
and U10752 (N_10752,N_9613,N_10066);
nand U10753 (N_10753,N_9708,N_10195);
nand U10754 (N_10754,N_10000,N_10348);
xnor U10755 (N_10755,N_9868,N_9918);
and U10756 (N_10756,N_9786,N_9870);
or U10757 (N_10757,N_9812,N_9784);
xor U10758 (N_10758,N_9791,N_10086);
or U10759 (N_10759,N_10253,N_9769);
or U10760 (N_10760,N_10187,N_9820);
nand U10761 (N_10761,N_9866,N_10044);
and U10762 (N_10762,N_10332,N_9625);
or U10763 (N_10763,N_10147,N_10166);
nand U10764 (N_10764,N_10239,N_10099);
nand U10765 (N_10765,N_10298,N_10258);
nor U10766 (N_10766,N_9895,N_9857);
xnor U10767 (N_10767,N_10012,N_10387);
and U10768 (N_10768,N_9802,N_10144);
nand U10769 (N_10769,N_10212,N_9974);
or U10770 (N_10770,N_9889,N_10123);
nor U10771 (N_10771,N_10341,N_9888);
nand U10772 (N_10772,N_10162,N_10149);
nor U10773 (N_10773,N_9669,N_10210);
or U10774 (N_10774,N_10218,N_9631);
nor U10775 (N_10775,N_10397,N_9694);
nor U10776 (N_10776,N_9683,N_10037);
xor U10777 (N_10777,N_9601,N_10021);
and U10778 (N_10778,N_10022,N_10085);
nor U10779 (N_10779,N_10130,N_9621);
nand U10780 (N_10780,N_10300,N_10333);
or U10781 (N_10781,N_9846,N_9671);
and U10782 (N_10782,N_10236,N_9733);
or U10783 (N_10783,N_10288,N_10388);
or U10784 (N_10784,N_10027,N_10380);
and U10785 (N_10785,N_10065,N_10153);
xor U10786 (N_10786,N_9681,N_10116);
nand U10787 (N_10787,N_9874,N_10285);
nand U10788 (N_10788,N_10033,N_9963);
nor U10789 (N_10789,N_10016,N_10084);
nor U10790 (N_10790,N_9623,N_9901);
xnor U10791 (N_10791,N_10280,N_9685);
and U10792 (N_10792,N_9712,N_9687);
and U10793 (N_10793,N_9893,N_9899);
xnor U10794 (N_10794,N_9879,N_10356);
xor U10795 (N_10795,N_10048,N_10108);
or U10796 (N_10796,N_10386,N_10109);
xor U10797 (N_10797,N_9816,N_9783);
or U10798 (N_10798,N_9831,N_10240);
nor U10799 (N_10799,N_9844,N_10364);
nor U10800 (N_10800,N_10240,N_9893);
or U10801 (N_10801,N_10235,N_10332);
nand U10802 (N_10802,N_9842,N_10246);
or U10803 (N_10803,N_9970,N_9688);
and U10804 (N_10804,N_9986,N_10091);
or U10805 (N_10805,N_10299,N_10288);
or U10806 (N_10806,N_9858,N_9909);
xnor U10807 (N_10807,N_9626,N_9955);
or U10808 (N_10808,N_10261,N_10327);
and U10809 (N_10809,N_10184,N_9803);
or U10810 (N_10810,N_10217,N_9618);
nor U10811 (N_10811,N_9717,N_9924);
nand U10812 (N_10812,N_9680,N_10173);
nand U10813 (N_10813,N_9784,N_10387);
and U10814 (N_10814,N_9954,N_9608);
nor U10815 (N_10815,N_10180,N_9922);
and U10816 (N_10816,N_9694,N_9764);
nor U10817 (N_10817,N_9709,N_10374);
xnor U10818 (N_10818,N_9702,N_9818);
xor U10819 (N_10819,N_9843,N_9819);
nand U10820 (N_10820,N_9734,N_10147);
nor U10821 (N_10821,N_9778,N_10395);
nor U10822 (N_10822,N_10155,N_9850);
xnor U10823 (N_10823,N_10172,N_10352);
or U10824 (N_10824,N_9982,N_10343);
and U10825 (N_10825,N_10152,N_10187);
xor U10826 (N_10826,N_9945,N_10109);
nor U10827 (N_10827,N_9758,N_9952);
or U10828 (N_10828,N_9838,N_10037);
nor U10829 (N_10829,N_10177,N_10396);
nand U10830 (N_10830,N_10126,N_10115);
nand U10831 (N_10831,N_10273,N_9869);
and U10832 (N_10832,N_9789,N_10108);
or U10833 (N_10833,N_9900,N_10306);
nand U10834 (N_10834,N_10086,N_10239);
nand U10835 (N_10835,N_10026,N_9984);
nor U10836 (N_10836,N_9692,N_10364);
xnor U10837 (N_10837,N_10163,N_10397);
and U10838 (N_10838,N_9954,N_9994);
nor U10839 (N_10839,N_10393,N_10306);
and U10840 (N_10840,N_9813,N_9742);
nor U10841 (N_10841,N_9936,N_10343);
or U10842 (N_10842,N_10133,N_10084);
and U10843 (N_10843,N_9714,N_10059);
nand U10844 (N_10844,N_9796,N_9754);
nand U10845 (N_10845,N_9816,N_9821);
or U10846 (N_10846,N_10253,N_9643);
and U10847 (N_10847,N_9791,N_10247);
xor U10848 (N_10848,N_9952,N_10121);
xnor U10849 (N_10849,N_10293,N_10133);
xor U10850 (N_10850,N_10307,N_9724);
nor U10851 (N_10851,N_10266,N_9602);
xnor U10852 (N_10852,N_9910,N_10074);
and U10853 (N_10853,N_10169,N_9862);
and U10854 (N_10854,N_10144,N_10179);
xnor U10855 (N_10855,N_9858,N_9833);
and U10856 (N_10856,N_10263,N_9868);
xor U10857 (N_10857,N_10016,N_9988);
nor U10858 (N_10858,N_10039,N_10061);
nand U10859 (N_10859,N_10141,N_9919);
and U10860 (N_10860,N_9681,N_10341);
xor U10861 (N_10861,N_9645,N_9698);
or U10862 (N_10862,N_9906,N_9898);
xnor U10863 (N_10863,N_9658,N_9745);
and U10864 (N_10864,N_9990,N_10064);
nor U10865 (N_10865,N_9936,N_10007);
nor U10866 (N_10866,N_10045,N_10398);
xnor U10867 (N_10867,N_9779,N_10173);
xnor U10868 (N_10868,N_10273,N_9611);
and U10869 (N_10869,N_10168,N_10075);
nand U10870 (N_10870,N_9682,N_9700);
and U10871 (N_10871,N_9754,N_9740);
nand U10872 (N_10872,N_9736,N_10110);
and U10873 (N_10873,N_10332,N_9771);
or U10874 (N_10874,N_9924,N_9757);
nand U10875 (N_10875,N_10385,N_10240);
and U10876 (N_10876,N_10156,N_9759);
nor U10877 (N_10877,N_9973,N_9725);
nand U10878 (N_10878,N_10082,N_10314);
or U10879 (N_10879,N_9947,N_9646);
xnor U10880 (N_10880,N_10010,N_10275);
nand U10881 (N_10881,N_10252,N_9799);
or U10882 (N_10882,N_9605,N_10003);
nor U10883 (N_10883,N_9888,N_10055);
xor U10884 (N_10884,N_10016,N_9608);
and U10885 (N_10885,N_10172,N_10283);
and U10886 (N_10886,N_9895,N_10315);
and U10887 (N_10887,N_10183,N_10069);
and U10888 (N_10888,N_10321,N_9908);
and U10889 (N_10889,N_9913,N_9630);
and U10890 (N_10890,N_9610,N_10368);
nand U10891 (N_10891,N_10399,N_10117);
or U10892 (N_10892,N_9909,N_10035);
or U10893 (N_10893,N_9901,N_10217);
or U10894 (N_10894,N_9965,N_9621);
nor U10895 (N_10895,N_10284,N_10368);
nor U10896 (N_10896,N_10036,N_9895);
or U10897 (N_10897,N_9651,N_10389);
or U10898 (N_10898,N_9862,N_10094);
nor U10899 (N_10899,N_9653,N_9823);
and U10900 (N_10900,N_9900,N_9807);
nand U10901 (N_10901,N_9791,N_9672);
xor U10902 (N_10902,N_10120,N_10076);
xnor U10903 (N_10903,N_10065,N_10338);
nor U10904 (N_10904,N_10230,N_9754);
and U10905 (N_10905,N_9736,N_10009);
nor U10906 (N_10906,N_9631,N_9735);
or U10907 (N_10907,N_9932,N_9916);
and U10908 (N_10908,N_10340,N_9855);
nand U10909 (N_10909,N_9826,N_10121);
and U10910 (N_10910,N_9967,N_9813);
or U10911 (N_10911,N_10397,N_10381);
nand U10912 (N_10912,N_9610,N_10394);
and U10913 (N_10913,N_10173,N_9659);
or U10914 (N_10914,N_10287,N_9981);
nand U10915 (N_10915,N_10002,N_10087);
and U10916 (N_10916,N_10064,N_9856);
nor U10917 (N_10917,N_9892,N_10306);
or U10918 (N_10918,N_9977,N_10148);
nand U10919 (N_10919,N_10252,N_10181);
and U10920 (N_10920,N_10061,N_10107);
and U10921 (N_10921,N_9927,N_10140);
nor U10922 (N_10922,N_9967,N_9667);
xor U10923 (N_10923,N_10398,N_10251);
and U10924 (N_10924,N_9832,N_10050);
nand U10925 (N_10925,N_10240,N_9955);
and U10926 (N_10926,N_10314,N_9996);
or U10927 (N_10927,N_10238,N_10285);
and U10928 (N_10928,N_10206,N_9918);
and U10929 (N_10929,N_9756,N_10213);
or U10930 (N_10930,N_10369,N_9929);
nand U10931 (N_10931,N_9847,N_9764);
or U10932 (N_10932,N_9600,N_10372);
or U10933 (N_10933,N_10244,N_9794);
nand U10934 (N_10934,N_9624,N_10358);
and U10935 (N_10935,N_9603,N_9968);
nor U10936 (N_10936,N_10305,N_10226);
or U10937 (N_10937,N_10274,N_9854);
nand U10938 (N_10938,N_9754,N_10197);
and U10939 (N_10939,N_10221,N_10052);
or U10940 (N_10940,N_9982,N_10391);
and U10941 (N_10941,N_9668,N_9619);
nor U10942 (N_10942,N_9885,N_10339);
nand U10943 (N_10943,N_10121,N_9606);
nor U10944 (N_10944,N_10386,N_9802);
xnor U10945 (N_10945,N_9966,N_9807);
and U10946 (N_10946,N_9615,N_10044);
or U10947 (N_10947,N_10250,N_10016);
nor U10948 (N_10948,N_10297,N_9885);
or U10949 (N_10949,N_10293,N_9617);
and U10950 (N_10950,N_10041,N_10057);
xor U10951 (N_10951,N_9752,N_9672);
and U10952 (N_10952,N_10361,N_9681);
and U10953 (N_10953,N_10334,N_10277);
nor U10954 (N_10954,N_10029,N_10368);
nor U10955 (N_10955,N_10183,N_10339);
nand U10956 (N_10956,N_9872,N_10146);
xor U10957 (N_10957,N_10383,N_10113);
nor U10958 (N_10958,N_9927,N_9618);
or U10959 (N_10959,N_10117,N_10207);
xnor U10960 (N_10960,N_10320,N_9632);
nor U10961 (N_10961,N_10214,N_9665);
or U10962 (N_10962,N_9700,N_9824);
and U10963 (N_10963,N_10367,N_10073);
nor U10964 (N_10964,N_9718,N_9607);
nand U10965 (N_10965,N_10143,N_10276);
or U10966 (N_10966,N_9847,N_10350);
xnor U10967 (N_10967,N_10016,N_10285);
nor U10968 (N_10968,N_9659,N_10120);
and U10969 (N_10969,N_10125,N_9646);
xnor U10970 (N_10970,N_9813,N_9847);
nand U10971 (N_10971,N_9853,N_9637);
or U10972 (N_10972,N_9719,N_9819);
nand U10973 (N_10973,N_10226,N_10079);
nand U10974 (N_10974,N_9945,N_9604);
or U10975 (N_10975,N_9813,N_9610);
and U10976 (N_10976,N_9655,N_10287);
or U10977 (N_10977,N_10275,N_9763);
xnor U10978 (N_10978,N_9965,N_9871);
or U10979 (N_10979,N_10382,N_10049);
or U10980 (N_10980,N_9875,N_9607);
or U10981 (N_10981,N_9714,N_9852);
or U10982 (N_10982,N_10309,N_10050);
nor U10983 (N_10983,N_10210,N_10395);
xnor U10984 (N_10984,N_9739,N_10023);
nand U10985 (N_10985,N_10228,N_10229);
nand U10986 (N_10986,N_10326,N_9982);
nand U10987 (N_10987,N_10354,N_10119);
or U10988 (N_10988,N_9744,N_9914);
nand U10989 (N_10989,N_9731,N_10189);
or U10990 (N_10990,N_9965,N_9906);
nor U10991 (N_10991,N_9628,N_9788);
nor U10992 (N_10992,N_9828,N_9800);
nor U10993 (N_10993,N_10255,N_9644);
nor U10994 (N_10994,N_10399,N_9815);
or U10995 (N_10995,N_9603,N_9610);
nor U10996 (N_10996,N_9789,N_10002);
nand U10997 (N_10997,N_10232,N_10211);
nor U10998 (N_10998,N_9779,N_10017);
nor U10999 (N_10999,N_9807,N_10152);
nor U11000 (N_11000,N_10120,N_10277);
or U11001 (N_11001,N_10259,N_10396);
nor U11002 (N_11002,N_9635,N_9812);
xor U11003 (N_11003,N_10153,N_10276);
and U11004 (N_11004,N_9954,N_9978);
or U11005 (N_11005,N_10360,N_9895);
nor U11006 (N_11006,N_10374,N_9993);
xnor U11007 (N_11007,N_9658,N_10064);
nor U11008 (N_11008,N_10057,N_10258);
or U11009 (N_11009,N_9614,N_10281);
xnor U11010 (N_11010,N_9984,N_9606);
nor U11011 (N_11011,N_10323,N_10273);
nand U11012 (N_11012,N_9677,N_10080);
or U11013 (N_11013,N_9610,N_9942);
nand U11014 (N_11014,N_10388,N_9635);
xnor U11015 (N_11015,N_10304,N_9872);
xnor U11016 (N_11016,N_10008,N_9677);
nand U11017 (N_11017,N_10057,N_10018);
nand U11018 (N_11018,N_9795,N_9938);
nor U11019 (N_11019,N_9712,N_10326);
and U11020 (N_11020,N_10332,N_9763);
and U11021 (N_11021,N_9870,N_9711);
xnor U11022 (N_11022,N_10101,N_9657);
and U11023 (N_11023,N_10118,N_9736);
nor U11024 (N_11024,N_10191,N_9705);
and U11025 (N_11025,N_10342,N_9651);
or U11026 (N_11026,N_9744,N_10373);
nor U11027 (N_11027,N_9808,N_9983);
nand U11028 (N_11028,N_10025,N_9781);
nor U11029 (N_11029,N_9968,N_9839);
nor U11030 (N_11030,N_10390,N_9828);
or U11031 (N_11031,N_9705,N_9650);
xnor U11032 (N_11032,N_9801,N_9895);
nand U11033 (N_11033,N_10350,N_9677);
nor U11034 (N_11034,N_9709,N_10257);
and U11035 (N_11035,N_10235,N_9791);
or U11036 (N_11036,N_10269,N_10304);
nand U11037 (N_11037,N_10081,N_10354);
nand U11038 (N_11038,N_10129,N_9841);
and U11039 (N_11039,N_9784,N_9815);
nand U11040 (N_11040,N_9753,N_10029);
or U11041 (N_11041,N_10384,N_10291);
and U11042 (N_11042,N_9776,N_10398);
nand U11043 (N_11043,N_10133,N_10108);
or U11044 (N_11044,N_10177,N_10061);
or U11045 (N_11045,N_9922,N_9736);
nand U11046 (N_11046,N_9705,N_10045);
or U11047 (N_11047,N_10139,N_10318);
and U11048 (N_11048,N_10171,N_10192);
nand U11049 (N_11049,N_10395,N_10086);
or U11050 (N_11050,N_9983,N_10066);
or U11051 (N_11051,N_10128,N_10250);
xor U11052 (N_11052,N_10023,N_10228);
or U11053 (N_11053,N_9731,N_9878);
or U11054 (N_11054,N_9603,N_10043);
nor U11055 (N_11055,N_9771,N_10016);
xnor U11056 (N_11056,N_9741,N_10235);
and U11057 (N_11057,N_10391,N_10371);
or U11058 (N_11058,N_9993,N_10135);
nand U11059 (N_11059,N_9892,N_10294);
xor U11060 (N_11060,N_10144,N_10326);
or U11061 (N_11061,N_9619,N_9733);
nand U11062 (N_11062,N_10350,N_9814);
nor U11063 (N_11063,N_9762,N_9697);
nand U11064 (N_11064,N_9753,N_10059);
nand U11065 (N_11065,N_9654,N_10287);
xnor U11066 (N_11066,N_9940,N_9788);
xnor U11067 (N_11067,N_10245,N_10007);
xor U11068 (N_11068,N_9680,N_10288);
xor U11069 (N_11069,N_10136,N_9827);
and U11070 (N_11070,N_10302,N_9734);
nor U11071 (N_11071,N_9957,N_9811);
nor U11072 (N_11072,N_10055,N_10342);
nor U11073 (N_11073,N_10236,N_10353);
nor U11074 (N_11074,N_9887,N_10047);
or U11075 (N_11075,N_10308,N_9956);
xor U11076 (N_11076,N_10274,N_9850);
and U11077 (N_11077,N_10385,N_9925);
nand U11078 (N_11078,N_10189,N_10374);
and U11079 (N_11079,N_10367,N_9753);
or U11080 (N_11080,N_10140,N_10253);
or U11081 (N_11081,N_10255,N_10279);
xor U11082 (N_11082,N_9622,N_10278);
nor U11083 (N_11083,N_9833,N_10352);
xnor U11084 (N_11084,N_10294,N_9935);
and U11085 (N_11085,N_10352,N_10199);
nand U11086 (N_11086,N_10144,N_10143);
nand U11087 (N_11087,N_9999,N_9739);
nor U11088 (N_11088,N_10132,N_10172);
and U11089 (N_11089,N_10104,N_9787);
nand U11090 (N_11090,N_10087,N_10036);
xor U11091 (N_11091,N_9789,N_9908);
xnor U11092 (N_11092,N_10331,N_10237);
or U11093 (N_11093,N_10061,N_9865);
nor U11094 (N_11094,N_10376,N_9958);
nor U11095 (N_11095,N_10324,N_9755);
nor U11096 (N_11096,N_9865,N_9798);
or U11097 (N_11097,N_10021,N_10060);
nor U11098 (N_11098,N_9739,N_10285);
nor U11099 (N_11099,N_10010,N_9650);
nand U11100 (N_11100,N_9764,N_10322);
xor U11101 (N_11101,N_9711,N_10005);
xnor U11102 (N_11102,N_10073,N_10273);
or U11103 (N_11103,N_10337,N_10155);
or U11104 (N_11104,N_9763,N_10310);
xnor U11105 (N_11105,N_9901,N_9791);
nand U11106 (N_11106,N_9945,N_9792);
and U11107 (N_11107,N_10065,N_9857);
nand U11108 (N_11108,N_10283,N_9822);
nand U11109 (N_11109,N_9950,N_9744);
nor U11110 (N_11110,N_10147,N_10228);
xor U11111 (N_11111,N_9709,N_9926);
nor U11112 (N_11112,N_9916,N_10018);
nand U11113 (N_11113,N_10052,N_10007);
nor U11114 (N_11114,N_9889,N_9897);
and U11115 (N_11115,N_9647,N_9621);
or U11116 (N_11116,N_9760,N_9654);
and U11117 (N_11117,N_10228,N_10389);
or U11118 (N_11118,N_9937,N_10098);
nor U11119 (N_11119,N_9749,N_10072);
xnor U11120 (N_11120,N_9780,N_10199);
xnor U11121 (N_11121,N_10217,N_10248);
nand U11122 (N_11122,N_9775,N_9980);
xnor U11123 (N_11123,N_9962,N_9741);
or U11124 (N_11124,N_9664,N_10166);
xnor U11125 (N_11125,N_10373,N_9979);
or U11126 (N_11126,N_10235,N_10317);
xnor U11127 (N_11127,N_9991,N_10334);
nand U11128 (N_11128,N_9814,N_10333);
nor U11129 (N_11129,N_10072,N_9768);
nand U11130 (N_11130,N_10221,N_9734);
nor U11131 (N_11131,N_9778,N_9748);
xnor U11132 (N_11132,N_9674,N_10148);
nand U11133 (N_11133,N_9714,N_9651);
and U11134 (N_11134,N_9746,N_9818);
xor U11135 (N_11135,N_9663,N_10155);
and U11136 (N_11136,N_9788,N_10280);
and U11137 (N_11137,N_9669,N_10341);
or U11138 (N_11138,N_9818,N_9692);
or U11139 (N_11139,N_10025,N_10080);
nor U11140 (N_11140,N_10368,N_10206);
xor U11141 (N_11141,N_9891,N_9930);
or U11142 (N_11142,N_10098,N_10120);
nor U11143 (N_11143,N_9955,N_9976);
xor U11144 (N_11144,N_10102,N_9828);
xnor U11145 (N_11145,N_9783,N_10210);
and U11146 (N_11146,N_9608,N_10001);
xor U11147 (N_11147,N_10158,N_10295);
and U11148 (N_11148,N_9704,N_10313);
or U11149 (N_11149,N_9746,N_10227);
nor U11150 (N_11150,N_10149,N_10111);
and U11151 (N_11151,N_9769,N_10079);
nor U11152 (N_11152,N_9791,N_9685);
nor U11153 (N_11153,N_10093,N_9867);
and U11154 (N_11154,N_9731,N_10152);
xnor U11155 (N_11155,N_10259,N_9705);
xnor U11156 (N_11156,N_10106,N_10107);
xor U11157 (N_11157,N_9654,N_9852);
nor U11158 (N_11158,N_9859,N_10307);
nor U11159 (N_11159,N_10391,N_9752);
or U11160 (N_11160,N_9865,N_10121);
xnor U11161 (N_11161,N_9653,N_9839);
nand U11162 (N_11162,N_9926,N_9850);
and U11163 (N_11163,N_9862,N_9898);
and U11164 (N_11164,N_10018,N_10311);
or U11165 (N_11165,N_10185,N_10292);
xnor U11166 (N_11166,N_10267,N_9616);
or U11167 (N_11167,N_10293,N_10361);
and U11168 (N_11168,N_9730,N_9726);
nor U11169 (N_11169,N_10242,N_9977);
and U11170 (N_11170,N_10218,N_10321);
nor U11171 (N_11171,N_9997,N_10054);
and U11172 (N_11172,N_9879,N_9866);
or U11173 (N_11173,N_10289,N_10379);
and U11174 (N_11174,N_9927,N_9806);
or U11175 (N_11175,N_10004,N_9954);
nand U11176 (N_11176,N_9870,N_10001);
or U11177 (N_11177,N_9876,N_10153);
or U11178 (N_11178,N_10051,N_9617);
or U11179 (N_11179,N_9900,N_9632);
or U11180 (N_11180,N_10294,N_10276);
nand U11181 (N_11181,N_10217,N_10307);
nand U11182 (N_11182,N_9651,N_9858);
nor U11183 (N_11183,N_10063,N_9613);
or U11184 (N_11184,N_9757,N_9721);
and U11185 (N_11185,N_9644,N_9826);
nor U11186 (N_11186,N_9863,N_10102);
nand U11187 (N_11187,N_10339,N_9976);
and U11188 (N_11188,N_10297,N_9690);
nand U11189 (N_11189,N_10379,N_9636);
nand U11190 (N_11190,N_9614,N_10153);
and U11191 (N_11191,N_9891,N_10190);
and U11192 (N_11192,N_10147,N_9978);
xnor U11193 (N_11193,N_9764,N_9952);
xnor U11194 (N_11194,N_9924,N_9973);
and U11195 (N_11195,N_9992,N_9600);
nand U11196 (N_11196,N_10330,N_10175);
or U11197 (N_11197,N_9819,N_10087);
nor U11198 (N_11198,N_10218,N_10308);
nor U11199 (N_11199,N_9740,N_10268);
nand U11200 (N_11200,N_10549,N_10908);
nor U11201 (N_11201,N_10761,N_10779);
or U11202 (N_11202,N_10925,N_10659);
xnor U11203 (N_11203,N_11087,N_10976);
and U11204 (N_11204,N_11055,N_11089);
nand U11205 (N_11205,N_11173,N_10461);
nor U11206 (N_11206,N_10489,N_10810);
or U11207 (N_11207,N_10467,N_11106);
xnor U11208 (N_11208,N_10463,N_11133);
or U11209 (N_11209,N_10838,N_10726);
or U11210 (N_11210,N_11049,N_10930);
nor U11211 (N_11211,N_11141,N_10451);
nor U11212 (N_11212,N_11154,N_10892);
and U11213 (N_11213,N_10718,N_10952);
xnor U11214 (N_11214,N_10992,N_10860);
xnor U11215 (N_11215,N_10437,N_10427);
xnor U11216 (N_11216,N_10788,N_11018);
nand U11217 (N_11217,N_10864,N_10614);
nand U11218 (N_11218,N_11083,N_10510);
nand U11219 (N_11219,N_10604,N_11136);
xor U11220 (N_11220,N_10502,N_10826);
nand U11221 (N_11221,N_11109,N_10770);
nand U11222 (N_11222,N_10784,N_10883);
or U11223 (N_11223,N_10571,N_10420);
and U11224 (N_11224,N_10792,N_11027);
xor U11225 (N_11225,N_11071,N_10492);
nand U11226 (N_11226,N_11054,N_11004);
or U11227 (N_11227,N_10818,N_11131);
nand U11228 (N_11228,N_10589,N_11061);
nand U11229 (N_11229,N_10532,N_10528);
nor U11230 (N_11230,N_11093,N_10503);
nor U11231 (N_11231,N_10591,N_10416);
or U11232 (N_11232,N_10945,N_10763);
nand U11233 (N_11233,N_11091,N_10939);
nand U11234 (N_11234,N_10547,N_10491);
xor U11235 (N_11235,N_10505,N_11129);
or U11236 (N_11236,N_10683,N_10853);
nor U11237 (N_11237,N_10628,N_10795);
and U11238 (N_11238,N_10508,N_10612);
xor U11239 (N_11239,N_10641,N_11074);
nor U11240 (N_11240,N_10872,N_11188);
nor U11241 (N_11241,N_11149,N_10756);
xnor U11242 (N_11242,N_10432,N_10671);
xnor U11243 (N_11243,N_11166,N_10592);
xnor U11244 (N_11244,N_11104,N_10704);
nor U11245 (N_11245,N_10520,N_10941);
nor U11246 (N_11246,N_10744,N_10724);
xor U11247 (N_11247,N_10819,N_10972);
nor U11248 (N_11248,N_10686,N_10710);
or U11249 (N_11249,N_10550,N_10652);
nor U11250 (N_11250,N_10938,N_10760);
or U11251 (N_11251,N_10982,N_10450);
and U11252 (N_11252,N_10643,N_10880);
nand U11253 (N_11253,N_11044,N_10858);
xor U11254 (N_11254,N_10986,N_10736);
or U11255 (N_11255,N_10924,N_10702);
nor U11256 (N_11256,N_10906,N_10768);
or U11257 (N_11257,N_10501,N_11148);
nor U11258 (N_11258,N_10757,N_10919);
xor U11259 (N_11259,N_10431,N_10595);
nand U11260 (N_11260,N_10722,N_10603);
nand U11261 (N_11261,N_10854,N_11099);
xor U11262 (N_11262,N_10961,N_11058);
nand U11263 (N_11263,N_10588,N_11028);
nand U11264 (N_11264,N_11130,N_10587);
nand U11265 (N_11265,N_10645,N_10633);
nor U11266 (N_11266,N_10500,N_10511);
and U11267 (N_11267,N_10829,N_10994);
or U11268 (N_11268,N_10566,N_10968);
or U11269 (N_11269,N_11017,N_10476);
nor U11270 (N_11270,N_10447,N_10861);
and U11271 (N_11271,N_10676,N_10749);
xor U11272 (N_11272,N_11118,N_10949);
nor U11273 (N_11273,N_10727,N_10490);
nand U11274 (N_11274,N_10609,N_10765);
and U11275 (N_11275,N_10890,N_10552);
nor U11276 (N_11276,N_10443,N_10921);
nand U11277 (N_11277,N_10781,N_10617);
or U11278 (N_11278,N_10891,N_10421);
nand U11279 (N_11279,N_10873,N_10980);
xor U11280 (N_11280,N_11177,N_10742);
xor U11281 (N_11281,N_11035,N_10651);
xor U11282 (N_11282,N_10855,N_10869);
xnor U11283 (N_11283,N_10573,N_11047);
xor U11284 (N_11284,N_10464,N_10579);
or U11285 (N_11285,N_10808,N_10750);
xnor U11286 (N_11286,N_10732,N_11075);
or U11287 (N_11287,N_10964,N_10600);
xor U11288 (N_11288,N_10851,N_10907);
and U11289 (N_11289,N_10835,N_10663);
xor U11290 (N_11290,N_10755,N_10885);
and U11291 (N_11291,N_10745,N_10785);
or U11292 (N_11292,N_10905,N_10739);
or U11293 (N_11293,N_10405,N_11060);
and U11294 (N_11294,N_11165,N_10418);
and U11295 (N_11295,N_10478,N_10911);
nand U11296 (N_11296,N_10606,N_10965);
and U11297 (N_11297,N_10556,N_10767);
nand U11298 (N_11298,N_10916,N_11011);
nand U11299 (N_11299,N_10404,N_10996);
or U11300 (N_11300,N_10735,N_10632);
nor U11301 (N_11301,N_10967,N_11102);
nor U11302 (N_11302,N_10626,N_10569);
nand U11303 (N_11303,N_10894,N_10498);
nor U11304 (N_11304,N_11142,N_10553);
nand U11305 (N_11305,N_10936,N_10586);
xor U11306 (N_11306,N_10811,N_11006);
and U11307 (N_11307,N_11101,N_11079);
and U11308 (N_11308,N_10828,N_10960);
nor U11309 (N_11309,N_10773,N_10910);
nor U11310 (N_11310,N_11000,N_11037);
xnor U11311 (N_11311,N_11114,N_10513);
xnor U11312 (N_11312,N_11170,N_11103);
or U11313 (N_11313,N_11191,N_11120);
and U11314 (N_11314,N_10474,N_10769);
or U11315 (N_11315,N_10630,N_10809);
xor U11316 (N_11316,N_11072,N_10725);
or U11317 (N_11317,N_10407,N_11023);
nor U11318 (N_11318,N_10954,N_10422);
nor U11319 (N_11319,N_10413,N_10687);
nand U11320 (N_11320,N_10530,N_10867);
or U11321 (N_11321,N_10608,N_10680);
nor U11322 (N_11322,N_11157,N_11124);
nand U11323 (N_11323,N_10578,N_10408);
xor U11324 (N_11324,N_10636,N_11171);
and U11325 (N_11325,N_10805,N_10665);
and U11326 (N_11326,N_10682,N_10694);
xnor U11327 (N_11327,N_10902,N_10555);
nor U11328 (N_11328,N_10497,N_10793);
or U11329 (N_11329,N_10615,N_11150);
or U11330 (N_11330,N_10804,N_10777);
and U11331 (N_11331,N_10874,N_10535);
or U11332 (N_11332,N_11098,N_11179);
nand U11333 (N_11333,N_10570,N_11151);
and U11334 (N_11334,N_11056,N_11084);
or U11335 (N_11335,N_10841,N_10973);
or U11336 (N_11336,N_11122,N_10542);
and U11337 (N_11337,N_10951,N_10944);
nor U11338 (N_11338,N_10563,N_10822);
nand U11339 (N_11339,N_10425,N_10806);
xnor U11340 (N_11340,N_10700,N_10649);
nand U11341 (N_11341,N_10582,N_10848);
and U11342 (N_11342,N_10488,N_10657);
and U11343 (N_11343,N_10823,N_11010);
nand U11344 (N_11344,N_10584,N_10844);
or U11345 (N_11345,N_10813,N_10993);
and U11346 (N_11346,N_10743,N_10758);
nor U11347 (N_11347,N_10449,N_10714);
xnor U11348 (N_11348,N_10875,N_10529);
and U11349 (N_11349,N_10560,N_10821);
or U11350 (N_11350,N_10803,N_11070);
nor U11351 (N_11351,N_10983,N_10509);
nand U11352 (N_11352,N_10526,N_10729);
nand U11353 (N_11353,N_10624,N_11155);
xnor U11354 (N_11354,N_10877,N_10523);
nor U11355 (N_11355,N_11192,N_10791);
xor U11356 (N_11356,N_11057,N_10562);
and U11357 (N_11357,N_10507,N_11126);
xnor U11358 (N_11358,N_10666,N_10977);
or U11359 (N_11359,N_10470,N_10898);
nand U11360 (N_11360,N_10981,N_10471);
or U11361 (N_11361,N_10780,N_11042);
and U11362 (N_11362,N_10575,N_11117);
nand U11363 (N_11363,N_11040,N_10538);
xnor U11364 (N_11364,N_10667,N_10524);
or U11365 (N_11365,N_10479,N_10688);
nand U11366 (N_11366,N_11045,N_10846);
nand U11367 (N_11367,N_11076,N_10863);
or U11368 (N_11368,N_11196,N_10602);
or U11369 (N_11369,N_10912,N_10441);
nand U11370 (N_11370,N_10879,N_10857);
nor U11371 (N_11371,N_11147,N_10436);
xor U11372 (N_11372,N_10419,N_11167);
nor U11373 (N_11373,N_10859,N_11145);
nand U11374 (N_11374,N_11041,N_10827);
nor U11375 (N_11375,N_10889,N_11100);
and U11376 (N_11376,N_10786,N_10856);
or U11377 (N_11377,N_11143,N_10928);
nor U11378 (N_11378,N_10955,N_10519);
or U11379 (N_11379,N_10896,N_10620);
or U11380 (N_11380,N_10782,N_10653);
nor U11381 (N_11381,N_11024,N_10915);
xnor U11382 (N_11382,N_11080,N_10929);
or U11383 (N_11383,N_10635,N_10650);
nand U11384 (N_11384,N_11088,N_10454);
nor U11385 (N_11385,N_11163,N_10927);
or U11386 (N_11386,N_10695,N_10494);
xnor U11387 (N_11387,N_10473,N_10920);
or U11388 (N_11388,N_11134,N_10868);
xor U11389 (N_11389,N_10815,N_10487);
nor U11390 (N_11390,N_11046,N_10544);
nor U11391 (N_11391,N_11043,N_10581);
nand U11392 (N_11392,N_10751,N_11097);
nor U11393 (N_11393,N_10878,N_10747);
nor U11394 (N_11394,N_10692,N_11199);
and U11395 (N_11395,N_10833,N_10577);
and U11396 (N_11396,N_10886,N_10715);
or U11397 (N_11397,N_11069,N_10409);
and U11398 (N_11398,N_10995,N_10506);
nor U11399 (N_11399,N_10631,N_10897);
or U11400 (N_11400,N_10400,N_10537);
and U11401 (N_11401,N_11197,N_10654);
and U11402 (N_11402,N_11195,N_11032);
or U11403 (N_11403,N_10895,N_11025);
nor U11404 (N_11404,N_10825,N_10871);
or U11405 (N_11405,N_10596,N_10406);
nor U11406 (N_11406,N_10677,N_10623);
and U11407 (N_11407,N_10966,N_11115);
or U11408 (N_11408,N_10551,N_10881);
nand U11409 (N_11409,N_10696,N_11002);
xnor U11410 (N_11410,N_11036,N_10574);
nor U11411 (N_11411,N_10884,N_10797);
xnor U11412 (N_11412,N_11059,N_10459);
nand U11413 (N_11413,N_10598,N_10482);
or U11414 (N_11414,N_11034,N_11014);
xor U11415 (N_11415,N_10799,N_10716);
xnor U11416 (N_11416,N_11020,N_10963);
nor U11417 (N_11417,N_10947,N_10787);
nor U11418 (N_11418,N_11053,N_10618);
nand U11419 (N_11419,N_10764,N_10918);
nand U11420 (N_11420,N_11105,N_10644);
xnor U11421 (N_11421,N_10723,N_11193);
xor U11422 (N_11422,N_10728,N_10539);
nand U11423 (N_11423,N_10439,N_10748);
or U11424 (N_11424,N_10801,N_11113);
or U11425 (N_11425,N_10621,N_10655);
and U11426 (N_11426,N_10658,N_11095);
or U11427 (N_11427,N_10824,N_10440);
xnor U11428 (N_11428,N_10417,N_10517);
nand U11429 (N_11429,N_11050,N_10412);
nand U11430 (N_11430,N_10990,N_10865);
nand U11431 (N_11431,N_10568,N_11162);
xnor U11432 (N_11432,N_10888,N_10933);
xor U11433 (N_11433,N_10627,N_10985);
xnor U11434 (N_11434,N_10625,N_10935);
nor U11435 (N_11435,N_11082,N_11063);
nor U11436 (N_11436,N_10814,N_10672);
nand U11437 (N_11437,N_10931,N_10903);
nor U11438 (N_11438,N_10932,N_10675);
and U11439 (N_11439,N_10446,N_11138);
nor U11440 (N_11440,N_11068,N_10734);
and U11441 (N_11441,N_10975,N_11039);
and U11442 (N_11442,N_10946,N_10882);
nand U11443 (N_11443,N_11013,N_11185);
and U11444 (N_11444,N_10738,N_10515);
nand U11445 (N_11445,N_10411,N_10789);
xnor U11446 (N_11446,N_10557,N_10776);
xnor U11447 (N_11447,N_11096,N_10428);
and U11448 (N_11448,N_11190,N_10594);
xor U11449 (N_11449,N_10564,N_10711);
nor U11450 (N_11450,N_10540,N_10546);
nand U11451 (N_11451,N_10599,N_10434);
nor U11452 (N_11452,N_11137,N_10640);
or U11453 (N_11453,N_10590,N_10998);
nor U11454 (N_11454,N_10458,N_11033);
and U11455 (N_11455,N_11094,N_10812);
nand U11456 (N_11456,N_10698,N_11176);
nand U11457 (N_11457,N_11183,N_10634);
and U11458 (N_11458,N_10759,N_11132);
or U11459 (N_11459,N_10518,N_10469);
and U11460 (N_11460,N_10610,N_10834);
nand U11461 (N_11461,N_11153,N_10934);
nand U11462 (N_11462,N_10798,N_10772);
nand U11463 (N_11463,N_10962,N_11086);
nor U11464 (N_11464,N_10455,N_10438);
xnor U11465 (N_11465,N_10703,N_11194);
nor U11466 (N_11466,N_10558,N_10691);
and U11467 (N_11467,N_10597,N_10401);
nor U11468 (N_11468,N_11123,N_10984);
and U11469 (N_11469,N_10456,N_10836);
nand U11470 (N_11470,N_10426,N_11015);
and U11471 (N_11471,N_11112,N_10585);
nor U11472 (N_11472,N_11172,N_10712);
xnor U11473 (N_11473,N_10430,N_10746);
nor U11474 (N_11474,N_10790,N_11186);
or U11475 (N_11475,N_10820,N_10926);
xor U11476 (N_11476,N_10685,N_10678);
nor U11477 (N_11477,N_11077,N_11139);
xnor U11478 (N_11478,N_10561,N_11108);
xor U11479 (N_11479,N_10521,N_10567);
nor U11480 (N_11480,N_10796,N_10783);
nand U11481 (N_11481,N_10847,N_10771);
xor U11482 (N_11482,N_10840,N_10737);
xor U11483 (N_11483,N_11189,N_10495);
and U11484 (N_11484,N_10646,N_10648);
xnor U11485 (N_11485,N_11164,N_10415);
nor U11486 (N_11486,N_11016,N_11169);
nor U11487 (N_11487,N_11073,N_10534);
nor U11488 (N_11488,N_10713,N_10849);
nor U11489 (N_11489,N_10802,N_10904);
and U11490 (N_11490,N_10842,N_11140);
and U11491 (N_11491,N_10572,N_11062);
and U11492 (N_11492,N_10991,N_10429);
and U11493 (N_11493,N_10611,N_10622);
xor U11494 (N_11494,N_10778,N_10901);
nor U11495 (N_11495,N_10457,N_10942);
or U11496 (N_11496,N_10762,N_11135);
nor U11497 (N_11497,N_10580,N_10970);
nor U11498 (N_11498,N_10839,N_11066);
or U11499 (N_11499,N_11160,N_10527);
nor U11500 (N_11500,N_10484,N_10870);
xnor U11501 (N_11501,N_10923,N_11107);
nand U11502 (N_11502,N_11003,N_10832);
nor U11503 (N_11503,N_11156,N_11001);
or U11504 (N_11504,N_10472,N_10496);
or U11505 (N_11505,N_10775,N_11127);
and U11506 (N_11506,N_11110,N_10673);
nand U11507 (N_11507,N_10485,N_10697);
nor U11508 (N_11508,N_10403,N_10499);
or U11509 (N_11509,N_10493,N_11009);
xnor U11510 (N_11510,N_10721,N_11022);
or U11511 (N_11511,N_10477,N_10629);
nor U11512 (N_11512,N_10706,N_10483);
nor U11513 (N_11513,N_10554,N_10843);
or U11514 (N_11514,N_10674,N_10731);
nor U11515 (N_11515,N_10800,N_11178);
nor U11516 (N_11516,N_10708,N_11081);
nor U11517 (N_11517,N_10900,N_11026);
or U11518 (N_11518,N_11198,N_10979);
nand U11519 (N_11519,N_10670,N_11019);
xnor U11520 (N_11520,N_10943,N_10619);
nand U11521 (N_11521,N_10679,N_10444);
nand U11522 (N_11522,N_10605,N_10956);
nand U11523 (N_11523,N_10950,N_10435);
xnor U11524 (N_11524,N_10794,N_10922);
and U11525 (N_11525,N_10937,N_10424);
nor U11526 (N_11526,N_10565,N_10548);
xnor U11527 (N_11527,N_10753,N_11128);
or U11528 (N_11528,N_10637,N_10699);
or U11529 (N_11529,N_11090,N_10452);
nand U11530 (N_11530,N_10453,N_10583);
xnor U11531 (N_11531,N_11161,N_11065);
xor U11532 (N_11532,N_10607,N_10720);
and U11533 (N_11533,N_10638,N_11030);
nor U11534 (N_11534,N_10642,N_10774);
nor U11535 (N_11535,N_10514,N_11187);
nor U11536 (N_11536,N_10766,N_10817);
xor U11537 (N_11537,N_11078,N_11182);
nand U11538 (N_11538,N_10465,N_10730);
nand U11539 (N_11539,N_10543,N_10958);
xnor U11540 (N_11540,N_10536,N_10999);
nor U11541 (N_11541,N_10669,N_10689);
and U11542 (N_11542,N_10953,N_11180);
nand U11543 (N_11543,N_10664,N_10940);
xnor U11544 (N_11544,N_10987,N_10899);
nor U11545 (N_11545,N_11168,N_10959);
or U11546 (N_11546,N_11085,N_10830);
nand U11547 (N_11547,N_11005,N_10522);
or U11548 (N_11548,N_10733,N_10917);
nor U11549 (N_11549,N_11181,N_10541);
xor U11550 (N_11550,N_10576,N_11144);
nand U11551 (N_11551,N_10662,N_10852);
and U11552 (N_11552,N_10909,N_10656);
and U11553 (N_11553,N_10613,N_10462);
nor U11554 (N_11554,N_11064,N_10668);
nor U11555 (N_11555,N_10831,N_10516);
xor U11556 (N_11556,N_10971,N_10410);
or U11557 (N_11557,N_11092,N_10647);
nand U11558 (N_11558,N_10402,N_10693);
or U11559 (N_11559,N_10709,N_10887);
or U11560 (N_11560,N_10601,N_11008);
and U11561 (N_11561,N_10850,N_10717);
xor U11562 (N_11562,N_10639,N_10701);
nor U11563 (N_11563,N_10754,N_10480);
and U11564 (N_11564,N_11175,N_11184);
xor U11565 (N_11565,N_10876,N_10837);
or U11566 (N_11566,N_11007,N_10974);
xnor U11567 (N_11567,N_10914,N_10414);
and U11568 (N_11568,N_10660,N_10741);
or U11569 (N_11569,N_10481,N_10988);
xnor U11570 (N_11570,N_10948,N_11038);
and U11571 (N_11571,N_10445,N_10807);
or U11572 (N_11572,N_10442,N_10423);
and U11573 (N_11573,N_10740,N_10862);
nand U11574 (N_11574,N_11121,N_11111);
nor U11575 (N_11575,N_10893,N_11116);
xor U11576 (N_11576,N_10593,N_10512);
and U11577 (N_11577,N_10866,N_11048);
nand U11578 (N_11578,N_10533,N_11152);
xor U11579 (N_11579,N_11158,N_11029);
nor U11580 (N_11580,N_10486,N_11021);
xor U11581 (N_11581,N_10989,N_10448);
and U11582 (N_11582,N_10468,N_10681);
and U11583 (N_11583,N_10957,N_10719);
nand U11584 (N_11584,N_11146,N_10816);
and U11585 (N_11585,N_10997,N_11012);
and U11586 (N_11586,N_10616,N_10545);
and U11587 (N_11587,N_10752,N_11119);
nand U11588 (N_11588,N_10433,N_10705);
or U11589 (N_11589,N_10504,N_10690);
xor U11590 (N_11590,N_10460,N_11051);
nand U11591 (N_11591,N_10707,N_11174);
nor U11592 (N_11592,N_10845,N_10913);
nor U11593 (N_11593,N_10475,N_10684);
nand U11594 (N_11594,N_11052,N_10559);
nand U11595 (N_11595,N_11125,N_10531);
nor U11596 (N_11596,N_11159,N_10466);
nor U11597 (N_11597,N_10525,N_10978);
xnor U11598 (N_11598,N_11067,N_10969);
or U11599 (N_11599,N_11031,N_10661);
or U11600 (N_11600,N_10632,N_10641);
xnor U11601 (N_11601,N_11077,N_10430);
and U11602 (N_11602,N_10545,N_10544);
nand U11603 (N_11603,N_11119,N_10951);
xor U11604 (N_11604,N_10438,N_10901);
nand U11605 (N_11605,N_11085,N_10531);
xor U11606 (N_11606,N_10471,N_10863);
and U11607 (N_11607,N_10998,N_11099);
or U11608 (N_11608,N_11066,N_10835);
xnor U11609 (N_11609,N_10459,N_10508);
xor U11610 (N_11610,N_10410,N_10870);
nor U11611 (N_11611,N_10567,N_10638);
and U11612 (N_11612,N_10462,N_11146);
nor U11613 (N_11613,N_10915,N_10662);
and U11614 (N_11614,N_10741,N_10585);
nand U11615 (N_11615,N_11047,N_10743);
or U11616 (N_11616,N_10749,N_10514);
and U11617 (N_11617,N_10483,N_10865);
and U11618 (N_11618,N_10942,N_10754);
xnor U11619 (N_11619,N_10870,N_10673);
nor U11620 (N_11620,N_10712,N_10588);
xor U11621 (N_11621,N_10528,N_11008);
nand U11622 (N_11622,N_10528,N_11130);
nor U11623 (N_11623,N_11136,N_10607);
nand U11624 (N_11624,N_10408,N_10411);
xor U11625 (N_11625,N_10973,N_10988);
nand U11626 (N_11626,N_10783,N_10692);
and U11627 (N_11627,N_11147,N_11073);
xnor U11628 (N_11628,N_10590,N_10572);
and U11629 (N_11629,N_10644,N_10604);
nor U11630 (N_11630,N_10675,N_10956);
and U11631 (N_11631,N_10433,N_10895);
or U11632 (N_11632,N_11155,N_10530);
xnor U11633 (N_11633,N_10483,N_11023);
and U11634 (N_11634,N_10644,N_11019);
xnor U11635 (N_11635,N_10464,N_10998);
and U11636 (N_11636,N_10924,N_11024);
nor U11637 (N_11637,N_10400,N_10694);
and U11638 (N_11638,N_10885,N_10429);
nor U11639 (N_11639,N_10721,N_10593);
nor U11640 (N_11640,N_10536,N_10499);
nor U11641 (N_11641,N_10420,N_10448);
nor U11642 (N_11642,N_10726,N_10944);
xor U11643 (N_11643,N_10574,N_11157);
and U11644 (N_11644,N_10453,N_10672);
and U11645 (N_11645,N_11152,N_10430);
and U11646 (N_11646,N_11069,N_11132);
nand U11647 (N_11647,N_10752,N_10883);
nand U11648 (N_11648,N_10738,N_10502);
or U11649 (N_11649,N_10892,N_10829);
nand U11650 (N_11650,N_10945,N_10996);
nand U11651 (N_11651,N_10550,N_10538);
nor U11652 (N_11652,N_10815,N_10590);
xor U11653 (N_11653,N_10600,N_10421);
nand U11654 (N_11654,N_10445,N_10698);
xnor U11655 (N_11655,N_11197,N_10592);
xnor U11656 (N_11656,N_10462,N_10692);
xnor U11657 (N_11657,N_10792,N_10679);
or U11658 (N_11658,N_10571,N_11082);
xor U11659 (N_11659,N_10886,N_10854);
xor U11660 (N_11660,N_10867,N_10950);
nor U11661 (N_11661,N_11097,N_10902);
nor U11662 (N_11662,N_11064,N_10473);
nand U11663 (N_11663,N_10429,N_10823);
xor U11664 (N_11664,N_10927,N_10816);
or U11665 (N_11665,N_10569,N_10591);
nor U11666 (N_11666,N_10839,N_10408);
and U11667 (N_11667,N_10494,N_10442);
xnor U11668 (N_11668,N_10624,N_10752);
nor U11669 (N_11669,N_11138,N_10528);
or U11670 (N_11670,N_10697,N_10512);
or U11671 (N_11671,N_10666,N_10418);
nand U11672 (N_11672,N_10515,N_10536);
or U11673 (N_11673,N_10920,N_10583);
and U11674 (N_11674,N_10953,N_11186);
nand U11675 (N_11675,N_10964,N_11185);
xnor U11676 (N_11676,N_10646,N_10562);
nand U11677 (N_11677,N_10532,N_10747);
and U11678 (N_11678,N_10619,N_11044);
or U11679 (N_11679,N_10854,N_10689);
xor U11680 (N_11680,N_10782,N_10992);
and U11681 (N_11681,N_10804,N_10457);
or U11682 (N_11682,N_10458,N_11024);
and U11683 (N_11683,N_10878,N_11083);
nor U11684 (N_11684,N_11084,N_11109);
nor U11685 (N_11685,N_10440,N_10547);
or U11686 (N_11686,N_11041,N_10778);
nor U11687 (N_11687,N_10660,N_10988);
or U11688 (N_11688,N_10819,N_10532);
xor U11689 (N_11689,N_10525,N_10458);
or U11690 (N_11690,N_10856,N_11039);
xnor U11691 (N_11691,N_10750,N_10680);
nand U11692 (N_11692,N_10638,N_10640);
nand U11693 (N_11693,N_10443,N_11145);
and U11694 (N_11694,N_10540,N_10690);
nor U11695 (N_11695,N_10820,N_10415);
xnor U11696 (N_11696,N_10784,N_10957);
nand U11697 (N_11697,N_10842,N_11118);
nand U11698 (N_11698,N_10554,N_10715);
and U11699 (N_11699,N_10647,N_10545);
xor U11700 (N_11700,N_11117,N_10429);
xor U11701 (N_11701,N_10977,N_11184);
nor U11702 (N_11702,N_11145,N_11048);
nand U11703 (N_11703,N_10436,N_10488);
nand U11704 (N_11704,N_10410,N_10773);
nand U11705 (N_11705,N_10525,N_10645);
nand U11706 (N_11706,N_10479,N_10556);
and U11707 (N_11707,N_10819,N_10410);
xnor U11708 (N_11708,N_10539,N_10815);
xnor U11709 (N_11709,N_11018,N_11090);
nor U11710 (N_11710,N_10435,N_10529);
nor U11711 (N_11711,N_10556,N_10422);
and U11712 (N_11712,N_10913,N_11048);
nor U11713 (N_11713,N_10717,N_10991);
nor U11714 (N_11714,N_11198,N_10663);
nor U11715 (N_11715,N_10961,N_10768);
xor U11716 (N_11716,N_10451,N_11190);
or U11717 (N_11717,N_11095,N_10924);
nand U11718 (N_11718,N_10521,N_10708);
nand U11719 (N_11719,N_10993,N_11042);
and U11720 (N_11720,N_10906,N_10821);
or U11721 (N_11721,N_10737,N_10785);
and U11722 (N_11722,N_10423,N_11174);
and U11723 (N_11723,N_10851,N_10789);
and U11724 (N_11724,N_10795,N_10786);
xnor U11725 (N_11725,N_10599,N_10559);
nand U11726 (N_11726,N_10530,N_11195);
nor U11727 (N_11727,N_10420,N_10854);
xnor U11728 (N_11728,N_10501,N_10918);
nand U11729 (N_11729,N_10851,N_10575);
xor U11730 (N_11730,N_10462,N_10720);
or U11731 (N_11731,N_10733,N_10795);
nor U11732 (N_11732,N_10449,N_10826);
nor U11733 (N_11733,N_10442,N_10520);
or U11734 (N_11734,N_10650,N_11090);
xnor U11735 (N_11735,N_10958,N_10512);
nand U11736 (N_11736,N_10624,N_10625);
xor U11737 (N_11737,N_10468,N_11089);
and U11738 (N_11738,N_10503,N_10706);
or U11739 (N_11739,N_10762,N_10917);
xor U11740 (N_11740,N_10688,N_10535);
or U11741 (N_11741,N_11046,N_10837);
xnor U11742 (N_11742,N_10789,N_10506);
or U11743 (N_11743,N_10852,N_10438);
xor U11744 (N_11744,N_10775,N_10559);
and U11745 (N_11745,N_10902,N_10617);
xor U11746 (N_11746,N_10991,N_10827);
and U11747 (N_11747,N_10679,N_11198);
nand U11748 (N_11748,N_10914,N_10571);
or U11749 (N_11749,N_11102,N_11003);
or U11750 (N_11750,N_10575,N_11055);
nand U11751 (N_11751,N_10431,N_10413);
xnor U11752 (N_11752,N_10778,N_10494);
nand U11753 (N_11753,N_10603,N_10434);
and U11754 (N_11754,N_11102,N_10585);
and U11755 (N_11755,N_10634,N_10545);
or U11756 (N_11756,N_10705,N_10911);
nor U11757 (N_11757,N_10757,N_10937);
nand U11758 (N_11758,N_10721,N_10462);
and U11759 (N_11759,N_11117,N_11159);
or U11760 (N_11760,N_10992,N_10568);
nand U11761 (N_11761,N_10925,N_10634);
nor U11762 (N_11762,N_10428,N_10798);
nand U11763 (N_11763,N_10423,N_11162);
nor U11764 (N_11764,N_10728,N_10821);
nor U11765 (N_11765,N_11121,N_11042);
xor U11766 (N_11766,N_11071,N_10690);
or U11767 (N_11767,N_10497,N_10839);
or U11768 (N_11768,N_10679,N_11022);
nand U11769 (N_11769,N_11075,N_10985);
and U11770 (N_11770,N_10873,N_10740);
or U11771 (N_11771,N_10499,N_10640);
nand U11772 (N_11772,N_11038,N_10916);
xor U11773 (N_11773,N_10498,N_10824);
nor U11774 (N_11774,N_10876,N_10733);
xnor U11775 (N_11775,N_10441,N_11150);
or U11776 (N_11776,N_10612,N_10594);
xor U11777 (N_11777,N_11187,N_10909);
xor U11778 (N_11778,N_11078,N_10676);
or U11779 (N_11779,N_10751,N_10747);
nor U11780 (N_11780,N_10493,N_11024);
and U11781 (N_11781,N_10807,N_11019);
nor U11782 (N_11782,N_10964,N_11177);
and U11783 (N_11783,N_11008,N_11025);
or U11784 (N_11784,N_10463,N_10829);
nor U11785 (N_11785,N_10600,N_10694);
or U11786 (N_11786,N_10725,N_11079);
nor U11787 (N_11787,N_11147,N_11163);
nand U11788 (N_11788,N_10445,N_10705);
nand U11789 (N_11789,N_10666,N_10772);
and U11790 (N_11790,N_10808,N_10785);
xnor U11791 (N_11791,N_10910,N_10902);
and U11792 (N_11792,N_10961,N_10997);
nor U11793 (N_11793,N_10774,N_10546);
or U11794 (N_11794,N_10575,N_10457);
and U11795 (N_11795,N_10847,N_10893);
and U11796 (N_11796,N_10672,N_11059);
nor U11797 (N_11797,N_10496,N_10874);
xor U11798 (N_11798,N_10779,N_10950);
nor U11799 (N_11799,N_10842,N_10931);
nand U11800 (N_11800,N_11089,N_10978);
or U11801 (N_11801,N_10936,N_10516);
or U11802 (N_11802,N_10524,N_10623);
and U11803 (N_11803,N_10905,N_10879);
nand U11804 (N_11804,N_10576,N_10738);
nor U11805 (N_11805,N_10538,N_10440);
and U11806 (N_11806,N_10487,N_11118);
nor U11807 (N_11807,N_10585,N_11033);
and U11808 (N_11808,N_10544,N_10663);
and U11809 (N_11809,N_11118,N_10506);
and U11810 (N_11810,N_10582,N_10899);
or U11811 (N_11811,N_11190,N_10931);
nand U11812 (N_11812,N_10906,N_10664);
nor U11813 (N_11813,N_11058,N_10725);
and U11814 (N_11814,N_10478,N_11040);
nor U11815 (N_11815,N_11072,N_10702);
xor U11816 (N_11816,N_10782,N_10923);
xor U11817 (N_11817,N_11132,N_10946);
or U11818 (N_11818,N_10918,N_10408);
nand U11819 (N_11819,N_10620,N_10503);
or U11820 (N_11820,N_10423,N_11199);
or U11821 (N_11821,N_10598,N_10809);
or U11822 (N_11822,N_10760,N_10734);
xnor U11823 (N_11823,N_10850,N_10938);
or U11824 (N_11824,N_10977,N_10520);
nor U11825 (N_11825,N_10974,N_10488);
and U11826 (N_11826,N_10525,N_10998);
and U11827 (N_11827,N_10952,N_10750);
nand U11828 (N_11828,N_10765,N_10881);
nand U11829 (N_11829,N_10989,N_10753);
nor U11830 (N_11830,N_10544,N_10494);
or U11831 (N_11831,N_10527,N_11164);
nor U11832 (N_11832,N_11003,N_10924);
nand U11833 (N_11833,N_11057,N_11191);
and U11834 (N_11834,N_10510,N_11014);
or U11835 (N_11835,N_10827,N_10875);
nor U11836 (N_11836,N_10946,N_10924);
nand U11837 (N_11837,N_10603,N_10646);
xor U11838 (N_11838,N_10669,N_10525);
or U11839 (N_11839,N_10450,N_10442);
or U11840 (N_11840,N_11059,N_10776);
xnor U11841 (N_11841,N_10840,N_10678);
nand U11842 (N_11842,N_11082,N_11076);
and U11843 (N_11843,N_10893,N_11063);
nand U11844 (N_11844,N_10520,N_10675);
nand U11845 (N_11845,N_11129,N_10799);
or U11846 (N_11846,N_10930,N_10695);
xor U11847 (N_11847,N_10588,N_11019);
nor U11848 (N_11848,N_10748,N_10827);
xnor U11849 (N_11849,N_11157,N_11132);
nand U11850 (N_11850,N_11045,N_11034);
xnor U11851 (N_11851,N_11113,N_10694);
nor U11852 (N_11852,N_10883,N_10876);
nand U11853 (N_11853,N_10960,N_10895);
nor U11854 (N_11854,N_11155,N_10759);
and U11855 (N_11855,N_10603,N_10811);
nor U11856 (N_11856,N_10846,N_10488);
or U11857 (N_11857,N_11096,N_10951);
nand U11858 (N_11858,N_10691,N_10670);
and U11859 (N_11859,N_10874,N_10611);
nor U11860 (N_11860,N_10915,N_11179);
xor U11861 (N_11861,N_11113,N_10520);
and U11862 (N_11862,N_10964,N_10464);
xnor U11863 (N_11863,N_10809,N_11068);
nand U11864 (N_11864,N_11099,N_11035);
nand U11865 (N_11865,N_10738,N_10494);
nor U11866 (N_11866,N_10867,N_10851);
and U11867 (N_11867,N_10457,N_11070);
or U11868 (N_11868,N_11182,N_10630);
or U11869 (N_11869,N_10449,N_11113);
and U11870 (N_11870,N_10980,N_10710);
xnor U11871 (N_11871,N_10817,N_10496);
xnor U11872 (N_11872,N_10572,N_10536);
nor U11873 (N_11873,N_11173,N_10797);
or U11874 (N_11874,N_10413,N_11095);
nand U11875 (N_11875,N_11157,N_10995);
or U11876 (N_11876,N_10679,N_10766);
nand U11877 (N_11877,N_10927,N_11038);
or U11878 (N_11878,N_10797,N_11117);
and U11879 (N_11879,N_10874,N_10623);
nand U11880 (N_11880,N_10574,N_10996);
xor U11881 (N_11881,N_10469,N_10566);
nand U11882 (N_11882,N_10590,N_10579);
xnor U11883 (N_11883,N_11196,N_11104);
nor U11884 (N_11884,N_10699,N_10630);
or U11885 (N_11885,N_11150,N_10670);
nand U11886 (N_11886,N_10656,N_10952);
nor U11887 (N_11887,N_10900,N_10863);
or U11888 (N_11888,N_10875,N_10495);
xnor U11889 (N_11889,N_10537,N_10683);
nor U11890 (N_11890,N_10974,N_10805);
or U11891 (N_11891,N_10824,N_11187);
or U11892 (N_11892,N_11106,N_10653);
or U11893 (N_11893,N_10559,N_10661);
or U11894 (N_11894,N_11002,N_11148);
xnor U11895 (N_11895,N_10915,N_11028);
nor U11896 (N_11896,N_11156,N_10816);
xnor U11897 (N_11897,N_10407,N_10948);
xor U11898 (N_11898,N_10572,N_10902);
and U11899 (N_11899,N_10555,N_11015);
or U11900 (N_11900,N_10554,N_10828);
and U11901 (N_11901,N_10409,N_10402);
or U11902 (N_11902,N_10600,N_10883);
and U11903 (N_11903,N_10641,N_10503);
xnor U11904 (N_11904,N_10458,N_11082);
or U11905 (N_11905,N_10602,N_10701);
nor U11906 (N_11906,N_10552,N_10997);
nor U11907 (N_11907,N_10989,N_11172);
or U11908 (N_11908,N_10549,N_10680);
or U11909 (N_11909,N_11000,N_10922);
nand U11910 (N_11910,N_10774,N_11093);
nor U11911 (N_11911,N_11136,N_10814);
xor U11912 (N_11912,N_10519,N_10434);
or U11913 (N_11913,N_10607,N_10536);
and U11914 (N_11914,N_11144,N_11069);
nor U11915 (N_11915,N_11003,N_10528);
nor U11916 (N_11916,N_10584,N_11110);
or U11917 (N_11917,N_10505,N_11031);
nand U11918 (N_11918,N_10893,N_10510);
nand U11919 (N_11919,N_10510,N_10749);
nor U11920 (N_11920,N_10667,N_10864);
xnor U11921 (N_11921,N_10410,N_10634);
xnor U11922 (N_11922,N_10773,N_11054);
and U11923 (N_11923,N_10890,N_10759);
and U11924 (N_11924,N_10648,N_10627);
and U11925 (N_11925,N_10962,N_10772);
or U11926 (N_11926,N_11171,N_10820);
and U11927 (N_11927,N_10660,N_10831);
or U11928 (N_11928,N_10684,N_10608);
nor U11929 (N_11929,N_10581,N_11162);
nand U11930 (N_11930,N_11096,N_10788);
and U11931 (N_11931,N_10704,N_10832);
xor U11932 (N_11932,N_10477,N_10498);
xor U11933 (N_11933,N_10466,N_10405);
xnor U11934 (N_11934,N_10568,N_10434);
or U11935 (N_11935,N_10553,N_10971);
and U11936 (N_11936,N_10468,N_10909);
nor U11937 (N_11937,N_10451,N_10572);
xnor U11938 (N_11938,N_10858,N_10954);
and U11939 (N_11939,N_10658,N_11053);
xor U11940 (N_11940,N_11148,N_10685);
or U11941 (N_11941,N_10617,N_10560);
nor U11942 (N_11942,N_10789,N_10681);
nor U11943 (N_11943,N_10480,N_10980);
or U11944 (N_11944,N_10939,N_10816);
and U11945 (N_11945,N_10581,N_10591);
nand U11946 (N_11946,N_10677,N_10896);
or U11947 (N_11947,N_10415,N_11001);
nand U11948 (N_11948,N_10753,N_10529);
nor U11949 (N_11949,N_11050,N_10551);
nor U11950 (N_11950,N_10482,N_10620);
and U11951 (N_11951,N_11183,N_10694);
nand U11952 (N_11952,N_11065,N_11154);
nand U11953 (N_11953,N_11024,N_10998);
xor U11954 (N_11954,N_11129,N_11049);
nor U11955 (N_11955,N_11180,N_11158);
nand U11956 (N_11956,N_11170,N_10646);
nor U11957 (N_11957,N_10931,N_11183);
nor U11958 (N_11958,N_11098,N_10700);
nand U11959 (N_11959,N_10482,N_11076);
xnor U11960 (N_11960,N_10409,N_10536);
xnor U11961 (N_11961,N_10640,N_10730);
and U11962 (N_11962,N_10960,N_10413);
xnor U11963 (N_11963,N_11166,N_11084);
and U11964 (N_11964,N_10479,N_10647);
and U11965 (N_11965,N_10573,N_10561);
or U11966 (N_11966,N_10834,N_10689);
or U11967 (N_11967,N_11082,N_10965);
xnor U11968 (N_11968,N_10902,N_10648);
or U11969 (N_11969,N_10947,N_10583);
or U11970 (N_11970,N_10940,N_10608);
xor U11971 (N_11971,N_11147,N_10726);
nor U11972 (N_11972,N_11115,N_10736);
nand U11973 (N_11973,N_10990,N_11042);
xor U11974 (N_11974,N_10847,N_10811);
nor U11975 (N_11975,N_10704,N_11143);
or U11976 (N_11976,N_10510,N_11024);
nand U11977 (N_11977,N_10978,N_10611);
nand U11978 (N_11978,N_10673,N_10608);
xnor U11979 (N_11979,N_10605,N_10721);
nor U11980 (N_11980,N_10593,N_10972);
xnor U11981 (N_11981,N_10936,N_10856);
or U11982 (N_11982,N_10500,N_10579);
xnor U11983 (N_11983,N_11036,N_11091);
nand U11984 (N_11984,N_11180,N_11008);
or U11985 (N_11985,N_10950,N_10789);
nand U11986 (N_11986,N_11193,N_10920);
nand U11987 (N_11987,N_11168,N_10923);
and U11988 (N_11988,N_10930,N_10561);
xnor U11989 (N_11989,N_10515,N_10427);
and U11990 (N_11990,N_10497,N_10470);
and U11991 (N_11991,N_10510,N_10676);
nor U11992 (N_11992,N_10682,N_11008);
nand U11993 (N_11993,N_10728,N_11161);
and U11994 (N_11994,N_10610,N_10847);
nor U11995 (N_11995,N_10871,N_10538);
xnor U11996 (N_11996,N_10488,N_10653);
nor U11997 (N_11997,N_10405,N_11079);
xnor U11998 (N_11998,N_10463,N_10984);
nand U11999 (N_11999,N_11119,N_10957);
xor U12000 (N_12000,N_11847,N_11490);
nor U12001 (N_12001,N_11496,N_11544);
or U12002 (N_12002,N_11231,N_11462);
xnor U12003 (N_12003,N_11829,N_11521);
nand U12004 (N_12004,N_11629,N_11283);
xnor U12005 (N_12005,N_11694,N_11926);
nand U12006 (N_12006,N_11279,N_11662);
or U12007 (N_12007,N_11667,N_11232);
or U12008 (N_12008,N_11796,N_11583);
nor U12009 (N_12009,N_11359,N_11921);
or U12010 (N_12010,N_11513,N_11930);
or U12011 (N_12011,N_11449,N_11611);
nor U12012 (N_12012,N_11377,N_11246);
nand U12013 (N_12013,N_11242,N_11207);
nor U12014 (N_12014,N_11789,N_11491);
xor U12015 (N_12015,N_11946,N_11965);
and U12016 (N_12016,N_11392,N_11675);
xor U12017 (N_12017,N_11226,N_11233);
or U12018 (N_12018,N_11515,N_11944);
nand U12019 (N_12019,N_11707,N_11722);
or U12020 (N_12020,N_11618,N_11399);
and U12021 (N_12021,N_11769,N_11969);
nor U12022 (N_12022,N_11940,N_11428);
or U12023 (N_12023,N_11295,N_11846);
or U12024 (N_12024,N_11748,N_11976);
and U12025 (N_12025,N_11455,N_11656);
nand U12026 (N_12026,N_11645,N_11451);
and U12027 (N_12027,N_11999,N_11585);
nor U12028 (N_12028,N_11660,N_11463);
or U12029 (N_12029,N_11784,N_11743);
and U12030 (N_12030,N_11948,N_11519);
xor U12031 (N_12031,N_11209,N_11783);
and U12032 (N_12032,N_11276,N_11813);
nand U12033 (N_12033,N_11894,N_11863);
nand U12034 (N_12034,N_11270,N_11693);
nand U12035 (N_12035,N_11380,N_11958);
nor U12036 (N_12036,N_11872,N_11402);
and U12037 (N_12037,N_11875,N_11573);
xor U12038 (N_12038,N_11814,N_11736);
and U12039 (N_12039,N_11354,N_11827);
or U12040 (N_12040,N_11838,N_11775);
xor U12041 (N_12041,N_11780,N_11841);
nor U12042 (N_12042,N_11897,N_11777);
and U12043 (N_12043,N_11746,N_11737);
nand U12044 (N_12044,N_11826,N_11729);
nand U12045 (N_12045,N_11211,N_11772);
or U12046 (N_12046,N_11401,N_11778);
nand U12047 (N_12047,N_11365,N_11333);
nand U12048 (N_12048,N_11712,N_11981);
nand U12049 (N_12049,N_11773,N_11854);
or U12050 (N_12050,N_11507,N_11447);
xnor U12051 (N_12051,N_11351,N_11297);
nand U12052 (N_12052,N_11364,N_11692);
nand U12053 (N_12053,N_11408,N_11832);
nand U12054 (N_12054,N_11835,N_11326);
xnor U12055 (N_12055,N_11749,N_11934);
and U12056 (N_12056,N_11711,N_11222);
nor U12057 (N_12057,N_11882,N_11848);
and U12058 (N_12058,N_11388,N_11757);
nand U12059 (N_12059,N_11661,N_11484);
and U12060 (N_12060,N_11240,N_11298);
nand U12061 (N_12061,N_11717,N_11954);
and U12062 (N_12062,N_11918,N_11208);
and U12063 (N_12063,N_11422,N_11497);
nor U12064 (N_12064,N_11895,N_11337);
and U12065 (N_12065,N_11723,N_11647);
xor U12066 (N_12066,N_11836,N_11349);
and U12067 (N_12067,N_11517,N_11459);
xor U12068 (N_12068,N_11753,N_11621);
nor U12069 (N_12069,N_11372,N_11433);
or U12070 (N_12070,N_11442,N_11239);
or U12071 (N_12071,N_11443,N_11458);
nand U12072 (N_12072,N_11676,N_11902);
and U12073 (N_12073,N_11465,N_11395);
or U12074 (N_12074,N_11911,N_11810);
nand U12075 (N_12075,N_11523,N_11935);
xnor U12076 (N_12076,N_11642,N_11899);
nand U12077 (N_12077,N_11236,N_11672);
and U12078 (N_12078,N_11527,N_11261);
nor U12079 (N_12079,N_11464,N_11360);
or U12080 (N_12080,N_11310,N_11986);
nor U12081 (N_12081,N_11452,N_11390);
nor U12082 (N_12082,N_11367,N_11885);
nor U12083 (N_12083,N_11213,N_11909);
or U12084 (N_12084,N_11529,N_11924);
nand U12085 (N_12085,N_11602,N_11557);
nand U12086 (N_12086,N_11430,N_11329);
xnor U12087 (N_12087,N_11851,N_11666);
xnor U12088 (N_12088,N_11738,N_11649);
xor U12089 (N_12089,N_11331,N_11570);
or U12090 (N_12090,N_11963,N_11330);
xor U12091 (N_12091,N_11925,N_11845);
xor U12092 (N_12092,N_11795,N_11368);
nand U12093 (N_12093,N_11339,N_11237);
or U12094 (N_12094,N_11514,N_11375);
nor U12095 (N_12095,N_11785,N_11385);
xnor U12096 (N_12096,N_11949,N_11891);
xnor U12097 (N_12097,N_11244,N_11959);
xnor U12098 (N_12098,N_11866,N_11929);
nor U12099 (N_12099,N_11831,N_11639);
nor U12100 (N_12100,N_11302,N_11679);
xnor U12101 (N_12101,N_11830,N_11467);
nand U12102 (N_12102,N_11724,N_11898);
or U12103 (N_12103,N_11334,N_11598);
xor U12104 (N_12104,N_11290,N_11445);
or U12105 (N_12105,N_11821,N_11210);
and U12106 (N_12106,N_11892,N_11366);
or U12107 (N_12107,N_11828,N_11426);
xor U12108 (N_12108,N_11665,N_11802);
and U12109 (N_12109,N_11411,N_11284);
nor U12110 (N_12110,N_11977,N_11238);
and U12111 (N_12111,N_11914,N_11271);
xor U12112 (N_12112,N_11945,N_11254);
or U12113 (N_12113,N_11609,N_11912);
and U12114 (N_12114,N_11974,N_11715);
xnor U12115 (N_12115,N_11750,N_11747);
nor U12116 (N_12116,N_11876,N_11384);
nand U12117 (N_12117,N_11413,N_11460);
nand U12118 (N_12118,N_11640,N_11506);
and U12119 (N_12119,N_11528,N_11868);
xnor U12120 (N_12120,N_11584,N_11241);
nand U12121 (N_12121,N_11325,N_11978);
xnor U12122 (N_12122,N_11985,N_11774);
or U12123 (N_12123,N_11601,N_11561);
xor U12124 (N_12124,N_11691,N_11708);
nand U12125 (N_12125,N_11476,N_11756);
nor U12126 (N_12126,N_11684,N_11670);
or U12127 (N_12127,N_11296,N_11355);
and U12128 (N_12128,N_11989,N_11888);
xnor U12129 (N_12129,N_11352,N_11531);
and U12130 (N_12130,N_11904,N_11568);
or U12131 (N_12131,N_11713,N_11923);
xor U12132 (N_12132,N_11417,N_11424);
and U12133 (N_12133,N_11804,N_11571);
nand U12134 (N_12134,N_11590,N_11993);
xnor U12135 (N_12135,N_11627,N_11504);
nor U12136 (N_12136,N_11951,N_11732);
nand U12137 (N_12137,N_11794,N_11663);
xnor U12138 (N_12138,N_11953,N_11908);
nand U12139 (N_12139,N_11274,N_11341);
nand U12140 (N_12140,N_11674,N_11499);
nand U12141 (N_12141,N_11805,N_11867);
nor U12142 (N_12142,N_11555,N_11658);
nor U12143 (N_12143,N_11710,N_11536);
and U12144 (N_12144,N_11538,N_11787);
nand U12145 (N_12145,N_11577,N_11525);
xor U12146 (N_12146,N_11680,N_11450);
nor U12147 (N_12147,N_11806,N_11797);
xnor U12148 (N_12148,N_11346,N_11520);
nor U12149 (N_12149,N_11503,N_11644);
nand U12150 (N_12150,N_11281,N_11980);
nor U12151 (N_12151,N_11473,N_11509);
nand U12152 (N_12152,N_11324,N_11861);
nand U12153 (N_12153,N_11540,N_11630);
or U12154 (N_12154,N_11358,N_11235);
nor U12155 (N_12155,N_11628,N_11441);
and U12156 (N_12156,N_11219,N_11637);
nand U12157 (N_12157,N_11900,N_11403);
nand U12158 (N_12158,N_11860,N_11466);
xor U12159 (N_12159,N_11728,N_11825);
xnor U12160 (N_12160,N_11396,N_11816);
nor U12161 (N_12161,N_11356,N_11734);
or U12162 (N_12162,N_11952,N_11489);
nor U12163 (N_12163,N_11942,N_11698);
xnor U12164 (N_12164,N_11970,N_11842);
nand U12165 (N_12165,N_11225,N_11664);
xnor U12166 (N_12166,N_11881,N_11361);
and U12167 (N_12167,N_11655,N_11852);
nand U12168 (N_12168,N_11532,N_11652);
nor U12169 (N_12169,N_11688,N_11456);
and U12170 (N_12170,N_11543,N_11487);
nor U12171 (N_12171,N_11457,N_11500);
nand U12172 (N_12172,N_11932,N_11376);
and U12173 (N_12173,N_11409,N_11558);
or U12174 (N_12174,N_11414,N_11906);
nor U12175 (N_12175,N_11947,N_11307);
xnor U12176 (N_12176,N_11844,N_11379);
nand U12177 (N_12177,N_11956,N_11579);
nand U12178 (N_12178,N_11998,N_11311);
nand U12179 (N_12179,N_11799,N_11893);
and U12180 (N_12180,N_11335,N_11471);
nor U12181 (N_12181,N_11404,N_11511);
or U12182 (N_12182,N_11348,N_11393);
nor U12183 (N_12183,N_11595,N_11291);
and U12184 (N_12184,N_11822,N_11766);
or U12185 (N_12185,N_11927,N_11982);
nand U12186 (N_12186,N_11420,N_11478);
nor U12187 (N_12187,N_11383,N_11870);
xnor U12188 (N_12188,N_11322,N_11243);
or U12189 (N_12189,N_11771,N_11586);
nand U12190 (N_12190,N_11542,N_11735);
xor U12191 (N_12191,N_11683,N_11770);
xnor U12192 (N_12192,N_11318,N_11480);
nor U12193 (N_12193,N_11634,N_11622);
xor U12194 (N_12194,N_11287,N_11559);
nand U12195 (N_12195,N_11865,N_11481);
or U12196 (N_12196,N_11657,N_11537);
nand U12197 (N_12197,N_11915,N_11943);
nand U12198 (N_12198,N_11305,N_11839);
xor U12199 (N_12199,N_11338,N_11938);
nor U12200 (N_12200,N_11321,N_11421);
xor U12201 (N_12201,N_11916,N_11488);
nor U12202 (N_12202,N_11883,N_11817);
or U12203 (N_12203,N_11887,N_11397);
and U12204 (N_12204,N_11638,N_11907);
nand U12205 (N_12205,N_11438,N_11505);
nand U12206 (N_12206,N_11415,N_11823);
nand U12207 (N_12207,N_11964,N_11607);
nand U12208 (N_12208,N_11873,N_11782);
nor U12209 (N_12209,N_11919,N_11435);
or U12210 (N_12210,N_11840,N_11314);
nand U12211 (N_12211,N_11858,N_11896);
nand U12212 (N_12212,N_11556,N_11398);
or U12213 (N_12213,N_11603,N_11578);
or U12214 (N_12214,N_11502,N_11546);
nor U12215 (N_12215,N_11687,N_11850);
and U12216 (N_12216,N_11880,N_11677);
or U12217 (N_12217,N_11790,N_11686);
nand U12218 (N_12218,N_11400,N_11535);
and U12219 (N_12219,N_11701,N_11234);
xnor U12220 (N_12220,N_11983,N_11461);
or U12221 (N_12221,N_11522,N_11328);
and U12222 (N_12222,N_11988,N_11903);
or U12223 (N_12223,N_11220,N_11316);
xor U12224 (N_12224,N_11575,N_11760);
and U12225 (N_12225,N_11597,N_11751);
or U12226 (N_12226,N_11659,N_11574);
xnor U12227 (N_12227,N_11215,N_11886);
xor U12228 (N_12228,N_11793,N_11263);
or U12229 (N_12229,N_11987,N_11444);
xor U12230 (N_12230,N_11494,N_11669);
or U12231 (N_12231,N_11569,N_11306);
xnor U12232 (N_12232,N_11961,N_11257);
or U12233 (N_12233,N_11262,N_11347);
xor U12234 (N_12234,N_11733,N_11648);
nand U12235 (N_12235,N_11332,N_11572);
or U12236 (N_12236,N_11937,N_11275);
nand U12237 (N_12237,N_11716,N_11779);
or U12238 (N_12238,N_11317,N_11820);
nor U12239 (N_12239,N_11800,N_11418);
nand U12240 (N_12240,N_11984,N_11495);
xnor U12241 (N_12241,N_11624,N_11615);
xnor U12242 (N_12242,N_11991,N_11264);
xnor U12243 (N_12243,N_11690,N_11289);
xor U12244 (N_12244,N_11957,N_11250);
nor U12245 (N_12245,N_11931,N_11801);
nor U12246 (N_12246,N_11541,N_11371);
nor U12247 (N_12247,N_11253,N_11510);
xnor U12248 (N_12248,N_11437,N_11255);
xnor U12249 (N_12249,N_11706,N_11547);
nand U12250 (N_12250,N_11619,N_11620);
and U12251 (N_12251,N_11812,N_11973);
and U12252 (N_12252,N_11752,N_11968);
or U12253 (N_12253,N_11268,N_11990);
nor U12254 (N_12254,N_11596,N_11350);
and U12255 (N_12255,N_11767,N_11285);
nor U12256 (N_12256,N_11608,N_11551);
nand U12257 (N_12257,N_11612,N_11200);
and U12258 (N_12258,N_11901,N_11533);
nor U12259 (N_12259,N_11224,N_11763);
or U12260 (N_12260,N_11731,N_11299);
nand U12261 (N_12261,N_11212,N_11266);
nand U12262 (N_12262,N_11997,N_11636);
nor U12263 (N_12263,N_11327,N_11292);
nand U12264 (N_12264,N_11563,N_11834);
nor U12265 (N_12265,N_11580,N_11759);
nand U12266 (N_12266,N_11933,N_11249);
nor U12267 (N_12267,N_11439,N_11248);
xor U12268 (N_12268,N_11277,N_11631);
xnor U12269 (N_12269,N_11966,N_11524);
nor U12270 (N_12270,N_11434,N_11600);
xnor U12271 (N_12271,N_11781,N_11995);
and U12272 (N_12272,N_11792,N_11941);
xnor U12273 (N_12273,N_11604,N_11576);
nand U12274 (N_12274,N_11626,N_11971);
xor U12275 (N_12275,N_11389,N_11501);
xor U12276 (N_12276,N_11227,N_11344);
and U12277 (N_12277,N_11381,N_11319);
and U12278 (N_12278,N_11407,N_11718);
or U12279 (N_12279,N_11764,N_11856);
nor U12280 (N_12280,N_11641,N_11725);
nand U12281 (N_12281,N_11755,N_11996);
or U12282 (N_12282,N_11431,N_11218);
nor U12283 (N_12283,N_11689,N_11593);
and U12284 (N_12284,N_11553,N_11857);
and U12285 (N_12285,N_11837,N_11278);
and U12286 (N_12286,N_11623,N_11405);
nand U12287 (N_12287,N_11651,N_11229);
and U12288 (N_12288,N_11486,N_11475);
and U12289 (N_12289,N_11740,N_11599);
xnor U12290 (N_12290,N_11862,N_11758);
xnor U12291 (N_12291,N_11654,N_11653);
and U12292 (N_12292,N_11345,N_11703);
nand U12293 (N_12293,N_11591,N_11343);
nor U12294 (N_12294,N_11681,N_11765);
or U12295 (N_12295,N_11228,N_11362);
or U12296 (N_12296,N_11286,N_11960);
nor U12297 (N_12297,N_11745,N_11616);
nor U12298 (N_12298,N_11429,N_11482);
xnor U12299 (N_12299,N_11550,N_11582);
nand U12300 (N_12300,N_11453,N_11419);
nor U12301 (N_12301,N_11518,N_11288);
nand U12302 (N_12302,N_11606,N_11633);
xnor U12303 (N_12303,N_11992,N_11762);
xor U12304 (N_12304,N_11394,N_11472);
xor U12305 (N_12305,N_11313,N_11245);
nor U12306 (N_12306,N_11741,N_11920);
nor U12307 (N_12307,N_11632,N_11205);
and U12308 (N_12308,N_11259,N_11512);
and U12309 (N_12309,N_11548,N_11280);
xnor U12310 (N_12310,N_11468,N_11353);
or U12311 (N_12311,N_11849,N_11539);
nand U12312 (N_12312,N_11605,N_11391);
and U12313 (N_12313,N_11357,N_11855);
nor U12314 (N_12314,N_11614,N_11962);
and U12315 (N_12315,N_11878,N_11410);
xnor U12316 (N_12316,N_11217,N_11699);
nand U12317 (N_12317,N_11566,N_11534);
nand U12318 (N_12318,N_11833,N_11650);
and U12319 (N_12319,N_11871,N_11809);
and U12320 (N_12320,N_11483,N_11702);
or U12321 (N_12321,N_11309,N_11416);
nand U12322 (N_12322,N_11877,N_11776);
nand U12323 (N_12323,N_11294,N_11386);
xnor U12324 (N_12324,N_11247,N_11204);
or U12325 (N_12325,N_11979,N_11214);
and U12326 (N_12326,N_11588,N_11440);
xnor U12327 (N_12327,N_11251,N_11719);
or U12328 (N_12328,N_11492,N_11587);
nand U12329 (N_12329,N_11890,N_11202);
nor U12330 (N_12330,N_11387,N_11721);
or U12331 (N_12331,N_11552,N_11549);
and U12332 (N_12332,N_11530,N_11554);
nand U12333 (N_12333,N_11293,N_11859);
or U12334 (N_12334,N_11269,N_11673);
and U12335 (N_12335,N_11370,N_11581);
or U12336 (N_12336,N_11695,N_11788);
nand U12337 (N_12337,N_11267,N_11206);
xor U12338 (N_12338,N_11252,N_11742);
xnor U12339 (N_12339,N_11798,N_11709);
and U12340 (N_12340,N_11905,N_11373);
nand U12341 (N_12341,N_11625,N_11950);
and U12342 (N_12342,N_11260,N_11646);
and U12343 (N_12343,N_11939,N_11432);
nand U12344 (N_12344,N_11994,N_11273);
and U12345 (N_12345,N_11975,N_11913);
xnor U12346 (N_12346,N_11714,N_11594);
nor U12347 (N_12347,N_11589,N_11282);
or U12348 (N_12348,N_11223,N_11678);
nand U12349 (N_12349,N_11300,N_11374);
and U12350 (N_12350,N_11696,N_11425);
xor U12351 (N_12351,N_11312,N_11922);
or U12352 (N_12352,N_11727,N_11869);
or U12353 (N_12353,N_11843,N_11363);
xor U12354 (N_12354,N_11791,N_11704);
and U12355 (N_12355,N_11808,N_11508);
or U12356 (N_12356,N_11336,N_11203);
nand U12357 (N_12357,N_11201,N_11617);
xor U12358 (N_12358,N_11955,N_11256);
nand U12359 (N_12359,N_11744,N_11272);
nor U12360 (N_12360,N_11526,N_11342);
nand U12361 (N_12361,N_11315,N_11567);
nor U12362 (N_12362,N_11884,N_11382);
nor U12363 (N_12363,N_11889,N_11967);
or U12364 (N_12364,N_11671,N_11448);
or U12365 (N_12365,N_11697,N_11928);
nand U12366 (N_12366,N_11720,N_11485);
xor U12367 (N_12367,N_11910,N_11824);
nor U12368 (N_12368,N_11864,N_11564);
or U12369 (N_12369,N_11516,N_11436);
xnor U12370 (N_12370,N_11807,N_11560);
nor U12371 (N_12371,N_11216,N_11754);
nor U12372 (N_12372,N_11423,N_11304);
and U12373 (N_12373,N_11972,N_11454);
or U12374 (N_12374,N_11545,N_11221);
and U12375 (N_12375,N_11320,N_11768);
and U12376 (N_12376,N_11562,N_11668);
nor U12377 (N_12377,N_11879,N_11258);
nor U12378 (N_12378,N_11479,N_11303);
or U12379 (N_12379,N_11761,N_11739);
xor U12380 (N_12380,N_11786,N_11301);
nor U12381 (N_12381,N_11635,N_11493);
xor U12382 (N_12382,N_11323,N_11936);
nor U12383 (N_12383,N_11815,N_11498);
xor U12384 (N_12384,N_11378,N_11474);
xnor U12385 (N_12385,N_11470,N_11726);
xnor U12386 (N_12386,N_11811,N_11685);
nor U12387 (N_12387,N_11874,N_11700);
nor U12388 (N_12388,N_11917,N_11682);
nand U12389 (N_12389,N_11819,N_11406);
and U12390 (N_12390,N_11610,N_11308);
xor U12391 (N_12391,N_11592,N_11565);
and U12392 (N_12392,N_11643,N_11803);
or U12393 (N_12393,N_11818,N_11265);
nor U12394 (N_12394,N_11477,N_11369);
xnor U12395 (N_12395,N_11446,N_11469);
nand U12396 (N_12396,N_11613,N_11340);
nand U12397 (N_12397,N_11230,N_11412);
xor U12398 (N_12398,N_11853,N_11705);
nand U12399 (N_12399,N_11730,N_11427);
xor U12400 (N_12400,N_11982,N_11459);
nor U12401 (N_12401,N_11790,N_11531);
nand U12402 (N_12402,N_11875,N_11864);
nor U12403 (N_12403,N_11813,N_11480);
xor U12404 (N_12404,N_11284,N_11716);
xnor U12405 (N_12405,N_11307,N_11657);
nand U12406 (N_12406,N_11221,N_11530);
and U12407 (N_12407,N_11487,N_11350);
nand U12408 (N_12408,N_11708,N_11936);
nand U12409 (N_12409,N_11846,N_11377);
and U12410 (N_12410,N_11471,N_11939);
or U12411 (N_12411,N_11580,N_11270);
xor U12412 (N_12412,N_11299,N_11980);
nor U12413 (N_12413,N_11622,N_11901);
nand U12414 (N_12414,N_11785,N_11576);
and U12415 (N_12415,N_11205,N_11792);
and U12416 (N_12416,N_11603,N_11649);
and U12417 (N_12417,N_11748,N_11893);
nand U12418 (N_12418,N_11757,N_11955);
nor U12419 (N_12419,N_11732,N_11381);
xnor U12420 (N_12420,N_11975,N_11761);
or U12421 (N_12421,N_11538,N_11237);
or U12422 (N_12422,N_11555,N_11714);
nor U12423 (N_12423,N_11653,N_11638);
nor U12424 (N_12424,N_11341,N_11788);
or U12425 (N_12425,N_11934,N_11353);
xor U12426 (N_12426,N_11441,N_11967);
nand U12427 (N_12427,N_11757,N_11205);
and U12428 (N_12428,N_11348,N_11984);
nand U12429 (N_12429,N_11929,N_11387);
and U12430 (N_12430,N_11222,N_11493);
nor U12431 (N_12431,N_11926,N_11838);
or U12432 (N_12432,N_11222,N_11660);
or U12433 (N_12433,N_11687,N_11206);
and U12434 (N_12434,N_11290,N_11998);
or U12435 (N_12435,N_11426,N_11959);
xnor U12436 (N_12436,N_11764,N_11227);
nand U12437 (N_12437,N_11754,N_11293);
xor U12438 (N_12438,N_11832,N_11779);
or U12439 (N_12439,N_11668,N_11969);
nand U12440 (N_12440,N_11525,N_11332);
nand U12441 (N_12441,N_11809,N_11814);
xnor U12442 (N_12442,N_11865,N_11659);
or U12443 (N_12443,N_11453,N_11367);
and U12444 (N_12444,N_11599,N_11304);
xnor U12445 (N_12445,N_11569,N_11356);
nand U12446 (N_12446,N_11598,N_11202);
or U12447 (N_12447,N_11297,N_11726);
and U12448 (N_12448,N_11274,N_11807);
or U12449 (N_12449,N_11392,N_11305);
and U12450 (N_12450,N_11459,N_11729);
or U12451 (N_12451,N_11845,N_11293);
xnor U12452 (N_12452,N_11287,N_11852);
nor U12453 (N_12453,N_11377,N_11664);
nor U12454 (N_12454,N_11430,N_11896);
and U12455 (N_12455,N_11550,N_11284);
nor U12456 (N_12456,N_11930,N_11481);
or U12457 (N_12457,N_11515,N_11849);
and U12458 (N_12458,N_11284,N_11812);
nor U12459 (N_12459,N_11465,N_11442);
xor U12460 (N_12460,N_11681,N_11489);
nand U12461 (N_12461,N_11473,N_11386);
and U12462 (N_12462,N_11439,N_11368);
xnor U12463 (N_12463,N_11505,N_11352);
or U12464 (N_12464,N_11850,N_11869);
or U12465 (N_12465,N_11635,N_11509);
xnor U12466 (N_12466,N_11435,N_11321);
nand U12467 (N_12467,N_11937,N_11531);
or U12468 (N_12468,N_11547,N_11347);
xnor U12469 (N_12469,N_11412,N_11268);
or U12470 (N_12470,N_11621,N_11774);
nand U12471 (N_12471,N_11390,N_11774);
nor U12472 (N_12472,N_11567,N_11687);
nor U12473 (N_12473,N_11690,N_11360);
nor U12474 (N_12474,N_11287,N_11364);
and U12475 (N_12475,N_11748,N_11367);
and U12476 (N_12476,N_11484,N_11937);
nand U12477 (N_12477,N_11211,N_11777);
xnor U12478 (N_12478,N_11416,N_11305);
nand U12479 (N_12479,N_11407,N_11804);
nor U12480 (N_12480,N_11542,N_11559);
or U12481 (N_12481,N_11209,N_11383);
or U12482 (N_12482,N_11775,N_11356);
xnor U12483 (N_12483,N_11632,N_11481);
or U12484 (N_12484,N_11571,N_11246);
nand U12485 (N_12485,N_11399,N_11479);
nand U12486 (N_12486,N_11899,N_11908);
nand U12487 (N_12487,N_11505,N_11534);
or U12488 (N_12488,N_11793,N_11403);
or U12489 (N_12489,N_11539,N_11896);
nand U12490 (N_12490,N_11383,N_11761);
xor U12491 (N_12491,N_11959,N_11395);
xnor U12492 (N_12492,N_11445,N_11764);
nand U12493 (N_12493,N_11743,N_11920);
xor U12494 (N_12494,N_11347,N_11734);
and U12495 (N_12495,N_11296,N_11329);
nor U12496 (N_12496,N_11396,N_11773);
nor U12497 (N_12497,N_11510,N_11297);
and U12498 (N_12498,N_11991,N_11289);
nor U12499 (N_12499,N_11823,N_11575);
or U12500 (N_12500,N_11349,N_11365);
and U12501 (N_12501,N_11784,N_11261);
and U12502 (N_12502,N_11636,N_11388);
xor U12503 (N_12503,N_11600,N_11998);
xor U12504 (N_12504,N_11874,N_11886);
nand U12505 (N_12505,N_11799,N_11964);
and U12506 (N_12506,N_11850,N_11486);
and U12507 (N_12507,N_11404,N_11966);
or U12508 (N_12508,N_11843,N_11207);
nand U12509 (N_12509,N_11242,N_11951);
nand U12510 (N_12510,N_11255,N_11248);
xor U12511 (N_12511,N_11765,N_11220);
and U12512 (N_12512,N_11219,N_11367);
nand U12513 (N_12513,N_11964,N_11466);
xnor U12514 (N_12514,N_11209,N_11638);
xor U12515 (N_12515,N_11210,N_11287);
and U12516 (N_12516,N_11783,N_11332);
and U12517 (N_12517,N_11812,N_11472);
or U12518 (N_12518,N_11904,N_11282);
and U12519 (N_12519,N_11925,N_11273);
and U12520 (N_12520,N_11888,N_11678);
and U12521 (N_12521,N_11949,N_11429);
nor U12522 (N_12522,N_11860,N_11508);
or U12523 (N_12523,N_11955,N_11505);
xnor U12524 (N_12524,N_11408,N_11991);
nor U12525 (N_12525,N_11650,N_11572);
xnor U12526 (N_12526,N_11940,N_11290);
nor U12527 (N_12527,N_11497,N_11920);
nand U12528 (N_12528,N_11736,N_11416);
nor U12529 (N_12529,N_11868,N_11249);
and U12530 (N_12530,N_11485,N_11343);
nand U12531 (N_12531,N_11531,N_11822);
xnor U12532 (N_12532,N_11523,N_11471);
xor U12533 (N_12533,N_11956,N_11514);
and U12534 (N_12534,N_11850,N_11217);
nand U12535 (N_12535,N_11286,N_11853);
or U12536 (N_12536,N_11696,N_11230);
nand U12537 (N_12537,N_11463,N_11661);
xor U12538 (N_12538,N_11422,N_11592);
and U12539 (N_12539,N_11790,N_11784);
xor U12540 (N_12540,N_11244,N_11697);
nand U12541 (N_12541,N_11219,N_11857);
or U12542 (N_12542,N_11357,N_11466);
or U12543 (N_12543,N_11664,N_11706);
or U12544 (N_12544,N_11350,N_11435);
xor U12545 (N_12545,N_11328,N_11972);
nand U12546 (N_12546,N_11622,N_11757);
nor U12547 (N_12547,N_11755,N_11487);
and U12548 (N_12548,N_11547,N_11673);
nand U12549 (N_12549,N_11692,N_11578);
nand U12550 (N_12550,N_11381,N_11630);
or U12551 (N_12551,N_11338,N_11501);
nor U12552 (N_12552,N_11580,N_11879);
xnor U12553 (N_12553,N_11421,N_11212);
xor U12554 (N_12554,N_11641,N_11214);
or U12555 (N_12555,N_11718,N_11890);
nand U12556 (N_12556,N_11256,N_11642);
and U12557 (N_12557,N_11228,N_11364);
and U12558 (N_12558,N_11474,N_11871);
and U12559 (N_12559,N_11693,N_11510);
nor U12560 (N_12560,N_11269,N_11913);
nor U12561 (N_12561,N_11210,N_11320);
nor U12562 (N_12562,N_11761,N_11485);
nand U12563 (N_12563,N_11979,N_11892);
nor U12564 (N_12564,N_11619,N_11908);
xnor U12565 (N_12565,N_11351,N_11532);
and U12566 (N_12566,N_11547,N_11773);
xor U12567 (N_12567,N_11531,N_11583);
xor U12568 (N_12568,N_11376,N_11357);
nor U12569 (N_12569,N_11978,N_11764);
or U12570 (N_12570,N_11945,N_11748);
and U12571 (N_12571,N_11426,N_11356);
and U12572 (N_12572,N_11767,N_11281);
nand U12573 (N_12573,N_11520,N_11295);
nand U12574 (N_12574,N_11316,N_11460);
and U12575 (N_12575,N_11787,N_11933);
or U12576 (N_12576,N_11627,N_11570);
nor U12577 (N_12577,N_11725,N_11472);
or U12578 (N_12578,N_11686,N_11821);
nor U12579 (N_12579,N_11518,N_11598);
and U12580 (N_12580,N_11914,N_11915);
and U12581 (N_12581,N_11877,N_11735);
xor U12582 (N_12582,N_11529,N_11231);
nand U12583 (N_12583,N_11619,N_11586);
nor U12584 (N_12584,N_11565,N_11674);
xor U12585 (N_12585,N_11260,N_11809);
nand U12586 (N_12586,N_11573,N_11277);
xor U12587 (N_12587,N_11279,N_11434);
nand U12588 (N_12588,N_11208,N_11894);
nand U12589 (N_12589,N_11739,N_11724);
nand U12590 (N_12590,N_11428,N_11352);
nand U12591 (N_12591,N_11697,N_11999);
nor U12592 (N_12592,N_11976,N_11250);
or U12593 (N_12593,N_11527,N_11537);
xnor U12594 (N_12594,N_11611,N_11732);
xnor U12595 (N_12595,N_11693,N_11696);
nand U12596 (N_12596,N_11531,N_11877);
xor U12597 (N_12597,N_11955,N_11269);
nand U12598 (N_12598,N_11967,N_11262);
and U12599 (N_12599,N_11893,N_11454);
or U12600 (N_12600,N_11646,N_11952);
or U12601 (N_12601,N_11715,N_11475);
nor U12602 (N_12602,N_11835,N_11911);
or U12603 (N_12603,N_11382,N_11786);
and U12604 (N_12604,N_11715,N_11392);
or U12605 (N_12605,N_11379,N_11943);
and U12606 (N_12606,N_11808,N_11606);
and U12607 (N_12607,N_11224,N_11814);
and U12608 (N_12608,N_11515,N_11561);
xnor U12609 (N_12609,N_11784,N_11730);
nor U12610 (N_12610,N_11286,N_11749);
nor U12611 (N_12611,N_11386,N_11803);
or U12612 (N_12612,N_11243,N_11970);
or U12613 (N_12613,N_11887,N_11679);
xor U12614 (N_12614,N_11460,N_11357);
and U12615 (N_12615,N_11333,N_11226);
or U12616 (N_12616,N_11444,N_11717);
or U12617 (N_12617,N_11853,N_11647);
nor U12618 (N_12618,N_11654,N_11438);
xor U12619 (N_12619,N_11815,N_11601);
or U12620 (N_12620,N_11202,N_11264);
or U12621 (N_12621,N_11809,N_11408);
nor U12622 (N_12622,N_11632,N_11526);
nand U12623 (N_12623,N_11548,N_11661);
nand U12624 (N_12624,N_11738,N_11372);
and U12625 (N_12625,N_11610,N_11700);
or U12626 (N_12626,N_11819,N_11415);
nor U12627 (N_12627,N_11763,N_11735);
and U12628 (N_12628,N_11668,N_11824);
xor U12629 (N_12629,N_11701,N_11298);
nand U12630 (N_12630,N_11959,N_11943);
nor U12631 (N_12631,N_11801,N_11871);
nor U12632 (N_12632,N_11361,N_11376);
nor U12633 (N_12633,N_11812,N_11554);
xnor U12634 (N_12634,N_11875,N_11380);
or U12635 (N_12635,N_11978,N_11742);
nor U12636 (N_12636,N_11627,N_11980);
nand U12637 (N_12637,N_11892,N_11925);
xnor U12638 (N_12638,N_11273,N_11319);
xnor U12639 (N_12639,N_11562,N_11793);
or U12640 (N_12640,N_11440,N_11393);
or U12641 (N_12641,N_11621,N_11961);
or U12642 (N_12642,N_11512,N_11958);
nor U12643 (N_12643,N_11293,N_11473);
nand U12644 (N_12644,N_11806,N_11881);
xnor U12645 (N_12645,N_11272,N_11626);
nor U12646 (N_12646,N_11762,N_11415);
nand U12647 (N_12647,N_11866,N_11622);
and U12648 (N_12648,N_11766,N_11762);
nand U12649 (N_12649,N_11302,N_11343);
nor U12650 (N_12650,N_11424,N_11859);
and U12651 (N_12651,N_11657,N_11464);
or U12652 (N_12652,N_11365,N_11304);
nor U12653 (N_12653,N_11217,N_11894);
nor U12654 (N_12654,N_11318,N_11674);
nand U12655 (N_12655,N_11752,N_11209);
nor U12656 (N_12656,N_11791,N_11547);
xnor U12657 (N_12657,N_11519,N_11381);
xor U12658 (N_12658,N_11630,N_11285);
xnor U12659 (N_12659,N_11390,N_11356);
nand U12660 (N_12660,N_11728,N_11971);
nor U12661 (N_12661,N_11522,N_11363);
nand U12662 (N_12662,N_11639,N_11435);
nor U12663 (N_12663,N_11759,N_11277);
nor U12664 (N_12664,N_11246,N_11763);
nand U12665 (N_12665,N_11332,N_11368);
and U12666 (N_12666,N_11333,N_11295);
xor U12667 (N_12667,N_11878,N_11355);
nor U12668 (N_12668,N_11879,N_11581);
nand U12669 (N_12669,N_11531,N_11821);
and U12670 (N_12670,N_11338,N_11297);
or U12671 (N_12671,N_11475,N_11342);
nand U12672 (N_12672,N_11335,N_11454);
xor U12673 (N_12673,N_11646,N_11854);
and U12674 (N_12674,N_11554,N_11553);
nor U12675 (N_12675,N_11307,N_11265);
nand U12676 (N_12676,N_11889,N_11338);
nand U12677 (N_12677,N_11666,N_11804);
and U12678 (N_12678,N_11544,N_11826);
nor U12679 (N_12679,N_11956,N_11625);
and U12680 (N_12680,N_11222,N_11898);
xnor U12681 (N_12681,N_11878,N_11294);
and U12682 (N_12682,N_11890,N_11586);
or U12683 (N_12683,N_11547,N_11889);
nand U12684 (N_12684,N_11889,N_11642);
nand U12685 (N_12685,N_11318,N_11993);
and U12686 (N_12686,N_11331,N_11668);
nor U12687 (N_12687,N_11360,N_11934);
xor U12688 (N_12688,N_11780,N_11897);
xnor U12689 (N_12689,N_11354,N_11285);
nand U12690 (N_12690,N_11546,N_11966);
and U12691 (N_12691,N_11649,N_11630);
nand U12692 (N_12692,N_11665,N_11927);
and U12693 (N_12693,N_11694,N_11311);
nor U12694 (N_12694,N_11339,N_11420);
or U12695 (N_12695,N_11874,N_11303);
nand U12696 (N_12696,N_11506,N_11843);
nor U12697 (N_12697,N_11308,N_11928);
and U12698 (N_12698,N_11431,N_11302);
and U12699 (N_12699,N_11646,N_11593);
and U12700 (N_12700,N_11370,N_11416);
xnor U12701 (N_12701,N_11314,N_11472);
nand U12702 (N_12702,N_11316,N_11604);
or U12703 (N_12703,N_11525,N_11793);
and U12704 (N_12704,N_11946,N_11556);
or U12705 (N_12705,N_11988,N_11686);
nor U12706 (N_12706,N_11216,N_11371);
xor U12707 (N_12707,N_11331,N_11993);
xor U12708 (N_12708,N_11442,N_11529);
xor U12709 (N_12709,N_11308,N_11430);
nor U12710 (N_12710,N_11205,N_11602);
or U12711 (N_12711,N_11288,N_11329);
and U12712 (N_12712,N_11338,N_11842);
nand U12713 (N_12713,N_11204,N_11930);
nor U12714 (N_12714,N_11541,N_11941);
or U12715 (N_12715,N_11434,N_11335);
and U12716 (N_12716,N_11616,N_11404);
nor U12717 (N_12717,N_11896,N_11313);
nor U12718 (N_12718,N_11513,N_11795);
nor U12719 (N_12719,N_11364,N_11347);
nand U12720 (N_12720,N_11957,N_11904);
nor U12721 (N_12721,N_11511,N_11674);
xnor U12722 (N_12722,N_11813,N_11501);
nor U12723 (N_12723,N_11877,N_11725);
xor U12724 (N_12724,N_11936,N_11490);
and U12725 (N_12725,N_11398,N_11284);
nor U12726 (N_12726,N_11352,N_11368);
and U12727 (N_12727,N_11678,N_11868);
nor U12728 (N_12728,N_11453,N_11913);
nor U12729 (N_12729,N_11963,N_11488);
nor U12730 (N_12730,N_11525,N_11481);
nand U12731 (N_12731,N_11551,N_11650);
xnor U12732 (N_12732,N_11948,N_11218);
nand U12733 (N_12733,N_11876,N_11404);
xnor U12734 (N_12734,N_11370,N_11729);
and U12735 (N_12735,N_11481,N_11472);
and U12736 (N_12736,N_11957,N_11736);
xnor U12737 (N_12737,N_11397,N_11207);
and U12738 (N_12738,N_11854,N_11492);
nand U12739 (N_12739,N_11583,N_11799);
and U12740 (N_12740,N_11485,N_11214);
xor U12741 (N_12741,N_11726,N_11705);
and U12742 (N_12742,N_11824,N_11434);
nand U12743 (N_12743,N_11928,N_11377);
xnor U12744 (N_12744,N_11258,N_11844);
xnor U12745 (N_12745,N_11355,N_11836);
xor U12746 (N_12746,N_11624,N_11805);
nor U12747 (N_12747,N_11373,N_11804);
or U12748 (N_12748,N_11261,N_11693);
xor U12749 (N_12749,N_11434,N_11266);
and U12750 (N_12750,N_11722,N_11816);
and U12751 (N_12751,N_11235,N_11560);
xnor U12752 (N_12752,N_11410,N_11953);
or U12753 (N_12753,N_11316,N_11684);
or U12754 (N_12754,N_11528,N_11450);
and U12755 (N_12755,N_11324,N_11625);
or U12756 (N_12756,N_11360,N_11842);
and U12757 (N_12757,N_11487,N_11423);
xnor U12758 (N_12758,N_11657,N_11808);
and U12759 (N_12759,N_11572,N_11544);
or U12760 (N_12760,N_11473,N_11697);
nor U12761 (N_12761,N_11483,N_11832);
nor U12762 (N_12762,N_11915,N_11882);
nor U12763 (N_12763,N_11324,N_11796);
and U12764 (N_12764,N_11794,N_11434);
xnor U12765 (N_12765,N_11236,N_11950);
xnor U12766 (N_12766,N_11611,N_11916);
nor U12767 (N_12767,N_11388,N_11407);
xnor U12768 (N_12768,N_11219,N_11895);
or U12769 (N_12769,N_11746,N_11433);
or U12770 (N_12770,N_11447,N_11713);
nor U12771 (N_12771,N_11566,N_11365);
nor U12772 (N_12772,N_11813,N_11392);
nand U12773 (N_12773,N_11911,N_11514);
xor U12774 (N_12774,N_11436,N_11947);
xnor U12775 (N_12775,N_11451,N_11670);
or U12776 (N_12776,N_11993,N_11881);
or U12777 (N_12777,N_11878,N_11663);
and U12778 (N_12778,N_11775,N_11764);
nand U12779 (N_12779,N_11919,N_11867);
or U12780 (N_12780,N_11212,N_11390);
xor U12781 (N_12781,N_11700,N_11887);
xnor U12782 (N_12782,N_11482,N_11529);
nand U12783 (N_12783,N_11434,N_11242);
and U12784 (N_12784,N_11802,N_11295);
nor U12785 (N_12785,N_11853,N_11688);
nor U12786 (N_12786,N_11790,N_11555);
nor U12787 (N_12787,N_11726,N_11359);
nand U12788 (N_12788,N_11911,N_11201);
xor U12789 (N_12789,N_11505,N_11328);
nand U12790 (N_12790,N_11233,N_11922);
nand U12791 (N_12791,N_11336,N_11799);
nand U12792 (N_12792,N_11903,N_11215);
nor U12793 (N_12793,N_11964,N_11272);
or U12794 (N_12794,N_11379,N_11875);
xnor U12795 (N_12795,N_11367,N_11916);
or U12796 (N_12796,N_11870,N_11898);
nor U12797 (N_12797,N_11284,N_11404);
nand U12798 (N_12798,N_11765,N_11974);
nand U12799 (N_12799,N_11796,N_11459);
nor U12800 (N_12800,N_12437,N_12703);
or U12801 (N_12801,N_12371,N_12537);
and U12802 (N_12802,N_12355,N_12126);
or U12803 (N_12803,N_12638,N_12533);
xnor U12804 (N_12804,N_12406,N_12688);
and U12805 (N_12805,N_12786,N_12682);
xnor U12806 (N_12806,N_12395,N_12030);
and U12807 (N_12807,N_12214,N_12404);
and U12808 (N_12808,N_12462,N_12439);
or U12809 (N_12809,N_12665,N_12446);
or U12810 (N_12810,N_12747,N_12066);
or U12811 (N_12811,N_12149,N_12575);
or U12812 (N_12812,N_12620,N_12087);
nor U12813 (N_12813,N_12448,N_12675);
nand U12814 (N_12814,N_12139,N_12231);
nand U12815 (N_12815,N_12138,N_12586);
nor U12816 (N_12816,N_12483,N_12491);
nor U12817 (N_12817,N_12543,N_12497);
nor U12818 (N_12818,N_12168,N_12315);
nand U12819 (N_12819,N_12085,N_12051);
or U12820 (N_12820,N_12579,N_12768);
or U12821 (N_12821,N_12242,N_12245);
and U12822 (N_12822,N_12608,N_12523);
nand U12823 (N_12823,N_12131,N_12719);
or U12824 (N_12824,N_12727,N_12607);
nand U12825 (N_12825,N_12362,N_12076);
nand U12826 (N_12826,N_12264,N_12686);
nor U12827 (N_12827,N_12271,N_12558);
xor U12828 (N_12828,N_12623,N_12295);
nand U12829 (N_12829,N_12089,N_12503);
nand U12830 (N_12830,N_12380,N_12210);
and U12831 (N_12831,N_12609,N_12552);
and U12832 (N_12832,N_12018,N_12148);
or U12833 (N_12833,N_12755,N_12602);
and U12834 (N_12834,N_12181,N_12211);
nor U12835 (N_12835,N_12464,N_12673);
and U12836 (N_12836,N_12569,N_12123);
nand U12837 (N_12837,N_12254,N_12618);
nor U12838 (N_12838,N_12449,N_12068);
or U12839 (N_12839,N_12538,N_12162);
nor U12840 (N_12840,N_12300,N_12329);
or U12841 (N_12841,N_12041,N_12289);
or U12842 (N_12842,N_12209,N_12370);
and U12843 (N_12843,N_12457,N_12422);
xor U12844 (N_12844,N_12029,N_12026);
and U12845 (N_12845,N_12434,N_12224);
nand U12846 (N_12846,N_12384,N_12695);
nand U12847 (N_12847,N_12304,N_12606);
and U12848 (N_12848,N_12206,N_12482);
nand U12849 (N_12849,N_12494,N_12561);
or U12850 (N_12850,N_12364,N_12173);
nor U12851 (N_12851,N_12180,N_12325);
or U12852 (N_12852,N_12192,N_12310);
xnor U12853 (N_12853,N_12440,N_12101);
nor U12854 (N_12854,N_12146,N_12647);
and U12855 (N_12855,N_12738,N_12614);
or U12856 (N_12856,N_12518,N_12689);
nand U12857 (N_12857,N_12700,N_12277);
nand U12858 (N_12858,N_12657,N_12611);
nor U12859 (N_12859,N_12486,N_12770);
xor U12860 (N_12860,N_12221,N_12723);
nand U12861 (N_12861,N_12145,N_12567);
nand U12862 (N_12862,N_12565,N_12474);
and U12863 (N_12863,N_12798,N_12322);
or U12864 (N_12864,N_12663,N_12791);
nor U12865 (N_12865,N_12200,N_12487);
xnor U12866 (N_12866,N_12504,N_12674);
and U12867 (N_12867,N_12094,N_12118);
or U12868 (N_12868,N_12658,N_12296);
and U12869 (N_12869,N_12568,N_12635);
or U12870 (N_12870,N_12025,N_12141);
nand U12871 (N_12871,N_12704,N_12511);
or U12872 (N_12872,N_12773,N_12754);
nand U12873 (N_12873,N_12392,N_12001);
xor U12874 (N_12874,N_12220,N_12515);
and U12875 (N_12875,N_12637,N_12328);
nor U12876 (N_12876,N_12326,N_12044);
or U12877 (N_12877,N_12357,N_12456);
nor U12878 (N_12878,N_12293,N_12728);
nand U12879 (N_12879,N_12130,N_12281);
nor U12880 (N_12880,N_12681,N_12778);
nand U12881 (N_12881,N_12365,N_12722);
or U12882 (N_12882,N_12083,N_12527);
nor U12883 (N_12883,N_12246,N_12046);
xnor U12884 (N_12884,N_12797,N_12276);
or U12885 (N_12885,N_12072,N_12591);
nand U12886 (N_12886,N_12369,N_12147);
nor U12887 (N_12887,N_12261,N_12429);
or U12888 (N_12888,N_12302,N_12493);
xor U12889 (N_12889,N_12646,N_12115);
xor U12890 (N_12890,N_12283,N_12223);
nor U12891 (N_12891,N_12438,N_12102);
nand U12892 (N_12892,N_12366,N_12400);
xnor U12893 (N_12893,N_12507,N_12153);
nor U12894 (N_12894,N_12705,N_12498);
xnor U12895 (N_12895,N_12485,N_12622);
or U12896 (N_12896,N_12667,N_12331);
or U12897 (N_12897,N_12426,N_12521);
and U12898 (N_12898,N_12780,N_12117);
xor U12899 (N_12899,N_12671,N_12536);
nand U12900 (N_12900,N_12396,N_12069);
or U12901 (N_12901,N_12539,N_12104);
nor U12902 (N_12902,N_12109,N_12441);
xnor U12903 (N_12903,N_12556,N_12772);
nand U12904 (N_12904,N_12269,N_12090);
and U12905 (N_12905,N_12458,N_12161);
nand U12906 (N_12906,N_12559,N_12359);
xor U12907 (N_12907,N_12154,N_12764);
xor U12908 (N_12908,N_12307,N_12430);
or U12909 (N_12909,N_12524,N_12035);
or U12910 (N_12910,N_12783,N_12151);
xnor U12911 (N_12911,N_12297,N_12012);
nor U12912 (N_12912,N_12240,N_12022);
and U12913 (N_12913,N_12460,N_12061);
nand U12914 (N_12914,N_12444,N_12428);
or U12915 (N_12915,N_12234,N_12553);
nor U12916 (N_12916,N_12381,N_12793);
and U12917 (N_12917,N_12170,N_12034);
nand U12918 (N_12918,N_12699,N_12582);
nor U12919 (N_12919,N_12306,N_12262);
nor U12920 (N_12920,N_12495,N_12758);
nand U12921 (N_12921,N_12016,N_12407);
and U12922 (N_12922,N_12387,N_12335);
nor U12923 (N_12923,N_12229,N_12230);
nor U12924 (N_12924,N_12191,N_12279);
and U12925 (N_12925,N_12557,N_12047);
or U12926 (N_12926,N_12160,N_12048);
nand U12927 (N_12927,N_12420,N_12749);
nor U12928 (N_12928,N_12787,N_12063);
xnor U12929 (N_12929,N_12742,N_12626);
and U12930 (N_12930,N_12019,N_12415);
nand U12931 (N_12931,N_12776,N_12767);
nand U12932 (N_12932,N_12436,N_12106);
nor U12933 (N_12933,N_12572,N_12452);
nand U12934 (N_12934,N_12733,N_12484);
and U12935 (N_12935,N_12795,N_12394);
nand U12936 (N_12936,N_12455,N_12236);
nand U12937 (N_12937,N_12120,N_12459);
xor U12938 (N_12938,N_12379,N_12055);
nand U12939 (N_12939,N_12583,N_12654);
nor U12940 (N_12940,N_12207,N_12368);
xnor U12941 (N_12941,N_12159,N_12137);
and U12942 (N_12942,N_12725,N_12711);
nor U12943 (N_12943,N_12259,N_12642);
xnor U12944 (N_12944,N_12040,N_12519);
nor U12945 (N_12945,N_12488,N_12166);
xnor U12946 (N_12946,N_12062,N_12454);
nand U12947 (N_12947,N_12111,N_12530);
or U12948 (N_12948,N_12303,N_12666);
or U12949 (N_12949,N_12480,N_12756);
xor U12950 (N_12950,N_12706,N_12363);
xor U12951 (N_12951,N_12172,N_12361);
or U12952 (N_12952,N_12785,N_12215);
xor U12953 (N_12953,N_12774,N_12045);
or U12954 (N_12954,N_12332,N_12112);
nand U12955 (N_12955,N_12476,N_12470);
and U12956 (N_12956,N_12550,N_12348);
nor U12957 (N_12957,N_12571,N_12188);
or U12958 (N_12958,N_12508,N_12746);
and U12959 (N_12959,N_12634,N_12648);
nand U12960 (N_12960,N_12416,N_12757);
nand U12961 (N_12961,N_12714,N_12453);
nand U12962 (N_12962,N_12517,N_12251);
xor U12963 (N_12963,N_12391,N_12472);
nor U12964 (N_12964,N_12077,N_12761);
nor U12965 (N_12965,N_12082,N_12114);
nand U12966 (N_12966,N_12610,N_12630);
nor U12967 (N_12967,N_12128,N_12334);
nand U12968 (N_12968,N_12427,N_12378);
and U12969 (N_12969,N_12321,N_12021);
xor U12970 (N_12970,N_12652,N_12140);
and U12971 (N_12971,N_12253,N_12350);
nor U12972 (N_12972,N_12752,N_12718);
nor U12973 (N_12973,N_12250,N_12678);
nor U12974 (N_12974,N_12475,N_12197);
and U12975 (N_12975,N_12445,N_12411);
nor U12976 (N_12976,N_12032,N_12133);
xnor U12977 (N_12977,N_12177,N_12008);
and U12978 (N_12978,N_12268,N_12292);
nand U12979 (N_12979,N_12313,N_12672);
and U12980 (N_12980,N_12093,N_12218);
nand U12981 (N_12981,N_12701,N_12528);
nor U12982 (N_12982,N_12463,N_12466);
nor U12983 (N_12983,N_12238,N_12564);
and U12984 (N_12984,N_12726,N_12011);
xor U12985 (N_12985,N_12375,N_12717);
xor U12986 (N_12986,N_12272,N_12401);
and U12987 (N_12987,N_12351,N_12595);
xnor U12988 (N_12988,N_12339,N_12002);
and U12989 (N_12989,N_12057,N_12651);
and U12990 (N_12990,N_12258,N_12547);
nor U12991 (N_12991,N_12419,N_12766);
or U12992 (N_12992,N_12353,N_12053);
xnor U12993 (N_12993,N_12433,N_12078);
nor U12994 (N_12994,N_12636,N_12525);
or U12995 (N_12995,N_12374,N_12064);
nor U12996 (N_12996,N_12244,N_12447);
nand U12997 (N_12997,N_12431,N_12341);
xor U12998 (N_12998,N_12732,N_12156);
xnor U12999 (N_12999,N_12782,N_12222);
or U13000 (N_13000,N_12314,N_12205);
and U13001 (N_13001,N_12081,N_12096);
nand U13002 (N_13002,N_12645,N_12604);
nor U13003 (N_13003,N_12668,N_12171);
nor U13004 (N_13004,N_12540,N_12043);
xor U13005 (N_13005,N_12799,N_12639);
and U13006 (N_13006,N_12372,N_12257);
and U13007 (N_13007,N_12006,N_12769);
nor U13008 (N_13008,N_12263,N_12065);
nor U13009 (N_13009,N_12619,N_12054);
nor U13010 (N_13010,N_12390,N_12551);
xor U13011 (N_13011,N_12009,N_12033);
nor U13012 (N_13012,N_12183,N_12169);
nor U13013 (N_13013,N_12203,N_12039);
nor U13014 (N_13014,N_12301,N_12080);
nand U13015 (N_13015,N_12165,N_12256);
nand U13016 (N_13016,N_12763,N_12513);
or U13017 (N_13017,N_12603,N_12270);
xnor U13018 (N_13018,N_12435,N_12684);
nor U13019 (N_13019,N_12189,N_12481);
xor U13020 (N_13020,N_12070,N_12724);
or U13021 (N_13021,N_12038,N_12692);
or U13022 (N_13022,N_12580,N_12745);
xor U13023 (N_13023,N_12278,N_12185);
nor U13024 (N_13024,N_12336,N_12095);
nor U13025 (N_13025,N_12590,N_12058);
and U13026 (N_13026,N_12598,N_12237);
and U13027 (N_13027,N_12576,N_12105);
nor U13028 (N_13028,N_12158,N_12509);
nand U13029 (N_13029,N_12534,N_12195);
or U13030 (N_13030,N_12290,N_12627);
or U13031 (N_13031,N_12702,N_12024);
xor U13032 (N_13032,N_12318,N_12157);
nor U13033 (N_13033,N_12142,N_12386);
or U13034 (N_13034,N_12562,N_12349);
xor U13035 (N_13035,N_12228,N_12125);
nor U13036 (N_13036,N_12584,N_12134);
and U13037 (N_13037,N_12176,N_12554);
xor U13038 (N_13038,N_12743,N_12653);
nand U13039 (N_13039,N_12641,N_12333);
and U13040 (N_13040,N_12589,N_12629);
xnor U13041 (N_13041,N_12252,N_12592);
nor U13042 (N_13042,N_12028,N_12621);
nor U13043 (N_13043,N_12740,N_12298);
nor U13044 (N_13044,N_12669,N_12649);
or U13045 (N_13045,N_12760,N_12338);
or U13046 (N_13046,N_12255,N_12526);
nor U13047 (N_13047,N_12577,N_12730);
xor U13048 (N_13048,N_12074,N_12337);
and U13049 (N_13049,N_12144,N_12015);
nor U13050 (N_13050,N_12599,N_12587);
xor U13051 (N_13051,N_12204,N_12650);
and U13052 (N_13052,N_12103,N_12317);
or U13053 (N_13053,N_12052,N_12327);
and U13054 (N_13054,N_12687,N_12036);
and U13055 (N_13055,N_12690,N_12656);
xor U13056 (N_13056,N_12425,N_12477);
and U13057 (N_13057,N_12037,N_12182);
nor U13058 (N_13058,N_12108,N_12367);
nor U13059 (N_13059,N_12010,N_12685);
and U13060 (N_13060,N_12305,N_12432);
and U13061 (N_13061,N_12679,N_12249);
and U13062 (N_13062,N_12116,N_12007);
and U13063 (N_13063,N_12492,N_12496);
nand U13064 (N_13064,N_12541,N_12152);
and U13065 (N_13065,N_12091,N_12414);
and U13066 (N_13066,N_12285,N_12136);
nand U13067 (N_13067,N_12088,N_12319);
xnor U13068 (N_13068,N_12461,N_12383);
xnor U13069 (N_13069,N_12529,N_12049);
or U13070 (N_13070,N_12683,N_12267);
nand U13071 (N_13071,N_12013,N_12469);
nand U13072 (N_13072,N_12178,N_12403);
nand U13073 (N_13073,N_12199,N_12573);
and U13074 (N_13074,N_12710,N_12594);
or U13075 (N_13075,N_12275,N_12624);
nand U13076 (N_13076,N_12164,N_12499);
or U13077 (N_13077,N_12605,N_12190);
nor U13078 (N_13078,N_12597,N_12753);
or U13079 (N_13079,N_12232,N_12708);
or U13080 (N_13080,N_12465,N_12119);
or U13081 (N_13081,N_12186,N_12280);
and U13082 (N_13082,N_12122,N_12545);
xor U13083 (N_13083,N_12284,N_12409);
nor U13084 (N_13084,N_12729,N_12003);
and U13085 (N_13085,N_12092,N_12516);
xnor U13086 (N_13086,N_12243,N_12691);
nor U13087 (N_13087,N_12777,N_12004);
nor U13088 (N_13088,N_12451,N_12377);
or U13089 (N_13089,N_12309,N_12748);
and U13090 (N_13090,N_12184,N_12548);
and U13091 (N_13091,N_12625,N_12388);
and U13092 (N_13092,N_12789,N_12342);
nand U13093 (N_13093,N_12709,N_12471);
and U13094 (N_13094,N_12467,N_12071);
or U13095 (N_13095,N_12417,N_12099);
or U13096 (N_13096,N_12023,N_12288);
or U13097 (N_13097,N_12697,N_12633);
or U13098 (N_13098,N_12241,N_12788);
xnor U13099 (N_13099,N_12343,N_12751);
nor U13100 (N_13100,N_12385,N_12020);
nand U13101 (N_13101,N_12347,N_12716);
xnor U13102 (N_13102,N_12059,N_12792);
nor U13103 (N_13103,N_12737,N_12050);
and U13104 (N_13104,N_12585,N_12312);
or U13105 (N_13105,N_12179,N_12399);
or U13106 (N_13106,N_12212,N_12693);
and U13107 (N_13107,N_12031,N_12555);
xor U13108 (N_13108,N_12512,N_12311);
nand U13109 (N_13109,N_12124,N_12316);
nor U13110 (N_13110,N_12680,N_12219);
nor U13111 (N_13111,N_12442,N_12389);
nand U13112 (N_13112,N_12424,N_12593);
nor U13113 (N_13113,N_12382,N_12187);
or U13114 (N_13114,N_12616,N_12287);
nor U13115 (N_13115,N_12274,N_12110);
nor U13116 (N_13116,N_12617,N_12060);
and U13117 (N_13117,N_12632,N_12739);
and U13118 (N_13118,N_12771,N_12413);
or U13119 (N_13119,N_12659,N_12143);
nand U13120 (N_13120,N_12794,N_12479);
or U13121 (N_13121,N_12563,N_12696);
nor U13122 (N_13122,N_12356,N_12216);
nor U13123 (N_13123,N_12079,N_12354);
nand U13124 (N_13124,N_12588,N_12505);
xor U13125 (N_13125,N_12779,N_12500);
nand U13126 (N_13126,N_12744,N_12520);
and U13127 (N_13127,N_12225,N_12781);
and U13128 (N_13128,N_12468,N_12397);
or U13129 (N_13129,N_12502,N_12360);
xnor U13130 (N_13130,N_12660,N_12405);
or U13131 (N_13131,N_12402,N_12075);
and U13132 (N_13132,N_12736,N_12601);
xor U13133 (N_13133,N_12631,N_12473);
nand U13134 (N_13134,N_12193,N_12600);
and U13135 (N_13135,N_12490,N_12664);
nor U13136 (N_13136,N_12741,N_12640);
nand U13137 (N_13137,N_12412,N_12410);
and U13138 (N_13138,N_12421,N_12163);
nand U13139 (N_13139,N_12299,N_12514);
nand U13140 (N_13140,N_12345,N_12127);
nor U13141 (N_13141,N_12418,N_12084);
xor U13142 (N_13142,N_12073,N_12358);
or U13143 (N_13143,N_12107,N_12612);
and U13144 (N_13144,N_12014,N_12150);
nor U13145 (N_13145,N_12097,N_12765);
nor U13146 (N_13146,N_12294,N_12544);
xor U13147 (N_13147,N_12132,N_12644);
or U13148 (N_13148,N_12489,N_12775);
xor U13149 (N_13149,N_12790,N_12735);
and U13150 (N_13150,N_12000,N_12340);
or U13151 (N_13151,N_12239,N_12506);
or U13152 (N_13152,N_12643,N_12155);
xnor U13153 (N_13153,N_12086,N_12194);
xnor U13154 (N_13154,N_12248,N_12694);
xnor U13155 (N_13155,N_12217,N_12227);
and U13156 (N_13156,N_12712,N_12330);
nor U13157 (N_13157,N_12067,N_12167);
nor U13158 (N_13158,N_12017,N_12282);
nand U13159 (N_13159,N_12566,N_12762);
xnor U13160 (N_13160,N_12398,N_12535);
or U13161 (N_13161,N_12129,N_12574);
xnor U13162 (N_13162,N_12273,N_12056);
and U13163 (N_13163,N_12198,N_12613);
nor U13164 (N_13164,N_12260,N_12734);
nor U13165 (N_13165,N_12662,N_12100);
xor U13166 (N_13166,N_12720,N_12202);
and U13167 (N_13167,N_12226,N_12784);
and U13168 (N_13168,N_12113,N_12042);
xnor U13169 (N_13169,N_12707,N_12759);
nor U13170 (N_13170,N_12135,N_12731);
or U13171 (N_13171,N_12655,N_12373);
nor U13172 (N_13172,N_12393,N_12546);
and U13173 (N_13173,N_12510,N_12323);
or U13174 (N_13174,N_12578,N_12713);
or U13175 (N_13175,N_12208,N_12522);
nor U13176 (N_13176,N_12570,N_12628);
nand U13177 (N_13177,N_12698,N_12750);
nor U13178 (N_13178,N_12121,N_12098);
and U13179 (N_13179,N_12265,N_12542);
or U13180 (N_13180,N_12676,N_12308);
or U13181 (N_13181,N_12266,N_12677);
nand U13182 (N_13182,N_12596,N_12721);
or U13183 (N_13183,N_12670,N_12320);
nor U13184 (N_13184,N_12247,N_12423);
and U13185 (N_13185,N_12661,N_12196);
and U13186 (N_13186,N_12346,N_12201);
or U13187 (N_13187,N_12352,N_12174);
or U13188 (N_13188,N_12005,N_12213);
nand U13189 (N_13189,N_12286,N_12532);
nand U13190 (N_13190,N_12443,N_12501);
xor U13191 (N_13191,N_12450,N_12344);
nand U13192 (N_13192,N_12581,N_12324);
and U13193 (N_13193,N_12027,N_12291);
nand U13194 (N_13194,N_12376,N_12233);
xnor U13195 (N_13195,N_12235,N_12478);
nand U13196 (N_13196,N_12796,N_12531);
xor U13197 (N_13197,N_12560,N_12615);
nand U13198 (N_13198,N_12715,N_12175);
nor U13199 (N_13199,N_12408,N_12549);
and U13200 (N_13200,N_12044,N_12481);
nand U13201 (N_13201,N_12013,N_12477);
nor U13202 (N_13202,N_12001,N_12219);
xor U13203 (N_13203,N_12451,N_12260);
nand U13204 (N_13204,N_12173,N_12459);
nor U13205 (N_13205,N_12692,N_12540);
and U13206 (N_13206,N_12467,N_12691);
or U13207 (N_13207,N_12513,N_12161);
and U13208 (N_13208,N_12227,N_12196);
xnor U13209 (N_13209,N_12795,N_12111);
nand U13210 (N_13210,N_12783,N_12303);
nand U13211 (N_13211,N_12173,N_12326);
nand U13212 (N_13212,N_12374,N_12452);
xor U13213 (N_13213,N_12186,N_12523);
or U13214 (N_13214,N_12614,N_12458);
or U13215 (N_13215,N_12327,N_12368);
and U13216 (N_13216,N_12684,N_12718);
or U13217 (N_13217,N_12402,N_12568);
nor U13218 (N_13218,N_12498,N_12659);
nor U13219 (N_13219,N_12314,N_12537);
or U13220 (N_13220,N_12568,N_12315);
xnor U13221 (N_13221,N_12065,N_12770);
xnor U13222 (N_13222,N_12523,N_12512);
nor U13223 (N_13223,N_12485,N_12004);
and U13224 (N_13224,N_12498,N_12779);
or U13225 (N_13225,N_12299,N_12266);
xnor U13226 (N_13226,N_12177,N_12301);
and U13227 (N_13227,N_12508,N_12050);
nor U13228 (N_13228,N_12229,N_12219);
nand U13229 (N_13229,N_12795,N_12258);
nand U13230 (N_13230,N_12210,N_12236);
nand U13231 (N_13231,N_12364,N_12469);
nand U13232 (N_13232,N_12650,N_12646);
nand U13233 (N_13233,N_12539,N_12448);
xnor U13234 (N_13234,N_12701,N_12491);
or U13235 (N_13235,N_12107,N_12163);
and U13236 (N_13236,N_12341,N_12592);
nand U13237 (N_13237,N_12076,N_12758);
nor U13238 (N_13238,N_12713,N_12096);
or U13239 (N_13239,N_12080,N_12231);
xnor U13240 (N_13240,N_12205,N_12412);
nor U13241 (N_13241,N_12037,N_12277);
nor U13242 (N_13242,N_12503,N_12219);
xnor U13243 (N_13243,N_12168,N_12143);
nand U13244 (N_13244,N_12659,N_12174);
or U13245 (N_13245,N_12339,N_12037);
xor U13246 (N_13246,N_12742,N_12026);
xor U13247 (N_13247,N_12139,N_12423);
nor U13248 (N_13248,N_12497,N_12572);
and U13249 (N_13249,N_12347,N_12092);
xnor U13250 (N_13250,N_12376,N_12577);
nor U13251 (N_13251,N_12508,N_12411);
or U13252 (N_13252,N_12389,N_12419);
nand U13253 (N_13253,N_12746,N_12006);
nand U13254 (N_13254,N_12165,N_12667);
or U13255 (N_13255,N_12080,N_12050);
nand U13256 (N_13256,N_12320,N_12621);
nand U13257 (N_13257,N_12472,N_12332);
xor U13258 (N_13258,N_12032,N_12492);
or U13259 (N_13259,N_12690,N_12422);
and U13260 (N_13260,N_12522,N_12749);
or U13261 (N_13261,N_12396,N_12425);
nor U13262 (N_13262,N_12075,N_12495);
or U13263 (N_13263,N_12706,N_12451);
and U13264 (N_13264,N_12499,N_12272);
and U13265 (N_13265,N_12751,N_12649);
nand U13266 (N_13266,N_12000,N_12024);
xnor U13267 (N_13267,N_12569,N_12225);
nand U13268 (N_13268,N_12317,N_12779);
xor U13269 (N_13269,N_12311,N_12624);
nand U13270 (N_13270,N_12122,N_12476);
nor U13271 (N_13271,N_12156,N_12139);
nand U13272 (N_13272,N_12644,N_12471);
or U13273 (N_13273,N_12747,N_12446);
xor U13274 (N_13274,N_12391,N_12166);
nor U13275 (N_13275,N_12547,N_12398);
or U13276 (N_13276,N_12063,N_12472);
or U13277 (N_13277,N_12128,N_12457);
xor U13278 (N_13278,N_12657,N_12531);
nand U13279 (N_13279,N_12136,N_12326);
and U13280 (N_13280,N_12316,N_12728);
or U13281 (N_13281,N_12587,N_12376);
xor U13282 (N_13282,N_12060,N_12024);
xor U13283 (N_13283,N_12069,N_12185);
nand U13284 (N_13284,N_12449,N_12020);
nand U13285 (N_13285,N_12074,N_12305);
and U13286 (N_13286,N_12010,N_12049);
or U13287 (N_13287,N_12750,N_12462);
nor U13288 (N_13288,N_12578,N_12482);
xnor U13289 (N_13289,N_12171,N_12239);
xnor U13290 (N_13290,N_12623,N_12448);
nor U13291 (N_13291,N_12768,N_12401);
xnor U13292 (N_13292,N_12298,N_12048);
nand U13293 (N_13293,N_12157,N_12642);
nand U13294 (N_13294,N_12626,N_12528);
or U13295 (N_13295,N_12681,N_12224);
xor U13296 (N_13296,N_12658,N_12413);
xnor U13297 (N_13297,N_12081,N_12632);
and U13298 (N_13298,N_12210,N_12270);
nand U13299 (N_13299,N_12590,N_12466);
and U13300 (N_13300,N_12481,N_12565);
nor U13301 (N_13301,N_12660,N_12731);
nand U13302 (N_13302,N_12444,N_12487);
nor U13303 (N_13303,N_12450,N_12635);
or U13304 (N_13304,N_12157,N_12127);
nand U13305 (N_13305,N_12147,N_12462);
and U13306 (N_13306,N_12689,N_12263);
and U13307 (N_13307,N_12085,N_12062);
or U13308 (N_13308,N_12095,N_12683);
nor U13309 (N_13309,N_12488,N_12098);
nand U13310 (N_13310,N_12567,N_12542);
nand U13311 (N_13311,N_12286,N_12723);
nand U13312 (N_13312,N_12535,N_12112);
xnor U13313 (N_13313,N_12254,N_12327);
nor U13314 (N_13314,N_12462,N_12622);
xor U13315 (N_13315,N_12452,N_12061);
nor U13316 (N_13316,N_12263,N_12640);
xor U13317 (N_13317,N_12172,N_12363);
nand U13318 (N_13318,N_12313,N_12056);
nand U13319 (N_13319,N_12648,N_12376);
nor U13320 (N_13320,N_12689,N_12150);
nor U13321 (N_13321,N_12230,N_12776);
or U13322 (N_13322,N_12772,N_12560);
or U13323 (N_13323,N_12503,N_12535);
and U13324 (N_13324,N_12664,N_12386);
or U13325 (N_13325,N_12570,N_12748);
nand U13326 (N_13326,N_12170,N_12704);
or U13327 (N_13327,N_12580,N_12434);
nor U13328 (N_13328,N_12741,N_12442);
xor U13329 (N_13329,N_12474,N_12048);
nor U13330 (N_13330,N_12334,N_12612);
nor U13331 (N_13331,N_12497,N_12646);
nand U13332 (N_13332,N_12286,N_12799);
or U13333 (N_13333,N_12106,N_12627);
and U13334 (N_13334,N_12458,N_12566);
xor U13335 (N_13335,N_12397,N_12751);
nand U13336 (N_13336,N_12220,N_12091);
nand U13337 (N_13337,N_12068,N_12298);
nor U13338 (N_13338,N_12492,N_12070);
nor U13339 (N_13339,N_12670,N_12060);
xnor U13340 (N_13340,N_12285,N_12336);
nand U13341 (N_13341,N_12520,N_12093);
xnor U13342 (N_13342,N_12773,N_12238);
or U13343 (N_13343,N_12394,N_12562);
and U13344 (N_13344,N_12396,N_12599);
xnor U13345 (N_13345,N_12216,N_12486);
nor U13346 (N_13346,N_12680,N_12582);
and U13347 (N_13347,N_12020,N_12029);
nor U13348 (N_13348,N_12270,N_12178);
nor U13349 (N_13349,N_12708,N_12038);
xnor U13350 (N_13350,N_12503,N_12411);
nor U13351 (N_13351,N_12062,N_12519);
nor U13352 (N_13352,N_12376,N_12526);
nand U13353 (N_13353,N_12203,N_12622);
nor U13354 (N_13354,N_12420,N_12589);
xor U13355 (N_13355,N_12575,N_12246);
and U13356 (N_13356,N_12072,N_12637);
nor U13357 (N_13357,N_12454,N_12276);
nand U13358 (N_13358,N_12120,N_12521);
xor U13359 (N_13359,N_12308,N_12703);
nor U13360 (N_13360,N_12696,N_12264);
and U13361 (N_13361,N_12182,N_12283);
xnor U13362 (N_13362,N_12583,N_12749);
nand U13363 (N_13363,N_12218,N_12447);
nor U13364 (N_13364,N_12203,N_12183);
xor U13365 (N_13365,N_12159,N_12585);
and U13366 (N_13366,N_12452,N_12552);
xnor U13367 (N_13367,N_12329,N_12723);
or U13368 (N_13368,N_12717,N_12697);
and U13369 (N_13369,N_12678,N_12095);
or U13370 (N_13370,N_12137,N_12534);
nand U13371 (N_13371,N_12092,N_12597);
nand U13372 (N_13372,N_12691,N_12061);
nor U13373 (N_13373,N_12345,N_12787);
or U13374 (N_13374,N_12522,N_12752);
nor U13375 (N_13375,N_12299,N_12697);
xnor U13376 (N_13376,N_12555,N_12643);
or U13377 (N_13377,N_12709,N_12680);
nand U13378 (N_13378,N_12213,N_12413);
and U13379 (N_13379,N_12799,N_12755);
xor U13380 (N_13380,N_12407,N_12708);
nor U13381 (N_13381,N_12739,N_12793);
xor U13382 (N_13382,N_12635,N_12614);
nand U13383 (N_13383,N_12690,N_12509);
xor U13384 (N_13384,N_12242,N_12677);
or U13385 (N_13385,N_12168,N_12299);
or U13386 (N_13386,N_12277,N_12126);
nand U13387 (N_13387,N_12090,N_12668);
and U13388 (N_13388,N_12091,N_12186);
nand U13389 (N_13389,N_12775,N_12328);
xnor U13390 (N_13390,N_12532,N_12183);
xor U13391 (N_13391,N_12242,N_12585);
xnor U13392 (N_13392,N_12013,N_12380);
nand U13393 (N_13393,N_12434,N_12799);
xnor U13394 (N_13394,N_12381,N_12262);
or U13395 (N_13395,N_12662,N_12304);
xnor U13396 (N_13396,N_12239,N_12323);
or U13397 (N_13397,N_12185,N_12569);
nand U13398 (N_13398,N_12381,N_12617);
and U13399 (N_13399,N_12783,N_12403);
xnor U13400 (N_13400,N_12144,N_12370);
nor U13401 (N_13401,N_12218,N_12281);
nor U13402 (N_13402,N_12157,N_12261);
and U13403 (N_13403,N_12668,N_12368);
nor U13404 (N_13404,N_12189,N_12249);
nand U13405 (N_13405,N_12413,N_12271);
and U13406 (N_13406,N_12356,N_12133);
nand U13407 (N_13407,N_12309,N_12146);
nor U13408 (N_13408,N_12282,N_12636);
nor U13409 (N_13409,N_12250,N_12713);
nor U13410 (N_13410,N_12567,N_12564);
nand U13411 (N_13411,N_12350,N_12155);
and U13412 (N_13412,N_12634,N_12793);
nand U13413 (N_13413,N_12336,N_12164);
nor U13414 (N_13414,N_12775,N_12601);
or U13415 (N_13415,N_12555,N_12101);
xor U13416 (N_13416,N_12013,N_12621);
nand U13417 (N_13417,N_12601,N_12413);
nand U13418 (N_13418,N_12046,N_12732);
nor U13419 (N_13419,N_12285,N_12775);
xnor U13420 (N_13420,N_12342,N_12205);
xnor U13421 (N_13421,N_12544,N_12573);
nand U13422 (N_13422,N_12447,N_12616);
and U13423 (N_13423,N_12473,N_12407);
nor U13424 (N_13424,N_12325,N_12560);
and U13425 (N_13425,N_12265,N_12755);
and U13426 (N_13426,N_12194,N_12370);
nand U13427 (N_13427,N_12301,N_12514);
nor U13428 (N_13428,N_12731,N_12500);
or U13429 (N_13429,N_12622,N_12210);
nor U13430 (N_13430,N_12604,N_12352);
nand U13431 (N_13431,N_12346,N_12034);
and U13432 (N_13432,N_12008,N_12577);
and U13433 (N_13433,N_12699,N_12235);
and U13434 (N_13434,N_12727,N_12508);
or U13435 (N_13435,N_12454,N_12300);
and U13436 (N_13436,N_12154,N_12477);
or U13437 (N_13437,N_12648,N_12382);
and U13438 (N_13438,N_12460,N_12133);
nand U13439 (N_13439,N_12242,N_12599);
nand U13440 (N_13440,N_12075,N_12042);
or U13441 (N_13441,N_12736,N_12190);
or U13442 (N_13442,N_12272,N_12385);
and U13443 (N_13443,N_12093,N_12631);
nor U13444 (N_13444,N_12226,N_12169);
xnor U13445 (N_13445,N_12295,N_12104);
or U13446 (N_13446,N_12236,N_12191);
nor U13447 (N_13447,N_12490,N_12670);
and U13448 (N_13448,N_12206,N_12468);
xor U13449 (N_13449,N_12359,N_12344);
and U13450 (N_13450,N_12197,N_12021);
or U13451 (N_13451,N_12556,N_12555);
nor U13452 (N_13452,N_12462,N_12547);
nand U13453 (N_13453,N_12337,N_12122);
nand U13454 (N_13454,N_12589,N_12657);
xor U13455 (N_13455,N_12756,N_12107);
nand U13456 (N_13456,N_12031,N_12068);
and U13457 (N_13457,N_12220,N_12525);
or U13458 (N_13458,N_12491,N_12670);
nor U13459 (N_13459,N_12763,N_12268);
nand U13460 (N_13460,N_12499,N_12037);
and U13461 (N_13461,N_12181,N_12054);
nor U13462 (N_13462,N_12738,N_12257);
or U13463 (N_13463,N_12633,N_12134);
and U13464 (N_13464,N_12540,N_12517);
xor U13465 (N_13465,N_12298,N_12798);
nand U13466 (N_13466,N_12128,N_12721);
or U13467 (N_13467,N_12364,N_12216);
xnor U13468 (N_13468,N_12576,N_12155);
nand U13469 (N_13469,N_12307,N_12798);
nand U13470 (N_13470,N_12592,N_12655);
nand U13471 (N_13471,N_12424,N_12664);
nor U13472 (N_13472,N_12657,N_12112);
xor U13473 (N_13473,N_12194,N_12374);
nand U13474 (N_13474,N_12381,N_12790);
nand U13475 (N_13475,N_12437,N_12341);
xnor U13476 (N_13476,N_12683,N_12742);
or U13477 (N_13477,N_12625,N_12248);
or U13478 (N_13478,N_12039,N_12467);
xor U13479 (N_13479,N_12562,N_12043);
or U13480 (N_13480,N_12539,N_12786);
xnor U13481 (N_13481,N_12404,N_12551);
nand U13482 (N_13482,N_12317,N_12404);
nand U13483 (N_13483,N_12711,N_12400);
xor U13484 (N_13484,N_12136,N_12590);
nor U13485 (N_13485,N_12439,N_12360);
xor U13486 (N_13486,N_12147,N_12206);
xor U13487 (N_13487,N_12560,N_12025);
or U13488 (N_13488,N_12188,N_12239);
nand U13489 (N_13489,N_12796,N_12002);
or U13490 (N_13490,N_12317,N_12018);
or U13491 (N_13491,N_12645,N_12717);
nor U13492 (N_13492,N_12304,N_12298);
xnor U13493 (N_13493,N_12081,N_12391);
or U13494 (N_13494,N_12204,N_12365);
nand U13495 (N_13495,N_12332,N_12623);
xnor U13496 (N_13496,N_12754,N_12082);
xnor U13497 (N_13497,N_12341,N_12543);
nor U13498 (N_13498,N_12013,N_12766);
xnor U13499 (N_13499,N_12482,N_12173);
or U13500 (N_13500,N_12449,N_12436);
xor U13501 (N_13501,N_12028,N_12689);
and U13502 (N_13502,N_12739,N_12105);
or U13503 (N_13503,N_12648,N_12258);
nor U13504 (N_13504,N_12617,N_12288);
xnor U13505 (N_13505,N_12341,N_12471);
nand U13506 (N_13506,N_12312,N_12447);
nand U13507 (N_13507,N_12716,N_12797);
nand U13508 (N_13508,N_12180,N_12682);
and U13509 (N_13509,N_12404,N_12291);
and U13510 (N_13510,N_12098,N_12733);
xnor U13511 (N_13511,N_12066,N_12698);
nor U13512 (N_13512,N_12641,N_12594);
xnor U13513 (N_13513,N_12072,N_12688);
or U13514 (N_13514,N_12502,N_12742);
xnor U13515 (N_13515,N_12737,N_12425);
or U13516 (N_13516,N_12381,N_12541);
and U13517 (N_13517,N_12262,N_12785);
or U13518 (N_13518,N_12294,N_12146);
xnor U13519 (N_13519,N_12777,N_12760);
xnor U13520 (N_13520,N_12296,N_12010);
nand U13521 (N_13521,N_12028,N_12762);
nor U13522 (N_13522,N_12243,N_12432);
xnor U13523 (N_13523,N_12693,N_12749);
xnor U13524 (N_13524,N_12731,N_12779);
and U13525 (N_13525,N_12377,N_12557);
xor U13526 (N_13526,N_12781,N_12093);
nand U13527 (N_13527,N_12772,N_12463);
nand U13528 (N_13528,N_12174,N_12270);
or U13529 (N_13529,N_12598,N_12266);
and U13530 (N_13530,N_12129,N_12465);
nand U13531 (N_13531,N_12100,N_12019);
xnor U13532 (N_13532,N_12393,N_12519);
nor U13533 (N_13533,N_12627,N_12112);
nor U13534 (N_13534,N_12575,N_12684);
and U13535 (N_13535,N_12716,N_12475);
xor U13536 (N_13536,N_12147,N_12048);
and U13537 (N_13537,N_12548,N_12076);
nand U13538 (N_13538,N_12675,N_12344);
or U13539 (N_13539,N_12580,N_12189);
xor U13540 (N_13540,N_12051,N_12484);
xor U13541 (N_13541,N_12026,N_12257);
and U13542 (N_13542,N_12763,N_12662);
or U13543 (N_13543,N_12005,N_12256);
or U13544 (N_13544,N_12305,N_12164);
and U13545 (N_13545,N_12109,N_12415);
nand U13546 (N_13546,N_12658,N_12728);
xor U13547 (N_13547,N_12378,N_12719);
and U13548 (N_13548,N_12791,N_12691);
and U13549 (N_13549,N_12799,N_12514);
nand U13550 (N_13550,N_12445,N_12750);
or U13551 (N_13551,N_12180,N_12731);
nor U13552 (N_13552,N_12760,N_12060);
xor U13553 (N_13553,N_12298,N_12633);
xnor U13554 (N_13554,N_12036,N_12243);
xor U13555 (N_13555,N_12667,N_12018);
nand U13556 (N_13556,N_12242,N_12257);
and U13557 (N_13557,N_12563,N_12741);
nand U13558 (N_13558,N_12388,N_12005);
nor U13559 (N_13559,N_12532,N_12702);
xnor U13560 (N_13560,N_12491,N_12577);
nor U13561 (N_13561,N_12098,N_12467);
xor U13562 (N_13562,N_12139,N_12286);
and U13563 (N_13563,N_12713,N_12635);
nand U13564 (N_13564,N_12216,N_12385);
and U13565 (N_13565,N_12101,N_12712);
and U13566 (N_13566,N_12203,N_12270);
nor U13567 (N_13567,N_12745,N_12255);
nand U13568 (N_13568,N_12416,N_12118);
nand U13569 (N_13569,N_12080,N_12514);
or U13570 (N_13570,N_12594,N_12650);
or U13571 (N_13571,N_12335,N_12002);
xor U13572 (N_13572,N_12495,N_12755);
xnor U13573 (N_13573,N_12232,N_12744);
nand U13574 (N_13574,N_12105,N_12341);
and U13575 (N_13575,N_12417,N_12798);
or U13576 (N_13576,N_12180,N_12617);
or U13577 (N_13577,N_12709,N_12510);
or U13578 (N_13578,N_12610,N_12334);
nor U13579 (N_13579,N_12089,N_12439);
nand U13580 (N_13580,N_12268,N_12097);
and U13581 (N_13581,N_12714,N_12258);
nand U13582 (N_13582,N_12733,N_12386);
nand U13583 (N_13583,N_12408,N_12140);
nor U13584 (N_13584,N_12257,N_12612);
and U13585 (N_13585,N_12417,N_12502);
nor U13586 (N_13586,N_12557,N_12553);
nor U13587 (N_13587,N_12530,N_12323);
nor U13588 (N_13588,N_12177,N_12522);
nand U13589 (N_13589,N_12289,N_12474);
xnor U13590 (N_13590,N_12030,N_12507);
and U13591 (N_13591,N_12231,N_12269);
and U13592 (N_13592,N_12203,N_12213);
or U13593 (N_13593,N_12416,N_12617);
xor U13594 (N_13594,N_12784,N_12033);
and U13595 (N_13595,N_12124,N_12381);
xnor U13596 (N_13596,N_12202,N_12534);
or U13597 (N_13597,N_12414,N_12611);
xnor U13598 (N_13598,N_12509,N_12377);
xor U13599 (N_13599,N_12407,N_12566);
nand U13600 (N_13600,N_13178,N_12812);
or U13601 (N_13601,N_12841,N_12995);
nor U13602 (N_13602,N_13057,N_13274);
and U13603 (N_13603,N_13070,N_13088);
nor U13604 (N_13604,N_13453,N_13023);
xnor U13605 (N_13605,N_13193,N_13579);
nand U13606 (N_13606,N_12899,N_12938);
or U13607 (N_13607,N_12910,N_13234);
and U13608 (N_13608,N_12956,N_13233);
and U13609 (N_13609,N_12907,N_13464);
and U13610 (N_13610,N_13498,N_12887);
nor U13611 (N_13611,N_13039,N_12829);
nand U13612 (N_13612,N_13374,N_13383);
nand U13613 (N_13613,N_13147,N_13034);
or U13614 (N_13614,N_13235,N_13211);
and U13615 (N_13615,N_13053,N_12916);
and U13616 (N_13616,N_12889,N_13093);
nor U13617 (N_13617,N_13550,N_13240);
xor U13618 (N_13618,N_13592,N_13359);
xor U13619 (N_13619,N_12953,N_13494);
and U13620 (N_13620,N_12882,N_12923);
and U13621 (N_13621,N_13575,N_13058);
nand U13622 (N_13622,N_13414,N_13185);
or U13623 (N_13623,N_13388,N_12984);
nand U13624 (N_13624,N_12885,N_13378);
nand U13625 (N_13625,N_13109,N_12978);
xnor U13626 (N_13626,N_12964,N_13462);
nand U13627 (N_13627,N_12981,N_13106);
nand U13628 (N_13628,N_12855,N_13283);
and U13629 (N_13629,N_13141,N_13294);
xnor U13630 (N_13630,N_13144,N_13328);
nand U13631 (N_13631,N_13167,N_13082);
xor U13632 (N_13632,N_13408,N_13430);
or U13633 (N_13633,N_13480,N_13543);
and U13634 (N_13634,N_13248,N_13124);
nor U13635 (N_13635,N_13073,N_12962);
nor U13636 (N_13636,N_12993,N_12965);
xor U13637 (N_13637,N_13570,N_13333);
xor U13638 (N_13638,N_12853,N_13249);
xnor U13639 (N_13639,N_13346,N_12818);
and U13640 (N_13640,N_13165,N_13561);
nor U13641 (N_13641,N_13028,N_13064);
nor U13642 (N_13642,N_13368,N_13020);
nor U13643 (N_13643,N_13369,N_13087);
and U13644 (N_13644,N_12991,N_12897);
nor U13645 (N_13645,N_13254,N_12821);
or U13646 (N_13646,N_13531,N_13499);
nand U13647 (N_13647,N_12846,N_13560);
xor U13648 (N_13648,N_13330,N_12968);
nand U13649 (N_13649,N_13176,N_13491);
nand U13650 (N_13650,N_13139,N_13195);
xnor U13651 (N_13651,N_13012,N_13025);
and U13652 (N_13652,N_12931,N_12982);
xor U13653 (N_13653,N_13126,N_13341);
and U13654 (N_13654,N_13246,N_13078);
or U13655 (N_13655,N_13018,N_13121);
and U13656 (N_13656,N_13594,N_13214);
nand U13657 (N_13657,N_13415,N_12972);
or U13658 (N_13658,N_12960,N_13492);
nor U13659 (N_13659,N_13559,N_13345);
nor U13660 (N_13660,N_13272,N_12876);
xnor U13661 (N_13661,N_13544,N_13514);
xnor U13662 (N_13662,N_13271,N_13596);
nand U13663 (N_13663,N_13143,N_13382);
xor U13664 (N_13664,N_13385,N_13405);
nor U13665 (N_13665,N_13479,N_13556);
and U13666 (N_13666,N_12918,N_13355);
nor U13667 (N_13667,N_13273,N_12800);
nor U13668 (N_13668,N_12936,N_13171);
or U13669 (N_13669,N_13392,N_13302);
xnor U13670 (N_13670,N_13452,N_13595);
xor U13671 (N_13671,N_12900,N_12950);
nor U13672 (N_13672,N_12831,N_13298);
or U13673 (N_13673,N_13091,N_13587);
xor U13674 (N_13674,N_13136,N_13542);
and U13675 (N_13675,N_13197,N_12961);
xor U13676 (N_13676,N_13243,N_12994);
nor U13677 (N_13677,N_13125,N_13068);
nor U13678 (N_13678,N_13004,N_13168);
xor U13679 (N_13679,N_13140,N_13473);
or U13680 (N_13680,N_13315,N_13558);
and U13681 (N_13681,N_13280,N_13072);
nor U13682 (N_13682,N_13324,N_13047);
and U13683 (N_13683,N_13554,N_13578);
xnor U13684 (N_13684,N_13376,N_13213);
and U13685 (N_13685,N_13201,N_13401);
xor U13686 (N_13686,N_13236,N_13276);
and U13687 (N_13687,N_13067,N_13005);
nor U13688 (N_13688,N_13353,N_13089);
or U13689 (N_13689,N_13375,N_13512);
nand U13690 (N_13690,N_13164,N_13112);
or U13691 (N_13691,N_13312,N_13119);
or U13692 (N_13692,N_13541,N_13299);
nor U13693 (N_13693,N_12830,N_13501);
nor U13694 (N_13694,N_12904,N_13268);
and U13695 (N_13695,N_12898,N_13242);
or U13696 (N_13696,N_12801,N_12838);
and U13697 (N_13697,N_12850,N_13557);
and U13698 (N_13698,N_13503,N_13520);
nand U13699 (N_13699,N_13253,N_13370);
xnor U13700 (N_13700,N_13244,N_12976);
nand U13701 (N_13701,N_13426,N_13413);
nand U13702 (N_13702,N_12934,N_13419);
and U13703 (N_13703,N_13535,N_13311);
and U13704 (N_13704,N_13526,N_13502);
or U13705 (N_13705,N_12975,N_13161);
or U13706 (N_13706,N_13154,N_13237);
or U13707 (N_13707,N_12822,N_13478);
nor U13708 (N_13708,N_12854,N_13371);
or U13709 (N_13709,N_13133,N_13245);
and U13710 (N_13710,N_13303,N_13270);
or U13711 (N_13711,N_13216,N_13313);
or U13712 (N_13712,N_12827,N_13349);
and U13713 (N_13713,N_13537,N_13517);
nand U13714 (N_13714,N_13116,N_12902);
or U13715 (N_13715,N_13577,N_12852);
nand U13716 (N_13716,N_12868,N_13493);
and U13717 (N_13717,N_12947,N_13040);
and U13718 (N_13718,N_13463,N_13555);
or U13719 (N_13719,N_13564,N_13580);
and U13720 (N_13720,N_12870,N_12840);
nor U13721 (N_13721,N_13122,N_13568);
nand U13722 (N_13722,N_12983,N_13460);
nand U13723 (N_13723,N_12939,N_12913);
nor U13724 (N_13724,N_13199,N_13402);
nand U13725 (N_13725,N_13000,N_13159);
and U13726 (N_13726,N_13200,N_13016);
nor U13727 (N_13727,N_13207,N_12871);
or U13728 (N_13728,N_13284,N_12941);
xnor U13729 (N_13729,N_13048,N_13196);
or U13730 (N_13730,N_12844,N_13033);
nor U13731 (N_13731,N_13467,N_13038);
xor U13732 (N_13732,N_13437,N_13425);
nand U13733 (N_13733,N_13314,N_12928);
xor U13734 (N_13734,N_13160,N_13008);
and U13735 (N_13735,N_12869,N_13525);
or U13736 (N_13736,N_12826,N_13098);
xor U13737 (N_13737,N_13574,N_13230);
or U13738 (N_13738,N_12967,N_12815);
and U13739 (N_13739,N_13186,N_13553);
and U13740 (N_13740,N_12839,N_12945);
nor U13741 (N_13741,N_13343,N_13538);
and U13742 (N_13742,N_13055,N_13552);
nor U13743 (N_13743,N_12903,N_13336);
nor U13744 (N_13744,N_13198,N_12988);
or U13745 (N_13745,N_12933,N_12864);
or U13746 (N_13746,N_13377,N_12863);
nand U13747 (N_13747,N_12861,N_13562);
or U13748 (N_13748,N_13316,N_13009);
and U13749 (N_13749,N_13340,N_13454);
nand U13750 (N_13750,N_13032,N_13044);
xnor U13751 (N_13751,N_13458,N_12865);
xor U13752 (N_13752,N_12894,N_13434);
xnor U13753 (N_13753,N_13476,N_12880);
nor U13754 (N_13754,N_13128,N_13412);
nand U13755 (N_13755,N_12985,N_13582);
and U13756 (N_13756,N_13471,N_12998);
or U13757 (N_13757,N_13361,N_13518);
xnor U13758 (N_13758,N_13086,N_13175);
nand U13759 (N_13759,N_13059,N_13002);
xnor U13760 (N_13760,N_13074,N_13468);
nand U13761 (N_13761,N_12872,N_13380);
nand U13762 (N_13762,N_13567,N_13267);
and U13763 (N_13763,N_13290,N_13540);
or U13764 (N_13764,N_13599,N_13507);
and U13765 (N_13765,N_13563,N_13096);
nand U13766 (N_13766,N_13591,N_13181);
or U13767 (N_13767,N_13046,N_13572);
and U13768 (N_13768,N_13351,N_13277);
nor U13769 (N_13769,N_13465,N_12929);
or U13770 (N_13770,N_13588,N_13417);
and U13771 (N_13771,N_13108,N_13505);
xnor U13772 (N_13772,N_13241,N_13151);
or U13773 (N_13773,N_13321,N_13327);
nor U13774 (N_13774,N_13508,N_13584);
and U13775 (N_13775,N_13305,N_13308);
xnor U13776 (N_13776,N_13451,N_13571);
or U13777 (N_13777,N_13118,N_12873);
or U13778 (N_13778,N_13352,N_13256);
or U13779 (N_13779,N_13338,N_13158);
or U13780 (N_13780,N_13206,N_13485);
nor U13781 (N_13781,N_12803,N_13566);
xor U13782 (N_13782,N_12859,N_12875);
nor U13783 (N_13783,N_13084,N_13329);
nand U13784 (N_13784,N_13372,N_13427);
and U13785 (N_13785,N_13325,N_13318);
and U13786 (N_13786,N_12959,N_13202);
nand U13787 (N_13787,N_13079,N_13569);
nand U13788 (N_13788,N_13062,N_13010);
nand U13789 (N_13789,N_13509,N_13483);
nor U13790 (N_13790,N_13285,N_13212);
and U13791 (N_13791,N_13429,N_13286);
nand U13792 (N_13792,N_13527,N_12977);
and U13793 (N_13793,N_13111,N_13477);
nand U13794 (N_13794,N_13042,N_13519);
xor U13795 (N_13795,N_13130,N_13344);
or U13796 (N_13796,N_13428,N_13386);
nor U13797 (N_13797,N_13162,N_13482);
xor U13798 (N_13798,N_12878,N_13061);
nand U13799 (N_13799,N_13472,N_13251);
or U13800 (N_13800,N_12808,N_13179);
nand U13801 (N_13801,N_13115,N_12908);
nor U13802 (N_13802,N_13443,N_13506);
and U13803 (N_13803,N_13598,N_13281);
nand U13804 (N_13804,N_13539,N_12817);
xor U13805 (N_13805,N_12819,N_13177);
nor U13806 (N_13806,N_12948,N_13263);
nor U13807 (N_13807,N_12834,N_13085);
xnor U13808 (N_13808,N_13152,N_12832);
nor U13809 (N_13809,N_13297,N_13049);
and U13810 (N_13810,N_13585,N_13306);
xnor U13811 (N_13811,N_13546,N_13037);
and U13812 (N_13812,N_12874,N_13100);
or U13813 (N_13813,N_13332,N_13204);
and U13814 (N_13814,N_13489,N_12946);
nor U13815 (N_13815,N_13586,N_13265);
nand U13816 (N_13816,N_13275,N_13365);
or U13817 (N_13817,N_13123,N_12940);
nand U13818 (N_13818,N_13228,N_13014);
xor U13819 (N_13819,N_13410,N_12997);
nand U13820 (N_13820,N_13229,N_13183);
xnor U13821 (N_13821,N_13250,N_12809);
and U13822 (N_13822,N_13384,N_12820);
and U13823 (N_13823,N_12858,N_12914);
nand U13824 (N_13824,N_13515,N_13225);
nand U13825 (N_13825,N_12892,N_13261);
and U13826 (N_13826,N_13455,N_13247);
nand U13827 (N_13827,N_13219,N_13348);
xor U13828 (N_13828,N_13565,N_13022);
nor U13829 (N_13829,N_13440,N_13120);
nor U13830 (N_13830,N_12963,N_13169);
nand U13831 (N_13831,N_13222,N_12802);
and U13832 (N_13832,N_13545,N_13192);
xor U13833 (N_13833,N_13232,N_13547);
nor U13834 (N_13834,N_13356,N_13013);
nand U13835 (N_13835,N_13105,N_13576);
xnor U13836 (N_13836,N_12806,N_13532);
nand U13837 (N_13837,N_13094,N_13409);
or U13838 (N_13838,N_13194,N_12805);
nand U13839 (N_13839,N_12987,N_13052);
and U13840 (N_13840,N_13036,N_12814);
nor U13841 (N_13841,N_13533,N_12906);
and U13842 (N_13842,N_13269,N_13069);
xor U13843 (N_13843,N_13031,N_13583);
nor U13844 (N_13844,N_13528,N_13357);
or U13845 (N_13845,N_13081,N_13593);
and U13846 (N_13846,N_12925,N_13347);
nand U13847 (N_13847,N_13404,N_13182);
and U13848 (N_13848,N_13011,N_13447);
nand U13849 (N_13849,N_13400,N_12917);
xor U13850 (N_13850,N_13050,N_12851);
and U13851 (N_13851,N_13063,N_12952);
nor U13852 (N_13852,N_12810,N_12891);
or U13853 (N_13853,N_13362,N_13466);
nor U13854 (N_13854,N_13135,N_12884);
xnor U13855 (N_13855,N_12986,N_13307);
or U13856 (N_13856,N_13231,N_13342);
xor U13857 (N_13857,N_13296,N_12969);
and U13858 (N_13858,N_12816,N_12856);
nor U13859 (N_13859,N_13390,N_13487);
or U13860 (N_13860,N_13043,N_12862);
nand U13861 (N_13861,N_13155,N_13080);
xnor U13862 (N_13862,N_13449,N_13497);
or U13863 (N_13863,N_13548,N_13054);
or U13864 (N_13864,N_13331,N_12999);
or U13865 (N_13865,N_13132,N_13260);
nor U13866 (N_13866,N_13524,N_13335);
and U13867 (N_13867,N_13310,N_13549);
nor U13868 (N_13868,N_13397,N_13102);
or U13869 (N_13869,N_13334,N_13522);
nand U13870 (N_13870,N_13490,N_13252);
or U13871 (N_13871,N_12954,N_13187);
or U13872 (N_13872,N_13027,N_12905);
or U13873 (N_13873,N_13536,N_13075);
nand U13874 (N_13874,N_13099,N_12837);
nor U13875 (N_13875,N_13205,N_13350);
or U13876 (N_13876,N_13190,N_13282);
and U13877 (N_13877,N_13045,N_13076);
and U13878 (N_13878,N_13258,N_13156);
or U13879 (N_13879,N_13148,N_13209);
and U13880 (N_13880,N_12958,N_13470);
or U13881 (N_13881,N_12990,N_13238);
or U13882 (N_13882,N_13516,N_12860);
xnor U13883 (N_13883,N_13090,N_12842);
nor U13884 (N_13884,N_13398,N_13157);
xor U13885 (N_13885,N_13424,N_13217);
nor U13886 (N_13886,N_13262,N_12825);
nand U13887 (N_13887,N_13418,N_12893);
xor U13888 (N_13888,N_13597,N_12807);
xor U13889 (N_13889,N_12881,N_13015);
xnor U13890 (N_13890,N_12823,N_13457);
or U13891 (N_13891,N_13304,N_12811);
and U13892 (N_13892,N_12974,N_13589);
nand U13893 (N_13893,N_13003,N_13113);
xor U13894 (N_13894,N_13289,N_13393);
nor U13895 (N_13895,N_13188,N_12924);
nand U13896 (N_13896,N_12970,N_13264);
nor U13897 (N_13897,N_13446,N_13104);
nand U13898 (N_13898,N_13373,N_13326);
and U13899 (N_13899,N_13092,N_13529);
or U13900 (N_13900,N_13117,N_13363);
nand U13901 (N_13901,N_12979,N_13030);
nand U13902 (N_13902,N_13066,N_13131);
xnor U13903 (N_13903,N_13300,N_13389);
nor U13904 (N_13904,N_13295,N_13530);
or U13905 (N_13905,N_13259,N_13077);
nand U13906 (N_13906,N_13189,N_12877);
xnor U13907 (N_13907,N_12867,N_13301);
or U13908 (N_13908,N_12927,N_13395);
xor U13909 (N_13909,N_13534,N_13215);
or U13910 (N_13910,N_13394,N_13435);
nor U13911 (N_13911,N_13172,N_13484);
xnor U13912 (N_13912,N_13024,N_13019);
xnor U13913 (N_13913,N_12921,N_13438);
or U13914 (N_13914,N_13445,N_12942);
xor U13915 (N_13915,N_12888,N_12890);
nor U13916 (N_13916,N_12804,N_13403);
nor U13917 (N_13917,N_13224,N_13442);
nand U13918 (N_13918,N_13051,N_12915);
nand U13919 (N_13919,N_13510,N_13288);
nor U13920 (N_13920,N_13354,N_13432);
and U13921 (N_13921,N_13496,N_12901);
or U13922 (N_13922,N_13218,N_13504);
and U13923 (N_13923,N_12937,N_13166);
nor U13924 (N_13924,N_12971,N_13227);
nor U13925 (N_13925,N_12895,N_13221);
nor U13926 (N_13926,N_13358,N_13391);
nor U13927 (N_13927,N_13551,N_13323);
nand U13928 (N_13928,N_13461,N_13337);
or U13929 (N_13929,N_13456,N_13339);
or U13930 (N_13930,N_12920,N_12911);
nand U13931 (N_13931,N_13056,N_13180);
and U13932 (N_13932,N_13291,N_13007);
xnor U13933 (N_13933,N_12843,N_13486);
and U13934 (N_13934,N_13083,N_13153);
or U13935 (N_13935,N_13142,N_13026);
nor U13936 (N_13936,N_13450,N_13266);
or U13937 (N_13937,N_13210,N_13590);
or U13938 (N_13938,N_13322,N_13444);
xnor U13939 (N_13939,N_13097,N_13114);
xnor U13940 (N_13940,N_12909,N_13060);
nor U13941 (N_13941,N_13399,N_12857);
and U13942 (N_13942,N_12955,N_12848);
xor U13943 (N_13943,N_13420,N_12866);
nand U13944 (N_13944,N_13223,N_12879);
and U13945 (N_13945,N_12896,N_12883);
or U13946 (N_13946,N_12949,N_12922);
and U13947 (N_13947,N_13459,N_13523);
or U13948 (N_13948,N_12992,N_13220);
or U13949 (N_13949,N_13071,N_13511);
xnor U13950 (N_13950,N_13257,N_12828);
or U13951 (N_13951,N_13278,N_13170);
xor U13952 (N_13952,N_12919,N_13411);
and U13953 (N_13953,N_13441,N_13255);
or U13954 (N_13954,N_12836,N_12926);
nand U13955 (N_13955,N_13107,N_13110);
nand U13956 (N_13956,N_13239,N_13366);
nand U13957 (N_13957,N_13226,N_13367);
nand U13958 (N_13958,N_13309,N_12845);
xnor U13959 (N_13959,N_13521,N_12944);
nor U13960 (N_13960,N_13319,N_12824);
or U13961 (N_13961,N_13021,N_12973);
and U13962 (N_13962,N_13292,N_13173);
nand U13963 (N_13963,N_13396,N_13029);
and U13964 (N_13964,N_13317,N_13191);
nor U13965 (N_13965,N_13573,N_12989);
xnor U13966 (N_13966,N_12957,N_12996);
nand U13967 (N_13967,N_13581,N_13001);
nand U13968 (N_13968,N_13381,N_13163);
and U13969 (N_13969,N_13149,N_12943);
xnor U13970 (N_13970,N_13475,N_12951);
xor U13971 (N_13971,N_13203,N_13320);
or U13972 (N_13972,N_13433,N_12932);
and U13973 (N_13973,N_12835,N_13127);
xnor U13974 (N_13974,N_12849,N_13287);
and U13975 (N_13975,N_13137,N_13101);
nand U13976 (N_13976,N_13387,N_13500);
nor U13977 (N_13977,N_13423,N_12980);
nor U13978 (N_13978,N_13469,N_13006);
or U13979 (N_13979,N_12813,N_13146);
or U13980 (N_13980,N_13360,N_13174);
or U13981 (N_13981,N_13035,N_13017);
or U13982 (N_13982,N_13448,N_13436);
or U13983 (N_13983,N_13293,N_13379);
and U13984 (N_13984,N_12833,N_12935);
nand U13985 (N_13985,N_13439,N_13208);
nand U13986 (N_13986,N_12966,N_13407);
nand U13987 (N_13987,N_13474,N_13095);
xnor U13988 (N_13988,N_13495,N_12930);
nand U13989 (N_13989,N_13184,N_13513);
xor U13990 (N_13990,N_13065,N_12886);
nor U13991 (N_13991,N_13041,N_13129);
nor U13992 (N_13992,N_13406,N_13416);
nand U13993 (N_13993,N_13134,N_13145);
nor U13994 (N_13994,N_13279,N_13422);
xnor U13995 (N_13995,N_13421,N_13431);
or U13996 (N_13996,N_13364,N_12912);
nor U13997 (N_13997,N_13488,N_12847);
xor U13998 (N_13998,N_13103,N_13138);
nor U13999 (N_13999,N_13481,N_13150);
xnor U14000 (N_14000,N_13370,N_13422);
nand U14001 (N_14001,N_13489,N_13058);
nand U14002 (N_14002,N_13250,N_13376);
nor U14003 (N_14003,N_13327,N_13295);
nor U14004 (N_14004,N_13069,N_13368);
nor U14005 (N_14005,N_13070,N_13375);
and U14006 (N_14006,N_13553,N_12845);
nor U14007 (N_14007,N_13156,N_13377);
xor U14008 (N_14008,N_13581,N_13593);
nor U14009 (N_14009,N_12879,N_12884);
or U14010 (N_14010,N_12832,N_13506);
nand U14011 (N_14011,N_13578,N_12841);
nand U14012 (N_14012,N_13111,N_12909);
and U14013 (N_14013,N_13430,N_13435);
nor U14014 (N_14014,N_13286,N_13019);
or U14015 (N_14015,N_13343,N_13407);
or U14016 (N_14016,N_13264,N_13093);
xnor U14017 (N_14017,N_12814,N_13585);
or U14018 (N_14018,N_13507,N_13020);
xor U14019 (N_14019,N_13546,N_13520);
xnor U14020 (N_14020,N_13300,N_13519);
xnor U14021 (N_14021,N_13348,N_13011);
or U14022 (N_14022,N_13314,N_12915);
nor U14023 (N_14023,N_13230,N_13077);
or U14024 (N_14024,N_13226,N_13010);
and U14025 (N_14025,N_13177,N_13450);
xor U14026 (N_14026,N_13225,N_13223);
nand U14027 (N_14027,N_12885,N_12951);
and U14028 (N_14028,N_13248,N_12907);
or U14029 (N_14029,N_13079,N_13333);
or U14030 (N_14030,N_12959,N_13454);
and U14031 (N_14031,N_13570,N_12970);
nand U14032 (N_14032,N_12833,N_13547);
or U14033 (N_14033,N_13073,N_13227);
xor U14034 (N_14034,N_13117,N_13224);
nand U14035 (N_14035,N_12916,N_12965);
or U14036 (N_14036,N_13471,N_13100);
nand U14037 (N_14037,N_12851,N_12855);
and U14038 (N_14038,N_13091,N_12953);
nor U14039 (N_14039,N_13559,N_13261);
and U14040 (N_14040,N_13567,N_13469);
xnor U14041 (N_14041,N_12857,N_13336);
nand U14042 (N_14042,N_13104,N_13507);
and U14043 (N_14043,N_13394,N_13376);
xnor U14044 (N_14044,N_13226,N_13127);
and U14045 (N_14045,N_13098,N_13415);
xor U14046 (N_14046,N_13338,N_13296);
xnor U14047 (N_14047,N_12844,N_13390);
xor U14048 (N_14048,N_13492,N_13050);
nand U14049 (N_14049,N_13030,N_13008);
or U14050 (N_14050,N_13530,N_13388);
nand U14051 (N_14051,N_12961,N_12914);
nand U14052 (N_14052,N_13508,N_13145);
nand U14053 (N_14053,N_12843,N_13267);
xor U14054 (N_14054,N_13312,N_12944);
and U14055 (N_14055,N_13373,N_13485);
nand U14056 (N_14056,N_13368,N_13135);
and U14057 (N_14057,N_12867,N_13597);
nand U14058 (N_14058,N_13060,N_12842);
xor U14059 (N_14059,N_12934,N_12911);
nor U14060 (N_14060,N_13115,N_13353);
and U14061 (N_14061,N_13585,N_13556);
or U14062 (N_14062,N_13558,N_13181);
nor U14063 (N_14063,N_13270,N_12948);
and U14064 (N_14064,N_13442,N_13360);
nand U14065 (N_14065,N_13204,N_13263);
nor U14066 (N_14066,N_13461,N_13557);
nor U14067 (N_14067,N_13506,N_13193);
and U14068 (N_14068,N_13035,N_13337);
xor U14069 (N_14069,N_13056,N_13005);
nor U14070 (N_14070,N_13113,N_12821);
and U14071 (N_14071,N_13308,N_13342);
and U14072 (N_14072,N_12860,N_13046);
nand U14073 (N_14073,N_13078,N_12941);
and U14074 (N_14074,N_13503,N_13301);
or U14075 (N_14075,N_13063,N_12837);
and U14076 (N_14076,N_13126,N_13456);
and U14077 (N_14077,N_13330,N_13285);
nor U14078 (N_14078,N_13471,N_13537);
xnor U14079 (N_14079,N_13293,N_13213);
nand U14080 (N_14080,N_13227,N_13391);
xnor U14081 (N_14081,N_12856,N_13391);
and U14082 (N_14082,N_13352,N_13555);
and U14083 (N_14083,N_12960,N_13489);
xnor U14084 (N_14084,N_13512,N_13224);
or U14085 (N_14085,N_13167,N_13065);
xnor U14086 (N_14086,N_13278,N_13577);
nand U14087 (N_14087,N_13291,N_13506);
or U14088 (N_14088,N_13075,N_13547);
nor U14089 (N_14089,N_12918,N_13041);
nor U14090 (N_14090,N_13140,N_12928);
nor U14091 (N_14091,N_13446,N_13449);
or U14092 (N_14092,N_13189,N_13100);
xor U14093 (N_14093,N_13122,N_12829);
nor U14094 (N_14094,N_13560,N_13569);
xor U14095 (N_14095,N_13525,N_13263);
and U14096 (N_14096,N_13563,N_13254);
or U14097 (N_14097,N_13071,N_13255);
nor U14098 (N_14098,N_13420,N_13296);
and U14099 (N_14099,N_12997,N_13327);
nor U14100 (N_14100,N_13339,N_13420);
or U14101 (N_14101,N_12813,N_13247);
xor U14102 (N_14102,N_13226,N_13437);
nor U14103 (N_14103,N_13234,N_13443);
nand U14104 (N_14104,N_13398,N_12978);
nor U14105 (N_14105,N_12847,N_12932);
and U14106 (N_14106,N_12951,N_13252);
nand U14107 (N_14107,N_13518,N_13589);
nor U14108 (N_14108,N_13366,N_12890);
or U14109 (N_14109,N_13347,N_12856);
nand U14110 (N_14110,N_13446,N_13198);
or U14111 (N_14111,N_13092,N_13224);
or U14112 (N_14112,N_12910,N_13250);
and U14113 (N_14113,N_13426,N_13226);
nand U14114 (N_14114,N_13283,N_13274);
or U14115 (N_14115,N_13119,N_12932);
nand U14116 (N_14116,N_13580,N_13379);
and U14117 (N_14117,N_13043,N_13253);
or U14118 (N_14118,N_13163,N_12840);
or U14119 (N_14119,N_12940,N_13040);
and U14120 (N_14120,N_13418,N_13296);
or U14121 (N_14121,N_13548,N_13152);
and U14122 (N_14122,N_13318,N_13441);
or U14123 (N_14123,N_13102,N_13130);
and U14124 (N_14124,N_12812,N_13448);
nor U14125 (N_14125,N_13083,N_13159);
xnor U14126 (N_14126,N_12945,N_13375);
or U14127 (N_14127,N_13583,N_13537);
xor U14128 (N_14128,N_13315,N_13252);
and U14129 (N_14129,N_13332,N_13206);
nand U14130 (N_14130,N_13146,N_13078);
or U14131 (N_14131,N_12984,N_13599);
nor U14132 (N_14132,N_13389,N_13347);
or U14133 (N_14133,N_12890,N_13489);
nand U14134 (N_14134,N_12881,N_13269);
nor U14135 (N_14135,N_13382,N_13598);
and U14136 (N_14136,N_13525,N_12912);
and U14137 (N_14137,N_13533,N_13220);
nor U14138 (N_14138,N_13353,N_13255);
xnor U14139 (N_14139,N_13353,N_13372);
nor U14140 (N_14140,N_13187,N_12948);
or U14141 (N_14141,N_12986,N_12850);
nand U14142 (N_14142,N_12800,N_12929);
and U14143 (N_14143,N_13086,N_13008);
and U14144 (N_14144,N_13070,N_13404);
and U14145 (N_14145,N_13418,N_13183);
or U14146 (N_14146,N_13297,N_13009);
nor U14147 (N_14147,N_13051,N_13472);
nor U14148 (N_14148,N_13145,N_13399);
nor U14149 (N_14149,N_13056,N_13150);
nor U14150 (N_14150,N_13137,N_13504);
xnor U14151 (N_14151,N_13398,N_13288);
nand U14152 (N_14152,N_13155,N_12992);
xnor U14153 (N_14153,N_13505,N_13178);
and U14154 (N_14154,N_13475,N_13321);
nand U14155 (N_14155,N_13277,N_12992);
nor U14156 (N_14156,N_13065,N_12817);
nor U14157 (N_14157,N_13034,N_12984);
xnor U14158 (N_14158,N_13558,N_13199);
nand U14159 (N_14159,N_13428,N_12808);
or U14160 (N_14160,N_13134,N_12937);
nor U14161 (N_14161,N_13125,N_12846);
nor U14162 (N_14162,N_13013,N_13043);
nor U14163 (N_14163,N_13508,N_13140);
and U14164 (N_14164,N_13108,N_13558);
nor U14165 (N_14165,N_13419,N_13557);
and U14166 (N_14166,N_13169,N_12996);
xnor U14167 (N_14167,N_13035,N_13003);
nand U14168 (N_14168,N_13153,N_13508);
nor U14169 (N_14169,N_12878,N_13327);
nor U14170 (N_14170,N_13173,N_13076);
nor U14171 (N_14171,N_13547,N_13291);
nor U14172 (N_14172,N_13388,N_12910);
nor U14173 (N_14173,N_13568,N_13254);
nand U14174 (N_14174,N_13336,N_13217);
xor U14175 (N_14175,N_13290,N_13266);
xor U14176 (N_14176,N_12944,N_13530);
and U14177 (N_14177,N_13537,N_13499);
nor U14178 (N_14178,N_12931,N_13132);
or U14179 (N_14179,N_13556,N_13180);
and U14180 (N_14180,N_13596,N_12910);
or U14181 (N_14181,N_13552,N_12993);
nand U14182 (N_14182,N_12964,N_13319);
and U14183 (N_14183,N_12987,N_13264);
xnor U14184 (N_14184,N_13498,N_13576);
and U14185 (N_14185,N_13220,N_13429);
xnor U14186 (N_14186,N_13021,N_13237);
nor U14187 (N_14187,N_13067,N_12982);
and U14188 (N_14188,N_13411,N_13499);
and U14189 (N_14189,N_13335,N_13004);
and U14190 (N_14190,N_13330,N_12844);
nand U14191 (N_14191,N_13563,N_13520);
or U14192 (N_14192,N_13044,N_13148);
or U14193 (N_14193,N_13352,N_13222);
nor U14194 (N_14194,N_13381,N_13317);
xnor U14195 (N_14195,N_13014,N_13302);
nand U14196 (N_14196,N_13093,N_12810);
and U14197 (N_14197,N_13465,N_12849);
nor U14198 (N_14198,N_12876,N_13571);
nand U14199 (N_14199,N_12824,N_12869);
nand U14200 (N_14200,N_13233,N_13466);
and U14201 (N_14201,N_13379,N_13052);
nand U14202 (N_14202,N_13313,N_13044);
and U14203 (N_14203,N_13021,N_13418);
or U14204 (N_14204,N_13347,N_13219);
or U14205 (N_14205,N_12815,N_12840);
nand U14206 (N_14206,N_13069,N_13162);
and U14207 (N_14207,N_13498,N_12880);
and U14208 (N_14208,N_12815,N_13291);
or U14209 (N_14209,N_12982,N_13502);
xnor U14210 (N_14210,N_13071,N_13265);
nor U14211 (N_14211,N_13471,N_12900);
and U14212 (N_14212,N_13341,N_13397);
nand U14213 (N_14213,N_13081,N_13485);
xor U14214 (N_14214,N_13231,N_13026);
nor U14215 (N_14215,N_12977,N_13127);
xor U14216 (N_14216,N_12836,N_13341);
xnor U14217 (N_14217,N_13065,N_13231);
and U14218 (N_14218,N_13538,N_13519);
nand U14219 (N_14219,N_13037,N_13154);
nand U14220 (N_14220,N_13121,N_13481);
nand U14221 (N_14221,N_13223,N_12851);
xor U14222 (N_14222,N_13284,N_13348);
nand U14223 (N_14223,N_13599,N_12874);
xor U14224 (N_14224,N_13335,N_13112);
and U14225 (N_14225,N_12942,N_13213);
nand U14226 (N_14226,N_13297,N_13243);
xnor U14227 (N_14227,N_13452,N_13177);
and U14228 (N_14228,N_13472,N_13287);
xor U14229 (N_14229,N_13056,N_13168);
xnor U14230 (N_14230,N_13162,N_13501);
nor U14231 (N_14231,N_13391,N_12825);
nand U14232 (N_14232,N_13307,N_13166);
or U14233 (N_14233,N_12931,N_13182);
nand U14234 (N_14234,N_13036,N_13172);
nor U14235 (N_14235,N_12810,N_13413);
xor U14236 (N_14236,N_13547,N_12879);
and U14237 (N_14237,N_13200,N_13392);
and U14238 (N_14238,N_12960,N_13393);
nand U14239 (N_14239,N_13233,N_13027);
and U14240 (N_14240,N_13432,N_13584);
xnor U14241 (N_14241,N_12935,N_12897);
nand U14242 (N_14242,N_13349,N_12933);
nand U14243 (N_14243,N_13509,N_12821);
nand U14244 (N_14244,N_13557,N_13390);
nand U14245 (N_14245,N_13534,N_12919);
xnor U14246 (N_14246,N_12824,N_13457);
or U14247 (N_14247,N_12803,N_12989);
nand U14248 (N_14248,N_13542,N_13487);
or U14249 (N_14249,N_13314,N_13014);
nand U14250 (N_14250,N_13391,N_13434);
nor U14251 (N_14251,N_12879,N_13291);
xor U14252 (N_14252,N_13487,N_13106);
or U14253 (N_14253,N_13200,N_13105);
nor U14254 (N_14254,N_13117,N_13367);
nand U14255 (N_14255,N_13127,N_13166);
or U14256 (N_14256,N_13568,N_13574);
and U14257 (N_14257,N_13004,N_13182);
nand U14258 (N_14258,N_13488,N_13144);
nor U14259 (N_14259,N_12890,N_12934);
and U14260 (N_14260,N_13048,N_13125);
xor U14261 (N_14261,N_13596,N_13378);
xor U14262 (N_14262,N_13278,N_13349);
and U14263 (N_14263,N_13478,N_13420);
xnor U14264 (N_14264,N_13494,N_13340);
and U14265 (N_14265,N_13334,N_13393);
nand U14266 (N_14266,N_13325,N_13575);
nor U14267 (N_14267,N_13563,N_12938);
xor U14268 (N_14268,N_13010,N_13011);
nor U14269 (N_14269,N_13233,N_13069);
xnor U14270 (N_14270,N_12887,N_12909);
and U14271 (N_14271,N_13458,N_13472);
nand U14272 (N_14272,N_13259,N_13246);
nand U14273 (N_14273,N_13069,N_13147);
nor U14274 (N_14274,N_12827,N_13194);
xnor U14275 (N_14275,N_13056,N_13314);
nor U14276 (N_14276,N_12851,N_12844);
nor U14277 (N_14277,N_13504,N_12939);
and U14278 (N_14278,N_12996,N_13276);
or U14279 (N_14279,N_13460,N_13425);
xor U14280 (N_14280,N_13328,N_12895);
and U14281 (N_14281,N_13014,N_13537);
and U14282 (N_14282,N_13164,N_13373);
nor U14283 (N_14283,N_13437,N_13583);
and U14284 (N_14284,N_13044,N_12999);
xor U14285 (N_14285,N_13559,N_13138);
and U14286 (N_14286,N_13530,N_12908);
xnor U14287 (N_14287,N_13346,N_13464);
and U14288 (N_14288,N_13491,N_13399);
nor U14289 (N_14289,N_12883,N_13376);
nor U14290 (N_14290,N_13272,N_12968);
nand U14291 (N_14291,N_13096,N_13021);
nor U14292 (N_14292,N_13128,N_12881);
nor U14293 (N_14293,N_13263,N_13508);
nand U14294 (N_14294,N_13560,N_13067);
nor U14295 (N_14295,N_13019,N_12984);
and U14296 (N_14296,N_13454,N_13043);
nand U14297 (N_14297,N_13396,N_13254);
nor U14298 (N_14298,N_13338,N_13343);
nor U14299 (N_14299,N_13373,N_13253);
nand U14300 (N_14300,N_13237,N_13471);
or U14301 (N_14301,N_13453,N_13034);
nand U14302 (N_14302,N_13210,N_13401);
nand U14303 (N_14303,N_13254,N_12880);
nand U14304 (N_14304,N_12815,N_12923);
nor U14305 (N_14305,N_13111,N_13130);
xnor U14306 (N_14306,N_12934,N_13360);
and U14307 (N_14307,N_12823,N_13293);
nor U14308 (N_14308,N_12850,N_12943);
xnor U14309 (N_14309,N_13458,N_13002);
nand U14310 (N_14310,N_12811,N_13330);
or U14311 (N_14311,N_12996,N_13209);
nor U14312 (N_14312,N_13361,N_13183);
nand U14313 (N_14313,N_12892,N_13538);
xnor U14314 (N_14314,N_13250,N_13557);
xor U14315 (N_14315,N_12914,N_13552);
xor U14316 (N_14316,N_13362,N_13179);
xnor U14317 (N_14317,N_13133,N_13370);
nand U14318 (N_14318,N_12820,N_12878);
xor U14319 (N_14319,N_13249,N_12992);
and U14320 (N_14320,N_13180,N_13365);
xor U14321 (N_14321,N_13350,N_13073);
or U14322 (N_14322,N_13461,N_12808);
and U14323 (N_14323,N_13377,N_13070);
nor U14324 (N_14324,N_13216,N_13513);
and U14325 (N_14325,N_12978,N_13346);
and U14326 (N_14326,N_12918,N_13459);
and U14327 (N_14327,N_13212,N_13218);
and U14328 (N_14328,N_13484,N_13115);
xor U14329 (N_14329,N_13580,N_13221);
xnor U14330 (N_14330,N_13599,N_13475);
nor U14331 (N_14331,N_12815,N_12898);
nand U14332 (N_14332,N_13327,N_12853);
nor U14333 (N_14333,N_13278,N_13580);
and U14334 (N_14334,N_12881,N_13296);
xor U14335 (N_14335,N_12828,N_13211);
xor U14336 (N_14336,N_13002,N_13423);
and U14337 (N_14337,N_13510,N_12870);
and U14338 (N_14338,N_13125,N_13146);
nand U14339 (N_14339,N_12869,N_12819);
nand U14340 (N_14340,N_13481,N_12878);
and U14341 (N_14341,N_12995,N_13208);
nand U14342 (N_14342,N_13176,N_13436);
nor U14343 (N_14343,N_13023,N_13581);
xnor U14344 (N_14344,N_12959,N_12826);
nand U14345 (N_14345,N_13110,N_13288);
xor U14346 (N_14346,N_13576,N_13225);
nor U14347 (N_14347,N_13308,N_13497);
nand U14348 (N_14348,N_13157,N_13367);
or U14349 (N_14349,N_12927,N_13239);
nand U14350 (N_14350,N_13008,N_13323);
or U14351 (N_14351,N_13048,N_13092);
and U14352 (N_14352,N_13029,N_13551);
xnor U14353 (N_14353,N_13049,N_13472);
nor U14354 (N_14354,N_13431,N_13012);
nor U14355 (N_14355,N_13181,N_13285);
nand U14356 (N_14356,N_13573,N_13165);
nor U14357 (N_14357,N_12823,N_13102);
nor U14358 (N_14358,N_12994,N_13458);
and U14359 (N_14359,N_13043,N_13218);
xnor U14360 (N_14360,N_12866,N_13087);
xor U14361 (N_14361,N_13116,N_13114);
and U14362 (N_14362,N_13479,N_12870);
nand U14363 (N_14363,N_13066,N_13566);
xnor U14364 (N_14364,N_13118,N_13032);
xor U14365 (N_14365,N_13550,N_13099);
nand U14366 (N_14366,N_13417,N_13436);
or U14367 (N_14367,N_13133,N_13257);
nor U14368 (N_14368,N_13413,N_12887);
nor U14369 (N_14369,N_13069,N_12920);
and U14370 (N_14370,N_12997,N_12861);
xor U14371 (N_14371,N_13389,N_13176);
xnor U14372 (N_14372,N_13234,N_13487);
nor U14373 (N_14373,N_13507,N_12822);
and U14374 (N_14374,N_12888,N_12951);
or U14375 (N_14375,N_13429,N_12942);
nor U14376 (N_14376,N_13589,N_12991);
xnor U14377 (N_14377,N_13238,N_13422);
or U14378 (N_14378,N_13121,N_13398);
xnor U14379 (N_14379,N_13339,N_13279);
and U14380 (N_14380,N_13295,N_13591);
nor U14381 (N_14381,N_13396,N_12845);
or U14382 (N_14382,N_13095,N_12994);
nand U14383 (N_14383,N_12894,N_12960);
nor U14384 (N_14384,N_12818,N_13501);
and U14385 (N_14385,N_13574,N_12883);
or U14386 (N_14386,N_12875,N_12817);
nand U14387 (N_14387,N_13329,N_12989);
or U14388 (N_14388,N_13305,N_12853);
or U14389 (N_14389,N_13444,N_13381);
nand U14390 (N_14390,N_13210,N_13558);
xnor U14391 (N_14391,N_13357,N_13147);
or U14392 (N_14392,N_13517,N_13412);
nor U14393 (N_14393,N_13286,N_12999);
and U14394 (N_14394,N_12884,N_13598);
xnor U14395 (N_14395,N_13004,N_13414);
and U14396 (N_14396,N_13418,N_13540);
xnor U14397 (N_14397,N_13148,N_13482);
nand U14398 (N_14398,N_13188,N_12807);
xnor U14399 (N_14399,N_13305,N_13425);
or U14400 (N_14400,N_14017,N_14160);
and U14401 (N_14401,N_14230,N_14047);
and U14402 (N_14402,N_14080,N_13664);
xnor U14403 (N_14403,N_13946,N_14092);
or U14404 (N_14404,N_13990,N_13941);
nor U14405 (N_14405,N_14114,N_13957);
xnor U14406 (N_14406,N_13892,N_14390);
and U14407 (N_14407,N_13956,N_14016);
and U14408 (N_14408,N_13783,N_13913);
nor U14409 (N_14409,N_13944,N_13991);
nor U14410 (N_14410,N_13795,N_14136);
xor U14411 (N_14411,N_14144,N_14165);
xor U14412 (N_14412,N_13730,N_13888);
and U14413 (N_14413,N_14188,N_13665);
or U14414 (N_14414,N_14349,N_13942);
and U14415 (N_14415,N_14151,N_14350);
and U14416 (N_14416,N_14302,N_13756);
and U14417 (N_14417,N_14061,N_13692);
nand U14418 (N_14418,N_14204,N_13971);
nand U14419 (N_14419,N_14170,N_13858);
nand U14420 (N_14420,N_13828,N_14276);
nand U14421 (N_14421,N_14185,N_14056);
nand U14422 (N_14422,N_13840,N_13886);
xor U14423 (N_14423,N_13959,N_14281);
nor U14424 (N_14424,N_14389,N_13898);
xor U14425 (N_14425,N_13698,N_14308);
or U14426 (N_14426,N_14316,N_14266);
nor U14427 (N_14427,N_13667,N_13878);
nand U14428 (N_14428,N_13845,N_14196);
nand U14429 (N_14429,N_14096,N_14026);
and U14430 (N_14430,N_13853,N_14053);
nand U14431 (N_14431,N_14384,N_13741);
nand U14432 (N_14432,N_13856,N_13843);
and U14433 (N_14433,N_13643,N_13639);
or U14434 (N_14434,N_13661,N_13775);
and U14435 (N_14435,N_14296,N_13790);
and U14436 (N_14436,N_13953,N_13686);
xor U14437 (N_14437,N_13960,N_14381);
nor U14438 (N_14438,N_14356,N_14270);
or U14439 (N_14439,N_14152,N_13640);
nand U14440 (N_14440,N_14089,N_14127);
nand U14441 (N_14441,N_14087,N_14262);
nand U14442 (N_14442,N_14365,N_13810);
and U14443 (N_14443,N_14298,N_14139);
or U14444 (N_14444,N_13601,N_13937);
xnor U14445 (N_14445,N_13987,N_13777);
nor U14446 (N_14446,N_13964,N_13890);
nand U14447 (N_14447,N_13945,N_13762);
nand U14448 (N_14448,N_13879,N_13785);
xor U14449 (N_14449,N_13757,N_14081);
nand U14450 (N_14450,N_13802,N_14135);
nor U14451 (N_14451,N_13862,N_14202);
nand U14452 (N_14452,N_13723,N_14201);
nand U14453 (N_14453,N_13715,N_14077);
nand U14454 (N_14454,N_13935,N_14210);
nor U14455 (N_14455,N_14271,N_13712);
and U14456 (N_14456,N_13928,N_13763);
and U14457 (N_14457,N_13829,N_14035);
nand U14458 (N_14458,N_13706,N_13826);
nand U14459 (N_14459,N_13974,N_13770);
nand U14460 (N_14460,N_14231,N_14304);
nor U14461 (N_14461,N_13732,N_14293);
nand U14462 (N_14462,N_13659,N_13710);
and U14463 (N_14463,N_14004,N_13678);
or U14464 (N_14464,N_13847,N_14237);
nand U14465 (N_14465,N_13656,N_14387);
nor U14466 (N_14466,N_13815,N_14297);
xor U14467 (N_14467,N_14086,N_13984);
nor U14468 (N_14468,N_14166,N_14383);
and U14469 (N_14469,N_14221,N_14070);
or U14470 (N_14470,N_14343,N_14377);
and U14471 (N_14471,N_13700,N_13615);
xor U14472 (N_14472,N_14357,N_13871);
nor U14473 (N_14473,N_13827,N_14124);
and U14474 (N_14474,N_14208,N_13868);
or U14475 (N_14475,N_14300,N_13649);
xor U14476 (N_14476,N_14184,N_14279);
and U14477 (N_14477,N_13824,N_13830);
xor U14478 (N_14478,N_14075,N_14267);
and U14479 (N_14479,N_13943,N_13839);
xnor U14480 (N_14480,N_13663,N_13895);
and U14481 (N_14481,N_13658,N_13893);
or U14482 (N_14482,N_14321,N_14031);
or U14483 (N_14483,N_14030,N_14015);
or U14484 (N_14484,N_13743,N_13719);
and U14485 (N_14485,N_13911,N_13816);
nor U14486 (N_14486,N_13778,N_13642);
xor U14487 (N_14487,N_14288,N_13823);
or U14488 (N_14488,N_13767,N_13746);
nor U14489 (N_14489,N_13747,N_13889);
or U14490 (N_14490,N_13764,N_13855);
or U14491 (N_14491,N_13891,N_13672);
nor U14492 (N_14492,N_14173,N_13780);
or U14493 (N_14493,N_13836,N_13820);
nor U14494 (N_14494,N_14039,N_13948);
and U14495 (N_14495,N_14312,N_14146);
nor U14496 (N_14496,N_14244,N_13818);
nand U14497 (N_14497,N_13854,N_14046);
nand U14498 (N_14498,N_14223,N_13704);
nand U14499 (N_14499,N_13752,N_14337);
nor U14500 (N_14500,N_14339,N_13917);
or U14501 (N_14501,N_14088,N_13771);
and U14502 (N_14502,N_14023,N_14049);
or U14503 (N_14503,N_14100,N_13859);
nand U14504 (N_14504,N_13981,N_13821);
and U14505 (N_14505,N_14175,N_13793);
xor U14506 (N_14506,N_13671,N_14380);
or U14507 (N_14507,N_13654,N_14189);
nand U14508 (N_14508,N_13896,N_14001);
nand U14509 (N_14509,N_13994,N_13628);
xor U14510 (N_14510,N_13835,N_14118);
nand U14511 (N_14511,N_13860,N_14005);
nor U14512 (N_14512,N_13701,N_13967);
xnor U14513 (N_14513,N_13600,N_14248);
and U14514 (N_14514,N_13992,N_14050);
nand U14515 (N_14515,N_14022,N_14029);
nor U14516 (N_14516,N_14059,N_13753);
or U14517 (N_14517,N_14191,N_13958);
or U14518 (N_14518,N_14102,N_13884);
and U14519 (N_14519,N_14199,N_13765);
nor U14520 (N_14520,N_14363,N_13651);
and U14521 (N_14521,N_14299,N_13633);
and U14522 (N_14522,N_13936,N_14283);
and U14523 (N_14523,N_14095,N_13660);
and U14524 (N_14524,N_13690,N_13782);
nand U14525 (N_14525,N_13726,N_13852);
nand U14526 (N_14526,N_13922,N_13813);
or U14527 (N_14527,N_13982,N_14240);
or U14528 (N_14528,N_14093,N_14067);
and U14529 (N_14529,N_14251,N_13973);
and U14530 (N_14530,N_13697,N_14216);
or U14531 (N_14531,N_13625,N_14317);
or U14532 (N_14532,N_14280,N_14256);
xor U14533 (N_14533,N_13784,N_14111);
or U14534 (N_14534,N_13648,N_14252);
xnor U14535 (N_14535,N_14180,N_14024);
nor U14536 (N_14536,N_14368,N_14195);
nand U14537 (N_14537,N_14013,N_14370);
nand U14538 (N_14538,N_14048,N_13629);
xor U14539 (N_14539,N_13803,N_14028);
nand U14540 (N_14540,N_14141,N_13989);
nand U14541 (N_14541,N_14131,N_13833);
and U14542 (N_14542,N_14161,N_14206);
nand U14543 (N_14543,N_14328,N_13965);
nand U14544 (N_14544,N_14187,N_13761);
nor U14545 (N_14545,N_13605,N_14083);
or U14546 (N_14546,N_14305,N_14287);
nor U14547 (N_14547,N_13617,N_13621);
xor U14548 (N_14548,N_14174,N_13977);
xor U14549 (N_14549,N_14386,N_14018);
or U14550 (N_14550,N_13720,N_13685);
and U14551 (N_14551,N_13800,N_14218);
nor U14552 (N_14552,N_14063,N_13614);
and U14553 (N_14553,N_13910,N_13609);
or U14554 (N_14554,N_13923,N_13857);
nand U14555 (N_14555,N_14239,N_13787);
nand U14556 (N_14556,N_13729,N_13657);
nor U14557 (N_14557,N_14132,N_14398);
nor U14558 (N_14558,N_13819,N_14133);
or U14559 (N_14559,N_14392,N_14097);
and U14560 (N_14560,N_13993,N_14183);
xor U14561 (N_14561,N_13736,N_13679);
xnor U14562 (N_14562,N_14181,N_13724);
nand U14563 (N_14563,N_13972,N_13834);
nor U14564 (N_14564,N_14197,N_14130);
xnor U14565 (N_14565,N_14309,N_13655);
nand U14566 (N_14566,N_13718,N_14369);
xnor U14567 (N_14567,N_14007,N_13644);
nor U14568 (N_14568,N_14071,N_13637);
xor U14569 (N_14569,N_14045,N_13817);
or U14570 (N_14570,N_13635,N_14106);
and U14571 (N_14571,N_14385,N_13603);
nand U14572 (N_14572,N_13769,N_14113);
or U14573 (N_14573,N_13755,N_13900);
xnor U14574 (N_14574,N_14198,N_13880);
and U14575 (N_14575,N_14396,N_14027);
and U14576 (N_14576,N_13630,N_13636);
and U14577 (N_14577,N_14143,N_14224);
nand U14578 (N_14578,N_13662,N_13955);
nor U14579 (N_14579,N_14044,N_14294);
nor U14580 (N_14580,N_13885,N_13652);
or U14581 (N_14581,N_13675,N_14153);
nand U14582 (N_14582,N_14065,N_14324);
nand U14583 (N_14583,N_14145,N_14333);
or U14584 (N_14584,N_14043,N_13722);
xor U14585 (N_14585,N_13695,N_13882);
nand U14586 (N_14586,N_14213,N_13924);
or U14587 (N_14587,N_14278,N_14074);
and U14588 (N_14588,N_14104,N_13645);
nand U14589 (N_14589,N_14099,N_14229);
and U14590 (N_14590,N_14238,N_14259);
and U14591 (N_14591,N_13745,N_14137);
nand U14592 (N_14592,N_13939,N_14091);
nor U14593 (N_14593,N_13702,N_14362);
or U14594 (N_14594,N_13985,N_13738);
or U14595 (N_14595,N_13731,N_13687);
xor U14596 (N_14596,N_13613,N_14162);
xnor U14597 (N_14597,N_13750,N_14110);
nor U14598 (N_14598,N_13807,N_13804);
xnor U14599 (N_14599,N_14397,N_13930);
or U14600 (N_14600,N_14225,N_13708);
nand U14601 (N_14601,N_13799,N_14227);
and U14602 (N_14602,N_13934,N_14084);
nor U14603 (N_14603,N_14108,N_14042);
nand U14604 (N_14604,N_14179,N_14203);
nand U14605 (N_14605,N_13949,N_14395);
nand U14606 (N_14606,N_13768,N_14212);
and U14607 (N_14607,N_14347,N_14361);
and U14608 (N_14608,N_14066,N_14319);
nor U14609 (N_14609,N_14177,N_13773);
nand U14610 (N_14610,N_13986,N_13717);
nor U14611 (N_14611,N_13809,N_14032);
or U14612 (N_14612,N_14076,N_14372);
or U14613 (N_14613,N_14058,N_13881);
xor U14614 (N_14614,N_13808,N_13842);
nor U14615 (N_14615,N_14282,N_13838);
nand U14616 (N_14616,N_14090,N_13919);
nor U14617 (N_14617,N_14103,N_13801);
nor U14618 (N_14618,N_14354,N_13906);
nand U14619 (N_14619,N_14115,N_14375);
xnor U14620 (N_14620,N_13861,N_13734);
nand U14621 (N_14621,N_13754,N_14382);
xor U14622 (N_14622,N_14338,N_13618);
nand U14623 (N_14623,N_13760,N_14344);
nand U14624 (N_14624,N_13901,N_13647);
or U14625 (N_14625,N_13641,N_13844);
nand U14626 (N_14626,N_14054,N_14254);
nand U14627 (N_14627,N_13849,N_13608);
xnor U14628 (N_14628,N_13791,N_14192);
nor U14629 (N_14629,N_13980,N_14364);
or U14630 (N_14630,N_14117,N_14009);
nor U14631 (N_14631,N_13611,N_14399);
xor U14632 (N_14632,N_14352,N_14220);
nor U14633 (N_14633,N_13950,N_14391);
or U14634 (N_14634,N_14351,N_13966);
or U14635 (N_14635,N_14068,N_13962);
and U14636 (N_14636,N_13759,N_14367);
or U14637 (N_14637,N_14359,N_13669);
and U14638 (N_14638,N_14311,N_14335);
or U14639 (N_14639,N_13707,N_13694);
nand U14640 (N_14640,N_13899,N_14277);
nand U14641 (N_14641,N_13999,N_13825);
nand U14642 (N_14642,N_13794,N_13997);
nor U14643 (N_14643,N_14138,N_14329);
nand U14644 (N_14644,N_14261,N_14057);
nand U14645 (N_14645,N_13869,N_14129);
and U14646 (N_14646,N_14034,N_13622);
xnor U14647 (N_14647,N_14194,N_14322);
xor U14648 (N_14648,N_14010,N_13742);
xnor U14649 (N_14649,N_13875,N_14393);
or U14650 (N_14650,N_14025,N_13766);
nor U14651 (N_14651,N_13797,N_14082);
nor U14652 (N_14652,N_14353,N_14275);
xor U14653 (N_14653,N_14012,N_13902);
and U14654 (N_14654,N_14250,N_13607);
and U14655 (N_14655,N_13739,N_13716);
and U14656 (N_14656,N_13908,N_14167);
xnor U14657 (N_14657,N_13634,N_13968);
or U14658 (N_14658,N_13713,N_14006);
nand U14659 (N_14659,N_13865,N_13925);
nor U14660 (N_14660,N_14258,N_14011);
and U14661 (N_14661,N_14169,N_13872);
nor U14662 (N_14662,N_14209,N_14008);
xor U14663 (N_14663,N_14072,N_14182);
or U14664 (N_14664,N_14242,N_14348);
and U14665 (N_14665,N_14318,N_14320);
nand U14666 (N_14666,N_13931,N_13979);
xnor U14667 (N_14667,N_14323,N_13748);
or U14668 (N_14668,N_14085,N_14014);
or U14669 (N_14669,N_13866,N_13749);
and U14670 (N_14670,N_14388,N_13638);
xnor U14671 (N_14671,N_13699,N_14303);
or U14672 (N_14672,N_13626,N_14255);
nor U14673 (N_14673,N_13711,N_13619);
xnor U14674 (N_14674,N_14345,N_13867);
xor U14675 (N_14675,N_13788,N_14150);
or U14676 (N_14676,N_14268,N_14286);
xor U14677 (N_14677,N_14163,N_14306);
nand U14678 (N_14678,N_14079,N_14157);
xor U14679 (N_14679,N_14101,N_13848);
nor U14680 (N_14680,N_14078,N_14332);
xor U14681 (N_14681,N_13650,N_13926);
nand U14682 (N_14682,N_13932,N_13933);
xor U14683 (N_14683,N_14264,N_14128);
nand U14684 (N_14684,N_13796,N_14330);
nand U14685 (N_14685,N_13627,N_14284);
nor U14686 (N_14686,N_14155,N_14265);
or U14687 (N_14687,N_13689,N_14245);
or U14688 (N_14688,N_14219,N_13873);
or U14689 (N_14689,N_13954,N_14291);
or U14690 (N_14690,N_13863,N_14178);
or U14691 (N_14691,N_14314,N_13680);
or U14692 (N_14692,N_14358,N_13673);
nor U14693 (N_14693,N_14374,N_13894);
or U14694 (N_14694,N_13915,N_13846);
or U14695 (N_14695,N_13947,N_14315);
xnor U14696 (N_14696,N_14186,N_14215);
and U14697 (N_14697,N_13681,N_14217);
or U14698 (N_14698,N_13904,N_14378);
nor U14699 (N_14699,N_14147,N_13806);
xnor U14700 (N_14700,N_13912,N_13996);
xor U14701 (N_14701,N_14341,N_13975);
nand U14702 (N_14702,N_14064,N_13610);
and U14703 (N_14703,N_14257,N_14109);
xor U14704 (N_14704,N_13805,N_14292);
or U14705 (N_14705,N_13721,N_13666);
nand U14706 (N_14706,N_14360,N_14123);
and U14707 (N_14707,N_13837,N_13668);
nand U14708 (N_14708,N_14234,N_13612);
xor U14709 (N_14709,N_14289,N_13693);
xor U14710 (N_14710,N_13674,N_14355);
or U14711 (N_14711,N_13909,N_14326);
nor U14712 (N_14712,N_14062,N_14313);
nor U14713 (N_14713,N_13653,N_14346);
and U14714 (N_14714,N_13705,N_13887);
or U14715 (N_14715,N_14290,N_13940);
nand U14716 (N_14716,N_13918,N_13604);
xnor U14717 (N_14717,N_13876,N_13631);
xor U14718 (N_14718,N_13798,N_13779);
nor U14719 (N_14719,N_14060,N_13677);
nand U14720 (N_14720,N_14373,N_13851);
and U14721 (N_14721,N_13983,N_14200);
xnor U14722 (N_14722,N_13792,N_14207);
xor U14723 (N_14723,N_13850,N_13624);
xor U14724 (N_14724,N_14134,N_13976);
nand U14725 (N_14725,N_14325,N_14094);
xnor U14726 (N_14726,N_13623,N_13751);
nand U14727 (N_14727,N_13870,N_13874);
and U14728 (N_14728,N_14069,N_13728);
nor U14729 (N_14729,N_14263,N_14211);
nor U14730 (N_14730,N_14122,N_14222);
nor U14731 (N_14731,N_14020,N_14260);
and U14732 (N_14732,N_14371,N_13927);
and U14733 (N_14733,N_14107,N_13744);
xnor U14734 (N_14734,N_14190,N_14285);
xnor U14735 (N_14735,N_14176,N_13914);
and U14736 (N_14736,N_13877,N_13988);
and U14737 (N_14737,N_13737,N_13602);
xnor U14738 (N_14738,N_14140,N_14214);
or U14739 (N_14739,N_14394,N_13952);
nand U14740 (N_14740,N_14243,N_14051);
or U14741 (N_14741,N_13725,N_14098);
nand U14742 (N_14742,N_14233,N_14021);
or U14743 (N_14743,N_13995,N_14164);
xor U14744 (N_14744,N_14159,N_13907);
nand U14745 (N_14745,N_14126,N_13632);
nand U14746 (N_14746,N_14274,N_13814);
nor U14747 (N_14747,N_14002,N_13864);
and U14748 (N_14748,N_14331,N_14295);
or U14749 (N_14749,N_13606,N_14000);
and U14750 (N_14750,N_14158,N_14336);
nor U14751 (N_14751,N_13616,N_14040);
nand U14752 (N_14752,N_13897,N_13812);
xnor U14753 (N_14753,N_14205,N_14105);
xnor U14754 (N_14754,N_13714,N_14241);
xor U14755 (N_14755,N_14376,N_13691);
nand U14756 (N_14756,N_13929,N_14003);
or U14757 (N_14757,N_13916,N_14142);
or U14758 (N_14758,N_14366,N_13789);
or U14759 (N_14759,N_13772,N_14269);
and U14760 (N_14760,N_13920,N_14172);
nor U14761 (N_14761,N_14379,N_13905);
nor U14762 (N_14762,N_14340,N_14154);
nand U14763 (N_14763,N_14037,N_13727);
nor U14764 (N_14764,N_13688,N_14148);
xor U14765 (N_14765,N_14116,N_13670);
xor U14766 (N_14766,N_13703,N_13841);
or U14767 (N_14767,N_13963,N_14273);
nand U14768 (N_14768,N_13938,N_14156);
nor U14769 (N_14769,N_14228,N_14121);
xnor U14770 (N_14770,N_14168,N_13646);
nor U14771 (N_14771,N_13620,N_14236);
and U14772 (N_14772,N_14272,N_14149);
or U14773 (N_14773,N_14249,N_14307);
or U14774 (N_14774,N_13883,N_14310);
or U14775 (N_14775,N_14342,N_14327);
or U14776 (N_14776,N_14247,N_13733);
nand U14777 (N_14777,N_13822,N_13781);
nor U14778 (N_14778,N_13998,N_14119);
nand U14779 (N_14779,N_14235,N_13776);
nor U14780 (N_14780,N_14125,N_14055);
nor U14781 (N_14781,N_14193,N_13978);
or U14782 (N_14782,N_13696,N_13774);
or U14783 (N_14783,N_13951,N_13831);
or U14784 (N_14784,N_14041,N_14334);
nand U14785 (N_14785,N_13709,N_13903);
or U14786 (N_14786,N_14246,N_14301);
xor U14787 (N_14787,N_14052,N_13811);
nor U14788 (N_14788,N_14019,N_13682);
and U14789 (N_14789,N_14112,N_14073);
nor U14790 (N_14790,N_14171,N_14232);
nand U14791 (N_14791,N_13970,N_13683);
nor U14792 (N_14792,N_14226,N_13735);
or U14793 (N_14793,N_13786,N_13676);
nor U14794 (N_14794,N_13969,N_14038);
or U14795 (N_14795,N_13921,N_13832);
nor U14796 (N_14796,N_13740,N_13684);
or U14797 (N_14797,N_14036,N_14033);
and U14798 (N_14798,N_13758,N_14120);
nor U14799 (N_14799,N_13961,N_14253);
nor U14800 (N_14800,N_14226,N_14229);
or U14801 (N_14801,N_13873,N_13744);
or U14802 (N_14802,N_13840,N_14069);
and U14803 (N_14803,N_14318,N_13656);
and U14804 (N_14804,N_14095,N_13876);
nand U14805 (N_14805,N_14224,N_14239);
nor U14806 (N_14806,N_13796,N_14187);
xor U14807 (N_14807,N_14071,N_14026);
nor U14808 (N_14808,N_13690,N_14151);
nand U14809 (N_14809,N_14022,N_14105);
xnor U14810 (N_14810,N_14348,N_13701);
xnor U14811 (N_14811,N_13648,N_13821);
and U14812 (N_14812,N_14218,N_14078);
nor U14813 (N_14813,N_13774,N_13988);
nand U14814 (N_14814,N_13656,N_14088);
xnor U14815 (N_14815,N_14049,N_13695);
and U14816 (N_14816,N_14212,N_14399);
nand U14817 (N_14817,N_14178,N_14245);
xnor U14818 (N_14818,N_14014,N_14108);
or U14819 (N_14819,N_14357,N_13980);
or U14820 (N_14820,N_13679,N_14325);
xor U14821 (N_14821,N_14295,N_13841);
xor U14822 (N_14822,N_13973,N_14256);
xor U14823 (N_14823,N_13726,N_13739);
nor U14824 (N_14824,N_13798,N_13922);
and U14825 (N_14825,N_14066,N_13652);
nor U14826 (N_14826,N_13809,N_13647);
xor U14827 (N_14827,N_13887,N_13633);
nand U14828 (N_14828,N_14209,N_14360);
or U14829 (N_14829,N_14187,N_13924);
nor U14830 (N_14830,N_14047,N_14190);
and U14831 (N_14831,N_14308,N_13630);
and U14832 (N_14832,N_13720,N_13818);
and U14833 (N_14833,N_14334,N_13727);
or U14834 (N_14834,N_13870,N_13883);
xnor U14835 (N_14835,N_14148,N_14333);
xnor U14836 (N_14836,N_14024,N_14032);
xor U14837 (N_14837,N_14374,N_13958);
nand U14838 (N_14838,N_13895,N_14026);
nand U14839 (N_14839,N_14229,N_14321);
nand U14840 (N_14840,N_14092,N_14213);
nor U14841 (N_14841,N_14098,N_14313);
nor U14842 (N_14842,N_14293,N_13813);
nor U14843 (N_14843,N_13666,N_13992);
nand U14844 (N_14844,N_13974,N_13694);
nor U14845 (N_14845,N_14397,N_13845);
xor U14846 (N_14846,N_14392,N_13959);
and U14847 (N_14847,N_14188,N_13973);
and U14848 (N_14848,N_13778,N_13703);
and U14849 (N_14849,N_14069,N_14046);
xor U14850 (N_14850,N_14057,N_13756);
nor U14851 (N_14851,N_14370,N_13896);
or U14852 (N_14852,N_13741,N_13712);
and U14853 (N_14853,N_14352,N_13720);
and U14854 (N_14854,N_14041,N_13907);
xnor U14855 (N_14855,N_13992,N_14103);
and U14856 (N_14856,N_14386,N_13621);
or U14857 (N_14857,N_14198,N_13953);
or U14858 (N_14858,N_13978,N_14259);
and U14859 (N_14859,N_14262,N_14323);
nor U14860 (N_14860,N_13638,N_14172);
nand U14861 (N_14861,N_14138,N_14144);
and U14862 (N_14862,N_14135,N_14249);
or U14863 (N_14863,N_14258,N_14157);
nor U14864 (N_14864,N_13981,N_13722);
and U14865 (N_14865,N_14014,N_14169);
nor U14866 (N_14866,N_13813,N_13733);
nand U14867 (N_14867,N_14338,N_14265);
xor U14868 (N_14868,N_14286,N_13881);
nor U14869 (N_14869,N_14070,N_14364);
and U14870 (N_14870,N_13899,N_14398);
or U14871 (N_14871,N_14105,N_14234);
nand U14872 (N_14872,N_14198,N_13887);
and U14873 (N_14873,N_14084,N_14381);
xnor U14874 (N_14874,N_14066,N_13739);
xor U14875 (N_14875,N_14097,N_13879);
or U14876 (N_14876,N_13983,N_13851);
nor U14877 (N_14877,N_13953,N_14266);
and U14878 (N_14878,N_14398,N_14040);
nand U14879 (N_14879,N_14211,N_13840);
nor U14880 (N_14880,N_13626,N_14025);
xor U14881 (N_14881,N_13656,N_13852);
or U14882 (N_14882,N_14103,N_14061);
nor U14883 (N_14883,N_14361,N_14398);
or U14884 (N_14884,N_13973,N_13707);
xnor U14885 (N_14885,N_14191,N_13917);
xor U14886 (N_14886,N_14128,N_14022);
and U14887 (N_14887,N_14321,N_14126);
nand U14888 (N_14888,N_13665,N_14114);
and U14889 (N_14889,N_13754,N_14346);
and U14890 (N_14890,N_13981,N_14077);
nand U14891 (N_14891,N_14104,N_14129);
and U14892 (N_14892,N_14066,N_13982);
xor U14893 (N_14893,N_14013,N_13600);
or U14894 (N_14894,N_13830,N_14057);
nor U14895 (N_14895,N_13601,N_14175);
or U14896 (N_14896,N_14134,N_14245);
xnor U14897 (N_14897,N_14369,N_13750);
or U14898 (N_14898,N_14163,N_14195);
nand U14899 (N_14899,N_14156,N_14249);
or U14900 (N_14900,N_14115,N_13653);
and U14901 (N_14901,N_13968,N_13842);
or U14902 (N_14902,N_13978,N_14296);
or U14903 (N_14903,N_14051,N_13916);
or U14904 (N_14904,N_14347,N_13970);
nor U14905 (N_14905,N_14141,N_14322);
nor U14906 (N_14906,N_14066,N_14372);
nand U14907 (N_14907,N_13835,N_14169);
or U14908 (N_14908,N_13698,N_13735);
or U14909 (N_14909,N_14057,N_14225);
or U14910 (N_14910,N_13866,N_14115);
nor U14911 (N_14911,N_13738,N_13811);
or U14912 (N_14912,N_14220,N_14083);
and U14913 (N_14913,N_14126,N_14344);
nor U14914 (N_14914,N_14160,N_14374);
xnor U14915 (N_14915,N_13884,N_13657);
nand U14916 (N_14916,N_14362,N_13921);
nor U14917 (N_14917,N_14334,N_13937);
nor U14918 (N_14918,N_13917,N_13640);
or U14919 (N_14919,N_13636,N_14373);
xnor U14920 (N_14920,N_14245,N_14258);
nor U14921 (N_14921,N_14098,N_13920);
nor U14922 (N_14922,N_13960,N_14032);
or U14923 (N_14923,N_14331,N_14395);
or U14924 (N_14924,N_14308,N_14250);
nor U14925 (N_14925,N_13804,N_14233);
nand U14926 (N_14926,N_14057,N_14311);
nand U14927 (N_14927,N_13872,N_13867);
nor U14928 (N_14928,N_14027,N_13727);
nor U14929 (N_14929,N_14065,N_13844);
or U14930 (N_14930,N_14043,N_13767);
nor U14931 (N_14931,N_14273,N_13846);
and U14932 (N_14932,N_13852,N_13771);
or U14933 (N_14933,N_13989,N_13661);
and U14934 (N_14934,N_14325,N_14024);
and U14935 (N_14935,N_14162,N_13791);
or U14936 (N_14936,N_13913,N_13717);
xnor U14937 (N_14937,N_13688,N_13951);
or U14938 (N_14938,N_13871,N_14004);
xor U14939 (N_14939,N_13758,N_14322);
or U14940 (N_14940,N_14367,N_14265);
or U14941 (N_14941,N_14392,N_13672);
nor U14942 (N_14942,N_13916,N_13831);
nor U14943 (N_14943,N_14287,N_13839);
or U14944 (N_14944,N_13908,N_14271);
and U14945 (N_14945,N_13843,N_14209);
nor U14946 (N_14946,N_14202,N_13939);
xnor U14947 (N_14947,N_14230,N_13673);
nor U14948 (N_14948,N_13890,N_14300);
nor U14949 (N_14949,N_14197,N_13948);
or U14950 (N_14950,N_13902,N_13848);
and U14951 (N_14951,N_14398,N_13603);
or U14952 (N_14952,N_14124,N_13800);
nand U14953 (N_14953,N_13870,N_13742);
xor U14954 (N_14954,N_14179,N_13820);
or U14955 (N_14955,N_13823,N_13802);
and U14956 (N_14956,N_14131,N_13823);
xor U14957 (N_14957,N_14379,N_14046);
or U14958 (N_14958,N_14103,N_13775);
nor U14959 (N_14959,N_13839,N_14356);
or U14960 (N_14960,N_13852,N_14292);
or U14961 (N_14961,N_13950,N_14059);
and U14962 (N_14962,N_13756,N_13636);
or U14963 (N_14963,N_13952,N_13914);
and U14964 (N_14964,N_14112,N_13818);
nand U14965 (N_14965,N_14317,N_14180);
xnor U14966 (N_14966,N_14010,N_13770);
nand U14967 (N_14967,N_13705,N_13832);
and U14968 (N_14968,N_13836,N_14302);
or U14969 (N_14969,N_14298,N_14148);
xor U14970 (N_14970,N_13828,N_14188);
nand U14971 (N_14971,N_14005,N_13692);
nand U14972 (N_14972,N_14256,N_14356);
nand U14973 (N_14973,N_13838,N_13989);
xor U14974 (N_14974,N_13954,N_14394);
nor U14975 (N_14975,N_13978,N_14127);
xnor U14976 (N_14976,N_13724,N_13669);
nor U14977 (N_14977,N_13745,N_14367);
nand U14978 (N_14978,N_13748,N_13605);
and U14979 (N_14979,N_13922,N_13713);
nor U14980 (N_14980,N_14205,N_14165);
nor U14981 (N_14981,N_13761,N_14376);
nand U14982 (N_14982,N_14081,N_13733);
nand U14983 (N_14983,N_14135,N_14021);
nor U14984 (N_14984,N_13939,N_13626);
and U14985 (N_14985,N_13676,N_13711);
nor U14986 (N_14986,N_14192,N_13740);
and U14987 (N_14987,N_14079,N_13750);
nand U14988 (N_14988,N_14249,N_13778);
nand U14989 (N_14989,N_14330,N_14228);
or U14990 (N_14990,N_14016,N_14004);
xnor U14991 (N_14991,N_13892,N_13955);
and U14992 (N_14992,N_13821,N_13808);
and U14993 (N_14993,N_14363,N_13665);
and U14994 (N_14994,N_14358,N_14145);
nand U14995 (N_14995,N_13858,N_13857);
or U14996 (N_14996,N_14067,N_13969);
and U14997 (N_14997,N_14315,N_13817);
nor U14998 (N_14998,N_13750,N_13927);
and U14999 (N_14999,N_13828,N_13736);
nand U15000 (N_15000,N_14262,N_13692);
nand U15001 (N_15001,N_14398,N_13962);
nor U15002 (N_15002,N_14216,N_14072);
nand U15003 (N_15003,N_13662,N_14176);
and U15004 (N_15004,N_14298,N_13832);
nand U15005 (N_15005,N_13730,N_13866);
or U15006 (N_15006,N_13959,N_13615);
or U15007 (N_15007,N_14042,N_13897);
or U15008 (N_15008,N_14284,N_14157);
nor U15009 (N_15009,N_14061,N_13958);
nor U15010 (N_15010,N_13726,N_14171);
nor U15011 (N_15011,N_14075,N_14102);
or U15012 (N_15012,N_13967,N_13822);
and U15013 (N_15013,N_13667,N_13693);
or U15014 (N_15014,N_13959,N_13797);
nand U15015 (N_15015,N_14015,N_13924);
and U15016 (N_15016,N_13967,N_14192);
nand U15017 (N_15017,N_13725,N_13802);
nor U15018 (N_15018,N_13609,N_13622);
xor U15019 (N_15019,N_14357,N_14310);
xnor U15020 (N_15020,N_14308,N_13743);
nor U15021 (N_15021,N_13666,N_14045);
and U15022 (N_15022,N_14344,N_13990);
nor U15023 (N_15023,N_14127,N_14212);
nand U15024 (N_15024,N_13637,N_14380);
nor U15025 (N_15025,N_14092,N_13663);
xor U15026 (N_15026,N_14108,N_13995);
nor U15027 (N_15027,N_14324,N_13819);
nand U15028 (N_15028,N_13705,N_14328);
nand U15029 (N_15029,N_13755,N_14239);
nand U15030 (N_15030,N_14118,N_13842);
or U15031 (N_15031,N_14141,N_14330);
and U15032 (N_15032,N_14004,N_14243);
or U15033 (N_15033,N_14219,N_13825);
nor U15034 (N_15034,N_14372,N_14145);
or U15035 (N_15035,N_14067,N_13730);
and U15036 (N_15036,N_14022,N_14380);
nand U15037 (N_15037,N_14300,N_13922);
nor U15038 (N_15038,N_14228,N_14181);
nand U15039 (N_15039,N_13732,N_14030);
xnor U15040 (N_15040,N_13956,N_14333);
or U15041 (N_15041,N_14015,N_14129);
nor U15042 (N_15042,N_14273,N_14059);
or U15043 (N_15043,N_13835,N_13727);
nor U15044 (N_15044,N_13735,N_14106);
or U15045 (N_15045,N_13826,N_14147);
and U15046 (N_15046,N_14167,N_13720);
nand U15047 (N_15047,N_14128,N_14294);
and U15048 (N_15048,N_13638,N_13964);
or U15049 (N_15049,N_14366,N_14092);
nand U15050 (N_15050,N_13841,N_13918);
xnor U15051 (N_15051,N_13812,N_13930);
or U15052 (N_15052,N_13630,N_13773);
nor U15053 (N_15053,N_13894,N_13997);
nor U15054 (N_15054,N_14347,N_13863);
nand U15055 (N_15055,N_14151,N_14368);
and U15056 (N_15056,N_13774,N_14396);
nand U15057 (N_15057,N_13654,N_14045);
xor U15058 (N_15058,N_13715,N_13995);
nor U15059 (N_15059,N_13832,N_14033);
nor U15060 (N_15060,N_13751,N_13691);
nor U15061 (N_15061,N_14055,N_14193);
and U15062 (N_15062,N_13857,N_14125);
and U15063 (N_15063,N_13675,N_14195);
nor U15064 (N_15064,N_14312,N_14245);
xor U15065 (N_15065,N_14149,N_13889);
or U15066 (N_15066,N_14253,N_14194);
xnor U15067 (N_15067,N_13960,N_14334);
or U15068 (N_15068,N_14076,N_13862);
or U15069 (N_15069,N_13826,N_14098);
or U15070 (N_15070,N_14035,N_13931);
or U15071 (N_15071,N_14082,N_13935);
nand U15072 (N_15072,N_14169,N_14204);
and U15073 (N_15073,N_14229,N_14065);
and U15074 (N_15074,N_13995,N_14278);
and U15075 (N_15075,N_13991,N_13737);
or U15076 (N_15076,N_14004,N_14003);
nor U15077 (N_15077,N_14259,N_13713);
and U15078 (N_15078,N_13642,N_14074);
or U15079 (N_15079,N_14266,N_14118);
nor U15080 (N_15080,N_13715,N_13835);
nand U15081 (N_15081,N_13701,N_13749);
or U15082 (N_15082,N_14067,N_14149);
nand U15083 (N_15083,N_14200,N_14321);
or U15084 (N_15084,N_14225,N_14251);
xor U15085 (N_15085,N_14039,N_14316);
nor U15086 (N_15086,N_13769,N_13659);
nor U15087 (N_15087,N_13812,N_13670);
or U15088 (N_15088,N_14309,N_14325);
xnor U15089 (N_15089,N_13988,N_14125);
and U15090 (N_15090,N_14215,N_13693);
nor U15091 (N_15091,N_13825,N_14263);
nand U15092 (N_15092,N_13892,N_13607);
nor U15093 (N_15093,N_13964,N_14005);
nor U15094 (N_15094,N_14293,N_14278);
xor U15095 (N_15095,N_14193,N_13744);
nand U15096 (N_15096,N_13839,N_14388);
and U15097 (N_15097,N_13931,N_14227);
and U15098 (N_15098,N_13954,N_14331);
nand U15099 (N_15099,N_13906,N_13623);
and U15100 (N_15100,N_14157,N_13686);
nor U15101 (N_15101,N_13863,N_14398);
nor U15102 (N_15102,N_13933,N_14142);
and U15103 (N_15103,N_14082,N_14047);
xnor U15104 (N_15104,N_13681,N_14396);
nand U15105 (N_15105,N_14193,N_14152);
nand U15106 (N_15106,N_13724,N_14178);
xnor U15107 (N_15107,N_14115,N_14085);
and U15108 (N_15108,N_14268,N_13671);
or U15109 (N_15109,N_13877,N_13850);
and U15110 (N_15110,N_14376,N_13877);
or U15111 (N_15111,N_14297,N_13873);
or U15112 (N_15112,N_13656,N_13965);
xnor U15113 (N_15113,N_13632,N_13668);
nor U15114 (N_15114,N_13829,N_14152);
and U15115 (N_15115,N_13865,N_14145);
and U15116 (N_15116,N_13741,N_14068);
xor U15117 (N_15117,N_14209,N_14033);
xnor U15118 (N_15118,N_13883,N_14101);
nor U15119 (N_15119,N_14088,N_13624);
xor U15120 (N_15120,N_13991,N_14037);
xor U15121 (N_15121,N_14142,N_14327);
or U15122 (N_15122,N_13868,N_14056);
xnor U15123 (N_15123,N_13747,N_14328);
nand U15124 (N_15124,N_13688,N_13830);
xor U15125 (N_15125,N_14347,N_13632);
nand U15126 (N_15126,N_13965,N_14053);
xnor U15127 (N_15127,N_14066,N_13618);
and U15128 (N_15128,N_13743,N_13842);
nand U15129 (N_15129,N_13748,N_14016);
and U15130 (N_15130,N_13932,N_14123);
xnor U15131 (N_15131,N_13883,N_13694);
nand U15132 (N_15132,N_14364,N_13770);
nor U15133 (N_15133,N_14070,N_14115);
and U15134 (N_15134,N_13835,N_14033);
and U15135 (N_15135,N_14009,N_14391);
or U15136 (N_15136,N_13725,N_13899);
or U15137 (N_15137,N_13645,N_13681);
or U15138 (N_15138,N_14178,N_14000);
nand U15139 (N_15139,N_14174,N_13943);
nor U15140 (N_15140,N_14277,N_14159);
xnor U15141 (N_15141,N_13711,N_14355);
nor U15142 (N_15142,N_13847,N_14067);
or U15143 (N_15143,N_14293,N_14234);
or U15144 (N_15144,N_13947,N_14363);
or U15145 (N_15145,N_13992,N_14115);
or U15146 (N_15146,N_13785,N_14053);
and U15147 (N_15147,N_13742,N_14061);
nand U15148 (N_15148,N_14063,N_13967);
nor U15149 (N_15149,N_13837,N_13633);
or U15150 (N_15150,N_14150,N_14121);
xor U15151 (N_15151,N_13945,N_13838);
nor U15152 (N_15152,N_13798,N_14029);
xnor U15153 (N_15153,N_13659,N_13810);
or U15154 (N_15154,N_14330,N_13674);
or U15155 (N_15155,N_14287,N_13930);
and U15156 (N_15156,N_13852,N_14118);
and U15157 (N_15157,N_14153,N_14347);
and U15158 (N_15158,N_13999,N_14157);
xnor U15159 (N_15159,N_14076,N_13746);
nor U15160 (N_15160,N_13870,N_14218);
or U15161 (N_15161,N_14088,N_14245);
nand U15162 (N_15162,N_13637,N_14059);
nand U15163 (N_15163,N_14067,N_13972);
xor U15164 (N_15164,N_14373,N_13791);
and U15165 (N_15165,N_13821,N_14398);
or U15166 (N_15166,N_13887,N_14074);
nand U15167 (N_15167,N_13743,N_14103);
nor U15168 (N_15168,N_14387,N_14120);
and U15169 (N_15169,N_13969,N_13905);
xor U15170 (N_15170,N_14053,N_13797);
xor U15171 (N_15171,N_14279,N_14128);
xor U15172 (N_15172,N_14006,N_14117);
or U15173 (N_15173,N_13774,N_14252);
or U15174 (N_15174,N_13817,N_13651);
or U15175 (N_15175,N_13731,N_14134);
and U15176 (N_15176,N_13691,N_13749);
nor U15177 (N_15177,N_13675,N_13848);
and U15178 (N_15178,N_13989,N_14327);
nor U15179 (N_15179,N_14294,N_13639);
or U15180 (N_15180,N_14366,N_14296);
xor U15181 (N_15181,N_14283,N_13882);
nand U15182 (N_15182,N_14266,N_13858);
nor U15183 (N_15183,N_13931,N_14004);
nor U15184 (N_15184,N_13639,N_14270);
nand U15185 (N_15185,N_13828,N_13727);
nor U15186 (N_15186,N_14200,N_14184);
nor U15187 (N_15187,N_14356,N_14358);
nand U15188 (N_15188,N_14043,N_14050);
nand U15189 (N_15189,N_14304,N_14344);
or U15190 (N_15190,N_14079,N_14003);
nor U15191 (N_15191,N_13911,N_13616);
nand U15192 (N_15192,N_14155,N_14271);
or U15193 (N_15193,N_13931,N_14169);
nand U15194 (N_15194,N_14306,N_14027);
xnor U15195 (N_15195,N_14011,N_13771);
nor U15196 (N_15196,N_14000,N_13683);
and U15197 (N_15197,N_13952,N_13610);
nand U15198 (N_15198,N_14257,N_14146);
nor U15199 (N_15199,N_13962,N_14145);
nand U15200 (N_15200,N_14664,N_14491);
nor U15201 (N_15201,N_14711,N_15174);
nor U15202 (N_15202,N_15062,N_14731);
nand U15203 (N_15203,N_14983,N_14428);
xnor U15204 (N_15204,N_15118,N_15141);
or U15205 (N_15205,N_14508,N_14586);
or U15206 (N_15206,N_14478,N_15074);
xor U15207 (N_15207,N_14781,N_14774);
xor U15208 (N_15208,N_14997,N_14492);
nand U15209 (N_15209,N_14582,N_14990);
nor U15210 (N_15210,N_14622,N_15083);
nand U15211 (N_15211,N_14653,N_14797);
or U15212 (N_15212,N_14982,N_14724);
nor U15213 (N_15213,N_15167,N_14457);
nand U15214 (N_15214,N_14544,N_15137);
nand U15215 (N_15215,N_15047,N_14908);
or U15216 (N_15216,N_14907,N_14896);
nand U15217 (N_15217,N_14688,N_14686);
xor U15218 (N_15218,N_14779,N_14580);
nand U15219 (N_15219,N_14537,N_14937);
nor U15220 (N_15220,N_14723,N_15182);
and U15221 (N_15221,N_14803,N_14490);
or U15222 (N_15222,N_14484,N_14528);
nor U15223 (N_15223,N_14561,N_14941);
or U15224 (N_15224,N_15034,N_15181);
and U15225 (N_15225,N_15040,N_14634);
and U15226 (N_15226,N_15091,N_15070);
or U15227 (N_15227,N_14863,N_14577);
xnor U15228 (N_15228,N_14898,N_15159);
or U15229 (N_15229,N_14402,N_14851);
nand U15230 (N_15230,N_14887,N_14871);
nor U15231 (N_15231,N_14938,N_14600);
or U15232 (N_15232,N_14575,N_14784);
or U15233 (N_15233,N_15188,N_15116);
nand U15234 (N_15234,N_15021,N_14764);
nand U15235 (N_15235,N_14595,N_14917);
or U15236 (N_15236,N_14685,N_15196);
xnor U15237 (N_15237,N_14864,N_15102);
nand U15238 (N_15238,N_14885,N_15162);
nor U15239 (N_15239,N_14444,N_15052);
nand U15240 (N_15240,N_15148,N_14429);
nand U15241 (N_15241,N_15095,N_14909);
nor U15242 (N_15242,N_14737,N_15146);
or U15243 (N_15243,N_14424,N_14667);
nor U15244 (N_15244,N_15061,N_15123);
and U15245 (N_15245,N_14465,N_14649);
or U15246 (N_15246,N_15112,N_14924);
and U15247 (N_15247,N_14981,N_15036);
or U15248 (N_15248,N_14999,N_14929);
or U15249 (N_15249,N_15059,N_15066);
xor U15250 (N_15250,N_14963,N_15176);
xor U15251 (N_15251,N_14936,N_14785);
nor U15252 (N_15252,N_14902,N_14692);
xnor U15253 (N_15253,N_15084,N_14472);
or U15254 (N_15254,N_14978,N_14827);
nand U15255 (N_15255,N_14921,N_14932);
or U15256 (N_15256,N_14629,N_14609);
and U15257 (N_15257,N_14900,N_14624);
or U15258 (N_15258,N_14494,N_15138);
or U15259 (N_15259,N_14670,N_14695);
nor U15260 (N_15260,N_15120,N_15111);
and U15261 (N_15261,N_14651,N_14893);
or U15262 (N_15262,N_15145,N_14509);
nor U15263 (N_15263,N_14862,N_15004);
or U15264 (N_15264,N_15133,N_15071);
nor U15265 (N_15265,N_14989,N_14748);
or U15266 (N_15266,N_15173,N_14480);
xnor U15267 (N_15267,N_15177,N_14733);
and U15268 (N_15268,N_15122,N_14794);
or U15269 (N_15269,N_14698,N_15086);
or U15270 (N_15270,N_15101,N_15092);
and U15271 (N_15271,N_14845,N_14534);
nand U15272 (N_15272,N_14466,N_14625);
xor U15273 (N_15273,N_15171,N_14881);
and U15274 (N_15274,N_14884,N_14880);
nand U15275 (N_15275,N_15183,N_14599);
nor U15276 (N_15276,N_14959,N_14601);
nor U15277 (N_15277,N_15073,N_14894);
nor U15278 (N_15278,N_14957,N_15000);
nor U15279 (N_15279,N_14975,N_14713);
and U15280 (N_15280,N_14453,N_15166);
and U15281 (N_15281,N_15158,N_15128);
or U15282 (N_15282,N_15168,N_14955);
and U15283 (N_15283,N_15076,N_14858);
nand U15284 (N_15284,N_15081,N_14883);
nand U15285 (N_15285,N_14861,N_14451);
nand U15286 (N_15286,N_14886,N_14656);
nand U15287 (N_15287,N_15117,N_14801);
xor U15288 (N_15288,N_14627,N_15089);
and U15289 (N_15289,N_14942,N_15178);
nor U15290 (N_15290,N_14571,N_15078);
xor U15291 (N_15291,N_14765,N_14931);
nand U15292 (N_15292,N_15015,N_14682);
or U15293 (N_15293,N_14901,N_14510);
or U15294 (N_15294,N_14549,N_14523);
nand U15295 (N_15295,N_14842,N_14768);
or U15296 (N_15296,N_14565,N_14888);
and U15297 (N_15297,N_14965,N_15119);
xnor U15298 (N_15298,N_14538,N_14507);
xor U15299 (N_15299,N_15053,N_14837);
nor U15300 (N_15300,N_14690,N_14714);
or U15301 (N_15301,N_14977,N_14961);
nand U15302 (N_15302,N_14469,N_14805);
and U15303 (N_15303,N_15049,N_14721);
or U15304 (N_15304,N_15050,N_14922);
and U15305 (N_15305,N_14436,N_14889);
xnor U15306 (N_15306,N_15014,N_14743);
nor U15307 (N_15307,N_15032,N_15115);
nor U15308 (N_15308,N_14503,N_14758);
nand U15309 (N_15309,N_14694,N_14705);
and U15310 (N_15310,N_14786,N_14432);
xor U15311 (N_15311,N_15063,N_14867);
or U15312 (N_15312,N_14829,N_14587);
nand U15313 (N_15313,N_14869,N_15189);
and U15314 (N_15314,N_14822,N_14573);
or U15315 (N_15315,N_14590,N_14488);
xor U15316 (N_15316,N_15008,N_14811);
xnor U15317 (N_15317,N_15108,N_14594);
and U15318 (N_15318,N_14497,N_14952);
or U15319 (N_15319,N_15184,N_15042);
nand U15320 (N_15320,N_14521,N_14654);
and U15321 (N_15321,N_14736,N_14915);
xnor U15322 (N_15322,N_14584,N_15194);
nand U15323 (N_15323,N_14740,N_14415);
nor U15324 (N_15324,N_14559,N_14495);
xor U15325 (N_15325,N_15025,N_14400);
xor U15326 (N_15326,N_15067,N_15163);
xor U15327 (N_15327,N_14772,N_14535);
and U15328 (N_15328,N_14671,N_14461);
and U15329 (N_15329,N_14430,N_14483);
xor U15330 (N_15330,N_14669,N_14854);
nor U15331 (N_15331,N_15124,N_14683);
nand U15332 (N_15332,N_14536,N_15149);
or U15333 (N_15333,N_14789,N_14741);
nor U15334 (N_15334,N_14834,N_14940);
nand U15335 (N_15335,N_14707,N_14646);
nor U15336 (N_15336,N_14993,N_15097);
and U15337 (N_15337,N_14603,N_14852);
xor U15338 (N_15338,N_14767,N_15153);
nand U15339 (N_15339,N_14916,N_14447);
xnor U15340 (N_15340,N_15191,N_14673);
and U15341 (N_15341,N_14910,N_14550);
xor U15342 (N_15342,N_15035,N_15164);
and U15343 (N_15343,N_14529,N_14793);
or U15344 (N_15344,N_14579,N_14742);
nand U15345 (N_15345,N_14712,N_14663);
xnor U15346 (N_15346,N_14477,N_15170);
and U15347 (N_15347,N_14404,N_14820);
and U15348 (N_15348,N_14816,N_14652);
nor U15349 (N_15349,N_14882,N_14807);
nor U15350 (N_15350,N_14558,N_15156);
xnor U15351 (N_15351,N_14876,N_14897);
nor U15352 (N_15352,N_14605,N_15033);
or U15353 (N_15353,N_15088,N_15020);
nand U15354 (N_15354,N_14496,N_14514);
nand U15355 (N_15355,N_14914,N_14847);
and U15356 (N_15356,N_14833,N_14777);
nand U15357 (N_15357,N_14425,N_15093);
and U15358 (N_15358,N_14499,N_14744);
and U15359 (N_15359,N_15130,N_14527);
nor U15360 (N_15360,N_15131,N_15142);
nor U15361 (N_15361,N_14419,N_14979);
or U15362 (N_15362,N_14788,N_14623);
and U15363 (N_15363,N_15030,N_14524);
or U15364 (N_15364,N_15151,N_14420);
nand U15365 (N_15365,N_15085,N_15022);
nor U15366 (N_15366,N_14546,N_14417);
or U15367 (N_15367,N_15126,N_14968);
nor U15368 (N_15368,N_15127,N_14626);
nand U15369 (N_15369,N_14679,N_15080);
and U15370 (N_15370,N_14530,N_14870);
and U15371 (N_15371,N_14872,N_14589);
nor U15372 (N_15372,N_14762,N_14776);
nand U15373 (N_15373,N_14442,N_14591);
and U15374 (N_15374,N_14541,N_14547);
xor U15375 (N_15375,N_14554,N_14895);
or U15376 (N_15376,N_14645,N_14746);
xor U15377 (N_15377,N_14439,N_14734);
or U15378 (N_15378,N_14855,N_14755);
and U15379 (N_15379,N_14440,N_15024);
xnor U15380 (N_15380,N_14951,N_15099);
and U15381 (N_15381,N_15185,N_15154);
and U15382 (N_15382,N_14602,N_14569);
nand U15383 (N_15383,N_14906,N_14452);
nand U15384 (N_15384,N_14630,N_14966);
nand U15385 (N_15385,N_14751,N_14944);
and U15386 (N_15386,N_15140,N_15028);
xnor U15387 (N_15387,N_14504,N_14403);
xor U15388 (N_15388,N_14726,N_14771);
nor U15389 (N_15389,N_14703,N_15172);
xor U15390 (N_15390,N_14641,N_14954);
or U15391 (N_15391,N_14681,N_14747);
or U15392 (N_15392,N_14950,N_14552);
and U15393 (N_15393,N_14572,N_14502);
and U15394 (N_15394,N_15079,N_14735);
xnor U15395 (N_15395,N_14775,N_14581);
xor U15396 (N_15396,N_14819,N_14874);
or U15397 (N_15397,N_14647,N_14435);
or U15398 (N_15398,N_14935,N_15017);
nor U15399 (N_15399,N_15075,N_14865);
nor U15400 (N_15400,N_14574,N_14866);
nand U15401 (N_15401,N_14525,N_15143);
or U15402 (N_15402,N_14891,N_14700);
and U15403 (N_15403,N_14610,N_14505);
and U15404 (N_15404,N_14551,N_14918);
nor U15405 (N_15405,N_14704,N_14548);
xor U15406 (N_15406,N_14640,N_14405);
and U15407 (N_15407,N_14782,N_14846);
xor U15408 (N_15408,N_15106,N_14970);
or U15409 (N_15409,N_14719,N_14680);
and U15410 (N_15410,N_14443,N_15011);
nor U15411 (N_15411,N_15013,N_14543);
or U15412 (N_15412,N_14516,N_14665);
nand U15413 (N_15413,N_14976,N_15002);
nor U15414 (N_15414,N_14542,N_14621);
nand U15415 (N_15415,N_14754,N_14716);
and U15416 (N_15416,N_14696,N_15190);
or U15417 (N_15417,N_14556,N_14658);
xnor U15418 (N_15418,N_14446,N_14585);
nand U15419 (N_15419,N_14596,N_14564);
nor U15420 (N_15420,N_14422,N_14994);
nand U15421 (N_15421,N_15056,N_14969);
and U15422 (N_15422,N_14826,N_14953);
nand U15423 (N_15423,N_14738,N_15039);
or U15424 (N_15424,N_14401,N_15057);
nand U15425 (N_15425,N_14838,N_14661);
and U15426 (N_15426,N_14974,N_15087);
nand U15427 (N_15427,N_15121,N_14848);
xnor U15428 (N_15428,N_14947,N_14956);
and U15429 (N_15429,N_14410,N_14701);
nand U15430 (N_15430,N_14666,N_14433);
nand U15431 (N_15431,N_14455,N_14449);
and U15432 (N_15432,N_14583,N_14844);
xnor U15433 (N_15433,N_14821,N_14780);
and U15434 (N_15434,N_14948,N_14482);
nor U15435 (N_15435,N_14612,N_14412);
nand U15436 (N_15436,N_14857,N_15027);
and U15437 (N_15437,N_14684,N_15179);
xor U15438 (N_15438,N_15150,N_14792);
xor U15439 (N_15439,N_14506,N_15100);
and U15440 (N_15440,N_14644,N_14557);
or U15441 (N_15441,N_14739,N_15007);
and U15442 (N_15442,N_15187,N_14729);
and U15443 (N_15443,N_14973,N_14423);
nand U15444 (N_15444,N_14642,N_14562);
nand U15445 (N_15445,N_14568,N_14996);
or U15446 (N_15446,N_14710,N_14843);
nand U15447 (N_15447,N_14464,N_15051);
nor U15448 (N_15448,N_15136,N_14806);
nand U15449 (N_15449,N_14725,N_15135);
nand U15450 (N_15450,N_14840,N_14905);
nor U15451 (N_15451,N_14759,N_14727);
xor U15452 (N_15452,N_14409,N_15103);
nand U15453 (N_15453,N_14745,N_14998);
nor U15454 (N_15454,N_14675,N_14836);
xnor U15455 (N_15455,N_14462,N_14824);
nor U15456 (N_15456,N_14413,N_14615);
and U15457 (N_15457,N_15038,N_14613);
and U15458 (N_15458,N_14949,N_14408);
nand U15459 (N_15459,N_14835,N_14545);
xor U15460 (N_15460,N_14431,N_14791);
and U15461 (N_15461,N_14459,N_14945);
or U15462 (N_15462,N_14672,N_15110);
or U15463 (N_15463,N_14454,N_14643);
and U15464 (N_15464,N_15068,N_14414);
or U15465 (N_15465,N_14407,N_15144);
xor U15466 (N_15466,N_14783,N_14438);
nor U15467 (N_15467,N_14606,N_14512);
and U15468 (N_15468,N_14798,N_15105);
xor U15469 (N_15469,N_14511,N_14814);
and U15470 (N_15470,N_14920,N_14912);
and U15471 (N_15471,N_15160,N_14849);
nor U15472 (N_15472,N_14540,N_14567);
xnor U15473 (N_15473,N_14728,N_15104);
nand U15474 (N_15474,N_15003,N_14992);
nand U15475 (N_15475,N_14892,N_14850);
or U15476 (N_15476,N_14608,N_14445);
nand U15477 (N_15477,N_14639,N_14633);
xnor U15478 (N_15478,N_15109,N_14533);
nor U15479 (N_15479,N_14632,N_14971);
or U15480 (N_15480,N_14903,N_14720);
xnor U15481 (N_15481,N_14563,N_15058);
and U15482 (N_15482,N_15046,N_15195);
and U15483 (N_15483,N_14611,N_14578);
and U15484 (N_15484,N_15029,N_14810);
nand U15485 (N_15485,N_14473,N_14750);
nand U15486 (N_15486,N_14717,N_14927);
nor U15487 (N_15487,N_15044,N_14987);
or U15488 (N_15488,N_14986,N_14868);
nand U15489 (N_15489,N_14732,N_15129);
or U15490 (N_15490,N_14487,N_14699);
nor U15491 (N_15491,N_14925,N_14839);
or U15492 (N_15492,N_15125,N_14479);
nor U15493 (N_15493,N_15082,N_14662);
and U15494 (N_15494,N_14617,N_14962);
nand U15495 (N_15495,N_14809,N_15005);
xnor U15496 (N_15496,N_15037,N_14448);
nand U15497 (N_15497,N_14458,N_15114);
xnor U15498 (N_15498,N_14718,N_14702);
and U15499 (N_15499,N_15113,N_15175);
nand U15500 (N_15500,N_14481,N_14756);
nand U15501 (N_15501,N_14960,N_14598);
nand U15502 (N_15502,N_14877,N_14566);
xnor U15503 (N_15503,N_14856,N_14800);
or U15504 (N_15504,N_15077,N_15098);
and U15505 (N_15505,N_15090,N_14620);
and U15506 (N_15506,N_14946,N_14830);
or U15507 (N_15507,N_15161,N_14531);
and U15508 (N_15508,N_14486,N_14787);
xnor U15509 (N_15509,N_14468,N_14674);
nor U15510 (N_15510,N_14657,N_14539);
or U15511 (N_15511,N_14555,N_14919);
and U15512 (N_15512,N_14763,N_15019);
xnor U15513 (N_15513,N_14678,N_14501);
and U15514 (N_15514,N_15147,N_14616);
xor U15515 (N_15515,N_15169,N_14930);
xor U15516 (N_15516,N_14655,N_15043);
or U15517 (N_15517,N_14676,N_15016);
or U15518 (N_15518,N_15155,N_14752);
nor U15519 (N_15519,N_14796,N_14689);
and U15520 (N_15520,N_14421,N_14463);
or U15521 (N_15521,N_15107,N_14709);
nor U15522 (N_15522,N_14708,N_14722);
nand U15523 (N_15523,N_14493,N_14899);
nand U15524 (N_15524,N_14434,N_14437);
nand U15525 (N_15525,N_14659,N_14697);
nand U15526 (N_15526,N_14770,N_15134);
and U15527 (N_15527,N_15165,N_15199);
and U15528 (N_15528,N_14532,N_14879);
nor U15529 (N_15529,N_15031,N_14456);
nor U15530 (N_15530,N_14753,N_14964);
nor U15531 (N_15531,N_14677,N_14660);
nor U15532 (N_15532,N_14831,N_15193);
xnor U15533 (N_15533,N_14985,N_14650);
nor U15534 (N_15534,N_15152,N_14859);
nand U15535 (N_15535,N_14878,N_14607);
or U15536 (N_15536,N_15055,N_14825);
nor U15537 (N_15537,N_15197,N_14904);
xor U15538 (N_15538,N_14967,N_14687);
and U15539 (N_15539,N_14778,N_14635);
nor U15540 (N_15540,N_14873,N_14604);
nor U15541 (N_15541,N_14426,N_15069);
or U15542 (N_15542,N_14588,N_15054);
xor U15543 (N_15543,N_14790,N_14757);
nor U15544 (N_15544,N_14513,N_14991);
xor U15545 (N_15545,N_14766,N_14812);
nand U15546 (N_15546,N_15010,N_14926);
and U15547 (N_15547,N_15009,N_14933);
or U15548 (N_15548,N_14911,N_15139);
nand U15549 (N_15549,N_14648,N_14485);
nand U15550 (N_15550,N_14804,N_14406);
nand U15551 (N_15551,N_14972,N_15018);
or U15552 (N_15552,N_14934,N_14560);
or U15553 (N_15553,N_15023,N_15048);
nand U15554 (N_15554,N_14853,N_14637);
or U15555 (N_15555,N_14619,N_14427);
and U15556 (N_15556,N_14636,N_14470);
or U15557 (N_15557,N_14411,N_15012);
or U15558 (N_15558,N_14795,N_14693);
or U15559 (N_15559,N_14988,N_14519);
xor U15560 (N_15560,N_14761,N_14802);
or U15561 (N_15561,N_14614,N_14730);
nor U15562 (N_15562,N_14517,N_15072);
and U15563 (N_15563,N_14691,N_14769);
nand U15564 (N_15564,N_15192,N_14943);
nor U15565 (N_15565,N_14832,N_14441);
nand U15566 (N_15566,N_14489,N_14498);
or U15567 (N_15567,N_15041,N_14749);
or U15568 (N_15568,N_15180,N_15064);
or U15569 (N_15569,N_14875,N_15096);
and U15570 (N_15570,N_15026,N_14476);
or U15571 (N_15571,N_14467,N_14841);
nor U15572 (N_15572,N_14576,N_14815);
or U15573 (N_15573,N_14474,N_15132);
nand U15574 (N_15574,N_15186,N_14631);
nor U15575 (N_15575,N_14773,N_14418);
and U15576 (N_15576,N_14518,N_14760);
xnor U15577 (N_15577,N_14939,N_14823);
or U15578 (N_15578,N_14475,N_14553);
xor U15579 (N_15579,N_15060,N_14416);
and U15580 (N_15580,N_14923,N_14715);
and U15581 (N_15581,N_15065,N_14913);
and U15582 (N_15582,N_14860,N_14799);
nand U15583 (N_15583,N_14628,N_14618);
nor U15584 (N_15584,N_14593,N_14500);
xnor U15585 (N_15585,N_15157,N_14980);
xnor U15586 (N_15586,N_14928,N_15001);
nor U15587 (N_15587,N_14808,N_15198);
nor U15588 (N_15588,N_14818,N_14813);
xnor U15589 (N_15589,N_14471,N_14597);
nand U15590 (N_15590,N_14890,N_14668);
and U15591 (N_15591,N_14526,N_14706);
nor U15592 (N_15592,N_14570,N_14958);
nand U15593 (N_15593,N_14592,N_14460);
xnor U15594 (N_15594,N_14450,N_14995);
nor U15595 (N_15595,N_15045,N_15006);
nand U15596 (N_15596,N_14520,N_14638);
nand U15597 (N_15597,N_14984,N_14522);
xor U15598 (N_15598,N_14817,N_14515);
xor U15599 (N_15599,N_14828,N_15094);
nor U15600 (N_15600,N_14620,N_15025);
and U15601 (N_15601,N_14749,N_14830);
nor U15602 (N_15602,N_14556,N_14520);
nand U15603 (N_15603,N_14458,N_15142);
nand U15604 (N_15604,N_14593,N_14621);
nor U15605 (N_15605,N_14596,N_14753);
nor U15606 (N_15606,N_14799,N_14499);
and U15607 (N_15607,N_14632,N_14442);
xor U15608 (N_15608,N_14824,N_14613);
xor U15609 (N_15609,N_15092,N_15021);
xor U15610 (N_15610,N_15104,N_15137);
xor U15611 (N_15611,N_15069,N_15061);
nor U15612 (N_15612,N_14428,N_14405);
nand U15613 (N_15613,N_15140,N_14433);
and U15614 (N_15614,N_15145,N_14678);
nand U15615 (N_15615,N_14982,N_15010);
nand U15616 (N_15616,N_14475,N_15185);
nor U15617 (N_15617,N_14428,N_14739);
xnor U15618 (N_15618,N_14501,N_14715);
nand U15619 (N_15619,N_14984,N_14519);
nand U15620 (N_15620,N_15106,N_14956);
nand U15621 (N_15621,N_14479,N_15158);
or U15622 (N_15622,N_14939,N_14650);
and U15623 (N_15623,N_14863,N_14576);
and U15624 (N_15624,N_14851,N_14578);
nand U15625 (N_15625,N_15059,N_15122);
nand U15626 (N_15626,N_15046,N_14791);
nor U15627 (N_15627,N_14870,N_15114);
xnor U15628 (N_15628,N_14722,N_15114);
and U15629 (N_15629,N_14648,N_14723);
xnor U15630 (N_15630,N_15160,N_14722);
nor U15631 (N_15631,N_15054,N_14582);
and U15632 (N_15632,N_14464,N_14960);
xor U15633 (N_15633,N_15128,N_15117);
nand U15634 (N_15634,N_15134,N_15030);
or U15635 (N_15635,N_15012,N_14414);
and U15636 (N_15636,N_14789,N_14882);
or U15637 (N_15637,N_15120,N_14907);
or U15638 (N_15638,N_14742,N_14854);
or U15639 (N_15639,N_14651,N_15078);
xor U15640 (N_15640,N_14790,N_14811);
or U15641 (N_15641,N_14932,N_15013);
nand U15642 (N_15642,N_14572,N_14642);
or U15643 (N_15643,N_14724,N_14818);
nand U15644 (N_15644,N_14517,N_14872);
nor U15645 (N_15645,N_14638,N_14631);
nor U15646 (N_15646,N_14681,N_14452);
nand U15647 (N_15647,N_14546,N_14407);
nand U15648 (N_15648,N_14894,N_14714);
nand U15649 (N_15649,N_14714,N_14408);
nor U15650 (N_15650,N_14721,N_15108);
nand U15651 (N_15651,N_14809,N_15064);
xor U15652 (N_15652,N_14714,N_14553);
nor U15653 (N_15653,N_14557,N_14540);
xor U15654 (N_15654,N_14644,N_14797);
nand U15655 (N_15655,N_14583,N_14760);
and U15656 (N_15656,N_15049,N_14920);
and U15657 (N_15657,N_15004,N_14886);
xor U15658 (N_15658,N_14876,N_14966);
or U15659 (N_15659,N_14668,N_15084);
xnor U15660 (N_15660,N_14570,N_14438);
xor U15661 (N_15661,N_14860,N_14967);
nand U15662 (N_15662,N_14691,N_15077);
xor U15663 (N_15663,N_14914,N_14628);
or U15664 (N_15664,N_14710,N_15141);
and U15665 (N_15665,N_14529,N_14648);
xor U15666 (N_15666,N_14417,N_15010);
and U15667 (N_15667,N_14740,N_15081);
nand U15668 (N_15668,N_14426,N_14945);
xor U15669 (N_15669,N_14941,N_14501);
xnor U15670 (N_15670,N_14821,N_14848);
nor U15671 (N_15671,N_14993,N_14882);
nor U15672 (N_15672,N_14422,N_14883);
nor U15673 (N_15673,N_14423,N_14681);
and U15674 (N_15674,N_14663,N_14614);
or U15675 (N_15675,N_15136,N_14736);
or U15676 (N_15676,N_14487,N_14868);
or U15677 (N_15677,N_15177,N_14740);
nand U15678 (N_15678,N_15035,N_14434);
nand U15679 (N_15679,N_15148,N_14624);
nand U15680 (N_15680,N_14975,N_14532);
or U15681 (N_15681,N_15041,N_14639);
and U15682 (N_15682,N_14876,N_14651);
or U15683 (N_15683,N_14715,N_14778);
xnor U15684 (N_15684,N_15039,N_14629);
and U15685 (N_15685,N_14549,N_15009);
or U15686 (N_15686,N_15084,N_14982);
xor U15687 (N_15687,N_14993,N_14713);
xor U15688 (N_15688,N_14797,N_14648);
xor U15689 (N_15689,N_14986,N_14643);
nand U15690 (N_15690,N_14804,N_14777);
and U15691 (N_15691,N_14967,N_14905);
xor U15692 (N_15692,N_15107,N_14493);
and U15693 (N_15693,N_14624,N_14779);
xor U15694 (N_15694,N_14664,N_14662);
nor U15695 (N_15695,N_15092,N_15064);
nor U15696 (N_15696,N_14904,N_15003);
nor U15697 (N_15697,N_14834,N_14806);
nand U15698 (N_15698,N_14995,N_14514);
xnor U15699 (N_15699,N_14622,N_15150);
and U15700 (N_15700,N_14693,N_14845);
nor U15701 (N_15701,N_14859,N_14501);
nor U15702 (N_15702,N_14967,N_14483);
xor U15703 (N_15703,N_14802,N_14678);
nand U15704 (N_15704,N_15123,N_14440);
xnor U15705 (N_15705,N_14576,N_14948);
or U15706 (N_15706,N_14725,N_14744);
or U15707 (N_15707,N_14855,N_15064);
and U15708 (N_15708,N_14870,N_14747);
nand U15709 (N_15709,N_14529,N_14938);
nor U15710 (N_15710,N_14788,N_14506);
nand U15711 (N_15711,N_15012,N_15051);
nor U15712 (N_15712,N_14913,N_14876);
nand U15713 (N_15713,N_14412,N_15169);
and U15714 (N_15714,N_15061,N_15016);
or U15715 (N_15715,N_15129,N_14705);
nand U15716 (N_15716,N_15058,N_14468);
and U15717 (N_15717,N_14732,N_14783);
or U15718 (N_15718,N_14577,N_14609);
nand U15719 (N_15719,N_14728,N_14718);
and U15720 (N_15720,N_14607,N_14499);
xnor U15721 (N_15721,N_14994,N_14483);
xor U15722 (N_15722,N_14974,N_14955);
nand U15723 (N_15723,N_14787,N_15020);
or U15724 (N_15724,N_14916,N_15131);
nor U15725 (N_15725,N_14694,N_15138);
or U15726 (N_15726,N_15165,N_14433);
and U15727 (N_15727,N_14746,N_14804);
nand U15728 (N_15728,N_15039,N_14418);
xnor U15729 (N_15729,N_15139,N_15100);
nor U15730 (N_15730,N_15101,N_14769);
or U15731 (N_15731,N_14685,N_14872);
or U15732 (N_15732,N_14790,N_14759);
nand U15733 (N_15733,N_14764,N_14759);
or U15734 (N_15734,N_14401,N_14472);
xnor U15735 (N_15735,N_15070,N_15111);
and U15736 (N_15736,N_14542,N_14403);
and U15737 (N_15737,N_14513,N_14982);
nor U15738 (N_15738,N_14830,N_15155);
xor U15739 (N_15739,N_14799,N_14730);
and U15740 (N_15740,N_15114,N_14808);
nor U15741 (N_15741,N_14670,N_14646);
nand U15742 (N_15742,N_14471,N_15184);
xnor U15743 (N_15743,N_14711,N_15166);
nand U15744 (N_15744,N_14441,N_14576);
and U15745 (N_15745,N_14772,N_14673);
and U15746 (N_15746,N_14849,N_15086);
nor U15747 (N_15747,N_14556,N_14942);
nand U15748 (N_15748,N_14587,N_14846);
nand U15749 (N_15749,N_15109,N_14408);
xnor U15750 (N_15750,N_14986,N_14718);
nand U15751 (N_15751,N_14441,N_14743);
nor U15752 (N_15752,N_15026,N_14613);
nor U15753 (N_15753,N_14879,N_14454);
nor U15754 (N_15754,N_14615,N_14742);
or U15755 (N_15755,N_14509,N_15138);
or U15756 (N_15756,N_14509,N_14617);
nand U15757 (N_15757,N_14772,N_14835);
or U15758 (N_15758,N_14889,N_14820);
and U15759 (N_15759,N_15195,N_14493);
nand U15760 (N_15760,N_15086,N_14466);
xor U15761 (N_15761,N_15136,N_14410);
xnor U15762 (N_15762,N_14719,N_15198);
and U15763 (N_15763,N_14440,N_14505);
xnor U15764 (N_15764,N_14473,N_14426);
or U15765 (N_15765,N_14953,N_14768);
or U15766 (N_15766,N_14643,N_15184);
and U15767 (N_15767,N_15130,N_14612);
nor U15768 (N_15768,N_14874,N_14842);
nor U15769 (N_15769,N_14904,N_14725);
nand U15770 (N_15770,N_15037,N_15072);
xnor U15771 (N_15771,N_15001,N_15090);
nor U15772 (N_15772,N_15135,N_15027);
and U15773 (N_15773,N_14959,N_14516);
and U15774 (N_15774,N_14811,N_15052);
nand U15775 (N_15775,N_14700,N_14602);
xor U15776 (N_15776,N_14438,N_14874);
nand U15777 (N_15777,N_14613,N_14664);
or U15778 (N_15778,N_14414,N_15169);
nor U15779 (N_15779,N_14713,N_14458);
xor U15780 (N_15780,N_15088,N_14952);
and U15781 (N_15781,N_15057,N_15174);
xnor U15782 (N_15782,N_14969,N_15063);
or U15783 (N_15783,N_15044,N_14408);
and U15784 (N_15784,N_14808,N_15068);
and U15785 (N_15785,N_14714,N_14956);
and U15786 (N_15786,N_15174,N_14876);
nor U15787 (N_15787,N_15194,N_15006);
or U15788 (N_15788,N_14725,N_14799);
and U15789 (N_15789,N_15087,N_14754);
or U15790 (N_15790,N_14837,N_14562);
xnor U15791 (N_15791,N_14922,N_14463);
nor U15792 (N_15792,N_14868,N_14451);
nor U15793 (N_15793,N_14588,N_14713);
nor U15794 (N_15794,N_14869,N_15135);
and U15795 (N_15795,N_14498,N_14862);
or U15796 (N_15796,N_14904,N_14824);
xor U15797 (N_15797,N_14764,N_14615);
xnor U15798 (N_15798,N_14943,N_14875);
nand U15799 (N_15799,N_15063,N_14753);
and U15800 (N_15800,N_14985,N_14756);
nor U15801 (N_15801,N_14670,N_14417);
nand U15802 (N_15802,N_15142,N_14474);
xnor U15803 (N_15803,N_15188,N_14991);
nor U15804 (N_15804,N_14478,N_14402);
nor U15805 (N_15805,N_14949,N_14419);
and U15806 (N_15806,N_14418,N_14556);
nor U15807 (N_15807,N_14413,N_14517);
nand U15808 (N_15808,N_15174,N_14824);
xnor U15809 (N_15809,N_14565,N_14811);
nor U15810 (N_15810,N_15171,N_14860);
or U15811 (N_15811,N_14431,N_14677);
nand U15812 (N_15812,N_14519,N_15167);
xnor U15813 (N_15813,N_14588,N_14949);
nor U15814 (N_15814,N_15012,N_14442);
and U15815 (N_15815,N_14816,N_14857);
nor U15816 (N_15816,N_15120,N_14876);
xnor U15817 (N_15817,N_14625,N_14672);
xor U15818 (N_15818,N_14538,N_15097);
xor U15819 (N_15819,N_15166,N_14655);
and U15820 (N_15820,N_14437,N_14539);
nor U15821 (N_15821,N_14440,N_14460);
or U15822 (N_15822,N_14832,N_15149);
xnor U15823 (N_15823,N_15097,N_14557);
or U15824 (N_15824,N_15069,N_14695);
nor U15825 (N_15825,N_14428,N_14660);
or U15826 (N_15826,N_14896,N_14921);
nand U15827 (N_15827,N_15041,N_14518);
nand U15828 (N_15828,N_15165,N_15109);
and U15829 (N_15829,N_15001,N_14506);
nor U15830 (N_15830,N_14720,N_15112);
nor U15831 (N_15831,N_15003,N_14775);
xor U15832 (N_15832,N_14433,N_14626);
xor U15833 (N_15833,N_14485,N_15188);
xnor U15834 (N_15834,N_15140,N_14904);
xor U15835 (N_15835,N_14460,N_15143);
xnor U15836 (N_15836,N_14987,N_15015);
or U15837 (N_15837,N_14519,N_14941);
nor U15838 (N_15838,N_15092,N_14565);
xor U15839 (N_15839,N_14895,N_14932);
xor U15840 (N_15840,N_14518,N_14943);
nor U15841 (N_15841,N_15011,N_14958);
nor U15842 (N_15842,N_14881,N_15048);
xor U15843 (N_15843,N_14419,N_14814);
nand U15844 (N_15844,N_14822,N_14808);
xor U15845 (N_15845,N_14429,N_14901);
and U15846 (N_15846,N_15033,N_14669);
xor U15847 (N_15847,N_15115,N_14608);
xnor U15848 (N_15848,N_14985,N_15062);
and U15849 (N_15849,N_14462,N_14526);
and U15850 (N_15850,N_14859,N_14497);
nand U15851 (N_15851,N_14609,N_14683);
xnor U15852 (N_15852,N_14666,N_14612);
nand U15853 (N_15853,N_14925,N_14947);
nand U15854 (N_15854,N_14445,N_14418);
and U15855 (N_15855,N_14836,N_14935);
nand U15856 (N_15856,N_14824,N_14617);
xor U15857 (N_15857,N_14684,N_15099);
and U15858 (N_15858,N_14930,N_15013);
and U15859 (N_15859,N_14532,N_14631);
nor U15860 (N_15860,N_14480,N_14776);
and U15861 (N_15861,N_15111,N_14771);
nand U15862 (N_15862,N_14976,N_14404);
xor U15863 (N_15863,N_15008,N_14631);
nor U15864 (N_15864,N_15166,N_14654);
and U15865 (N_15865,N_14402,N_14483);
nor U15866 (N_15866,N_14476,N_15021);
xor U15867 (N_15867,N_14535,N_14823);
nand U15868 (N_15868,N_14854,N_14921);
or U15869 (N_15869,N_15134,N_14989);
xor U15870 (N_15870,N_14618,N_14652);
nor U15871 (N_15871,N_14452,N_14546);
and U15872 (N_15872,N_15129,N_14618);
nor U15873 (N_15873,N_14877,N_14636);
xor U15874 (N_15874,N_14578,N_14610);
and U15875 (N_15875,N_14907,N_14531);
and U15876 (N_15876,N_14803,N_14417);
nor U15877 (N_15877,N_14420,N_15035);
and U15878 (N_15878,N_14860,N_14832);
nand U15879 (N_15879,N_14493,N_15028);
and U15880 (N_15880,N_14841,N_14679);
xor U15881 (N_15881,N_14618,N_15135);
xor U15882 (N_15882,N_14602,N_15144);
or U15883 (N_15883,N_15084,N_14490);
or U15884 (N_15884,N_14532,N_14943);
nand U15885 (N_15885,N_15019,N_14422);
nand U15886 (N_15886,N_15023,N_14875);
or U15887 (N_15887,N_14656,N_14924);
xor U15888 (N_15888,N_14555,N_14409);
xor U15889 (N_15889,N_14447,N_14743);
and U15890 (N_15890,N_14505,N_14954);
nand U15891 (N_15891,N_15034,N_14828);
nor U15892 (N_15892,N_14848,N_14578);
nor U15893 (N_15893,N_15060,N_14450);
xnor U15894 (N_15894,N_14761,N_15066);
or U15895 (N_15895,N_14517,N_14685);
and U15896 (N_15896,N_15096,N_15182);
xor U15897 (N_15897,N_15059,N_14846);
nor U15898 (N_15898,N_14903,N_15099);
nand U15899 (N_15899,N_14497,N_15085);
xnor U15900 (N_15900,N_14446,N_15064);
nand U15901 (N_15901,N_14614,N_14654);
nand U15902 (N_15902,N_14778,N_14836);
nor U15903 (N_15903,N_15089,N_14672);
nand U15904 (N_15904,N_14558,N_15181);
and U15905 (N_15905,N_14949,N_14491);
nand U15906 (N_15906,N_14639,N_14585);
xor U15907 (N_15907,N_15005,N_14729);
nor U15908 (N_15908,N_15150,N_14878);
xnor U15909 (N_15909,N_14964,N_14895);
and U15910 (N_15910,N_15053,N_15091);
xnor U15911 (N_15911,N_14688,N_14656);
nand U15912 (N_15912,N_14577,N_15136);
or U15913 (N_15913,N_14492,N_14669);
nand U15914 (N_15914,N_14498,N_14556);
nor U15915 (N_15915,N_14690,N_14729);
nor U15916 (N_15916,N_14942,N_14862);
nand U15917 (N_15917,N_14955,N_14402);
nor U15918 (N_15918,N_14630,N_14550);
nand U15919 (N_15919,N_15078,N_15189);
nor U15920 (N_15920,N_15099,N_14763);
nand U15921 (N_15921,N_14760,N_14434);
or U15922 (N_15922,N_14461,N_14876);
nor U15923 (N_15923,N_15132,N_15164);
and U15924 (N_15924,N_14716,N_15168);
or U15925 (N_15925,N_14490,N_15139);
nand U15926 (N_15926,N_14805,N_14699);
and U15927 (N_15927,N_15025,N_14646);
nand U15928 (N_15928,N_15004,N_15186);
nand U15929 (N_15929,N_14519,N_14505);
xor U15930 (N_15930,N_15185,N_15093);
nand U15931 (N_15931,N_14667,N_14803);
and U15932 (N_15932,N_14801,N_14736);
xor U15933 (N_15933,N_14606,N_14922);
nor U15934 (N_15934,N_14565,N_14516);
nor U15935 (N_15935,N_14993,N_14568);
nand U15936 (N_15936,N_14450,N_14848);
or U15937 (N_15937,N_15121,N_14732);
nor U15938 (N_15938,N_14672,N_14712);
nor U15939 (N_15939,N_14615,N_15143);
nand U15940 (N_15940,N_15096,N_14828);
xor U15941 (N_15941,N_15113,N_15086);
and U15942 (N_15942,N_14411,N_15002);
or U15943 (N_15943,N_15152,N_15078);
and U15944 (N_15944,N_14545,N_15111);
xnor U15945 (N_15945,N_15192,N_14565);
nand U15946 (N_15946,N_14885,N_14790);
nand U15947 (N_15947,N_14446,N_14463);
nor U15948 (N_15948,N_15064,N_14499);
nand U15949 (N_15949,N_14715,N_14429);
nor U15950 (N_15950,N_14991,N_14490);
nand U15951 (N_15951,N_14457,N_14453);
or U15952 (N_15952,N_14653,N_14496);
or U15953 (N_15953,N_14459,N_14781);
nand U15954 (N_15954,N_14841,N_14528);
nand U15955 (N_15955,N_14584,N_14728);
and U15956 (N_15956,N_15062,N_15099);
nor U15957 (N_15957,N_14765,N_15080);
and U15958 (N_15958,N_14475,N_14755);
nand U15959 (N_15959,N_14834,N_14599);
and U15960 (N_15960,N_14603,N_14629);
and U15961 (N_15961,N_14484,N_14772);
and U15962 (N_15962,N_14618,N_15062);
or U15963 (N_15963,N_14889,N_14586);
nand U15964 (N_15964,N_14453,N_15168);
nor U15965 (N_15965,N_15109,N_15085);
nor U15966 (N_15966,N_15001,N_14769);
nand U15967 (N_15967,N_14497,N_14940);
nand U15968 (N_15968,N_14862,N_15125);
or U15969 (N_15969,N_14427,N_14825);
and U15970 (N_15970,N_14628,N_14644);
nor U15971 (N_15971,N_14556,N_14516);
nand U15972 (N_15972,N_14639,N_14859);
or U15973 (N_15973,N_15040,N_15084);
and U15974 (N_15974,N_14562,N_15118);
and U15975 (N_15975,N_14867,N_14820);
and U15976 (N_15976,N_14984,N_14521);
nand U15977 (N_15977,N_14600,N_14438);
xnor U15978 (N_15978,N_14763,N_14591);
nor U15979 (N_15979,N_14884,N_14885);
or U15980 (N_15980,N_15077,N_14828);
xnor U15981 (N_15981,N_14919,N_14725);
and U15982 (N_15982,N_14679,N_14603);
xnor U15983 (N_15983,N_15176,N_14600);
and U15984 (N_15984,N_14927,N_14512);
xor U15985 (N_15985,N_15141,N_14484);
nand U15986 (N_15986,N_15081,N_14458);
nor U15987 (N_15987,N_15172,N_14674);
nand U15988 (N_15988,N_14464,N_15001);
xnor U15989 (N_15989,N_14444,N_14674);
or U15990 (N_15990,N_14980,N_14701);
xnor U15991 (N_15991,N_14885,N_14697);
and U15992 (N_15992,N_14429,N_14527);
nand U15993 (N_15993,N_14477,N_15061);
nand U15994 (N_15994,N_14400,N_15068);
and U15995 (N_15995,N_14781,N_14772);
nand U15996 (N_15996,N_15135,N_14610);
nor U15997 (N_15997,N_14732,N_14621);
nand U15998 (N_15998,N_15181,N_14862);
xnor U15999 (N_15999,N_14899,N_14914);
nor U16000 (N_16000,N_15424,N_15514);
nand U16001 (N_16001,N_15441,N_15554);
nand U16002 (N_16002,N_15314,N_15332);
nor U16003 (N_16003,N_15216,N_15523);
nand U16004 (N_16004,N_15460,N_15617);
nor U16005 (N_16005,N_15716,N_15833);
and U16006 (N_16006,N_15267,N_15822);
and U16007 (N_16007,N_15603,N_15682);
nand U16008 (N_16008,N_15852,N_15732);
xnor U16009 (N_16009,N_15551,N_15610);
and U16010 (N_16010,N_15395,N_15359);
nand U16011 (N_16011,N_15507,N_15742);
xnor U16012 (N_16012,N_15647,N_15672);
xor U16013 (N_16013,N_15527,N_15317);
nand U16014 (N_16014,N_15336,N_15687);
nor U16015 (N_16015,N_15780,N_15338);
nor U16016 (N_16016,N_15434,N_15204);
nand U16017 (N_16017,N_15401,N_15646);
nor U16018 (N_16018,N_15391,N_15686);
nand U16019 (N_16019,N_15818,N_15711);
xor U16020 (N_16020,N_15693,N_15995);
and U16021 (N_16021,N_15209,N_15276);
and U16022 (N_16022,N_15524,N_15817);
nand U16023 (N_16023,N_15779,N_15439);
xnor U16024 (N_16024,N_15989,N_15713);
and U16025 (N_16025,N_15973,N_15270);
nor U16026 (N_16026,N_15960,N_15924);
and U16027 (N_16027,N_15616,N_15600);
nor U16028 (N_16028,N_15367,N_15839);
and U16029 (N_16029,N_15774,N_15325);
or U16030 (N_16030,N_15504,N_15476);
nand U16031 (N_16031,N_15882,N_15720);
nor U16032 (N_16032,N_15393,N_15668);
nor U16033 (N_16033,N_15411,N_15951);
nand U16034 (N_16034,N_15457,N_15928);
nand U16035 (N_16035,N_15806,N_15225);
nand U16036 (N_16036,N_15629,N_15784);
and U16037 (N_16037,N_15837,N_15258);
xor U16038 (N_16038,N_15447,N_15654);
and U16039 (N_16039,N_15811,N_15416);
nand U16040 (N_16040,N_15362,N_15678);
and U16041 (N_16041,N_15714,N_15268);
xor U16042 (N_16042,N_15203,N_15509);
or U16043 (N_16043,N_15583,N_15351);
nand U16044 (N_16044,N_15581,N_15635);
nand U16045 (N_16045,N_15517,N_15501);
and U16046 (N_16046,N_15880,N_15612);
nand U16047 (N_16047,N_15883,N_15731);
or U16048 (N_16048,N_15214,N_15915);
or U16049 (N_16049,N_15316,N_15881);
or U16050 (N_16050,N_15488,N_15718);
or U16051 (N_16051,N_15508,N_15838);
xnor U16052 (N_16052,N_15243,N_15418);
nand U16053 (N_16053,N_15993,N_15749);
nand U16054 (N_16054,N_15226,N_15237);
and U16055 (N_16055,N_15927,N_15277);
nand U16056 (N_16056,N_15631,N_15894);
xnor U16057 (N_16057,N_15475,N_15233);
nor U16058 (N_16058,N_15566,N_15285);
xnor U16059 (N_16059,N_15405,N_15260);
or U16060 (N_16060,N_15483,N_15620);
nor U16061 (N_16061,N_15354,N_15502);
or U16062 (N_16062,N_15522,N_15433);
and U16063 (N_16063,N_15322,N_15804);
or U16064 (N_16064,N_15375,N_15933);
xor U16065 (N_16065,N_15823,N_15762);
nand U16066 (N_16066,N_15584,N_15492);
xnor U16067 (N_16067,N_15201,N_15529);
or U16068 (N_16068,N_15294,N_15248);
or U16069 (N_16069,N_15795,N_15482);
or U16070 (N_16070,N_15572,N_15750);
or U16071 (N_16071,N_15900,N_15472);
or U16072 (N_16072,N_15931,N_15790);
and U16073 (N_16073,N_15957,N_15704);
and U16074 (N_16074,N_15884,N_15499);
nand U16075 (N_16075,N_15988,N_15318);
xnor U16076 (N_16076,N_15675,N_15444);
or U16077 (N_16077,N_15985,N_15305);
nand U16078 (N_16078,N_15613,N_15343);
nor U16079 (N_16079,N_15295,N_15885);
xor U16080 (N_16080,N_15478,N_15220);
nand U16081 (N_16081,N_15281,N_15679);
and U16082 (N_16082,N_15311,N_15320);
xnor U16083 (N_16083,N_15841,N_15601);
and U16084 (N_16084,N_15717,N_15752);
nand U16085 (N_16085,N_15813,N_15775);
xor U16086 (N_16086,N_15531,N_15453);
nand U16087 (N_16087,N_15681,N_15490);
or U16088 (N_16088,N_15596,N_15550);
or U16089 (N_16089,N_15563,N_15286);
xnor U16090 (N_16090,N_15432,N_15794);
or U16091 (N_16091,N_15990,N_15280);
xor U16092 (N_16092,N_15473,N_15764);
or U16093 (N_16093,N_15385,N_15471);
or U16094 (N_16094,N_15796,N_15575);
and U16095 (N_16095,N_15648,N_15339);
and U16096 (N_16096,N_15803,N_15602);
or U16097 (N_16097,N_15234,N_15710);
nor U16098 (N_16098,N_15854,N_15886);
and U16099 (N_16099,N_15866,N_15878);
and U16100 (N_16100,N_15673,N_15573);
nand U16101 (N_16101,N_15862,N_15458);
xnor U16102 (N_16102,N_15505,N_15525);
xnor U16103 (N_16103,N_15848,N_15558);
nor U16104 (N_16104,N_15728,N_15218);
nand U16105 (N_16105,N_15403,N_15279);
xnor U16106 (N_16106,N_15419,N_15217);
and U16107 (N_16107,N_15656,N_15970);
xor U16108 (N_16108,N_15491,N_15944);
nand U16109 (N_16109,N_15628,N_15435);
xnor U16110 (N_16110,N_15956,N_15980);
nor U16111 (N_16111,N_15816,N_15879);
nand U16112 (N_16112,N_15992,N_15388);
nand U16113 (N_16113,N_15858,N_15589);
and U16114 (N_16114,N_15569,N_15567);
or U16115 (N_16115,N_15913,N_15776);
and U16116 (N_16116,N_15251,N_15983);
and U16117 (N_16117,N_15863,N_15291);
xnor U16118 (N_16118,N_15534,N_15238);
nor U16119 (N_16119,N_15308,N_15560);
and U16120 (N_16120,N_15977,N_15827);
nand U16121 (N_16121,N_15363,N_15850);
nor U16122 (N_16122,N_15208,N_15239);
or U16123 (N_16123,N_15431,N_15366);
and U16124 (N_16124,N_15451,N_15495);
nand U16125 (N_16125,N_15422,N_15799);
xnor U16126 (N_16126,N_15530,N_15369);
or U16127 (N_16127,N_15765,N_15709);
nor U16128 (N_16128,N_15864,N_15987);
nand U16129 (N_16129,N_15831,N_15228);
xnor U16130 (N_16130,N_15415,N_15727);
xnor U16131 (N_16131,N_15734,N_15443);
xnor U16132 (N_16132,N_15872,N_15740);
nand U16133 (N_16133,N_15936,N_15333);
and U16134 (N_16134,N_15556,N_15702);
nand U16135 (N_16135,N_15737,N_15697);
and U16136 (N_16136,N_15334,N_15296);
and U16137 (N_16137,N_15290,N_15917);
nor U16138 (N_16138,N_15386,N_15341);
nor U16139 (N_16139,N_15300,N_15412);
or U16140 (N_16140,N_15748,N_15708);
xor U16141 (N_16141,N_15907,N_15825);
or U16142 (N_16142,N_15874,N_15743);
or U16143 (N_16143,N_15259,N_15969);
or U16144 (N_16144,N_15759,N_15684);
and U16145 (N_16145,N_15979,N_15414);
xor U16146 (N_16146,N_15851,N_15479);
and U16147 (N_16147,N_15515,N_15398);
xor U16148 (N_16148,N_15946,N_15725);
nand U16149 (N_16149,N_15899,N_15356);
or U16150 (N_16150,N_15500,N_15565);
or U16151 (N_16151,N_15543,N_15426);
xor U16152 (N_16152,N_15221,N_15814);
nand U16153 (N_16153,N_15691,N_15767);
nor U16154 (N_16154,N_15521,N_15658);
xor U16155 (N_16155,N_15723,N_15562);
xnor U16156 (N_16156,N_15440,N_15446);
and U16157 (N_16157,N_15622,N_15206);
or U16158 (N_16158,N_15739,N_15898);
or U16159 (N_16159,N_15568,N_15901);
and U16160 (N_16160,N_15891,N_15706);
or U16161 (N_16161,N_15820,N_15834);
nor U16162 (N_16162,N_15427,N_15452);
and U16163 (N_16163,N_15760,N_15381);
nand U16164 (N_16164,N_15511,N_15288);
xnor U16165 (N_16165,N_15981,N_15489);
nand U16166 (N_16166,N_15746,N_15921);
or U16167 (N_16167,N_15906,N_15344);
xnor U16168 (N_16168,N_15758,N_15669);
xnor U16169 (N_16169,N_15402,N_15496);
nand U16170 (N_16170,N_15284,N_15413);
or U16171 (N_16171,N_15417,N_15470);
or U16172 (N_16172,N_15655,N_15577);
xnor U16173 (N_16173,N_15802,N_15809);
xor U16174 (N_16174,N_15399,N_15370);
xor U16175 (N_16175,N_15379,N_15662);
xnor U16176 (N_16176,N_15663,N_15867);
xor U16177 (N_16177,N_15461,N_15497);
nor U16178 (N_16178,N_15494,N_15657);
xor U16179 (N_16179,N_15778,N_15950);
xnor U16180 (N_16180,N_15598,N_15212);
or U16181 (N_16181,N_15735,N_15348);
nand U16182 (N_16182,N_15408,N_15614);
xor U16183 (N_16183,N_15597,N_15254);
xnor U16184 (N_16184,N_15604,N_15798);
xnor U16185 (N_16185,N_15219,N_15557);
and U16186 (N_16186,N_15637,N_15309);
xor U16187 (N_16187,N_15892,N_15832);
xnor U16188 (N_16188,N_15861,N_15469);
and U16189 (N_16189,N_15605,N_15241);
nand U16190 (N_16190,N_15474,N_15783);
or U16191 (N_16191,N_15207,N_15539);
xor U16192 (N_16192,N_15346,N_15299);
and U16193 (N_16193,N_15485,N_15893);
nor U16194 (N_16194,N_15707,N_15321);
nand U16195 (N_16195,N_15213,N_15671);
nand U16196 (N_16196,N_15585,N_15922);
xnor U16197 (N_16197,N_15896,N_15694);
or U16198 (N_16198,N_15968,N_15700);
nand U16199 (N_16199,N_15283,N_15755);
nand U16200 (N_16200,N_15683,N_15215);
nand U16201 (N_16201,N_15741,N_15559);
xnor U16202 (N_16202,N_15302,N_15571);
or U16203 (N_16203,N_15676,N_15293);
and U16204 (N_16204,N_15397,N_15463);
xnor U16205 (N_16205,N_15910,N_15312);
xnor U16206 (N_16206,N_15916,N_15540);
and U16207 (N_16207,N_15394,N_15786);
nand U16208 (N_16208,N_15210,N_15624);
or U16209 (N_16209,N_15670,N_15340);
nor U16210 (N_16210,N_15769,N_15705);
nand U16211 (N_16211,N_15926,N_15365);
xnor U16212 (N_16212,N_15952,N_15480);
nand U16213 (N_16213,N_15653,N_15660);
xnor U16214 (N_16214,N_15730,N_15615);
nor U16215 (N_16215,N_15904,N_15692);
or U16216 (N_16216,N_15328,N_15448);
nor U16217 (N_16217,N_15756,N_15587);
or U16218 (N_16218,N_15590,N_15919);
or U16219 (N_16219,N_15244,N_15249);
xnor U16220 (N_16220,N_15287,N_15227);
or U16221 (N_16221,N_15357,N_15954);
nor U16222 (N_16222,N_15247,N_15819);
and U16223 (N_16223,N_15877,N_15680);
nand U16224 (N_16224,N_15326,N_15580);
or U16225 (N_16225,N_15961,N_15410);
or U16226 (N_16226,N_15908,N_15352);
or U16227 (N_16227,N_15998,N_15666);
and U16228 (N_16228,N_15271,N_15939);
and U16229 (N_16229,N_15930,N_15406);
nand U16230 (N_16230,N_15689,N_15310);
and U16231 (N_16231,N_15947,N_15840);
xor U16232 (N_16232,N_15766,N_15736);
xor U16233 (N_16233,N_15532,N_15611);
nand U16234 (N_16234,N_15235,N_15262);
and U16235 (N_16235,N_15315,N_15856);
and U16236 (N_16236,N_15526,N_15889);
and U16237 (N_16237,N_15763,N_15329);
nor U16238 (N_16238,N_15518,N_15396);
xor U16239 (N_16239,N_15782,N_15645);
nor U16240 (N_16240,N_15223,N_15703);
or U16241 (N_16241,N_15425,N_15205);
nand U16242 (N_16242,N_15800,N_15230);
nor U16243 (N_16243,N_15619,N_15246);
nand U16244 (N_16244,N_15757,N_15327);
nand U16245 (N_16245,N_15273,N_15593);
and U16246 (N_16246,N_15875,N_15630);
and U16247 (N_16247,N_15943,N_15791);
xor U16248 (N_16248,N_15506,N_15378);
or U16249 (N_16249,N_15701,N_15512);
nor U16250 (N_16250,N_15516,N_15888);
or U16251 (N_16251,N_15510,N_15436);
xnor U16252 (N_16252,N_15224,N_15963);
nand U16253 (N_16253,N_15430,N_15665);
or U16254 (N_16254,N_15618,N_15229);
nor U16255 (N_16255,N_15345,N_15382);
and U16256 (N_16256,N_15785,N_15659);
or U16257 (N_16257,N_15905,N_15652);
and U16258 (N_16258,N_15971,N_15719);
nand U16259 (N_16259,N_15842,N_15738);
or U16260 (N_16260,N_15984,N_15297);
nand U16261 (N_16261,N_15942,N_15633);
and U16262 (N_16262,N_15955,N_15726);
xnor U16263 (N_16263,N_15211,N_15450);
nand U16264 (N_16264,N_15781,N_15642);
nand U16265 (N_16265,N_15876,N_15869);
and U16266 (N_16266,N_15753,N_15384);
nor U16267 (N_16267,N_15976,N_15627);
or U16268 (N_16268,N_15812,N_15555);
nor U16269 (N_16269,N_15400,N_15256);
nor U16270 (N_16270,N_15996,N_15360);
xor U16271 (N_16271,N_15549,N_15390);
or U16272 (N_16272,N_15389,N_15644);
xor U16273 (N_16273,N_15787,N_15528);
nor U16274 (N_16274,N_15634,N_15751);
or U16275 (N_16275,N_15978,N_15538);
xnor U16276 (N_16276,N_15591,N_15263);
nand U16277 (N_16277,N_15324,N_15421);
and U16278 (N_16278,N_15552,N_15773);
and U16279 (N_16279,N_15909,N_15487);
or U16280 (N_16280,N_15242,N_15253);
or U16281 (N_16281,N_15771,N_15661);
nand U16282 (N_16282,N_15912,N_15292);
xor U16283 (N_16283,N_15377,N_15744);
or U16284 (N_16284,N_15865,N_15965);
xor U16285 (N_16285,N_15306,N_15940);
nand U16286 (N_16286,N_15546,N_15690);
xnor U16287 (N_16287,N_15964,N_15592);
nand U16288 (N_16288,N_15307,N_15349);
nand U16289 (N_16289,N_15625,N_15846);
nor U16290 (N_16290,N_15793,N_15313);
or U16291 (N_16291,N_15200,N_15994);
xor U16292 (N_16292,N_15859,N_15202);
nor U16293 (N_16293,N_15364,N_15582);
xnor U16294 (N_16294,N_15438,N_15576);
nor U16295 (N_16295,N_15437,N_15853);
nor U16296 (N_16296,N_15456,N_15586);
and U16297 (N_16297,N_15358,N_15807);
or U16298 (N_16298,N_15949,N_15974);
nor U16299 (N_16299,N_15513,N_15935);
and U16300 (N_16300,N_15278,N_15371);
nand U16301 (N_16301,N_15698,N_15636);
nand U16302 (N_16302,N_15932,N_15594);
nand U16303 (N_16303,N_15815,N_15409);
xor U16304 (N_16304,N_15257,N_15423);
nand U16305 (N_16305,N_15464,N_15383);
nor U16306 (N_16306,N_15442,N_15805);
or U16307 (N_16307,N_15467,N_15982);
xnor U16308 (N_16308,N_15975,N_15959);
and U16309 (N_16309,N_15824,N_15967);
xor U16310 (N_16310,N_15772,N_15849);
xor U16311 (N_16311,N_15887,N_15997);
and U16312 (N_16312,N_15588,N_15368);
or U16313 (N_16313,N_15484,N_15564);
nor U16314 (N_16314,N_15897,N_15929);
nand U16315 (N_16315,N_15252,N_15699);
and U16316 (N_16316,N_15948,N_15761);
or U16317 (N_16317,N_15374,N_15330);
or U16318 (N_16318,N_15918,N_15466);
or U16319 (N_16319,N_15685,N_15607);
nor U16320 (N_16320,N_15938,N_15331);
xnor U16321 (N_16321,N_15953,N_15533);
nand U16322 (N_16322,N_15845,N_15266);
nor U16323 (N_16323,N_15455,N_15609);
nand U16324 (N_16324,N_15542,N_15301);
or U16325 (N_16325,N_15724,N_15844);
xnor U16326 (N_16326,N_15621,N_15570);
nand U16327 (N_16327,N_15733,N_15945);
xnor U16328 (N_16328,N_15925,N_15553);
xnor U16329 (N_16329,N_15274,N_15650);
nor U16330 (N_16330,N_15319,N_15372);
nand U16331 (N_16331,N_15232,N_15498);
and U16332 (N_16332,N_15289,N_15747);
xnor U16333 (N_16333,N_15873,N_15355);
and U16334 (N_16334,N_15941,N_15608);
nor U16335 (N_16335,N_15643,N_15688);
nor U16336 (N_16336,N_15595,N_15855);
and U16337 (N_16337,N_15250,N_15407);
and U16338 (N_16338,N_15847,N_15792);
nand U16339 (N_16339,N_15911,N_15579);
or U16340 (N_16340,N_15477,N_15768);
nor U16341 (N_16341,N_15828,N_15275);
xor U16342 (N_16342,N_15826,N_15641);
xnor U16343 (N_16343,N_15677,N_15361);
nor U16344 (N_16344,N_15754,N_15303);
nand U16345 (N_16345,N_15626,N_15420);
xnor U16346 (N_16346,N_15895,N_15265);
xor U16347 (N_16347,N_15871,N_15937);
or U16348 (N_16348,N_15578,N_15870);
or U16349 (N_16349,N_15404,N_15449);
or U16350 (N_16350,N_15547,N_15298);
and U16351 (N_16351,N_15664,N_15712);
and U16352 (N_16352,N_15667,N_15323);
nor U16353 (N_16353,N_15903,N_15914);
or U16354 (N_16354,N_15373,N_15715);
xor U16355 (N_16355,N_15245,N_15337);
nor U16356 (N_16356,N_15860,N_15623);
xor U16357 (N_16357,N_15923,N_15638);
or U16358 (N_16358,N_15272,N_15639);
and U16359 (N_16359,N_15745,N_15468);
or U16360 (N_16360,N_15651,N_15902);
and U16361 (N_16361,N_15574,N_15342);
and U16362 (N_16362,N_15606,N_15541);
nand U16363 (N_16363,N_15729,N_15429);
and U16364 (N_16364,N_15836,N_15770);
and U16365 (N_16365,N_15843,N_15777);
nor U16366 (N_16366,N_15599,N_15958);
or U16367 (N_16367,N_15459,N_15986);
or U16368 (N_16368,N_15353,N_15966);
xnor U16369 (N_16369,N_15544,N_15486);
or U16370 (N_16370,N_15493,N_15821);
nand U16371 (N_16371,N_15535,N_15222);
nor U16372 (N_16372,N_15920,N_15721);
or U16373 (N_16373,N_15810,N_15537);
xor U16374 (N_16374,N_15465,N_15462);
nand U16375 (N_16375,N_15255,N_15545);
and U16376 (N_16376,N_15649,N_15376);
nor U16377 (N_16377,N_15890,N_15261);
nand U16378 (N_16378,N_15835,N_15387);
and U16379 (N_16379,N_15695,N_15304);
and U16380 (N_16380,N_15991,N_15264);
and U16381 (N_16381,N_15829,N_15548);
or U16382 (N_16382,N_15520,N_15350);
nand U16383 (N_16383,N_15445,N_15519);
and U16384 (N_16384,N_15392,N_15962);
xnor U16385 (N_16385,N_15972,N_15428);
and U16386 (N_16386,N_15808,N_15696);
nor U16387 (N_16387,N_15380,N_15561);
nand U16388 (N_16388,N_15722,N_15240);
nor U16389 (N_16389,N_15347,N_15632);
or U16390 (N_16390,N_15830,N_15640);
or U16391 (N_16391,N_15934,N_15789);
or U16392 (N_16392,N_15536,N_15857);
nor U16393 (N_16393,N_15999,N_15282);
xor U16394 (N_16394,N_15674,N_15454);
nor U16395 (N_16395,N_15801,N_15236);
nor U16396 (N_16396,N_15269,N_15788);
xnor U16397 (N_16397,N_15335,N_15481);
or U16398 (N_16398,N_15503,N_15797);
xnor U16399 (N_16399,N_15868,N_15231);
nand U16400 (N_16400,N_15403,N_15613);
or U16401 (N_16401,N_15231,N_15591);
nor U16402 (N_16402,N_15879,N_15482);
nand U16403 (N_16403,N_15926,N_15262);
nand U16404 (N_16404,N_15334,N_15241);
and U16405 (N_16405,N_15389,N_15922);
nor U16406 (N_16406,N_15449,N_15510);
and U16407 (N_16407,N_15859,N_15933);
or U16408 (N_16408,N_15603,N_15397);
or U16409 (N_16409,N_15815,N_15848);
or U16410 (N_16410,N_15994,N_15209);
nor U16411 (N_16411,N_15447,N_15819);
and U16412 (N_16412,N_15507,N_15209);
nor U16413 (N_16413,N_15473,N_15683);
or U16414 (N_16414,N_15966,N_15677);
nor U16415 (N_16415,N_15305,N_15898);
nor U16416 (N_16416,N_15696,N_15961);
nor U16417 (N_16417,N_15522,N_15367);
xnor U16418 (N_16418,N_15253,N_15348);
and U16419 (N_16419,N_15505,N_15328);
and U16420 (N_16420,N_15642,N_15662);
xnor U16421 (N_16421,N_15502,N_15677);
nand U16422 (N_16422,N_15768,N_15366);
xnor U16423 (N_16423,N_15360,N_15685);
nor U16424 (N_16424,N_15441,N_15299);
xor U16425 (N_16425,N_15918,N_15644);
xor U16426 (N_16426,N_15583,N_15550);
nand U16427 (N_16427,N_15849,N_15921);
nand U16428 (N_16428,N_15797,N_15394);
nor U16429 (N_16429,N_15645,N_15979);
nand U16430 (N_16430,N_15837,N_15944);
nand U16431 (N_16431,N_15858,N_15771);
nand U16432 (N_16432,N_15417,N_15628);
nor U16433 (N_16433,N_15600,N_15258);
and U16434 (N_16434,N_15221,N_15826);
and U16435 (N_16435,N_15464,N_15919);
or U16436 (N_16436,N_15533,N_15902);
xnor U16437 (N_16437,N_15864,N_15511);
nand U16438 (N_16438,N_15242,N_15519);
and U16439 (N_16439,N_15905,N_15958);
xor U16440 (N_16440,N_15519,N_15600);
nand U16441 (N_16441,N_15883,N_15971);
and U16442 (N_16442,N_15788,N_15508);
nand U16443 (N_16443,N_15360,N_15744);
or U16444 (N_16444,N_15981,N_15426);
nor U16445 (N_16445,N_15327,N_15718);
nor U16446 (N_16446,N_15216,N_15372);
or U16447 (N_16447,N_15673,N_15678);
nand U16448 (N_16448,N_15833,N_15445);
or U16449 (N_16449,N_15805,N_15219);
nand U16450 (N_16450,N_15488,N_15971);
nand U16451 (N_16451,N_15713,N_15524);
nand U16452 (N_16452,N_15231,N_15941);
nand U16453 (N_16453,N_15761,N_15247);
or U16454 (N_16454,N_15556,N_15515);
xnor U16455 (N_16455,N_15641,N_15817);
and U16456 (N_16456,N_15960,N_15290);
or U16457 (N_16457,N_15334,N_15832);
and U16458 (N_16458,N_15581,N_15939);
and U16459 (N_16459,N_15999,N_15495);
nor U16460 (N_16460,N_15381,N_15449);
nor U16461 (N_16461,N_15729,N_15724);
xor U16462 (N_16462,N_15866,N_15497);
or U16463 (N_16463,N_15602,N_15428);
xnor U16464 (N_16464,N_15843,N_15549);
or U16465 (N_16465,N_15409,N_15778);
nand U16466 (N_16466,N_15941,N_15852);
nor U16467 (N_16467,N_15817,N_15734);
nand U16468 (N_16468,N_15896,N_15516);
or U16469 (N_16469,N_15687,N_15765);
nand U16470 (N_16470,N_15709,N_15879);
xnor U16471 (N_16471,N_15484,N_15607);
xor U16472 (N_16472,N_15451,N_15456);
nor U16473 (N_16473,N_15949,N_15626);
nand U16474 (N_16474,N_15633,N_15790);
or U16475 (N_16475,N_15760,N_15538);
nand U16476 (N_16476,N_15362,N_15350);
or U16477 (N_16477,N_15690,N_15443);
or U16478 (N_16478,N_15938,N_15460);
or U16479 (N_16479,N_15367,N_15976);
or U16480 (N_16480,N_15457,N_15295);
nor U16481 (N_16481,N_15576,N_15208);
or U16482 (N_16482,N_15835,N_15646);
nor U16483 (N_16483,N_15240,N_15667);
and U16484 (N_16484,N_15998,N_15582);
nand U16485 (N_16485,N_15324,N_15209);
or U16486 (N_16486,N_15531,N_15554);
xnor U16487 (N_16487,N_15234,N_15732);
and U16488 (N_16488,N_15334,N_15371);
nor U16489 (N_16489,N_15798,N_15950);
or U16490 (N_16490,N_15765,N_15862);
or U16491 (N_16491,N_15499,N_15463);
xor U16492 (N_16492,N_15475,N_15634);
and U16493 (N_16493,N_15869,N_15565);
and U16494 (N_16494,N_15716,N_15781);
and U16495 (N_16495,N_15238,N_15596);
nor U16496 (N_16496,N_15998,N_15334);
or U16497 (N_16497,N_15963,N_15425);
nand U16498 (N_16498,N_15337,N_15952);
and U16499 (N_16499,N_15845,N_15543);
nor U16500 (N_16500,N_15939,N_15396);
and U16501 (N_16501,N_15777,N_15607);
xnor U16502 (N_16502,N_15720,N_15750);
and U16503 (N_16503,N_15892,N_15937);
xor U16504 (N_16504,N_15200,N_15795);
or U16505 (N_16505,N_15307,N_15732);
and U16506 (N_16506,N_15326,N_15870);
nand U16507 (N_16507,N_15762,N_15247);
nand U16508 (N_16508,N_15898,N_15921);
or U16509 (N_16509,N_15700,N_15380);
and U16510 (N_16510,N_15843,N_15469);
nor U16511 (N_16511,N_15607,N_15989);
and U16512 (N_16512,N_15917,N_15294);
and U16513 (N_16513,N_15993,N_15495);
nor U16514 (N_16514,N_15669,N_15840);
xnor U16515 (N_16515,N_15906,N_15952);
or U16516 (N_16516,N_15400,N_15697);
or U16517 (N_16517,N_15743,N_15733);
and U16518 (N_16518,N_15743,N_15943);
xnor U16519 (N_16519,N_15298,N_15458);
nand U16520 (N_16520,N_15411,N_15805);
xor U16521 (N_16521,N_15744,N_15875);
or U16522 (N_16522,N_15357,N_15811);
or U16523 (N_16523,N_15427,N_15967);
and U16524 (N_16524,N_15821,N_15806);
nor U16525 (N_16525,N_15416,N_15699);
nand U16526 (N_16526,N_15516,N_15937);
nor U16527 (N_16527,N_15959,N_15932);
xor U16528 (N_16528,N_15652,N_15215);
or U16529 (N_16529,N_15602,N_15407);
or U16530 (N_16530,N_15699,N_15217);
nor U16531 (N_16531,N_15625,N_15663);
and U16532 (N_16532,N_15581,N_15414);
nand U16533 (N_16533,N_15505,N_15419);
xor U16534 (N_16534,N_15247,N_15593);
nand U16535 (N_16535,N_15322,N_15500);
and U16536 (N_16536,N_15239,N_15848);
and U16537 (N_16537,N_15495,N_15276);
nand U16538 (N_16538,N_15679,N_15705);
nand U16539 (N_16539,N_15969,N_15784);
nor U16540 (N_16540,N_15318,N_15446);
xnor U16541 (N_16541,N_15711,N_15328);
nor U16542 (N_16542,N_15964,N_15916);
or U16543 (N_16543,N_15777,N_15237);
nand U16544 (N_16544,N_15410,N_15623);
nor U16545 (N_16545,N_15353,N_15637);
or U16546 (N_16546,N_15911,N_15675);
and U16547 (N_16547,N_15709,N_15297);
or U16548 (N_16548,N_15729,N_15998);
nand U16549 (N_16549,N_15465,N_15327);
and U16550 (N_16550,N_15842,N_15939);
or U16551 (N_16551,N_15614,N_15300);
nand U16552 (N_16552,N_15996,N_15332);
or U16553 (N_16553,N_15525,N_15779);
and U16554 (N_16554,N_15343,N_15361);
nor U16555 (N_16555,N_15674,N_15963);
xnor U16556 (N_16556,N_15384,N_15781);
or U16557 (N_16557,N_15788,N_15332);
and U16558 (N_16558,N_15297,N_15382);
or U16559 (N_16559,N_15973,N_15365);
or U16560 (N_16560,N_15822,N_15845);
xor U16561 (N_16561,N_15899,N_15470);
and U16562 (N_16562,N_15295,N_15786);
or U16563 (N_16563,N_15826,N_15467);
nor U16564 (N_16564,N_15743,N_15979);
nor U16565 (N_16565,N_15384,N_15953);
and U16566 (N_16566,N_15646,N_15611);
nor U16567 (N_16567,N_15992,N_15480);
nor U16568 (N_16568,N_15908,N_15373);
nand U16569 (N_16569,N_15823,N_15491);
or U16570 (N_16570,N_15870,N_15794);
nand U16571 (N_16571,N_15965,N_15892);
xor U16572 (N_16572,N_15513,N_15910);
or U16573 (N_16573,N_15746,N_15893);
or U16574 (N_16574,N_15386,N_15921);
xor U16575 (N_16575,N_15521,N_15412);
and U16576 (N_16576,N_15274,N_15788);
xnor U16577 (N_16577,N_15809,N_15393);
nor U16578 (N_16578,N_15973,N_15751);
nand U16579 (N_16579,N_15620,N_15468);
nor U16580 (N_16580,N_15784,N_15506);
nand U16581 (N_16581,N_15396,N_15770);
or U16582 (N_16582,N_15811,N_15609);
and U16583 (N_16583,N_15693,N_15275);
or U16584 (N_16584,N_15783,N_15516);
or U16585 (N_16585,N_15793,N_15344);
or U16586 (N_16586,N_15706,N_15281);
nor U16587 (N_16587,N_15992,N_15667);
xor U16588 (N_16588,N_15468,N_15456);
nor U16589 (N_16589,N_15860,N_15983);
nand U16590 (N_16590,N_15777,N_15840);
xor U16591 (N_16591,N_15585,N_15582);
and U16592 (N_16592,N_15458,N_15686);
nand U16593 (N_16593,N_15984,N_15951);
or U16594 (N_16594,N_15610,N_15771);
or U16595 (N_16595,N_15813,N_15525);
nand U16596 (N_16596,N_15351,N_15240);
xnor U16597 (N_16597,N_15926,N_15453);
or U16598 (N_16598,N_15241,N_15321);
nor U16599 (N_16599,N_15590,N_15346);
nand U16600 (N_16600,N_15597,N_15995);
and U16601 (N_16601,N_15670,N_15729);
or U16602 (N_16602,N_15563,N_15936);
nor U16603 (N_16603,N_15217,N_15999);
nand U16604 (N_16604,N_15724,N_15424);
and U16605 (N_16605,N_15443,N_15257);
xnor U16606 (N_16606,N_15496,N_15354);
xnor U16607 (N_16607,N_15226,N_15655);
nand U16608 (N_16608,N_15793,N_15752);
or U16609 (N_16609,N_15975,N_15542);
xnor U16610 (N_16610,N_15812,N_15932);
nand U16611 (N_16611,N_15950,N_15678);
xnor U16612 (N_16612,N_15472,N_15740);
and U16613 (N_16613,N_15465,N_15649);
or U16614 (N_16614,N_15347,N_15200);
xnor U16615 (N_16615,N_15778,N_15816);
and U16616 (N_16616,N_15400,N_15662);
xor U16617 (N_16617,N_15580,N_15553);
xnor U16618 (N_16618,N_15528,N_15260);
or U16619 (N_16619,N_15961,N_15750);
nor U16620 (N_16620,N_15670,N_15924);
xnor U16621 (N_16621,N_15729,N_15350);
nor U16622 (N_16622,N_15718,N_15489);
xor U16623 (N_16623,N_15535,N_15859);
and U16624 (N_16624,N_15654,N_15985);
nor U16625 (N_16625,N_15935,N_15780);
and U16626 (N_16626,N_15719,N_15635);
nor U16627 (N_16627,N_15863,N_15664);
or U16628 (N_16628,N_15649,N_15745);
nand U16629 (N_16629,N_15308,N_15730);
or U16630 (N_16630,N_15462,N_15393);
or U16631 (N_16631,N_15339,N_15914);
nand U16632 (N_16632,N_15766,N_15500);
nand U16633 (N_16633,N_15383,N_15735);
xor U16634 (N_16634,N_15361,N_15488);
nor U16635 (N_16635,N_15614,N_15846);
nand U16636 (N_16636,N_15731,N_15838);
xnor U16637 (N_16637,N_15749,N_15459);
or U16638 (N_16638,N_15605,N_15955);
nand U16639 (N_16639,N_15512,N_15640);
and U16640 (N_16640,N_15320,N_15728);
xnor U16641 (N_16641,N_15464,N_15573);
or U16642 (N_16642,N_15431,N_15793);
or U16643 (N_16643,N_15876,N_15628);
and U16644 (N_16644,N_15586,N_15888);
nand U16645 (N_16645,N_15284,N_15685);
xor U16646 (N_16646,N_15431,N_15616);
nand U16647 (N_16647,N_15790,N_15796);
nor U16648 (N_16648,N_15931,N_15642);
xor U16649 (N_16649,N_15268,N_15270);
or U16650 (N_16650,N_15811,N_15817);
xnor U16651 (N_16651,N_15443,N_15673);
nand U16652 (N_16652,N_15290,N_15327);
xnor U16653 (N_16653,N_15500,N_15883);
xor U16654 (N_16654,N_15498,N_15314);
xnor U16655 (N_16655,N_15323,N_15268);
and U16656 (N_16656,N_15600,N_15871);
xor U16657 (N_16657,N_15813,N_15764);
or U16658 (N_16658,N_15753,N_15586);
nor U16659 (N_16659,N_15537,N_15804);
xor U16660 (N_16660,N_15952,N_15806);
xnor U16661 (N_16661,N_15786,N_15807);
nand U16662 (N_16662,N_15583,N_15891);
nand U16663 (N_16663,N_15878,N_15305);
xnor U16664 (N_16664,N_15240,N_15719);
nor U16665 (N_16665,N_15414,N_15537);
nand U16666 (N_16666,N_15640,N_15780);
and U16667 (N_16667,N_15931,N_15316);
nand U16668 (N_16668,N_15250,N_15846);
nand U16669 (N_16669,N_15810,N_15639);
nand U16670 (N_16670,N_15237,N_15966);
or U16671 (N_16671,N_15707,N_15875);
nor U16672 (N_16672,N_15753,N_15648);
nand U16673 (N_16673,N_15478,N_15570);
nand U16674 (N_16674,N_15867,N_15945);
xnor U16675 (N_16675,N_15385,N_15890);
nand U16676 (N_16676,N_15237,N_15643);
nor U16677 (N_16677,N_15843,N_15262);
and U16678 (N_16678,N_15597,N_15464);
or U16679 (N_16679,N_15857,N_15909);
nand U16680 (N_16680,N_15229,N_15763);
xor U16681 (N_16681,N_15906,N_15345);
or U16682 (N_16682,N_15727,N_15873);
and U16683 (N_16683,N_15223,N_15528);
nor U16684 (N_16684,N_15721,N_15454);
nor U16685 (N_16685,N_15358,N_15802);
nor U16686 (N_16686,N_15731,N_15588);
and U16687 (N_16687,N_15947,N_15775);
nand U16688 (N_16688,N_15241,N_15886);
or U16689 (N_16689,N_15686,N_15564);
and U16690 (N_16690,N_15535,N_15340);
xnor U16691 (N_16691,N_15852,N_15337);
nor U16692 (N_16692,N_15358,N_15920);
xnor U16693 (N_16693,N_15551,N_15205);
xnor U16694 (N_16694,N_15787,N_15401);
nor U16695 (N_16695,N_15449,N_15482);
and U16696 (N_16696,N_15367,N_15448);
or U16697 (N_16697,N_15863,N_15544);
xor U16698 (N_16698,N_15628,N_15656);
and U16699 (N_16699,N_15261,N_15741);
and U16700 (N_16700,N_15388,N_15716);
nand U16701 (N_16701,N_15494,N_15478);
and U16702 (N_16702,N_15561,N_15680);
nor U16703 (N_16703,N_15268,N_15526);
nor U16704 (N_16704,N_15836,N_15625);
or U16705 (N_16705,N_15474,N_15904);
nor U16706 (N_16706,N_15306,N_15221);
and U16707 (N_16707,N_15644,N_15600);
nand U16708 (N_16708,N_15304,N_15915);
nor U16709 (N_16709,N_15785,N_15912);
nor U16710 (N_16710,N_15891,N_15795);
nor U16711 (N_16711,N_15210,N_15638);
or U16712 (N_16712,N_15421,N_15653);
xnor U16713 (N_16713,N_15848,N_15889);
and U16714 (N_16714,N_15343,N_15782);
xnor U16715 (N_16715,N_15767,N_15863);
or U16716 (N_16716,N_15792,N_15902);
and U16717 (N_16717,N_15200,N_15860);
or U16718 (N_16718,N_15262,N_15497);
nor U16719 (N_16719,N_15436,N_15450);
xor U16720 (N_16720,N_15571,N_15774);
nor U16721 (N_16721,N_15954,N_15457);
nand U16722 (N_16722,N_15668,N_15553);
nor U16723 (N_16723,N_15409,N_15436);
nand U16724 (N_16724,N_15513,N_15420);
xor U16725 (N_16725,N_15309,N_15267);
nand U16726 (N_16726,N_15561,N_15555);
and U16727 (N_16727,N_15289,N_15766);
and U16728 (N_16728,N_15798,N_15209);
nand U16729 (N_16729,N_15393,N_15439);
and U16730 (N_16730,N_15753,N_15948);
and U16731 (N_16731,N_15340,N_15280);
or U16732 (N_16732,N_15463,N_15707);
nand U16733 (N_16733,N_15275,N_15667);
and U16734 (N_16734,N_15428,N_15670);
nand U16735 (N_16735,N_15815,N_15505);
nand U16736 (N_16736,N_15623,N_15631);
nand U16737 (N_16737,N_15287,N_15740);
and U16738 (N_16738,N_15772,N_15864);
xnor U16739 (N_16739,N_15246,N_15634);
and U16740 (N_16740,N_15244,N_15418);
or U16741 (N_16741,N_15645,N_15475);
or U16742 (N_16742,N_15810,N_15888);
nor U16743 (N_16743,N_15265,N_15405);
xor U16744 (N_16744,N_15999,N_15606);
or U16745 (N_16745,N_15376,N_15608);
and U16746 (N_16746,N_15654,N_15973);
and U16747 (N_16747,N_15936,N_15477);
nand U16748 (N_16748,N_15597,N_15299);
and U16749 (N_16749,N_15567,N_15949);
nand U16750 (N_16750,N_15268,N_15937);
nor U16751 (N_16751,N_15976,N_15241);
or U16752 (N_16752,N_15489,N_15996);
xnor U16753 (N_16753,N_15724,N_15874);
nand U16754 (N_16754,N_15264,N_15700);
nand U16755 (N_16755,N_15352,N_15851);
nor U16756 (N_16756,N_15683,N_15825);
nor U16757 (N_16757,N_15221,N_15768);
and U16758 (N_16758,N_15459,N_15233);
xnor U16759 (N_16759,N_15303,N_15289);
or U16760 (N_16760,N_15462,N_15455);
nand U16761 (N_16761,N_15441,N_15399);
nand U16762 (N_16762,N_15313,N_15753);
xnor U16763 (N_16763,N_15838,N_15719);
or U16764 (N_16764,N_15967,N_15543);
and U16765 (N_16765,N_15684,N_15773);
or U16766 (N_16766,N_15456,N_15552);
nor U16767 (N_16767,N_15816,N_15558);
or U16768 (N_16768,N_15599,N_15329);
xor U16769 (N_16769,N_15861,N_15837);
nand U16770 (N_16770,N_15557,N_15954);
nor U16771 (N_16771,N_15522,N_15722);
xor U16772 (N_16772,N_15218,N_15957);
xnor U16773 (N_16773,N_15437,N_15356);
xor U16774 (N_16774,N_15820,N_15934);
or U16775 (N_16775,N_15698,N_15816);
nand U16776 (N_16776,N_15811,N_15205);
and U16777 (N_16777,N_15703,N_15211);
or U16778 (N_16778,N_15789,N_15741);
xnor U16779 (N_16779,N_15995,N_15250);
xnor U16780 (N_16780,N_15963,N_15240);
or U16781 (N_16781,N_15836,N_15236);
nand U16782 (N_16782,N_15261,N_15884);
or U16783 (N_16783,N_15618,N_15402);
xnor U16784 (N_16784,N_15515,N_15207);
or U16785 (N_16785,N_15855,N_15491);
and U16786 (N_16786,N_15673,N_15754);
or U16787 (N_16787,N_15245,N_15825);
nand U16788 (N_16788,N_15396,N_15334);
nand U16789 (N_16789,N_15496,N_15273);
xor U16790 (N_16790,N_15507,N_15411);
nand U16791 (N_16791,N_15413,N_15633);
or U16792 (N_16792,N_15597,N_15488);
nand U16793 (N_16793,N_15244,N_15679);
and U16794 (N_16794,N_15940,N_15654);
xnor U16795 (N_16795,N_15749,N_15884);
nand U16796 (N_16796,N_15905,N_15428);
or U16797 (N_16797,N_15307,N_15891);
nand U16798 (N_16798,N_15707,N_15856);
and U16799 (N_16799,N_15308,N_15686);
and U16800 (N_16800,N_16223,N_16768);
and U16801 (N_16801,N_16058,N_16230);
xor U16802 (N_16802,N_16427,N_16143);
nand U16803 (N_16803,N_16241,N_16140);
xor U16804 (N_16804,N_16454,N_16262);
and U16805 (N_16805,N_16261,N_16560);
nor U16806 (N_16806,N_16209,N_16554);
and U16807 (N_16807,N_16666,N_16690);
or U16808 (N_16808,N_16721,N_16305);
or U16809 (N_16809,N_16071,N_16180);
xor U16810 (N_16810,N_16777,N_16108);
nand U16811 (N_16811,N_16270,N_16611);
nor U16812 (N_16812,N_16088,N_16333);
or U16813 (N_16813,N_16064,N_16439);
nor U16814 (N_16814,N_16050,N_16582);
and U16815 (N_16815,N_16158,N_16066);
or U16816 (N_16816,N_16102,N_16380);
nand U16817 (N_16817,N_16431,N_16299);
and U16818 (N_16818,N_16092,N_16199);
or U16819 (N_16819,N_16580,N_16406);
xnor U16820 (N_16820,N_16404,N_16649);
xnor U16821 (N_16821,N_16485,N_16292);
nand U16822 (N_16822,N_16515,N_16166);
nor U16823 (N_16823,N_16113,N_16222);
and U16824 (N_16824,N_16687,N_16033);
and U16825 (N_16825,N_16310,N_16403);
nand U16826 (N_16826,N_16449,N_16274);
xnor U16827 (N_16827,N_16095,N_16795);
nand U16828 (N_16828,N_16749,N_16324);
xor U16829 (N_16829,N_16120,N_16481);
nand U16830 (N_16830,N_16225,N_16119);
nand U16831 (N_16831,N_16667,N_16326);
nand U16832 (N_16832,N_16383,N_16765);
nor U16833 (N_16833,N_16148,N_16249);
nand U16834 (N_16834,N_16542,N_16437);
xor U16835 (N_16835,N_16693,N_16503);
and U16836 (N_16836,N_16268,N_16609);
nor U16837 (N_16837,N_16060,N_16643);
xnor U16838 (N_16838,N_16679,N_16364);
and U16839 (N_16839,N_16188,N_16207);
nand U16840 (N_16840,N_16743,N_16189);
and U16841 (N_16841,N_16365,N_16137);
xor U16842 (N_16842,N_16085,N_16239);
and U16843 (N_16843,N_16685,N_16699);
or U16844 (N_16844,N_16297,N_16208);
and U16845 (N_16845,N_16183,N_16116);
nand U16846 (N_16846,N_16564,N_16584);
or U16847 (N_16847,N_16368,N_16078);
nor U16848 (N_16848,N_16349,N_16311);
and U16849 (N_16849,N_16520,N_16316);
nand U16850 (N_16850,N_16613,N_16484);
xnor U16851 (N_16851,N_16659,N_16414);
xnor U16852 (N_16852,N_16125,N_16417);
nand U16853 (N_16853,N_16450,N_16797);
xor U16854 (N_16854,N_16110,N_16791);
nand U16855 (N_16855,N_16312,N_16157);
or U16856 (N_16856,N_16232,N_16196);
or U16857 (N_16857,N_16602,N_16635);
or U16858 (N_16858,N_16793,N_16764);
nand U16859 (N_16859,N_16395,N_16746);
nand U16860 (N_16860,N_16546,N_16354);
and U16861 (N_16861,N_16151,N_16363);
nor U16862 (N_16862,N_16422,N_16592);
and U16863 (N_16863,N_16553,N_16537);
nand U16864 (N_16864,N_16424,N_16769);
and U16865 (N_16865,N_16736,N_16000);
nand U16866 (N_16866,N_16074,N_16195);
and U16867 (N_16867,N_16750,N_16692);
nor U16868 (N_16868,N_16250,N_16547);
xor U16869 (N_16869,N_16455,N_16615);
or U16870 (N_16870,N_16676,N_16341);
or U16871 (N_16871,N_16393,N_16696);
nor U16872 (N_16872,N_16475,N_16339);
nand U16873 (N_16873,N_16723,N_16130);
or U16874 (N_16874,N_16751,N_16012);
and U16875 (N_16875,N_16641,N_16224);
nand U16876 (N_16876,N_16147,N_16030);
and U16877 (N_16877,N_16488,N_16366);
nor U16878 (N_16878,N_16570,N_16680);
and U16879 (N_16879,N_16303,N_16332);
xor U16880 (N_16880,N_16080,N_16522);
nand U16881 (N_16881,N_16718,N_16678);
xnor U16882 (N_16882,N_16251,N_16445);
nand U16883 (N_16883,N_16145,N_16487);
nand U16884 (N_16884,N_16519,N_16565);
nand U16885 (N_16885,N_16356,N_16319);
nor U16886 (N_16886,N_16122,N_16440);
or U16887 (N_16887,N_16501,N_16556);
nor U16888 (N_16888,N_16744,N_16294);
nor U16889 (N_16889,N_16205,N_16523);
and U16890 (N_16890,N_16355,N_16098);
and U16891 (N_16891,N_16174,N_16229);
xor U16892 (N_16892,N_16541,N_16379);
xnor U16893 (N_16893,N_16049,N_16351);
nor U16894 (N_16894,N_16083,N_16630);
and U16895 (N_16895,N_16430,N_16720);
nor U16896 (N_16896,N_16226,N_16682);
nand U16897 (N_16897,N_16260,N_16367);
nor U16898 (N_16898,N_16134,N_16684);
xor U16899 (N_16899,N_16650,N_16664);
or U16900 (N_16900,N_16272,N_16442);
xnor U16901 (N_16901,N_16287,N_16182);
nor U16902 (N_16902,N_16082,N_16127);
or U16903 (N_16903,N_16001,N_16415);
nor U16904 (N_16904,N_16518,N_16533);
or U16905 (N_16905,N_16105,N_16621);
or U16906 (N_16906,N_16253,N_16674);
or U16907 (N_16907,N_16638,N_16628);
nor U16908 (N_16908,N_16357,N_16639);
or U16909 (N_16909,N_16426,N_16799);
and U16910 (N_16910,N_16179,N_16571);
and U16911 (N_16911,N_16123,N_16551);
nand U16912 (N_16912,N_16604,N_16017);
and U16913 (N_16913,N_16173,N_16007);
nor U16914 (N_16914,N_16063,N_16087);
nand U16915 (N_16915,N_16405,N_16606);
nand U16916 (N_16916,N_16474,N_16375);
and U16917 (N_16917,N_16138,N_16315);
nand U16918 (N_16918,N_16771,N_16708);
and U16919 (N_16919,N_16069,N_16091);
nor U16920 (N_16920,N_16322,N_16766);
xnor U16921 (N_16921,N_16651,N_16745);
nand U16922 (N_16922,N_16524,N_16040);
or U16923 (N_16923,N_16727,N_16192);
or U16924 (N_16924,N_16053,N_16348);
nor U16925 (N_16925,N_16478,N_16742);
and U16926 (N_16926,N_16645,N_16489);
nand U16927 (N_16927,N_16735,N_16291);
and U16928 (N_16928,N_16335,N_16644);
and U16929 (N_16929,N_16280,N_16569);
or U16930 (N_16930,N_16656,N_16707);
or U16931 (N_16931,N_16008,N_16117);
and U16932 (N_16932,N_16257,N_16300);
xor U16933 (N_16933,N_16121,N_16394);
nand U16934 (N_16934,N_16586,N_16516);
nand U16935 (N_16935,N_16231,N_16539);
nand U16936 (N_16936,N_16616,N_16675);
nand U16937 (N_16937,N_16374,N_16234);
xor U16938 (N_16938,N_16614,N_16309);
nor U16939 (N_16939,N_16115,N_16730);
xnor U16940 (N_16940,N_16778,N_16217);
or U16941 (N_16941,N_16558,N_16329);
nand U16942 (N_16942,N_16384,N_16468);
nand U16943 (N_16943,N_16411,N_16453);
nand U16944 (N_16944,N_16480,N_16052);
nor U16945 (N_16945,N_16005,N_16323);
or U16946 (N_16946,N_16055,N_16617);
nor U16947 (N_16947,N_16711,N_16794);
xnor U16948 (N_16948,N_16107,N_16267);
or U16949 (N_16949,N_16704,N_16047);
xnor U16950 (N_16950,N_16298,N_16725);
nor U16951 (N_16951,N_16245,N_16197);
nand U16952 (N_16952,N_16677,N_16446);
xnor U16953 (N_16953,N_16510,N_16779);
nor U16954 (N_16954,N_16304,N_16695);
nor U16955 (N_16955,N_16671,N_16263);
and U16956 (N_16956,N_16076,N_16773);
xnor U16957 (N_16957,N_16248,N_16738);
nor U16958 (N_16958,N_16511,N_16663);
xnor U16959 (N_16959,N_16443,N_16529);
xor U16960 (N_16960,N_16737,N_16572);
or U16961 (N_16961,N_16376,N_16447);
nor U16962 (N_16962,N_16763,N_16201);
and U16963 (N_16963,N_16461,N_16798);
or U16964 (N_16964,N_16715,N_16026);
nand U16965 (N_16965,N_16061,N_16096);
or U16966 (N_16966,N_16466,N_16728);
nor U16967 (N_16967,N_16072,N_16184);
xor U16968 (N_16968,N_16203,N_16264);
and U16969 (N_16969,N_16330,N_16200);
and U16970 (N_16970,N_16160,N_16540);
nor U16971 (N_16971,N_16494,N_16101);
nor U16972 (N_16972,N_16528,N_16691);
xnor U16973 (N_16973,N_16290,N_16109);
xnor U16974 (N_16974,N_16390,N_16792);
nand U16975 (N_16975,N_16697,N_16362);
nor U16976 (N_16976,N_16118,N_16787);
nand U16977 (N_16977,N_16521,N_16103);
nand U16978 (N_16978,N_16788,N_16077);
xnor U16979 (N_16979,N_16626,N_16552);
xor U16980 (N_16980,N_16549,N_16607);
nand U16981 (N_16981,N_16086,N_16283);
or U16982 (N_16982,N_16458,N_16227);
xnor U16983 (N_16983,N_16509,N_16465);
nor U16984 (N_16984,N_16590,N_16605);
xor U16985 (N_16985,N_16396,N_16451);
and U16986 (N_16986,N_16497,N_16416);
xnor U16987 (N_16987,N_16579,N_16653);
and U16988 (N_16988,N_16634,N_16289);
xor U16989 (N_16989,N_16716,N_16350);
xnor U16990 (N_16990,N_16618,N_16670);
and U16991 (N_16991,N_16421,N_16486);
or U16992 (N_16992,N_16002,N_16022);
or U16993 (N_16993,N_16345,N_16097);
nor U16994 (N_16994,N_16563,N_16473);
or U16995 (N_16995,N_16006,N_16432);
nand U16996 (N_16996,N_16700,N_16627);
or U16997 (N_16997,N_16555,N_16194);
xnor U16998 (N_16998,N_16504,N_16392);
nand U16999 (N_16999,N_16048,N_16469);
xnor U17000 (N_17000,N_16386,N_16093);
or U17001 (N_17001,N_16610,N_16713);
nand U17002 (N_17002,N_16597,N_16100);
nand U17003 (N_17003,N_16531,N_16202);
nor U17004 (N_17004,N_16023,N_16191);
and U17005 (N_17005,N_16028,N_16419);
or U17006 (N_17006,N_16039,N_16265);
or U17007 (N_17007,N_16652,N_16598);
nand U17008 (N_17008,N_16576,N_16429);
nor U17009 (N_17009,N_16133,N_16544);
and U17010 (N_17010,N_16789,N_16508);
nor U17011 (N_17011,N_16758,N_16709);
xnor U17012 (N_17012,N_16067,N_16428);
nand U17013 (N_17013,N_16400,N_16233);
nor U17014 (N_17014,N_16654,N_16438);
xnor U17015 (N_17015,N_16694,N_16658);
and U17016 (N_17016,N_16075,N_16178);
nand U17017 (N_17017,N_16517,N_16661);
xnor U17018 (N_17018,N_16464,N_16433);
nor U17019 (N_17019,N_16318,N_16276);
or U17020 (N_17020,N_16593,N_16009);
nand U17021 (N_17021,N_16741,N_16284);
and U17022 (N_17022,N_16603,N_16373);
or U17023 (N_17023,N_16084,N_16471);
xor U17024 (N_17024,N_16360,N_16612);
nand U17025 (N_17025,N_16702,N_16514);
xor U17026 (N_17026,N_16279,N_16631);
and U17027 (N_17027,N_16770,N_16470);
xnor U17028 (N_17028,N_16755,N_16689);
nand U17029 (N_17029,N_16046,N_16371);
or U17030 (N_17030,N_16408,N_16600);
xor U17031 (N_17031,N_16124,N_16314);
or U17032 (N_17032,N_16215,N_16623);
or U17033 (N_17033,N_16206,N_16459);
nor U17034 (N_17034,N_16062,N_16035);
or U17035 (N_17035,N_16479,N_16247);
nand U17036 (N_17036,N_16759,N_16218);
or U17037 (N_17037,N_16352,N_16171);
nor U17038 (N_17038,N_16266,N_16167);
nor U17039 (N_17039,N_16477,N_16338);
xor U17040 (N_17040,N_16038,N_16242);
or U17041 (N_17041,N_16633,N_16211);
xor U17042 (N_17042,N_16003,N_16672);
nand U17043 (N_17043,N_16296,N_16244);
xnor U17044 (N_17044,N_16104,N_16307);
and U17045 (N_17045,N_16129,N_16513);
or U17046 (N_17046,N_16594,N_16328);
and U17047 (N_17047,N_16648,N_16657);
and U17048 (N_17048,N_16293,N_16629);
xnor U17049 (N_17049,N_16646,N_16169);
or U17050 (N_17050,N_16387,N_16347);
xor U17051 (N_17051,N_16783,N_16669);
and U17052 (N_17052,N_16302,N_16668);
xnor U17053 (N_17053,N_16340,N_16756);
xnor U17054 (N_17054,N_16595,N_16212);
and U17055 (N_17055,N_16165,N_16334);
or U17056 (N_17056,N_16252,N_16761);
or U17057 (N_17057,N_16505,N_16624);
xnor U17058 (N_17058,N_16220,N_16089);
xor U17059 (N_17059,N_16378,N_16647);
nor U17060 (N_17060,N_16562,N_16295);
and U17061 (N_17061,N_16767,N_16136);
or U17062 (N_17062,N_16757,N_16754);
or U17063 (N_17063,N_16021,N_16536);
xor U17064 (N_17064,N_16271,N_16237);
nor U17065 (N_17065,N_16216,N_16389);
nand U17066 (N_17066,N_16559,N_16482);
nand U17067 (N_17067,N_16775,N_16583);
xnor U17068 (N_17068,N_16156,N_16094);
or U17069 (N_17069,N_16495,N_16079);
nor U17070 (N_17070,N_16784,N_16512);
nand U17071 (N_17071,N_16402,N_16043);
or U17072 (N_17072,N_16398,N_16506);
or U17073 (N_17073,N_16436,N_16031);
nor U17074 (N_17074,N_16620,N_16139);
nand U17075 (N_17075,N_16385,N_16032);
nand U17076 (N_17076,N_16126,N_16144);
xnor U17077 (N_17077,N_16152,N_16254);
or U17078 (N_17078,N_16181,N_16710);
nand U17079 (N_17079,N_16543,N_16278);
nor U17080 (N_17080,N_16774,N_16114);
nand U17081 (N_17081,N_16014,N_16492);
or U17082 (N_17082,N_16409,N_16327);
nor U17083 (N_17083,N_16753,N_16420);
xnor U17084 (N_17084,N_16567,N_16587);
nor U17085 (N_17085,N_16441,N_16573);
and U17086 (N_17086,N_16381,N_16412);
nand U17087 (N_17087,N_16397,N_16591);
xnor U17088 (N_17088,N_16219,N_16719);
nor U17089 (N_17089,N_16016,N_16752);
and U17090 (N_17090,N_16187,N_16256);
or U17091 (N_17091,N_16051,N_16632);
and U17092 (N_17092,N_16705,N_16281);
and U17093 (N_17093,N_16286,N_16342);
xor U17094 (N_17094,N_16235,N_16472);
or U17095 (N_17095,N_16457,N_16068);
nand U17096 (N_17096,N_16146,N_16153);
or U17097 (N_17097,N_16308,N_16739);
or U17098 (N_17098,N_16065,N_16163);
nor U17099 (N_17099,N_16301,N_16525);
or U17100 (N_17100,N_16683,N_16059);
and U17101 (N_17101,N_16325,N_16177);
xor U17102 (N_17102,N_16336,N_16785);
xor U17103 (N_17103,N_16714,N_16681);
or U17104 (N_17104,N_16724,N_16285);
nor U17105 (N_17105,N_16729,N_16204);
or U17106 (N_17106,N_16535,N_16019);
or U17107 (N_17107,N_16269,N_16010);
and U17108 (N_17108,N_16476,N_16135);
nor U17109 (N_17109,N_16154,N_16673);
nand U17110 (N_17110,N_16526,N_16185);
xnor U17111 (N_17111,N_16637,N_16460);
xnor U17112 (N_17112,N_16013,N_16159);
nor U17113 (N_17113,N_16545,N_16796);
or U17114 (N_17114,N_16642,N_16150);
nor U17115 (N_17115,N_16141,N_16575);
and U17116 (N_17116,N_16243,N_16550);
xor U17117 (N_17117,N_16561,N_16036);
and U17118 (N_17118,N_16106,N_16186);
or U17119 (N_17119,N_16391,N_16423);
nand U17120 (N_17120,N_16740,N_16034);
xor U17121 (N_17121,N_16527,N_16377);
xor U17122 (N_17122,N_16131,N_16321);
and U17123 (N_17123,N_16660,N_16372);
or U17124 (N_17124,N_16090,N_16162);
and U17125 (N_17125,N_16772,N_16566);
nor U17126 (N_17126,N_16240,N_16747);
nor U17127 (N_17127,N_16112,N_16491);
and U17128 (N_17128,N_16780,N_16399);
and U17129 (N_17129,N_16410,N_16760);
nor U17130 (N_17130,N_16734,N_16640);
nand U17131 (N_17131,N_16782,N_16258);
nor U17132 (N_17132,N_16011,N_16568);
nor U17133 (N_17133,N_16712,N_16331);
nand U17134 (N_17134,N_16306,N_16425);
xor U17135 (N_17135,N_16732,N_16155);
xnor U17136 (N_17136,N_16132,N_16548);
or U17137 (N_17137,N_16221,N_16731);
and U17138 (N_17138,N_16282,N_16081);
xor U17139 (N_17139,N_16238,N_16588);
nor U17140 (N_17140,N_16037,N_16161);
and U17141 (N_17141,N_16320,N_16717);
nor U17142 (N_17142,N_16577,N_16190);
nor U17143 (N_17143,N_16701,N_16498);
or U17144 (N_17144,N_16596,N_16622);
or U17145 (N_17145,N_16198,N_16070);
nand U17146 (N_17146,N_16149,N_16142);
or U17147 (N_17147,N_16246,N_16128);
or U17148 (N_17148,N_16175,N_16686);
xor U17149 (N_17149,N_16413,N_16214);
nand U17150 (N_17150,N_16168,N_16790);
or U17151 (N_17151,N_16722,N_16407);
or U17152 (N_17152,N_16361,N_16703);
nor U17153 (N_17153,N_16236,N_16493);
nand U17154 (N_17154,N_16530,N_16359);
or U17155 (N_17155,N_16589,N_16502);
and U17156 (N_17156,N_16255,N_16557);
nor U17157 (N_17157,N_16499,N_16655);
xnor U17158 (N_17158,N_16004,N_16020);
nand U17159 (N_17159,N_16057,N_16277);
xor U17160 (N_17160,N_16581,N_16490);
nor U17161 (N_17161,N_16353,N_16313);
and U17162 (N_17162,N_16369,N_16636);
and U17163 (N_17163,N_16688,N_16574);
nand U17164 (N_17164,N_16273,N_16601);
nand U17165 (N_17165,N_16358,N_16213);
nor U17166 (N_17166,N_16288,N_16467);
nand U17167 (N_17167,N_16073,N_16054);
nand U17168 (N_17168,N_16444,N_16462);
and U17169 (N_17169,N_16388,N_16176);
xor U17170 (N_17170,N_16344,N_16228);
nand U17171 (N_17171,N_16015,N_16210);
and U17172 (N_17172,N_16483,N_16698);
or U17173 (N_17173,N_16056,N_16042);
or U17174 (N_17174,N_16041,N_16111);
nor U17175 (N_17175,N_16029,N_16172);
nand U17176 (N_17176,N_16625,N_16578);
nor U17177 (N_17177,N_16786,N_16027);
nor U17178 (N_17178,N_16500,N_16025);
nand U17179 (N_17179,N_16418,N_16507);
nor U17180 (N_17180,N_16317,N_16164);
nand U17181 (N_17181,N_16538,N_16706);
and U17182 (N_17182,N_16733,N_16337);
xnor U17183 (N_17183,N_16193,N_16456);
nor U17184 (N_17184,N_16382,N_16599);
xor U17185 (N_17185,N_16452,N_16463);
or U17186 (N_17186,N_16343,N_16534);
nor U17187 (N_17187,N_16762,N_16585);
or U17188 (N_17188,N_16448,N_16776);
or U17189 (N_17189,N_16608,N_16496);
and U17190 (N_17190,N_16370,N_16044);
nor U17191 (N_17191,N_16662,N_16045);
and U17192 (N_17192,N_16435,N_16018);
nand U17193 (N_17193,N_16532,N_16401);
xor U17194 (N_17194,N_16434,N_16346);
nand U17195 (N_17195,N_16665,N_16275);
nor U17196 (N_17196,N_16259,N_16748);
and U17197 (N_17197,N_16619,N_16099);
or U17198 (N_17198,N_16170,N_16726);
xor U17199 (N_17199,N_16024,N_16781);
or U17200 (N_17200,N_16609,N_16772);
xnor U17201 (N_17201,N_16298,N_16202);
nand U17202 (N_17202,N_16149,N_16467);
xnor U17203 (N_17203,N_16692,N_16260);
and U17204 (N_17204,N_16698,N_16390);
nand U17205 (N_17205,N_16581,N_16287);
nor U17206 (N_17206,N_16484,N_16236);
xor U17207 (N_17207,N_16304,N_16688);
xnor U17208 (N_17208,N_16432,N_16729);
xnor U17209 (N_17209,N_16074,N_16170);
nor U17210 (N_17210,N_16527,N_16075);
xnor U17211 (N_17211,N_16311,N_16625);
nand U17212 (N_17212,N_16500,N_16794);
xnor U17213 (N_17213,N_16581,N_16025);
nand U17214 (N_17214,N_16289,N_16475);
nand U17215 (N_17215,N_16151,N_16663);
nor U17216 (N_17216,N_16696,N_16770);
nand U17217 (N_17217,N_16295,N_16169);
nand U17218 (N_17218,N_16515,N_16798);
or U17219 (N_17219,N_16289,N_16699);
xor U17220 (N_17220,N_16207,N_16412);
xnor U17221 (N_17221,N_16231,N_16017);
xor U17222 (N_17222,N_16534,N_16681);
and U17223 (N_17223,N_16455,N_16183);
or U17224 (N_17224,N_16543,N_16181);
nor U17225 (N_17225,N_16472,N_16588);
xnor U17226 (N_17226,N_16091,N_16359);
or U17227 (N_17227,N_16315,N_16755);
and U17228 (N_17228,N_16054,N_16739);
nor U17229 (N_17229,N_16004,N_16420);
nand U17230 (N_17230,N_16083,N_16449);
and U17231 (N_17231,N_16731,N_16372);
and U17232 (N_17232,N_16742,N_16074);
nor U17233 (N_17233,N_16246,N_16794);
and U17234 (N_17234,N_16411,N_16097);
or U17235 (N_17235,N_16731,N_16291);
nor U17236 (N_17236,N_16253,N_16339);
or U17237 (N_17237,N_16025,N_16458);
or U17238 (N_17238,N_16351,N_16535);
xnor U17239 (N_17239,N_16100,N_16588);
nand U17240 (N_17240,N_16685,N_16741);
nand U17241 (N_17241,N_16400,N_16013);
nand U17242 (N_17242,N_16411,N_16535);
nor U17243 (N_17243,N_16378,N_16621);
nor U17244 (N_17244,N_16278,N_16262);
nand U17245 (N_17245,N_16400,N_16346);
xor U17246 (N_17246,N_16350,N_16033);
and U17247 (N_17247,N_16276,N_16786);
xor U17248 (N_17248,N_16088,N_16263);
xnor U17249 (N_17249,N_16156,N_16322);
and U17250 (N_17250,N_16204,N_16357);
or U17251 (N_17251,N_16645,N_16214);
nor U17252 (N_17252,N_16574,N_16206);
xnor U17253 (N_17253,N_16506,N_16294);
nor U17254 (N_17254,N_16416,N_16326);
or U17255 (N_17255,N_16234,N_16687);
and U17256 (N_17256,N_16510,N_16544);
or U17257 (N_17257,N_16232,N_16757);
nand U17258 (N_17258,N_16490,N_16659);
and U17259 (N_17259,N_16360,N_16708);
or U17260 (N_17260,N_16470,N_16511);
nor U17261 (N_17261,N_16630,N_16760);
or U17262 (N_17262,N_16265,N_16021);
xnor U17263 (N_17263,N_16019,N_16300);
xnor U17264 (N_17264,N_16295,N_16115);
xor U17265 (N_17265,N_16759,N_16459);
nand U17266 (N_17266,N_16724,N_16792);
xor U17267 (N_17267,N_16011,N_16495);
nor U17268 (N_17268,N_16453,N_16461);
xnor U17269 (N_17269,N_16607,N_16551);
or U17270 (N_17270,N_16663,N_16374);
and U17271 (N_17271,N_16175,N_16583);
or U17272 (N_17272,N_16257,N_16116);
nand U17273 (N_17273,N_16444,N_16443);
and U17274 (N_17274,N_16438,N_16337);
and U17275 (N_17275,N_16222,N_16378);
and U17276 (N_17276,N_16603,N_16024);
nand U17277 (N_17277,N_16299,N_16221);
or U17278 (N_17278,N_16308,N_16754);
xor U17279 (N_17279,N_16650,N_16060);
xor U17280 (N_17280,N_16428,N_16095);
or U17281 (N_17281,N_16758,N_16430);
nand U17282 (N_17282,N_16176,N_16782);
nand U17283 (N_17283,N_16283,N_16658);
nand U17284 (N_17284,N_16296,N_16213);
xor U17285 (N_17285,N_16332,N_16695);
and U17286 (N_17286,N_16549,N_16285);
nand U17287 (N_17287,N_16391,N_16723);
and U17288 (N_17288,N_16456,N_16585);
nor U17289 (N_17289,N_16559,N_16646);
nand U17290 (N_17290,N_16684,N_16251);
or U17291 (N_17291,N_16579,N_16739);
xnor U17292 (N_17292,N_16334,N_16054);
nor U17293 (N_17293,N_16365,N_16100);
xor U17294 (N_17294,N_16684,N_16431);
or U17295 (N_17295,N_16121,N_16483);
or U17296 (N_17296,N_16471,N_16531);
nand U17297 (N_17297,N_16647,N_16155);
or U17298 (N_17298,N_16439,N_16731);
or U17299 (N_17299,N_16185,N_16091);
nor U17300 (N_17300,N_16221,N_16059);
nand U17301 (N_17301,N_16007,N_16273);
nand U17302 (N_17302,N_16040,N_16359);
or U17303 (N_17303,N_16257,N_16328);
or U17304 (N_17304,N_16450,N_16696);
or U17305 (N_17305,N_16380,N_16695);
and U17306 (N_17306,N_16712,N_16626);
and U17307 (N_17307,N_16113,N_16314);
xnor U17308 (N_17308,N_16085,N_16419);
and U17309 (N_17309,N_16522,N_16375);
nor U17310 (N_17310,N_16330,N_16315);
xor U17311 (N_17311,N_16102,N_16444);
xnor U17312 (N_17312,N_16253,N_16519);
nand U17313 (N_17313,N_16757,N_16204);
xnor U17314 (N_17314,N_16319,N_16046);
and U17315 (N_17315,N_16768,N_16640);
and U17316 (N_17316,N_16480,N_16466);
and U17317 (N_17317,N_16385,N_16271);
nand U17318 (N_17318,N_16128,N_16092);
nand U17319 (N_17319,N_16092,N_16461);
nor U17320 (N_17320,N_16796,N_16132);
nor U17321 (N_17321,N_16095,N_16241);
xnor U17322 (N_17322,N_16154,N_16123);
xnor U17323 (N_17323,N_16430,N_16658);
or U17324 (N_17324,N_16209,N_16157);
or U17325 (N_17325,N_16192,N_16282);
nor U17326 (N_17326,N_16096,N_16090);
or U17327 (N_17327,N_16760,N_16263);
nand U17328 (N_17328,N_16209,N_16238);
nor U17329 (N_17329,N_16056,N_16275);
or U17330 (N_17330,N_16576,N_16280);
and U17331 (N_17331,N_16684,N_16304);
nor U17332 (N_17332,N_16186,N_16783);
xnor U17333 (N_17333,N_16716,N_16113);
or U17334 (N_17334,N_16797,N_16465);
nand U17335 (N_17335,N_16295,N_16732);
and U17336 (N_17336,N_16479,N_16290);
or U17337 (N_17337,N_16229,N_16552);
nand U17338 (N_17338,N_16322,N_16068);
nand U17339 (N_17339,N_16175,N_16596);
xnor U17340 (N_17340,N_16266,N_16731);
or U17341 (N_17341,N_16466,N_16051);
xnor U17342 (N_17342,N_16028,N_16052);
nand U17343 (N_17343,N_16260,N_16118);
or U17344 (N_17344,N_16503,N_16627);
and U17345 (N_17345,N_16264,N_16315);
nand U17346 (N_17346,N_16017,N_16026);
nand U17347 (N_17347,N_16546,N_16184);
and U17348 (N_17348,N_16607,N_16186);
or U17349 (N_17349,N_16238,N_16661);
and U17350 (N_17350,N_16648,N_16410);
or U17351 (N_17351,N_16298,N_16231);
and U17352 (N_17352,N_16706,N_16055);
or U17353 (N_17353,N_16463,N_16022);
xnor U17354 (N_17354,N_16120,N_16139);
nand U17355 (N_17355,N_16632,N_16092);
and U17356 (N_17356,N_16372,N_16598);
and U17357 (N_17357,N_16767,N_16676);
and U17358 (N_17358,N_16106,N_16438);
nor U17359 (N_17359,N_16323,N_16459);
xor U17360 (N_17360,N_16020,N_16152);
and U17361 (N_17361,N_16275,N_16717);
nand U17362 (N_17362,N_16719,N_16671);
nand U17363 (N_17363,N_16649,N_16102);
xor U17364 (N_17364,N_16420,N_16519);
nor U17365 (N_17365,N_16762,N_16079);
or U17366 (N_17366,N_16160,N_16469);
xnor U17367 (N_17367,N_16151,N_16579);
and U17368 (N_17368,N_16638,N_16735);
nand U17369 (N_17369,N_16457,N_16036);
and U17370 (N_17370,N_16216,N_16270);
nand U17371 (N_17371,N_16528,N_16580);
or U17372 (N_17372,N_16053,N_16754);
nand U17373 (N_17373,N_16296,N_16575);
or U17374 (N_17374,N_16658,N_16367);
and U17375 (N_17375,N_16729,N_16614);
or U17376 (N_17376,N_16628,N_16635);
xor U17377 (N_17377,N_16282,N_16555);
nor U17378 (N_17378,N_16252,N_16798);
nand U17379 (N_17379,N_16375,N_16655);
xor U17380 (N_17380,N_16262,N_16291);
and U17381 (N_17381,N_16646,N_16351);
nand U17382 (N_17382,N_16629,N_16518);
nor U17383 (N_17383,N_16241,N_16130);
and U17384 (N_17384,N_16314,N_16653);
xor U17385 (N_17385,N_16493,N_16450);
nand U17386 (N_17386,N_16515,N_16152);
nor U17387 (N_17387,N_16144,N_16467);
or U17388 (N_17388,N_16509,N_16504);
or U17389 (N_17389,N_16533,N_16290);
nor U17390 (N_17390,N_16735,N_16776);
nand U17391 (N_17391,N_16342,N_16736);
or U17392 (N_17392,N_16208,N_16198);
or U17393 (N_17393,N_16378,N_16182);
nand U17394 (N_17394,N_16499,N_16533);
or U17395 (N_17395,N_16789,N_16546);
and U17396 (N_17396,N_16743,N_16660);
or U17397 (N_17397,N_16290,N_16666);
or U17398 (N_17398,N_16055,N_16732);
or U17399 (N_17399,N_16229,N_16160);
xor U17400 (N_17400,N_16161,N_16555);
and U17401 (N_17401,N_16006,N_16783);
xnor U17402 (N_17402,N_16049,N_16727);
nand U17403 (N_17403,N_16660,N_16356);
nand U17404 (N_17404,N_16004,N_16189);
nor U17405 (N_17405,N_16715,N_16407);
and U17406 (N_17406,N_16193,N_16534);
xor U17407 (N_17407,N_16227,N_16753);
and U17408 (N_17408,N_16636,N_16022);
nor U17409 (N_17409,N_16147,N_16575);
or U17410 (N_17410,N_16763,N_16658);
nand U17411 (N_17411,N_16444,N_16193);
and U17412 (N_17412,N_16167,N_16350);
xnor U17413 (N_17413,N_16774,N_16590);
and U17414 (N_17414,N_16762,N_16695);
xor U17415 (N_17415,N_16770,N_16119);
nor U17416 (N_17416,N_16313,N_16129);
nand U17417 (N_17417,N_16660,N_16093);
or U17418 (N_17418,N_16088,N_16210);
nand U17419 (N_17419,N_16536,N_16129);
and U17420 (N_17420,N_16755,N_16067);
nor U17421 (N_17421,N_16155,N_16037);
or U17422 (N_17422,N_16183,N_16191);
nor U17423 (N_17423,N_16751,N_16384);
and U17424 (N_17424,N_16740,N_16788);
and U17425 (N_17425,N_16256,N_16666);
xor U17426 (N_17426,N_16761,N_16070);
or U17427 (N_17427,N_16406,N_16414);
nand U17428 (N_17428,N_16432,N_16629);
nand U17429 (N_17429,N_16612,N_16706);
nor U17430 (N_17430,N_16706,N_16154);
nor U17431 (N_17431,N_16374,N_16324);
nand U17432 (N_17432,N_16766,N_16363);
and U17433 (N_17433,N_16245,N_16631);
and U17434 (N_17434,N_16731,N_16322);
nor U17435 (N_17435,N_16098,N_16759);
xor U17436 (N_17436,N_16470,N_16539);
and U17437 (N_17437,N_16400,N_16452);
nor U17438 (N_17438,N_16449,N_16372);
xnor U17439 (N_17439,N_16518,N_16237);
xor U17440 (N_17440,N_16636,N_16325);
and U17441 (N_17441,N_16069,N_16589);
nor U17442 (N_17442,N_16231,N_16527);
and U17443 (N_17443,N_16600,N_16049);
nand U17444 (N_17444,N_16041,N_16259);
nand U17445 (N_17445,N_16421,N_16434);
xor U17446 (N_17446,N_16170,N_16691);
nand U17447 (N_17447,N_16142,N_16724);
and U17448 (N_17448,N_16594,N_16063);
nor U17449 (N_17449,N_16668,N_16477);
xnor U17450 (N_17450,N_16535,N_16782);
nor U17451 (N_17451,N_16139,N_16412);
and U17452 (N_17452,N_16135,N_16732);
nand U17453 (N_17453,N_16776,N_16316);
and U17454 (N_17454,N_16224,N_16045);
nor U17455 (N_17455,N_16256,N_16160);
nor U17456 (N_17456,N_16258,N_16473);
xor U17457 (N_17457,N_16764,N_16440);
and U17458 (N_17458,N_16431,N_16134);
and U17459 (N_17459,N_16221,N_16468);
nor U17460 (N_17460,N_16170,N_16217);
and U17461 (N_17461,N_16607,N_16452);
and U17462 (N_17462,N_16391,N_16238);
or U17463 (N_17463,N_16341,N_16417);
nor U17464 (N_17464,N_16159,N_16696);
and U17465 (N_17465,N_16345,N_16327);
xnor U17466 (N_17466,N_16597,N_16402);
xnor U17467 (N_17467,N_16226,N_16717);
or U17468 (N_17468,N_16520,N_16328);
xnor U17469 (N_17469,N_16709,N_16033);
and U17470 (N_17470,N_16602,N_16012);
nand U17471 (N_17471,N_16771,N_16105);
or U17472 (N_17472,N_16362,N_16439);
nand U17473 (N_17473,N_16209,N_16555);
and U17474 (N_17474,N_16734,N_16546);
nor U17475 (N_17475,N_16485,N_16602);
xor U17476 (N_17476,N_16270,N_16721);
and U17477 (N_17477,N_16401,N_16434);
nor U17478 (N_17478,N_16471,N_16194);
and U17479 (N_17479,N_16526,N_16730);
or U17480 (N_17480,N_16420,N_16792);
xor U17481 (N_17481,N_16357,N_16183);
nor U17482 (N_17482,N_16055,N_16135);
nor U17483 (N_17483,N_16191,N_16636);
or U17484 (N_17484,N_16607,N_16333);
nand U17485 (N_17485,N_16728,N_16346);
xnor U17486 (N_17486,N_16758,N_16270);
nor U17487 (N_17487,N_16106,N_16413);
or U17488 (N_17488,N_16704,N_16656);
nor U17489 (N_17489,N_16580,N_16412);
xor U17490 (N_17490,N_16100,N_16145);
and U17491 (N_17491,N_16081,N_16021);
and U17492 (N_17492,N_16027,N_16367);
or U17493 (N_17493,N_16085,N_16465);
nor U17494 (N_17494,N_16024,N_16011);
xor U17495 (N_17495,N_16357,N_16154);
or U17496 (N_17496,N_16369,N_16471);
and U17497 (N_17497,N_16497,N_16057);
xnor U17498 (N_17498,N_16762,N_16380);
and U17499 (N_17499,N_16662,N_16027);
nor U17500 (N_17500,N_16461,N_16309);
and U17501 (N_17501,N_16227,N_16705);
nand U17502 (N_17502,N_16571,N_16451);
nand U17503 (N_17503,N_16036,N_16554);
xor U17504 (N_17504,N_16674,N_16138);
nor U17505 (N_17505,N_16049,N_16252);
nand U17506 (N_17506,N_16264,N_16293);
and U17507 (N_17507,N_16686,N_16244);
or U17508 (N_17508,N_16363,N_16050);
nand U17509 (N_17509,N_16787,N_16029);
xor U17510 (N_17510,N_16118,N_16456);
nand U17511 (N_17511,N_16343,N_16270);
nand U17512 (N_17512,N_16193,N_16138);
nand U17513 (N_17513,N_16380,N_16005);
or U17514 (N_17514,N_16285,N_16731);
xnor U17515 (N_17515,N_16064,N_16464);
nor U17516 (N_17516,N_16523,N_16066);
nor U17517 (N_17517,N_16313,N_16411);
nand U17518 (N_17518,N_16097,N_16033);
nand U17519 (N_17519,N_16499,N_16329);
nor U17520 (N_17520,N_16394,N_16334);
xnor U17521 (N_17521,N_16582,N_16678);
or U17522 (N_17522,N_16449,N_16287);
nor U17523 (N_17523,N_16049,N_16372);
nor U17524 (N_17524,N_16597,N_16143);
nand U17525 (N_17525,N_16500,N_16017);
nor U17526 (N_17526,N_16144,N_16013);
and U17527 (N_17527,N_16051,N_16007);
and U17528 (N_17528,N_16223,N_16628);
xor U17529 (N_17529,N_16519,N_16090);
nand U17530 (N_17530,N_16687,N_16177);
nand U17531 (N_17531,N_16591,N_16177);
nor U17532 (N_17532,N_16479,N_16274);
and U17533 (N_17533,N_16520,N_16713);
or U17534 (N_17534,N_16004,N_16467);
nand U17535 (N_17535,N_16123,N_16053);
xor U17536 (N_17536,N_16307,N_16697);
nor U17537 (N_17537,N_16056,N_16276);
and U17538 (N_17538,N_16023,N_16357);
nand U17539 (N_17539,N_16122,N_16219);
xor U17540 (N_17540,N_16053,N_16649);
nand U17541 (N_17541,N_16709,N_16057);
nor U17542 (N_17542,N_16162,N_16741);
or U17543 (N_17543,N_16258,N_16390);
nor U17544 (N_17544,N_16599,N_16131);
xnor U17545 (N_17545,N_16130,N_16486);
nor U17546 (N_17546,N_16625,N_16726);
nand U17547 (N_17547,N_16664,N_16773);
nand U17548 (N_17548,N_16367,N_16716);
xor U17549 (N_17549,N_16374,N_16207);
and U17550 (N_17550,N_16610,N_16205);
xor U17551 (N_17551,N_16499,N_16079);
nor U17552 (N_17552,N_16232,N_16097);
nor U17553 (N_17553,N_16174,N_16580);
xor U17554 (N_17554,N_16286,N_16133);
nand U17555 (N_17555,N_16613,N_16579);
and U17556 (N_17556,N_16147,N_16361);
nand U17557 (N_17557,N_16103,N_16533);
and U17558 (N_17558,N_16516,N_16420);
nand U17559 (N_17559,N_16242,N_16332);
xor U17560 (N_17560,N_16736,N_16157);
and U17561 (N_17561,N_16248,N_16556);
and U17562 (N_17562,N_16215,N_16424);
nor U17563 (N_17563,N_16743,N_16601);
xor U17564 (N_17564,N_16177,N_16700);
nand U17565 (N_17565,N_16383,N_16745);
nand U17566 (N_17566,N_16396,N_16444);
nor U17567 (N_17567,N_16345,N_16116);
nand U17568 (N_17568,N_16685,N_16790);
or U17569 (N_17569,N_16598,N_16601);
or U17570 (N_17570,N_16489,N_16366);
and U17571 (N_17571,N_16099,N_16571);
or U17572 (N_17572,N_16427,N_16613);
nand U17573 (N_17573,N_16263,N_16504);
and U17574 (N_17574,N_16348,N_16095);
and U17575 (N_17575,N_16507,N_16496);
or U17576 (N_17576,N_16616,N_16162);
or U17577 (N_17577,N_16121,N_16423);
or U17578 (N_17578,N_16604,N_16179);
nor U17579 (N_17579,N_16738,N_16394);
nand U17580 (N_17580,N_16659,N_16680);
and U17581 (N_17581,N_16542,N_16558);
and U17582 (N_17582,N_16579,N_16689);
or U17583 (N_17583,N_16199,N_16019);
xor U17584 (N_17584,N_16163,N_16325);
xnor U17585 (N_17585,N_16575,N_16756);
nand U17586 (N_17586,N_16668,N_16436);
nand U17587 (N_17587,N_16663,N_16437);
nand U17588 (N_17588,N_16017,N_16251);
xor U17589 (N_17589,N_16071,N_16612);
or U17590 (N_17590,N_16276,N_16411);
nor U17591 (N_17591,N_16377,N_16659);
and U17592 (N_17592,N_16095,N_16000);
nor U17593 (N_17593,N_16347,N_16540);
and U17594 (N_17594,N_16417,N_16638);
nand U17595 (N_17595,N_16221,N_16145);
or U17596 (N_17596,N_16166,N_16023);
xnor U17597 (N_17597,N_16230,N_16457);
or U17598 (N_17598,N_16471,N_16520);
and U17599 (N_17599,N_16242,N_16063);
and U17600 (N_17600,N_17444,N_16819);
nand U17601 (N_17601,N_17085,N_17520);
nand U17602 (N_17602,N_16858,N_17031);
and U17603 (N_17603,N_16887,N_17409);
nor U17604 (N_17604,N_17076,N_16910);
nand U17605 (N_17605,N_17326,N_17412);
and U17606 (N_17606,N_17257,N_17224);
or U17607 (N_17607,N_17228,N_17267);
nand U17608 (N_17608,N_17423,N_17499);
or U17609 (N_17609,N_17103,N_16845);
and U17610 (N_17610,N_17390,N_17157);
or U17611 (N_17611,N_16982,N_17160);
nor U17612 (N_17612,N_16876,N_17335);
xor U17613 (N_17613,N_16963,N_17402);
xor U17614 (N_17614,N_17300,N_17020);
xor U17615 (N_17615,N_17133,N_17273);
or U17616 (N_17616,N_17355,N_17029);
nor U17617 (N_17617,N_17285,N_16960);
nand U17618 (N_17618,N_16864,N_16968);
xor U17619 (N_17619,N_17045,N_17361);
xnor U17620 (N_17620,N_17012,N_17465);
nor U17621 (N_17621,N_17459,N_17496);
nor U17622 (N_17622,N_17566,N_17422);
and U17623 (N_17623,N_17225,N_17147);
nor U17624 (N_17624,N_16824,N_16911);
and U17625 (N_17625,N_17251,N_17275);
or U17626 (N_17626,N_17396,N_17044);
nand U17627 (N_17627,N_17311,N_16892);
xnor U17628 (N_17628,N_17407,N_17441);
or U17629 (N_17629,N_17420,N_17097);
nand U17630 (N_17630,N_17486,N_17101);
and U17631 (N_17631,N_17377,N_17120);
nand U17632 (N_17632,N_16801,N_17021);
and U17633 (N_17633,N_16987,N_17122);
xnor U17634 (N_17634,N_17127,N_17540);
or U17635 (N_17635,N_16804,N_17589);
nor U17636 (N_17636,N_16961,N_17588);
or U17637 (N_17637,N_16934,N_17027);
or U17638 (N_17638,N_17202,N_17568);
nor U17639 (N_17639,N_17339,N_17107);
xor U17640 (N_17640,N_17570,N_17585);
xor U17641 (N_17641,N_17388,N_17395);
xor U17642 (N_17642,N_17450,N_16909);
and U17643 (N_17643,N_17093,N_17091);
and U17644 (N_17644,N_17517,N_17236);
nand U17645 (N_17645,N_16886,N_16991);
xnor U17646 (N_17646,N_17515,N_17479);
and U17647 (N_17647,N_17067,N_16998);
nand U17648 (N_17648,N_16914,N_16924);
or U17649 (N_17649,N_16955,N_17200);
nand U17650 (N_17650,N_17382,N_17197);
or U17651 (N_17651,N_17293,N_17469);
nor U17652 (N_17652,N_17130,N_16931);
nor U17653 (N_17653,N_17061,N_17146);
nand U17654 (N_17654,N_17211,N_17424);
or U17655 (N_17655,N_17547,N_17064);
nor U17656 (N_17656,N_16832,N_16981);
or U17657 (N_17657,N_17221,N_17204);
nand U17658 (N_17658,N_17456,N_17095);
nand U17659 (N_17659,N_17105,N_16994);
nor U17660 (N_17660,N_16992,N_16975);
xor U17661 (N_17661,N_17266,N_17309);
and U17662 (N_17662,N_17244,N_17381);
xor U17663 (N_17663,N_17449,N_17043);
xor U17664 (N_17664,N_17376,N_16962);
or U17665 (N_17665,N_16965,N_17360);
xnor U17666 (N_17666,N_16927,N_17239);
nand U17667 (N_17667,N_16812,N_17063);
xnor U17668 (N_17668,N_17528,N_16966);
nor U17669 (N_17669,N_17443,N_17233);
nand U17670 (N_17670,N_17324,N_17089);
xnor U17671 (N_17671,N_17578,N_17159);
xnor U17672 (N_17672,N_17128,N_16802);
nand U17673 (N_17673,N_16875,N_16890);
xnor U17674 (N_17674,N_16995,N_17158);
and U17675 (N_17675,N_16907,N_17037);
nand U17676 (N_17676,N_17370,N_17113);
nor U17677 (N_17677,N_17596,N_17576);
nand U17678 (N_17678,N_16929,N_17018);
and U17679 (N_17679,N_17425,N_17152);
xor U17680 (N_17680,N_17172,N_17003);
nor U17681 (N_17681,N_17271,N_17489);
nand U17682 (N_17682,N_17567,N_16850);
nand U17683 (N_17683,N_17183,N_16888);
nor U17684 (N_17684,N_17561,N_16808);
or U17685 (N_17685,N_17374,N_17321);
xor U17686 (N_17686,N_16904,N_17344);
and U17687 (N_17687,N_17419,N_17332);
nor U17688 (N_17688,N_17573,N_17303);
nor U17689 (N_17689,N_17090,N_16996);
nor U17690 (N_17690,N_17312,N_16879);
or U17691 (N_17691,N_17306,N_17587);
and U17692 (N_17692,N_17473,N_17041);
or U17693 (N_17693,N_17060,N_16997);
or U17694 (N_17694,N_16829,N_17535);
and U17695 (N_17695,N_17357,N_16868);
nor U17696 (N_17696,N_17466,N_17206);
xnor U17697 (N_17697,N_17119,N_16811);
nand U17698 (N_17698,N_17592,N_17294);
or U17699 (N_17699,N_17049,N_16878);
and U17700 (N_17700,N_17560,N_17070);
and U17701 (N_17701,N_17546,N_17150);
xor U17702 (N_17702,N_17416,N_17401);
nor U17703 (N_17703,N_16843,N_17558);
xnor U17704 (N_17704,N_17557,N_17284);
nand U17705 (N_17705,N_17028,N_16990);
or U17706 (N_17706,N_17171,N_17092);
nor U17707 (N_17707,N_17391,N_17350);
nor U17708 (N_17708,N_17077,N_16932);
and U17709 (N_17709,N_17575,N_17565);
or U17710 (N_17710,N_17156,N_17138);
nor U17711 (N_17711,N_17212,N_17081);
nor U17712 (N_17712,N_17252,N_17518);
nor U17713 (N_17713,N_16891,N_16857);
or U17714 (N_17714,N_17161,N_17162);
or U17715 (N_17715,N_17265,N_17563);
nor U17716 (N_17716,N_17232,N_17347);
xnor U17717 (N_17717,N_17590,N_17203);
nand U17718 (N_17718,N_17214,N_17322);
nand U17719 (N_17719,N_17551,N_16814);
or U17720 (N_17720,N_16984,N_17166);
nand U17721 (N_17721,N_17512,N_17054);
nand U17722 (N_17722,N_16815,N_17259);
and U17723 (N_17723,N_16828,N_17522);
nor U17724 (N_17724,N_17510,N_17210);
xor U17725 (N_17725,N_17421,N_17414);
nand U17726 (N_17726,N_17559,N_17231);
nand U17727 (N_17727,N_17383,N_17562);
nor U17728 (N_17728,N_17513,N_17554);
or U17729 (N_17729,N_17485,N_17073);
xnor U17730 (N_17730,N_17436,N_17190);
or U17731 (N_17731,N_17291,N_17249);
or U17732 (N_17732,N_17051,N_17597);
and U17733 (N_17733,N_17532,N_17218);
nand U17734 (N_17734,N_17536,N_17223);
or U17735 (N_17735,N_17329,N_16883);
nand U17736 (N_17736,N_17062,N_17142);
or U17737 (N_17737,N_17181,N_17048);
or U17738 (N_17738,N_17507,N_16822);
and U17739 (N_17739,N_17296,N_17386);
or U17740 (N_17740,N_16851,N_17487);
and U17741 (N_17741,N_17253,N_16936);
nor U17742 (N_17742,N_17032,N_17235);
xor U17743 (N_17743,N_17299,N_17505);
xor U17744 (N_17744,N_17534,N_17539);
xnor U17745 (N_17745,N_17508,N_17277);
nand U17746 (N_17746,N_17019,N_17433);
xnor U17747 (N_17747,N_16830,N_17581);
nand U17748 (N_17748,N_17470,N_16841);
xnor U17749 (N_17749,N_17260,N_17272);
xnor U17750 (N_17750,N_16947,N_17006);
and U17751 (N_17751,N_17036,N_16921);
nand U17752 (N_17752,N_17217,N_17030);
nand U17753 (N_17753,N_16977,N_17055);
xnor U17754 (N_17754,N_17213,N_17178);
or U17755 (N_17755,N_17179,N_17463);
and U17756 (N_17756,N_17230,N_17106);
xor U17757 (N_17757,N_16827,N_17112);
xnor U17758 (N_17758,N_16948,N_17325);
nor U17759 (N_17759,N_17102,N_16854);
nor U17760 (N_17760,N_17464,N_17298);
xor U17761 (N_17761,N_16897,N_17504);
or U17762 (N_17762,N_17269,N_17279);
and U17763 (N_17763,N_17186,N_17410);
or U17764 (N_17764,N_17569,N_17083);
nor U17765 (N_17765,N_16835,N_17457);
xor U17766 (N_17766,N_17593,N_17368);
nand U17767 (N_17767,N_17509,N_16809);
and U17768 (N_17768,N_17313,N_17109);
xor U17769 (N_17769,N_17201,N_16923);
xnor U17770 (N_17770,N_17584,N_16976);
or U17771 (N_17771,N_17553,N_16860);
xor U17772 (N_17772,N_16800,N_17154);
and U17773 (N_17773,N_17008,N_17595);
nor U17774 (N_17774,N_16951,N_17448);
and U17775 (N_17775,N_17022,N_16874);
and U17776 (N_17776,N_17319,N_16944);
xnor U17777 (N_17777,N_16908,N_17148);
nand U17778 (N_17778,N_16949,N_16870);
xnor U17779 (N_17779,N_16837,N_17174);
nand U17780 (N_17780,N_17490,N_17367);
and U17781 (N_17781,N_17432,N_17491);
or U17782 (N_17782,N_17538,N_17187);
xnor U17783 (N_17783,N_17256,N_16928);
xor U17784 (N_17784,N_16872,N_17115);
xnor U17785 (N_17785,N_17582,N_16983);
and U17786 (N_17786,N_17346,N_17591);
nor U17787 (N_17787,N_17488,N_17276);
and U17788 (N_17788,N_17192,N_17164);
nand U17789 (N_17789,N_16861,N_17058);
nor U17790 (N_17790,N_17482,N_17389);
and U17791 (N_17791,N_17379,N_16852);
nand U17792 (N_17792,N_17467,N_17461);
xor U17793 (N_17793,N_16974,N_17431);
nand U17794 (N_17794,N_17086,N_17384);
xor U17795 (N_17795,N_17428,N_17042);
or U17796 (N_17796,N_16865,N_17140);
nand U17797 (N_17797,N_17177,N_16902);
nand U17798 (N_17798,N_16894,N_17435);
and U17799 (N_17799,N_16853,N_17168);
nand U17800 (N_17800,N_17182,N_17193);
xnor U17801 (N_17801,N_17046,N_17352);
nand U17802 (N_17802,N_17100,N_17413);
or U17803 (N_17803,N_16935,N_17264);
and U17804 (N_17804,N_17438,N_17365);
xnor U17805 (N_17805,N_17574,N_16958);
xnor U17806 (N_17806,N_17447,N_17243);
and U17807 (N_17807,N_17359,N_17246);
or U17808 (N_17808,N_17472,N_17088);
and U17809 (N_17809,N_16825,N_17380);
xor U17810 (N_17810,N_16986,N_17184);
xor U17811 (N_17811,N_17098,N_17007);
xor U17812 (N_17812,N_17503,N_16813);
xor U17813 (N_17813,N_17533,N_17572);
and U17814 (N_17814,N_17351,N_16880);
and U17815 (N_17815,N_17282,N_17023);
xor U17816 (N_17816,N_16964,N_17445);
or U17817 (N_17817,N_17278,N_17337);
xor U17818 (N_17818,N_17238,N_17016);
or U17819 (N_17819,N_16871,N_16940);
nand U17820 (N_17820,N_17286,N_17247);
xnor U17821 (N_17821,N_17564,N_17366);
and U17822 (N_17822,N_16922,N_17069);
nand U17823 (N_17823,N_17579,N_17341);
nand U17824 (N_17824,N_16877,N_17288);
and U17825 (N_17825,N_17394,N_17099);
and U17826 (N_17826,N_17427,N_17111);
nor U17827 (N_17827,N_16846,N_16945);
and U17828 (N_17828,N_17501,N_17129);
and U17829 (N_17829,N_17270,N_16941);
or U17830 (N_17830,N_17011,N_16919);
nand U17831 (N_17831,N_17527,N_16988);
or U17832 (N_17832,N_16950,N_16842);
nor U17833 (N_17833,N_17400,N_17010);
nor U17834 (N_17834,N_17072,N_17516);
nand U17835 (N_17835,N_17417,N_17131);
or U17836 (N_17836,N_17132,N_16836);
nand U17837 (N_17837,N_17580,N_17118);
or U17838 (N_17838,N_16896,N_17263);
xnor U17839 (N_17839,N_17050,N_17369);
nor U17840 (N_17840,N_17245,N_16859);
and U17841 (N_17841,N_16839,N_17544);
xor U17842 (N_17842,N_17255,N_17362);
nand U17843 (N_17843,N_16920,N_16959);
and U17844 (N_17844,N_17453,N_17340);
nor U17845 (N_17845,N_17468,N_17378);
or U17846 (N_17846,N_17336,N_16834);
and U17847 (N_17847,N_17316,N_16985);
and U17848 (N_17848,N_16942,N_16937);
nor U17849 (N_17849,N_17583,N_16863);
xor U17850 (N_17850,N_17451,N_17165);
xor U17851 (N_17851,N_17258,N_17145);
nand U17852 (N_17852,N_17180,N_16993);
nand U17853 (N_17853,N_17458,N_17078);
and U17854 (N_17854,N_16957,N_16946);
or U17855 (N_17855,N_17219,N_17096);
or U17856 (N_17856,N_17004,N_17195);
nand U17857 (N_17857,N_17215,N_17545);
nor U17858 (N_17858,N_17552,N_17220);
or U17859 (N_17859,N_17025,N_17483);
xnor U17860 (N_17860,N_17477,N_17302);
or U17861 (N_17861,N_17297,N_16972);
and U17862 (N_17862,N_16905,N_16895);
xor U17863 (N_17863,N_16882,N_17139);
or U17864 (N_17864,N_17492,N_17429);
xor U17865 (N_17865,N_17209,N_17250);
nor U17866 (N_17866,N_17315,N_17471);
xnor U17867 (N_17867,N_16881,N_17082);
or U17868 (N_17868,N_17530,N_16806);
xnor U17869 (N_17869,N_17399,N_17017);
or U17870 (N_17870,N_17191,N_17135);
nand U17871 (N_17871,N_17354,N_17405);
or U17872 (N_17872,N_17393,N_17013);
nor U17873 (N_17873,N_17506,N_17542);
or U17874 (N_17874,N_17334,N_17514);
and U17875 (N_17875,N_17480,N_16873);
nand U17876 (N_17876,N_17525,N_16954);
or U17877 (N_17877,N_17434,N_17262);
or U17878 (N_17878,N_16915,N_17571);
and U17879 (N_17879,N_17207,N_17015);
and U17880 (N_17880,N_17363,N_16807);
xor U17881 (N_17881,N_17242,N_17343);
xnor U17882 (N_17882,N_17327,N_17241);
and U17883 (N_17883,N_16979,N_17068);
xor U17884 (N_17884,N_17307,N_17155);
nand U17885 (N_17885,N_16869,N_17353);
nor U17886 (N_17886,N_17124,N_17108);
and U17887 (N_17887,N_17261,N_16840);
or U17888 (N_17888,N_16938,N_17189);
nor U17889 (N_17889,N_16918,N_17053);
nand U17890 (N_17890,N_17455,N_16926);
or U17891 (N_17891,N_17153,N_17237);
nand U17892 (N_17892,N_17454,N_17500);
xor U17893 (N_17893,N_17356,N_17170);
and U17894 (N_17894,N_17196,N_17331);
or U17895 (N_17895,N_17074,N_17310);
and U17896 (N_17896,N_17493,N_17446);
xor U17897 (N_17897,N_17198,N_16884);
nand U17898 (N_17898,N_17033,N_17084);
xnor U17899 (N_17899,N_17372,N_16818);
nand U17900 (N_17900,N_17452,N_16805);
and U17901 (N_17901,N_17439,N_17476);
xnor U17902 (N_17902,N_17586,N_16916);
nor U17903 (N_17903,N_17460,N_17289);
xnor U17904 (N_17904,N_17462,N_17163);
xor U17905 (N_17905,N_17283,N_17349);
and U17906 (N_17906,N_17080,N_16889);
nand U17907 (N_17907,N_17038,N_17397);
and U17908 (N_17908,N_17126,N_16844);
and U17909 (N_17909,N_17328,N_17079);
xnor U17910 (N_17910,N_17556,N_17134);
nor U17911 (N_17911,N_16848,N_17408);
nand U17912 (N_17912,N_17104,N_17281);
nand U17913 (N_17913,N_17136,N_17137);
nand U17914 (N_17914,N_17549,N_17254);
nor U17915 (N_17915,N_17087,N_16900);
xor U17916 (N_17916,N_17317,N_17000);
xnor U17917 (N_17917,N_17066,N_17205);
nand U17918 (N_17918,N_16978,N_16943);
nand U17919 (N_17919,N_17226,N_17039);
or U17920 (N_17920,N_17345,N_17519);
xor U17921 (N_17921,N_17009,N_17308);
nand U17922 (N_17922,N_16898,N_17268);
nor U17923 (N_17923,N_17348,N_17199);
and U17924 (N_17924,N_17005,N_16856);
nand U17925 (N_17925,N_17599,N_17323);
or U17926 (N_17926,N_17474,N_16803);
nand U17927 (N_17927,N_17176,N_16817);
xnor U17928 (N_17928,N_17065,N_17437);
nand U17929 (N_17929,N_16973,N_17229);
nand U17930 (N_17930,N_16989,N_17149);
and U17931 (N_17931,N_17292,N_17598);
nand U17932 (N_17932,N_17555,N_17398);
and U17933 (N_17933,N_17531,N_17498);
nand U17934 (N_17934,N_16862,N_17222);
xnor U17935 (N_17935,N_16925,N_16906);
xnor U17936 (N_17936,N_17364,N_17358);
nor U17937 (N_17937,N_17143,N_17144);
nor U17938 (N_17938,N_17047,N_17318);
nor U17939 (N_17939,N_17342,N_17442);
or U17940 (N_17940,N_17418,N_17001);
and U17941 (N_17941,N_17175,N_16971);
and U17942 (N_17942,N_17526,N_17484);
xor U17943 (N_17943,N_17123,N_16952);
nor U17944 (N_17944,N_17034,N_17524);
or U17945 (N_17945,N_16838,N_17026);
or U17946 (N_17946,N_17333,N_17537);
nand U17947 (N_17947,N_17295,N_17071);
nand U17948 (N_17948,N_17495,N_17002);
nand U17949 (N_17949,N_17375,N_16912);
nor U17950 (N_17950,N_16820,N_16849);
and U17951 (N_17951,N_17387,N_16866);
nand U17952 (N_17952,N_16826,N_17094);
or U17953 (N_17953,N_17594,N_16999);
nor U17954 (N_17954,N_16953,N_16833);
nor U17955 (N_17955,N_17548,N_17497);
nor U17956 (N_17956,N_16831,N_17114);
nand U17957 (N_17957,N_16810,N_17440);
or U17958 (N_17958,N_17024,N_17415);
or U17959 (N_17959,N_17481,N_16969);
nor U17960 (N_17960,N_16967,N_17392);
and U17961 (N_17961,N_17301,N_16867);
nand U17962 (N_17962,N_17404,N_17116);
or U17963 (N_17963,N_16933,N_16816);
xor U17964 (N_17964,N_17173,N_16913);
xnor U17965 (N_17965,N_16821,N_17304);
nand U17966 (N_17966,N_17550,N_17511);
xnor U17967 (N_17967,N_16855,N_16917);
nor U17968 (N_17968,N_17371,N_16930);
nand U17969 (N_17969,N_17075,N_17475);
or U17970 (N_17970,N_17234,N_16899);
xnor U17971 (N_17971,N_17330,N_17478);
or U17972 (N_17972,N_17403,N_17194);
or U17973 (N_17973,N_17117,N_17248);
nor U17974 (N_17974,N_17577,N_17529);
nand U17975 (N_17975,N_16970,N_16885);
xor U17976 (N_17976,N_17274,N_17151);
nand U17977 (N_17977,N_16956,N_17287);
nand U17978 (N_17978,N_17385,N_17110);
xor U17979 (N_17979,N_17040,N_17227);
xnor U17980 (N_17980,N_16823,N_17014);
or U17981 (N_17981,N_16980,N_17141);
or U17982 (N_17982,N_16939,N_17167);
or U17983 (N_17983,N_17541,N_17185);
xor U17984 (N_17984,N_17056,N_17502);
xnor U17985 (N_17985,N_17430,N_17035);
nor U17986 (N_17986,N_17320,N_17059);
nand U17987 (N_17987,N_17216,N_17338);
nor U17988 (N_17988,N_17426,N_16847);
or U17989 (N_17989,N_17543,N_16903);
nand U17990 (N_17990,N_17494,N_17240);
nand U17991 (N_17991,N_17121,N_17406);
or U17992 (N_17992,N_17305,N_17523);
or U17993 (N_17993,N_16893,N_17052);
xor U17994 (N_17994,N_17411,N_17125);
and U17995 (N_17995,N_17280,N_17314);
xor U17996 (N_17996,N_17290,N_17057);
or U17997 (N_17997,N_17188,N_17521);
or U17998 (N_17998,N_17208,N_16901);
and U17999 (N_17999,N_17373,N_17169);
xnor U18000 (N_18000,N_17487,N_17032);
nand U18001 (N_18001,N_17425,N_17313);
and U18002 (N_18002,N_17333,N_17099);
or U18003 (N_18003,N_17107,N_17437);
or U18004 (N_18004,N_17364,N_16920);
or U18005 (N_18005,N_16870,N_16948);
and U18006 (N_18006,N_16883,N_17297);
nor U18007 (N_18007,N_16868,N_17081);
nor U18008 (N_18008,N_17356,N_17298);
xor U18009 (N_18009,N_16909,N_17381);
and U18010 (N_18010,N_16894,N_17148);
nand U18011 (N_18011,N_17097,N_17338);
nor U18012 (N_18012,N_16854,N_16839);
xnor U18013 (N_18013,N_16864,N_17132);
xor U18014 (N_18014,N_17551,N_17116);
and U18015 (N_18015,N_17503,N_17498);
nor U18016 (N_18016,N_17261,N_17011);
nor U18017 (N_18017,N_17368,N_16867);
and U18018 (N_18018,N_17343,N_16826);
xor U18019 (N_18019,N_16827,N_17566);
nand U18020 (N_18020,N_16854,N_17305);
xnor U18021 (N_18021,N_16882,N_17267);
xor U18022 (N_18022,N_17036,N_17274);
xor U18023 (N_18023,N_17095,N_17270);
nor U18024 (N_18024,N_17335,N_17213);
xnor U18025 (N_18025,N_17422,N_16990);
or U18026 (N_18026,N_17021,N_17332);
nand U18027 (N_18027,N_17027,N_17231);
nor U18028 (N_18028,N_17110,N_16867);
nor U18029 (N_18029,N_17025,N_17352);
nor U18030 (N_18030,N_17154,N_16815);
nor U18031 (N_18031,N_17125,N_17177);
nand U18032 (N_18032,N_17585,N_17530);
or U18033 (N_18033,N_17135,N_16998);
nand U18034 (N_18034,N_16921,N_17308);
nor U18035 (N_18035,N_16813,N_17099);
and U18036 (N_18036,N_17058,N_17581);
nand U18037 (N_18037,N_17250,N_17527);
nor U18038 (N_18038,N_17126,N_17423);
xor U18039 (N_18039,N_17493,N_17241);
nand U18040 (N_18040,N_17120,N_17000);
or U18041 (N_18041,N_17158,N_17494);
nor U18042 (N_18042,N_16967,N_16850);
xor U18043 (N_18043,N_17066,N_17408);
and U18044 (N_18044,N_17484,N_17211);
and U18045 (N_18045,N_17147,N_17328);
nor U18046 (N_18046,N_17005,N_17328);
or U18047 (N_18047,N_17117,N_17280);
and U18048 (N_18048,N_17401,N_17447);
nor U18049 (N_18049,N_17259,N_16858);
nand U18050 (N_18050,N_17542,N_17499);
nor U18051 (N_18051,N_17047,N_17261);
or U18052 (N_18052,N_17196,N_17507);
and U18053 (N_18053,N_17425,N_17067);
xor U18054 (N_18054,N_17265,N_16969);
or U18055 (N_18055,N_17228,N_17570);
or U18056 (N_18056,N_17167,N_17232);
xor U18057 (N_18057,N_17229,N_17283);
and U18058 (N_18058,N_17263,N_16872);
nor U18059 (N_18059,N_17529,N_17524);
nor U18060 (N_18060,N_17509,N_17560);
or U18061 (N_18061,N_17123,N_17197);
or U18062 (N_18062,N_16808,N_16973);
nand U18063 (N_18063,N_17172,N_17260);
nand U18064 (N_18064,N_17251,N_16812);
and U18065 (N_18065,N_17242,N_17405);
nand U18066 (N_18066,N_17458,N_17089);
or U18067 (N_18067,N_17486,N_17118);
or U18068 (N_18068,N_16819,N_17566);
nor U18069 (N_18069,N_17161,N_16849);
nor U18070 (N_18070,N_17026,N_17295);
and U18071 (N_18071,N_17016,N_16970);
nand U18072 (N_18072,N_16920,N_17284);
and U18073 (N_18073,N_17191,N_17339);
nand U18074 (N_18074,N_17314,N_17083);
and U18075 (N_18075,N_17421,N_17130);
and U18076 (N_18076,N_16884,N_17384);
xor U18077 (N_18077,N_16894,N_17152);
xor U18078 (N_18078,N_17266,N_16919);
nor U18079 (N_18079,N_16898,N_16972);
or U18080 (N_18080,N_17259,N_16847);
and U18081 (N_18081,N_17301,N_17185);
or U18082 (N_18082,N_17425,N_17188);
and U18083 (N_18083,N_17210,N_17129);
xor U18084 (N_18084,N_17161,N_16861);
or U18085 (N_18085,N_17380,N_17525);
and U18086 (N_18086,N_16922,N_17054);
nand U18087 (N_18087,N_17528,N_17060);
or U18088 (N_18088,N_17317,N_16943);
nor U18089 (N_18089,N_17523,N_17063);
nor U18090 (N_18090,N_17302,N_17410);
xnor U18091 (N_18091,N_17542,N_16973);
nand U18092 (N_18092,N_17088,N_16910);
nor U18093 (N_18093,N_17106,N_17143);
nand U18094 (N_18094,N_17200,N_17347);
nor U18095 (N_18095,N_16939,N_16901);
nand U18096 (N_18096,N_17524,N_17129);
nor U18097 (N_18097,N_17100,N_17126);
nand U18098 (N_18098,N_16947,N_16813);
nand U18099 (N_18099,N_17121,N_17517);
or U18100 (N_18100,N_17358,N_17354);
nand U18101 (N_18101,N_17321,N_17015);
xor U18102 (N_18102,N_17352,N_17119);
xor U18103 (N_18103,N_16915,N_17427);
nor U18104 (N_18104,N_16806,N_17441);
or U18105 (N_18105,N_17049,N_16994);
and U18106 (N_18106,N_17554,N_17185);
nor U18107 (N_18107,N_16898,N_17459);
nor U18108 (N_18108,N_17398,N_16967);
or U18109 (N_18109,N_17285,N_17390);
or U18110 (N_18110,N_17064,N_17216);
and U18111 (N_18111,N_17497,N_17287);
nor U18112 (N_18112,N_16974,N_17410);
xnor U18113 (N_18113,N_17367,N_17542);
and U18114 (N_18114,N_17372,N_17042);
nor U18115 (N_18115,N_17177,N_17557);
nor U18116 (N_18116,N_17151,N_16874);
or U18117 (N_18117,N_17570,N_17229);
nor U18118 (N_18118,N_17084,N_17491);
xor U18119 (N_18119,N_16872,N_17142);
xor U18120 (N_18120,N_17051,N_17168);
and U18121 (N_18121,N_17489,N_17353);
nor U18122 (N_18122,N_17070,N_17224);
or U18123 (N_18123,N_17360,N_17385);
nand U18124 (N_18124,N_16825,N_17343);
and U18125 (N_18125,N_17526,N_17028);
nor U18126 (N_18126,N_17149,N_17199);
and U18127 (N_18127,N_16939,N_17439);
xor U18128 (N_18128,N_17452,N_17289);
and U18129 (N_18129,N_17270,N_16979);
or U18130 (N_18130,N_17577,N_16864);
and U18131 (N_18131,N_17380,N_17338);
nand U18132 (N_18132,N_17138,N_16898);
and U18133 (N_18133,N_17387,N_17383);
xor U18134 (N_18134,N_16879,N_17070);
nand U18135 (N_18135,N_16979,N_17176);
nor U18136 (N_18136,N_17491,N_17560);
xnor U18137 (N_18137,N_17169,N_17460);
or U18138 (N_18138,N_17479,N_17326);
or U18139 (N_18139,N_17487,N_16853);
and U18140 (N_18140,N_17034,N_17039);
nand U18141 (N_18141,N_17494,N_17322);
xnor U18142 (N_18142,N_16957,N_17168);
nor U18143 (N_18143,N_17587,N_16948);
or U18144 (N_18144,N_16814,N_16916);
or U18145 (N_18145,N_17495,N_17401);
nor U18146 (N_18146,N_17529,N_17597);
xor U18147 (N_18147,N_16870,N_17564);
and U18148 (N_18148,N_16971,N_17545);
xnor U18149 (N_18149,N_17492,N_17435);
xor U18150 (N_18150,N_17094,N_17401);
nor U18151 (N_18151,N_16821,N_17443);
nor U18152 (N_18152,N_17203,N_17044);
nor U18153 (N_18153,N_17458,N_17295);
nor U18154 (N_18154,N_17308,N_16805);
or U18155 (N_18155,N_17507,N_16995);
xor U18156 (N_18156,N_17374,N_17014);
or U18157 (N_18157,N_17078,N_17558);
and U18158 (N_18158,N_17152,N_17066);
or U18159 (N_18159,N_17174,N_17119);
nor U18160 (N_18160,N_17314,N_16813);
nand U18161 (N_18161,N_16887,N_17490);
nand U18162 (N_18162,N_17196,N_17593);
nand U18163 (N_18163,N_17276,N_17339);
or U18164 (N_18164,N_17405,N_17549);
nor U18165 (N_18165,N_17578,N_17133);
nand U18166 (N_18166,N_17228,N_17105);
and U18167 (N_18167,N_17319,N_17268);
xor U18168 (N_18168,N_17230,N_17244);
or U18169 (N_18169,N_17557,N_17153);
and U18170 (N_18170,N_16857,N_17373);
and U18171 (N_18171,N_16970,N_17429);
xnor U18172 (N_18172,N_17391,N_17577);
nor U18173 (N_18173,N_16843,N_16809);
nand U18174 (N_18174,N_17447,N_17287);
and U18175 (N_18175,N_17048,N_17270);
xor U18176 (N_18176,N_17009,N_17010);
nor U18177 (N_18177,N_16892,N_17212);
and U18178 (N_18178,N_17417,N_16827);
or U18179 (N_18179,N_17594,N_17322);
nand U18180 (N_18180,N_17491,N_17177);
or U18181 (N_18181,N_16982,N_16873);
and U18182 (N_18182,N_17191,N_17546);
nand U18183 (N_18183,N_17492,N_16883);
and U18184 (N_18184,N_16929,N_17115);
nand U18185 (N_18185,N_16886,N_17444);
xnor U18186 (N_18186,N_17592,N_17105);
nor U18187 (N_18187,N_17237,N_17059);
nand U18188 (N_18188,N_17455,N_17450);
and U18189 (N_18189,N_17563,N_17207);
nand U18190 (N_18190,N_17007,N_17413);
nand U18191 (N_18191,N_17476,N_16803);
nor U18192 (N_18192,N_17120,N_17266);
or U18193 (N_18193,N_16962,N_17377);
or U18194 (N_18194,N_17337,N_17420);
nand U18195 (N_18195,N_17194,N_17404);
nor U18196 (N_18196,N_17166,N_17280);
nor U18197 (N_18197,N_17443,N_16864);
nand U18198 (N_18198,N_17509,N_17106);
nor U18199 (N_18199,N_17598,N_17137);
xor U18200 (N_18200,N_16947,N_17384);
nor U18201 (N_18201,N_17207,N_17350);
nand U18202 (N_18202,N_16851,N_17078);
and U18203 (N_18203,N_17288,N_17555);
and U18204 (N_18204,N_17321,N_17354);
nor U18205 (N_18205,N_17020,N_16823);
and U18206 (N_18206,N_17192,N_16964);
xnor U18207 (N_18207,N_17033,N_16999);
and U18208 (N_18208,N_17483,N_17406);
and U18209 (N_18209,N_17248,N_17571);
xnor U18210 (N_18210,N_16831,N_17263);
and U18211 (N_18211,N_17502,N_17328);
or U18212 (N_18212,N_17356,N_17495);
nand U18213 (N_18213,N_17306,N_16997);
nor U18214 (N_18214,N_16821,N_16965);
and U18215 (N_18215,N_17506,N_16919);
xor U18216 (N_18216,N_16967,N_17541);
and U18217 (N_18217,N_17182,N_17562);
xnor U18218 (N_18218,N_17317,N_16856);
nor U18219 (N_18219,N_17435,N_17312);
nor U18220 (N_18220,N_17286,N_17306);
nand U18221 (N_18221,N_16850,N_17527);
nor U18222 (N_18222,N_17227,N_17216);
or U18223 (N_18223,N_17092,N_16954);
nor U18224 (N_18224,N_16827,N_17175);
or U18225 (N_18225,N_16994,N_16906);
xnor U18226 (N_18226,N_16912,N_16919);
or U18227 (N_18227,N_17152,N_16885);
nor U18228 (N_18228,N_17038,N_16993);
or U18229 (N_18229,N_17443,N_17456);
or U18230 (N_18230,N_17434,N_16861);
nand U18231 (N_18231,N_16990,N_17207);
nor U18232 (N_18232,N_17513,N_17176);
and U18233 (N_18233,N_16853,N_17152);
and U18234 (N_18234,N_17406,N_17430);
nor U18235 (N_18235,N_17168,N_17107);
nand U18236 (N_18236,N_17458,N_17432);
nor U18237 (N_18237,N_17054,N_17206);
xnor U18238 (N_18238,N_17166,N_17147);
or U18239 (N_18239,N_17537,N_17439);
nand U18240 (N_18240,N_17252,N_16940);
or U18241 (N_18241,N_17374,N_17144);
nand U18242 (N_18242,N_17193,N_16849);
or U18243 (N_18243,N_17024,N_16874);
and U18244 (N_18244,N_17330,N_17261);
or U18245 (N_18245,N_17500,N_16993);
xnor U18246 (N_18246,N_17342,N_17179);
or U18247 (N_18247,N_16997,N_17066);
nand U18248 (N_18248,N_17453,N_17316);
nor U18249 (N_18249,N_17067,N_16996);
xnor U18250 (N_18250,N_17289,N_17430);
nor U18251 (N_18251,N_16822,N_17492);
nand U18252 (N_18252,N_16953,N_17004);
and U18253 (N_18253,N_17119,N_17050);
xnor U18254 (N_18254,N_17302,N_16831);
nor U18255 (N_18255,N_17220,N_16884);
nand U18256 (N_18256,N_17089,N_17499);
and U18257 (N_18257,N_17369,N_17520);
xnor U18258 (N_18258,N_16962,N_17188);
or U18259 (N_18259,N_17066,N_17439);
and U18260 (N_18260,N_17268,N_16851);
and U18261 (N_18261,N_17153,N_17137);
nor U18262 (N_18262,N_17098,N_17273);
xor U18263 (N_18263,N_17446,N_16903);
nor U18264 (N_18264,N_17584,N_17240);
nand U18265 (N_18265,N_17593,N_17201);
nand U18266 (N_18266,N_17321,N_17569);
nor U18267 (N_18267,N_17389,N_16825);
or U18268 (N_18268,N_17098,N_17263);
and U18269 (N_18269,N_17523,N_17164);
nor U18270 (N_18270,N_17277,N_17334);
and U18271 (N_18271,N_17456,N_17488);
and U18272 (N_18272,N_17337,N_17153);
or U18273 (N_18273,N_17170,N_17406);
nand U18274 (N_18274,N_17056,N_17251);
or U18275 (N_18275,N_17290,N_17262);
or U18276 (N_18276,N_17307,N_17096);
nor U18277 (N_18277,N_17592,N_16829);
xor U18278 (N_18278,N_17589,N_17341);
and U18279 (N_18279,N_17314,N_16938);
and U18280 (N_18280,N_17540,N_17227);
nor U18281 (N_18281,N_17256,N_17469);
and U18282 (N_18282,N_16985,N_16860);
nand U18283 (N_18283,N_17396,N_17294);
nand U18284 (N_18284,N_17424,N_17155);
nor U18285 (N_18285,N_16921,N_17202);
nor U18286 (N_18286,N_17169,N_17398);
nand U18287 (N_18287,N_17258,N_17407);
nor U18288 (N_18288,N_17356,N_17303);
or U18289 (N_18289,N_17139,N_17263);
and U18290 (N_18290,N_16894,N_17578);
nor U18291 (N_18291,N_16881,N_17598);
and U18292 (N_18292,N_17095,N_17101);
xor U18293 (N_18293,N_16837,N_17467);
xnor U18294 (N_18294,N_17486,N_17169);
and U18295 (N_18295,N_17183,N_17431);
or U18296 (N_18296,N_16809,N_16913);
nor U18297 (N_18297,N_17186,N_17158);
xnor U18298 (N_18298,N_16804,N_16935);
xor U18299 (N_18299,N_17151,N_17404);
xnor U18300 (N_18300,N_17007,N_17412);
nor U18301 (N_18301,N_17110,N_17461);
xnor U18302 (N_18302,N_17543,N_16873);
nor U18303 (N_18303,N_17072,N_17218);
xor U18304 (N_18304,N_17038,N_17139);
nand U18305 (N_18305,N_17352,N_16910);
xnor U18306 (N_18306,N_17366,N_17409);
or U18307 (N_18307,N_16982,N_16979);
xor U18308 (N_18308,N_17092,N_17111);
or U18309 (N_18309,N_17050,N_17000);
and U18310 (N_18310,N_17254,N_17199);
and U18311 (N_18311,N_17246,N_17559);
nand U18312 (N_18312,N_17563,N_17094);
nor U18313 (N_18313,N_17307,N_17504);
or U18314 (N_18314,N_17044,N_16826);
or U18315 (N_18315,N_16927,N_17294);
nand U18316 (N_18316,N_17417,N_17205);
xnor U18317 (N_18317,N_17241,N_17414);
nand U18318 (N_18318,N_17332,N_17315);
xnor U18319 (N_18319,N_17458,N_17408);
nand U18320 (N_18320,N_16903,N_16998);
nor U18321 (N_18321,N_17172,N_16827);
and U18322 (N_18322,N_17223,N_17318);
xnor U18323 (N_18323,N_17205,N_17342);
nand U18324 (N_18324,N_16819,N_16902);
nor U18325 (N_18325,N_17376,N_16975);
nor U18326 (N_18326,N_16816,N_17203);
and U18327 (N_18327,N_17448,N_17230);
or U18328 (N_18328,N_17057,N_16840);
xor U18329 (N_18329,N_17381,N_16958);
nor U18330 (N_18330,N_17488,N_16882);
xor U18331 (N_18331,N_17417,N_17474);
or U18332 (N_18332,N_17475,N_17426);
nor U18333 (N_18333,N_16998,N_16973);
nand U18334 (N_18334,N_16964,N_17203);
or U18335 (N_18335,N_17391,N_17354);
and U18336 (N_18336,N_16906,N_17392);
nor U18337 (N_18337,N_17462,N_17094);
nand U18338 (N_18338,N_16885,N_16889);
or U18339 (N_18339,N_17292,N_17448);
xor U18340 (N_18340,N_16938,N_16878);
nand U18341 (N_18341,N_17183,N_16814);
xnor U18342 (N_18342,N_16850,N_17339);
or U18343 (N_18343,N_16891,N_16970);
and U18344 (N_18344,N_17293,N_17339);
nor U18345 (N_18345,N_16865,N_17378);
or U18346 (N_18346,N_16977,N_17076);
nand U18347 (N_18347,N_17440,N_17002);
and U18348 (N_18348,N_17134,N_16844);
or U18349 (N_18349,N_17069,N_17429);
xnor U18350 (N_18350,N_17441,N_16904);
and U18351 (N_18351,N_17486,N_17313);
or U18352 (N_18352,N_17094,N_17297);
xnor U18353 (N_18353,N_17154,N_17476);
xor U18354 (N_18354,N_17475,N_16847);
nor U18355 (N_18355,N_16949,N_16877);
nor U18356 (N_18356,N_17063,N_17554);
xor U18357 (N_18357,N_16923,N_17245);
nand U18358 (N_18358,N_17255,N_17097);
and U18359 (N_18359,N_17195,N_17295);
xor U18360 (N_18360,N_17246,N_17315);
nand U18361 (N_18361,N_17159,N_17573);
and U18362 (N_18362,N_16951,N_17423);
or U18363 (N_18363,N_17541,N_17126);
or U18364 (N_18364,N_16990,N_17200);
and U18365 (N_18365,N_17596,N_17118);
xor U18366 (N_18366,N_17006,N_17140);
and U18367 (N_18367,N_16808,N_17396);
nor U18368 (N_18368,N_17353,N_16882);
xnor U18369 (N_18369,N_17303,N_17549);
or U18370 (N_18370,N_17544,N_17234);
or U18371 (N_18371,N_17445,N_17141);
nand U18372 (N_18372,N_17184,N_17236);
or U18373 (N_18373,N_16894,N_16915);
xor U18374 (N_18374,N_17176,N_17287);
or U18375 (N_18375,N_17111,N_17028);
nor U18376 (N_18376,N_17009,N_17058);
and U18377 (N_18377,N_17166,N_17238);
nor U18378 (N_18378,N_17000,N_16958);
and U18379 (N_18379,N_16914,N_17330);
xor U18380 (N_18380,N_17352,N_17180);
nor U18381 (N_18381,N_16831,N_17153);
and U18382 (N_18382,N_17368,N_17508);
or U18383 (N_18383,N_17535,N_17467);
or U18384 (N_18384,N_17226,N_17403);
and U18385 (N_18385,N_16923,N_16833);
or U18386 (N_18386,N_17417,N_17595);
or U18387 (N_18387,N_17168,N_16952);
and U18388 (N_18388,N_17299,N_16856);
or U18389 (N_18389,N_17428,N_17088);
or U18390 (N_18390,N_16835,N_17586);
nor U18391 (N_18391,N_17340,N_17443);
or U18392 (N_18392,N_17374,N_17213);
nor U18393 (N_18393,N_17441,N_17122);
nand U18394 (N_18394,N_17456,N_17584);
xnor U18395 (N_18395,N_17233,N_17508);
or U18396 (N_18396,N_16858,N_17578);
nor U18397 (N_18397,N_17592,N_17374);
nand U18398 (N_18398,N_17521,N_16983);
nand U18399 (N_18399,N_17346,N_17485);
and U18400 (N_18400,N_17946,N_17840);
xnor U18401 (N_18401,N_17770,N_18200);
or U18402 (N_18402,N_17646,N_18132);
and U18403 (N_18403,N_18316,N_17959);
nor U18404 (N_18404,N_17615,N_18210);
and U18405 (N_18405,N_17967,N_17939);
nor U18406 (N_18406,N_17837,N_18113);
or U18407 (N_18407,N_18269,N_18130);
nor U18408 (N_18408,N_17645,N_18299);
and U18409 (N_18409,N_18103,N_18123);
nor U18410 (N_18410,N_18312,N_17714);
nor U18411 (N_18411,N_18260,N_18191);
nor U18412 (N_18412,N_17659,N_18195);
or U18413 (N_18413,N_18389,N_17920);
xor U18414 (N_18414,N_18071,N_18031);
nor U18415 (N_18415,N_18270,N_18214);
and U18416 (N_18416,N_17649,N_18151);
nand U18417 (N_18417,N_17652,N_17816);
and U18418 (N_18418,N_17826,N_18285);
nor U18419 (N_18419,N_18057,N_17685);
and U18420 (N_18420,N_18093,N_18266);
and U18421 (N_18421,N_17728,N_17688);
and U18422 (N_18422,N_17634,N_18264);
xnor U18423 (N_18423,N_18334,N_18176);
or U18424 (N_18424,N_18361,N_17830);
nor U18425 (N_18425,N_17867,N_17934);
nor U18426 (N_18426,N_17968,N_17705);
or U18427 (N_18427,N_18115,N_18314);
xor U18428 (N_18428,N_17846,N_18188);
or U18429 (N_18429,N_17948,N_17774);
and U18430 (N_18430,N_18090,N_18294);
nor U18431 (N_18431,N_18075,N_18338);
nor U18432 (N_18432,N_17859,N_18356);
xnor U18433 (N_18433,N_17924,N_18366);
or U18434 (N_18434,N_17881,N_18351);
or U18435 (N_18435,N_17760,N_17677);
nand U18436 (N_18436,N_18136,N_18142);
and U18437 (N_18437,N_17779,N_18359);
nand U18438 (N_18438,N_17813,N_18357);
and U18439 (N_18439,N_17608,N_18078);
nor U18440 (N_18440,N_18282,N_18331);
or U18441 (N_18441,N_18126,N_17710);
and U18442 (N_18442,N_17702,N_18379);
nor U18443 (N_18443,N_18313,N_17869);
xnor U18444 (N_18444,N_17777,N_18208);
xor U18445 (N_18445,N_17928,N_18001);
and U18446 (N_18446,N_18028,N_18398);
or U18447 (N_18447,N_18372,N_17986);
or U18448 (N_18448,N_17616,N_17641);
or U18449 (N_18449,N_18102,N_18112);
or U18450 (N_18450,N_17648,N_18088);
and U18451 (N_18451,N_17684,N_17681);
or U18452 (N_18452,N_17970,N_17619);
or U18453 (N_18453,N_18399,N_17925);
or U18454 (N_18454,N_17804,N_17895);
or U18455 (N_18455,N_18207,N_18201);
nand U18456 (N_18456,N_17679,N_17889);
xor U18457 (N_18457,N_18107,N_17734);
or U18458 (N_18458,N_18169,N_17696);
nor U18459 (N_18459,N_18301,N_17611);
nand U18460 (N_18460,N_18383,N_18375);
or U18461 (N_18461,N_17871,N_18307);
and U18462 (N_18462,N_18240,N_17656);
and U18463 (N_18463,N_17717,N_18165);
and U18464 (N_18464,N_17772,N_18012);
or U18465 (N_18465,N_18013,N_17942);
and U18466 (N_18466,N_17692,N_17806);
and U18467 (N_18467,N_17730,N_17627);
or U18468 (N_18468,N_17757,N_17839);
and U18469 (N_18469,N_18295,N_18309);
or U18470 (N_18470,N_17762,N_17899);
nor U18471 (N_18471,N_18009,N_17953);
or U18472 (N_18472,N_17686,N_17810);
or U18473 (N_18473,N_18087,N_18127);
and U18474 (N_18474,N_17628,N_18129);
nor U18475 (N_18475,N_18277,N_18327);
nor U18476 (N_18476,N_18058,N_17817);
nand U18477 (N_18477,N_17820,N_17625);
and U18478 (N_18478,N_18175,N_17747);
nor U18479 (N_18479,N_18106,N_17614);
or U18480 (N_18480,N_17680,N_18336);
nor U18481 (N_18481,N_18304,N_18074);
and U18482 (N_18482,N_18043,N_17910);
xor U18483 (N_18483,N_17778,N_18380);
and U18484 (N_18484,N_17745,N_18373);
nor U18485 (N_18485,N_17907,N_17913);
or U18486 (N_18486,N_18382,N_18180);
or U18487 (N_18487,N_17700,N_18154);
or U18488 (N_18488,N_18155,N_17694);
and U18489 (N_18489,N_17850,N_18344);
or U18490 (N_18490,N_18203,N_18051);
xnor U18491 (N_18491,N_18086,N_17971);
nand U18492 (N_18492,N_18147,N_18163);
xnor U18493 (N_18493,N_18026,N_18273);
nor U18494 (N_18494,N_17888,N_18350);
and U18495 (N_18495,N_18215,N_17610);
xor U18496 (N_18496,N_17812,N_17731);
xor U18497 (N_18497,N_18118,N_17626);
nand U18498 (N_18498,N_17936,N_17974);
nand U18499 (N_18499,N_18092,N_17632);
xnor U18500 (N_18500,N_18381,N_17849);
nor U18501 (N_18501,N_18385,N_17739);
xnor U18502 (N_18502,N_18306,N_17941);
nand U18503 (N_18503,N_18072,N_17987);
xor U18504 (N_18504,N_18183,N_18164);
or U18505 (N_18505,N_18248,N_17997);
nor U18506 (N_18506,N_18021,N_18292);
nand U18507 (N_18507,N_17665,N_18345);
nand U18508 (N_18508,N_17638,N_17769);
nor U18509 (N_18509,N_18326,N_17961);
or U18510 (N_18510,N_17896,N_17980);
nor U18511 (N_18511,N_18333,N_17780);
nand U18512 (N_18512,N_18288,N_17995);
nand U18513 (N_18513,N_17944,N_17744);
nand U18514 (N_18514,N_17723,N_18287);
nor U18515 (N_18515,N_17984,N_17751);
xor U18516 (N_18516,N_17624,N_18347);
or U18517 (N_18517,N_17786,N_18048);
or U18518 (N_18518,N_17722,N_17758);
nand U18519 (N_18519,N_17797,N_18190);
or U18520 (N_18520,N_17977,N_18014);
or U18521 (N_18521,N_18003,N_18000);
or U18522 (N_18522,N_18109,N_18241);
xnor U18523 (N_18523,N_17658,N_17719);
xnor U18524 (N_18524,N_17919,N_18230);
and U18525 (N_18525,N_17799,N_17622);
or U18526 (N_18526,N_18308,N_18284);
xor U18527 (N_18527,N_18140,N_18302);
xnor U18528 (N_18528,N_18197,N_18050);
and U18529 (N_18529,N_18049,N_17633);
or U18530 (N_18530,N_17922,N_18089);
xnor U18531 (N_18531,N_17711,N_17651);
and U18532 (N_18532,N_17636,N_17932);
and U18533 (N_18533,N_18388,N_18256);
nand U18534 (N_18534,N_18186,N_17732);
and U18535 (N_18535,N_17661,N_18289);
and U18536 (N_18536,N_18038,N_18220);
xor U18537 (N_18537,N_18394,N_18293);
and U18538 (N_18538,N_17976,N_17654);
or U18539 (N_18539,N_17706,N_18077);
xnor U18540 (N_18540,N_18348,N_17943);
nand U18541 (N_18541,N_17918,N_17955);
nor U18542 (N_18542,N_18393,N_17882);
or U18543 (N_18543,N_18070,N_18296);
and U18544 (N_18544,N_18276,N_18252);
and U18545 (N_18545,N_18173,N_18167);
xor U18546 (N_18546,N_18387,N_18137);
xor U18547 (N_18547,N_18213,N_17873);
xor U18548 (N_18548,N_17958,N_18303);
and U18549 (N_18549,N_18209,N_17855);
and U18550 (N_18550,N_17668,N_17682);
or U18551 (N_18551,N_18337,N_17891);
xor U18552 (N_18552,N_18119,N_17742);
nor U18553 (N_18553,N_17979,N_17950);
or U18554 (N_18554,N_17897,N_17653);
nor U18555 (N_18555,N_18390,N_17848);
and U18556 (N_18556,N_17911,N_18145);
nor U18557 (N_18557,N_18365,N_17704);
nand U18558 (N_18558,N_18233,N_18286);
xnor U18559 (N_18559,N_17885,N_18039);
nand U18560 (N_18560,N_17727,N_17814);
and U18561 (N_18561,N_17858,N_18291);
or U18562 (N_18562,N_17715,N_17767);
or U18563 (N_18563,N_18108,N_18310);
nand U18564 (N_18564,N_18105,N_17612);
nor U18565 (N_18565,N_17992,N_18073);
nor U18566 (N_18566,N_18221,N_18297);
nor U18567 (N_18567,N_17975,N_17879);
xor U18568 (N_18568,N_18300,N_18275);
and U18569 (N_18569,N_18280,N_18247);
and U18570 (N_18570,N_18272,N_18152);
nand U18571 (N_18571,N_17993,N_18219);
and U18572 (N_18572,N_18052,N_17945);
or U18573 (N_18573,N_17916,N_18358);
nand U18574 (N_18574,N_18224,N_17667);
and U18575 (N_18575,N_17740,N_18133);
nor U18576 (N_18576,N_17738,N_17713);
xor U18577 (N_18577,N_18011,N_18143);
and U18578 (N_18578,N_18114,N_17796);
nand U18579 (N_18579,N_18332,N_18234);
xnor U18580 (N_18580,N_17834,N_18060);
and U18581 (N_18581,N_18352,N_18202);
xnor U18582 (N_18582,N_18042,N_17629);
nand U18583 (N_18583,N_18135,N_18251);
nor U18584 (N_18584,N_18311,N_18010);
or U18585 (N_18585,N_18037,N_17785);
or U18586 (N_18586,N_17947,N_18063);
xor U18587 (N_18587,N_18198,N_17712);
nor U18588 (N_18588,N_18218,N_17908);
nor U18589 (N_18589,N_17662,N_18329);
or U18590 (N_18590,N_18053,N_17841);
nor U18591 (N_18591,N_18149,N_17673);
xnor U18592 (N_18592,N_17736,N_17784);
or U18593 (N_18593,N_18177,N_17793);
nand U18594 (N_18594,N_18259,N_17860);
nor U18595 (N_18595,N_18392,N_17726);
and U18596 (N_18596,N_17802,N_18024);
nand U18597 (N_18597,N_18305,N_18020);
xnor U18598 (N_18598,N_17672,N_17824);
nor U18599 (N_18599,N_18315,N_18171);
nor U18600 (N_18600,N_17909,N_18255);
or U18601 (N_18601,N_17821,N_18232);
and U18602 (N_18602,N_18267,N_17754);
and U18603 (N_18603,N_18015,N_18298);
or U18604 (N_18604,N_17866,N_17852);
xor U18605 (N_18605,N_17914,N_17842);
xnor U18606 (N_18606,N_17605,N_17695);
xor U18607 (N_18607,N_17683,N_18189);
xor U18608 (N_18608,N_18002,N_17725);
and U18609 (N_18609,N_18341,N_17701);
xnor U18610 (N_18610,N_17776,N_17838);
nor U18611 (N_18611,N_17966,N_18146);
nand U18612 (N_18612,N_17666,N_18018);
or U18613 (N_18613,N_17602,N_17829);
or U18614 (N_18614,N_18085,N_18322);
nor U18615 (N_18615,N_18239,N_17721);
nor U18616 (N_18616,N_18150,N_18355);
or U18617 (N_18617,N_17905,N_18159);
and U18618 (N_18618,N_17828,N_18033);
nor U18619 (N_18619,N_18076,N_18371);
nand U18620 (N_18620,N_18228,N_18242);
and U18621 (N_18621,N_18320,N_18179);
nor U18622 (N_18622,N_18317,N_18004);
nand U18623 (N_18623,N_18116,N_18323);
and U18624 (N_18624,N_17601,N_18254);
nor U18625 (N_18625,N_18216,N_18046);
nor U18626 (N_18626,N_18091,N_18244);
xor U18627 (N_18627,N_18279,N_17874);
and U18628 (N_18628,N_18229,N_17900);
xnor U18629 (N_18629,N_17833,N_17775);
and U18630 (N_18630,N_17815,N_18170);
xnor U18631 (N_18631,N_18066,N_18141);
or U18632 (N_18632,N_17861,N_17854);
xnor U18633 (N_18633,N_18378,N_18231);
xor U18634 (N_18634,N_17748,N_17631);
and U18635 (N_18635,N_18121,N_18391);
nand U18636 (N_18636,N_18364,N_18369);
nor U18637 (N_18637,N_17781,N_18206);
and U18638 (N_18638,N_18153,N_18237);
xor U18639 (N_18639,N_17844,N_18061);
xnor U18640 (N_18640,N_18040,N_17877);
and U18641 (N_18641,N_18339,N_17892);
nor U18642 (N_18642,N_18016,N_18395);
nand U18643 (N_18643,N_18027,N_18217);
nand U18644 (N_18644,N_17825,N_17956);
nand U18645 (N_18645,N_17808,N_17604);
and U18646 (N_18646,N_18022,N_18253);
nor U18647 (N_18647,N_17724,N_18257);
or U18648 (N_18648,N_17880,N_17978);
nor U18649 (N_18649,N_18187,N_17707);
or U18650 (N_18650,N_17752,N_18168);
nor U18651 (N_18651,N_17674,N_18098);
or U18652 (N_18652,N_17782,N_18328);
or U18653 (N_18653,N_17960,N_18367);
xnor U18654 (N_18654,N_17853,N_17836);
xnor U18655 (N_18655,N_18174,N_18128);
nand U18656 (N_18656,N_17949,N_17963);
nand U18657 (N_18657,N_17832,N_17801);
or U18658 (N_18658,N_17693,N_18156);
nor U18659 (N_18659,N_18342,N_17964);
xnor U18660 (N_18660,N_18261,N_17994);
nor U18661 (N_18661,N_18268,N_17893);
or U18662 (N_18662,N_18099,N_18065);
nand U18663 (N_18663,N_17663,N_17735);
or U18664 (N_18664,N_18377,N_17898);
or U18665 (N_18665,N_17639,N_18192);
nand U18666 (N_18666,N_17635,N_18181);
and U18667 (N_18667,N_18222,N_17805);
nand U18668 (N_18668,N_18321,N_18030);
nor U18669 (N_18669,N_18249,N_17720);
nor U18670 (N_18670,N_18184,N_17856);
nor U18671 (N_18671,N_17988,N_17937);
nand U18672 (N_18672,N_18250,N_17794);
or U18673 (N_18673,N_17951,N_17894);
nand U18674 (N_18674,N_17903,N_17613);
or U18675 (N_18675,N_17765,N_18059);
xnor U18676 (N_18676,N_17687,N_17904);
xnor U18677 (N_18677,N_17851,N_18212);
nor U18678 (N_18678,N_18335,N_18162);
or U18679 (N_18679,N_18111,N_17931);
and U18680 (N_18680,N_17708,N_17835);
xor U18681 (N_18681,N_17827,N_18110);
or U18682 (N_18682,N_17862,N_17886);
and U18683 (N_18683,N_18124,N_17737);
xor U18684 (N_18684,N_18082,N_18069);
or U18685 (N_18685,N_18097,N_17809);
and U18686 (N_18686,N_18161,N_17965);
and U18687 (N_18687,N_17981,N_17691);
nand U18688 (N_18688,N_18023,N_17999);
and U18689 (N_18689,N_18083,N_18067);
nor U18690 (N_18690,N_17643,N_17985);
or U18691 (N_18691,N_17972,N_18226);
xor U18692 (N_18692,N_17753,N_18258);
or U18693 (N_18693,N_18283,N_18199);
nand U18694 (N_18694,N_17831,N_18263);
nand U18695 (N_18695,N_18343,N_17697);
nand U18696 (N_18696,N_17716,N_17623);
and U18697 (N_18697,N_17845,N_17800);
xnor U18698 (N_18698,N_17878,N_18144);
or U18699 (N_18699,N_18196,N_17771);
nand U18700 (N_18700,N_18035,N_17803);
and U18701 (N_18701,N_17930,N_18349);
or U18702 (N_18702,N_18397,N_17609);
and U18703 (N_18703,N_17990,N_18243);
and U18704 (N_18704,N_18054,N_18084);
or U18705 (N_18705,N_17933,N_18120);
nor U18706 (N_18706,N_17669,N_18318);
and U18707 (N_18707,N_17620,N_17675);
or U18708 (N_18708,N_18148,N_18225);
nand U18709 (N_18709,N_17890,N_17872);
nor U18710 (N_18710,N_18125,N_17921);
and U18711 (N_18711,N_17901,N_18006);
nand U18712 (N_18712,N_17883,N_17923);
nor U18713 (N_18713,N_18062,N_18117);
or U18714 (N_18714,N_18265,N_18368);
nor U18715 (N_18715,N_17822,N_17690);
xnor U18716 (N_18716,N_17991,N_18081);
nand U18717 (N_18717,N_17902,N_17733);
xnor U18718 (N_18718,N_18353,N_18235);
nor U18719 (N_18719,N_18138,N_18360);
nand U18720 (N_18720,N_18172,N_17759);
or U18721 (N_18721,N_18278,N_17863);
or U18722 (N_18722,N_17670,N_18019);
or U18723 (N_18723,N_17741,N_18036);
or U18724 (N_18724,N_18182,N_18017);
and U18725 (N_18725,N_18271,N_17671);
xor U18726 (N_18726,N_17768,N_18056);
nand U18727 (N_18727,N_18122,N_18047);
nor U18728 (N_18728,N_17969,N_17887);
and U18729 (N_18729,N_17600,N_18274);
nor U18730 (N_18730,N_17660,N_17790);
nor U18731 (N_18731,N_18384,N_17819);
or U18732 (N_18732,N_18374,N_17621);
or U18733 (N_18733,N_17847,N_18095);
nand U18734 (N_18734,N_17935,N_18363);
and U18735 (N_18735,N_18205,N_18104);
nand U18736 (N_18736,N_18005,N_17929);
nor U18737 (N_18737,N_18025,N_17698);
nand U18738 (N_18738,N_17843,N_18236);
xnor U18739 (N_18739,N_18100,N_17749);
nand U18740 (N_18740,N_18370,N_17915);
nand U18741 (N_18741,N_18041,N_18376);
and U18742 (N_18742,N_18068,N_17655);
nand U18743 (N_18743,N_17743,N_18166);
nor U18744 (N_18744,N_17865,N_17761);
nor U18745 (N_18745,N_17607,N_17630);
or U18746 (N_18746,N_17689,N_17764);
or U18747 (N_18747,N_17998,N_18045);
xor U18748 (N_18748,N_18246,N_17795);
nor U18749 (N_18749,N_17783,N_17983);
or U18750 (N_18750,N_18079,N_17617);
or U18751 (N_18751,N_17938,N_17906);
xnor U18752 (N_18752,N_17811,N_17750);
and U18753 (N_18753,N_17940,N_17746);
nor U18754 (N_18754,N_17884,N_18096);
and U18755 (N_18755,N_17703,N_18290);
or U18756 (N_18756,N_18194,N_17644);
nand U18757 (N_18757,N_18055,N_18185);
xnor U18758 (N_18758,N_18080,N_18094);
nand U18759 (N_18759,N_17798,N_17876);
nand U18760 (N_18760,N_17709,N_17756);
and U18761 (N_18761,N_17766,N_18245);
and U18762 (N_18762,N_18101,N_17864);
nor U18763 (N_18763,N_17642,N_17926);
nand U18764 (N_18764,N_18325,N_17868);
nand U18765 (N_18765,N_17870,N_17807);
nor U18766 (N_18766,N_17773,N_18007);
and U18767 (N_18767,N_18044,N_18281);
nand U18768 (N_18768,N_18362,N_18193);
and U18769 (N_18769,N_17927,N_17647);
nor U18770 (N_18770,N_17664,N_18238);
nor U18771 (N_18771,N_18034,N_18330);
xor U18772 (N_18772,N_18178,N_17954);
xnor U18773 (N_18773,N_18223,N_17763);
xor U18774 (N_18774,N_17755,N_18211);
and U18775 (N_18775,N_18157,N_17912);
nand U18776 (N_18776,N_18396,N_18134);
xor U18777 (N_18777,N_18227,N_18008);
and U18778 (N_18778,N_17699,N_17678);
nand U18779 (N_18779,N_17982,N_17640);
xor U18780 (N_18780,N_17788,N_17637);
xnor U18781 (N_18781,N_18386,N_17917);
and U18782 (N_18782,N_18158,N_17818);
or U18783 (N_18783,N_18204,N_18032);
xnor U18784 (N_18784,N_17787,N_18160);
nor U18785 (N_18785,N_17973,N_18064);
and U18786 (N_18786,N_17650,N_17792);
and U18787 (N_18787,N_18354,N_18346);
xor U18788 (N_18788,N_17857,N_17823);
and U18789 (N_18789,N_17657,N_18319);
and U18790 (N_18790,N_17875,N_18340);
and U18791 (N_18791,N_18324,N_17603);
xor U18792 (N_18792,N_18131,N_17789);
nor U18793 (N_18793,N_18262,N_17676);
xnor U18794 (N_18794,N_18139,N_17989);
or U18795 (N_18795,N_17962,N_17996);
nor U18796 (N_18796,N_17718,N_17606);
xor U18797 (N_18797,N_17729,N_17957);
and U18798 (N_18798,N_17791,N_17952);
nor U18799 (N_18799,N_18029,N_17618);
and U18800 (N_18800,N_18138,N_17778);
and U18801 (N_18801,N_17952,N_18044);
nor U18802 (N_18802,N_17813,N_18082);
nand U18803 (N_18803,N_17847,N_18276);
nor U18804 (N_18804,N_18299,N_18394);
and U18805 (N_18805,N_17720,N_17896);
nand U18806 (N_18806,N_18206,N_17826);
nand U18807 (N_18807,N_18075,N_18238);
and U18808 (N_18808,N_18086,N_17610);
xor U18809 (N_18809,N_18299,N_17855);
and U18810 (N_18810,N_17878,N_18040);
and U18811 (N_18811,N_18041,N_18354);
xnor U18812 (N_18812,N_17931,N_18191);
nand U18813 (N_18813,N_17657,N_17834);
and U18814 (N_18814,N_18212,N_18065);
nor U18815 (N_18815,N_18333,N_18141);
xor U18816 (N_18816,N_17916,N_17915);
xnor U18817 (N_18817,N_18221,N_17836);
or U18818 (N_18818,N_18138,N_17645);
nand U18819 (N_18819,N_17612,N_17703);
xnor U18820 (N_18820,N_18296,N_17918);
and U18821 (N_18821,N_18010,N_18354);
nand U18822 (N_18822,N_17732,N_17974);
nand U18823 (N_18823,N_17836,N_17740);
nor U18824 (N_18824,N_18262,N_17688);
and U18825 (N_18825,N_18196,N_17975);
xor U18826 (N_18826,N_17733,N_17947);
and U18827 (N_18827,N_17631,N_17615);
nor U18828 (N_18828,N_18009,N_17755);
nand U18829 (N_18829,N_17719,N_17698);
nor U18830 (N_18830,N_17775,N_17614);
and U18831 (N_18831,N_17619,N_18192);
and U18832 (N_18832,N_17984,N_18136);
or U18833 (N_18833,N_17787,N_17621);
nand U18834 (N_18834,N_18028,N_18323);
and U18835 (N_18835,N_18203,N_17984);
or U18836 (N_18836,N_17612,N_17915);
or U18837 (N_18837,N_18105,N_17819);
nor U18838 (N_18838,N_18330,N_18035);
nor U18839 (N_18839,N_18003,N_17808);
nor U18840 (N_18840,N_17781,N_18020);
xor U18841 (N_18841,N_18051,N_17934);
and U18842 (N_18842,N_18145,N_18275);
and U18843 (N_18843,N_17949,N_18198);
or U18844 (N_18844,N_17738,N_18382);
nand U18845 (N_18845,N_17651,N_17956);
nor U18846 (N_18846,N_17684,N_17844);
xnor U18847 (N_18847,N_18005,N_17696);
xor U18848 (N_18848,N_17896,N_17983);
nor U18849 (N_18849,N_17904,N_18167);
or U18850 (N_18850,N_17730,N_18274);
nor U18851 (N_18851,N_17860,N_18005);
nand U18852 (N_18852,N_18271,N_17973);
xor U18853 (N_18853,N_18246,N_18098);
and U18854 (N_18854,N_17866,N_18183);
and U18855 (N_18855,N_18355,N_18210);
nand U18856 (N_18856,N_18142,N_18389);
nor U18857 (N_18857,N_18388,N_18009);
xor U18858 (N_18858,N_18130,N_17873);
xor U18859 (N_18859,N_18124,N_17833);
nor U18860 (N_18860,N_17820,N_18130);
and U18861 (N_18861,N_17884,N_17605);
nor U18862 (N_18862,N_17812,N_18324);
or U18863 (N_18863,N_18123,N_18111);
nor U18864 (N_18864,N_17734,N_18218);
or U18865 (N_18865,N_18069,N_18084);
or U18866 (N_18866,N_17648,N_18254);
xor U18867 (N_18867,N_17970,N_18206);
or U18868 (N_18868,N_18050,N_17971);
nand U18869 (N_18869,N_18371,N_18288);
and U18870 (N_18870,N_17674,N_18216);
nor U18871 (N_18871,N_17922,N_18076);
xor U18872 (N_18872,N_17978,N_18382);
or U18873 (N_18873,N_18221,N_17904);
xnor U18874 (N_18874,N_18343,N_18251);
xnor U18875 (N_18875,N_18281,N_18126);
xor U18876 (N_18876,N_18089,N_18270);
nor U18877 (N_18877,N_17790,N_18037);
xnor U18878 (N_18878,N_18335,N_18258);
nand U18879 (N_18879,N_17989,N_17719);
nand U18880 (N_18880,N_18005,N_17872);
and U18881 (N_18881,N_18053,N_18249);
xor U18882 (N_18882,N_17936,N_18392);
nor U18883 (N_18883,N_18068,N_17605);
nor U18884 (N_18884,N_17833,N_18117);
nand U18885 (N_18885,N_17618,N_18150);
nand U18886 (N_18886,N_17639,N_18343);
xnor U18887 (N_18887,N_18226,N_17906);
nand U18888 (N_18888,N_18383,N_17935);
xnor U18889 (N_18889,N_18319,N_17683);
and U18890 (N_18890,N_18382,N_17778);
and U18891 (N_18891,N_17862,N_17933);
nand U18892 (N_18892,N_18365,N_18368);
and U18893 (N_18893,N_17792,N_18317);
nor U18894 (N_18894,N_18251,N_17724);
nor U18895 (N_18895,N_17863,N_17621);
or U18896 (N_18896,N_17690,N_18022);
xor U18897 (N_18897,N_18244,N_18240);
or U18898 (N_18898,N_18378,N_17761);
and U18899 (N_18899,N_18224,N_17834);
nor U18900 (N_18900,N_17871,N_18134);
nand U18901 (N_18901,N_18181,N_17966);
or U18902 (N_18902,N_18071,N_17780);
and U18903 (N_18903,N_17656,N_18164);
xor U18904 (N_18904,N_18341,N_18269);
and U18905 (N_18905,N_17795,N_17745);
and U18906 (N_18906,N_18318,N_18039);
and U18907 (N_18907,N_18131,N_17695);
or U18908 (N_18908,N_18363,N_17686);
xnor U18909 (N_18909,N_18343,N_17694);
nand U18910 (N_18910,N_18390,N_17763);
nor U18911 (N_18911,N_18337,N_17961);
or U18912 (N_18912,N_18289,N_18180);
or U18913 (N_18913,N_17956,N_17983);
nor U18914 (N_18914,N_18094,N_18067);
or U18915 (N_18915,N_17726,N_18315);
and U18916 (N_18916,N_18257,N_18244);
nor U18917 (N_18917,N_17893,N_18103);
and U18918 (N_18918,N_18388,N_18139);
and U18919 (N_18919,N_17679,N_17969);
nor U18920 (N_18920,N_18168,N_17681);
nand U18921 (N_18921,N_17961,N_17906);
or U18922 (N_18922,N_17689,N_18044);
or U18923 (N_18923,N_18202,N_17696);
or U18924 (N_18924,N_17926,N_17872);
nand U18925 (N_18925,N_18172,N_17965);
nor U18926 (N_18926,N_18196,N_17677);
and U18927 (N_18927,N_18185,N_18012);
and U18928 (N_18928,N_18286,N_18023);
nor U18929 (N_18929,N_17944,N_18229);
nor U18930 (N_18930,N_17680,N_18016);
or U18931 (N_18931,N_18269,N_18196);
nor U18932 (N_18932,N_18298,N_18258);
or U18933 (N_18933,N_18211,N_17900);
and U18934 (N_18934,N_18183,N_18390);
nand U18935 (N_18935,N_18393,N_18379);
nand U18936 (N_18936,N_17631,N_18319);
nor U18937 (N_18937,N_17995,N_18253);
nor U18938 (N_18938,N_18266,N_17682);
nor U18939 (N_18939,N_18210,N_17950);
or U18940 (N_18940,N_18083,N_17971);
and U18941 (N_18941,N_18092,N_18101);
nor U18942 (N_18942,N_18054,N_18396);
xnor U18943 (N_18943,N_18174,N_18366);
xor U18944 (N_18944,N_17978,N_17802);
and U18945 (N_18945,N_18227,N_17970);
and U18946 (N_18946,N_18201,N_17748);
and U18947 (N_18947,N_18151,N_17658);
or U18948 (N_18948,N_17821,N_17886);
nand U18949 (N_18949,N_17828,N_18309);
or U18950 (N_18950,N_17860,N_17629);
nor U18951 (N_18951,N_18140,N_18161);
or U18952 (N_18952,N_17860,N_17673);
and U18953 (N_18953,N_17609,N_17650);
xnor U18954 (N_18954,N_17825,N_17629);
xnor U18955 (N_18955,N_18202,N_17616);
nor U18956 (N_18956,N_18294,N_18065);
xor U18957 (N_18957,N_18196,N_17958);
nor U18958 (N_18958,N_17992,N_18290);
and U18959 (N_18959,N_17833,N_18331);
nand U18960 (N_18960,N_18011,N_17873);
and U18961 (N_18961,N_18208,N_18274);
xnor U18962 (N_18962,N_17740,N_17718);
nor U18963 (N_18963,N_17982,N_17905);
nor U18964 (N_18964,N_17922,N_18110);
xor U18965 (N_18965,N_17974,N_18175);
xor U18966 (N_18966,N_17629,N_17849);
or U18967 (N_18967,N_18197,N_18054);
and U18968 (N_18968,N_17789,N_18152);
or U18969 (N_18969,N_18315,N_17645);
xnor U18970 (N_18970,N_17604,N_18372);
xor U18971 (N_18971,N_17948,N_17900);
nand U18972 (N_18972,N_17981,N_17704);
nor U18973 (N_18973,N_17675,N_17773);
xnor U18974 (N_18974,N_18255,N_17986);
or U18975 (N_18975,N_17775,N_18326);
and U18976 (N_18976,N_17841,N_17859);
or U18977 (N_18977,N_18360,N_17885);
xnor U18978 (N_18978,N_18399,N_17879);
or U18979 (N_18979,N_17907,N_18002);
nor U18980 (N_18980,N_18010,N_18245);
or U18981 (N_18981,N_18064,N_17934);
nor U18982 (N_18982,N_17870,N_17885);
nor U18983 (N_18983,N_17935,N_17814);
or U18984 (N_18984,N_18369,N_17686);
nand U18985 (N_18985,N_17664,N_17792);
xor U18986 (N_18986,N_17600,N_17824);
xnor U18987 (N_18987,N_17755,N_17725);
nand U18988 (N_18988,N_17667,N_18009);
nand U18989 (N_18989,N_17935,N_17745);
or U18990 (N_18990,N_18084,N_18266);
nand U18991 (N_18991,N_17756,N_17808);
nand U18992 (N_18992,N_17930,N_18272);
nor U18993 (N_18993,N_17749,N_18349);
xor U18994 (N_18994,N_17699,N_17700);
or U18995 (N_18995,N_18091,N_17756);
and U18996 (N_18996,N_17682,N_17686);
nand U18997 (N_18997,N_17863,N_17789);
and U18998 (N_18998,N_18261,N_18232);
nor U18999 (N_18999,N_18010,N_17830);
nor U19000 (N_19000,N_17881,N_17618);
nand U19001 (N_19001,N_17608,N_17919);
xor U19002 (N_19002,N_18187,N_17601);
and U19003 (N_19003,N_18106,N_17762);
nand U19004 (N_19004,N_18297,N_18128);
nand U19005 (N_19005,N_18371,N_17603);
nor U19006 (N_19006,N_17813,N_17600);
nand U19007 (N_19007,N_18110,N_18014);
xor U19008 (N_19008,N_18365,N_18197);
nand U19009 (N_19009,N_18377,N_18142);
or U19010 (N_19010,N_18081,N_18083);
nand U19011 (N_19011,N_17745,N_17838);
nor U19012 (N_19012,N_17608,N_17949);
nand U19013 (N_19013,N_18006,N_17845);
or U19014 (N_19014,N_17905,N_18378);
or U19015 (N_19015,N_17654,N_18057);
nand U19016 (N_19016,N_17605,N_17911);
nand U19017 (N_19017,N_17959,N_18182);
xor U19018 (N_19018,N_17645,N_17683);
and U19019 (N_19019,N_18045,N_18392);
or U19020 (N_19020,N_18163,N_18363);
nor U19021 (N_19021,N_17875,N_17723);
and U19022 (N_19022,N_18364,N_18233);
xor U19023 (N_19023,N_18312,N_17694);
or U19024 (N_19024,N_17999,N_18321);
or U19025 (N_19025,N_17847,N_17614);
xnor U19026 (N_19026,N_18394,N_17719);
nor U19027 (N_19027,N_18215,N_18290);
or U19028 (N_19028,N_17783,N_18183);
or U19029 (N_19029,N_17679,N_18067);
xor U19030 (N_19030,N_17976,N_17851);
xor U19031 (N_19031,N_17749,N_17638);
nand U19032 (N_19032,N_17632,N_17768);
xnor U19033 (N_19033,N_17968,N_17664);
nand U19034 (N_19034,N_18205,N_18348);
nand U19035 (N_19035,N_18178,N_17625);
and U19036 (N_19036,N_17926,N_17958);
or U19037 (N_19037,N_18135,N_17804);
and U19038 (N_19038,N_18049,N_17732);
nand U19039 (N_19039,N_17702,N_17957);
and U19040 (N_19040,N_17977,N_18185);
or U19041 (N_19041,N_17818,N_17766);
nand U19042 (N_19042,N_18329,N_17819);
or U19043 (N_19043,N_18062,N_17999);
and U19044 (N_19044,N_17859,N_17799);
xor U19045 (N_19045,N_18182,N_17923);
xnor U19046 (N_19046,N_17664,N_18024);
nand U19047 (N_19047,N_18325,N_18185);
nand U19048 (N_19048,N_17856,N_17949);
xnor U19049 (N_19049,N_17900,N_17683);
nor U19050 (N_19050,N_18298,N_17922);
nand U19051 (N_19051,N_17823,N_18361);
or U19052 (N_19052,N_18222,N_17900);
nor U19053 (N_19053,N_18062,N_17675);
nor U19054 (N_19054,N_17783,N_18155);
nor U19055 (N_19055,N_18121,N_18252);
nand U19056 (N_19056,N_17818,N_18340);
nor U19057 (N_19057,N_18087,N_18339);
nand U19058 (N_19058,N_18376,N_18046);
and U19059 (N_19059,N_17681,N_18067);
nand U19060 (N_19060,N_17957,N_18350);
or U19061 (N_19061,N_18197,N_17962);
and U19062 (N_19062,N_18297,N_18080);
nand U19063 (N_19063,N_18129,N_18173);
or U19064 (N_19064,N_17886,N_17853);
and U19065 (N_19065,N_17931,N_18140);
xor U19066 (N_19066,N_18269,N_18004);
xor U19067 (N_19067,N_18351,N_18232);
or U19068 (N_19068,N_18268,N_17812);
xor U19069 (N_19069,N_17603,N_18143);
or U19070 (N_19070,N_18133,N_17997);
xor U19071 (N_19071,N_17871,N_17643);
or U19072 (N_19072,N_18213,N_17887);
xor U19073 (N_19073,N_18148,N_18365);
nor U19074 (N_19074,N_17936,N_18395);
xor U19075 (N_19075,N_18105,N_18233);
xnor U19076 (N_19076,N_17641,N_17605);
nand U19077 (N_19077,N_18138,N_17795);
or U19078 (N_19078,N_17614,N_17960);
nor U19079 (N_19079,N_17952,N_17637);
and U19080 (N_19080,N_18290,N_18386);
xnor U19081 (N_19081,N_17763,N_17911);
nand U19082 (N_19082,N_18143,N_18336);
nor U19083 (N_19083,N_18372,N_18068);
nand U19084 (N_19084,N_18223,N_18216);
or U19085 (N_19085,N_18399,N_17924);
nor U19086 (N_19086,N_17849,N_17782);
nand U19087 (N_19087,N_18252,N_17766);
or U19088 (N_19088,N_18139,N_17725);
and U19089 (N_19089,N_17939,N_18162);
or U19090 (N_19090,N_17835,N_17855);
or U19091 (N_19091,N_18271,N_17652);
and U19092 (N_19092,N_18207,N_17895);
and U19093 (N_19093,N_18015,N_17706);
nand U19094 (N_19094,N_18262,N_17605);
or U19095 (N_19095,N_18261,N_18212);
or U19096 (N_19096,N_18357,N_18367);
nand U19097 (N_19097,N_17948,N_18147);
nand U19098 (N_19098,N_17901,N_18222);
nand U19099 (N_19099,N_18157,N_17798);
nor U19100 (N_19100,N_18241,N_18224);
nor U19101 (N_19101,N_18258,N_18267);
nor U19102 (N_19102,N_17968,N_17884);
nor U19103 (N_19103,N_18178,N_17743);
or U19104 (N_19104,N_17983,N_18337);
nor U19105 (N_19105,N_18358,N_17829);
nand U19106 (N_19106,N_17679,N_18096);
nor U19107 (N_19107,N_17665,N_18099);
nor U19108 (N_19108,N_18167,N_17983);
xnor U19109 (N_19109,N_17687,N_17772);
or U19110 (N_19110,N_18020,N_17926);
or U19111 (N_19111,N_18324,N_18155);
nand U19112 (N_19112,N_18379,N_18359);
nand U19113 (N_19113,N_17786,N_17604);
and U19114 (N_19114,N_17743,N_18001);
nand U19115 (N_19115,N_18140,N_18205);
nand U19116 (N_19116,N_18340,N_18226);
nand U19117 (N_19117,N_18304,N_18081);
nor U19118 (N_19118,N_17616,N_18080);
and U19119 (N_19119,N_17702,N_18217);
or U19120 (N_19120,N_18118,N_18006);
nor U19121 (N_19121,N_17852,N_17674);
xor U19122 (N_19122,N_18064,N_17953);
and U19123 (N_19123,N_18264,N_18253);
xor U19124 (N_19124,N_18218,N_18185);
and U19125 (N_19125,N_18303,N_18365);
nor U19126 (N_19126,N_17992,N_17612);
nor U19127 (N_19127,N_18382,N_17765);
nand U19128 (N_19128,N_18194,N_18368);
nor U19129 (N_19129,N_18127,N_17884);
or U19130 (N_19130,N_17964,N_18077);
nor U19131 (N_19131,N_18362,N_18038);
xnor U19132 (N_19132,N_18169,N_18261);
nand U19133 (N_19133,N_18306,N_17760);
nand U19134 (N_19134,N_18394,N_17825);
nor U19135 (N_19135,N_18330,N_18308);
or U19136 (N_19136,N_17915,N_17973);
and U19137 (N_19137,N_17638,N_17741);
xnor U19138 (N_19138,N_17777,N_18314);
or U19139 (N_19139,N_17637,N_17941);
xnor U19140 (N_19140,N_17717,N_17635);
xnor U19141 (N_19141,N_17819,N_18036);
or U19142 (N_19142,N_18148,N_17997);
and U19143 (N_19143,N_17763,N_17631);
and U19144 (N_19144,N_17864,N_18197);
or U19145 (N_19145,N_18136,N_17703);
xnor U19146 (N_19146,N_17622,N_17962);
and U19147 (N_19147,N_18228,N_17969);
nor U19148 (N_19148,N_17892,N_18115);
nand U19149 (N_19149,N_17892,N_18310);
xnor U19150 (N_19150,N_17647,N_17960);
xnor U19151 (N_19151,N_17835,N_17941);
or U19152 (N_19152,N_18164,N_17905);
and U19153 (N_19153,N_18056,N_17787);
nor U19154 (N_19154,N_18218,N_18112);
xor U19155 (N_19155,N_17960,N_17915);
nor U19156 (N_19156,N_17840,N_17940);
and U19157 (N_19157,N_17895,N_18123);
or U19158 (N_19158,N_18009,N_17669);
and U19159 (N_19159,N_18341,N_18119);
and U19160 (N_19160,N_18193,N_18258);
or U19161 (N_19161,N_17895,N_18010);
nor U19162 (N_19162,N_17710,N_18238);
xor U19163 (N_19163,N_17737,N_17883);
nor U19164 (N_19164,N_17793,N_17818);
nor U19165 (N_19165,N_18205,N_17939);
or U19166 (N_19166,N_18276,N_18270);
xor U19167 (N_19167,N_17946,N_18091);
nor U19168 (N_19168,N_17862,N_17793);
nand U19169 (N_19169,N_18184,N_17677);
nor U19170 (N_19170,N_17686,N_17653);
and U19171 (N_19171,N_18239,N_17998);
xnor U19172 (N_19172,N_18352,N_18079);
or U19173 (N_19173,N_18367,N_18101);
and U19174 (N_19174,N_18119,N_18115);
nor U19175 (N_19175,N_18152,N_17865);
or U19176 (N_19176,N_18239,N_18338);
or U19177 (N_19177,N_18245,N_18180);
and U19178 (N_19178,N_17841,N_18119);
or U19179 (N_19179,N_18295,N_18142);
nand U19180 (N_19180,N_18146,N_17736);
and U19181 (N_19181,N_18265,N_17983);
and U19182 (N_19182,N_17619,N_17677);
nand U19183 (N_19183,N_17621,N_17927);
nand U19184 (N_19184,N_17729,N_18077);
and U19185 (N_19185,N_18256,N_17734);
nand U19186 (N_19186,N_17730,N_18343);
and U19187 (N_19187,N_18067,N_18240);
nor U19188 (N_19188,N_18062,N_18203);
or U19189 (N_19189,N_17810,N_17728);
xor U19190 (N_19190,N_18359,N_17715);
xor U19191 (N_19191,N_18340,N_17657);
xor U19192 (N_19192,N_18139,N_18313);
or U19193 (N_19193,N_17858,N_18005);
xor U19194 (N_19194,N_18326,N_17790);
and U19195 (N_19195,N_18063,N_18099);
nand U19196 (N_19196,N_18263,N_18308);
xor U19197 (N_19197,N_18141,N_17812);
and U19198 (N_19198,N_18024,N_17806);
or U19199 (N_19199,N_17879,N_17716);
or U19200 (N_19200,N_18763,N_18924);
or U19201 (N_19201,N_18582,N_18693);
nor U19202 (N_19202,N_18847,N_18903);
xor U19203 (N_19203,N_19071,N_18932);
and U19204 (N_19204,N_18865,N_19054);
xor U19205 (N_19205,N_18635,N_18850);
and U19206 (N_19206,N_18420,N_18674);
xor U19207 (N_19207,N_18422,N_18836);
xor U19208 (N_19208,N_19097,N_18948);
or U19209 (N_19209,N_19057,N_18411);
or U19210 (N_19210,N_19168,N_18942);
or U19211 (N_19211,N_19144,N_18528);
nand U19212 (N_19212,N_18658,N_19034);
or U19213 (N_19213,N_18487,N_19065);
xor U19214 (N_19214,N_18559,N_18637);
nand U19215 (N_19215,N_18401,N_18634);
nor U19216 (N_19216,N_18825,N_19199);
or U19217 (N_19217,N_19187,N_18921);
or U19218 (N_19218,N_18426,N_18553);
nor U19219 (N_19219,N_19102,N_18897);
nand U19220 (N_19220,N_19149,N_19181);
or U19221 (N_19221,N_18834,N_18419);
nand U19222 (N_19222,N_18476,N_19021);
nand U19223 (N_19223,N_18887,N_18937);
or U19224 (N_19224,N_18703,N_19083);
nand U19225 (N_19225,N_18599,N_18681);
and U19226 (N_19226,N_18661,N_18782);
nor U19227 (N_19227,N_18550,N_18931);
and U19228 (N_19228,N_19018,N_18460);
nand U19229 (N_19229,N_18985,N_18779);
nand U19230 (N_19230,N_18767,N_18575);
or U19231 (N_19231,N_18520,N_18452);
nor U19232 (N_19232,N_18955,N_18702);
nor U19233 (N_19233,N_19066,N_19177);
or U19234 (N_19234,N_18894,N_18527);
and U19235 (N_19235,N_19082,N_19027);
nor U19236 (N_19236,N_18480,N_18765);
and U19237 (N_19237,N_19129,N_18477);
and U19238 (N_19238,N_19009,N_18730);
nand U19239 (N_19239,N_18977,N_18900);
or U19240 (N_19240,N_18745,N_18835);
nor U19241 (N_19241,N_19006,N_18416);
nor U19242 (N_19242,N_18882,N_18901);
and U19243 (N_19243,N_18868,N_18874);
nand U19244 (N_19244,N_18475,N_19108);
and U19245 (N_19245,N_19158,N_18594);
xor U19246 (N_19246,N_18579,N_19157);
xor U19247 (N_19247,N_18572,N_18859);
nor U19248 (N_19248,N_18498,N_19182);
nand U19249 (N_19249,N_18772,N_18538);
xnor U19250 (N_19250,N_18562,N_18896);
xnor U19251 (N_19251,N_18983,N_18967);
or U19252 (N_19252,N_18766,N_18666);
nor U19253 (N_19253,N_18543,N_18727);
or U19254 (N_19254,N_19039,N_18953);
or U19255 (N_19255,N_18536,N_18642);
and U19256 (N_19256,N_18628,N_18793);
or U19257 (N_19257,N_19164,N_18971);
nor U19258 (N_19258,N_18406,N_18534);
and U19259 (N_19259,N_18610,N_18537);
xnor U19260 (N_19260,N_18884,N_18996);
or U19261 (N_19261,N_18928,N_19038);
nand U19262 (N_19262,N_18925,N_18524);
and U19263 (N_19263,N_18851,N_18690);
xor U19264 (N_19264,N_19002,N_18731);
nor U19265 (N_19265,N_18907,N_18962);
or U19266 (N_19266,N_18551,N_18555);
nor U19267 (N_19267,N_18784,N_18866);
nand U19268 (N_19268,N_18984,N_19194);
or U19269 (N_19269,N_18875,N_18747);
xnor U19270 (N_19270,N_18603,N_18873);
or U19271 (N_19271,N_18697,N_18744);
nor U19272 (N_19272,N_18604,N_18783);
and U19273 (N_19273,N_18624,N_18467);
and U19274 (N_19274,N_18516,N_18799);
and U19275 (N_19275,N_19025,N_18876);
nand U19276 (N_19276,N_18701,N_18620);
nor U19277 (N_19277,N_18933,N_18877);
and U19278 (N_19278,N_19089,N_18789);
or U19279 (N_19279,N_19030,N_18811);
and U19280 (N_19280,N_18507,N_19175);
and U19281 (N_19281,N_18795,N_18732);
and U19282 (N_19282,N_18770,N_19188);
and U19283 (N_19283,N_19036,N_18807);
nor U19284 (N_19284,N_19074,N_19167);
nand U19285 (N_19285,N_19063,N_18797);
or U19286 (N_19286,N_19058,N_18404);
or U19287 (N_19287,N_18991,N_18899);
xnor U19288 (N_19288,N_18539,N_19145);
nor U19289 (N_19289,N_18695,N_19107);
xnor U19290 (N_19290,N_18472,N_18429);
nor U19291 (N_19291,N_18918,N_19026);
nand U19292 (N_19292,N_18490,N_18653);
and U19293 (N_19293,N_18801,N_18706);
nand U19294 (N_19294,N_18934,N_18821);
and U19295 (N_19295,N_18717,N_18410);
xor U19296 (N_19296,N_18437,N_19046);
or U19297 (N_19297,N_18454,N_19010);
and U19298 (N_19298,N_19163,N_19121);
and U19299 (N_19299,N_18427,N_18966);
xnor U19300 (N_19300,N_19007,N_18776);
xnor U19301 (N_19301,N_18643,N_18492);
xor U19302 (N_19302,N_19067,N_18616);
and U19303 (N_19303,N_18905,N_18692);
xor U19304 (N_19304,N_18682,N_19091);
nand U19305 (N_19305,N_18584,N_18707);
or U19306 (N_19306,N_18812,N_19012);
nand U19307 (N_19307,N_18672,N_18407);
nand U19308 (N_19308,N_18623,N_18506);
nor U19309 (N_19309,N_19170,N_18418);
nor U19310 (N_19310,N_19048,N_18423);
xor U19311 (N_19311,N_18483,N_19062);
xor U19312 (N_19312,N_18968,N_19195);
xnor U19313 (N_19313,N_18842,N_18758);
or U19314 (N_19314,N_18961,N_19041);
xor U19315 (N_19315,N_18815,N_18833);
xor U19316 (N_19316,N_18400,N_19073);
nand U19317 (N_19317,N_18940,N_18714);
or U19318 (N_19318,N_19176,N_18614);
and U19319 (N_19319,N_18529,N_19172);
or U19320 (N_19320,N_18872,N_18880);
nor U19321 (N_19321,N_19135,N_18436);
nand U19322 (N_19322,N_19161,N_18949);
or U19323 (N_19323,N_18606,N_18951);
xor U19324 (N_19324,N_19136,N_19100);
xor U19325 (N_19325,N_19120,N_19092);
nand U19326 (N_19326,N_18451,N_18558);
and U19327 (N_19327,N_18626,N_18891);
nand U19328 (N_19328,N_18699,N_18595);
xnor U19329 (N_19329,N_18790,N_18573);
nor U19330 (N_19330,N_18839,N_18540);
nor U19331 (N_19331,N_18561,N_19037);
nor U19332 (N_19332,N_18916,N_19109);
xor U19333 (N_19333,N_18669,N_18496);
nor U19334 (N_19334,N_19053,N_18771);
and U19335 (N_19335,N_18627,N_19116);
nor U19336 (N_19336,N_18456,N_19070);
xor U19337 (N_19337,N_18578,N_19189);
or U19338 (N_19338,N_18974,N_18522);
and U19339 (N_19339,N_18554,N_18638);
nor U19340 (N_19340,N_18650,N_18945);
nor U19341 (N_19341,N_19019,N_19094);
and U19342 (N_19342,N_19140,N_18781);
xor U19343 (N_19343,N_18863,N_18656);
xnor U19344 (N_19344,N_19130,N_18752);
nand U19345 (N_19345,N_18412,N_18530);
xnor U19346 (N_19346,N_18959,N_18587);
nor U19347 (N_19347,N_18816,N_18533);
nand U19348 (N_19348,N_18769,N_18568);
and U19349 (N_19349,N_18618,N_18890);
or U19350 (N_19350,N_18660,N_18640);
nor U19351 (N_19351,N_18719,N_19064);
xnor U19352 (N_19352,N_19069,N_19015);
and U19353 (N_19353,N_19031,N_18557);
and U19354 (N_19354,N_19183,N_18929);
xnor U19355 (N_19355,N_18946,N_19079);
or U19356 (N_19356,N_18999,N_18408);
nand U19357 (N_19357,N_19084,N_19127);
and U19358 (N_19358,N_18488,N_18489);
nor U19359 (N_19359,N_18691,N_18957);
and U19360 (N_19360,N_18560,N_19098);
nor U19361 (N_19361,N_18685,N_18440);
and U19362 (N_19362,N_18800,N_18739);
nand U19363 (N_19363,N_19191,N_18670);
nand U19364 (N_19364,N_19081,N_18886);
or U19365 (N_19365,N_18756,N_18421);
xnor U19366 (N_19366,N_19190,N_19016);
xor U19367 (N_19367,N_18556,N_18671);
nor U19368 (N_19368,N_18935,N_18808);
nor U19369 (N_19369,N_19128,N_18822);
and U19370 (N_19370,N_18910,N_18917);
nand U19371 (N_19371,N_18571,N_18485);
and U19372 (N_19372,N_18950,N_18827);
and U19373 (N_19373,N_18857,N_18545);
nand U19374 (N_19374,N_18619,N_18810);
xor U19375 (N_19375,N_19068,N_18523);
nand U19376 (N_19376,N_18519,N_18469);
and U19377 (N_19377,N_19143,N_18673);
nor U19378 (N_19378,N_18775,N_18424);
nor U19379 (N_19379,N_19060,N_19117);
or U19380 (N_19380,N_18631,N_18878);
nand U19381 (N_19381,N_18952,N_18831);
and U19382 (N_19382,N_19011,N_18652);
nor U19383 (N_19383,N_18570,N_19196);
xnor U19384 (N_19384,N_18823,N_18751);
nor U19385 (N_19385,N_18405,N_19008);
nor U19386 (N_19386,N_18546,N_18592);
xnor U19387 (N_19387,N_18838,N_19033);
or U19388 (N_19388,N_19134,N_18486);
nor U19389 (N_19389,N_18657,N_18438);
nor U19390 (N_19390,N_19138,N_18497);
and U19391 (N_19391,N_18860,N_19162);
or U19392 (N_19392,N_19141,N_19197);
nand U19393 (N_19393,N_18773,N_18668);
or U19394 (N_19394,N_18402,N_18885);
xor U19395 (N_19395,N_19169,N_18694);
nand U19396 (N_19396,N_19159,N_18446);
or U19397 (N_19397,N_19111,N_19137);
nor U19398 (N_19398,N_18893,N_18943);
nand U19399 (N_19399,N_18755,N_19131);
nand U19400 (N_19400,N_18700,N_18826);
or U19401 (N_19401,N_18915,N_18647);
or U19402 (N_19402,N_19080,N_18787);
xnor U19403 (N_19403,N_18923,N_18960);
and U19404 (N_19404,N_18774,N_18721);
nor U19405 (N_19405,N_18414,N_18531);
and U19406 (N_19406,N_18500,N_18636);
xnor U19407 (N_19407,N_18457,N_18740);
xnor U19408 (N_19408,N_19184,N_18493);
xor U19409 (N_19409,N_19017,N_19032);
and U19410 (N_19410,N_18566,N_18780);
and U19411 (N_19411,N_19051,N_18442);
or U19412 (N_19412,N_19014,N_18499);
nor U19413 (N_19413,N_18802,N_19024);
xnor U19414 (N_19414,N_18818,N_18710);
xor U19415 (N_19415,N_18549,N_18908);
nand U19416 (N_19416,N_18728,N_18646);
nand U19417 (N_19417,N_18686,N_18704);
xor U19418 (N_19418,N_18501,N_18805);
nor U19419 (N_19419,N_18806,N_19088);
nor U19420 (N_19420,N_18513,N_19192);
xnor U19421 (N_19421,N_19166,N_18723);
xnor U19422 (N_19422,N_19052,N_18517);
nor U19423 (N_19423,N_18509,N_18849);
xor U19424 (N_19424,N_18995,N_18510);
or U19425 (N_19425,N_18435,N_19152);
and U19426 (N_19426,N_19044,N_18982);
nor U19427 (N_19427,N_19104,N_18737);
nor U19428 (N_19428,N_18845,N_18969);
xor U19429 (N_19429,N_19122,N_18632);
and U19430 (N_19430,N_18978,N_18864);
nor U19431 (N_19431,N_18667,N_18430);
and U19432 (N_19432,N_19118,N_18432);
or U19433 (N_19433,N_18963,N_18904);
or U19434 (N_19434,N_19179,N_18709);
and U19435 (N_19435,N_18439,N_18854);
and U19436 (N_19436,N_18824,N_18503);
xnor U19437 (N_19437,N_19099,N_18830);
and U19438 (N_19438,N_18413,N_19173);
xnor U19439 (N_19439,N_18846,N_18941);
xor U19440 (N_19440,N_18589,N_18871);
and U19441 (N_19441,N_18986,N_18518);
nor U19442 (N_19442,N_18746,N_18742);
or U19443 (N_19443,N_18841,N_18581);
or U19444 (N_19444,N_18683,N_18803);
or U19445 (N_19445,N_18708,N_18852);
nand U19446 (N_19446,N_19093,N_19154);
or U19447 (N_19447,N_19075,N_18663);
and U19448 (N_19448,N_18768,N_18869);
nor U19449 (N_19449,N_18761,N_18688);
nand U19450 (N_19450,N_18757,N_18712);
nand U19451 (N_19451,N_19174,N_18753);
and U19452 (N_19452,N_18856,N_18526);
nand U19453 (N_19453,N_19101,N_19119);
nor U19454 (N_19454,N_18881,N_18630);
nand U19455 (N_19455,N_19139,N_18861);
or U19456 (N_19456,N_19035,N_18569);
and U19457 (N_19457,N_18724,N_19055);
xor U19458 (N_19458,N_18615,N_18645);
or U19459 (N_19459,N_18461,N_18463);
and U19460 (N_19460,N_19077,N_19126);
or U19461 (N_19461,N_18919,N_18920);
and U19462 (N_19462,N_19153,N_18639);
nor U19463 (N_19463,N_18759,N_19056);
and U19464 (N_19464,N_19023,N_18633);
xor U19465 (N_19465,N_18936,N_18468);
xor U19466 (N_19466,N_18725,N_18458);
nor U19467 (N_19467,N_18926,N_18544);
or U19468 (N_19468,N_18798,N_18649);
or U19469 (N_19469,N_18711,N_19147);
or U19470 (N_19470,N_18804,N_18947);
nand U19471 (N_19471,N_19020,N_18607);
or U19472 (N_19472,N_18895,N_18979);
nor U19473 (N_19473,N_18590,N_19198);
or U19474 (N_19474,N_18902,N_18591);
xor U19475 (N_19475,N_18409,N_18445);
nand U19476 (N_19476,N_18862,N_19043);
nand U19477 (N_19477,N_18892,N_18809);
and U19478 (N_19478,N_18525,N_18720);
nand U19479 (N_19479,N_18867,N_18914);
or U19480 (N_19480,N_18611,N_19180);
and U19481 (N_19481,N_18598,N_18898);
or U19482 (N_19482,N_18705,N_18840);
xor U19483 (N_19483,N_18883,N_19003);
xnor U19484 (N_19484,N_18738,N_18450);
nand U19485 (N_19485,N_18567,N_19047);
and U19486 (N_19486,N_18814,N_19156);
xor U19487 (N_19487,N_18735,N_18478);
xnor U19488 (N_19488,N_18855,N_18444);
and U19489 (N_19489,N_19132,N_18989);
and U19490 (N_19490,N_19133,N_19105);
or U19491 (N_19491,N_18588,N_18481);
nor U19492 (N_19492,N_18532,N_18586);
and U19493 (N_19493,N_18482,N_18617);
and U19494 (N_19494,N_19113,N_18684);
or U19495 (N_19495,N_18625,N_18448);
and U19496 (N_19496,N_18484,N_19090);
nor U19497 (N_19497,N_19150,N_19001);
or U19498 (N_19498,N_18565,N_18583);
and U19499 (N_19499,N_18813,N_19045);
xnor U19500 (N_19500,N_18913,N_18596);
or U19501 (N_19501,N_18718,N_19114);
nor U19502 (N_19502,N_18508,N_19186);
nor U19503 (N_19503,N_18754,N_18741);
and U19504 (N_19504,N_19124,N_19013);
or U19505 (N_19505,N_18664,N_18428);
nand U19506 (N_19506,N_19096,N_18972);
and U19507 (N_19507,N_18796,N_18729);
xor U19508 (N_19508,N_18687,N_18655);
and U19509 (N_19509,N_18675,N_18612);
nor U19510 (N_19510,N_18749,N_18858);
xnor U19511 (N_19511,N_18563,N_18662);
and U19512 (N_19512,N_18734,N_18791);
or U19513 (N_19513,N_19123,N_18786);
nor U19514 (N_19514,N_18552,N_19072);
nor U19515 (N_19515,N_19112,N_18988);
and U19516 (N_19516,N_18843,N_18785);
and U19517 (N_19517,N_18512,N_18479);
and U19518 (N_19518,N_18449,N_19103);
and U19519 (N_19519,N_18879,N_18605);
or U19520 (N_19520,N_18608,N_18515);
xnor U19521 (N_19521,N_18777,N_19005);
xnor U19522 (N_19522,N_18521,N_18998);
nor U19523 (N_19523,N_18629,N_18930);
or U19524 (N_19524,N_18609,N_18980);
nand U19525 (N_19525,N_18542,N_19165);
nor U19526 (N_19526,N_18722,N_18441);
and U19527 (N_19527,N_18778,N_18621);
or U19528 (N_19528,N_18679,N_18853);
xnor U19529 (N_19529,N_19029,N_18689);
or U19530 (N_19530,N_18415,N_19155);
xnor U19531 (N_19531,N_18641,N_18944);
xor U19532 (N_19532,N_18970,N_18547);
or U19533 (N_19533,N_19040,N_18504);
nor U19534 (N_19534,N_18748,N_19049);
and U19535 (N_19535,N_18535,N_18992);
nand U19536 (N_19536,N_18993,N_19148);
or U19537 (N_19537,N_18987,N_18462);
nor U19538 (N_19538,N_19193,N_18927);
xnor U19539 (N_19539,N_18580,N_18473);
or U19540 (N_19540,N_18403,N_18911);
nor U19541 (N_19541,N_18597,N_18654);
and U19542 (N_19542,N_18848,N_18417);
xor U19543 (N_19543,N_18495,N_18514);
nand U19544 (N_19544,N_18466,N_18651);
nand U19545 (N_19545,N_18677,N_18443);
or U19546 (N_19546,N_18494,N_19004);
nand U19547 (N_19547,N_18794,N_18820);
and U19548 (N_19548,N_18976,N_19059);
nor U19549 (N_19549,N_18909,N_19110);
nand U19550 (N_19550,N_18593,N_19185);
nor U19551 (N_19551,N_18792,N_18760);
nor U19552 (N_19552,N_18888,N_19115);
and U19553 (N_19553,N_18958,N_19000);
nand U19554 (N_19554,N_18505,N_18828);
and U19555 (N_19555,N_19085,N_18447);
xnor U19556 (N_19556,N_19087,N_19061);
xor U19557 (N_19557,N_18600,N_19151);
and U19558 (N_19558,N_18938,N_18470);
and U19559 (N_19559,N_18453,N_18602);
and U19560 (N_19560,N_19125,N_19178);
and U19561 (N_19561,N_18680,N_19171);
and U19562 (N_19562,N_18648,N_18817);
nor U19563 (N_19563,N_18990,N_18574);
nand U19564 (N_19564,N_18511,N_18678);
nand U19565 (N_19565,N_18922,N_18906);
nor U19566 (N_19566,N_18912,N_18541);
nand U19567 (N_19567,N_18665,N_18954);
nor U19568 (N_19568,N_18965,N_18696);
nor U19569 (N_19569,N_19086,N_18750);
or U19570 (N_19570,N_18465,N_18464);
xor U19571 (N_19571,N_19050,N_18433);
and U19572 (N_19572,N_19022,N_18829);
nor U19573 (N_19573,N_19095,N_18764);
xor U19574 (N_19574,N_18474,N_18459);
xnor U19575 (N_19575,N_18455,N_18577);
and U19576 (N_19576,N_19028,N_18975);
xnor U19577 (N_19577,N_18698,N_18870);
xnor U19578 (N_19578,N_18548,N_19042);
and U19579 (N_19579,N_18837,N_18964);
nand U19580 (N_19580,N_18716,N_18832);
and U19581 (N_19581,N_19078,N_18889);
nor U19582 (N_19582,N_18431,N_18434);
xnor U19583 (N_19583,N_18762,N_18956);
nor U19584 (N_19584,N_19106,N_18973);
nor U19585 (N_19585,N_18819,N_18715);
xnor U19586 (N_19586,N_18743,N_19076);
and U19587 (N_19587,N_18713,N_18997);
nand U19588 (N_19588,N_18491,N_19160);
nand U19589 (N_19589,N_18471,N_18564);
and U19590 (N_19590,N_19146,N_18659);
xnor U19591 (N_19591,N_18601,N_18736);
nand U19592 (N_19592,N_18676,N_18939);
nor U19593 (N_19593,N_18844,N_19142);
nand U19594 (N_19594,N_18733,N_18585);
and U19595 (N_19595,N_18788,N_18613);
nand U19596 (N_19596,N_18622,N_18726);
and U19597 (N_19597,N_18502,N_18576);
nor U19598 (N_19598,N_18981,N_18425);
xor U19599 (N_19599,N_18994,N_18644);
nand U19600 (N_19600,N_18692,N_18622);
xor U19601 (N_19601,N_18797,N_19016);
nand U19602 (N_19602,N_18827,N_18605);
nor U19603 (N_19603,N_18929,N_18491);
and U19604 (N_19604,N_18433,N_18964);
and U19605 (N_19605,N_18702,N_18577);
nand U19606 (N_19606,N_18978,N_18660);
nand U19607 (N_19607,N_18407,N_18983);
nand U19608 (N_19608,N_18792,N_18630);
xor U19609 (N_19609,N_18669,N_18748);
or U19610 (N_19610,N_18786,N_18848);
nand U19611 (N_19611,N_18774,N_19021);
or U19612 (N_19612,N_18803,N_18688);
or U19613 (N_19613,N_18570,N_18817);
xor U19614 (N_19614,N_18562,N_18407);
nand U19615 (N_19615,N_18446,N_18498);
xor U19616 (N_19616,N_18807,N_18550);
or U19617 (N_19617,N_18688,N_18512);
nor U19618 (N_19618,N_18456,N_18927);
xnor U19619 (N_19619,N_18548,N_18614);
or U19620 (N_19620,N_18729,N_18722);
nor U19621 (N_19621,N_19023,N_18814);
nor U19622 (N_19622,N_19165,N_19026);
or U19623 (N_19623,N_19197,N_18796);
or U19624 (N_19624,N_18498,N_18655);
xor U19625 (N_19625,N_18776,N_18661);
or U19626 (N_19626,N_19017,N_18715);
and U19627 (N_19627,N_18878,N_18431);
and U19628 (N_19628,N_19156,N_19132);
and U19629 (N_19629,N_18551,N_19068);
and U19630 (N_19630,N_18888,N_18833);
nand U19631 (N_19631,N_18780,N_18702);
and U19632 (N_19632,N_18901,N_19031);
and U19633 (N_19633,N_18491,N_18406);
xnor U19634 (N_19634,N_18577,N_18588);
and U19635 (N_19635,N_18700,N_18520);
xnor U19636 (N_19636,N_18689,N_19136);
and U19637 (N_19637,N_18945,N_18839);
and U19638 (N_19638,N_19192,N_18537);
and U19639 (N_19639,N_18526,N_18583);
or U19640 (N_19640,N_18674,N_18401);
nand U19641 (N_19641,N_18975,N_18793);
nand U19642 (N_19642,N_18830,N_18988);
or U19643 (N_19643,N_18882,N_19074);
or U19644 (N_19644,N_19065,N_18405);
nor U19645 (N_19645,N_19147,N_18872);
nor U19646 (N_19646,N_18798,N_18595);
nand U19647 (N_19647,N_19165,N_18900);
nand U19648 (N_19648,N_19005,N_18559);
xor U19649 (N_19649,N_18928,N_19014);
xor U19650 (N_19650,N_18873,N_18615);
xnor U19651 (N_19651,N_18627,N_18630);
xnor U19652 (N_19652,N_19057,N_18510);
nand U19653 (N_19653,N_18476,N_18802);
or U19654 (N_19654,N_18850,N_18975);
or U19655 (N_19655,N_18886,N_18452);
nand U19656 (N_19656,N_18818,N_19014);
nand U19657 (N_19657,N_18831,N_18589);
or U19658 (N_19658,N_19052,N_18996);
or U19659 (N_19659,N_18787,N_18953);
or U19660 (N_19660,N_19173,N_18639);
and U19661 (N_19661,N_18593,N_18452);
nor U19662 (N_19662,N_18619,N_19053);
and U19663 (N_19663,N_18708,N_18461);
and U19664 (N_19664,N_18657,N_19054);
nand U19665 (N_19665,N_19025,N_18508);
nand U19666 (N_19666,N_18494,N_18421);
nor U19667 (N_19667,N_19144,N_18965);
nand U19668 (N_19668,N_18976,N_18484);
or U19669 (N_19669,N_18563,N_18622);
or U19670 (N_19670,N_19000,N_18616);
or U19671 (N_19671,N_18782,N_19054);
or U19672 (N_19672,N_18555,N_18661);
nor U19673 (N_19673,N_19043,N_18947);
or U19674 (N_19674,N_18683,N_18798);
nor U19675 (N_19675,N_19026,N_18450);
nand U19676 (N_19676,N_18802,N_18879);
nand U19677 (N_19677,N_19131,N_18779);
xor U19678 (N_19678,N_18698,N_18605);
and U19679 (N_19679,N_18634,N_19029);
nor U19680 (N_19680,N_18430,N_18554);
or U19681 (N_19681,N_18432,N_18995);
nand U19682 (N_19682,N_19132,N_18875);
or U19683 (N_19683,N_18683,N_18599);
nand U19684 (N_19684,N_18615,N_19146);
nor U19685 (N_19685,N_18678,N_19087);
nand U19686 (N_19686,N_19090,N_18902);
xnor U19687 (N_19687,N_18881,N_18569);
nand U19688 (N_19688,N_18536,N_18730);
or U19689 (N_19689,N_19049,N_19077);
nand U19690 (N_19690,N_19199,N_18977);
nor U19691 (N_19691,N_19106,N_18451);
or U19692 (N_19692,N_18984,N_18960);
xor U19693 (N_19693,N_18550,N_18667);
nand U19694 (N_19694,N_18697,N_18541);
and U19695 (N_19695,N_18554,N_18949);
or U19696 (N_19696,N_18470,N_19077);
nand U19697 (N_19697,N_18848,N_19029);
nor U19698 (N_19698,N_18406,N_18953);
and U19699 (N_19699,N_18420,N_18905);
nor U19700 (N_19700,N_18501,N_18443);
or U19701 (N_19701,N_18653,N_19153);
or U19702 (N_19702,N_18432,N_18824);
nand U19703 (N_19703,N_18581,N_19108);
and U19704 (N_19704,N_18642,N_18534);
nand U19705 (N_19705,N_18572,N_18442);
or U19706 (N_19706,N_19085,N_19156);
or U19707 (N_19707,N_19118,N_19109);
and U19708 (N_19708,N_18638,N_18903);
xnor U19709 (N_19709,N_18651,N_18739);
or U19710 (N_19710,N_18566,N_19023);
nand U19711 (N_19711,N_18494,N_18939);
nor U19712 (N_19712,N_18401,N_18488);
or U19713 (N_19713,N_18763,N_18903);
xor U19714 (N_19714,N_18474,N_18818);
or U19715 (N_19715,N_18823,N_18875);
xor U19716 (N_19716,N_18861,N_19029);
xor U19717 (N_19717,N_18477,N_19036);
or U19718 (N_19718,N_18506,N_18542);
and U19719 (N_19719,N_19186,N_18926);
xnor U19720 (N_19720,N_18750,N_19084);
nand U19721 (N_19721,N_19069,N_18892);
xnor U19722 (N_19722,N_19089,N_18464);
nor U19723 (N_19723,N_19018,N_18787);
nand U19724 (N_19724,N_18710,N_19180);
xnor U19725 (N_19725,N_19167,N_18449);
nand U19726 (N_19726,N_19116,N_18971);
nand U19727 (N_19727,N_18566,N_18676);
nor U19728 (N_19728,N_18405,N_18469);
nor U19729 (N_19729,N_18717,N_18853);
nor U19730 (N_19730,N_19151,N_18427);
and U19731 (N_19731,N_18535,N_18662);
or U19732 (N_19732,N_19084,N_19104);
nor U19733 (N_19733,N_19078,N_19154);
and U19734 (N_19734,N_19165,N_18951);
xnor U19735 (N_19735,N_19199,N_18416);
nor U19736 (N_19736,N_18485,N_18933);
or U19737 (N_19737,N_18762,N_18994);
or U19738 (N_19738,N_18532,N_18763);
nor U19739 (N_19739,N_18524,N_18635);
nor U19740 (N_19740,N_18807,N_18477);
nor U19741 (N_19741,N_18854,N_18955);
nor U19742 (N_19742,N_18787,N_18812);
nand U19743 (N_19743,N_19053,N_18869);
nand U19744 (N_19744,N_19071,N_18871);
nor U19745 (N_19745,N_18943,N_18735);
or U19746 (N_19746,N_18662,N_18987);
and U19747 (N_19747,N_18656,N_18680);
nand U19748 (N_19748,N_18419,N_18538);
nand U19749 (N_19749,N_18677,N_18642);
nor U19750 (N_19750,N_18988,N_18767);
or U19751 (N_19751,N_18841,N_18894);
nor U19752 (N_19752,N_18807,N_18567);
and U19753 (N_19753,N_18925,N_19023);
or U19754 (N_19754,N_18578,N_19078);
nor U19755 (N_19755,N_18479,N_19011);
nor U19756 (N_19756,N_18842,N_18599);
nand U19757 (N_19757,N_18750,N_18806);
nand U19758 (N_19758,N_18459,N_18539);
xor U19759 (N_19759,N_19177,N_18425);
nor U19760 (N_19760,N_18597,N_18631);
or U19761 (N_19761,N_18803,N_19054);
or U19762 (N_19762,N_18966,N_18981);
or U19763 (N_19763,N_18687,N_18957);
and U19764 (N_19764,N_18837,N_19164);
or U19765 (N_19765,N_19119,N_18988);
and U19766 (N_19766,N_18538,N_19013);
or U19767 (N_19767,N_18449,N_19186);
and U19768 (N_19768,N_18914,N_18854);
or U19769 (N_19769,N_18535,N_18748);
or U19770 (N_19770,N_18822,N_18808);
and U19771 (N_19771,N_18588,N_18988);
and U19772 (N_19772,N_18827,N_18652);
and U19773 (N_19773,N_19125,N_18992);
xnor U19774 (N_19774,N_19104,N_18610);
or U19775 (N_19775,N_18992,N_19001);
nand U19776 (N_19776,N_18784,N_18742);
nor U19777 (N_19777,N_18873,N_19036);
xor U19778 (N_19778,N_18405,N_18998);
nand U19779 (N_19779,N_18948,N_18703);
nand U19780 (N_19780,N_19111,N_18463);
and U19781 (N_19781,N_18473,N_18517);
nor U19782 (N_19782,N_18461,N_19071);
or U19783 (N_19783,N_18948,N_18785);
and U19784 (N_19784,N_18488,N_18485);
nand U19785 (N_19785,N_18724,N_18707);
nand U19786 (N_19786,N_19189,N_19103);
or U19787 (N_19787,N_19067,N_19134);
or U19788 (N_19788,N_18472,N_18408);
xor U19789 (N_19789,N_18865,N_19132);
nand U19790 (N_19790,N_18584,N_19150);
nor U19791 (N_19791,N_18435,N_19095);
xnor U19792 (N_19792,N_18492,N_19064);
and U19793 (N_19793,N_19024,N_18928);
and U19794 (N_19794,N_18948,N_18943);
xnor U19795 (N_19795,N_18969,N_18553);
nand U19796 (N_19796,N_18467,N_19107);
nand U19797 (N_19797,N_18630,N_19158);
and U19798 (N_19798,N_18873,N_18509);
xnor U19799 (N_19799,N_18680,N_18967);
and U19800 (N_19800,N_18700,N_18742);
and U19801 (N_19801,N_18514,N_19134);
or U19802 (N_19802,N_18874,N_18657);
or U19803 (N_19803,N_18680,N_18642);
xor U19804 (N_19804,N_18907,N_18814);
or U19805 (N_19805,N_18927,N_18876);
xnor U19806 (N_19806,N_19180,N_19195);
or U19807 (N_19807,N_18666,N_18712);
and U19808 (N_19808,N_18600,N_19075);
nand U19809 (N_19809,N_19033,N_18628);
and U19810 (N_19810,N_18484,N_18813);
nor U19811 (N_19811,N_18724,N_19191);
and U19812 (N_19812,N_18804,N_18571);
nand U19813 (N_19813,N_18463,N_18568);
xor U19814 (N_19814,N_18961,N_18697);
or U19815 (N_19815,N_18886,N_18537);
nor U19816 (N_19816,N_18500,N_19097);
and U19817 (N_19817,N_18869,N_18848);
nand U19818 (N_19818,N_19057,N_19172);
and U19819 (N_19819,N_18713,N_18821);
nor U19820 (N_19820,N_18501,N_18655);
and U19821 (N_19821,N_18790,N_18611);
xor U19822 (N_19822,N_19068,N_18930);
or U19823 (N_19823,N_19119,N_18881);
nor U19824 (N_19824,N_18885,N_18822);
xor U19825 (N_19825,N_18845,N_18480);
nor U19826 (N_19826,N_18776,N_18983);
and U19827 (N_19827,N_18692,N_18818);
nor U19828 (N_19828,N_18560,N_18614);
nor U19829 (N_19829,N_18645,N_19092);
xnor U19830 (N_19830,N_18694,N_19027);
nand U19831 (N_19831,N_18544,N_18801);
or U19832 (N_19832,N_18842,N_19017);
nand U19833 (N_19833,N_18902,N_18910);
xnor U19834 (N_19834,N_18730,N_18608);
nand U19835 (N_19835,N_18747,N_19172);
or U19836 (N_19836,N_19146,N_19111);
nor U19837 (N_19837,N_19165,N_18407);
nor U19838 (N_19838,N_19001,N_18914);
and U19839 (N_19839,N_19041,N_19068);
and U19840 (N_19840,N_18434,N_18733);
xnor U19841 (N_19841,N_18939,N_18537);
or U19842 (N_19842,N_18806,N_18963);
xor U19843 (N_19843,N_18974,N_18490);
xnor U19844 (N_19844,N_18576,N_18409);
and U19845 (N_19845,N_18694,N_19011);
nor U19846 (N_19846,N_19049,N_19119);
xnor U19847 (N_19847,N_18972,N_18561);
and U19848 (N_19848,N_18942,N_18813);
or U19849 (N_19849,N_18613,N_18706);
nor U19850 (N_19850,N_18511,N_18765);
nor U19851 (N_19851,N_18626,N_18852);
xnor U19852 (N_19852,N_19042,N_19199);
and U19853 (N_19853,N_19190,N_19052);
xnor U19854 (N_19854,N_19056,N_18559);
and U19855 (N_19855,N_18710,N_18769);
and U19856 (N_19856,N_18856,N_18907);
or U19857 (N_19857,N_18413,N_18565);
nor U19858 (N_19858,N_18911,N_18518);
nor U19859 (N_19859,N_18443,N_19046);
nand U19860 (N_19860,N_18450,N_18464);
or U19861 (N_19861,N_18442,N_18498);
nor U19862 (N_19862,N_18719,N_18457);
nor U19863 (N_19863,N_18517,N_18744);
or U19864 (N_19864,N_19123,N_18910);
nor U19865 (N_19865,N_19089,N_18531);
and U19866 (N_19866,N_19106,N_18722);
nand U19867 (N_19867,N_18849,N_18618);
nor U19868 (N_19868,N_19001,N_18742);
xnor U19869 (N_19869,N_18895,N_18490);
xor U19870 (N_19870,N_18732,N_19102);
nor U19871 (N_19871,N_18868,N_18872);
nor U19872 (N_19872,N_18553,N_18761);
nor U19873 (N_19873,N_18564,N_18892);
or U19874 (N_19874,N_18901,N_18670);
and U19875 (N_19875,N_18610,N_18654);
or U19876 (N_19876,N_18577,N_18443);
nand U19877 (N_19877,N_18741,N_18969);
nand U19878 (N_19878,N_18783,N_18578);
nand U19879 (N_19879,N_19175,N_18547);
and U19880 (N_19880,N_18553,N_18941);
xnor U19881 (N_19881,N_19198,N_18955);
xnor U19882 (N_19882,N_18743,N_18660);
and U19883 (N_19883,N_18780,N_18413);
and U19884 (N_19884,N_18537,N_18757);
nand U19885 (N_19885,N_18957,N_18884);
xor U19886 (N_19886,N_19095,N_18751);
or U19887 (N_19887,N_18633,N_18556);
or U19888 (N_19888,N_18439,N_18716);
xnor U19889 (N_19889,N_18843,N_18422);
nand U19890 (N_19890,N_18736,N_19163);
nor U19891 (N_19891,N_18609,N_18778);
nor U19892 (N_19892,N_18838,N_19027);
xor U19893 (N_19893,N_18602,N_19118);
nand U19894 (N_19894,N_19124,N_18868);
xnor U19895 (N_19895,N_18970,N_18936);
xnor U19896 (N_19896,N_18415,N_18645);
and U19897 (N_19897,N_18707,N_18508);
nor U19898 (N_19898,N_18977,N_18527);
and U19899 (N_19899,N_19037,N_18880);
and U19900 (N_19900,N_19071,N_18745);
and U19901 (N_19901,N_18734,N_18592);
or U19902 (N_19902,N_18744,N_18911);
nor U19903 (N_19903,N_19190,N_18995);
nor U19904 (N_19904,N_19125,N_18876);
and U19905 (N_19905,N_18781,N_18750);
nor U19906 (N_19906,N_18423,N_18431);
nand U19907 (N_19907,N_18763,N_18426);
nand U19908 (N_19908,N_18819,N_18598);
xnor U19909 (N_19909,N_19112,N_18438);
and U19910 (N_19910,N_18488,N_18754);
nor U19911 (N_19911,N_18411,N_18440);
and U19912 (N_19912,N_18833,N_19066);
and U19913 (N_19913,N_19031,N_18528);
xnor U19914 (N_19914,N_18427,N_18524);
nor U19915 (N_19915,N_19111,N_19097);
or U19916 (N_19916,N_19113,N_19021);
or U19917 (N_19917,N_18769,N_18626);
nand U19918 (N_19918,N_19196,N_18711);
nor U19919 (N_19919,N_18710,N_18529);
or U19920 (N_19920,N_18853,N_18812);
and U19921 (N_19921,N_18965,N_18653);
xnor U19922 (N_19922,N_19114,N_19078);
or U19923 (N_19923,N_18856,N_18837);
nor U19924 (N_19924,N_19037,N_18470);
nand U19925 (N_19925,N_18492,N_19109);
or U19926 (N_19926,N_18953,N_18945);
xor U19927 (N_19927,N_18645,N_18555);
or U19928 (N_19928,N_19099,N_18424);
nand U19929 (N_19929,N_18955,N_18618);
nand U19930 (N_19930,N_18519,N_18638);
nor U19931 (N_19931,N_19159,N_18636);
and U19932 (N_19932,N_18561,N_18766);
and U19933 (N_19933,N_19062,N_18477);
nand U19934 (N_19934,N_18840,N_18911);
and U19935 (N_19935,N_18891,N_18673);
nor U19936 (N_19936,N_18640,N_19124);
nand U19937 (N_19937,N_18527,N_18610);
xor U19938 (N_19938,N_18977,N_18537);
xor U19939 (N_19939,N_18543,N_18760);
and U19940 (N_19940,N_18576,N_18468);
nor U19941 (N_19941,N_19062,N_18692);
xnor U19942 (N_19942,N_18613,N_18671);
nor U19943 (N_19943,N_18733,N_18943);
and U19944 (N_19944,N_19141,N_18453);
xnor U19945 (N_19945,N_19047,N_18494);
nor U19946 (N_19946,N_19106,N_18755);
nor U19947 (N_19947,N_18832,N_18698);
xor U19948 (N_19948,N_19088,N_19028);
nor U19949 (N_19949,N_18564,N_18638);
xnor U19950 (N_19950,N_19075,N_18895);
nor U19951 (N_19951,N_19178,N_19054);
nand U19952 (N_19952,N_18956,N_18748);
nor U19953 (N_19953,N_18737,N_18657);
nand U19954 (N_19954,N_18618,N_19148);
nand U19955 (N_19955,N_18632,N_18827);
or U19956 (N_19956,N_18737,N_18972);
or U19957 (N_19957,N_18453,N_19078);
xor U19958 (N_19958,N_18684,N_18938);
nand U19959 (N_19959,N_18905,N_18971);
or U19960 (N_19960,N_18923,N_18952);
xor U19961 (N_19961,N_18966,N_18594);
nand U19962 (N_19962,N_19118,N_18414);
nor U19963 (N_19963,N_18800,N_18738);
xnor U19964 (N_19964,N_19027,N_19040);
nor U19965 (N_19965,N_18479,N_19092);
nor U19966 (N_19966,N_18497,N_18745);
and U19967 (N_19967,N_18417,N_18977);
and U19968 (N_19968,N_18460,N_18638);
and U19969 (N_19969,N_18779,N_19113);
nor U19970 (N_19970,N_18510,N_18637);
or U19971 (N_19971,N_19169,N_19130);
nand U19972 (N_19972,N_19119,N_18831);
xnor U19973 (N_19973,N_19080,N_18697);
xor U19974 (N_19974,N_18603,N_18665);
and U19975 (N_19975,N_18804,N_18668);
nor U19976 (N_19976,N_18506,N_19035);
nor U19977 (N_19977,N_18969,N_19178);
xor U19978 (N_19978,N_18565,N_18818);
nor U19979 (N_19979,N_18493,N_18656);
or U19980 (N_19980,N_18703,N_18405);
xnor U19981 (N_19981,N_18436,N_18537);
xnor U19982 (N_19982,N_18538,N_18659);
nand U19983 (N_19983,N_19136,N_18828);
nor U19984 (N_19984,N_18566,N_18502);
nor U19985 (N_19985,N_18749,N_18595);
xor U19986 (N_19986,N_18588,N_19015);
or U19987 (N_19987,N_18885,N_18793);
and U19988 (N_19988,N_18623,N_19169);
and U19989 (N_19989,N_18419,N_18448);
nor U19990 (N_19990,N_19041,N_18979);
or U19991 (N_19991,N_18524,N_18655);
xor U19992 (N_19992,N_18898,N_19108);
nor U19993 (N_19993,N_18727,N_18406);
or U19994 (N_19994,N_18456,N_18613);
or U19995 (N_19995,N_18756,N_18665);
or U19996 (N_19996,N_18465,N_19048);
xnor U19997 (N_19997,N_18941,N_18684);
xnor U19998 (N_19998,N_18964,N_19006);
xnor U19999 (N_19999,N_19008,N_18840);
and UO_0 (O_0,N_19460,N_19834);
nand UO_1 (O_1,N_19390,N_19290);
or UO_2 (O_2,N_19853,N_19915);
and UO_3 (O_3,N_19407,N_19416);
nand UO_4 (O_4,N_19607,N_19908);
and UO_5 (O_5,N_19485,N_19897);
and UO_6 (O_6,N_19226,N_19224);
xnor UO_7 (O_7,N_19941,N_19274);
nand UO_8 (O_8,N_19272,N_19669);
nand UO_9 (O_9,N_19413,N_19910);
nor UO_10 (O_10,N_19999,N_19754);
and UO_11 (O_11,N_19928,N_19716);
nor UO_12 (O_12,N_19392,N_19775);
xor UO_13 (O_13,N_19449,N_19332);
nand UO_14 (O_14,N_19396,N_19538);
nand UO_15 (O_15,N_19267,N_19901);
nor UO_16 (O_16,N_19672,N_19540);
xnor UO_17 (O_17,N_19849,N_19277);
nand UO_18 (O_18,N_19599,N_19745);
or UO_19 (O_19,N_19785,N_19920);
xnor UO_20 (O_20,N_19596,N_19615);
or UO_21 (O_21,N_19931,N_19981);
and UO_22 (O_22,N_19674,N_19822);
xnor UO_23 (O_23,N_19621,N_19531);
or UO_24 (O_24,N_19682,N_19991);
and UO_25 (O_25,N_19735,N_19365);
or UO_26 (O_26,N_19911,N_19964);
xor UO_27 (O_27,N_19425,N_19927);
or UO_28 (O_28,N_19397,N_19287);
nor UO_29 (O_29,N_19270,N_19994);
and UO_30 (O_30,N_19547,N_19631);
xor UO_31 (O_31,N_19266,N_19329);
xor UO_32 (O_32,N_19595,N_19320);
nor UO_33 (O_33,N_19770,N_19393);
and UO_34 (O_34,N_19988,N_19213);
and UO_35 (O_35,N_19500,N_19658);
nor UO_36 (O_36,N_19537,N_19411);
and UO_37 (O_37,N_19781,N_19334);
nor UO_38 (O_38,N_19516,N_19526);
or UO_39 (O_39,N_19616,N_19482);
or UO_40 (O_40,N_19541,N_19656);
and UO_41 (O_41,N_19427,N_19786);
and UO_42 (O_42,N_19336,N_19456);
or UO_43 (O_43,N_19574,N_19326);
or UO_44 (O_44,N_19455,N_19493);
and UO_45 (O_45,N_19697,N_19255);
xor UO_46 (O_46,N_19844,N_19592);
nor UO_47 (O_47,N_19230,N_19861);
xor UO_48 (O_48,N_19661,N_19546);
and UO_49 (O_49,N_19652,N_19391);
and UO_50 (O_50,N_19798,N_19666);
and UO_51 (O_51,N_19622,N_19415);
nor UO_52 (O_52,N_19423,N_19344);
or UO_53 (O_53,N_19828,N_19569);
xor UO_54 (O_54,N_19657,N_19315);
xnor UO_55 (O_55,N_19986,N_19387);
or UO_56 (O_56,N_19896,N_19434);
or UO_57 (O_57,N_19231,N_19937);
and UO_58 (O_58,N_19247,N_19648);
and UO_59 (O_59,N_19576,N_19629);
or UO_60 (O_60,N_19761,N_19527);
or UO_61 (O_61,N_19588,N_19357);
or UO_62 (O_62,N_19635,N_19579);
nor UO_63 (O_63,N_19814,N_19550);
or UO_64 (O_64,N_19571,N_19771);
xnor UO_65 (O_65,N_19206,N_19474);
and UO_66 (O_66,N_19322,N_19330);
or UO_67 (O_67,N_19843,N_19203);
and UO_68 (O_68,N_19281,N_19860);
xnor UO_69 (O_69,N_19806,N_19829);
nand UO_70 (O_70,N_19204,N_19317);
and UO_71 (O_71,N_19842,N_19545);
and UO_72 (O_72,N_19762,N_19536);
or UO_73 (O_73,N_19637,N_19633);
nor UO_74 (O_74,N_19623,N_19659);
nand UO_75 (O_75,N_19712,N_19371);
or UO_76 (O_76,N_19519,N_19566);
nor UO_77 (O_77,N_19216,N_19401);
or UO_78 (O_78,N_19684,N_19318);
nor UO_79 (O_79,N_19891,N_19488);
nand UO_80 (O_80,N_19280,N_19951);
nand UO_81 (O_81,N_19900,N_19307);
and UO_82 (O_82,N_19740,N_19305);
and UO_83 (O_83,N_19398,N_19238);
nor UO_84 (O_84,N_19506,N_19992);
nor UO_85 (O_85,N_19608,N_19801);
or UO_86 (O_86,N_19732,N_19851);
xor UO_87 (O_87,N_19980,N_19211);
and UO_88 (O_88,N_19653,N_19877);
and UO_89 (O_89,N_19892,N_19314);
nand UO_90 (O_90,N_19587,N_19953);
or UO_91 (O_91,N_19966,N_19373);
nand UO_92 (O_92,N_19311,N_19580);
xor UO_93 (O_93,N_19403,N_19530);
nand UO_94 (O_94,N_19711,N_19495);
and UO_95 (O_95,N_19998,N_19993);
nor UO_96 (O_96,N_19225,N_19555);
nand UO_97 (O_97,N_19233,N_19219);
and UO_98 (O_98,N_19817,N_19810);
nand UO_99 (O_99,N_19708,N_19939);
nor UO_100 (O_100,N_19399,N_19405);
nand UO_101 (O_101,N_19421,N_19720);
or UO_102 (O_102,N_19959,N_19316);
and UO_103 (O_103,N_19300,N_19222);
nand UO_104 (O_104,N_19356,N_19288);
and UO_105 (O_105,N_19691,N_19729);
and UO_106 (O_106,N_19501,N_19207);
xor UO_107 (O_107,N_19543,N_19979);
and UO_108 (O_108,N_19972,N_19996);
nand UO_109 (O_109,N_19551,N_19960);
xnor UO_110 (O_110,N_19378,N_19780);
nor UO_111 (O_111,N_19848,N_19673);
or UO_112 (O_112,N_19492,N_19874);
nor UO_113 (O_113,N_19795,N_19563);
nand UO_114 (O_114,N_19593,N_19961);
nand UO_115 (O_115,N_19955,N_19406);
and UO_116 (O_116,N_19445,N_19809);
nand UO_117 (O_117,N_19723,N_19997);
nor UO_118 (O_118,N_19469,N_19757);
or UO_119 (O_119,N_19298,N_19384);
and UO_120 (O_120,N_19221,N_19451);
or UO_121 (O_121,N_19858,N_19328);
nand UO_122 (O_122,N_19889,N_19769);
nor UO_123 (O_123,N_19605,N_19251);
and UO_124 (O_124,N_19513,N_19971);
nor UO_125 (O_125,N_19505,N_19448);
nor UO_126 (O_126,N_19826,N_19995);
nand UO_127 (O_127,N_19907,N_19453);
nor UO_128 (O_128,N_19232,N_19544);
nor UO_129 (O_129,N_19480,N_19627);
nand UO_130 (O_130,N_19533,N_19949);
xor UO_131 (O_131,N_19856,N_19586);
or UO_132 (O_132,N_19778,N_19292);
and UO_133 (O_133,N_19787,N_19847);
or UO_134 (O_134,N_19701,N_19755);
or UO_135 (O_135,N_19581,N_19990);
xor UO_136 (O_136,N_19234,N_19278);
xor UO_137 (O_137,N_19218,N_19873);
nand UO_138 (O_138,N_19634,N_19525);
nand UO_139 (O_139,N_19952,N_19878);
and UO_140 (O_140,N_19630,N_19776);
and UO_141 (O_141,N_19763,N_19948);
nor UO_142 (O_142,N_19854,N_19369);
and UO_143 (O_143,N_19647,N_19906);
or UO_144 (O_144,N_19650,N_19839);
and UO_145 (O_145,N_19676,N_19268);
and UO_146 (O_146,N_19984,N_19575);
xnor UO_147 (O_147,N_19921,N_19313);
and UO_148 (O_148,N_19728,N_19283);
nand UO_149 (O_149,N_19804,N_19905);
xnor UO_150 (O_150,N_19982,N_19430);
nor UO_151 (O_151,N_19916,N_19613);
and UO_152 (O_152,N_19361,N_19976);
nand UO_153 (O_153,N_19700,N_19584);
and UO_154 (O_154,N_19514,N_19428);
or UO_155 (O_155,N_19417,N_19567);
and UO_156 (O_156,N_19954,N_19914);
and UO_157 (O_157,N_19259,N_19509);
and UO_158 (O_158,N_19523,N_19600);
nor UO_159 (O_159,N_19522,N_19515);
nand UO_160 (O_160,N_19335,N_19749);
or UO_161 (O_161,N_19899,N_19626);
and UO_162 (O_162,N_19699,N_19302);
xor UO_163 (O_163,N_19312,N_19375);
nor UO_164 (O_164,N_19840,N_19303);
nor UO_165 (O_165,N_19386,N_19866);
nor UO_166 (O_166,N_19667,N_19556);
or UO_167 (O_167,N_19675,N_19461);
or UO_168 (O_168,N_19855,N_19354);
nand UO_169 (O_169,N_19338,N_19765);
and UO_170 (O_170,N_19358,N_19802);
nor UO_171 (O_171,N_19671,N_19490);
or UO_172 (O_172,N_19202,N_19258);
nor UO_173 (O_173,N_19987,N_19632);
xnor UO_174 (O_174,N_19422,N_19459);
xor UO_175 (O_175,N_19904,N_19898);
nor UO_176 (O_176,N_19831,N_19929);
nor UO_177 (O_177,N_19465,N_19583);
and UO_178 (O_178,N_19282,N_19208);
nor UO_179 (O_179,N_19350,N_19731);
nand UO_180 (O_180,N_19558,N_19262);
nor UO_181 (O_181,N_19487,N_19337);
and UO_182 (O_182,N_19887,N_19341);
xor UO_183 (O_183,N_19524,N_19973);
xnor UO_184 (O_184,N_19252,N_19359);
or UO_185 (O_185,N_19240,N_19815);
xor UO_186 (O_186,N_19660,N_19850);
nor UO_187 (O_187,N_19510,N_19816);
nor UO_188 (O_188,N_19253,N_19707);
nand UO_189 (O_189,N_19228,N_19559);
nand UO_190 (O_190,N_19738,N_19958);
or UO_191 (O_191,N_19478,N_19823);
nor UO_192 (O_192,N_19894,N_19865);
nor UO_193 (O_193,N_19473,N_19590);
and UO_194 (O_194,N_19433,N_19805);
nor UO_195 (O_195,N_19670,N_19200);
xnor UO_196 (O_196,N_19760,N_19250);
or UO_197 (O_197,N_19962,N_19468);
nand UO_198 (O_198,N_19333,N_19343);
and UO_199 (O_199,N_19719,N_19265);
nor UO_200 (O_200,N_19681,N_19210);
xnor UO_201 (O_201,N_19420,N_19881);
nor UO_202 (O_202,N_19690,N_19394);
and UO_203 (O_203,N_19484,N_19870);
and UO_204 (O_204,N_19685,N_19943);
xor UO_205 (O_205,N_19883,N_19381);
and UO_206 (O_206,N_19746,N_19539);
and UO_207 (O_207,N_19419,N_19875);
xnor UO_208 (O_208,N_19467,N_19957);
or UO_209 (O_209,N_19969,N_19710);
and UO_210 (O_210,N_19886,N_19363);
xnor UO_211 (O_211,N_19466,N_19237);
and UO_212 (O_212,N_19938,N_19528);
nand UO_213 (O_213,N_19561,N_19662);
xor UO_214 (O_214,N_19665,N_19747);
xnor UO_215 (O_215,N_19404,N_19677);
nand UO_216 (O_216,N_19293,N_19871);
nor UO_217 (O_217,N_19367,N_19439);
or UO_218 (O_218,N_19447,N_19235);
xor UO_219 (O_219,N_19400,N_19863);
nor UO_220 (O_220,N_19612,N_19339);
or UO_221 (O_221,N_19926,N_19923);
nor UO_222 (O_222,N_19718,N_19717);
nand UO_223 (O_223,N_19263,N_19876);
nand UO_224 (O_224,N_19687,N_19748);
nand UO_225 (O_225,N_19601,N_19497);
xor UO_226 (O_226,N_19703,N_19560);
and UO_227 (O_227,N_19726,N_19520);
nand UO_228 (O_228,N_19442,N_19651);
and UO_229 (O_229,N_19783,N_19893);
and UO_230 (O_230,N_19903,N_19532);
or UO_231 (O_231,N_19784,N_19619);
and UO_232 (O_232,N_19970,N_19841);
xor UO_233 (O_233,N_19812,N_19846);
nand UO_234 (O_234,N_19680,N_19715);
nor UO_235 (O_235,N_19362,N_19435);
or UO_236 (O_236,N_19286,N_19909);
nor UO_237 (O_237,N_19800,N_19942);
xor UO_238 (O_238,N_19441,N_19734);
and UO_239 (O_239,N_19917,N_19888);
nor UO_240 (O_240,N_19838,N_19628);
xor UO_241 (O_241,N_19603,N_19779);
nand UO_242 (O_242,N_19248,N_19736);
xnor UO_243 (O_243,N_19985,N_19772);
nor UO_244 (O_244,N_19370,N_19645);
and UO_245 (O_245,N_19799,N_19742);
xor UO_246 (O_246,N_19773,N_19353);
nor UO_247 (O_247,N_19882,N_19796);
or UO_248 (O_248,N_19444,N_19217);
nand UO_249 (O_249,N_19975,N_19486);
xnor UO_250 (O_250,N_19534,N_19457);
nand UO_251 (O_251,N_19348,N_19688);
and UO_252 (O_252,N_19429,N_19827);
nand UO_253 (O_253,N_19963,N_19275);
or UO_254 (O_254,N_19242,N_19297);
and UO_255 (O_255,N_19852,N_19725);
and UO_256 (O_256,N_19436,N_19604);
or UO_257 (O_257,N_19377,N_19254);
and UO_258 (O_258,N_19777,N_19517);
xor UO_259 (O_259,N_19376,N_19935);
or UO_260 (O_260,N_19304,N_19368);
nand UO_261 (O_261,N_19807,N_19483);
or UO_262 (O_262,N_19884,N_19294);
xnor UO_263 (O_263,N_19643,N_19913);
or UO_264 (O_264,N_19830,N_19568);
nor UO_265 (O_265,N_19352,N_19241);
and UO_266 (O_266,N_19714,N_19945);
or UO_267 (O_267,N_19214,N_19331);
and UO_268 (O_268,N_19646,N_19296);
and UO_269 (O_269,N_19470,N_19562);
and UO_270 (O_270,N_19880,N_19789);
nand UO_271 (O_271,N_19950,N_19989);
or UO_272 (O_272,N_19744,N_19649);
xnor UO_273 (O_273,N_19983,N_19965);
nor UO_274 (O_274,N_19758,N_19803);
nor UO_275 (O_275,N_19790,N_19611);
and UO_276 (O_276,N_19458,N_19310);
nor UO_277 (O_277,N_19835,N_19788);
nand UO_278 (O_278,N_19751,N_19308);
or UO_279 (O_279,N_19602,N_19382);
xnor UO_280 (O_280,N_19836,N_19655);
nand UO_281 (O_281,N_19309,N_19557);
and UO_282 (O_282,N_19223,N_19625);
nand UO_283 (O_283,N_19733,N_19366);
nand UO_284 (O_284,N_19383,N_19380);
nor UO_285 (O_285,N_19479,N_19511);
and UO_286 (O_286,N_19437,N_19813);
nand UO_287 (O_287,N_19766,N_19295);
nor UO_288 (O_288,N_19349,N_19695);
xor UO_289 (O_289,N_19289,N_19974);
or UO_290 (O_290,N_19640,N_19597);
nor UO_291 (O_291,N_19654,N_19679);
nor UO_292 (O_292,N_19837,N_19934);
nand UO_293 (O_293,N_19491,N_19476);
xor UO_294 (O_294,N_19918,N_19229);
and UO_295 (O_295,N_19496,N_19782);
or UO_296 (O_296,N_19857,N_19440);
xor UO_297 (O_297,N_19489,N_19864);
or UO_298 (O_298,N_19610,N_19730);
nor UO_299 (O_299,N_19319,N_19885);
nand UO_300 (O_300,N_19768,N_19301);
nand UO_301 (O_301,N_19872,N_19347);
or UO_302 (O_302,N_19912,N_19614);
nand UO_303 (O_303,N_19832,N_19767);
and UO_304 (O_304,N_19535,N_19978);
and UO_305 (O_305,N_19323,N_19327);
nand UO_306 (O_306,N_19663,N_19269);
nand UO_307 (O_307,N_19351,N_19585);
or UO_308 (O_308,N_19573,N_19598);
xnor UO_309 (O_309,N_19578,N_19564);
xor UO_310 (O_310,N_19694,N_19220);
nor UO_311 (O_311,N_19862,N_19408);
nor UO_312 (O_312,N_19257,N_19925);
and UO_313 (O_313,N_19572,N_19845);
and UO_314 (O_314,N_19494,N_19209);
nand UO_315 (O_315,N_19821,N_19824);
nand UO_316 (O_316,N_19791,N_19818);
nand UO_317 (O_317,N_19529,N_19792);
nand UO_318 (O_318,N_19698,N_19412);
nand UO_319 (O_319,N_19683,N_19704);
and UO_320 (O_320,N_19753,N_19642);
nand UO_321 (O_321,N_19825,N_19774);
or UO_322 (O_322,N_19324,N_19678);
xor UO_323 (O_323,N_19325,N_19764);
or UO_324 (O_324,N_19379,N_19554);
or UO_325 (O_325,N_19750,N_19759);
or UO_326 (O_326,N_19245,N_19808);
nor UO_327 (O_327,N_19620,N_19276);
or UO_328 (O_328,N_19424,N_19724);
and UO_329 (O_329,N_19542,N_19504);
nand UO_330 (O_330,N_19752,N_19946);
or UO_331 (O_331,N_19705,N_19345);
xnor UO_332 (O_332,N_19552,N_19867);
xnor UO_333 (O_333,N_19285,N_19794);
nor UO_334 (O_334,N_19355,N_19342);
xor UO_335 (O_335,N_19236,N_19570);
or UO_336 (O_336,N_19689,N_19414);
or UO_337 (O_337,N_19922,N_19462);
nor UO_338 (O_338,N_19868,N_19833);
nand UO_339 (O_339,N_19264,N_19443);
xnor UO_340 (O_340,N_19246,N_19664);
or UO_341 (O_341,N_19284,N_19239);
and UO_342 (O_342,N_19895,N_19944);
nand UO_343 (O_343,N_19553,N_19243);
nand UO_344 (O_344,N_19279,N_19507);
or UO_345 (O_345,N_19869,N_19549);
or UO_346 (O_346,N_19638,N_19606);
nor UO_347 (O_347,N_19639,N_19548);
nand UO_348 (O_348,N_19977,N_19388);
xnor UO_349 (O_349,N_19932,N_19967);
nand UO_350 (O_350,N_19582,N_19686);
nand UO_351 (O_351,N_19340,N_19450);
nor UO_352 (O_352,N_19201,N_19956);
xnor UO_353 (O_353,N_19464,N_19260);
nand UO_354 (O_354,N_19409,N_19741);
nand UO_355 (O_355,N_19644,N_19215);
nand UO_356 (O_356,N_19636,N_19521);
nor UO_357 (O_357,N_19321,N_19709);
and UO_358 (O_358,N_19820,N_19793);
nor UO_359 (O_359,N_19936,N_19426);
nand UO_360 (O_360,N_19890,N_19609);
or UO_361 (O_361,N_19696,N_19261);
nand UO_362 (O_362,N_19692,N_19722);
or UO_363 (O_363,N_19299,N_19591);
xor UO_364 (O_364,N_19452,N_19518);
nor UO_365 (O_365,N_19727,N_19463);
and UO_366 (O_366,N_19498,N_19481);
xor UO_367 (O_367,N_19502,N_19212);
and UO_368 (O_368,N_19618,N_19589);
or UO_369 (O_369,N_19706,N_19306);
nand UO_370 (O_370,N_19244,N_19291);
or UO_371 (O_371,N_19713,N_19273);
xor UO_372 (O_372,N_19737,N_19902);
and UO_373 (O_373,N_19668,N_19819);
xnor UO_374 (O_374,N_19364,N_19432);
and UO_375 (O_375,N_19721,N_19471);
xnor UO_376 (O_376,N_19438,N_19508);
xnor UO_377 (O_377,N_19702,N_19271);
xnor UO_378 (O_378,N_19410,N_19811);
nor UO_379 (O_379,N_19879,N_19431);
xnor UO_380 (O_380,N_19249,N_19577);
nand UO_381 (O_381,N_19947,N_19503);
or UO_382 (O_382,N_19205,N_19940);
nor UO_383 (O_383,N_19924,N_19385);
or UO_384 (O_384,N_19693,N_19454);
nand UO_385 (O_385,N_19389,N_19499);
nand UO_386 (O_386,N_19346,N_19395);
and UO_387 (O_387,N_19797,N_19594);
or UO_388 (O_388,N_19374,N_19919);
nor UO_389 (O_389,N_19475,N_19227);
or UO_390 (O_390,N_19402,N_19933);
nand UO_391 (O_391,N_19360,N_19739);
nand UO_392 (O_392,N_19512,N_19256);
and UO_393 (O_393,N_19743,N_19641);
or UO_394 (O_394,N_19472,N_19930);
nand UO_395 (O_395,N_19477,N_19756);
nand UO_396 (O_396,N_19617,N_19624);
nor UO_397 (O_397,N_19968,N_19446);
and UO_398 (O_398,N_19859,N_19418);
nor UO_399 (O_399,N_19565,N_19372);
nor UO_400 (O_400,N_19381,N_19731);
xor UO_401 (O_401,N_19202,N_19410);
xor UO_402 (O_402,N_19973,N_19724);
and UO_403 (O_403,N_19697,N_19302);
nand UO_404 (O_404,N_19260,N_19869);
xor UO_405 (O_405,N_19487,N_19231);
or UO_406 (O_406,N_19245,N_19959);
nand UO_407 (O_407,N_19261,N_19769);
nor UO_408 (O_408,N_19215,N_19547);
nor UO_409 (O_409,N_19396,N_19583);
or UO_410 (O_410,N_19599,N_19991);
xor UO_411 (O_411,N_19864,N_19388);
nor UO_412 (O_412,N_19407,N_19253);
and UO_413 (O_413,N_19680,N_19982);
xor UO_414 (O_414,N_19286,N_19338);
nand UO_415 (O_415,N_19981,N_19491);
and UO_416 (O_416,N_19979,N_19770);
nand UO_417 (O_417,N_19264,N_19616);
and UO_418 (O_418,N_19372,N_19643);
nor UO_419 (O_419,N_19342,N_19651);
xnor UO_420 (O_420,N_19322,N_19245);
or UO_421 (O_421,N_19413,N_19664);
xor UO_422 (O_422,N_19608,N_19561);
nor UO_423 (O_423,N_19444,N_19916);
nor UO_424 (O_424,N_19398,N_19682);
or UO_425 (O_425,N_19894,N_19530);
nor UO_426 (O_426,N_19677,N_19530);
and UO_427 (O_427,N_19244,N_19946);
or UO_428 (O_428,N_19620,N_19515);
or UO_429 (O_429,N_19476,N_19202);
and UO_430 (O_430,N_19301,N_19407);
nor UO_431 (O_431,N_19566,N_19609);
or UO_432 (O_432,N_19848,N_19551);
xnor UO_433 (O_433,N_19781,N_19418);
xnor UO_434 (O_434,N_19391,N_19286);
or UO_435 (O_435,N_19474,N_19892);
or UO_436 (O_436,N_19635,N_19259);
and UO_437 (O_437,N_19914,N_19968);
or UO_438 (O_438,N_19299,N_19517);
or UO_439 (O_439,N_19619,N_19828);
or UO_440 (O_440,N_19206,N_19231);
xnor UO_441 (O_441,N_19989,N_19696);
and UO_442 (O_442,N_19568,N_19204);
nor UO_443 (O_443,N_19568,N_19471);
and UO_444 (O_444,N_19497,N_19893);
nand UO_445 (O_445,N_19274,N_19735);
nand UO_446 (O_446,N_19467,N_19863);
or UO_447 (O_447,N_19213,N_19814);
and UO_448 (O_448,N_19223,N_19881);
xor UO_449 (O_449,N_19344,N_19594);
nand UO_450 (O_450,N_19436,N_19229);
and UO_451 (O_451,N_19851,N_19341);
nor UO_452 (O_452,N_19558,N_19979);
or UO_453 (O_453,N_19726,N_19386);
and UO_454 (O_454,N_19420,N_19646);
xnor UO_455 (O_455,N_19401,N_19485);
or UO_456 (O_456,N_19878,N_19712);
nor UO_457 (O_457,N_19372,N_19645);
xor UO_458 (O_458,N_19210,N_19731);
nor UO_459 (O_459,N_19448,N_19638);
nor UO_460 (O_460,N_19251,N_19248);
and UO_461 (O_461,N_19499,N_19594);
xnor UO_462 (O_462,N_19265,N_19340);
nand UO_463 (O_463,N_19577,N_19587);
and UO_464 (O_464,N_19614,N_19868);
or UO_465 (O_465,N_19210,N_19978);
and UO_466 (O_466,N_19810,N_19916);
nand UO_467 (O_467,N_19966,N_19857);
nor UO_468 (O_468,N_19571,N_19231);
xnor UO_469 (O_469,N_19525,N_19921);
xnor UO_470 (O_470,N_19273,N_19790);
nand UO_471 (O_471,N_19903,N_19972);
and UO_472 (O_472,N_19575,N_19231);
or UO_473 (O_473,N_19954,N_19838);
xnor UO_474 (O_474,N_19929,N_19708);
nand UO_475 (O_475,N_19351,N_19704);
and UO_476 (O_476,N_19900,N_19359);
or UO_477 (O_477,N_19942,N_19601);
and UO_478 (O_478,N_19523,N_19967);
and UO_479 (O_479,N_19778,N_19379);
nor UO_480 (O_480,N_19554,N_19253);
nor UO_481 (O_481,N_19548,N_19315);
or UO_482 (O_482,N_19369,N_19218);
xnor UO_483 (O_483,N_19783,N_19317);
xnor UO_484 (O_484,N_19609,N_19628);
or UO_485 (O_485,N_19859,N_19497);
xnor UO_486 (O_486,N_19565,N_19240);
or UO_487 (O_487,N_19370,N_19933);
xor UO_488 (O_488,N_19783,N_19496);
xnor UO_489 (O_489,N_19229,N_19216);
xor UO_490 (O_490,N_19343,N_19666);
nor UO_491 (O_491,N_19417,N_19218);
or UO_492 (O_492,N_19243,N_19832);
xnor UO_493 (O_493,N_19665,N_19246);
nor UO_494 (O_494,N_19878,N_19937);
and UO_495 (O_495,N_19878,N_19900);
xnor UO_496 (O_496,N_19521,N_19510);
or UO_497 (O_497,N_19531,N_19352);
and UO_498 (O_498,N_19814,N_19668);
or UO_499 (O_499,N_19240,N_19306);
nand UO_500 (O_500,N_19879,N_19542);
and UO_501 (O_501,N_19755,N_19390);
nand UO_502 (O_502,N_19814,N_19841);
xor UO_503 (O_503,N_19538,N_19828);
nand UO_504 (O_504,N_19706,N_19992);
xnor UO_505 (O_505,N_19557,N_19551);
nor UO_506 (O_506,N_19606,N_19962);
or UO_507 (O_507,N_19856,N_19357);
nor UO_508 (O_508,N_19829,N_19725);
xnor UO_509 (O_509,N_19451,N_19610);
xor UO_510 (O_510,N_19962,N_19974);
nor UO_511 (O_511,N_19416,N_19539);
nor UO_512 (O_512,N_19315,N_19322);
xor UO_513 (O_513,N_19881,N_19930);
nand UO_514 (O_514,N_19523,N_19438);
or UO_515 (O_515,N_19735,N_19473);
nor UO_516 (O_516,N_19424,N_19627);
xor UO_517 (O_517,N_19231,N_19314);
xnor UO_518 (O_518,N_19524,N_19491);
nand UO_519 (O_519,N_19670,N_19875);
or UO_520 (O_520,N_19498,N_19663);
nand UO_521 (O_521,N_19911,N_19372);
nand UO_522 (O_522,N_19383,N_19880);
nor UO_523 (O_523,N_19998,N_19577);
and UO_524 (O_524,N_19414,N_19327);
and UO_525 (O_525,N_19262,N_19932);
nor UO_526 (O_526,N_19561,N_19823);
nand UO_527 (O_527,N_19672,N_19443);
and UO_528 (O_528,N_19937,N_19255);
nand UO_529 (O_529,N_19770,N_19389);
or UO_530 (O_530,N_19619,N_19348);
nand UO_531 (O_531,N_19727,N_19327);
or UO_532 (O_532,N_19653,N_19753);
xor UO_533 (O_533,N_19811,N_19659);
and UO_534 (O_534,N_19232,N_19319);
or UO_535 (O_535,N_19213,N_19570);
nor UO_536 (O_536,N_19874,N_19895);
nand UO_537 (O_537,N_19680,N_19718);
and UO_538 (O_538,N_19342,N_19896);
or UO_539 (O_539,N_19735,N_19598);
and UO_540 (O_540,N_19447,N_19704);
nand UO_541 (O_541,N_19574,N_19890);
or UO_542 (O_542,N_19832,N_19965);
and UO_543 (O_543,N_19770,N_19531);
xor UO_544 (O_544,N_19260,N_19576);
nand UO_545 (O_545,N_19490,N_19851);
nor UO_546 (O_546,N_19988,N_19535);
and UO_547 (O_547,N_19674,N_19534);
or UO_548 (O_548,N_19407,N_19373);
and UO_549 (O_549,N_19328,N_19481);
or UO_550 (O_550,N_19926,N_19916);
xor UO_551 (O_551,N_19461,N_19255);
or UO_552 (O_552,N_19940,N_19795);
or UO_553 (O_553,N_19696,N_19214);
and UO_554 (O_554,N_19825,N_19896);
or UO_555 (O_555,N_19418,N_19953);
xnor UO_556 (O_556,N_19583,N_19457);
and UO_557 (O_557,N_19550,N_19969);
or UO_558 (O_558,N_19992,N_19879);
and UO_559 (O_559,N_19744,N_19948);
and UO_560 (O_560,N_19239,N_19978);
or UO_561 (O_561,N_19801,N_19372);
and UO_562 (O_562,N_19452,N_19998);
or UO_563 (O_563,N_19340,N_19968);
and UO_564 (O_564,N_19345,N_19566);
nand UO_565 (O_565,N_19992,N_19750);
or UO_566 (O_566,N_19245,N_19608);
or UO_567 (O_567,N_19501,N_19540);
nor UO_568 (O_568,N_19414,N_19315);
and UO_569 (O_569,N_19792,N_19538);
nand UO_570 (O_570,N_19874,N_19213);
nor UO_571 (O_571,N_19330,N_19534);
nor UO_572 (O_572,N_19405,N_19557);
nand UO_573 (O_573,N_19612,N_19477);
or UO_574 (O_574,N_19523,N_19990);
nand UO_575 (O_575,N_19873,N_19909);
nor UO_576 (O_576,N_19365,N_19453);
and UO_577 (O_577,N_19305,N_19746);
nand UO_578 (O_578,N_19462,N_19561);
or UO_579 (O_579,N_19787,N_19348);
and UO_580 (O_580,N_19799,N_19748);
and UO_581 (O_581,N_19235,N_19310);
nor UO_582 (O_582,N_19971,N_19954);
xor UO_583 (O_583,N_19293,N_19275);
and UO_584 (O_584,N_19494,N_19205);
or UO_585 (O_585,N_19929,N_19487);
nand UO_586 (O_586,N_19605,N_19482);
nand UO_587 (O_587,N_19476,N_19334);
nor UO_588 (O_588,N_19927,N_19470);
or UO_589 (O_589,N_19733,N_19825);
nand UO_590 (O_590,N_19713,N_19710);
nor UO_591 (O_591,N_19374,N_19287);
or UO_592 (O_592,N_19710,N_19519);
nand UO_593 (O_593,N_19907,N_19237);
xor UO_594 (O_594,N_19510,N_19853);
xor UO_595 (O_595,N_19524,N_19997);
nor UO_596 (O_596,N_19209,N_19524);
nor UO_597 (O_597,N_19549,N_19672);
xnor UO_598 (O_598,N_19727,N_19489);
and UO_599 (O_599,N_19504,N_19604);
nor UO_600 (O_600,N_19205,N_19816);
nor UO_601 (O_601,N_19905,N_19832);
and UO_602 (O_602,N_19502,N_19737);
and UO_603 (O_603,N_19725,N_19286);
nand UO_604 (O_604,N_19406,N_19253);
xor UO_605 (O_605,N_19929,N_19646);
and UO_606 (O_606,N_19700,N_19695);
nand UO_607 (O_607,N_19350,N_19766);
nor UO_608 (O_608,N_19802,N_19690);
or UO_609 (O_609,N_19950,N_19458);
nand UO_610 (O_610,N_19488,N_19271);
and UO_611 (O_611,N_19368,N_19310);
xor UO_612 (O_612,N_19989,N_19574);
nand UO_613 (O_613,N_19879,N_19702);
or UO_614 (O_614,N_19552,N_19485);
xor UO_615 (O_615,N_19298,N_19459);
nand UO_616 (O_616,N_19842,N_19535);
nand UO_617 (O_617,N_19730,N_19939);
or UO_618 (O_618,N_19779,N_19390);
and UO_619 (O_619,N_19413,N_19344);
and UO_620 (O_620,N_19711,N_19412);
nand UO_621 (O_621,N_19524,N_19782);
nor UO_622 (O_622,N_19605,N_19965);
nor UO_623 (O_623,N_19678,N_19772);
xor UO_624 (O_624,N_19261,N_19427);
or UO_625 (O_625,N_19742,N_19843);
or UO_626 (O_626,N_19423,N_19661);
or UO_627 (O_627,N_19325,N_19644);
nand UO_628 (O_628,N_19667,N_19624);
and UO_629 (O_629,N_19660,N_19609);
nand UO_630 (O_630,N_19818,N_19981);
nor UO_631 (O_631,N_19632,N_19668);
xnor UO_632 (O_632,N_19985,N_19764);
nand UO_633 (O_633,N_19454,N_19632);
nand UO_634 (O_634,N_19525,N_19463);
and UO_635 (O_635,N_19589,N_19288);
nand UO_636 (O_636,N_19449,N_19589);
xor UO_637 (O_637,N_19683,N_19639);
and UO_638 (O_638,N_19995,N_19899);
xnor UO_639 (O_639,N_19811,N_19763);
nor UO_640 (O_640,N_19292,N_19542);
and UO_641 (O_641,N_19613,N_19867);
and UO_642 (O_642,N_19822,N_19724);
xnor UO_643 (O_643,N_19988,N_19731);
and UO_644 (O_644,N_19736,N_19743);
xnor UO_645 (O_645,N_19619,N_19302);
or UO_646 (O_646,N_19671,N_19349);
nand UO_647 (O_647,N_19609,N_19282);
nand UO_648 (O_648,N_19706,N_19235);
nor UO_649 (O_649,N_19980,N_19631);
xnor UO_650 (O_650,N_19588,N_19596);
nor UO_651 (O_651,N_19261,N_19551);
nand UO_652 (O_652,N_19487,N_19308);
xnor UO_653 (O_653,N_19649,N_19679);
nor UO_654 (O_654,N_19770,N_19206);
and UO_655 (O_655,N_19405,N_19611);
nand UO_656 (O_656,N_19290,N_19467);
nor UO_657 (O_657,N_19202,N_19511);
nor UO_658 (O_658,N_19910,N_19296);
nand UO_659 (O_659,N_19614,N_19560);
and UO_660 (O_660,N_19935,N_19310);
and UO_661 (O_661,N_19877,N_19712);
nand UO_662 (O_662,N_19658,N_19835);
nand UO_663 (O_663,N_19486,N_19829);
nand UO_664 (O_664,N_19735,N_19211);
nand UO_665 (O_665,N_19879,N_19425);
xnor UO_666 (O_666,N_19776,N_19248);
xor UO_667 (O_667,N_19930,N_19997);
nor UO_668 (O_668,N_19909,N_19944);
xnor UO_669 (O_669,N_19538,N_19912);
xnor UO_670 (O_670,N_19460,N_19586);
or UO_671 (O_671,N_19364,N_19350);
xnor UO_672 (O_672,N_19658,N_19268);
nand UO_673 (O_673,N_19566,N_19316);
xnor UO_674 (O_674,N_19292,N_19449);
or UO_675 (O_675,N_19529,N_19906);
and UO_676 (O_676,N_19446,N_19689);
nor UO_677 (O_677,N_19720,N_19292);
xor UO_678 (O_678,N_19234,N_19912);
xor UO_679 (O_679,N_19733,N_19756);
xnor UO_680 (O_680,N_19274,N_19319);
nand UO_681 (O_681,N_19387,N_19822);
nor UO_682 (O_682,N_19681,N_19817);
or UO_683 (O_683,N_19580,N_19300);
and UO_684 (O_684,N_19205,N_19322);
nor UO_685 (O_685,N_19455,N_19413);
xor UO_686 (O_686,N_19502,N_19906);
xnor UO_687 (O_687,N_19256,N_19334);
and UO_688 (O_688,N_19633,N_19917);
nor UO_689 (O_689,N_19439,N_19637);
or UO_690 (O_690,N_19771,N_19554);
nand UO_691 (O_691,N_19572,N_19991);
and UO_692 (O_692,N_19695,N_19809);
xnor UO_693 (O_693,N_19421,N_19906);
or UO_694 (O_694,N_19978,N_19948);
xor UO_695 (O_695,N_19249,N_19731);
or UO_696 (O_696,N_19478,N_19706);
and UO_697 (O_697,N_19352,N_19375);
xnor UO_698 (O_698,N_19419,N_19386);
xnor UO_699 (O_699,N_19935,N_19907);
and UO_700 (O_700,N_19409,N_19786);
or UO_701 (O_701,N_19277,N_19548);
nand UO_702 (O_702,N_19225,N_19873);
nor UO_703 (O_703,N_19818,N_19740);
nand UO_704 (O_704,N_19521,N_19667);
or UO_705 (O_705,N_19628,N_19469);
nor UO_706 (O_706,N_19732,N_19476);
and UO_707 (O_707,N_19267,N_19740);
and UO_708 (O_708,N_19376,N_19289);
nand UO_709 (O_709,N_19480,N_19220);
and UO_710 (O_710,N_19212,N_19576);
or UO_711 (O_711,N_19906,N_19584);
and UO_712 (O_712,N_19978,N_19853);
xor UO_713 (O_713,N_19259,N_19785);
and UO_714 (O_714,N_19501,N_19545);
or UO_715 (O_715,N_19759,N_19257);
nand UO_716 (O_716,N_19365,N_19344);
or UO_717 (O_717,N_19635,N_19320);
or UO_718 (O_718,N_19979,N_19917);
nand UO_719 (O_719,N_19215,N_19396);
nor UO_720 (O_720,N_19642,N_19652);
and UO_721 (O_721,N_19327,N_19361);
or UO_722 (O_722,N_19311,N_19553);
nor UO_723 (O_723,N_19657,N_19826);
and UO_724 (O_724,N_19994,N_19536);
xnor UO_725 (O_725,N_19865,N_19948);
xnor UO_726 (O_726,N_19832,N_19461);
nor UO_727 (O_727,N_19373,N_19746);
nand UO_728 (O_728,N_19925,N_19543);
and UO_729 (O_729,N_19617,N_19743);
nand UO_730 (O_730,N_19316,N_19419);
and UO_731 (O_731,N_19761,N_19721);
xnor UO_732 (O_732,N_19675,N_19947);
nand UO_733 (O_733,N_19431,N_19421);
xor UO_734 (O_734,N_19353,N_19235);
nor UO_735 (O_735,N_19375,N_19236);
nor UO_736 (O_736,N_19330,N_19669);
and UO_737 (O_737,N_19997,N_19891);
and UO_738 (O_738,N_19340,N_19235);
nor UO_739 (O_739,N_19551,N_19683);
or UO_740 (O_740,N_19789,N_19666);
nor UO_741 (O_741,N_19791,N_19357);
nor UO_742 (O_742,N_19493,N_19842);
or UO_743 (O_743,N_19223,N_19889);
and UO_744 (O_744,N_19262,N_19674);
and UO_745 (O_745,N_19591,N_19658);
xnor UO_746 (O_746,N_19348,N_19606);
or UO_747 (O_747,N_19405,N_19403);
or UO_748 (O_748,N_19481,N_19415);
and UO_749 (O_749,N_19485,N_19484);
or UO_750 (O_750,N_19716,N_19397);
nor UO_751 (O_751,N_19669,N_19684);
and UO_752 (O_752,N_19507,N_19428);
nor UO_753 (O_753,N_19881,N_19498);
or UO_754 (O_754,N_19316,N_19722);
nor UO_755 (O_755,N_19782,N_19631);
or UO_756 (O_756,N_19443,N_19259);
nor UO_757 (O_757,N_19605,N_19580);
and UO_758 (O_758,N_19870,N_19489);
and UO_759 (O_759,N_19567,N_19910);
and UO_760 (O_760,N_19811,N_19728);
or UO_761 (O_761,N_19908,N_19456);
or UO_762 (O_762,N_19449,N_19428);
or UO_763 (O_763,N_19904,N_19330);
nor UO_764 (O_764,N_19761,N_19491);
nand UO_765 (O_765,N_19370,N_19716);
xnor UO_766 (O_766,N_19462,N_19695);
and UO_767 (O_767,N_19981,N_19681);
nor UO_768 (O_768,N_19557,N_19646);
xnor UO_769 (O_769,N_19333,N_19429);
nand UO_770 (O_770,N_19879,N_19641);
and UO_771 (O_771,N_19250,N_19669);
nand UO_772 (O_772,N_19366,N_19362);
or UO_773 (O_773,N_19846,N_19298);
nor UO_774 (O_774,N_19599,N_19860);
nand UO_775 (O_775,N_19912,N_19574);
and UO_776 (O_776,N_19892,N_19907);
xnor UO_777 (O_777,N_19291,N_19970);
nand UO_778 (O_778,N_19634,N_19827);
nor UO_779 (O_779,N_19889,N_19340);
nor UO_780 (O_780,N_19299,N_19642);
xnor UO_781 (O_781,N_19251,N_19873);
xnor UO_782 (O_782,N_19345,N_19993);
xor UO_783 (O_783,N_19216,N_19291);
nor UO_784 (O_784,N_19903,N_19496);
or UO_785 (O_785,N_19203,N_19700);
nor UO_786 (O_786,N_19364,N_19374);
and UO_787 (O_787,N_19976,N_19331);
xnor UO_788 (O_788,N_19217,N_19450);
and UO_789 (O_789,N_19204,N_19878);
nand UO_790 (O_790,N_19241,N_19473);
and UO_791 (O_791,N_19377,N_19948);
xnor UO_792 (O_792,N_19438,N_19809);
or UO_793 (O_793,N_19343,N_19730);
nor UO_794 (O_794,N_19297,N_19632);
nor UO_795 (O_795,N_19920,N_19581);
xor UO_796 (O_796,N_19584,N_19478);
nand UO_797 (O_797,N_19345,N_19228);
xnor UO_798 (O_798,N_19394,N_19938);
xor UO_799 (O_799,N_19289,N_19406);
nand UO_800 (O_800,N_19798,N_19530);
xor UO_801 (O_801,N_19580,N_19205);
xor UO_802 (O_802,N_19275,N_19299);
and UO_803 (O_803,N_19634,N_19924);
nand UO_804 (O_804,N_19625,N_19431);
nor UO_805 (O_805,N_19705,N_19346);
nor UO_806 (O_806,N_19486,N_19402);
xor UO_807 (O_807,N_19580,N_19641);
and UO_808 (O_808,N_19768,N_19725);
and UO_809 (O_809,N_19310,N_19801);
xor UO_810 (O_810,N_19810,N_19947);
nand UO_811 (O_811,N_19311,N_19744);
nor UO_812 (O_812,N_19915,N_19290);
nor UO_813 (O_813,N_19379,N_19608);
nor UO_814 (O_814,N_19627,N_19915);
and UO_815 (O_815,N_19943,N_19746);
xnor UO_816 (O_816,N_19470,N_19365);
or UO_817 (O_817,N_19978,N_19355);
nor UO_818 (O_818,N_19709,N_19575);
xor UO_819 (O_819,N_19573,N_19649);
and UO_820 (O_820,N_19580,N_19573);
xnor UO_821 (O_821,N_19918,N_19920);
nor UO_822 (O_822,N_19823,N_19578);
nand UO_823 (O_823,N_19792,N_19523);
or UO_824 (O_824,N_19783,N_19895);
nand UO_825 (O_825,N_19842,N_19550);
or UO_826 (O_826,N_19577,N_19578);
nand UO_827 (O_827,N_19502,N_19645);
nand UO_828 (O_828,N_19784,N_19295);
nand UO_829 (O_829,N_19550,N_19739);
nor UO_830 (O_830,N_19739,N_19229);
nor UO_831 (O_831,N_19606,N_19299);
nor UO_832 (O_832,N_19650,N_19246);
nand UO_833 (O_833,N_19590,N_19531);
xnor UO_834 (O_834,N_19462,N_19772);
and UO_835 (O_835,N_19285,N_19528);
nor UO_836 (O_836,N_19829,N_19340);
and UO_837 (O_837,N_19482,N_19581);
or UO_838 (O_838,N_19864,N_19678);
nor UO_839 (O_839,N_19837,N_19442);
or UO_840 (O_840,N_19876,N_19227);
xnor UO_841 (O_841,N_19661,N_19455);
and UO_842 (O_842,N_19977,N_19716);
or UO_843 (O_843,N_19566,N_19239);
or UO_844 (O_844,N_19374,N_19778);
and UO_845 (O_845,N_19251,N_19221);
nand UO_846 (O_846,N_19566,N_19724);
nor UO_847 (O_847,N_19864,N_19553);
nor UO_848 (O_848,N_19764,N_19285);
xor UO_849 (O_849,N_19437,N_19927);
nand UO_850 (O_850,N_19237,N_19690);
and UO_851 (O_851,N_19577,N_19341);
nor UO_852 (O_852,N_19461,N_19478);
nand UO_853 (O_853,N_19772,N_19872);
and UO_854 (O_854,N_19924,N_19224);
and UO_855 (O_855,N_19498,N_19604);
xor UO_856 (O_856,N_19534,N_19888);
or UO_857 (O_857,N_19393,N_19228);
or UO_858 (O_858,N_19894,N_19891);
nand UO_859 (O_859,N_19433,N_19600);
nand UO_860 (O_860,N_19953,N_19978);
xor UO_861 (O_861,N_19481,N_19253);
and UO_862 (O_862,N_19358,N_19584);
and UO_863 (O_863,N_19406,N_19285);
or UO_864 (O_864,N_19202,N_19695);
xor UO_865 (O_865,N_19252,N_19961);
xnor UO_866 (O_866,N_19561,N_19877);
xnor UO_867 (O_867,N_19441,N_19605);
or UO_868 (O_868,N_19868,N_19538);
nand UO_869 (O_869,N_19515,N_19800);
or UO_870 (O_870,N_19793,N_19286);
or UO_871 (O_871,N_19445,N_19614);
xnor UO_872 (O_872,N_19858,N_19667);
and UO_873 (O_873,N_19903,N_19576);
xor UO_874 (O_874,N_19259,N_19750);
or UO_875 (O_875,N_19433,N_19294);
and UO_876 (O_876,N_19411,N_19690);
nor UO_877 (O_877,N_19612,N_19601);
xor UO_878 (O_878,N_19932,N_19864);
and UO_879 (O_879,N_19494,N_19897);
nand UO_880 (O_880,N_19238,N_19501);
xor UO_881 (O_881,N_19590,N_19657);
and UO_882 (O_882,N_19372,N_19539);
xnor UO_883 (O_883,N_19743,N_19460);
and UO_884 (O_884,N_19690,N_19621);
nor UO_885 (O_885,N_19955,N_19243);
nand UO_886 (O_886,N_19524,N_19656);
nor UO_887 (O_887,N_19344,N_19661);
nor UO_888 (O_888,N_19263,N_19967);
nor UO_889 (O_889,N_19487,N_19881);
xnor UO_890 (O_890,N_19360,N_19238);
and UO_891 (O_891,N_19292,N_19374);
nand UO_892 (O_892,N_19280,N_19861);
xor UO_893 (O_893,N_19204,N_19419);
and UO_894 (O_894,N_19203,N_19785);
xnor UO_895 (O_895,N_19765,N_19460);
nor UO_896 (O_896,N_19493,N_19958);
or UO_897 (O_897,N_19537,N_19557);
nor UO_898 (O_898,N_19489,N_19461);
xnor UO_899 (O_899,N_19306,N_19840);
xnor UO_900 (O_900,N_19731,N_19766);
xnor UO_901 (O_901,N_19351,N_19819);
nand UO_902 (O_902,N_19582,N_19631);
and UO_903 (O_903,N_19793,N_19928);
nor UO_904 (O_904,N_19771,N_19827);
or UO_905 (O_905,N_19903,N_19966);
nor UO_906 (O_906,N_19850,N_19570);
or UO_907 (O_907,N_19524,N_19536);
and UO_908 (O_908,N_19489,N_19562);
or UO_909 (O_909,N_19645,N_19781);
and UO_910 (O_910,N_19458,N_19670);
or UO_911 (O_911,N_19930,N_19336);
or UO_912 (O_912,N_19520,N_19571);
xor UO_913 (O_913,N_19639,N_19943);
and UO_914 (O_914,N_19726,N_19648);
nor UO_915 (O_915,N_19304,N_19666);
nand UO_916 (O_916,N_19219,N_19236);
or UO_917 (O_917,N_19611,N_19551);
xor UO_918 (O_918,N_19727,N_19495);
nor UO_919 (O_919,N_19856,N_19941);
or UO_920 (O_920,N_19603,N_19742);
and UO_921 (O_921,N_19476,N_19213);
nor UO_922 (O_922,N_19333,N_19553);
and UO_923 (O_923,N_19244,N_19684);
nand UO_924 (O_924,N_19559,N_19729);
or UO_925 (O_925,N_19670,N_19869);
nand UO_926 (O_926,N_19233,N_19477);
nor UO_927 (O_927,N_19761,N_19760);
or UO_928 (O_928,N_19732,N_19200);
and UO_929 (O_929,N_19909,N_19363);
nor UO_930 (O_930,N_19609,N_19230);
and UO_931 (O_931,N_19669,N_19549);
and UO_932 (O_932,N_19988,N_19657);
or UO_933 (O_933,N_19269,N_19829);
or UO_934 (O_934,N_19912,N_19670);
or UO_935 (O_935,N_19287,N_19756);
nor UO_936 (O_936,N_19885,N_19612);
nor UO_937 (O_937,N_19624,N_19729);
xnor UO_938 (O_938,N_19754,N_19562);
nand UO_939 (O_939,N_19913,N_19888);
and UO_940 (O_940,N_19250,N_19891);
and UO_941 (O_941,N_19319,N_19558);
and UO_942 (O_942,N_19848,N_19399);
nand UO_943 (O_943,N_19838,N_19966);
or UO_944 (O_944,N_19731,N_19801);
and UO_945 (O_945,N_19807,N_19626);
nor UO_946 (O_946,N_19264,N_19223);
nor UO_947 (O_947,N_19993,N_19438);
and UO_948 (O_948,N_19687,N_19378);
nor UO_949 (O_949,N_19981,N_19481);
nand UO_950 (O_950,N_19525,N_19568);
nand UO_951 (O_951,N_19817,N_19262);
nor UO_952 (O_952,N_19333,N_19863);
xnor UO_953 (O_953,N_19832,N_19930);
nand UO_954 (O_954,N_19692,N_19819);
xor UO_955 (O_955,N_19391,N_19441);
or UO_956 (O_956,N_19716,N_19502);
or UO_957 (O_957,N_19422,N_19354);
xnor UO_958 (O_958,N_19223,N_19909);
or UO_959 (O_959,N_19594,N_19313);
and UO_960 (O_960,N_19877,N_19724);
xnor UO_961 (O_961,N_19832,N_19609);
nand UO_962 (O_962,N_19559,N_19624);
or UO_963 (O_963,N_19256,N_19290);
nand UO_964 (O_964,N_19371,N_19569);
nand UO_965 (O_965,N_19209,N_19396);
or UO_966 (O_966,N_19782,N_19287);
and UO_967 (O_967,N_19328,N_19615);
xnor UO_968 (O_968,N_19868,N_19949);
and UO_969 (O_969,N_19270,N_19434);
or UO_970 (O_970,N_19584,N_19690);
or UO_971 (O_971,N_19851,N_19995);
nand UO_972 (O_972,N_19938,N_19833);
nor UO_973 (O_973,N_19481,N_19496);
nor UO_974 (O_974,N_19862,N_19986);
or UO_975 (O_975,N_19417,N_19219);
xnor UO_976 (O_976,N_19623,N_19806);
xnor UO_977 (O_977,N_19496,N_19385);
and UO_978 (O_978,N_19649,N_19968);
and UO_979 (O_979,N_19827,N_19447);
nor UO_980 (O_980,N_19693,N_19821);
nor UO_981 (O_981,N_19931,N_19370);
nand UO_982 (O_982,N_19813,N_19960);
nand UO_983 (O_983,N_19711,N_19319);
and UO_984 (O_984,N_19811,N_19502);
xor UO_985 (O_985,N_19623,N_19943);
or UO_986 (O_986,N_19975,N_19293);
or UO_987 (O_987,N_19536,N_19543);
nor UO_988 (O_988,N_19691,N_19954);
and UO_989 (O_989,N_19429,N_19366);
nand UO_990 (O_990,N_19361,N_19493);
and UO_991 (O_991,N_19971,N_19484);
and UO_992 (O_992,N_19853,N_19805);
and UO_993 (O_993,N_19934,N_19927);
or UO_994 (O_994,N_19288,N_19984);
or UO_995 (O_995,N_19502,N_19385);
nand UO_996 (O_996,N_19318,N_19695);
or UO_997 (O_997,N_19202,N_19844);
nand UO_998 (O_998,N_19454,N_19200);
nor UO_999 (O_999,N_19358,N_19745);
nand UO_1000 (O_1000,N_19766,N_19833);
nand UO_1001 (O_1001,N_19742,N_19237);
nor UO_1002 (O_1002,N_19752,N_19383);
and UO_1003 (O_1003,N_19900,N_19344);
nand UO_1004 (O_1004,N_19575,N_19561);
or UO_1005 (O_1005,N_19485,N_19743);
nand UO_1006 (O_1006,N_19402,N_19622);
nand UO_1007 (O_1007,N_19534,N_19334);
xnor UO_1008 (O_1008,N_19588,N_19639);
nor UO_1009 (O_1009,N_19983,N_19793);
nor UO_1010 (O_1010,N_19735,N_19718);
nor UO_1011 (O_1011,N_19836,N_19984);
xnor UO_1012 (O_1012,N_19329,N_19919);
nor UO_1013 (O_1013,N_19382,N_19405);
nor UO_1014 (O_1014,N_19960,N_19698);
nor UO_1015 (O_1015,N_19965,N_19376);
and UO_1016 (O_1016,N_19710,N_19772);
and UO_1017 (O_1017,N_19688,N_19548);
nand UO_1018 (O_1018,N_19300,N_19676);
and UO_1019 (O_1019,N_19464,N_19568);
or UO_1020 (O_1020,N_19805,N_19712);
xnor UO_1021 (O_1021,N_19334,N_19540);
xnor UO_1022 (O_1022,N_19692,N_19589);
nor UO_1023 (O_1023,N_19307,N_19391);
and UO_1024 (O_1024,N_19860,N_19256);
and UO_1025 (O_1025,N_19641,N_19935);
nor UO_1026 (O_1026,N_19528,N_19886);
nor UO_1027 (O_1027,N_19805,N_19979);
nand UO_1028 (O_1028,N_19563,N_19341);
nor UO_1029 (O_1029,N_19588,N_19262);
xnor UO_1030 (O_1030,N_19715,N_19306);
nand UO_1031 (O_1031,N_19267,N_19959);
xnor UO_1032 (O_1032,N_19965,N_19799);
nand UO_1033 (O_1033,N_19379,N_19277);
nor UO_1034 (O_1034,N_19912,N_19896);
and UO_1035 (O_1035,N_19908,N_19581);
nor UO_1036 (O_1036,N_19704,N_19603);
nand UO_1037 (O_1037,N_19472,N_19550);
nor UO_1038 (O_1038,N_19628,N_19407);
nand UO_1039 (O_1039,N_19326,N_19724);
and UO_1040 (O_1040,N_19783,N_19911);
xor UO_1041 (O_1041,N_19689,N_19225);
or UO_1042 (O_1042,N_19298,N_19376);
nor UO_1043 (O_1043,N_19807,N_19478);
and UO_1044 (O_1044,N_19839,N_19657);
nor UO_1045 (O_1045,N_19766,N_19940);
and UO_1046 (O_1046,N_19809,N_19650);
or UO_1047 (O_1047,N_19827,N_19531);
xnor UO_1048 (O_1048,N_19454,N_19432);
xor UO_1049 (O_1049,N_19207,N_19383);
and UO_1050 (O_1050,N_19232,N_19831);
xnor UO_1051 (O_1051,N_19391,N_19295);
nand UO_1052 (O_1052,N_19335,N_19275);
or UO_1053 (O_1053,N_19396,N_19909);
xnor UO_1054 (O_1054,N_19866,N_19509);
nor UO_1055 (O_1055,N_19745,N_19254);
xor UO_1056 (O_1056,N_19237,N_19867);
xnor UO_1057 (O_1057,N_19300,N_19320);
nor UO_1058 (O_1058,N_19759,N_19812);
or UO_1059 (O_1059,N_19834,N_19829);
nand UO_1060 (O_1060,N_19886,N_19720);
and UO_1061 (O_1061,N_19879,N_19334);
xor UO_1062 (O_1062,N_19806,N_19543);
or UO_1063 (O_1063,N_19580,N_19335);
nand UO_1064 (O_1064,N_19889,N_19500);
or UO_1065 (O_1065,N_19694,N_19232);
nand UO_1066 (O_1066,N_19391,N_19401);
or UO_1067 (O_1067,N_19573,N_19862);
xnor UO_1068 (O_1068,N_19875,N_19553);
xor UO_1069 (O_1069,N_19320,N_19930);
xnor UO_1070 (O_1070,N_19710,N_19338);
nor UO_1071 (O_1071,N_19729,N_19839);
nand UO_1072 (O_1072,N_19750,N_19577);
nand UO_1073 (O_1073,N_19807,N_19438);
and UO_1074 (O_1074,N_19843,N_19607);
nand UO_1075 (O_1075,N_19212,N_19409);
and UO_1076 (O_1076,N_19274,N_19688);
or UO_1077 (O_1077,N_19860,N_19793);
nand UO_1078 (O_1078,N_19744,N_19786);
or UO_1079 (O_1079,N_19359,N_19565);
and UO_1080 (O_1080,N_19535,N_19925);
or UO_1081 (O_1081,N_19764,N_19870);
nand UO_1082 (O_1082,N_19956,N_19363);
or UO_1083 (O_1083,N_19900,N_19601);
xor UO_1084 (O_1084,N_19550,N_19424);
and UO_1085 (O_1085,N_19721,N_19299);
nand UO_1086 (O_1086,N_19874,N_19720);
nor UO_1087 (O_1087,N_19569,N_19330);
nand UO_1088 (O_1088,N_19305,N_19920);
nand UO_1089 (O_1089,N_19698,N_19935);
xnor UO_1090 (O_1090,N_19712,N_19917);
nand UO_1091 (O_1091,N_19327,N_19585);
and UO_1092 (O_1092,N_19206,N_19454);
or UO_1093 (O_1093,N_19469,N_19283);
and UO_1094 (O_1094,N_19329,N_19451);
nand UO_1095 (O_1095,N_19813,N_19577);
nand UO_1096 (O_1096,N_19230,N_19613);
or UO_1097 (O_1097,N_19474,N_19734);
or UO_1098 (O_1098,N_19817,N_19476);
or UO_1099 (O_1099,N_19841,N_19782);
nor UO_1100 (O_1100,N_19815,N_19747);
nand UO_1101 (O_1101,N_19318,N_19624);
and UO_1102 (O_1102,N_19799,N_19497);
nor UO_1103 (O_1103,N_19526,N_19575);
nor UO_1104 (O_1104,N_19459,N_19503);
xnor UO_1105 (O_1105,N_19831,N_19541);
nand UO_1106 (O_1106,N_19540,N_19212);
xor UO_1107 (O_1107,N_19844,N_19965);
nand UO_1108 (O_1108,N_19592,N_19874);
or UO_1109 (O_1109,N_19399,N_19886);
and UO_1110 (O_1110,N_19455,N_19705);
xor UO_1111 (O_1111,N_19277,N_19209);
xnor UO_1112 (O_1112,N_19260,N_19434);
nor UO_1113 (O_1113,N_19674,N_19253);
and UO_1114 (O_1114,N_19859,N_19480);
nor UO_1115 (O_1115,N_19619,N_19396);
xnor UO_1116 (O_1116,N_19748,N_19441);
and UO_1117 (O_1117,N_19773,N_19328);
or UO_1118 (O_1118,N_19204,N_19609);
nand UO_1119 (O_1119,N_19251,N_19476);
nand UO_1120 (O_1120,N_19715,N_19869);
and UO_1121 (O_1121,N_19684,N_19984);
nor UO_1122 (O_1122,N_19222,N_19887);
nand UO_1123 (O_1123,N_19959,N_19698);
and UO_1124 (O_1124,N_19876,N_19236);
nor UO_1125 (O_1125,N_19314,N_19779);
nand UO_1126 (O_1126,N_19406,N_19792);
nor UO_1127 (O_1127,N_19570,N_19378);
nand UO_1128 (O_1128,N_19802,N_19774);
nand UO_1129 (O_1129,N_19595,N_19984);
xor UO_1130 (O_1130,N_19395,N_19926);
xor UO_1131 (O_1131,N_19438,N_19570);
xnor UO_1132 (O_1132,N_19371,N_19934);
xnor UO_1133 (O_1133,N_19788,N_19251);
nor UO_1134 (O_1134,N_19741,N_19917);
xor UO_1135 (O_1135,N_19255,N_19930);
xnor UO_1136 (O_1136,N_19400,N_19516);
nand UO_1137 (O_1137,N_19976,N_19395);
nor UO_1138 (O_1138,N_19717,N_19555);
or UO_1139 (O_1139,N_19720,N_19224);
nand UO_1140 (O_1140,N_19688,N_19896);
or UO_1141 (O_1141,N_19610,N_19965);
or UO_1142 (O_1142,N_19397,N_19509);
xor UO_1143 (O_1143,N_19538,N_19295);
xor UO_1144 (O_1144,N_19621,N_19634);
and UO_1145 (O_1145,N_19240,N_19597);
nor UO_1146 (O_1146,N_19655,N_19299);
xnor UO_1147 (O_1147,N_19430,N_19789);
and UO_1148 (O_1148,N_19391,N_19507);
and UO_1149 (O_1149,N_19850,N_19670);
nand UO_1150 (O_1150,N_19940,N_19466);
and UO_1151 (O_1151,N_19868,N_19549);
nand UO_1152 (O_1152,N_19927,N_19980);
and UO_1153 (O_1153,N_19812,N_19818);
nand UO_1154 (O_1154,N_19992,N_19908);
and UO_1155 (O_1155,N_19694,N_19749);
xor UO_1156 (O_1156,N_19444,N_19417);
nand UO_1157 (O_1157,N_19338,N_19738);
or UO_1158 (O_1158,N_19544,N_19480);
or UO_1159 (O_1159,N_19308,N_19407);
nand UO_1160 (O_1160,N_19660,N_19259);
and UO_1161 (O_1161,N_19373,N_19480);
and UO_1162 (O_1162,N_19439,N_19768);
or UO_1163 (O_1163,N_19966,N_19830);
or UO_1164 (O_1164,N_19237,N_19587);
and UO_1165 (O_1165,N_19992,N_19542);
nor UO_1166 (O_1166,N_19207,N_19735);
nor UO_1167 (O_1167,N_19399,N_19926);
or UO_1168 (O_1168,N_19898,N_19932);
nand UO_1169 (O_1169,N_19399,N_19703);
nor UO_1170 (O_1170,N_19453,N_19744);
and UO_1171 (O_1171,N_19231,N_19272);
or UO_1172 (O_1172,N_19585,N_19955);
xnor UO_1173 (O_1173,N_19970,N_19596);
nand UO_1174 (O_1174,N_19398,N_19555);
or UO_1175 (O_1175,N_19583,N_19604);
nand UO_1176 (O_1176,N_19276,N_19763);
xor UO_1177 (O_1177,N_19839,N_19643);
xor UO_1178 (O_1178,N_19857,N_19242);
nand UO_1179 (O_1179,N_19519,N_19621);
nand UO_1180 (O_1180,N_19588,N_19487);
xor UO_1181 (O_1181,N_19542,N_19594);
xnor UO_1182 (O_1182,N_19587,N_19939);
and UO_1183 (O_1183,N_19651,N_19737);
and UO_1184 (O_1184,N_19980,N_19525);
and UO_1185 (O_1185,N_19868,N_19285);
nor UO_1186 (O_1186,N_19314,N_19682);
xnor UO_1187 (O_1187,N_19608,N_19563);
and UO_1188 (O_1188,N_19623,N_19702);
and UO_1189 (O_1189,N_19473,N_19525);
nand UO_1190 (O_1190,N_19713,N_19765);
and UO_1191 (O_1191,N_19219,N_19545);
or UO_1192 (O_1192,N_19510,N_19377);
nor UO_1193 (O_1193,N_19210,N_19556);
nor UO_1194 (O_1194,N_19750,N_19266);
nand UO_1195 (O_1195,N_19526,N_19608);
nor UO_1196 (O_1196,N_19379,N_19598);
xor UO_1197 (O_1197,N_19357,N_19478);
and UO_1198 (O_1198,N_19745,N_19460);
nor UO_1199 (O_1199,N_19349,N_19441);
nand UO_1200 (O_1200,N_19874,N_19973);
nand UO_1201 (O_1201,N_19940,N_19253);
xnor UO_1202 (O_1202,N_19792,N_19682);
xnor UO_1203 (O_1203,N_19682,N_19876);
nor UO_1204 (O_1204,N_19593,N_19347);
or UO_1205 (O_1205,N_19528,N_19826);
or UO_1206 (O_1206,N_19964,N_19365);
nor UO_1207 (O_1207,N_19811,N_19575);
nand UO_1208 (O_1208,N_19252,N_19504);
and UO_1209 (O_1209,N_19825,N_19713);
or UO_1210 (O_1210,N_19751,N_19723);
or UO_1211 (O_1211,N_19428,N_19975);
and UO_1212 (O_1212,N_19367,N_19445);
and UO_1213 (O_1213,N_19549,N_19559);
and UO_1214 (O_1214,N_19687,N_19592);
xor UO_1215 (O_1215,N_19933,N_19494);
or UO_1216 (O_1216,N_19978,N_19493);
nand UO_1217 (O_1217,N_19972,N_19407);
nor UO_1218 (O_1218,N_19618,N_19998);
nand UO_1219 (O_1219,N_19730,N_19526);
nor UO_1220 (O_1220,N_19730,N_19721);
and UO_1221 (O_1221,N_19746,N_19691);
and UO_1222 (O_1222,N_19759,N_19600);
or UO_1223 (O_1223,N_19718,N_19754);
nor UO_1224 (O_1224,N_19810,N_19687);
nand UO_1225 (O_1225,N_19885,N_19792);
nand UO_1226 (O_1226,N_19758,N_19484);
and UO_1227 (O_1227,N_19765,N_19422);
and UO_1228 (O_1228,N_19788,N_19518);
nand UO_1229 (O_1229,N_19353,N_19893);
and UO_1230 (O_1230,N_19875,N_19334);
or UO_1231 (O_1231,N_19432,N_19409);
xnor UO_1232 (O_1232,N_19852,N_19894);
nor UO_1233 (O_1233,N_19405,N_19750);
and UO_1234 (O_1234,N_19233,N_19465);
xor UO_1235 (O_1235,N_19473,N_19386);
nand UO_1236 (O_1236,N_19523,N_19338);
and UO_1237 (O_1237,N_19842,N_19564);
nand UO_1238 (O_1238,N_19701,N_19295);
and UO_1239 (O_1239,N_19705,N_19945);
nor UO_1240 (O_1240,N_19659,N_19325);
nor UO_1241 (O_1241,N_19531,N_19388);
nor UO_1242 (O_1242,N_19816,N_19452);
and UO_1243 (O_1243,N_19432,N_19488);
nand UO_1244 (O_1244,N_19629,N_19869);
nand UO_1245 (O_1245,N_19512,N_19254);
nand UO_1246 (O_1246,N_19405,N_19554);
xnor UO_1247 (O_1247,N_19331,N_19630);
nand UO_1248 (O_1248,N_19862,N_19398);
and UO_1249 (O_1249,N_19857,N_19269);
or UO_1250 (O_1250,N_19976,N_19721);
nand UO_1251 (O_1251,N_19344,N_19580);
xnor UO_1252 (O_1252,N_19883,N_19370);
xor UO_1253 (O_1253,N_19658,N_19482);
and UO_1254 (O_1254,N_19486,N_19977);
and UO_1255 (O_1255,N_19562,N_19248);
and UO_1256 (O_1256,N_19871,N_19606);
xnor UO_1257 (O_1257,N_19542,N_19424);
or UO_1258 (O_1258,N_19744,N_19435);
and UO_1259 (O_1259,N_19913,N_19782);
nand UO_1260 (O_1260,N_19475,N_19368);
nor UO_1261 (O_1261,N_19348,N_19590);
nor UO_1262 (O_1262,N_19918,N_19820);
or UO_1263 (O_1263,N_19654,N_19779);
nand UO_1264 (O_1264,N_19770,N_19457);
nand UO_1265 (O_1265,N_19342,N_19497);
xor UO_1266 (O_1266,N_19386,N_19939);
or UO_1267 (O_1267,N_19265,N_19560);
nand UO_1268 (O_1268,N_19541,N_19683);
nand UO_1269 (O_1269,N_19820,N_19500);
nand UO_1270 (O_1270,N_19815,N_19843);
nand UO_1271 (O_1271,N_19776,N_19817);
nand UO_1272 (O_1272,N_19771,N_19685);
nand UO_1273 (O_1273,N_19530,N_19286);
or UO_1274 (O_1274,N_19421,N_19713);
nor UO_1275 (O_1275,N_19622,N_19353);
xor UO_1276 (O_1276,N_19233,N_19455);
and UO_1277 (O_1277,N_19362,N_19460);
xor UO_1278 (O_1278,N_19806,N_19250);
xor UO_1279 (O_1279,N_19920,N_19599);
nand UO_1280 (O_1280,N_19777,N_19551);
nor UO_1281 (O_1281,N_19738,N_19801);
nand UO_1282 (O_1282,N_19573,N_19333);
and UO_1283 (O_1283,N_19269,N_19805);
xnor UO_1284 (O_1284,N_19278,N_19886);
nand UO_1285 (O_1285,N_19927,N_19638);
and UO_1286 (O_1286,N_19880,N_19847);
nor UO_1287 (O_1287,N_19214,N_19913);
or UO_1288 (O_1288,N_19547,N_19961);
nor UO_1289 (O_1289,N_19749,N_19768);
or UO_1290 (O_1290,N_19658,N_19430);
xnor UO_1291 (O_1291,N_19414,N_19206);
and UO_1292 (O_1292,N_19338,N_19633);
nand UO_1293 (O_1293,N_19556,N_19537);
nor UO_1294 (O_1294,N_19933,N_19391);
or UO_1295 (O_1295,N_19789,N_19593);
or UO_1296 (O_1296,N_19870,N_19775);
nand UO_1297 (O_1297,N_19451,N_19613);
or UO_1298 (O_1298,N_19891,N_19844);
or UO_1299 (O_1299,N_19838,N_19353);
or UO_1300 (O_1300,N_19456,N_19552);
and UO_1301 (O_1301,N_19748,N_19666);
xnor UO_1302 (O_1302,N_19211,N_19374);
or UO_1303 (O_1303,N_19214,N_19271);
xnor UO_1304 (O_1304,N_19244,N_19936);
nor UO_1305 (O_1305,N_19480,N_19518);
nand UO_1306 (O_1306,N_19659,N_19717);
and UO_1307 (O_1307,N_19535,N_19310);
nand UO_1308 (O_1308,N_19636,N_19895);
xor UO_1309 (O_1309,N_19390,N_19505);
nor UO_1310 (O_1310,N_19804,N_19767);
nand UO_1311 (O_1311,N_19560,N_19963);
nor UO_1312 (O_1312,N_19823,N_19202);
or UO_1313 (O_1313,N_19303,N_19269);
or UO_1314 (O_1314,N_19495,N_19747);
and UO_1315 (O_1315,N_19880,N_19614);
or UO_1316 (O_1316,N_19752,N_19436);
or UO_1317 (O_1317,N_19266,N_19596);
nor UO_1318 (O_1318,N_19778,N_19410);
nor UO_1319 (O_1319,N_19421,N_19845);
nand UO_1320 (O_1320,N_19922,N_19537);
xnor UO_1321 (O_1321,N_19987,N_19843);
xor UO_1322 (O_1322,N_19288,N_19343);
and UO_1323 (O_1323,N_19621,N_19526);
nor UO_1324 (O_1324,N_19302,N_19872);
nor UO_1325 (O_1325,N_19304,N_19915);
nand UO_1326 (O_1326,N_19229,N_19543);
xnor UO_1327 (O_1327,N_19709,N_19396);
and UO_1328 (O_1328,N_19847,N_19684);
xor UO_1329 (O_1329,N_19554,N_19843);
xor UO_1330 (O_1330,N_19420,N_19824);
and UO_1331 (O_1331,N_19444,N_19878);
nor UO_1332 (O_1332,N_19629,N_19391);
or UO_1333 (O_1333,N_19675,N_19851);
nor UO_1334 (O_1334,N_19957,N_19688);
nor UO_1335 (O_1335,N_19402,N_19782);
or UO_1336 (O_1336,N_19705,N_19336);
nand UO_1337 (O_1337,N_19622,N_19616);
nor UO_1338 (O_1338,N_19341,N_19962);
and UO_1339 (O_1339,N_19611,N_19469);
nand UO_1340 (O_1340,N_19500,N_19966);
or UO_1341 (O_1341,N_19784,N_19621);
nand UO_1342 (O_1342,N_19641,N_19209);
or UO_1343 (O_1343,N_19752,N_19602);
and UO_1344 (O_1344,N_19224,N_19592);
or UO_1345 (O_1345,N_19990,N_19619);
or UO_1346 (O_1346,N_19751,N_19943);
xnor UO_1347 (O_1347,N_19918,N_19868);
nor UO_1348 (O_1348,N_19883,N_19230);
nor UO_1349 (O_1349,N_19853,N_19388);
xor UO_1350 (O_1350,N_19250,N_19890);
xor UO_1351 (O_1351,N_19394,N_19832);
nor UO_1352 (O_1352,N_19461,N_19385);
or UO_1353 (O_1353,N_19280,N_19568);
nand UO_1354 (O_1354,N_19604,N_19203);
or UO_1355 (O_1355,N_19522,N_19668);
and UO_1356 (O_1356,N_19214,N_19386);
or UO_1357 (O_1357,N_19462,N_19834);
nand UO_1358 (O_1358,N_19650,N_19286);
nand UO_1359 (O_1359,N_19436,N_19896);
nor UO_1360 (O_1360,N_19220,N_19386);
nand UO_1361 (O_1361,N_19376,N_19936);
nand UO_1362 (O_1362,N_19358,N_19976);
and UO_1363 (O_1363,N_19766,N_19299);
xor UO_1364 (O_1364,N_19885,N_19306);
xnor UO_1365 (O_1365,N_19330,N_19860);
or UO_1366 (O_1366,N_19651,N_19802);
xor UO_1367 (O_1367,N_19869,N_19993);
xor UO_1368 (O_1368,N_19762,N_19771);
and UO_1369 (O_1369,N_19907,N_19267);
xor UO_1370 (O_1370,N_19491,N_19330);
xnor UO_1371 (O_1371,N_19537,N_19440);
and UO_1372 (O_1372,N_19207,N_19685);
xnor UO_1373 (O_1373,N_19745,N_19662);
nand UO_1374 (O_1374,N_19976,N_19636);
and UO_1375 (O_1375,N_19247,N_19465);
nand UO_1376 (O_1376,N_19223,N_19903);
and UO_1377 (O_1377,N_19760,N_19304);
or UO_1378 (O_1378,N_19251,N_19936);
xnor UO_1379 (O_1379,N_19814,N_19825);
and UO_1380 (O_1380,N_19635,N_19916);
nand UO_1381 (O_1381,N_19239,N_19333);
or UO_1382 (O_1382,N_19799,N_19416);
and UO_1383 (O_1383,N_19433,N_19800);
or UO_1384 (O_1384,N_19405,N_19518);
nand UO_1385 (O_1385,N_19830,N_19883);
xnor UO_1386 (O_1386,N_19473,N_19579);
nand UO_1387 (O_1387,N_19865,N_19520);
xor UO_1388 (O_1388,N_19402,N_19252);
and UO_1389 (O_1389,N_19302,N_19261);
and UO_1390 (O_1390,N_19869,N_19935);
nand UO_1391 (O_1391,N_19761,N_19882);
and UO_1392 (O_1392,N_19215,N_19936);
nand UO_1393 (O_1393,N_19363,N_19673);
nor UO_1394 (O_1394,N_19314,N_19961);
xor UO_1395 (O_1395,N_19710,N_19457);
or UO_1396 (O_1396,N_19942,N_19206);
xnor UO_1397 (O_1397,N_19275,N_19939);
xnor UO_1398 (O_1398,N_19306,N_19593);
or UO_1399 (O_1399,N_19526,N_19345);
nor UO_1400 (O_1400,N_19567,N_19472);
xor UO_1401 (O_1401,N_19433,N_19441);
nand UO_1402 (O_1402,N_19283,N_19797);
xnor UO_1403 (O_1403,N_19360,N_19279);
nor UO_1404 (O_1404,N_19456,N_19900);
nand UO_1405 (O_1405,N_19349,N_19243);
or UO_1406 (O_1406,N_19588,N_19600);
nor UO_1407 (O_1407,N_19300,N_19792);
xnor UO_1408 (O_1408,N_19427,N_19956);
and UO_1409 (O_1409,N_19300,N_19416);
or UO_1410 (O_1410,N_19746,N_19626);
nor UO_1411 (O_1411,N_19918,N_19997);
nand UO_1412 (O_1412,N_19415,N_19299);
or UO_1413 (O_1413,N_19262,N_19329);
nand UO_1414 (O_1414,N_19968,N_19428);
nand UO_1415 (O_1415,N_19704,N_19558);
xnor UO_1416 (O_1416,N_19392,N_19458);
or UO_1417 (O_1417,N_19221,N_19580);
nor UO_1418 (O_1418,N_19388,N_19965);
nand UO_1419 (O_1419,N_19286,N_19245);
nand UO_1420 (O_1420,N_19990,N_19525);
nand UO_1421 (O_1421,N_19324,N_19727);
or UO_1422 (O_1422,N_19571,N_19803);
nand UO_1423 (O_1423,N_19683,N_19302);
nand UO_1424 (O_1424,N_19592,N_19275);
or UO_1425 (O_1425,N_19783,N_19553);
or UO_1426 (O_1426,N_19695,N_19933);
nand UO_1427 (O_1427,N_19658,N_19220);
nand UO_1428 (O_1428,N_19405,N_19627);
or UO_1429 (O_1429,N_19866,N_19288);
nand UO_1430 (O_1430,N_19497,N_19853);
and UO_1431 (O_1431,N_19321,N_19284);
and UO_1432 (O_1432,N_19598,N_19406);
xor UO_1433 (O_1433,N_19494,N_19380);
and UO_1434 (O_1434,N_19793,N_19782);
and UO_1435 (O_1435,N_19680,N_19634);
nor UO_1436 (O_1436,N_19866,N_19575);
nand UO_1437 (O_1437,N_19922,N_19726);
or UO_1438 (O_1438,N_19463,N_19657);
xor UO_1439 (O_1439,N_19553,N_19351);
xor UO_1440 (O_1440,N_19998,N_19757);
xor UO_1441 (O_1441,N_19417,N_19433);
xnor UO_1442 (O_1442,N_19877,N_19536);
and UO_1443 (O_1443,N_19432,N_19878);
or UO_1444 (O_1444,N_19624,N_19206);
nor UO_1445 (O_1445,N_19346,N_19839);
nor UO_1446 (O_1446,N_19328,N_19696);
nand UO_1447 (O_1447,N_19473,N_19400);
or UO_1448 (O_1448,N_19547,N_19592);
and UO_1449 (O_1449,N_19732,N_19508);
nand UO_1450 (O_1450,N_19430,N_19825);
nor UO_1451 (O_1451,N_19948,N_19612);
nand UO_1452 (O_1452,N_19986,N_19622);
or UO_1453 (O_1453,N_19547,N_19905);
or UO_1454 (O_1454,N_19317,N_19723);
xor UO_1455 (O_1455,N_19650,N_19261);
xnor UO_1456 (O_1456,N_19665,N_19673);
nor UO_1457 (O_1457,N_19504,N_19524);
nor UO_1458 (O_1458,N_19283,N_19433);
or UO_1459 (O_1459,N_19662,N_19728);
nand UO_1460 (O_1460,N_19506,N_19360);
xor UO_1461 (O_1461,N_19755,N_19760);
and UO_1462 (O_1462,N_19842,N_19305);
xor UO_1463 (O_1463,N_19207,N_19788);
or UO_1464 (O_1464,N_19450,N_19774);
or UO_1465 (O_1465,N_19651,N_19513);
nor UO_1466 (O_1466,N_19447,N_19581);
nand UO_1467 (O_1467,N_19502,N_19983);
nor UO_1468 (O_1468,N_19742,N_19236);
nand UO_1469 (O_1469,N_19494,N_19305);
and UO_1470 (O_1470,N_19562,N_19355);
nand UO_1471 (O_1471,N_19711,N_19467);
or UO_1472 (O_1472,N_19983,N_19333);
nand UO_1473 (O_1473,N_19440,N_19700);
nor UO_1474 (O_1474,N_19549,N_19793);
or UO_1475 (O_1475,N_19885,N_19772);
and UO_1476 (O_1476,N_19592,N_19285);
and UO_1477 (O_1477,N_19512,N_19382);
or UO_1478 (O_1478,N_19460,N_19878);
nand UO_1479 (O_1479,N_19993,N_19729);
and UO_1480 (O_1480,N_19224,N_19423);
nand UO_1481 (O_1481,N_19306,N_19731);
nor UO_1482 (O_1482,N_19669,N_19225);
xor UO_1483 (O_1483,N_19531,N_19443);
nand UO_1484 (O_1484,N_19967,N_19550);
nand UO_1485 (O_1485,N_19555,N_19457);
or UO_1486 (O_1486,N_19352,N_19961);
xor UO_1487 (O_1487,N_19342,N_19504);
nor UO_1488 (O_1488,N_19277,N_19284);
nand UO_1489 (O_1489,N_19229,N_19601);
or UO_1490 (O_1490,N_19720,N_19387);
nor UO_1491 (O_1491,N_19855,N_19522);
nor UO_1492 (O_1492,N_19203,N_19282);
xor UO_1493 (O_1493,N_19445,N_19557);
nand UO_1494 (O_1494,N_19460,N_19670);
nand UO_1495 (O_1495,N_19811,N_19808);
xnor UO_1496 (O_1496,N_19729,N_19228);
xor UO_1497 (O_1497,N_19405,N_19716);
nand UO_1498 (O_1498,N_19862,N_19596);
nor UO_1499 (O_1499,N_19674,N_19972);
and UO_1500 (O_1500,N_19642,N_19906);
nor UO_1501 (O_1501,N_19253,N_19774);
nand UO_1502 (O_1502,N_19288,N_19926);
and UO_1503 (O_1503,N_19636,N_19484);
nand UO_1504 (O_1504,N_19468,N_19709);
nor UO_1505 (O_1505,N_19866,N_19669);
or UO_1506 (O_1506,N_19809,N_19233);
nor UO_1507 (O_1507,N_19276,N_19830);
and UO_1508 (O_1508,N_19437,N_19844);
nand UO_1509 (O_1509,N_19291,N_19820);
and UO_1510 (O_1510,N_19906,N_19470);
and UO_1511 (O_1511,N_19952,N_19310);
or UO_1512 (O_1512,N_19680,N_19420);
nand UO_1513 (O_1513,N_19269,N_19293);
or UO_1514 (O_1514,N_19213,N_19239);
and UO_1515 (O_1515,N_19388,N_19553);
nor UO_1516 (O_1516,N_19704,N_19981);
nand UO_1517 (O_1517,N_19883,N_19887);
xor UO_1518 (O_1518,N_19769,N_19888);
and UO_1519 (O_1519,N_19447,N_19599);
and UO_1520 (O_1520,N_19985,N_19352);
and UO_1521 (O_1521,N_19747,N_19913);
and UO_1522 (O_1522,N_19444,N_19556);
nor UO_1523 (O_1523,N_19669,N_19747);
xor UO_1524 (O_1524,N_19925,N_19790);
and UO_1525 (O_1525,N_19254,N_19652);
and UO_1526 (O_1526,N_19624,N_19469);
nand UO_1527 (O_1527,N_19869,N_19908);
or UO_1528 (O_1528,N_19914,N_19840);
nor UO_1529 (O_1529,N_19617,N_19470);
nand UO_1530 (O_1530,N_19249,N_19565);
xor UO_1531 (O_1531,N_19705,N_19524);
and UO_1532 (O_1532,N_19318,N_19597);
and UO_1533 (O_1533,N_19250,N_19221);
nor UO_1534 (O_1534,N_19535,N_19946);
nand UO_1535 (O_1535,N_19244,N_19938);
and UO_1536 (O_1536,N_19957,N_19488);
or UO_1537 (O_1537,N_19548,N_19504);
nand UO_1538 (O_1538,N_19362,N_19527);
nor UO_1539 (O_1539,N_19683,N_19695);
or UO_1540 (O_1540,N_19778,N_19381);
nand UO_1541 (O_1541,N_19534,N_19238);
nand UO_1542 (O_1542,N_19250,N_19809);
nor UO_1543 (O_1543,N_19257,N_19411);
xnor UO_1544 (O_1544,N_19988,N_19263);
nand UO_1545 (O_1545,N_19475,N_19746);
and UO_1546 (O_1546,N_19854,N_19537);
nor UO_1547 (O_1547,N_19614,N_19886);
or UO_1548 (O_1548,N_19430,N_19422);
or UO_1549 (O_1549,N_19498,N_19222);
nor UO_1550 (O_1550,N_19379,N_19633);
and UO_1551 (O_1551,N_19683,N_19454);
and UO_1552 (O_1552,N_19688,N_19894);
xnor UO_1553 (O_1553,N_19347,N_19988);
or UO_1554 (O_1554,N_19799,N_19376);
xor UO_1555 (O_1555,N_19995,N_19479);
nor UO_1556 (O_1556,N_19722,N_19901);
and UO_1557 (O_1557,N_19391,N_19679);
xnor UO_1558 (O_1558,N_19484,N_19250);
and UO_1559 (O_1559,N_19461,N_19880);
and UO_1560 (O_1560,N_19630,N_19468);
nor UO_1561 (O_1561,N_19396,N_19969);
nor UO_1562 (O_1562,N_19561,N_19949);
nand UO_1563 (O_1563,N_19475,N_19973);
xnor UO_1564 (O_1564,N_19852,N_19731);
or UO_1565 (O_1565,N_19600,N_19595);
and UO_1566 (O_1566,N_19390,N_19550);
and UO_1567 (O_1567,N_19636,N_19842);
xnor UO_1568 (O_1568,N_19474,N_19852);
nor UO_1569 (O_1569,N_19218,N_19973);
xor UO_1570 (O_1570,N_19266,N_19918);
and UO_1571 (O_1571,N_19996,N_19414);
nor UO_1572 (O_1572,N_19706,N_19222);
nor UO_1573 (O_1573,N_19926,N_19313);
and UO_1574 (O_1574,N_19258,N_19808);
or UO_1575 (O_1575,N_19559,N_19733);
and UO_1576 (O_1576,N_19303,N_19812);
nor UO_1577 (O_1577,N_19770,N_19737);
or UO_1578 (O_1578,N_19375,N_19427);
and UO_1579 (O_1579,N_19243,N_19585);
nor UO_1580 (O_1580,N_19641,N_19335);
nand UO_1581 (O_1581,N_19577,N_19967);
nor UO_1582 (O_1582,N_19773,N_19884);
and UO_1583 (O_1583,N_19480,N_19547);
and UO_1584 (O_1584,N_19849,N_19578);
and UO_1585 (O_1585,N_19868,N_19723);
nor UO_1586 (O_1586,N_19320,N_19779);
and UO_1587 (O_1587,N_19857,N_19851);
or UO_1588 (O_1588,N_19757,N_19505);
xor UO_1589 (O_1589,N_19605,N_19648);
and UO_1590 (O_1590,N_19775,N_19476);
nand UO_1591 (O_1591,N_19967,N_19934);
nor UO_1592 (O_1592,N_19791,N_19335);
and UO_1593 (O_1593,N_19246,N_19254);
and UO_1594 (O_1594,N_19310,N_19320);
nand UO_1595 (O_1595,N_19545,N_19550);
nor UO_1596 (O_1596,N_19977,N_19641);
or UO_1597 (O_1597,N_19436,N_19944);
xnor UO_1598 (O_1598,N_19476,N_19862);
xor UO_1599 (O_1599,N_19454,N_19233);
nor UO_1600 (O_1600,N_19579,N_19843);
xor UO_1601 (O_1601,N_19824,N_19391);
xor UO_1602 (O_1602,N_19715,N_19339);
nor UO_1603 (O_1603,N_19483,N_19405);
nor UO_1604 (O_1604,N_19221,N_19265);
nor UO_1605 (O_1605,N_19225,N_19341);
nand UO_1606 (O_1606,N_19428,N_19709);
nand UO_1607 (O_1607,N_19227,N_19213);
nand UO_1608 (O_1608,N_19306,N_19869);
and UO_1609 (O_1609,N_19792,N_19583);
or UO_1610 (O_1610,N_19938,N_19313);
and UO_1611 (O_1611,N_19923,N_19919);
nand UO_1612 (O_1612,N_19582,N_19625);
or UO_1613 (O_1613,N_19892,N_19235);
nand UO_1614 (O_1614,N_19336,N_19953);
or UO_1615 (O_1615,N_19359,N_19972);
xor UO_1616 (O_1616,N_19820,N_19636);
xnor UO_1617 (O_1617,N_19666,N_19564);
and UO_1618 (O_1618,N_19382,N_19686);
nand UO_1619 (O_1619,N_19408,N_19456);
nand UO_1620 (O_1620,N_19595,N_19758);
and UO_1621 (O_1621,N_19976,N_19318);
nand UO_1622 (O_1622,N_19494,N_19953);
or UO_1623 (O_1623,N_19886,N_19866);
and UO_1624 (O_1624,N_19253,N_19716);
or UO_1625 (O_1625,N_19661,N_19385);
nand UO_1626 (O_1626,N_19682,N_19564);
nand UO_1627 (O_1627,N_19546,N_19650);
nand UO_1628 (O_1628,N_19985,N_19541);
and UO_1629 (O_1629,N_19644,N_19649);
xnor UO_1630 (O_1630,N_19435,N_19458);
nor UO_1631 (O_1631,N_19932,N_19361);
xor UO_1632 (O_1632,N_19544,N_19437);
xnor UO_1633 (O_1633,N_19554,N_19566);
xnor UO_1634 (O_1634,N_19349,N_19648);
and UO_1635 (O_1635,N_19242,N_19467);
nand UO_1636 (O_1636,N_19841,N_19919);
nor UO_1637 (O_1637,N_19698,N_19462);
nand UO_1638 (O_1638,N_19449,N_19631);
nand UO_1639 (O_1639,N_19824,N_19943);
nor UO_1640 (O_1640,N_19969,N_19367);
and UO_1641 (O_1641,N_19770,N_19694);
nand UO_1642 (O_1642,N_19539,N_19662);
xor UO_1643 (O_1643,N_19656,N_19970);
xor UO_1644 (O_1644,N_19500,N_19719);
and UO_1645 (O_1645,N_19553,N_19902);
or UO_1646 (O_1646,N_19602,N_19448);
nor UO_1647 (O_1647,N_19428,N_19275);
nand UO_1648 (O_1648,N_19828,N_19299);
and UO_1649 (O_1649,N_19439,N_19390);
nand UO_1650 (O_1650,N_19264,N_19710);
nor UO_1651 (O_1651,N_19584,N_19988);
nand UO_1652 (O_1652,N_19570,N_19632);
nand UO_1653 (O_1653,N_19691,N_19788);
nor UO_1654 (O_1654,N_19612,N_19260);
xor UO_1655 (O_1655,N_19970,N_19713);
nand UO_1656 (O_1656,N_19422,N_19996);
xor UO_1657 (O_1657,N_19923,N_19952);
nor UO_1658 (O_1658,N_19966,N_19937);
nor UO_1659 (O_1659,N_19860,N_19590);
nor UO_1660 (O_1660,N_19924,N_19750);
nor UO_1661 (O_1661,N_19404,N_19638);
nor UO_1662 (O_1662,N_19338,N_19466);
nor UO_1663 (O_1663,N_19712,N_19327);
or UO_1664 (O_1664,N_19866,N_19298);
or UO_1665 (O_1665,N_19473,N_19952);
nor UO_1666 (O_1666,N_19694,N_19308);
xor UO_1667 (O_1667,N_19929,N_19436);
xnor UO_1668 (O_1668,N_19996,N_19752);
and UO_1669 (O_1669,N_19700,N_19938);
and UO_1670 (O_1670,N_19993,N_19369);
nand UO_1671 (O_1671,N_19268,N_19401);
or UO_1672 (O_1672,N_19370,N_19877);
and UO_1673 (O_1673,N_19888,N_19828);
xor UO_1674 (O_1674,N_19894,N_19895);
xnor UO_1675 (O_1675,N_19630,N_19904);
nor UO_1676 (O_1676,N_19900,N_19219);
xor UO_1677 (O_1677,N_19359,N_19961);
or UO_1678 (O_1678,N_19799,N_19819);
nand UO_1679 (O_1679,N_19575,N_19690);
nand UO_1680 (O_1680,N_19441,N_19518);
and UO_1681 (O_1681,N_19250,N_19752);
or UO_1682 (O_1682,N_19762,N_19308);
nor UO_1683 (O_1683,N_19464,N_19779);
and UO_1684 (O_1684,N_19629,N_19444);
nand UO_1685 (O_1685,N_19429,N_19550);
xnor UO_1686 (O_1686,N_19339,N_19744);
nand UO_1687 (O_1687,N_19742,N_19614);
nand UO_1688 (O_1688,N_19749,N_19758);
or UO_1689 (O_1689,N_19414,N_19404);
nor UO_1690 (O_1690,N_19893,N_19772);
or UO_1691 (O_1691,N_19243,N_19575);
nor UO_1692 (O_1692,N_19781,N_19512);
xnor UO_1693 (O_1693,N_19402,N_19489);
nand UO_1694 (O_1694,N_19368,N_19484);
or UO_1695 (O_1695,N_19260,N_19417);
or UO_1696 (O_1696,N_19600,N_19798);
nor UO_1697 (O_1697,N_19395,N_19845);
and UO_1698 (O_1698,N_19767,N_19629);
nand UO_1699 (O_1699,N_19511,N_19839);
nand UO_1700 (O_1700,N_19545,N_19403);
nand UO_1701 (O_1701,N_19935,N_19811);
or UO_1702 (O_1702,N_19423,N_19847);
or UO_1703 (O_1703,N_19992,N_19396);
xor UO_1704 (O_1704,N_19367,N_19294);
xnor UO_1705 (O_1705,N_19283,N_19375);
nor UO_1706 (O_1706,N_19424,N_19862);
nor UO_1707 (O_1707,N_19219,N_19222);
or UO_1708 (O_1708,N_19825,N_19868);
xor UO_1709 (O_1709,N_19648,N_19616);
nand UO_1710 (O_1710,N_19807,N_19411);
and UO_1711 (O_1711,N_19510,N_19476);
nand UO_1712 (O_1712,N_19705,N_19915);
or UO_1713 (O_1713,N_19566,N_19751);
nand UO_1714 (O_1714,N_19237,N_19205);
nand UO_1715 (O_1715,N_19266,N_19273);
or UO_1716 (O_1716,N_19904,N_19346);
nor UO_1717 (O_1717,N_19408,N_19452);
xor UO_1718 (O_1718,N_19908,N_19918);
and UO_1719 (O_1719,N_19664,N_19500);
xnor UO_1720 (O_1720,N_19593,N_19389);
xor UO_1721 (O_1721,N_19448,N_19220);
nor UO_1722 (O_1722,N_19269,N_19262);
nor UO_1723 (O_1723,N_19301,N_19723);
nand UO_1724 (O_1724,N_19724,N_19867);
nand UO_1725 (O_1725,N_19465,N_19702);
and UO_1726 (O_1726,N_19572,N_19400);
and UO_1727 (O_1727,N_19581,N_19766);
nand UO_1728 (O_1728,N_19241,N_19465);
nand UO_1729 (O_1729,N_19424,N_19850);
or UO_1730 (O_1730,N_19568,N_19239);
xnor UO_1731 (O_1731,N_19975,N_19249);
nor UO_1732 (O_1732,N_19499,N_19480);
nand UO_1733 (O_1733,N_19416,N_19804);
or UO_1734 (O_1734,N_19324,N_19375);
nor UO_1735 (O_1735,N_19837,N_19802);
nand UO_1736 (O_1736,N_19335,N_19668);
or UO_1737 (O_1737,N_19636,N_19783);
nand UO_1738 (O_1738,N_19872,N_19439);
nor UO_1739 (O_1739,N_19209,N_19905);
nor UO_1740 (O_1740,N_19473,N_19709);
nand UO_1741 (O_1741,N_19592,N_19847);
nand UO_1742 (O_1742,N_19284,N_19389);
or UO_1743 (O_1743,N_19202,N_19875);
nand UO_1744 (O_1744,N_19906,N_19996);
xnor UO_1745 (O_1745,N_19452,N_19887);
nor UO_1746 (O_1746,N_19535,N_19324);
or UO_1747 (O_1747,N_19506,N_19343);
nand UO_1748 (O_1748,N_19975,N_19658);
nand UO_1749 (O_1749,N_19372,N_19411);
nand UO_1750 (O_1750,N_19264,N_19622);
xor UO_1751 (O_1751,N_19674,N_19775);
or UO_1752 (O_1752,N_19394,N_19943);
nor UO_1753 (O_1753,N_19958,N_19504);
nand UO_1754 (O_1754,N_19452,N_19776);
or UO_1755 (O_1755,N_19548,N_19589);
nand UO_1756 (O_1756,N_19287,N_19856);
or UO_1757 (O_1757,N_19200,N_19928);
and UO_1758 (O_1758,N_19802,N_19359);
xor UO_1759 (O_1759,N_19329,N_19453);
nand UO_1760 (O_1760,N_19913,N_19207);
xnor UO_1761 (O_1761,N_19543,N_19778);
nor UO_1762 (O_1762,N_19849,N_19877);
xnor UO_1763 (O_1763,N_19399,N_19212);
nand UO_1764 (O_1764,N_19688,N_19935);
or UO_1765 (O_1765,N_19783,N_19602);
nor UO_1766 (O_1766,N_19987,N_19523);
xnor UO_1767 (O_1767,N_19347,N_19664);
nand UO_1768 (O_1768,N_19575,N_19847);
and UO_1769 (O_1769,N_19844,N_19544);
nand UO_1770 (O_1770,N_19555,N_19787);
nor UO_1771 (O_1771,N_19862,N_19479);
or UO_1772 (O_1772,N_19949,N_19730);
xor UO_1773 (O_1773,N_19723,N_19302);
xnor UO_1774 (O_1774,N_19790,N_19289);
nand UO_1775 (O_1775,N_19336,N_19234);
and UO_1776 (O_1776,N_19437,N_19476);
nor UO_1777 (O_1777,N_19213,N_19205);
or UO_1778 (O_1778,N_19298,N_19415);
nor UO_1779 (O_1779,N_19435,N_19889);
xor UO_1780 (O_1780,N_19581,N_19648);
xnor UO_1781 (O_1781,N_19299,N_19382);
nor UO_1782 (O_1782,N_19645,N_19420);
nand UO_1783 (O_1783,N_19886,N_19409);
nor UO_1784 (O_1784,N_19301,N_19904);
nor UO_1785 (O_1785,N_19969,N_19852);
and UO_1786 (O_1786,N_19905,N_19795);
nand UO_1787 (O_1787,N_19937,N_19712);
nand UO_1788 (O_1788,N_19596,N_19502);
xor UO_1789 (O_1789,N_19201,N_19976);
and UO_1790 (O_1790,N_19275,N_19688);
xnor UO_1791 (O_1791,N_19525,N_19403);
and UO_1792 (O_1792,N_19287,N_19545);
nor UO_1793 (O_1793,N_19645,N_19349);
xnor UO_1794 (O_1794,N_19891,N_19414);
xor UO_1795 (O_1795,N_19586,N_19658);
or UO_1796 (O_1796,N_19596,N_19710);
nand UO_1797 (O_1797,N_19990,N_19902);
nand UO_1798 (O_1798,N_19309,N_19799);
or UO_1799 (O_1799,N_19803,N_19869);
nand UO_1800 (O_1800,N_19705,N_19553);
xor UO_1801 (O_1801,N_19380,N_19252);
and UO_1802 (O_1802,N_19414,N_19888);
and UO_1803 (O_1803,N_19797,N_19842);
nand UO_1804 (O_1804,N_19784,N_19928);
and UO_1805 (O_1805,N_19338,N_19879);
xor UO_1806 (O_1806,N_19705,N_19359);
nor UO_1807 (O_1807,N_19270,N_19277);
and UO_1808 (O_1808,N_19957,N_19807);
nand UO_1809 (O_1809,N_19516,N_19875);
or UO_1810 (O_1810,N_19820,N_19885);
and UO_1811 (O_1811,N_19637,N_19398);
nor UO_1812 (O_1812,N_19335,N_19333);
or UO_1813 (O_1813,N_19240,N_19392);
nor UO_1814 (O_1814,N_19806,N_19230);
nand UO_1815 (O_1815,N_19306,N_19323);
and UO_1816 (O_1816,N_19332,N_19630);
nand UO_1817 (O_1817,N_19744,N_19704);
nand UO_1818 (O_1818,N_19555,N_19561);
nand UO_1819 (O_1819,N_19750,N_19411);
and UO_1820 (O_1820,N_19203,N_19603);
and UO_1821 (O_1821,N_19226,N_19337);
nand UO_1822 (O_1822,N_19897,N_19338);
nor UO_1823 (O_1823,N_19967,N_19839);
or UO_1824 (O_1824,N_19644,N_19214);
nand UO_1825 (O_1825,N_19529,N_19678);
xnor UO_1826 (O_1826,N_19353,N_19473);
or UO_1827 (O_1827,N_19803,N_19851);
nor UO_1828 (O_1828,N_19728,N_19793);
or UO_1829 (O_1829,N_19888,N_19861);
xnor UO_1830 (O_1830,N_19881,N_19393);
nand UO_1831 (O_1831,N_19820,N_19975);
xor UO_1832 (O_1832,N_19420,N_19718);
nand UO_1833 (O_1833,N_19713,N_19367);
nand UO_1834 (O_1834,N_19568,N_19387);
and UO_1835 (O_1835,N_19284,N_19493);
nand UO_1836 (O_1836,N_19547,N_19223);
nor UO_1837 (O_1837,N_19657,N_19374);
nor UO_1838 (O_1838,N_19306,N_19862);
xnor UO_1839 (O_1839,N_19811,N_19385);
xnor UO_1840 (O_1840,N_19997,N_19661);
and UO_1841 (O_1841,N_19726,N_19486);
xnor UO_1842 (O_1842,N_19626,N_19821);
xnor UO_1843 (O_1843,N_19313,N_19277);
and UO_1844 (O_1844,N_19827,N_19969);
nor UO_1845 (O_1845,N_19811,N_19254);
and UO_1846 (O_1846,N_19723,N_19260);
nand UO_1847 (O_1847,N_19868,N_19752);
nor UO_1848 (O_1848,N_19595,N_19956);
and UO_1849 (O_1849,N_19394,N_19990);
or UO_1850 (O_1850,N_19673,N_19436);
and UO_1851 (O_1851,N_19954,N_19820);
nor UO_1852 (O_1852,N_19590,N_19481);
or UO_1853 (O_1853,N_19854,N_19501);
or UO_1854 (O_1854,N_19360,N_19433);
or UO_1855 (O_1855,N_19314,N_19293);
xnor UO_1856 (O_1856,N_19670,N_19876);
nand UO_1857 (O_1857,N_19244,N_19543);
nor UO_1858 (O_1858,N_19639,N_19539);
nor UO_1859 (O_1859,N_19742,N_19824);
or UO_1860 (O_1860,N_19756,N_19380);
nand UO_1861 (O_1861,N_19614,N_19903);
xor UO_1862 (O_1862,N_19807,N_19389);
or UO_1863 (O_1863,N_19794,N_19463);
or UO_1864 (O_1864,N_19746,N_19799);
xor UO_1865 (O_1865,N_19863,N_19366);
and UO_1866 (O_1866,N_19815,N_19633);
xnor UO_1867 (O_1867,N_19772,N_19247);
or UO_1868 (O_1868,N_19236,N_19345);
xnor UO_1869 (O_1869,N_19715,N_19298);
or UO_1870 (O_1870,N_19698,N_19367);
nor UO_1871 (O_1871,N_19425,N_19982);
xnor UO_1872 (O_1872,N_19397,N_19499);
nor UO_1873 (O_1873,N_19308,N_19418);
and UO_1874 (O_1874,N_19598,N_19658);
xor UO_1875 (O_1875,N_19284,N_19448);
nand UO_1876 (O_1876,N_19859,N_19335);
nor UO_1877 (O_1877,N_19377,N_19290);
xnor UO_1878 (O_1878,N_19938,N_19753);
nor UO_1879 (O_1879,N_19997,N_19489);
xnor UO_1880 (O_1880,N_19437,N_19521);
and UO_1881 (O_1881,N_19384,N_19445);
xor UO_1882 (O_1882,N_19374,N_19274);
xor UO_1883 (O_1883,N_19947,N_19570);
nor UO_1884 (O_1884,N_19668,N_19411);
or UO_1885 (O_1885,N_19398,N_19552);
or UO_1886 (O_1886,N_19295,N_19293);
and UO_1887 (O_1887,N_19314,N_19222);
or UO_1888 (O_1888,N_19874,N_19329);
or UO_1889 (O_1889,N_19822,N_19279);
nor UO_1890 (O_1890,N_19383,N_19769);
and UO_1891 (O_1891,N_19921,N_19657);
nor UO_1892 (O_1892,N_19785,N_19853);
nand UO_1893 (O_1893,N_19443,N_19302);
and UO_1894 (O_1894,N_19740,N_19690);
and UO_1895 (O_1895,N_19516,N_19916);
xnor UO_1896 (O_1896,N_19673,N_19963);
or UO_1897 (O_1897,N_19704,N_19674);
or UO_1898 (O_1898,N_19855,N_19383);
and UO_1899 (O_1899,N_19204,N_19703);
or UO_1900 (O_1900,N_19299,N_19905);
nand UO_1901 (O_1901,N_19472,N_19725);
xor UO_1902 (O_1902,N_19885,N_19466);
or UO_1903 (O_1903,N_19736,N_19938);
nor UO_1904 (O_1904,N_19647,N_19491);
nor UO_1905 (O_1905,N_19652,N_19783);
and UO_1906 (O_1906,N_19777,N_19931);
or UO_1907 (O_1907,N_19582,N_19946);
nor UO_1908 (O_1908,N_19910,N_19389);
or UO_1909 (O_1909,N_19395,N_19804);
or UO_1910 (O_1910,N_19981,N_19613);
and UO_1911 (O_1911,N_19828,N_19834);
nand UO_1912 (O_1912,N_19582,N_19953);
and UO_1913 (O_1913,N_19721,N_19929);
nand UO_1914 (O_1914,N_19748,N_19520);
or UO_1915 (O_1915,N_19240,N_19932);
nor UO_1916 (O_1916,N_19229,N_19383);
and UO_1917 (O_1917,N_19551,N_19605);
nor UO_1918 (O_1918,N_19265,N_19893);
nor UO_1919 (O_1919,N_19524,N_19718);
nor UO_1920 (O_1920,N_19472,N_19677);
or UO_1921 (O_1921,N_19541,N_19719);
and UO_1922 (O_1922,N_19846,N_19633);
nand UO_1923 (O_1923,N_19362,N_19932);
nor UO_1924 (O_1924,N_19378,N_19458);
nor UO_1925 (O_1925,N_19834,N_19374);
nor UO_1926 (O_1926,N_19624,N_19543);
xor UO_1927 (O_1927,N_19900,N_19834);
nand UO_1928 (O_1928,N_19843,N_19378);
or UO_1929 (O_1929,N_19499,N_19515);
or UO_1930 (O_1930,N_19920,N_19537);
nor UO_1931 (O_1931,N_19438,N_19619);
xnor UO_1932 (O_1932,N_19793,N_19655);
and UO_1933 (O_1933,N_19695,N_19611);
xnor UO_1934 (O_1934,N_19832,N_19838);
or UO_1935 (O_1935,N_19253,N_19842);
nand UO_1936 (O_1936,N_19474,N_19755);
or UO_1937 (O_1937,N_19742,N_19201);
nor UO_1938 (O_1938,N_19676,N_19467);
nor UO_1939 (O_1939,N_19617,N_19596);
and UO_1940 (O_1940,N_19310,N_19646);
or UO_1941 (O_1941,N_19850,N_19429);
xor UO_1942 (O_1942,N_19341,N_19262);
nor UO_1943 (O_1943,N_19989,N_19638);
or UO_1944 (O_1944,N_19987,N_19794);
or UO_1945 (O_1945,N_19371,N_19499);
xnor UO_1946 (O_1946,N_19932,N_19969);
nor UO_1947 (O_1947,N_19220,N_19306);
nand UO_1948 (O_1948,N_19830,N_19942);
and UO_1949 (O_1949,N_19872,N_19922);
and UO_1950 (O_1950,N_19679,N_19919);
xor UO_1951 (O_1951,N_19255,N_19441);
or UO_1952 (O_1952,N_19599,N_19530);
xnor UO_1953 (O_1953,N_19625,N_19610);
or UO_1954 (O_1954,N_19592,N_19205);
nand UO_1955 (O_1955,N_19576,N_19797);
or UO_1956 (O_1956,N_19749,N_19743);
xor UO_1957 (O_1957,N_19510,N_19207);
nand UO_1958 (O_1958,N_19756,N_19249);
and UO_1959 (O_1959,N_19752,N_19482);
or UO_1960 (O_1960,N_19711,N_19850);
nand UO_1961 (O_1961,N_19616,N_19838);
nor UO_1962 (O_1962,N_19959,N_19231);
and UO_1963 (O_1963,N_19759,N_19791);
or UO_1964 (O_1964,N_19381,N_19218);
or UO_1965 (O_1965,N_19838,N_19693);
and UO_1966 (O_1966,N_19384,N_19475);
and UO_1967 (O_1967,N_19220,N_19965);
nor UO_1968 (O_1968,N_19458,N_19930);
or UO_1969 (O_1969,N_19245,N_19929);
or UO_1970 (O_1970,N_19234,N_19326);
or UO_1971 (O_1971,N_19284,N_19370);
and UO_1972 (O_1972,N_19274,N_19562);
nand UO_1973 (O_1973,N_19554,N_19414);
or UO_1974 (O_1974,N_19608,N_19947);
or UO_1975 (O_1975,N_19215,N_19209);
nor UO_1976 (O_1976,N_19778,N_19475);
xnor UO_1977 (O_1977,N_19770,N_19714);
or UO_1978 (O_1978,N_19702,N_19964);
and UO_1979 (O_1979,N_19409,N_19803);
or UO_1980 (O_1980,N_19830,N_19489);
or UO_1981 (O_1981,N_19816,N_19300);
xnor UO_1982 (O_1982,N_19293,N_19461);
or UO_1983 (O_1983,N_19408,N_19387);
and UO_1984 (O_1984,N_19597,N_19636);
and UO_1985 (O_1985,N_19915,N_19888);
or UO_1986 (O_1986,N_19863,N_19425);
and UO_1987 (O_1987,N_19270,N_19741);
or UO_1988 (O_1988,N_19559,N_19556);
xnor UO_1989 (O_1989,N_19288,N_19411);
xnor UO_1990 (O_1990,N_19408,N_19353);
xor UO_1991 (O_1991,N_19412,N_19256);
nor UO_1992 (O_1992,N_19495,N_19602);
and UO_1993 (O_1993,N_19652,N_19311);
nand UO_1994 (O_1994,N_19989,N_19564);
or UO_1995 (O_1995,N_19515,N_19479);
nand UO_1996 (O_1996,N_19274,N_19525);
xnor UO_1997 (O_1997,N_19492,N_19961);
nand UO_1998 (O_1998,N_19673,N_19254);
xnor UO_1999 (O_1999,N_19738,N_19815);
nor UO_2000 (O_2000,N_19693,N_19694);
nand UO_2001 (O_2001,N_19602,N_19333);
xnor UO_2002 (O_2002,N_19215,N_19303);
nor UO_2003 (O_2003,N_19886,N_19595);
or UO_2004 (O_2004,N_19710,N_19438);
nor UO_2005 (O_2005,N_19771,N_19830);
or UO_2006 (O_2006,N_19500,N_19545);
and UO_2007 (O_2007,N_19701,N_19667);
xor UO_2008 (O_2008,N_19273,N_19461);
nor UO_2009 (O_2009,N_19647,N_19263);
and UO_2010 (O_2010,N_19508,N_19793);
and UO_2011 (O_2011,N_19829,N_19913);
nand UO_2012 (O_2012,N_19219,N_19650);
nor UO_2013 (O_2013,N_19338,N_19668);
nand UO_2014 (O_2014,N_19247,N_19891);
and UO_2015 (O_2015,N_19933,N_19708);
nor UO_2016 (O_2016,N_19723,N_19315);
or UO_2017 (O_2017,N_19875,N_19658);
and UO_2018 (O_2018,N_19655,N_19887);
or UO_2019 (O_2019,N_19767,N_19275);
or UO_2020 (O_2020,N_19236,N_19486);
and UO_2021 (O_2021,N_19276,N_19447);
or UO_2022 (O_2022,N_19407,N_19383);
nor UO_2023 (O_2023,N_19835,N_19580);
nor UO_2024 (O_2024,N_19876,N_19384);
or UO_2025 (O_2025,N_19537,N_19220);
or UO_2026 (O_2026,N_19544,N_19929);
or UO_2027 (O_2027,N_19909,N_19752);
nor UO_2028 (O_2028,N_19452,N_19280);
nor UO_2029 (O_2029,N_19387,N_19785);
xnor UO_2030 (O_2030,N_19746,N_19310);
xnor UO_2031 (O_2031,N_19301,N_19325);
xnor UO_2032 (O_2032,N_19580,N_19347);
xnor UO_2033 (O_2033,N_19950,N_19500);
xor UO_2034 (O_2034,N_19669,N_19824);
xor UO_2035 (O_2035,N_19558,N_19950);
nand UO_2036 (O_2036,N_19536,N_19405);
and UO_2037 (O_2037,N_19879,N_19765);
nor UO_2038 (O_2038,N_19759,N_19431);
xor UO_2039 (O_2039,N_19702,N_19302);
and UO_2040 (O_2040,N_19948,N_19495);
or UO_2041 (O_2041,N_19705,N_19289);
or UO_2042 (O_2042,N_19882,N_19267);
nor UO_2043 (O_2043,N_19486,N_19237);
and UO_2044 (O_2044,N_19298,N_19939);
or UO_2045 (O_2045,N_19412,N_19852);
or UO_2046 (O_2046,N_19212,N_19536);
and UO_2047 (O_2047,N_19571,N_19541);
nand UO_2048 (O_2048,N_19231,N_19322);
or UO_2049 (O_2049,N_19850,N_19646);
xor UO_2050 (O_2050,N_19548,N_19870);
or UO_2051 (O_2051,N_19603,N_19920);
xor UO_2052 (O_2052,N_19590,N_19712);
and UO_2053 (O_2053,N_19645,N_19815);
xor UO_2054 (O_2054,N_19774,N_19775);
and UO_2055 (O_2055,N_19966,N_19863);
nand UO_2056 (O_2056,N_19424,N_19549);
xor UO_2057 (O_2057,N_19293,N_19769);
and UO_2058 (O_2058,N_19327,N_19856);
nand UO_2059 (O_2059,N_19405,N_19225);
xor UO_2060 (O_2060,N_19864,N_19764);
nor UO_2061 (O_2061,N_19675,N_19948);
or UO_2062 (O_2062,N_19379,N_19553);
nand UO_2063 (O_2063,N_19740,N_19469);
nand UO_2064 (O_2064,N_19859,N_19662);
nor UO_2065 (O_2065,N_19933,N_19775);
or UO_2066 (O_2066,N_19338,N_19823);
or UO_2067 (O_2067,N_19898,N_19769);
xor UO_2068 (O_2068,N_19603,N_19311);
nand UO_2069 (O_2069,N_19844,N_19750);
or UO_2070 (O_2070,N_19552,N_19827);
or UO_2071 (O_2071,N_19874,N_19750);
nand UO_2072 (O_2072,N_19569,N_19764);
or UO_2073 (O_2073,N_19833,N_19963);
or UO_2074 (O_2074,N_19222,N_19754);
or UO_2075 (O_2075,N_19867,N_19756);
and UO_2076 (O_2076,N_19436,N_19927);
nor UO_2077 (O_2077,N_19753,N_19408);
xor UO_2078 (O_2078,N_19366,N_19201);
nor UO_2079 (O_2079,N_19235,N_19921);
or UO_2080 (O_2080,N_19837,N_19343);
xnor UO_2081 (O_2081,N_19604,N_19682);
and UO_2082 (O_2082,N_19749,N_19489);
nand UO_2083 (O_2083,N_19642,N_19976);
or UO_2084 (O_2084,N_19481,N_19589);
nor UO_2085 (O_2085,N_19936,N_19688);
nand UO_2086 (O_2086,N_19358,N_19634);
and UO_2087 (O_2087,N_19665,N_19676);
and UO_2088 (O_2088,N_19215,N_19212);
nand UO_2089 (O_2089,N_19712,N_19611);
or UO_2090 (O_2090,N_19640,N_19413);
nor UO_2091 (O_2091,N_19781,N_19247);
or UO_2092 (O_2092,N_19257,N_19394);
or UO_2093 (O_2093,N_19769,N_19664);
or UO_2094 (O_2094,N_19413,N_19749);
nor UO_2095 (O_2095,N_19686,N_19854);
nand UO_2096 (O_2096,N_19964,N_19809);
nand UO_2097 (O_2097,N_19367,N_19369);
or UO_2098 (O_2098,N_19482,N_19222);
xnor UO_2099 (O_2099,N_19694,N_19432);
nor UO_2100 (O_2100,N_19874,N_19647);
nor UO_2101 (O_2101,N_19966,N_19984);
or UO_2102 (O_2102,N_19901,N_19246);
nand UO_2103 (O_2103,N_19488,N_19977);
nand UO_2104 (O_2104,N_19625,N_19597);
xor UO_2105 (O_2105,N_19834,N_19883);
or UO_2106 (O_2106,N_19221,N_19428);
nand UO_2107 (O_2107,N_19887,N_19732);
or UO_2108 (O_2108,N_19842,N_19723);
xor UO_2109 (O_2109,N_19840,N_19723);
or UO_2110 (O_2110,N_19356,N_19516);
xor UO_2111 (O_2111,N_19739,N_19436);
xnor UO_2112 (O_2112,N_19973,N_19291);
and UO_2113 (O_2113,N_19997,N_19725);
xnor UO_2114 (O_2114,N_19505,N_19327);
xor UO_2115 (O_2115,N_19854,N_19552);
and UO_2116 (O_2116,N_19279,N_19339);
or UO_2117 (O_2117,N_19344,N_19658);
and UO_2118 (O_2118,N_19390,N_19706);
nand UO_2119 (O_2119,N_19411,N_19763);
nand UO_2120 (O_2120,N_19569,N_19835);
nor UO_2121 (O_2121,N_19430,N_19960);
xor UO_2122 (O_2122,N_19246,N_19525);
nor UO_2123 (O_2123,N_19635,N_19317);
and UO_2124 (O_2124,N_19785,N_19551);
xor UO_2125 (O_2125,N_19348,N_19552);
nand UO_2126 (O_2126,N_19850,N_19308);
xor UO_2127 (O_2127,N_19816,N_19356);
nand UO_2128 (O_2128,N_19987,N_19981);
and UO_2129 (O_2129,N_19767,N_19201);
nor UO_2130 (O_2130,N_19719,N_19862);
xor UO_2131 (O_2131,N_19398,N_19905);
or UO_2132 (O_2132,N_19656,N_19321);
xor UO_2133 (O_2133,N_19356,N_19700);
nand UO_2134 (O_2134,N_19768,N_19339);
or UO_2135 (O_2135,N_19239,N_19702);
nand UO_2136 (O_2136,N_19804,N_19934);
nand UO_2137 (O_2137,N_19790,N_19440);
and UO_2138 (O_2138,N_19560,N_19855);
xnor UO_2139 (O_2139,N_19325,N_19765);
nand UO_2140 (O_2140,N_19526,N_19665);
xnor UO_2141 (O_2141,N_19665,N_19978);
xor UO_2142 (O_2142,N_19367,N_19304);
xor UO_2143 (O_2143,N_19665,N_19669);
and UO_2144 (O_2144,N_19467,N_19369);
nor UO_2145 (O_2145,N_19937,N_19812);
nand UO_2146 (O_2146,N_19716,N_19416);
nor UO_2147 (O_2147,N_19349,N_19559);
xnor UO_2148 (O_2148,N_19678,N_19711);
or UO_2149 (O_2149,N_19485,N_19428);
nor UO_2150 (O_2150,N_19511,N_19498);
nand UO_2151 (O_2151,N_19227,N_19318);
nand UO_2152 (O_2152,N_19244,N_19382);
nor UO_2153 (O_2153,N_19327,N_19902);
nor UO_2154 (O_2154,N_19915,N_19966);
nor UO_2155 (O_2155,N_19204,N_19597);
and UO_2156 (O_2156,N_19791,N_19723);
nand UO_2157 (O_2157,N_19452,N_19587);
nand UO_2158 (O_2158,N_19859,N_19332);
nand UO_2159 (O_2159,N_19212,N_19592);
or UO_2160 (O_2160,N_19809,N_19271);
nor UO_2161 (O_2161,N_19454,N_19572);
nor UO_2162 (O_2162,N_19305,N_19267);
or UO_2163 (O_2163,N_19913,N_19659);
or UO_2164 (O_2164,N_19993,N_19631);
and UO_2165 (O_2165,N_19702,N_19619);
nand UO_2166 (O_2166,N_19278,N_19432);
and UO_2167 (O_2167,N_19206,N_19310);
xor UO_2168 (O_2168,N_19699,N_19813);
or UO_2169 (O_2169,N_19289,N_19748);
nand UO_2170 (O_2170,N_19328,N_19224);
or UO_2171 (O_2171,N_19564,N_19555);
and UO_2172 (O_2172,N_19887,N_19426);
nor UO_2173 (O_2173,N_19939,N_19961);
or UO_2174 (O_2174,N_19357,N_19911);
and UO_2175 (O_2175,N_19604,N_19978);
or UO_2176 (O_2176,N_19586,N_19996);
xnor UO_2177 (O_2177,N_19228,N_19372);
nor UO_2178 (O_2178,N_19742,N_19800);
or UO_2179 (O_2179,N_19717,N_19979);
nor UO_2180 (O_2180,N_19765,N_19365);
and UO_2181 (O_2181,N_19533,N_19695);
xor UO_2182 (O_2182,N_19227,N_19225);
xor UO_2183 (O_2183,N_19466,N_19793);
and UO_2184 (O_2184,N_19935,N_19848);
and UO_2185 (O_2185,N_19639,N_19886);
or UO_2186 (O_2186,N_19917,N_19940);
or UO_2187 (O_2187,N_19767,N_19653);
nand UO_2188 (O_2188,N_19446,N_19934);
and UO_2189 (O_2189,N_19381,N_19909);
nand UO_2190 (O_2190,N_19744,N_19941);
nor UO_2191 (O_2191,N_19694,N_19340);
xor UO_2192 (O_2192,N_19540,N_19460);
or UO_2193 (O_2193,N_19242,N_19416);
nor UO_2194 (O_2194,N_19638,N_19263);
nand UO_2195 (O_2195,N_19509,N_19598);
nor UO_2196 (O_2196,N_19966,N_19463);
or UO_2197 (O_2197,N_19761,N_19702);
nand UO_2198 (O_2198,N_19832,N_19728);
nand UO_2199 (O_2199,N_19634,N_19889);
xnor UO_2200 (O_2200,N_19379,N_19969);
nor UO_2201 (O_2201,N_19439,N_19939);
and UO_2202 (O_2202,N_19783,N_19757);
nand UO_2203 (O_2203,N_19567,N_19844);
xor UO_2204 (O_2204,N_19964,N_19610);
and UO_2205 (O_2205,N_19329,N_19544);
nand UO_2206 (O_2206,N_19405,N_19837);
or UO_2207 (O_2207,N_19774,N_19546);
nor UO_2208 (O_2208,N_19690,N_19611);
or UO_2209 (O_2209,N_19558,N_19999);
xor UO_2210 (O_2210,N_19566,N_19653);
xor UO_2211 (O_2211,N_19946,N_19452);
or UO_2212 (O_2212,N_19790,N_19469);
nor UO_2213 (O_2213,N_19806,N_19314);
nor UO_2214 (O_2214,N_19486,N_19822);
nor UO_2215 (O_2215,N_19290,N_19796);
nor UO_2216 (O_2216,N_19417,N_19511);
or UO_2217 (O_2217,N_19924,N_19892);
or UO_2218 (O_2218,N_19781,N_19541);
xor UO_2219 (O_2219,N_19855,N_19503);
or UO_2220 (O_2220,N_19886,N_19663);
and UO_2221 (O_2221,N_19648,N_19845);
or UO_2222 (O_2222,N_19627,N_19311);
xnor UO_2223 (O_2223,N_19597,N_19461);
xor UO_2224 (O_2224,N_19930,N_19778);
or UO_2225 (O_2225,N_19300,N_19988);
and UO_2226 (O_2226,N_19917,N_19368);
or UO_2227 (O_2227,N_19809,N_19400);
xnor UO_2228 (O_2228,N_19200,N_19783);
or UO_2229 (O_2229,N_19478,N_19956);
and UO_2230 (O_2230,N_19714,N_19360);
and UO_2231 (O_2231,N_19782,N_19748);
nand UO_2232 (O_2232,N_19689,N_19752);
and UO_2233 (O_2233,N_19376,N_19432);
or UO_2234 (O_2234,N_19793,N_19394);
nor UO_2235 (O_2235,N_19954,N_19910);
nor UO_2236 (O_2236,N_19918,N_19242);
and UO_2237 (O_2237,N_19784,N_19907);
and UO_2238 (O_2238,N_19761,N_19883);
or UO_2239 (O_2239,N_19307,N_19707);
or UO_2240 (O_2240,N_19912,N_19890);
nand UO_2241 (O_2241,N_19574,N_19427);
xor UO_2242 (O_2242,N_19246,N_19421);
nor UO_2243 (O_2243,N_19729,N_19506);
or UO_2244 (O_2244,N_19457,N_19672);
nor UO_2245 (O_2245,N_19370,N_19709);
and UO_2246 (O_2246,N_19662,N_19574);
nand UO_2247 (O_2247,N_19818,N_19710);
and UO_2248 (O_2248,N_19319,N_19349);
and UO_2249 (O_2249,N_19275,N_19628);
nor UO_2250 (O_2250,N_19357,N_19310);
and UO_2251 (O_2251,N_19319,N_19310);
or UO_2252 (O_2252,N_19978,N_19488);
or UO_2253 (O_2253,N_19814,N_19612);
xor UO_2254 (O_2254,N_19736,N_19210);
nor UO_2255 (O_2255,N_19895,N_19821);
or UO_2256 (O_2256,N_19690,N_19485);
nand UO_2257 (O_2257,N_19386,N_19265);
or UO_2258 (O_2258,N_19929,N_19393);
and UO_2259 (O_2259,N_19202,N_19839);
xnor UO_2260 (O_2260,N_19438,N_19694);
or UO_2261 (O_2261,N_19737,N_19556);
or UO_2262 (O_2262,N_19231,N_19744);
or UO_2263 (O_2263,N_19818,N_19623);
xnor UO_2264 (O_2264,N_19836,N_19491);
nand UO_2265 (O_2265,N_19893,N_19923);
or UO_2266 (O_2266,N_19399,N_19974);
xnor UO_2267 (O_2267,N_19429,N_19770);
nand UO_2268 (O_2268,N_19606,N_19314);
nor UO_2269 (O_2269,N_19969,N_19565);
nor UO_2270 (O_2270,N_19788,N_19894);
nor UO_2271 (O_2271,N_19794,N_19565);
xor UO_2272 (O_2272,N_19293,N_19990);
nor UO_2273 (O_2273,N_19847,N_19258);
nand UO_2274 (O_2274,N_19502,N_19525);
xor UO_2275 (O_2275,N_19861,N_19511);
nand UO_2276 (O_2276,N_19565,N_19317);
and UO_2277 (O_2277,N_19814,N_19360);
and UO_2278 (O_2278,N_19913,N_19810);
and UO_2279 (O_2279,N_19409,N_19752);
nand UO_2280 (O_2280,N_19588,N_19707);
xor UO_2281 (O_2281,N_19321,N_19590);
xnor UO_2282 (O_2282,N_19952,N_19742);
and UO_2283 (O_2283,N_19931,N_19927);
and UO_2284 (O_2284,N_19834,N_19704);
or UO_2285 (O_2285,N_19997,N_19507);
nor UO_2286 (O_2286,N_19479,N_19769);
nand UO_2287 (O_2287,N_19481,N_19283);
nand UO_2288 (O_2288,N_19899,N_19577);
xnor UO_2289 (O_2289,N_19560,N_19295);
or UO_2290 (O_2290,N_19431,N_19741);
xor UO_2291 (O_2291,N_19233,N_19905);
and UO_2292 (O_2292,N_19436,N_19801);
nand UO_2293 (O_2293,N_19896,N_19945);
or UO_2294 (O_2294,N_19591,N_19362);
xor UO_2295 (O_2295,N_19287,N_19683);
nand UO_2296 (O_2296,N_19216,N_19752);
xor UO_2297 (O_2297,N_19683,N_19418);
nor UO_2298 (O_2298,N_19426,N_19641);
nand UO_2299 (O_2299,N_19847,N_19342);
nor UO_2300 (O_2300,N_19606,N_19738);
xor UO_2301 (O_2301,N_19612,N_19293);
nand UO_2302 (O_2302,N_19282,N_19974);
nand UO_2303 (O_2303,N_19772,N_19218);
and UO_2304 (O_2304,N_19319,N_19922);
xor UO_2305 (O_2305,N_19901,N_19269);
nand UO_2306 (O_2306,N_19492,N_19537);
nand UO_2307 (O_2307,N_19750,N_19680);
nand UO_2308 (O_2308,N_19694,N_19627);
nand UO_2309 (O_2309,N_19869,N_19849);
or UO_2310 (O_2310,N_19588,N_19669);
nor UO_2311 (O_2311,N_19937,N_19269);
xnor UO_2312 (O_2312,N_19633,N_19276);
and UO_2313 (O_2313,N_19728,N_19358);
xnor UO_2314 (O_2314,N_19447,N_19345);
nand UO_2315 (O_2315,N_19769,N_19634);
nand UO_2316 (O_2316,N_19268,N_19485);
xor UO_2317 (O_2317,N_19646,N_19804);
or UO_2318 (O_2318,N_19822,N_19514);
nand UO_2319 (O_2319,N_19967,N_19791);
xor UO_2320 (O_2320,N_19895,N_19549);
and UO_2321 (O_2321,N_19479,N_19300);
and UO_2322 (O_2322,N_19925,N_19856);
xnor UO_2323 (O_2323,N_19402,N_19677);
and UO_2324 (O_2324,N_19990,N_19805);
and UO_2325 (O_2325,N_19942,N_19543);
or UO_2326 (O_2326,N_19430,N_19824);
xnor UO_2327 (O_2327,N_19505,N_19800);
xnor UO_2328 (O_2328,N_19447,N_19453);
and UO_2329 (O_2329,N_19663,N_19466);
and UO_2330 (O_2330,N_19903,N_19376);
xnor UO_2331 (O_2331,N_19687,N_19442);
nand UO_2332 (O_2332,N_19503,N_19845);
nand UO_2333 (O_2333,N_19461,N_19847);
xnor UO_2334 (O_2334,N_19415,N_19678);
nor UO_2335 (O_2335,N_19916,N_19525);
xnor UO_2336 (O_2336,N_19934,N_19377);
nor UO_2337 (O_2337,N_19553,N_19600);
xnor UO_2338 (O_2338,N_19685,N_19504);
nand UO_2339 (O_2339,N_19643,N_19316);
or UO_2340 (O_2340,N_19431,N_19964);
nor UO_2341 (O_2341,N_19873,N_19856);
or UO_2342 (O_2342,N_19355,N_19273);
xor UO_2343 (O_2343,N_19505,N_19731);
nand UO_2344 (O_2344,N_19762,N_19756);
and UO_2345 (O_2345,N_19348,N_19336);
and UO_2346 (O_2346,N_19333,N_19941);
or UO_2347 (O_2347,N_19727,N_19642);
nor UO_2348 (O_2348,N_19467,N_19939);
or UO_2349 (O_2349,N_19893,N_19389);
nand UO_2350 (O_2350,N_19258,N_19616);
nand UO_2351 (O_2351,N_19390,N_19543);
nand UO_2352 (O_2352,N_19829,N_19677);
nand UO_2353 (O_2353,N_19883,N_19953);
xor UO_2354 (O_2354,N_19789,N_19346);
nand UO_2355 (O_2355,N_19920,N_19981);
nand UO_2356 (O_2356,N_19514,N_19301);
xor UO_2357 (O_2357,N_19371,N_19805);
nor UO_2358 (O_2358,N_19806,N_19490);
xor UO_2359 (O_2359,N_19867,N_19299);
nor UO_2360 (O_2360,N_19212,N_19267);
xnor UO_2361 (O_2361,N_19713,N_19686);
xnor UO_2362 (O_2362,N_19763,N_19737);
nand UO_2363 (O_2363,N_19819,N_19434);
or UO_2364 (O_2364,N_19908,N_19295);
xor UO_2365 (O_2365,N_19340,N_19982);
nand UO_2366 (O_2366,N_19564,N_19725);
xnor UO_2367 (O_2367,N_19267,N_19701);
nor UO_2368 (O_2368,N_19634,N_19300);
xnor UO_2369 (O_2369,N_19590,N_19333);
nor UO_2370 (O_2370,N_19886,N_19602);
or UO_2371 (O_2371,N_19806,N_19865);
nand UO_2372 (O_2372,N_19989,N_19727);
nor UO_2373 (O_2373,N_19788,N_19959);
or UO_2374 (O_2374,N_19635,N_19943);
or UO_2375 (O_2375,N_19605,N_19388);
nand UO_2376 (O_2376,N_19945,N_19321);
nor UO_2377 (O_2377,N_19331,N_19737);
and UO_2378 (O_2378,N_19896,N_19506);
or UO_2379 (O_2379,N_19802,N_19563);
nand UO_2380 (O_2380,N_19263,N_19580);
nor UO_2381 (O_2381,N_19471,N_19407);
xor UO_2382 (O_2382,N_19814,N_19303);
xnor UO_2383 (O_2383,N_19248,N_19802);
nor UO_2384 (O_2384,N_19403,N_19910);
or UO_2385 (O_2385,N_19882,N_19986);
nor UO_2386 (O_2386,N_19754,N_19263);
and UO_2387 (O_2387,N_19735,N_19719);
nor UO_2388 (O_2388,N_19829,N_19536);
or UO_2389 (O_2389,N_19790,N_19521);
nor UO_2390 (O_2390,N_19711,N_19318);
or UO_2391 (O_2391,N_19440,N_19728);
or UO_2392 (O_2392,N_19965,N_19561);
xor UO_2393 (O_2393,N_19207,N_19741);
nand UO_2394 (O_2394,N_19460,N_19870);
nand UO_2395 (O_2395,N_19270,N_19378);
xor UO_2396 (O_2396,N_19286,N_19394);
nand UO_2397 (O_2397,N_19423,N_19803);
nand UO_2398 (O_2398,N_19281,N_19925);
xnor UO_2399 (O_2399,N_19636,N_19393);
nand UO_2400 (O_2400,N_19517,N_19757);
nand UO_2401 (O_2401,N_19598,N_19551);
and UO_2402 (O_2402,N_19450,N_19992);
or UO_2403 (O_2403,N_19682,N_19996);
nand UO_2404 (O_2404,N_19864,N_19312);
and UO_2405 (O_2405,N_19220,N_19764);
nor UO_2406 (O_2406,N_19861,N_19409);
or UO_2407 (O_2407,N_19777,N_19351);
or UO_2408 (O_2408,N_19530,N_19598);
or UO_2409 (O_2409,N_19906,N_19730);
and UO_2410 (O_2410,N_19603,N_19968);
or UO_2411 (O_2411,N_19532,N_19841);
or UO_2412 (O_2412,N_19392,N_19425);
and UO_2413 (O_2413,N_19925,N_19564);
nor UO_2414 (O_2414,N_19923,N_19965);
or UO_2415 (O_2415,N_19345,N_19618);
nor UO_2416 (O_2416,N_19998,N_19567);
nand UO_2417 (O_2417,N_19348,N_19640);
nand UO_2418 (O_2418,N_19358,N_19471);
or UO_2419 (O_2419,N_19326,N_19548);
nand UO_2420 (O_2420,N_19646,N_19879);
or UO_2421 (O_2421,N_19413,N_19768);
nor UO_2422 (O_2422,N_19444,N_19724);
nand UO_2423 (O_2423,N_19450,N_19712);
xor UO_2424 (O_2424,N_19278,N_19650);
nand UO_2425 (O_2425,N_19930,N_19890);
nor UO_2426 (O_2426,N_19975,N_19780);
nand UO_2427 (O_2427,N_19723,N_19879);
nand UO_2428 (O_2428,N_19818,N_19831);
nor UO_2429 (O_2429,N_19645,N_19492);
or UO_2430 (O_2430,N_19402,N_19235);
or UO_2431 (O_2431,N_19359,N_19238);
or UO_2432 (O_2432,N_19762,N_19352);
xor UO_2433 (O_2433,N_19736,N_19413);
nand UO_2434 (O_2434,N_19427,N_19510);
or UO_2435 (O_2435,N_19818,N_19860);
nand UO_2436 (O_2436,N_19408,N_19667);
or UO_2437 (O_2437,N_19631,N_19355);
and UO_2438 (O_2438,N_19376,N_19283);
xnor UO_2439 (O_2439,N_19863,N_19771);
nor UO_2440 (O_2440,N_19834,N_19835);
or UO_2441 (O_2441,N_19383,N_19284);
nand UO_2442 (O_2442,N_19949,N_19220);
nand UO_2443 (O_2443,N_19909,N_19949);
xnor UO_2444 (O_2444,N_19306,N_19473);
xor UO_2445 (O_2445,N_19286,N_19493);
and UO_2446 (O_2446,N_19588,N_19642);
xnor UO_2447 (O_2447,N_19890,N_19900);
or UO_2448 (O_2448,N_19802,N_19624);
and UO_2449 (O_2449,N_19909,N_19278);
nor UO_2450 (O_2450,N_19309,N_19950);
or UO_2451 (O_2451,N_19944,N_19756);
nand UO_2452 (O_2452,N_19281,N_19365);
nor UO_2453 (O_2453,N_19683,N_19582);
or UO_2454 (O_2454,N_19740,N_19517);
and UO_2455 (O_2455,N_19544,N_19312);
nor UO_2456 (O_2456,N_19688,N_19487);
or UO_2457 (O_2457,N_19244,N_19751);
or UO_2458 (O_2458,N_19878,N_19329);
xnor UO_2459 (O_2459,N_19686,N_19205);
xor UO_2460 (O_2460,N_19636,N_19451);
xnor UO_2461 (O_2461,N_19264,N_19740);
xor UO_2462 (O_2462,N_19794,N_19382);
nand UO_2463 (O_2463,N_19839,N_19499);
nand UO_2464 (O_2464,N_19756,N_19683);
nand UO_2465 (O_2465,N_19723,N_19359);
xnor UO_2466 (O_2466,N_19531,N_19806);
nand UO_2467 (O_2467,N_19647,N_19604);
or UO_2468 (O_2468,N_19919,N_19414);
nor UO_2469 (O_2469,N_19768,N_19449);
and UO_2470 (O_2470,N_19466,N_19393);
nand UO_2471 (O_2471,N_19557,N_19606);
nor UO_2472 (O_2472,N_19869,N_19723);
nor UO_2473 (O_2473,N_19437,N_19378);
and UO_2474 (O_2474,N_19241,N_19521);
nor UO_2475 (O_2475,N_19618,N_19710);
nor UO_2476 (O_2476,N_19776,N_19228);
nand UO_2477 (O_2477,N_19330,N_19406);
xnor UO_2478 (O_2478,N_19706,N_19556);
xor UO_2479 (O_2479,N_19496,N_19639);
and UO_2480 (O_2480,N_19923,N_19600);
xor UO_2481 (O_2481,N_19253,N_19999);
nand UO_2482 (O_2482,N_19218,N_19960);
xor UO_2483 (O_2483,N_19598,N_19244);
xnor UO_2484 (O_2484,N_19694,N_19322);
nor UO_2485 (O_2485,N_19840,N_19620);
nand UO_2486 (O_2486,N_19812,N_19229);
xnor UO_2487 (O_2487,N_19561,N_19903);
nand UO_2488 (O_2488,N_19545,N_19790);
and UO_2489 (O_2489,N_19586,N_19624);
or UO_2490 (O_2490,N_19511,N_19636);
xnor UO_2491 (O_2491,N_19649,N_19864);
and UO_2492 (O_2492,N_19951,N_19351);
or UO_2493 (O_2493,N_19853,N_19998);
nor UO_2494 (O_2494,N_19676,N_19925);
nand UO_2495 (O_2495,N_19705,N_19254);
and UO_2496 (O_2496,N_19320,N_19433);
nor UO_2497 (O_2497,N_19462,N_19880);
nand UO_2498 (O_2498,N_19325,N_19315);
and UO_2499 (O_2499,N_19958,N_19743);
endmodule