module basic_5000_50000_5000_25_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_2830,In_1368);
or U1 (N_1,In_3919,In_4154);
or U2 (N_2,In_3754,In_3523);
and U3 (N_3,In_1962,In_2184);
or U4 (N_4,In_2577,In_3413);
and U5 (N_5,In_546,In_1554);
xnor U6 (N_6,In_465,In_1216);
and U7 (N_7,In_464,In_3942);
and U8 (N_8,In_4663,In_4373);
nand U9 (N_9,In_335,In_72);
and U10 (N_10,In_2688,In_3908);
or U11 (N_11,In_4912,In_4699);
nand U12 (N_12,In_664,In_901);
and U13 (N_13,In_3612,In_2485);
nor U14 (N_14,In_543,In_1741);
nand U15 (N_15,In_1266,In_2095);
nand U16 (N_16,In_979,In_4956);
xnor U17 (N_17,In_324,In_2806);
nor U18 (N_18,In_3801,In_3780);
nand U19 (N_19,In_1691,In_4950);
and U20 (N_20,In_646,In_4113);
or U21 (N_21,In_3405,In_3731);
and U22 (N_22,In_2244,In_2356);
nor U23 (N_23,In_2934,In_2382);
and U24 (N_24,In_4039,In_1394);
and U25 (N_25,In_508,In_2080);
xor U26 (N_26,In_568,In_1870);
xor U27 (N_27,In_1446,In_2833);
xnor U28 (N_28,In_2372,In_3603);
nand U29 (N_29,In_331,In_751);
and U30 (N_30,In_4429,In_1518);
nor U31 (N_31,In_4733,In_1573);
and U32 (N_32,In_2627,In_2667);
xor U33 (N_33,In_4461,In_3417);
nor U34 (N_34,In_484,In_2735);
xor U35 (N_35,In_1708,In_174);
nor U36 (N_36,In_3890,In_3522);
xnor U37 (N_37,In_1445,In_4855);
nor U38 (N_38,In_2840,In_68);
nand U39 (N_39,In_4693,In_4169);
nor U40 (N_40,In_1560,In_303);
nor U41 (N_41,In_4451,In_2046);
nor U42 (N_42,In_2413,In_2314);
and U43 (N_43,In_4657,In_827);
or U44 (N_44,In_3727,In_1316);
nand U45 (N_45,In_1010,In_4807);
nor U46 (N_46,In_4999,In_24);
nor U47 (N_47,In_2203,In_349);
xor U48 (N_48,In_4653,In_551);
or U49 (N_49,In_3956,In_1537);
or U50 (N_50,In_2621,In_934);
nor U51 (N_51,In_559,In_1339);
xnor U52 (N_52,In_1855,In_826);
and U53 (N_53,In_1956,In_4862);
or U54 (N_54,In_169,In_2752);
and U55 (N_55,In_1884,In_1521);
and U56 (N_56,In_3006,In_1452);
and U57 (N_57,In_3810,In_3602);
nor U58 (N_58,In_4035,In_55);
xor U59 (N_59,In_3836,In_2994);
nor U60 (N_60,In_3569,In_3207);
nor U61 (N_61,In_2003,In_3001);
and U62 (N_62,In_1981,In_1584);
nor U63 (N_63,In_2072,In_986);
nor U64 (N_64,In_2373,In_3752);
nand U65 (N_65,In_812,In_3251);
and U66 (N_66,In_1666,In_4059);
and U67 (N_67,In_4412,In_645);
or U68 (N_68,In_4201,In_356);
or U69 (N_69,In_2639,In_1681);
nor U70 (N_70,In_2176,In_4055);
xnor U71 (N_71,In_1373,In_4941);
or U72 (N_72,In_696,In_4929);
nor U73 (N_73,In_2583,In_4215);
or U74 (N_74,In_1044,In_3667);
and U75 (N_75,In_2554,In_710);
nor U76 (N_76,In_1556,In_2034);
nor U77 (N_77,In_3005,In_1346);
nor U78 (N_78,In_2792,In_2324);
xor U79 (N_79,In_2596,In_3046);
nor U80 (N_80,In_4274,In_3357);
or U81 (N_81,In_3722,In_1916);
nor U82 (N_82,In_3802,In_2452);
and U83 (N_83,In_4625,In_4174);
xor U84 (N_84,In_872,In_1564);
and U85 (N_85,In_2993,In_2468);
nor U86 (N_86,In_4641,In_3600);
nand U87 (N_87,In_4046,In_4649);
and U88 (N_88,In_4462,In_3534);
and U89 (N_89,In_351,In_3305);
or U90 (N_90,In_3837,In_1931);
nand U91 (N_91,In_3137,In_563);
nor U92 (N_92,In_2855,In_1615);
or U93 (N_93,In_4435,In_3187);
or U94 (N_94,In_1866,In_1910);
or U95 (N_95,In_4717,In_1350);
and U96 (N_96,In_659,In_3293);
nor U97 (N_97,In_2876,In_1110);
xnor U98 (N_98,In_1430,In_4980);
nand U99 (N_99,In_1317,In_3394);
nand U100 (N_100,In_1811,In_3610);
and U101 (N_101,In_3817,In_3323);
and U102 (N_102,In_660,In_1798);
or U103 (N_103,In_1186,In_3396);
nor U104 (N_104,In_2676,In_3010);
nand U105 (N_105,In_4379,In_3247);
and U106 (N_106,In_3052,In_151);
nor U107 (N_107,In_1450,In_3376);
or U108 (N_108,In_126,In_3281);
nand U109 (N_109,In_3732,In_4193);
or U110 (N_110,In_435,In_1765);
nor U111 (N_111,In_760,In_565);
nand U112 (N_112,In_1619,In_1550);
or U113 (N_113,In_2649,In_238);
nand U114 (N_114,In_1248,In_658);
and U115 (N_115,In_3130,In_3432);
nand U116 (N_116,In_2817,In_3658);
and U117 (N_117,In_2240,In_3232);
nand U118 (N_118,In_2843,In_4425);
nor U119 (N_119,In_713,In_4365);
nor U120 (N_120,In_1764,In_3313);
or U121 (N_121,In_3133,In_4991);
nor U122 (N_122,In_2954,In_3451);
xnor U123 (N_123,In_1012,In_2943);
xnor U124 (N_124,In_1868,In_65);
nand U125 (N_125,In_2776,In_3548);
nor U126 (N_126,In_2499,In_4590);
and U127 (N_127,In_2559,In_4027);
or U128 (N_128,In_2337,In_2248);
or U129 (N_129,In_3079,In_130);
nor U130 (N_130,In_798,In_2063);
xnor U131 (N_131,In_1571,In_3123);
or U132 (N_132,In_4553,In_2487);
xor U133 (N_133,In_1008,In_813);
xor U134 (N_134,In_4220,In_3876);
xor U135 (N_135,In_572,In_1380);
nor U136 (N_136,In_1662,In_2055);
xor U137 (N_137,In_1586,In_1635);
nor U138 (N_138,In_3103,In_1502);
nor U139 (N_139,In_687,In_137);
or U140 (N_140,In_2174,In_3438);
nand U141 (N_141,In_2541,In_404);
nand U142 (N_142,In_1436,In_900);
nor U143 (N_143,In_866,In_4967);
or U144 (N_144,In_946,In_1228);
or U145 (N_145,In_3547,In_3389);
xnor U146 (N_146,In_1656,In_3974);
nor U147 (N_147,In_2040,In_433);
and U148 (N_148,In_1021,In_1014);
and U149 (N_149,In_3341,In_4995);
or U150 (N_150,In_4445,In_4253);
nor U151 (N_151,In_896,In_3833);
xnor U152 (N_152,In_1906,In_4575);
nor U153 (N_153,In_1355,In_3120);
nand U154 (N_154,In_2909,In_374);
nor U155 (N_155,In_2368,In_466);
xnor U156 (N_156,In_1019,In_4847);
xnor U157 (N_157,In_3820,In_4196);
nand U158 (N_158,In_4008,In_679);
nor U159 (N_159,In_53,In_4391);
or U160 (N_160,In_1908,In_3073);
xnor U161 (N_161,In_4987,In_3088);
xnor U162 (N_162,In_1041,In_66);
or U163 (N_163,In_4831,In_1678);
nand U164 (N_164,In_903,In_1877);
and U165 (N_165,In_67,In_4233);
nand U166 (N_166,In_3711,In_1623);
nand U167 (N_167,In_3664,In_3866);
nor U168 (N_168,In_3044,In_852);
and U169 (N_169,In_2326,In_4061);
xnor U170 (N_170,In_2210,In_2771);
nand U171 (N_171,In_1580,In_1022);
and U172 (N_172,In_2050,In_412);
or U173 (N_173,In_1152,In_4191);
xnor U174 (N_174,In_1314,In_109);
xor U175 (N_175,In_4030,In_1141);
nand U176 (N_176,In_2866,In_4789);
nor U177 (N_177,In_978,In_98);
or U178 (N_178,In_4014,In_1509);
or U179 (N_179,In_4994,In_69);
xnor U180 (N_180,In_1887,In_3984);
and U181 (N_181,In_1807,In_544);
nand U182 (N_182,In_792,In_4838);
and U183 (N_183,In_712,In_4514);
nor U184 (N_184,In_1092,In_3374);
and U185 (N_185,In_4845,In_614);
or U186 (N_186,In_3373,In_1304);
or U187 (N_187,In_3578,In_1805);
and U188 (N_188,In_2286,In_737);
and U189 (N_189,In_4841,In_384);
or U190 (N_190,In_796,In_3352);
or U191 (N_191,In_236,In_234);
or U192 (N_192,In_2344,In_1118);
or U193 (N_193,In_4345,In_2638);
nand U194 (N_194,In_4777,In_3690);
xor U195 (N_195,In_1082,In_4778);
and U196 (N_196,In_2364,In_4763);
or U197 (N_197,In_1832,In_319);
nor U198 (N_198,In_778,In_1786);
or U199 (N_199,In_592,In_3433);
nand U200 (N_200,In_2411,In_1453);
and U201 (N_201,In_3979,In_3440);
or U202 (N_202,In_2647,In_1848);
nor U203 (N_203,In_3470,In_2133);
xor U204 (N_204,In_4993,In_2572);
nor U205 (N_205,In_123,In_2762);
or U206 (N_206,In_164,In_3430);
or U207 (N_207,In_2631,In_1511);
nand U208 (N_208,In_1193,In_2233);
nor U209 (N_209,In_2673,In_3717);
xnor U210 (N_210,In_2699,In_4977);
or U211 (N_211,In_393,In_4892);
and U212 (N_212,In_1323,In_652);
and U213 (N_213,In_131,In_2228);
and U214 (N_214,In_266,In_36);
or U215 (N_215,In_3144,In_4604);
nor U216 (N_216,In_1361,In_4739);
or U217 (N_217,In_3228,In_4546);
xnor U218 (N_218,In_596,In_1227);
xor U219 (N_219,In_4137,In_3560);
or U220 (N_220,In_4949,In_283);
xor U221 (N_221,In_3962,In_3702);
or U222 (N_222,In_1169,In_4548);
nand U223 (N_223,In_2779,In_265);
nand U224 (N_224,In_275,In_3307);
or U225 (N_225,In_941,In_580);
nand U226 (N_226,In_537,In_341);
xnor U227 (N_227,In_4563,In_3925);
nand U228 (N_228,In_1559,In_4745);
or U229 (N_229,In_2440,In_2071);
xor U230 (N_230,In_3290,In_2462);
or U231 (N_231,In_3819,In_4818);
nor U232 (N_232,In_4923,In_4367);
nand U233 (N_233,In_2507,In_1555);
nand U234 (N_234,In_4782,In_401);
or U235 (N_235,In_4348,In_4051);
and U236 (N_236,In_110,In_322);
nor U237 (N_237,In_1828,In_2097);
nor U238 (N_238,In_761,In_4655);
and U239 (N_239,In_992,In_3544);
nor U240 (N_240,In_1911,In_2933);
nor U241 (N_241,In_2861,In_4427);
nand U242 (N_242,In_775,In_180);
or U243 (N_243,In_2802,In_3511);
nand U244 (N_244,In_663,In_1609);
nand U245 (N_245,In_1028,In_4695);
nand U246 (N_246,In_2006,In_133);
nand U247 (N_247,In_1922,In_4002);
xor U248 (N_248,In_945,In_420);
nor U249 (N_249,In_816,In_1163);
and U250 (N_250,In_3265,In_2796);
xor U251 (N_251,In_239,In_73);
and U252 (N_252,In_2092,In_1995);
and U253 (N_253,In_4869,In_529);
nand U254 (N_254,In_2813,In_1597);
xor U255 (N_255,In_3788,In_911);
nor U256 (N_256,In_1837,In_994);
xor U257 (N_257,In_2265,In_2053);
nor U258 (N_258,In_3277,In_1729);
or U259 (N_259,In_2982,In_2853);
nand U260 (N_260,In_3982,In_1204);
and U261 (N_261,In_3173,In_163);
nand U262 (N_262,In_3109,In_1064);
nand U263 (N_263,In_973,In_2508);
xnor U264 (N_264,In_116,In_4084);
and U265 (N_265,In_1326,In_121);
nor U266 (N_266,In_3528,In_1252);
xor U267 (N_267,In_2640,In_3028);
and U268 (N_268,In_2010,In_1347);
nor U269 (N_269,In_1251,In_286);
nand U270 (N_270,In_1410,In_860);
or U271 (N_271,In_3842,In_4765);
xnor U272 (N_272,In_4606,In_743);
nand U273 (N_273,In_1812,In_2293);
and U274 (N_274,In_897,In_4492);
or U275 (N_275,In_1234,In_1246);
nor U276 (N_276,In_918,In_1310);
and U277 (N_277,In_1171,In_3666);
nor U278 (N_278,In_1184,In_3991);
xor U279 (N_279,In_1257,In_4431);
or U280 (N_280,In_1864,In_959);
and U281 (N_281,In_4981,In_2295);
or U282 (N_282,In_3889,In_2680);
nand U283 (N_283,In_1135,In_2378);
xnor U284 (N_284,In_410,In_3827);
and U285 (N_285,In_3076,In_1481);
nand U286 (N_286,In_4172,In_1582);
xor U287 (N_287,In_666,In_2675);
and U288 (N_288,In_779,In_1224);
and U289 (N_289,In_253,In_617);
or U290 (N_290,In_2835,In_226);
and U291 (N_291,In_3695,In_1723);
or U292 (N_292,In_2886,In_2513);
nand U293 (N_293,In_357,In_1484);
nand U294 (N_294,In_667,In_1756);
or U295 (N_295,In_721,In_3342);
nor U296 (N_296,In_1005,In_2717);
xnor U297 (N_297,In_1682,In_746);
nand U298 (N_298,In_3682,In_2907);
and U299 (N_299,In_4735,In_3572);
nor U300 (N_300,In_2304,In_152);
or U301 (N_301,In_321,In_3983);
and U302 (N_302,In_2795,In_1414);
or U303 (N_303,In_561,In_1099);
or U304 (N_304,In_2266,In_1547);
or U305 (N_305,In_1567,In_3390);
nor U306 (N_306,In_8,In_78);
nor U307 (N_307,In_380,In_4226);
nand U308 (N_308,In_4293,In_2791);
nand U309 (N_309,In_3857,In_274);
xnor U310 (N_310,In_4885,In_1338);
nor U311 (N_311,In_2463,In_1267);
nor U312 (N_312,In_216,In_3096);
nand U313 (N_313,In_3854,In_3240);
nor U314 (N_314,In_719,In_3897);
and U315 (N_315,In_3038,In_558);
and U316 (N_316,In_367,In_1800);
xor U317 (N_317,In_4578,In_1164);
or U318 (N_318,In_183,In_1468);
and U319 (N_319,In_2536,In_2239);
and U320 (N_320,In_1492,In_280);
nand U321 (N_321,In_1987,In_4743);
nand U322 (N_322,In_2325,In_1102);
nor U323 (N_323,In_1989,In_241);
or U324 (N_324,In_1188,In_4296);
nor U325 (N_325,In_1083,In_2697);
or U326 (N_326,In_4985,In_1086);
or U327 (N_327,In_364,In_3315);
nand U328 (N_328,In_4775,In_1695);
nand U329 (N_329,In_4100,In_3985);
xor U330 (N_330,In_403,In_434);
nor U331 (N_331,In_1694,In_2575);
and U332 (N_332,In_201,In_947);
xnor U333 (N_333,In_3199,In_2571);
xnor U334 (N_334,In_2026,In_1401);
or U335 (N_335,In_1231,In_1552);
xor U336 (N_336,In_1944,In_2429);
and U337 (N_337,In_4132,In_3498);
xor U338 (N_338,In_2439,In_2610);
nor U339 (N_339,In_3204,In_2759);
nand U340 (N_340,In_3420,In_4727);
or U341 (N_341,In_3224,In_4890);
nor U342 (N_342,In_2051,In_505);
and U343 (N_343,In_974,In_1824);
nor U344 (N_344,In_1890,In_1668);
nor U345 (N_345,In_2637,In_4607);
and U346 (N_346,In_4957,In_2811);
nor U347 (N_347,In_2476,In_4840);
or U348 (N_348,In_37,In_4635);
and U349 (N_349,In_2885,In_103);
and U350 (N_350,In_79,In_4183);
nor U351 (N_351,In_962,In_2171);
xor U352 (N_352,In_542,In_1485);
or U353 (N_353,In_3512,In_4403);
and U354 (N_354,In_3351,In_2729);
and U355 (N_355,In_1438,In_379);
xnor U356 (N_356,In_3481,In_1624);
nand U357 (N_357,In_608,In_4126);
and U358 (N_358,In_1639,In_4009);
and U359 (N_359,In_1396,In_3720);
and U360 (N_360,In_2770,In_114);
nor U361 (N_361,In_4145,In_1979);
nor U362 (N_362,In_1035,In_2267);
and U363 (N_363,In_804,In_514);
nor U364 (N_364,In_1031,In_4134);
nand U365 (N_365,In_4698,In_3879);
xor U366 (N_366,In_3861,In_1051);
nand U367 (N_367,In_886,In_2854);
nand U368 (N_368,In_4013,In_3589);
xnor U369 (N_369,In_4438,In_1230);
xor U370 (N_370,In_1449,In_4771);
xor U371 (N_371,In_692,In_647);
or U372 (N_372,In_4263,In_1185);
xnor U373 (N_373,In_1200,In_200);
and U374 (N_374,In_3264,In_3607);
xor U375 (N_375,In_3410,In_2427);
xor U376 (N_376,In_4651,In_3742);
nand U377 (N_377,In_3852,In_522);
or U378 (N_378,In_1318,In_4023);
or U379 (N_379,In_2589,In_2607);
and U380 (N_380,In_1969,In_2951);
nand U381 (N_381,In_1149,In_4025);
nand U382 (N_382,In_2415,In_4407);
and U383 (N_383,In_28,In_4268);
or U384 (N_384,In_3118,In_377);
or U385 (N_385,In_1120,In_413);
and U386 (N_386,In_285,In_2871);
nand U387 (N_387,In_4768,In_2942);
and U388 (N_388,In_4489,In_1775);
or U389 (N_389,In_1545,In_656);
xnor U390 (N_390,In_3423,In_4910);
or U391 (N_391,In_3104,In_4908);
and U392 (N_392,In_1205,In_3762);
nor U393 (N_393,In_4754,In_3435);
nor U394 (N_394,In_988,In_3282);
xor U395 (N_395,In_3506,In_4372);
and U396 (N_396,In_1797,In_4654);
xnor U397 (N_397,In_3392,In_968);
nand U398 (N_398,In_1458,In_1050);
or U399 (N_399,In_2570,In_4378);
nor U400 (N_400,In_3053,In_3995);
nor U401 (N_401,In_156,In_3214);
nor U402 (N_402,In_52,In_4866);
or U403 (N_403,In_738,In_1264);
or U404 (N_404,In_553,In_125);
nor U405 (N_405,In_398,In_2135);
xnor U406 (N_406,In_995,In_540);
xor U407 (N_407,In_3625,In_4482);
or U408 (N_408,In_1148,In_2101);
nor U409 (N_409,In_1080,In_2319);
nor U410 (N_410,In_1535,In_1875);
or U411 (N_411,In_1119,In_1007);
nor U412 (N_412,In_4064,In_970);
nand U413 (N_413,In_1867,In_4404);
nand U414 (N_414,In_3441,In_936);
nor U415 (N_415,In_4617,In_1469);
xnor U416 (N_416,In_924,In_1479);
nand U417 (N_417,In_3507,In_4725);
or U418 (N_418,In_4110,In_1663);
xnor U419 (N_419,In_390,In_3784);
and U420 (N_420,In_3227,In_1651);
xor U421 (N_421,In_4162,In_3393);
or U422 (N_422,In_477,In_869);
and U423 (N_423,In_4012,In_459);
nand U424 (N_424,In_1829,In_3713);
nand U425 (N_425,In_0,In_248);
xnor U426 (N_426,In_3132,In_3310);
nand U427 (N_427,In_4401,In_1351);
xnor U428 (N_428,In_3851,In_2549);
or U429 (N_429,In_3475,In_4609);
and U430 (N_430,In_4481,In_1899);
and U431 (N_431,In_429,In_3673);
nand U432 (N_432,In_3508,In_1079);
nand U433 (N_433,In_2038,In_3033);
or U434 (N_434,In_4202,In_1255);
and U435 (N_435,In_1863,In_3346);
and U436 (N_436,In_3031,In_1871);
or U437 (N_437,In_1679,In_4082);
xnor U438 (N_438,In_2859,In_1094);
or U439 (N_439,In_4177,In_4670);
nand U440 (N_440,In_4779,In_3561);
xor U441 (N_441,In_4369,In_14);
and U442 (N_442,In_1256,In_2901);
or U443 (N_443,In_2446,In_4032);
nand U444 (N_444,In_4368,In_4581);
nand U445 (N_445,In_3609,In_3909);
nand U446 (N_446,In_925,In_2720);
xnor U447 (N_447,In_1690,In_832);
and U448 (N_448,In_3841,In_2109);
or U449 (N_449,In_2363,In_4095);
xor U450 (N_450,In_3447,In_2482);
nand U451 (N_451,In_651,In_2122);
and U452 (N_452,In_772,In_3409);
nor U453 (N_453,In_4219,In_727);
nand U454 (N_454,In_4668,In_1707);
nand U455 (N_455,In_1324,In_4824);
and U456 (N_456,In_4286,In_3115);
nand U457 (N_457,In_2355,In_3633);
xnor U458 (N_458,In_4120,In_4494);
nand U459 (N_459,In_2469,In_2067);
nand U460 (N_460,In_1773,In_1561);
xnor U461 (N_461,In_1375,In_1577);
or U462 (N_462,In_2312,In_3238);
and U463 (N_463,In_4602,In_3270);
xnor U464 (N_464,In_2810,In_4038);
xor U465 (N_465,In_1610,In_770);
nand U466 (N_466,In_823,In_4875);
or U467 (N_467,In_1980,In_3621);
and U468 (N_468,In_613,In_383);
nor U469 (N_469,In_1813,In_2851);
nor U470 (N_470,In_1293,In_2022);
xor U471 (N_471,In_1676,In_1859);
xnor U472 (N_472,In_4969,In_287);
nor U473 (N_473,In_4128,In_510);
xnor U474 (N_474,In_4229,In_209);
xor U475 (N_475,In_4280,In_528);
xor U476 (N_476,In_1857,In_310);
nor U477 (N_477,In_707,In_4246);
and U478 (N_478,In_3617,In_1287);
xnor U479 (N_479,In_3023,In_2609);
xor U480 (N_480,In_3198,In_3008);
nor U481 (N_481,In_1886,In_1367);
or U482 (N_482,In_3386,In_4351);
and U483 (N_483,In_399,In_3129);
or U484 (N_484,In_586,In_32);
xnor U485 (N_485,In_1942,In_2009);
xor U486 (N_486,In_2070,In_3733);
nor U487 (N_487,In_2908,In_2395);
or U488 (N_488,In_1596,In_744);
or U489 (N_489,In_352,In_175);
nand U490 (N_490,In_1958,In_3896);
nor U491 (N_491,In_2023,In_2564);
nor U492 (N_492,In_4256,In_601);
and U493 (N_493,In_439,In_4982);
or U494 (N_494,In_3941,In_2480);
nor U495 (N_495,In_2271,In_1229);
and U496 (N_496,In_4118,In_1054);
and U497 (N_497,In_1187,In_4135);
and U498 (N_498,In_3689,In_899);
xnor U499 (N_499,In_483,In_913);
and U500 (N_500,In_4886,In_576);
or U501 (N_501,In_1365,In_3099);
or U502 (N_502,In_1175,In_1476);
xor U503 (N_503,In_4676,In_1342);
nor U504 (N_504,In_3007,In_1661);
or U505 (N_505,In_1644,In_1312);
nand U506 (N_506,In_3233,In_4837);
nor U507 (N_507,In_1768,In_1011);
or U508 (N_508,In_3479,In_3808);
nor U509 (N_509,In_445,In_574);
and U510 (N_510,In_4466,In_2361);
or U511 (N_511,In_168,In_4340);
xor U512 (N_512,In_4021,In_4611);
nand U513 (N_513,In_488,In_4656);
or U514 (N_514,In_1751,In_1975);
nor U515 (N_515,In_1945,In_1512);
nand U516 (N_516,In_4488,In_3112);
nor U517 (N_517,In_3834,In_33);
xnor U518 (N_518,In_208,In_4562);
or U519 (N_519,In_2606,In_4976);
xor U520 (N_520,In_3904,In_2166);
nor U521 (N_521,In_3218,In_3627);
nand U522 (N_522,In_1904,In_4951);
and U523 (N_523,In_952,In_1387);
or U524 (N_524,In_3712,In_1563);
xor U525 (N_525,In_4070,In_1075);
or U526 (N_526,In_3935,In_3570);
or U527 (N_527,In_3710,In_550);
and U528 (N_528,In_961,In_402);
nand U529 (N_529,In_4278,In_1617);
and U530 (N_530,In_4496,In_3906);
nand U531 (N_531,In_2448,In_953);
nor U532 (N_532,In_3573,In_1456);
xnor U533 (N_533,In_837,In_3792);
nand U534 (N_534,In_2497,In_3697);
and U535 (N_535,In_780,In_10);
nand U536 (N_536,In_371,In_3737);
and U537 (N_537,In_754,In_4502);
and U538 (N_538,In_2490,In_2409);
and U539 (N_539,In_2535,In_4047);
and U540 (N_540,In_4130,In_683);
and U541 (N_541,In_4585,In_4330);
nor U542 (N_542,In_2927,In_1730);
xnor U543 (N_543,In_2175,In_942);
nand U544 (N_544,In_1898,In_346);
nand U545 (N_545,In_2626,In_3986);
nor U546 (N_546,In_495,In_3626);
and U547 (N_547,In_378,In_2658);
nor U548 (N_548,In_381,In_2595);
or U549 (N_549,In_2579,In_1631);
and U550 (N_550,In_4865,In_950);
or U551 (N_551,In_4190,In_1846);
nor U552 (N_552,In_4141,In_140);
or U553 (N_553,In_1745,In_1191);
nand U554 (N_554,In_3514,In_4323);
nor U555 (N_555,In_4127,In_4063);
xor U556 (N_556,In_1081,In_3895);
xor U557 (N_557,In_1687,In_2986);
nor U558 (N_558,In_1132,In_3442);
and U559 (N_559,In_4687,In_4769);
xnor U560 (N_560,In_931,In_1462);
and U561 (N_561,In_4241,In_222);
or U562 (N_562,In_3994,In_425);
nand U563 (N_563,In_1033,In_3755);
nand U564 (N_564,In_3158,In_2726);
and U565 (N_565,In_1091,In_1718);
or U566 (N_566,In_1974,In_2170);
nor U567 (N_567,In_3546,In_2785);
nand U568 (N_568,In_4747,In_2523);
nand U569 (N_569,In_636,In_2105);
or U570 (N_570,In_2212,In_2632);
or U571 (N_571,In_1024,In_4526);
and U572 (N_572,In_4097,In_44);
xor U573 (N_573,In_62,In_2450);
nand U574 (N_574,In_1771,In_4261);
nor U575 (N_575,In_4164,In_2090);
xor U576 (N_576,In_1814,In_4478);
or U577 (N_577,In_4983,In_300);
nand U578 (N_578,In_4920,In_722);
or U579 (N_579,In_2628,In_4473);
xor U580 (N_580,In_1105,In_2903);
nand U581 (N_581,In_4531,In_2689);
and U582 (N_582,In_3237,In_3131);
nor U583 (N_583,In_4123,In_2033);
and U584 (N_584,In_88,In_2983);
and U585 (N_585,In_2939,In_1461);
or U586 (N_586,In_1451,In_249);
and U587 (N_587,In_1540,In_1601);
nor U588 (N_588,In_142,In_2511);
and U589 (N_589,In_585,In_4092);
nor U590 (N_590,In_3778,In_2309);
and U591 (N_591,In_3964,In_785);
xor U592 (N_592,In_4416,In_874);
and U593 (N_593,In_3456,In_2397);
nand U594 (N_594,In_3723,In_1440);
and U595 (N_595,In_2459,In_276);
or U596 (N_596,In_1830,In_3165);
nor U597 (N_597,In_3990,In_4255);
or U598 (N_598,In_4387,In_4813);
xnor U599 (N_599,In_124,In_4895);
xnor U600 (N_600,In_1116,In_2617);
and U601 (N_601,In_1858,In_4458);
and U602 (N_602,In_3094,In_2932);
or U603 (N_603,In_3554,In_1850);
and U604 (N_604,In_3659,In_3358);
nand U605 (N_605,In_2576,In_2778);
and U606 (N_606,In_3337,In_1994);
and U607 (N_607,In_1499,In_2809);
nand U608 (N_608,In_2891,In_4393);
nand U609 (N_609,In_702,In_4307);
or U610 (N_610,In_3708,In_2527);
and U611 (N_611,In_4184,In_4430);
or U612 (N_612,In_4223,In_2844);
nand U613 (N_613,In_3412,In_626);
nand U614 (N_614,In_2352,In_2198);
nand U615 (N_615,In_1591,In_549);
or U616 (N_616,In_2117,In_1849);
and U617 (N_617,In_4103,In_4480);
nand U618 (N_618,In_1321,In_3947);
nor U619 (N_619,In_4005,In_1733);
nor U620 (N_620,In_4927,In_4195);
xnor U621 (N_621,In_1379,In_2371);
nand U622 (N_622,In_999,In_2310);
and U623 (N_623,In_1715,In_2916);
nor U624 (N_624,In_419,In_3243);
or U625 (N_625,In_417,In_4555);
or U626 (N_626,In_606,In_2831);
or U627 (N_627,In_3585,In_1608);
nor U628 (N_628,In_4102,In_1025);
and U629 (N_629,In_83,In_2426);
nand U630 (N_630,In_1195,In_4218);
xnor U631 (N_631,In_1125,In_1732);
or U632 (N_632,In_3744,In_4731);
nor U633 (N_633,In_2207,In_3495);
nand U634 (N_634,In_4400,In_1295);
nor U635 (N_635,In_1703,In_1717);
nand U636 (N_636,In_3699,In_1352);
and U637 (N_637,In_1793,In_975);
xnor U638 (N_638,In_3477,In_4);
nand U639 (N_639,In_1016,In_15);
nor U640 (N_640,In_4384,In_4689);
nor U641 (N_641,In_1762,In_3347);
and U642 (N_642,In_1434,In_2826);
or U643 (N_643,In_3147,In_2678);
xor U644 (N_644,In_1441,In_3380);
nor U645 (N_645,In_2522,In_4589);
xnor U646 (N_646,In_3004,In_3874);
xnor U647 (N_647,In_490,In_4650);
xnor U648 (N_648,In_3782,In_4138);
or U649 (N_649,In_1816,In_625);
xor U650 (N_650,In_4326,In_3930);
xnor U651 (N_651,In_3336,In_45);
and U652 (N_652,In_1085,In_590);
or U653 (N_653,In_4266,In_4342);
nor U654 (N_654,In_898,In_4091);
nand U655 (N_655,In_1930,In_3025);
xor U656 (N_656,In_1588,In_1932);
and U657 (N_657,In_395,In_4701);
or U658 (N_658,In_1455,In_2261);
nor U659 (N_659,In_3676,In_3789);
xnor U660 (N_660,In_4396,In_4382);
nor U661 (N_661,In_2313,In_210);
nand U662 (N_662,In_3678,In_1923);
xor U663 (N_663,In_2668,In_991);
or U664 (N_664,In_3296,In_690);
nor U665 (N_665,In_3036,In_366);
and U666 (N_666,In_1232,In_716);
and U667 (N_667,In_1167,In_182);
nand U668 (N_668,In_4251,In_2495);
nor U669 (N_669,In_2350,In_2157);
and U670 (N_670,In_2165,In_2366);
and U671 (N_671,In_1522,In_3849);
or U672 (N_672,In_2162,In_4536);
nand U673 (N_673,In_3966,In_2085);
nor U674 (N_674,In_1280,In_4108);
or U675 (N_675,In_2821,In_3927);
nor U676 (N_676,In_3840,In_3400);
nand U677 (N_677,In_4227,In_2190);
or U678 (N_678,In_2694,In_1378);
and U679 (N_679,In_3535,In_2149);
nor U680 (N_680,In_3899,In_845);
nand U681 (N_681,In_1675,In_161);
xor U682 (N_682,In_449,In_2199);
or U683 (N_683,In_2872,In_1968);
nor U684 (N_684,In_2912,In_2333);
xnor U685 (N_685,In_440,In_1693);
xor U686 (N_686,In_4426,In_3210);
or U687 (N_687,In_4664,In_3029);
nand U688 (N_688,In_739,In_4627);
and U689 (N_689,In_2311,In_2270);
xnor U690 (N_690,In_3940,In_3457);
xnor U691 (N_691,In_3369,In_4313);
and U692 (N_692,In_3579,In_777);
nand U693 (N_693,In_1202,In_1629);
nand U694 (N_694,In_4337,In_2924);
nor U695 (N_695,In_1124,In_3095);
nand U696 (N_696,In_2520,In_312);
nand U697 (N_697,In_541,In_1630);
or U698 (N_698,In_2547,In_2151);
nor U699 (N_699,In_1405,In_3252);
or U700 (N_700,In_1792,In_1178);
and U701 (N_701,In_1820,In_598);
nor U702 (N_702,In_2375,In_4225);
nor U703 (N_703,In_207,In_342);
and U704 (N_704,In_1976,In_3652);
xor U705 (N_705,In_1046,In_3743);
nand U706 (N_706,In_1743,In_2613);
xor U707 (N_707,In_3902,In_2211);
nand U708 (N_708,In_3020,In_887);
nor U709 (N_709,In_578,In_4946);
xnor U710 (N_710,In_2656,In_4358);
xnor U711 (N_711,In_1966,In_3701);
or U712 (N_712,In_1778,In_3992);
xor U713 (N_713,In_2173,In_3912);
or U714 (N_714,In_1004,In_4884);
or U715 (N_715,In_297,In_188);
or U716 (N_716,In_244,In_4405);
nand U717 (N_717,In_270,In_4235);
or U718 (N_718,In_1530,In_3872);
nor U719 (N_719,In_2042,In_1827);
nor U720 (N_720,In_4722,In_3704);
nor U721 (N_721,In_1826,In_2161);
nor U722 (N_722,In_1478,In_318);
or U723 (N_723,In_3783,In_2134);
nand U724 (N_724,In_2948,In_835);
nor U725 (N_725,In_4423,In_2728);
nor U726 (N_726,In_13,In_1363);
nor U727 (N_727,In_2048,In_4821);
nand U728 (N_728,In_2546,In_2327);
nor U729 (N_729,In_715,In_2249);
or U730 (N_730,In_1489,In_3041);
xnor U731 (N_731,In_1344,In_4350);
and U732 (N_732,In_4767,In_2692);
nand U733 (N_733,In_2018,In_2517);
or U734 (N_734,In_783,In_2622);
nor U735 (N_735,In_2618,In_2317);
nand U736 (N_736,In_2435,In_3739);
nand U737 (N_737,In_4799,In_741);
nand U738 (N_738,In_939,In_2603);
or U739 (N_739,In_2745,In_2292);
or U740 (N_740,In_2491,In_1421);
xor U741 (N_741,In_2185,In_763);
nand U742 (N_742,In_3549,In_1587);
nor U743 (N_743,In_4344,In_3830);
nor U744 (N_744,In_4756,In_3575);
and U745 (N_745,In_1795,In_16);
xor U746 (N_746,In_2205,In_2410);
xor U747 (N_747,In_2036,In_468);
xnor U748 (N_748,In_3034,In_4295);
xnor U749 (N_749,In_2938,In_634);
or U750 (N_750,In_3084,In_639);
or U751 (N_751,In_2347,In_3800);
xnor U752 (N_752,In_2178,In_3657);
or U753 (N_753,In_4069,In_1660);
or U754 (N_754,In_668,In_641);
nor U755 (N_755,In_640,In_260);
or U756 (N_756,In_3436,In_2614);
or U757 (N_757,In_2077,In_2661);
xor U758 (N_758,In_3868,In_531);
and U759 (N_759,In_1754,In_957);
and U760 (N_760,In_4835,In_1059);
xnor U761 (N_761,In_3735,In_1311);
nor U762 (N_762,In_4671,In_93);
nand U763 (N_763,In_2455,In_3623);
nor U764 (N_764,In_841,In_1600);
nand U765 (N_765,In_4587,In_3975);
nand U766 (N_766,In_3518,In_1428);
xnor U767 (N_767,In_4298,In_1638);
nor U768 (N_768,In_1117,In_2691);
nor U769 (N_769,In_1531,In_4321);
xor U770 (N_770,In_4690,In_2543);
nor U771 (N_771,In_2787,In_1454);
and U772 (N_772,In_2236,In_3091);
nand U773 (N_773,In_2136,In_3230);
nand U774 (N_774,In_2381,In_3371);
or U775 (N_775,In_2066,In_2918);
xor U776 (N_776,In_3359,In_628);
and U777 (N_777,In_1711,In_2322);
xnor U778 (N_778,In_4508,In_1860);
xor U779 (N_779,In_1912,In_793);
nand U780 (N_780,In_3847,In_4192);
or U781 (N_781,In_3225,In_4850);
or U782 (N_782,In_2803,In_1385);
and U783 (N_783,In_2284,In_3244);
nor U784 (N_784,In_3650,In_849);
xor U785 (N_785,In_4422,In_261);
or U786 (N_786,In_3703,In_1270);
and U787 (N_787,In_4017,In_3155);
or U788 (N_788,In_811,In_4207);
xor U789 (N_789,In_3388,In_1749);
nor U790 (N_790,In_1391,In_3060);
and U791 (N_791,In_4468,In_1985);
nand U792 (N_792,In_1173,In_3205);
and U793 (N_793,In_4889,In_1431);
xor U794 (N_794,In_604,In_4963);
nor U795 (N_795,In_1070,In_704);
and U796 (N_796,In_4054,In_2393);
or U797 (N_797,In_1645,In_2387);
nand U798 (N_798,In_1947,In_1517);
nand U799 (N_799,In_2091,In_2141);
xor U800 (N_800,In_4395,In_4570);
and U801 (N_801,In_3344,In_3646);
nand U802 (N_802,In_4870,In_2062);
or U803 (N_803,In_386,In_3149);
nand U804 (N_804,In_926,In_512);
or U805 (N_805,In_1061,In_2800);
and U806 (N_806,In_1382,In_4277);
xnor U807 (N_807,In_2082,In_3663);
or U808 (N_808,In_3870,In_220);
or U809 (N_809,In_2882,In_2425);
and U810 (N_810,In_2315,In_3855);
and U811 (N_811,In_905,In_2464);
nand U812 (N_812,In_1424,In_4397);
xnor U813 (N_813,In_2321,In_1894);
or U814 (N_814,In_3000,In_4748);
xor U815 (N_815,In_1594,In_3641);
and U816 (N_816,In_1685,In_4716);
and U817 (N_817,In_3068,In_4411);
nor U818 (N_818,In_577,In_2331);
xnor U819 (N_819,In_784,In_360);
nor U820 (N_820,In_642,In_2263);
and U821 (N_821,In_4052,In_2660);
and U822 (N_822,In_4907,In_4087);
nor U823 (N_823,In_4383,In_1043);
xor U824 (N_824,In_3350,In_326);
xnor U825 (N_825,In_2698,In_4188);
xnor U826 (N_826,In_662,In_4786);
or U827 (N_827,In_1978,In_2707);
nand U828 (N_828,In_3353,In_294);
and U829 (N_829,In_1726,In_4370);
nand U830 (N_830,In_4525,In_1140);
nor U831 (N_831,In_564,In_3064);
and U832 (N_832,In_3746,In_1155);
xor U833 (N_833,In_1714,In_4672);
nor U834 (N_834,In_1464,In_3584);
nor U835 (N_835,In_3937,In_4028);
nor U836 (N_836,In_3292,In_1993);
and U837 (N_837,In_1705,In_3159);
xor U838 (N_838,In_2769,In_1048);
or U839 (N_839,In_3749,In_4899);
nor U840 (N_840,In_2749,In_1472);
xor U841 (N_841,In_730,In_1398);
nor U842 (N_842,In_4544,In_3680);
nand U843 (N_843,In_296,In_1460);
xor U844 (N_844,In_3014,In_2408);
or U845 (N_845,In_3688,In_4564);
and U846 (N_846,In_1959,In_3563);
or U847 (N_847,In_3464,In_2581);
or U848 (N_848,In_2403,In_2598);
nand U849 (N_849,In_5,In_4958);
xnor U850 (N_850,In_3901,In_4424);
nor U851 (N_851,In_4491,In_2039);
or U852 (N_852,In_3042,In_3825);
xor U853 (N_853,In_4817,In_938);
nor U854 (N_854,In_861,In_302);
nand U855 (N_855,In_2301,In_2696);
xor U856 (N_856,In_4802,In_3162);
nand U857 (N_857,In_4186,In_3634);
nand U858 (N_858,In_2824,In_4909);
nor U859 (N_859,In_2197,In_166);
xor U860 (N_860,In_3309,In_4318);
and U861 (N_861,In_2037,In_2740);
or U862 (N_862,In_1207,In_314);
nand U863 (N_863,In_2693,In_1957);
or U864 (N_864,In_2259,In_2852);
or U865 (N_865,In_3471,In_2154);
or U866 (N_866,In_1960,In_2296);
xor U867 (N_867,In_1000,In_2519);
nand U868 (N_868,In_3012,In_2169);
xnor U869 (N_869,In_1746,In_1684);
xor U870 (N_870,In_159,In_3082);
xnor U871 (N_871,In_927,In_1034);
nand U872 (N_872,In_824,In_4463);
nand U873 (N_873,In_955,In_1590);
nand U874 (N_874,In_344,In_1636);
xnor U875 (N_875,In_2015,In_1641);
xor U876 (N_876,In_316,In_3107);
nand U877 (N_877,In_937,In_3171);
or U878 (N_878,In_1558,In_4554);
or U879 (N_879,In_3734,In_4530);
or U880 (N_880,In_2642,In_155);
or U881 (N_881,In_2760,In_3624);
nor U882 (N_882,In_3215,In_631);
nand U883 (N_883,In_4922,In_3080);
nand U884 (N_884,In_242,In_2731);
or U885 (N_885,In_1949,In_1426);
nor U886 (N_886,In_492,In_893);
xnor U887 (N_887,In_1296,In_30);
xor U888 (N_888,In_2690,In_4659);
or U889 (N_889,In_1157,In_3616);
or U890 (N_890,In_4694,In_1278);
or U891 (N_891,In_2129,In_638);
xor U892 (N_892,In_1928,In_1821);
nor U893 (N_893,In_768,In_4803);
xnor U894 (N_894,In_4565,In_1940);
and U895 (N_895,In_4541,In_4567);
or U896 (N_896,In_2929,In_4794);
nand U897 (N_897,In_2059,In_2416);
nand U898 (N_898,In_313,In_2574);
or U899 (N_899,In_3152,In_2121);
nor U900 (N_900,In_717,In_2021);
or U901 (N_901,In_2323,In_3);
xnor U902 (N_902,In_2104,In_1154);
or U903 (N_903,In_3952,In_4476);
nor U904 (N_904,In_1269,In_1965);
xnor U905 (N_905,In_3821,In_1306);
and U906 (N_906,In_2865,In_1390);
or U907 (N_907,In_1990,In_3209);
nand U908 (N_908,In_1605,In_4988);
or U909 (N_909,In_3484,In_1845);
and U910 (N_910,In_1392,In_1294);
or U911 (N_911,In_1247,In_4903);
nand U912 (N_912,In_1053,In_3030);
or U913 (N_913,In_4742,In_4335);
and U914 (N_914,In_4042,In_4242);
xor U915 (N_915,In_3108,In_4921);
nor U916 (N_916,In_734,In_480);
and U917 (N_917,In_2801,In_3674);
nor U918 (N_918,In_345,In_2914);
xor U919 (N_919,In_198,In_2703);
nand U920 (N_920,In_1853,In_2875);
xor U921 (N_921,In_623,In_2058);
or U922 (N_922,In_803,In_4804);
nor U923 (N_923,In_3196,In_627);
xnor U924 (N_924,In_4785,In_2889);
or U925 (N_925,In_2232,In_4965);
and U926 (N_926,In_871,In_745);
xnor U927 (N_927,In_2043,In_3426);
nor U928 (N_928,In_2489,In_4796);
xnor U929 (N_929,In_3963,In_1143);
xor U930 (N_930,In_2432,In_2187);
or U931 (N_931,In_4245,In_1277);
and U932 (N_932,In_358,In_4386);
xor U933 (N_933,In_1076,In_2585);
and U934 (N_934,In_189,In_4270);
xnor U935 (N_935,In_4471,In_3954);
nor U936 (N_936,In_2345,In_920);
and U937 (N_937,In_4591,In_23);
nor U938 (N_938,In_2981,In_4189);
nor U939 (N_939,In_143,In_1627);
nand U940 (N_940,In_64,In_491);
and U941 (N_941,In_977,In_251);
nor U942 (N_942,In_4580,In_3069);
and U943 (N_943,In_4450,In_2031);
nor U944 (N_944,In_473,In_3085);
nand U945 (N_945,In_2505,In_1712);
nor U946 (N_946,In_2978,In_3883);
nor U947 (N_947,In_1364,In_3473);
nor U948 (N_948,In_1406,In_3142);
nor U949 (N_949,In_3356,In_2213);
nand U950 (N_950,In_1179,In_4704);
nor U951 (N_951,In_4708,In_228);
xnor U952 (N_952,In_4031,In_534);
xor U953 (N_953,In_3024,In_4443);
nand U954 (N_954,In_49,In_1788);
or U955 (N_955,In_2417,In_4808);
xor U956 (N_956,In_3911,In_3378);
xor U957 (N_957,In_3338,In_3189);
and U958 (N_958,In_3040,In_4257);
xnor U959 (N_959,In_1766,In_26);
xnor U960 (N_960,In_1983,In_1151);
nor U961 (N_961,In_1265,In_2756);
nor U962 (N_962,In_2820,In_416);
and U963 (N_963,In_1952,In_3490);
xor U964 (N_964,In_620,In_255);
and U965 (N_965,In_1654,In_2475);
xor U966 (N_966,In_423,In_1503);
nand U967 (N_967,In_954,In_582);
xor U968 (N_968,In_4454,In_1842);
nor U969 (N_969,In_4436,In_3950);
and U970 (N_970,In_4718,In_767);
and U971 (N_971,In_3032,In_1138);
xnor U972 (N_972,In_4970,In_4954);
nand U973 (N_973,In_2624,In_862);
and U974 (N_974,In_1759,In_3718);
or U975 (N_975,In_4652,In_765);
xnor U976 (N_976,In_3804,In_3067);
and U977 (N_977,In_3027,In_4262);
nand U978 (N_978,In_290,In_3878);
xor U979 (N_979,In_1299,In_22);
and U980 (N_980,In_85,In_2884);
nand U981 (N_981,In_621,In_1847);
and U982 (N_982,In_1539,In_1716);
and U983 (N_983,In_1190,In_1551);
nor U984 (N_984,In_2936,In_29);
or U985 (N_985,In_104,In_4171);
xnor U986 (N_986,In_4303,In_4566);
and U987 (N_987,In_538,In_4271);
nand U988 (N_988,In_2238,In_3537);
and U989 (N_989,In_1239,In_3126);
nand U990 (N_990,In_1238,In_802);
or U991 (N_991,In_3611,In_3926);
nand U992 (N_992,In_3807,In_4679);
xnor U993 (N_993,In_1284,In_3764);
xor U994 (N_994,In_3269,In_3211);
or U995 (N_995,In_1527,In_673);
nor U996 (N_996,In_4750,In_1565);
nand U997 (N_997,In_2492,In_3987);
xnor U998 (N_998,In_822,In_2984);
xnor U999 (N_999,In_4622,In_2441);
nor U1000 (N_1000,In_3236,In_2548);
nor U1001 (N_1001,In_3884,In_1840);
nand U1002 (N_1002,In_1939,In_1374);
nand U1003 (N_1003,In_2167,In_814);
nand U1004 (N_1004,In_794,In_3932);
and U1005 (N_1005,In_3140,In_2078);
nand U1006 (N_1006,In_2103,In_2578);
xor U1007 (N_1007,In_4864,In_773);
or U1008 (N_1008,In_4234,In_725);
nand U1009 (N_1009,In_1292,In_158);
nand U1010 (N_1010,In_3087,In_193);
nand U1011 (N_1011,In_758,In_786);
xor U1012 (N_1012,In_4493,In_106);
xor U1013 (N_1013,In_224,In_4938);
xor U1014 (N_1014,In_2722,In_3787);
nand U1015 (N_1015,In_2320,In_4163);
and U1016 (N_1016,In_46,In_1700);
nor U1017 (N_1017,In_3061,In_1614);
or U1018 (N_1018,In_3151,In_2235);
xnor U1019 (N_1019,In_3959,In_4680);
xor U1020 (N_1020,In_2060,In_2945);
nand U1021 (N_1021,In_4883,In_4798);
nor U1022 (N_1022,In_3348,In_194);
xor U1023 (N_1023,In_605,In_771);
and U1024 (N_1024,In_3828,In_3175);
xor U1025 (N_1025,In_1308,In_1801);
xnor U1026 (N_1026,In_2880,In_806);
and U1027 (N_1027,In_2718,In_703);
nand U1028 (N_1028,In_3747,In_3192);
nor U1029 (N_1029,In_4352,In_2014);
nor U1030 (N_1030,In_4060,In_1728);
or U1031 (N_1031,In_1009,In_3515);
nor U1032 (N_1032,In_2841,In_2634);
xor U1033 (N_1033,In_4467,In_4758);
or U1034 (N_1034,In_396,In_2724);
nand U1035 (N_1035,In_4577,In_4197);
nor U1036 (N_1036,In_3125,In_1602);
nor U1037 (N_1037,In_2451,In_4485);
and U1038 (N_1038,In_2100,In_4228);
nand U1039 (N_1039,In_3488,In_3581);
and U1040 (N_1040,In_3349,In_317);
nor U1041 (N_1041,In_2930,In_1880);
xnor U1042 (N_1042,In_3062,In_3178);
nand U1043 (N_1043,In_4088,In_1856);
or U1044 (N_1044,In_2518,In_129);
and U1045 (N_1045,In_4610,In_1201);
nand U1046 (N_1046,In_2471,In_3049);
xor U1047 (N_1047,In_4248,In_2558);
or U1048 (N_1048,In_3303,In_3564);
and U1049 (N_1049,In_4879,In_3601);
and U1050 (N_1050,In_2781,In_3740);
nor U1051 (N_1051,In_4574,In_2002);
or U1052 (N_1052,In_3460,In_1158);
nor U1053 (N_1053,In_427,In_643);
or U1054 (N_1054,In_1972,In_1653);
xor U1055 (N_1055,In_2521,In_575);
and U1056 (N_1056,In_2599,In_4239);
xor U1057 (N_1057,In_3078,In_859);
nand U1058 (N_1058,In_3978,In_4428);
or U1059 (N_1059,In_4160,In_4336);
or U1060 (N_1060,In_499,In_54);
xor U1061 (N_1061,In_359,In_3670);
nor U1062 (N_1062,In_1781,In_4098);
nor U1063 (N_1063,In_2761,In_3288);
or U1064 (N_1064,In_3781,In_2254);
or U1065 (N_1065,In_3193,In_4868);
nand U1066 (N_1066,In_4830,In_1327);
or U1067 (N_1067,In_2962,In_4772);
xnor U1068 (N_1068,In_4971,In_436);
and U1069 (N_1069,In_1370,In_338);
xnor U1070 (N_1070,In_1137,In_2390);
nand U1071 (N_1071,In_2302,In_485);
and U1072 (N_1072,In_233,In_1680);
and U1073 (N_1073,In_1425,In_2977);
nor U1074 (N_1074,In_481,In_856);
and U1075 (N_1075,In_4285,In_82);
nand U1076 (N_1076,In_1557,In_834);
xor U1077 (N_1077,In_4500,In_4588);
or U1078 (N_1078,In_1891,In_3779);
xnor U1079 (N_1079,In_1348,In_4247);
and U1080 (N_1080,In_2089,In_362);
xnor U1081 (N_1081,In_1852,In_2290);
or U1082 (N_1082,In_2551,In_2216);
xor U1083 (N_1083,In_2965,In_2340);
and U1084 (N_1084,In_2988,In_1943);
nand U1085 (N_1085,In_2130,In_3379);
and U1086 (N_1086,In_4823,In_864);
nand U1087 (N_1087,In_3217,In_3768);
and U1088 (N_1088,In_4217,In_3811);
or U1089 (N_1089,In_3239,In_1017);
or U1090 (N_1090,In_689,In_2643);
nand U1091 (N_1091,In_3949,In_1647);
nand U1092 (N_1092,In_3767,In_2188);
xnor U1093 (N_1093,In_4208,In_987);
xor U1094 (N_1094,In_2496,In_2140);
xor U1095 (N_1095,In_394,In_1241);
or U1096 (N_1096,In_1254,In_2357);
and U1097 (N_1097,In_3999,In_560);
nand U1098 (N_1098,In_1649,In_2524);
and U1099 (N_1099,In_2786,In_2438);
xnor U1100 (N_1100,In_4881,In_2917);
xor U1101 (N_1101,In_1951,In_1970);
xor U1102 (N_1102,In_3972,In_4181);
nor U1103 (N_1103,In_2963,In_4001);
nand U1104 (N_1104,In_2113,In_677);
and U1105 (N_1105,In_3599,In_1785);
or U1106 (N_1106,In_4640,In_2181);
xor U1107 (N_1107,In_3910,In_3574);
nand U1108 (N_1108,In_2919,In_524);
or U1109 (N_1109,In_4896,In_3098);
xor U1110 (N_1110,In_2112,In_122);
nor U1111 (N_1111,In_2291,In_1825);
and U1112 (N_1112,In_2685,In_1794);
or U1113 (N_1113,In_1569,In_2110);
xor U1114 (N_1114,In_3093,In_4147);
or U1115 (N_1115,In_2020,In_3757);
xor U1116 (N_1116,In_956,In_2616);
nor U1117 (N_1117,In_2329,In_3971);
xnor U1118 (N_1118,In_2910,In_389);
or U1119 (N_1119,In_670,In_2531);
xor U1120 (N_1120,In_853,In_1341);
nand U1121 (N_1121,In_4914,In_482);
and U1122 (N_1122,In_4774,In_3145);
nor U1123 (N_1123,In_1896,In_3226);
or U1124 (N_1124,In_825,In_3968);
and U1125 (N_1125,In_2825,In_4300);
nand U1126 (N_1126,In_4446,In_4600);
nand U1127 (N_1127,In_4075,In_2592);
nor U1128 (N_1128,In_3797,In_2108);
nand U1129 (N_1129,In_257,In_3128);
nor U1130 (N_1130,In_4832,In_4081);
and U1131 (N_1131,In_2247,In_842);
nand U1132 (N_1132,In_320,In_4552);
or U1133 (N_1133,In_3724,In_762);
or U1134 (N_1134,In_4434,In_4159);
and U1135 (N_1135,In_150,In_2120);
xor U1136 (N_1136,In_2991,In_2877);
xnor U1137 (N_1137,In_2755,In_2753);
and U1138 (N_1138,In_1767,In_3110);
and U1139 (N_1139,In_4178,In_699);
nand U1140 (N_1140,In_442,In_2636);
or U1141 (N_1141,In_4791,In_4730);
nor U1142 (N_1142,In_3557,In_1);
nand U1143 (N_1143,In_2186,In_612);
and U1144 (N_1144,In_4026,In_2465);
nor U1145 (N_1145,In_107,In_600);
xor U1146 (N_1146,In_370,In_4267);
nand U1147 (N_1147,In_989,In_3311);
nand U1148 (N_1148,In_944,In_747);
and U1149 (N_1149,In_1194,In_4871);
or U1150 (N_1150,In_1895,In_4109);
nor U1151 (N_1151,In_81,In_2107);
and U1152 (N_1152,In_1376,In_2629);
nand U1153 (N_1153,In_4149,In_1787);
nand U1154 (N_1154,In_993,In_2710);
nor U1155 (N_1155,In_732,In_1538);
or U1156 (N_1156,In_4593,In_4806);
and U1157 (N_1157,In_2506,In_750);
xnor U1158 (N_1158,In_4643,In_1637);
nand U1159 (N_1159,In_848,In_4146);
and U1160 (N_1160,In_3047,In_2888);
nor U1161 (N_1161,In_1397,In_1362);
nor U1162 (N_1162,In_2780,In_4209);
or U1163 (N_1163,In_4801,In_2662);
nor U1164 (N_1164,In_3174,In_828);
and U1165 (N_1165,In_1704,In_4216);
nand U1166 (N_1166,In_552,In_2057);
or U1167 (N_1167,In_4448,In_1474);
xnor U1168 (N_1168,In_4518,In_108);
nor U1169 (N_1169,In_705,In_3399);
and U1170 (N_1170,In_611,In_1372);
xnor U1171 (N_1171,In_474,In_4511);
nor U1172 (N_1172,In_3397,In_2985);
nand U1173 (N_1173,In_1907,In_4018);
or U1174 (N_1174,In_2793,In_2545);
or U1175 (N_1175,In_3567,In_2604);
or U1176 (N_1176,In_4825,In_4144);
nand U1177 (N_1177,In_752,In_4952);
xnor U1178 (N_1178,In_2783,In_4619);
nor U1179 (N_1179,In_4829,In_2215);
or U1180 (N_1180,In_4465,In_594);
nor U1181 (N_1181,In_3016,In_3907);
nand U1182 (N_1182,In_1013,In_3760);
and U1183 (N_1183,In_176,In_1674);
xor U1184 (N_1184,In_4513,In_819);
nand U1185 (N_1185,In_4329,In_2377);
or U1186 (N_1186,In_3203,In_1166);
nor U1187 (N_1187,In_3592,In_4299);
nor U1188 (N_1188,In_2990,In_4083);
and U1189 (N_1189,In_2814,In_4741);
and U1190 (N_1190,In_1130,In_2915);
nor U1191 (N_1191,In_4646,In_4721);
xnor U1192 (N_1192,In_475,In_2137);
nor U1193 (N_1193,In_3274,In_3172);
nand U1194 (N_1194,In_723,In_4678);
nor U1195 (N_1195,In_4179,In_2816);
xnor U1196 (N_1196,In_3102,In_1084);
or U1197 (N_1197,In_3482,In_3018);
nor U1198 (N_1198,In_2219,In_1221);
or U1199 (N_1199,In_1997,In_1924);
xor U1200 (N_1200,In_3295,In_1506);
or U1201 (N_1201,In_757,In_3649);
or U1202 (N_1202,In_4029,In_3524);
nor U1203 (N_1203,In_674,In_3333);
and U1204 (N_1204,In_2510,In_3660);
and U1205 (N_1205,In_2845,In_1595);
nor U1206 (N_1206,In_4291,In_199);
and U1207 (N_1207,In_2504,In_2952);
nand U1208 (N_1208,In_2730,In_2208);
xnor U1209 (N_1209,In_1748,In_2257);
nand U1210 (N_1210,In_3513,In_2659);
nand U1211 (N_1211,In_1763,In_740);
and U1212 (N_1212,In_337,In_2600);
or U1213 (N_1213,In_99,In_1784);
nand U1214 (N_1214,In_4236,In_3302);
or U1215 (N_1215,In_157,In_4212);
nor U1216 (N_1216,In_2045,In_278);
nand U1217 (N_1217,In_3485,In_2354);
or U1218 (N_1218,In_4878,In_1946);
xor U1219 (N_1219,In_820,In_4037);
and U1220 (N_1220,In_2262,In_2971);
and U1221 (N_1221,In_4904,In_218);
nor U1222 (N_1222,In_4783,In_855);
nor U1223 (N_1223,In_4675,In_3914);
nand U1224 (N_1224,In_4170,In_469);
nor U1225 (N_1225,In_232,In_41);
xnor U1226 (N_1226,In_4873,In_1621);
nand U1227 (N_1227,In_4557,In_487);
xnor U1228 (N_1228,In_527,In_7);
nand U1229 (N_1229,In_1435,In_4880);
or U1230 (N_1230,In_2035,In_4076);
xnor U1231 (N_1231,In_1883,In_2473);
nand U1232 (N_1232,In_557,In_2353);
nand U1233 (N_1233,In_972,In_3871);
and U1234 (N_1234,In_881,In_4860);
or U1235 (N_1235,In_3262,In_2231);
nand U1236 (N_1236,In_1366,In_4151);
nor U1237 (N_1237,In_1210,In_3862);
and U1238 (N_1238,In_2380,In_2568);
xor U1239 (N_1239,In_2268,In_971);
and U1240 (N_1240,In_680,In_593);
nand U1241 (N_1241,In_4523,In_4560);
and U1242 (N_1242,In_4206,In_4437);
or U1243 (N_1243,In_711,In_3887);
and U1244 (N_1244,In_3445,In_3326);
nand U1245 (N_1245,In_3063,In_3539);
nor U1246 (N_1246,In_460,In_3586);
and U1247 (N_1247,In_279,In_2001);
nor U1248 (N_1248,In_2790,In_2808);
and U1249 (N_1249,In_2960,In_3136);
or U1250 (N_1250,In_4099,In_205);
nor U1251 (N_1251,In_1504,In_3958);
nand U1252 (N_1252,In_1702,In_4104);
and U1253 (N_1253,In_3831,In_2339);
or U1254 (N_1254,In_4238,In_3898);
nor U1255 (N_1255,In_172,In_3360);
xor U1256 (N_1256,In_1253,In_3961);
xor U1257 (N_1257,In_1477,In_4173);
nor U1258 (N_1258,In_2644,In_4974);
nand U1259 (N_1259,In_3437,In_2179);
and U1260 (N_1260,In_2000,In_330);
nor U1261 (N_1261,In_4067,In_548);
nor U1262 (N_1262,In_2148,In_3796);
or U1263 (N_1263,In_3568,In_2044);
and U1264 (N_1264,In_2474,In_4093);
and U1265 (N_1265,In_4935,In_2277);
nand U1266 (N_1266,In_1442,In_2941);
or U1267 (N_1267,In_171,In_1926);
nand U1268 (N_1268,In_583,In_844);
nand U1269 (N_1269,In_1160,In_4682);
nand U1270 (N_1270,In_1407,In_2719);
nand U1271 (N_1271,In_996,In_1519);
xnor U1272 (N_1272,In_3105,In_3846);
and U1273 (N_1273,In_4325,In_863);
nor U1274 (N_1274,In_801,In_2419);
and U1275 (N_1275,In_4706,In_3300);
and U1276 (N_1276,In_990,In_4842);
xnor U1277 (N_1277,In_983,In_1212);
and U1278 (N_1278,In_4684,In_4053);
nor U1279 (N_1279,In_2605,In_3517);
xnor U1280 (N_1280,In_2256,In_3707);
nor U1281 (N_1281,In_1273,In_3613);
nand U1282 (N_1282,In_4781,In_4015);
nor U1283 (N_1283,In_3055,In_3653);
nand U1284 (N_1284,In_4726,In_2777);
xor U1285 (N_1285,In_1507,In_2477);
nor U1286 (N_1286,In_787,In_2940);
nor U1287 (N_1287,In_2449,In_3462);
and U1288 (N_1288,In_3219,In_3157);
and U1289 (N_1289,In_4942,In_4510);
xor U1290 (N_1290,In_1740,In_4077);
nand U1291 (N_1291,In_478,In_1879);
and U1292 (N_1292,In_733,In_4260);
xor U1293 (N_1293,In_461,In_1671);
or U1294 (N_1294,In_4022,In_4156);
and U1295 (N_1295,In_1260,In_3208);
nor U1296 (N_1296,In_3222,In_3419);
nor U1297 (N_1297,In_850,In_875);
nor U1298 (N_1298,In_3501,In_3981);
xor U1299 (N_1299,In_1420,In_4691);
nand U1300 (N_1300,In_2922,In_2529);
and U1301 (N_1301,In_3525,In_1331);
nand U1302 (N_1302,In_521,In_3377);
nand U1303 (N_1303,In_3119,In_4780);
and U1304 (N_1304,In_1817,In_4931);
nor U1305 (N_1305,In_3681,In_3362);
and U1306 (N_1306,In_3499,In_904);
nand U1307 (N_1307,In_3086,In_500);
or U1308 (N_1308,In_4306,In_443);
or U1309 (N_1309,In_3771,In_4258);
and U1310 (N_1310,In_2493,In_2017);
xnor U1311 (N_1311,In_949,In_2858);
and U1312 (N_1312,In_4073,In_501);
nand U1313 (N_1313,In_3943,In_2561);
or U1314 (N_1314,In_2630,In_3594);
and U1315 (N_1315,In_1417,In_3421);
or U1316 (N_1316,In_1030,In_624);
or U1317 (N_1317,In_4596,In_3555);
and U1318 (N_1318,In_1289,In_347);
and U1319 (N_1319,In_2674,In_4858);
and U1320 (N_1320,In_1419,In_2457);
nor U1321 (N_1321,In_277,In_607);
or U1322 (N_1322,In_3997,In_3903);
nand U1323 (N_1323,In_2503,In_3150);
and U1324 (N_1324,In_3684,In_2196);
and U1325 (N_1325,In_2172,In_2705);
nor U1326 (N_1326,In_184,In_2958);
nor U1327 (N_1327,In_3531,In_2588);
or U1328 (N_1328,In_4793,In_1104);
nand U1329 (N_1329,In_2398,In_2807);
xor U1330 (N_1330,In_2863,In_1343);
nand U1331 (N_1331,In_916,In_1068);
nand U1332 (N_1332,In_701,In_4074);
xor U1333 (N_1333,In_2648,In_4532);
xnor U1334 (N_1334,In_3407,In_3213);
xnor U1335 (N_1335,In_1988,In_1156);
and U1336 (N_1336,In_4364,In_4642);
and U1337 (N_1337,In_127,In_3316);
nand U1338 (N_1338,In_2641,In_1467);
and U1339 (N_1339,In_1659,In_20);
nor U1340 (N_1340,In_92,In_3168);
xnor U1341 (N_1341,In_1144,In_4978);
and U1342 (N_1342,In_3838,In_4464);
xor U1343 (N_1343,In_4853,In_3424);
or U1344 (N_1344,In_4394,In_1836);
or U1345 (N_1345,In_3334,In_2374);
nor U1346 (N_1346,In_1213,In_4666);
xor U1347 (N_1347,In_3604,In_3973);
and U1348 (N_1348,In_3304,In_3478);
nor U1349 (N_1349,In_3186,In_4490);
and U1350 (N_1350,In_4413,In_1305);
nand U1351 (N_1351,In_4086,In_3686);
xnor U1352 (N_1352,In_2144,In_1098);
and U1353 (N_1353,In_3785,In_2358);
nor U1354 (N_1354,In_3458,In_4065);
xnor U1355 (N_1355,In_3860,In_3116);
and U1356 (N_1356,In_4573,In_1935);
or U1357 (N_1357,In_2307,In_4599);
or U1358 (N_1358,In_688,In_1950);
or U1359 (N_1359,In_2061,In_3299);
or U1360 (N_1360,In_1150,In_919);
nand U1361 (N_1361,In_672,In_1508);
xnor U1362 (N_1362,In_4790,In_4107);
xor U1363 (N_1363,In_2856,In_2539);
nand U1364 (N_1364,In_3298,In_3275);
and U1365 (N_1365,In_3153,In_2849);
nand U1366 (N_1366,In_2687,In_3070);
nand U1367 (N_1367,In_1686,In_753);
nand U1368 (N_1368,In_1648,In_1215);
xor U1369 (N_1369,In_2743,In_4062);
xor U1370 (N_1370,In_4734,In_90);
nor U1371 (N_1371,In_292,In_889);
nand U1372 (N_1372,In_4165,In_2281);
nor U1373 (N_1373,In_2873,In_4543);
xnor U1374 (N_1374,In_3541,In_976);
or U1375 (N_1375,In_3556,In_661);
nor U1376 (N_1376,In_295,In_2332);
and U1377 (N_1377,In_1710,In_197);
xnor U1378 (N_1378,In_4519,In_1074);
nor U1379 (N_1379,In_2798,In_4915);
and U1380 (N_1380,In_1818,In_3138);
nor U1381 (N_1381,In_982,In_3934);
nand U1382 (N_1382,In_3806,In_609);
or U1383 (N_1383,In_2767,In_1872);
nor U1384 (N_1384,In_4707,In_1165);
nand U1385 (N_1385,In_4150,In_1383);
and U1386 (N_1386,In_178,In_3184);
nand U1387 (N_1387,In_3526,In_3494);
xor U1388 (N_1388,In_2158,In_4213);
or U1389 (N_1389,In_2182,In_4673);
or U1390 (N_1390,In_4501,In_2812);
xnor U1391 (N_1391,In_3931,In_1220);
or U1392 (N_1392,In_4509,In_1303);
or U1393 (N_1393,In_4755,In_2992);
nand U1394 (N_1394,In_479,In_2047);
or U1395 (N_1395,In_556,In_1901);
nor U1396 (N_1396,In_35,In_2593);
nand U1397 (N_1397,In_3765,In_309);
or U1398 (N_1398,In_879,In_4180);
nand U1399 (N_1399,In_1963,In_4705);
and U1400 (N_1400,In_4182,In_4096);
nand U1401 (N_1401,In_3516,In_47);
nand U1402 (N_1402,In_3877,In_3559);
and U1403 (N_1403,In_870,In_3709);
or U1404 (N_1404,In_4854,In_1720);
nand U1405 (N_1405,In_1283,In_3543);
or U1406 (N_1406,In_1242,In_3121);
nand U1407 (N_1407,In_4990,In_4820);
nor U1408 (N_1408,In_1721,In_3212);
nor U1409 (N_1409,In_3202,In_2177);
nand U1410 (N_1410,In_2612,In_2217);
or U1411 (N_1411,In_839,In_678);
nor U1412 (N_1412,In_2949,In_2423);
nand U1413 (N_1413,In_4185,In_1330);
and U1414 (N_1414,In_4773,In_3364);
nor U1415 (N_1415,In_3996,In_411);
and U1416 (N_1416,In_2868,In_3815);
xor U1417 (N_1417,In_868,In_805);
or U1418 (N_1418,In_1040,In_3571);
nand U1419 (N_1419,In_4283,In_31);
or U1420 (N_1420,In_4316,In_3529);
nor U1421 (N_1421,In_1439,In_2712);
xor U1422 (N_1422,In_3576,In_4631);
nor U1423 (N_1423,In_458,In_298);
and U1424 (N_1424,In_4359,In_2083);
or U1425 (N_1425,In_4986,In_516);
and U1426 (N_1426,In_375,In_4787);
xor U1427 (N_1427,In_3848,In_1176);
nor U1428 (N_1428,In_902,In_2758);
xor U1429 (N_1429,In_2998,In_1616);
nor U1430 (N_1430,In_4551,In_2732);
and U1431 (N_1431,In_3864,In_1991);
xnor U1432 (N_1432,In_315,In_2396);
nor U1433 (N_1433,In_1770,In_306);
xor U1434 (N_1434,In_657,In_269);
xnor U1435 (N_1435,In_917,In_2434);
nor U1436 (N_1436,In_1429,In_4603);
nand U1437 (N_1437,In_3803,In_3583);
nor U1438 (N_1438,In_1927,In_2241);
or U1439 (N_1439,In_4214,In_2049);
xnor U1440 (N_1440,In_149,In_4304);
or U1441 (N_1441,In_958,In_1443);
nand U1442 (N_1442,In_2024,In_1542);
or U1443 (N_1443,In_2202,In_2088);
and U1444 (N_1444,In_1095,In_2542);
nand U1445 (N_1445,In_1466,In_2253);
or U1446 (N_1446,In_4444,In_1861);
and U1447 (N_1447,In_843,In_676);
nor U1448 (N_1448,In_365,In_4264);
and U1449 (N_1449,In_858,In_80);
and U1450 (N_1450,In_555,In_3790);
and U1451 (N_1451,In_892,In_457);
nor U1452 (N_1452,In_1815,In_517);
xor U1453 (N_1453,In_3015,In_1632);
nor U1454 (N_1454,In_2119,In_3111);
nand U1455 (N_1455,In_3960,In_2955);
nor U1456 (N_1456,In_3220,In_4647);
nor U1457 (N_1457,In_1356,In_1851);
xor U1458 (N_1458,In_2586,In_4360);
nand U1459 (N_1459,In_2666,In_3081);
nor U1460 (N_1460,In_2528,In_9);
or U1461 (N_1461,In_1533,In_4243);
or U1462 (N_1462,In_4292,In_415);
nor U1463 (N_1463,In_4749,In_177);
or U1464 (N_1464,In_1170,In_1709);
nor U1465 (N_1465,In_4381,In_2552);
nor U1466 (N_1466,In_731,In_766);
nand U1467 (N_1467,In_3814,In_3698);
nand U1468 (N_1468,In_4484,In_1688);
or U1469 (N_1469,In_3308,In_2394);
nor U1470 (N_1470,In_2822,In_3540);
nor U1471 (N_1471,In_997,In_4161);
xnor U1472 (N_1472,In_3383,In_3272);
and U1473 (N_1473,In_4681,In_2839);
and U1474 (N_1474,In_928,In_1755);
xor U1475 (N_1475,In_2143,In_1984);
xor U1476 (N_1476,In_4516,In_2763);
and U1477 (N_1477,In_1941,In_3335);
xnor U1478 (N_1478,In_1233,In_3916);
or U1479 (N_1479,In_2486,In_1734);
and U1480 (N_1480,In_948,In_414);
nand U1481 (N_1481,In_3206,In_202);
nand U1482 (N_1482,In_507,In_840);
or U1483 (N_1483,In_2997,In_3139);
or U1484 (N_1484,In_2298,In_1889);
or U1485 (N_1485,In_4487,In_3443);
or U1486 (N_1486,In_854,In_1667);
nor U1487 (N_1487,In_536,In_1885);
and U1488 (N_1488,In_3048,In_3900);
nand U1489 (N_1489,In_1698,In_3644);
nor U1490 (N_1490,In_1844,In_4933);
nand U1491 (N_1491,In_3881,In_447);
nand U1492 (N_1492,In_1353,In_1340);
or U1493 (N_1493,In_2657,In_4176);
or U1494 (N_1494,In_1514,In_1258);
nor U1495 (N_1495,In_821,In_1724);
and U1496 (N_1496,In_361,In_4409);
nand U1497 (N_1497,In_4882,In_2894);
or U1498 (N_1498,In_2966,In_1834);
or U1499 (N_1499,In_963,In_4992);
or U1500 (N_1500,In_34,In_3647);
nor U1501 (N_1501,In_4259,In_4934);
nor U1502 (N_1502,In_830,In_223);
nor U1503 (N_1503,In_3630,In_254);
xor U1504 (N_1504,In_4628,In_431);
nand U1505 (N_1505,In_4016,In_2670);
and U1506 (N_1506,In_2715,In_262);
nand U1507 (N_1507,In_3083,In_4960);
or U1508 (N_1508,In_448,In_1809);
xnor U1509 (N_1509,In_2700,In_3439);
or U1510 (N_1510,In_1300,In_229);
and U1511 (N_1511,In_1058,In_4863);
xor U1512 (N_1512,In_71,In_4237);
or U1513 (N_1513,In_4620,In_3809);
and U1514 (N_1514,In_3467,In_2682);
nand U1515 (N_1515,In_3278,In_494);
xnor U1516 (N_1516,In_3013,In_3385);
and U1517 (N_1517,In_4230,In_1982);
or U1518 (N_1518,In_4760,In_4943);
or U1519 (N_1519,In_736,In_4686);
or U1520 (N_1520,In_1133,In_2846);
nand U1521 (N_1521,In_1275,In_1459);
and U1522 (N_1522,In_3590,In_2766);
nor U1523 (N_1523,In_3587,In_6);
or U1524 (N_1524,In_4371,In_2269);
and U1525 (N_1525,In_2887,In_2970);
nand U1526 (N_1526,In_2389,In_817);
xnor U1527 (N_1527,In_1313,In_3320);
xor U1528 (N_1528,In_2501,In_3521);
or U1529 (N_1529,In_1006,In_2400);
or U1530 (N_1530,In_4597,In_3372);
nand U1531 (N_1531,In_4066,In_1288);
xor U1532 (N_1532,In_1523,In_463);
nand U1533 (N_1533,In_2560,In_1359);
nand U1534 (N_1534,In_2921,In_1413);
xor U1535 (N_1535,In_1128,In_530);
nor U1536 (N_1536,In_4198,In_3619);
nor U1537 (N_1537,In_3632,In_4702);
nand U1538 (N_1538,In_63,In_644);
or U1539 (N_1539,In_57,In_4856);
and U1540 (N_1540,In_1136,In_1146);
or U1541 (N_1541,In_1063,In_4968);
nor U1542 (N_1542,In_1510,In_4811);
xnor U1543 (N_1543,In_1902,In_1876);
or U1544 (N_1544,In_70,In_4639);
and U1545 (N_1545,In_2972,In_4155);
nor U1546 (N_1546,In_4874,In_1301);
or U1547 (N_1547,In_3402,In_4900);
and U1548 (N_1548,In_3257,In_2553);
or U1549 (N_1549,In_3694,In_2348);
nor U1550 (N_1550,In_40,In_1719);
xnor U1551 (N_1551,In_4529,In_610);
or U1552 (N_1552,In_1888,In_940);
xnor U1553 (N_1553,In_3448,In_4648);
or U1554 (N_1554,In_1400,In_1281);
xor U1555 (N_1555,In_1285,In_1108);
and U1556 (N_1556,In_95,In_3622);
or U1557 (N_1557,In_1174,In_4719);
or U1558 (N_1558,In_1395,In_196);
nand U1559 (N_1559,In_3552,In_3327);
nand U1560 (N_1560,In_3022,In_4795);
or U1561 (N_1561,In_1018,In_3366);
and U1562 (N_1562,In_120,In_569);
xor U1563 (N_1563,In_3706,In_4392);
nor U1564 (N_1564,In_4045,In_3466);
and U1565 (N_1565,In_4376,In_1309);
nor U1566 (N_1566,In_3577,In_1625);
nor U1567 (N_1567,In_3750,In_4168);
and U1568 (N_1568,In_1093,In_3953);
nor U1569 (N_1569,In_1498,In_476);
nor U1570 (N_1570,In_1203,In_38);
nand U1571 (N_1571,In_102,In_4402);
xnor U1572 (N_1572,In_3100,In_281);
nor U1573 (N_1573,In_4905,In_2260);
and U1574 (N_1574,In_4324,In_883);
or U1575 (N_1575,In_2867,In_3977);
or U1576 (N_1576,In_3161,In_1427);
xor U1577 (N_1577,In_1881,In_890);
xor U1578 (N_1578,In_160,In_3163);
or U1579 (N_1579,In_1002,In_4366);
and U1580 (N_1580,In_838,In_2736);
xor U1581 (N_1581,In_4050,In_2498);
and U1582 (N_1582,In_2069,In_2458);
and U1583 (N_1583,In_2926,In_3459);
nand U1584 (N_1584,In_2906,In_1706);
and U1585 (N_1585,In_2615,In_4346);
or U1586 (N_1586,In_847,In_437);
xnor U1587 (N_1587,In_1272,In_3700);
and U1588 (N_1588,In_237,In_4843);
nor U1589 (N_1589,In_1772,In_4953);
and U1590 (N_1590,In_3629,In_4469);
xnor U1591 (N_1591,In_1986,In_2671);
or U1592 (N_1592,In_3009,In_797);
nor U1593 (N_1593,In_3606,In_4729);
or U1594 (N_1594,In_4937,In_3845);
nor U1595 (N_1595,In_2566,In_884);
or U1596 (N_1596,In_3500,In_1572);
nand U1597 (N_1597,In_922,In_2099);
or U1598 (N_1598,In_3154,In_1606);
xnor U1599 (N_1599,In_2515,In_2706);
nor U1600 (N_1600,In_4902,In_3756);
nor U1601 (N_1601,In_2500,In_3918);
xor U1602 (N_1602,In_1903,In_141);
xor U1603 (N_1603,In_3185,In_3449);
xor U1604 (N_1604,In_4116,In_3945);
and U1605 (N_1605,In_343,In_2653);
xnor U1606 (N_1606,In_4964,In_4354);
xnor U1607 (N_1607,In_1892,In_430);
nor U1608 (N_1608,In_3026,In_1592);
nor U1609 (N_1609,In_4740,In_3805);
xor U1610 (N_1610,In_1823,In_2805);
and U1611 (N_1611,In_3074,In_3608);
nand U1612 (N_1612,In_2996,In_2318);
or U1613 (N_1613,In_4362,In_2282);
or U1614 (N_1614,In_1027,In_2229);
and U1615 (N_1615,In_1471,In_877);
xor U1616 (N_1616,In_2019,In_59);
and U1617 (N_1617,In_4101,In_1934);
xnor U1618 (N_1618,In_1416,In_2902);
and U1619 (N_1619,In_2479,In_2418);
and U1620 (N_1620,In_3124,In_3256);
nor U1621 (N_1621,In_4331,In_4667);
nand U1622 (N_1622,In_2818,In_4457);
nor U1623 (N_1623,In_1208,In_2402);
xnor U1624 (N_1624,In_515,In_3355);
or U1625 (N_1625,In_2246,In_2591);
nand U1626 (N_1626,In_4887,In_2273);
and U1627 (N_1627,In_1769,In_3429);
and U1628 (N_1628,In_1286,In_4932);
and U1629 (N_1629,In_4776,In_1077);
or U1630 (N_1630,In_2383,In_2306);
nor U1631 (N_1631,In_4669,In_2421);
nor U1632 (N_1632,In_2250,In_669);
and U1633 (N_1633,In_3329,In_3241);
nor U1634 (N_1634,In_3092,In_3117);
or U1635 (N_1635,In_1023,In_3566);
and U1636 (N_1636,In_873,In_1276);
nor U1637 (N_1637,In_637,In_616);
and U1638 (N_1638,In_3725,In_355);
and U1639 (N_1639,In_1549,In_2118);
or U1640 (N_1640,In_4089,In_4939);
xor U1641 (N_1641,In_329,In_3463);
nor U1642 (N_1642,In_2437,In_4320);
nor U1643 (N_1643,In_1657,In_4398);
xor U1644 (N_1644,In_2376,In_2714);
and U1645 (N_1645,In_3381,In_4524);
nand U1646 (N_1646,In_4535,In_1869);
xnor U1647 (N_1647,In_2881,In_708);
xnor U1648 (N_1648,In_1838,In_882);
or U1649 (N_1649,In_4826,In_2467);
and U1650 (N_1650,In_1302,In_2832);
or U1651 (N_1651,In_4327,In_2904);
or U1652 (N_1652,In_4119,In_4800);
nand U1653 (N_1653,In_2484,In_2672);
and U1654 (N_1654,In_4644,In_3580);
xor U1655 (N_1655,In_2460,In_1938);
nor U1656 (N_1656,In_2683,In_97);
nor U1657 (N_1657,In_3639,In_3638);
nand U1658 (N_1658,In_58,In_720);
xnor U1659 (N_1659,In_2723,In_3051);
nand U1660 (N_1660,In_1388,In_4314);
nor U1661 (N_1661,In_86,In_4626);
xnor U1662 (N_1662,In_4583,In_2789);
or U1663 (N_1663,In_4816,In_4559);
nand U1664 (N_1664,In_4576,In_4762);
or U1665 (N_1665,In_1078,In_1579);
and U1666 (N_1666,In_836,In_250);
nand U1667 (N_1667,In_3340,In_1727);
xnor U1668 (N_1668,In_618,In_4203);
nand U1669 (N_1669,In_3922,In_271);
or U1670 (N_1670,In_264,In_3929);
xnor U1671 (N_1671,In_3261,In_3651);
and U1672 (N_1672,In_4044,In_3453);
and U1673 (N_1673,In_3319,In_409);
nand U1674 (N_1674,In_145,In_3891);
and U1675 (N_1675,In_4753,In_3249);
xor U1676 (N_1676,In_1761,In_2937);
or U1677 (N_1677,In_498,In_566);
or U1678 (N_1678,In_2287,In_1015);
or U1679 (N_1679,In_2550,In_1918);
or U1680 (N_1680,In_4148,In_3141);
nor U1681 (N_1681,In_3059,In_2711);
nand U1682 (N_1682,In_3582,In_912);
or U1683 (N_1683,In_1528,In_2788);
and U1684 (N_1684,In_3993,In_305);
and U1685 (N_1685,In_1525,In_1333);
nor U1686 (N_1686,In_243,In_1713);
xor U1687 (N_1687,In_96,In_907);
and U1688 (N_1688,In_2765,In_4737);
nand U1689 (N_1689,In_3741,In_4979);
nor U1690 (N_1690,In_3294,In_2530);
xor U1691 (N_1691,In_2980,In_1574);
and U1692 (N_1692,In_1737,In_3188);
nand U1693 (N_1693,In_3998,In_94);
or U1694 (N_1694,In_1643,In_4616);
xor U1695 (N_1695,In_4688,In_4105);
xnor U1696 (N_1696,In_1470,In_2012);
xor U1697 (N_1697,In_3235,In_815);
xnor U1698 (N_1698,In_1620,In_3476);
and U1699 (N_1699,In_1802,In_615);
nor U1700 (N_1700,In_42,In_2509);
and U1701 (N_1701,In_1369,In_3258);
and U1702 (N_1702,In_4947,In_2096);
and U1703 (N_1703,In_2251,In_1214);
or U1704 (N_1704,In_1865,In_4432);
or U1705 (N_1705,In_2194,In_654);
xnor U1706 (N_1706,In_4312,In_144);
nor U1707 (N_1707,In_4685,In_2428);
or U1708 (N_1708,In_1909,In_1336);
or U1709 (N_1709,In_4928,In_3705);
nand U1710 (N_1710,In_4142,In_1235);
or U1711 (N_1711,In_2556,In_2470);
nor U1712 (N_1712,In_981,In_2454);
nand U1713 (N_1713,In_4284,In_1096);
or U1714 (N_1714,In_467,In_2619);
xnor U1715 (N_1715,In_923,In_4003);
nor U1716 (N_1716,In_3662,In_3301);
xnor U1717 (N_1717,In_2334,In_3375);
xnor U1718 (N_1718,In_3691,In_3254);
and U1719 (N_1719,In_258,In_1071);
xor U1720 (N_1720,In_4697,In_148);
nand U1721 (N_1721,In_4632,In_579);
and U1722 (N_1722,In_1097,In_1045);
nand U1723 (N_1723,In_1111,In_4112);
and U1724 (N_1724,In_4961,In_1658);
and U1725 (N_1725,In_2164,In_2620);
or U1726 (N_1726,In_2147,In_1501);
and U1727 (N_1727,In_2106,In_2747);
or U1728 (N_1728,In_1161,In_2804);
and U1729 (N_1729,In_4020,In_888);
and U1730 (N_1730,In_3231,In_1553);
nand U1731 (N_1731,In_2032,In_1496);
nand U1732 (N_1732,In_1839,In_2362);
xnor U1733 (N_1733,In_943,In_1131);
xnor U1734 (N_1734,In_2299,In_3816);
nor U1735 (N_1735,In_39,In_539);
xor U1736 (N_1736,In_3636,In_2116);
nand U1737 (N_1737,In_685,In_3597);
nand U1738 (N_1738,In_2878,In_1776);
xor U1739 (N_1739,In_1444,In_299);
xor U1740 (N_1740,In_4094,In_282);
nand U1741 (N_1741,In_694,In_1322);
or U1742 (N_1742,In_2651,In_4512);
xnor U1743 (N_1743,In_1913,In_4024);
xnor U1744 (N_1744,In_4527,In_1791);
or U1745 (N_1745,In_3221,In_348);
nor U1746 (N_1746,In_3487,In_2784);
nor U1747 (N_1747,In_2385,In_3774);
nand U1748 (N_1748,In_3011,In_1516);
nand U1749 (N_1749,In_170,In_4504);
xnor U1750 (N_1750,In_4728,In_509);
xor U1751 (N_1751,In_4624,In_3367);
and U1752 (N_1752,In_4153,In_3455);
nand U1753 (N_1753,In_2461,In_4534);
nand U1754 (N_1754,In_3928,In_2125);
and U1755 (N_1755,In_693,In_4579);
xnor U1756 (N_1756,In_3077,In_1123);
or U1757 (N_1757,In_1389,In_221);
nand U1758 (N_1758,In_4683,In_1411);
nor U1759 (N_1759,In_3596,In_4460);
xor U1760 (N_1760,In_1497,In_3643);
nand U1761 (N_1761,In_3260,In_4282);
xnor U1762 (N_1762,In_567,In_3562);
nand U1763 (N_1763,In_3823,In_1576);
and U1764 (N_1764,In_2028,In_4732);
nor U1765 (N_1765,In_4945,In_3182);
and U1766 (N_1766,In_1634,In_1664);
xor U1767 (N_1767,In_472,In_4078);
nand U1768 (N_1768,In_268,In_382);
xnor U1769 (N_1769,In_519,In_1613);
or U1770 (N_1770,In_3361,In_1328);
xnor U1771 (N_1771,In_1543,In_3325);
and U1772 (N_1772,In_1750,In_1291);
and U1773 (N_1773,In_776,In_2420);
nor U1774 (N_1774,In_4361,In_894);
xor U1775 (N_1775,In_809,In_4166);
nor U1776 (N_1776,In_2870,In_3245);
nand U1777 (N_1777,In_2829,In_4814);
nand U1778 (N_1778,In_3938,In_3770);
and U1779 (N_1779,In_4940,In_4276);
xor U1780 (N_1780,In_1893,In_2679);
nor U1781 (N_1781,In_1796,In_1799);
nor U1782 (N_1782,In_187,In_4049);
and U1783 (N_1783,In_2392,In_1067);
nor U1784 (N_1784,In_4959,In_289);
nand U1785 (N_1785,In_3892,In_518);
or U1786 (N_1786,In_3489,In_2815);
nand U1787 (N_1787,In_1237,In_4240);
nor U1788 (N_1788,In_363,In_1197);
nand U1789 (N_1789,In_2890,In_4975);
nor U1790 (N_1790,In_1052,In_3550);
xor U1791 (N_1791,In_1334,In_2445);
and U1792 (N_1792,In_2860,In_2369);
nor U1793 (N_1793,In_846,In_2041);
and U1794 (N_1794,In_3491,In_1121);
nand U1795 (N_1795,In_1757,In_4621);
xor U1796 (N_1796,In_1218,In_3976);
nor U1797 (N_1797,In_1689,In_1783);
xnor U1798 (N_1798,In_4477,In_1042);
nor U1799 (N_1799,In_3510,In_2654);
nor U1800 (N_1800,In_3465,In_2453);
xnor U1801 (N_1801,In_2923,In_1271);
xor U1802 (N_1802,In_2351,In_4374);
xnor U1803 (N_1803,In_2195,In_3519);
xor U1804 (N_1804,In_4408,In_714);
and U1805 (N_1805,In_2483,In_4674);
or U1806 (N_1806,In_3331,In_3640);
and U1807 (N_1807,In_2075,In_795);
nor U1808 (N_1808,In_50,In_1139);
or U1809 (N_1809,In_1920,In_2359);
and U1810 (N_1810,In_921,In_4085);
nand U1811 (N_1811,In_1760,In_2775);
nor U1812 (N_1812,In_2444,In_2623);
and U1813 (N_1813,In_4888,In_2442);
and U1814 (N_1814,In_4090,In_1532);
xor U1815 (N_1815,In_2224,In_2625);
or U1816 (N_1816,In_1038,In_4507);
nor U1817 (N_1817,In_1650,In_2481);
and U1818 (N_1818,In_2704,In_2608);
xor U1819 (N_1819,In_724,In_2478);
nor U1820 (N_1820,In_1412,In_1261);
and U1821 (N_1821,In_4205,In_3469);
nand U1822 (N_1822,In_1415,In_2008);
nor U1823 (N_1823,In_4308,In_2979);
and U1824 (N_1824,In_3234,In_3520);
or U1825 (N_1825,In_4595,In_2741);
nand U1826 (N_1826,In_4470,In_2365);
or U1827 (N_1827,In_2944,In_219);
or U1828 (N_1828,In_2280,In_2782);
or U1829 (N_1829,In_1752,In_2013);
and U1830 (N_1830,In_2925,In_4301);
and U1831 (N_1831,In_4827,In_3620);
xnor U1832 (N_1832,In_3772,In_3794);
or U1833 (N_1833,In_115,In_749);
xor U1834 (N_1834,In_1029,In_2582);
or U1835 (N_1835,In_729,In_4839);
nand U1836 (N_1836,In_4349,In_3598);
xor U1837 (N_1837,In_136,In_2399);
and U1838 (N_1838,In_1843,In_629);
nor U1839 (N_1839,In_2007,In_1189);
nand U1840 (N_1840,In_3693,In_3853);
or U1841 (N_1841,In_1536,In_113);
or U1842 (N_1842,In_3427,In_2677);
xnor U1843 (N_1843,In_4759,In_810);
nor U1844 (N_1844,In_665,In_146);
and U1845 (N_1845,In_2139,In_2959);
or U1846 (N_1846,In_4415,In_1106);
xor U1847 (N_1847,In_3980,In_2587);
nand U1848 (N_1848,In_327,In_441);
nand U1849 (N_1849,In_857,In_4289);
and U1850 (N_1850,In_230,In_964);
and U1851 (N_1851,In_1345,In_4418);
nor U1852 (N_1852,In_1992,In_4891);
nand U1853 (N_1853,In_526,In_3058);
xor U1854 (N_1854,In_1633,In_1381);
or U1855 (N_1855,In_2159,In_4200);
or U1856 (N_1856,In_2145,In_3856);
nor U1857 (N_1857,In_532,In_4311);
nor U1858 (N_1858,In_4861,In_706);
or U1859 (N_1859,In_3056,In_1114);
xnor U1860 (N_1860,In_4250,In_1332);
or U1861 (N_1861,In_4752,In_2879);
nor U1862 (N_1862,In_1069,In_2436);
or U1863 (N_1863,In_2750,In_2900);
xnor U1864 (N_1864,In_3763,In_3924);
or U1865 (N_1865,In_1360,In_1725);
nand U1866 (N_1866,In_726,In_3422);
xnor U1867 (N_1867,In_649,In_2920);
or U1868 (N_1868,In_446,In_3969);
nor U1869 (N_1869,In_2192,In_3127);
and U1870 (N_1870,In_1448,In_4723);
xor U1871 (N_1871,In_632,In_4601);
nand U1872 (N_1872,In_2384,In_2584);
nand U1873 (N_1873,In_4584,In_333);
nand U1874 (N_1874,In_1779,In_2773);
or U1875 (N_1875,In_2738,In_2709);
and U1876 (N_1876,In_633,In_89);
and U1877 (N_1877,In_1153,In_910);
nand U1878 (N_1878,In_4558,In_4356);
or U1879 (N_1879,In_4613,In_4542);
xnor U1880 (N_1880,In_4010,In_735);
nand U1881 (N_1881,In_3637,In_1226);
or U1882 (N_1882,In_2950,In_4549);
and U1883 (N_1883,In_2230,In_3395);
and U1884 (N_1884,In_3363,In_4805);
nor U1885 (N_1885,In_391,In_2379);
xor U1886 (N_1886,In_489,In_4341);
nand U1887 (N_1887,In_1964,In_4357);
and U1888 (N_1888,In_3160,In_1599);
and U1889 (N_1889,In_2029,In_3166);
nand U1890 (N_1890,In_3635,In_1819);
nand U1891 (N_1891,In_4231,In_4363);
and U1892 (N_1892,In_2565,In_2346);
xor U1893 (N_1893,In_3444,In_790);
nand U1894 (N_1894,In_4517,In_2532);
nand U1895 (N_1895,In_4948,In_535);
or U1896 (N_1896,In_4048,In_3593);
xor U1897 (N_1897,In_2695,In_1475);
or U1898 (N_1898,In_4665,In_2967);
and U1899 (N_1899,In_1180,In_686);
nand U1900 (N_1900,In_2494,In_2737);
and U1901 (N_1901,In_571,In_4538);
xnor U1902 (N_1902,In_307,In_1696);
or U1903 (N_1903,In_1103,In_4966);
xnor U1904 (N_1904,In_1955,In_909);
xnor U1905 (N_1905,In_1181,In_2975);
or U1906 (N_1906,In_2799,In_3411);
or U1907 (N_1907,In_759,In_2525);
xor U1908 (N_1908,In_1089,In_2928);
nor U1909 (N_1909,In_3253,In_3965);
or U1910 (N_1910,In_400,In_4455);
and U1911 (N_1911,In_4660,In_4877);
and U1912 (N_1912,In_1115,In_2754);
nand U1913 (N_1913,In_3542,In_3886);
nor U1914 (N_1914,In_3882,In_4143);
or U1915 (N_1915,In_3759,In_2702);
nor U1916 (N_1916,In_2533,In_2892);
nor U1917 (N_1917,In_3648,In_3330);
or U1918 (N_1918,In_584,In_4479);
xor U1919 (N_1919,In_1575,In_2127);
nor U1920 (N_1920,In_4441,In_181);
and U1921 (N_1921,In_2308,In_1408);
or U1922 (N_1922,In_2206,In_1422);
or U1923 (N_1923,In_829,In_190);
nand U1924 (N_1924,In_2114,In_1585);
and U1925 (N_1925,In_4815,In_3645);
xnor U1926 (N_1926,In_2073,In_878);
or U1927 (N_1927,In_2602,In_502);
and U1928 (N_1928,In_3285,In_581);
nand U1929 (N_1929,In_807,In_3019);
xor U1930 (N_1930,In_4167,In_4244);
xnor U1931 (N_1931,In_1652,In_4072);
and U1932 (N_1932,In_353,In_451);
nand U1933 (N_1933,In_1789,In_1032);
or U1934 (N_1934,In_4692,In_3075);
and U1935 (N_1935,In_1465,In_1996);
nand U1936 (N_1936,In_3859,In_1393);
xor U1937 (N_1937,In_1298,In_4204);
xnor U1938 (N_1938,In_1329,In_960);
nor U1939 (N_1939,In_2964,In_3955);
nor U1940 (N_1940,In_4764,In_3452);
or U1941 (N_1941,In_769,In_2220);
nand U1942 (N_1942,In_1742,In_4608);
and U1943 (N_1943,In_470,In_2163);
and U1944 (N_1944,In_1219,In_1337);
nor U1945 (N_1945,In_1611,In_291);
xnor U1946 (N_1946,In_3728,In_3291);
nor U1947 (N_1947,In_4634,In_3339);
xor U1948 (N_1948,In_4310,In_3588);
and U1949 (N_1949,In_4288,In_3656);
or U1950 (N_1950,In_354,In_2650);
xnor U1951 (N_1951,In_4924,In_4433);
and U1952 (N_1952,In_700,In_4058);
and U1953 (N_1953,In_4041,In_4380);
and U1954 (N_1954,In_3936,In_1998);
nor U1955 (N_1955,In_3279,In_1513);
nand U1956 (N_1956,In_4710,In_3324);
nand U1957 (N_1957,In_728,In_2819);
nand U1958 (N_1958,In_2973,In_2594);
or U1959 (N_1959,In_2947,In_336);
or U1960 (N_1960,In_1432,In_1168);
and U1961 (N_1961,In_2283,In_1001);
xnor U1962 (N_1962,In_675,In_4439);
nor U1963 (N_1963,In_1354,In_2004);
nand U1964 (N_1964,In_1953,In_4210);
or U1965 (N_1965,In_2713,In_3565);
xor U1966 (N_1966,In_4121,In_1921);
or U1967 (N_1967,In_3297,In_2969);
and U1968 (N_1968,In_4989,In_2225);
and U1969 (N_1969,In_1672,In_3200);
nand U1970 (N_1970,In_562,In_1206);
nor U1971 (N_1971,In_4784,In_3769);
nand U1972 (N_1972,In_4221,In_3431);
or U1973 (N_1973,In_4894,In_2316);
or U1974 (N_1974,In_3504,In_4757);
xor U1975 (N_1975,In_3035,In_876);
and U1976 (N_1976,In_709,In_304);
xnor U1977 (N_1977,In_2681,In_3106);
nor U1978 (N_1978,In_1490,In_4287);
nand U1979 (N_1979,In_1087,In_2214);
xnor U1980 (N_1980,In_2005,In_4472);
and U1981 (N_1981,In_4442,In_4857);
and U1982 (N_1982,In_3675,In_4389);
nand U1983 (N_1983,In_1669,In_998);
nand U1984 (N_1984,In_4926,In_2367);
or U1985 (N_1985,In_506,In_2957);
or U1986 (N_1986,In_1774,In_2544);
nor U1987 (N_1987,In_2294,In_3384);
and U1988 (N_1988,In_48,In_4319);
xor U1989 (N_1989,In_2540,In_3179);
nor U1990 (N_1990,In_1589,In_3321);
xnor U1991 (N_1991,In_1384,In_985);
or U1992 (N_1992,In_4079,In_4550);
and U1993 (N_1993,In_915,In_648);
nor U1994 (N_1994,In_3148,In_267);
nand U1995 (N_1995,In_2360,In_2567);
and U1996 (N_1996,In_3867,In_1744);
nand U1997 (N_1997,In_4568,In_4834);
and U1998 (N_1998,In_3017,In_1878);
or U1999 (N_1999,In_195,In_3267);
xnor U2000 (N_2000,N_1292,In_4615);
and U2001 (N_2001,In_2111,N_236);
xnor U2002 (N_2002,N_915,In_1049);
and U2003 (N_2003,N_1842,In_147);
nand U2004 (N_2004,N_1460,In_3263);
or U2005 (N_2005,N_1222,N_308);
nand U2006 (N_2006,In_891,N_844);
or U2007 (N_2007,N_562,N_198);
or U2008 (N_2008,In_4984,N_1283);
or U2009 (N_2009,N_1323,N_1567);
and U2010 (N_2010,In_3894,N_1949);
or U2011 (N_2011,N_654,In_851);
and U2012 (N_2012,In_1488,N_1582);
nand U2013 (N_2013,N_807,N_27);
or U2014 (N_2014,N_329,N_1766);
nor U2015 (N_2015,N_338,In_3368);
or U2016 (N_2016,N_760,N_1628);
or U2017 (N_2017,In_589,In_111);
xor U2018 (N_2018,N_1526,N_1458);
nor U2019 (N_2019,In_2857,N_1332);
and U2020 (N_2020,In_4533,N_511);
xor U2021 (N_2021,N_788,N_1330);
nor U2022 (N_2022,N_720,N_1340);
nand U2023 (N_2023,In_1122,N_349);
or U2024 (N_2024,N_1854,N_73);
xnor U2025 (N_2025,N_166,In_3468);
xor U2026 (N_2026,N_67,In_167);
and U2027 (N_2027,In_4944,N_1907);
and U2028 (N_2028,N_1378,N_361);
xnor U2029 (N_2029,N_1345,In_635);
xor U2030 (N_2030,N_846,N_1686);
nor U2031 (N_2031,N_140,In_2153);
nor U2032 (N_2032,N_1462,N_1835);
and U2033 (N_2033,N_974,In_3875);
or U2034 (N_2034,In_3813,In_2189);
and U2035 (N_2035,In_1057,N_417);
and U2036 (N_2036,In_4375,N_1825);
xor U2037 (N_2037,N_670,In_3496);
and U2038 (N_2038,In_4539,N_780);
nor U2039 (N_2039,In_4848,In_1409);
nand U2040 (N_2040,N_687,N_52);
xnor U2041 (N_2041,In_4406,N_21);
and U2042 (N_2042,N_1651,N_328);
or U2043 (N_2043,In_3492,N_115);
and U2044 (N_2044,N_255,N_1827);
or U2045 (N_2045,In_4377,N_1393);
nor U2046 (N_2046,N_191,N_304);
xor U2047 (N_2047,In_1790,N_1256);
xnor U2048 (N_2048,N_1273,N_958);
nand U2049 (N_2049,N_403,N_634);
or U2050 (N_2050,N_1897,N_681);
xor U2051 (N_2051,N_1068,N_596);
xnor U2052 (N_2052,N_1151,N_264);
and U2053 (N_2053,N_1685,In_4911);
or U2054 (N_2054,N_1851,N_1809);
nand U2055 (N_2055,In_2030,N_220);
and U2056 (N_2056,N_545,In_1290);
and U2057 (N_2057,N_1886,N_1317);
nand U2058 (N_2058,N_369,N_411);
nand U2059 (N_2059,In_1222,N_649);
xor U2060 (N_2060,N_663,N_1883);
xor U2061 (N_2061,N_109,N_1208);
or U2062 (N_2062,N_1972,N_1414);
and U2063 (N_2063,N_1565,N_307);
or U2064 (N_2064,N_898,N_997);
nand U2065 (N_2065,N_1060,In_2297);
xnor U2066 (N_2066,N_1621,In_1777);
and U2067 (N_2067,N_252,N_1138);
or U2068 (N_2068,N_449,In_980);
nor U2069 (N_2069,In_1274,N_1010);
nand U2070 (N_2070,In_2742,N_697);
xnor U2071 (N_2071,In_4333,In_969);
nand U2072 (N_2072,In_2422,In_1603);
xnor U2073 (N_2073,N_1871,In_1249);
and U2074 (N_2074,N_492,N_53);
and U2075 (N_2075,N_673,In_520);
nand U2076 (N_2076,In_1954,N_344);
or U2077 (N_2077,In_2953,N_1027);
nor U2078 (N_2078,In_1494,N_1302);
or U2079 (N_2079,N_1641,In_2946);
and U2080 (N_2080,N_409,N_1744);
or U2081 (N_2081,N_322,N_646);
nand U2082 (N_2082,N_1384,N_785);
or U2083 (N_2083,In_373,In_1520);
nor U2084 (N_2084,N_1404,In_4859);
nand U2085 (N_2085,N_1141,N_1596);
nor U2086 (N_2086,In_325,N_913);
or U2087 (N_2087,N_917,In_408);
nor U2088 (N_2088,N_1499,In_3483);
nor U2089 (N_2089,N_1855,N_540);
nand U2090 (N_2090,N_832,N_490);
nand U2091 (N_2091,N_20,N_1690);
nand U2092 (N_2092,N_1087,N_1626);
nor U2093 (N_2093,N_1609,N_139);
nand U2094 (N_2094,N_291,In_3773);
nand U2095 (N_2095,N_1610,In_117);
and U2096 (N_2096,N_1959,N_106);
and U2097 (N_2097,N_127,N_1576);
and U2098 (N_2098,In_227,In_3761);
and U2099 (N_2099,N_742,N_1356);
nand U2100 (N_2100,In_3786,N_566);
nor U2101 (N_2101,N_1873,N_1017);
xor U2102 (N_2102,N_143,In_211);
nand U2103 (N_2103,N_769,N_851);
nor U2104 (N_2104,N_1425,N_1718);
and U2105 (N_2105,N_1183,In_25);
nand U2106 (N_2106,N_1877,N_327);
xor U2107 (N_2107,N_239,N_1960);
nand U2108 (N_2108,N_1966,In_2913);
and U2109 (N_2109,N_721,In_831);
xor U2110 (N_2110,In_1977,N_1019);
xor U2111 (N_2111,In_3558,In_4000);
xor U2112 (N_2112,N_1599,In_4906);
or U2113 (N_2113,In_3917,In_4281);
or U2114 (N_2114,N_334,N_1798);
or U2115 (N_2115,N_1008,N_1494);
nor U2116 (N_2116,In_4766,N_521);
xor U2117 (N_2117,N_543,N_1857);
nor U2118 (N_2118,In_697,In_1377);
or U2119 (N_2119,In_3486,N_645);
or U2120 (N_2120,In_1250,In_4724);
or U2121 (N_2121,N_1900,N_96);
or U2122 (N_2122,N_1450,N_1901);
nand U2123 (N_2123,In_1905,In_2086);
and U2124 (N_2124,In_3839,In_3250);
and U2125 (N_2125,N_1716,In_2016);
nor U2126 (N_2126,In_2601,N_957);
or U2127 (N_2127,N_1220,N_394);
nand U2128 (N_2128,In_1810,N_1046);
nand U2129 (N_2129,N_847,In_3370);
nor U2130 (N_2130,N_1181,N_1354);
xnor U2131 (N_2131,N_964,In_1129);
xnor U2132 (N_2132,N_279,N_550);
nand U2133 (N_2133,In_2160,N_1074);
nor U2134 (N_2134,N_26,In_2221);
xor U2135 (N_2135,N_1627,N_1633);
nor U2136 (N_2136,N_1538,N_700);
or U2137 (N_2137,N_342,In_4043);
nor U2138 (N_2138,In_2665,N_850);
nand U2139 (N_2139,N_859,N_1575);
and U2140 (N_2140,N_909,N_1786);
nand U2141 (N_2141,N_454,In_3775);
nand U2142 (N_2142,In_2274,In_4770);
xor U2143 (N_2143,In_1101,In_3176);
nand U2144 (N_2144,N_1380,N_458);
or U2145 (N_2145,N_1693,N_1096);
nand U2146 (N_2146,N_1740,N_435);
nand U2147 (N_2147,In_3404,In_3671);
nor U2148 (N_2148,N_1615,N_1457);
and U2149 (N_2149,N_897,N_1915);
nand U2150 (N_2150,N_1142,N_1580);
nor U2151 (N_2151,N_1160,N_1926);
nor U2152 (N_2152,N_376,In_1758);
xor U2153 (N_2153,In_3605,N_1149);
or U2154 (N_2154,N_598,N_1466);
nor U2155 (N_2155,In_4122,In_1628);
nor U2156 (N_2156,In_4809,N_1469);
nand U2157 (N_2157,N_294,N_1122);
or U2158 (N_2158,In_339,N_1713);
nand U2159 (N_2159,N_426,N_1733);
or U2160 (N_2160,In_4007,In_3988);
nor U2161 (N_2161,N_740,N_1089);
xnor U2162 (N_2162,N_1334,In_1259);
and U2163 (N_2163,N_541,In_3039);
or U2164 (N_2164,N_714,N_331);
or U2165 (N_2165,N_158,In_588);
and U2166 (N_2166,In_3669,N_1105);
or U2167 (N_2167,N_612,N_1370);
and U2168 (N_2168,N_1824,N_1778);
or U2169 (N_2169,N_1416,In_3289);
and U2170 (N_2170,N_1171,N_65);
nor U2171 (N_2171,N_1903,N_980);
xor U2172 (N_2172,N_1773,In_2150);
nor U2173 (N_2173,In_2774,N_1263);
xnor U2174 (N_2174,N_1495,N_1026);
or U2175 (N_2175,N_1880,N_484);
nand U2176 (N_2176,In_2664,N_87);
xnor U2177 (N_2177,In_1245,In_4322);
xor U2178 (N_2178,In_908,N_23);
nand U2179 (N_2179,In_3714,N_1608);
or U2180 (N_2180,N_1318,N_1724);
and U2181 (N_2181,N_1412,In_4297);
and U2182 (N_2182,N_1396,N_1203);
nor U2183 (N_2183,In_2646,N_296);
nor U2184 (N_2184,N_1697,In_2976);
nand U2185 (N_2185,N_1107,N_1187);
or U2186 (N_2186,In_4420,N_1392);
or U2187 (N_2187,N_1422,N_93);
or U2188 (N_2188,In_2087,N_385);
or U2189 (N_2189,N_1209,In_3194);
or U2190 (N_2190,N_414,N_757);
or U2191 (N_2191,N_778,N_48);
and U2192 (N_2192,N_430,N_1573);
nor U2193 (N_2193,N_1213,N_1583);
and U2194 (N_2194,In_4962,N_1005);
nand U2195 (N_2195,In_2893,N_1849);
nor U2196 (N_2196,N_1401,N_767);
nor U2197 (N_2197,N_1435,N_1981);
nand U2198 (N_2198,In_493,N_1524);
and U2199 (N_2199,N_938,N_1834);
or U2200 (N_2200,In_1566,N_1612);
xnor U2201 (N_2201,N_130,In_1505);
or U2202 (N_2202,N_836,N_33);
nor U2203 (N_2203,N_708,N_1566);
xnor U2204 (N_2204,N_1359,N_639);
xor U2205 (N_2205,N_841,N_1048);
or U2206 (N_2206,N_928,N_1281);
xor U2207 (N_2207,In_2896,In_3826);
nor U2208 (N_2208,N_852,N_1833);
nand U2209 (N_2209,In_2234,N_1158);
nor U2210 (N_2210,N_422,N_315);
xnor U2211 (N_2211,N_1173,N_1982);
nand U2212 (N_2212,N_1182,In_503);
xor U2213 (N_2213,N_1073,N_1777);
nor U2214 (N_2214,N_1639,N_1682);
xnor U2215 (N_2215,In_781,N_886);
nand U2216 (N_2216,In_1581,In_3850);
nor U2217 (N_2217,N_386,In_2245);
or U2218 (N_2218,N_1124,N_1031);
xor U2219 (N_2219,In_19,In_3967);
or U2220 (N_2220,In_4537,In_2935);
or U2221 (N_2221,N_1063,In_3113);
or U2222 (N_2222,N_129,N_108);
or U2223 (N_2223,N_660,N_148);
xnor U2224 (N_2224,In_4712,In_418);
xnor U2225 (N_2225,N_513,In_2746);
xor U2226 (N_2226,N_683,N_819);
and U2227 (N_2227,In_3946,N_1109);
nand U2228 (N_2228,N_1887,In_984);
nor U2229 (N_2229,N_1348,N_1324);
nor U2230 (N_2230,N_734,N_230);
nor U2231 (N_2231,N_15,N_506);
nor U2232 (N_2232,N_1386,N_1398);
or U2233 (N_2233,In_4124,N_442);
nand U2234 (N_2234,N_1644,N_1658);
nor U2235 (N_2235,In_2748,N_337);
or U2236 (N_2236,In_3169,N_1968);
xor U2237 (N_2237,N_363,N_1817);
nand U2238 (N_2238,N_880,N_1705);
nor U2239 (N_2239,In_2974,In_272);
xor U2240 (N_2240,In_4897,N_515);
and U2241 (N_2241,In_56,N_1793);
xor U2242 (N_2242,N_1061,N_214);
or U2243 (N_2243,N_1315,N_1795);
xnor U2244 (N_2244,N_786,N_95);
and U2245 (N_2245,N_491,N_677);
nor U2246 (N_2246,N_514,In_4528);
nor U2247 (N_2247,In_2701,In_2081);
and U2248 (N_2248,N_893,N_16);
or U2249 (N_2249,N_1988,N_927);
and U2250 (N_2250,In_1183,N_494);
xnor U2251 (N_2251,In_1936,N_1092);
and U2252 (N_2252,In_1177,In_4872);
nand U2253 (N_2253,N_963,N_357);
nand U2254 (N_2254,N_1681,N_1975);
nor U2255 (N_2255,In_1835,N_1379);
nand U2256 (N_2256,In_3726,In_3921);
or U2257 (N_2257,In_3654,In_4997);
and U2258 (N_2258,N_1936,In_1753);
or U2259 (N_2259,In_3824,N_43);
nor U2260 (N_2260,In_3454,N_664);
xor U2261 (N_2261,In_1915,N_895);
xnor U2262 (N_2262,In_3527,N_621);
and U2263 (N_2263,In_3844,In_3873);
xor U2264 (N_2264,N_1179,N_1420);
nand U2265 (N_2265,In_1736,N_295);
xor U2266 (N_2266,N_1339,In_4272);
nor U2267 (N_2267,In_1073,N_476);
nand U2268 (N_2268,In_3818,In_1722);
or U2269 (N_2269,N_877,N_1542);
nor U2270 (N_2270,N_1042,N_485);
xnor U2271 (N_2271,N_1956,N_1030);
xnor U2272 (N_2272,N_172,In_3944);
and U2273 (N_2273,In_3685,In_3246);
and U2274 (N_2274,N_58,N_1312);
nor U2275 (N_2275,N_11,N_1440);
nand U2276 (N_2276,In_3354,In_3287);
nand U2277 (N_2277,In_2684,N_99);
and U2278 (N_2278,In_4474,In_1211);
nor U2279 (N_2279,N_1360,N_1207);
and U2280 (N_2280,N_1560,N_587);
or U2281 (N_2281,N_1168,In_2828);
nand U2282 (N_2282,N_419,In_369);
nand U2283 (N_2283,N_1298,In_328);
nand U2284 (N_2284,N_592,N_1590);
nor U2285 (N_2285,In_3538,In_782);
or U2286 (N_2286,In_4388,N_1328);
and U2287 (N_2287,N_1971,N_1050);
or U2288 (N_2288,In_3655,N_474);
nor U2289 (N_2289,N_178,In_4867);
xnor U2290 (N_2290,In_3893,In_4605);
nand U2291 (N_2291,N_1989,In_3721);
xor U2292 (N_2292,N_1625,N_5);
or U2293 (N_2293,In_4290,N_1876);
nor U2294 (N_2294,N_656,N_94);
xnor U2295 (N_2295,In_1056,N_1091);
xor U2296 (N_2296,N_246,In_2721);
or U2297 (N_2297,N_1372,N_1478);
nand U2298 (N_2298,N_795,N_1467);
nand U2299 (N_2299,In_1196,In_895);
xor U2300 (N_2300,N_354,N_1453);
or U2301 (N_2301,N_1976,N_584);
xnor U2302 (N_2302,In_4876,N_726);
xor U2303 (N_2303,In_1198,N_1243);
xnor U2304 (N_2304,In_4844,N_1572);
and U2305 (N_2305,In_2052,In_421);
nand U2306 (N_2306,N_1252,N_59);
nor U2307 (N_2307,N_838,N_512);
or U2308 (N_2308,In_1642,In_350);
nand U2309 (N_2309,N_270,N_215);
xnor U2310 (N_2310,N_1365,N_1133);
or U2311 (N_2311,N_450,In_2278);
nor U2312 (N_2312,N_642,N_370);
and U2313 (N_2313,N_273,In_3450);
nand U2314 (N_2314,N_1800,N_534);
or U2315 (N_2315,N_420,N_131);
or U2316 (N_2316,N_352,N_197);
or U2317 (N_2317,N_991,In_263);
nor U2318 (N_2318,N_168,In_2573);
nor U2319 (N_2319,N_1586,N_632);
and U2320 (N_2320,In_4955,N_472);
nor U2321 (N_2321,N_790,N_1523);
xnor U2322 (N_2322,N_1383,N_546);
and U2323 (N_2323,N_1593,N_1863);
xnor U2324 (N_2324,In_2146,N_1254);
and U2325 (N_2325,N_1210,N_1858);
xnor U2326 (N_2326,N_1659,N_1204);
nand U2327 (N_2327,N_339,In_4355);
nand U2328 (N_2328,N_1,N_1443);
nor U2329 (N_2329,In_4152,In_1107);
nand U2330 (N_2330,N_750,N_896);
xor U2331 (N_2331,N_1023,In_3758);
or U2332 (N_2332,N_1137,N_725);
or U2333 (N_2333,N_1251,In_2156);
or U2334 (N_2334,N_74,In_1423);
nand U2335 (N_2335,N_932,N_1922);
nor U2336 (N_2336,N_862,In_4916);
nand U2337 (N_2337,N_1902,In_4194);
and U2338 (N_2338,N_901,N_1121);
or U2339 (N_2339,N_1812,N_702);
and U2340 (N_2340,N_519,N_35);
nor U2341 (N_2341,N_288,N_1894);
xnor U2342 (N_2342,N_1914,In_4187);
xor U2343 (N_2343,In_2968,N_1941);
and U2344 (N_2344,In_2961,N_715);
nand U2345 (N_2345,N_1844,N_22);
xnor U2346 (N_2346,N_1135,In_3791);
nor U2347 (N_2347,N_1057,N_1081);
and U2348 (N_2348,N_812,In_4269);
nand U2349 (N_2349,N_1674,N_659);
nor U2350 (N_2350,In_75,N_589);
nor U2351 (N_2351,N_1634,In_4515);
xnor U2352 (N_2352,N_1226,N_865);
xnor U2353 (N_2353,N_696,In_1192);
and U2354 (N_2354,In_1925,In_3156);
nor U2355 (N_2355,In_932,N_855);
or U2356 (N_2356,In_3812,N_1299);
or U2357 (N_2357,In_2155,N_1369);
xnor U2358 (N_2358,In_3642,N_1022);
nor U2359 (N_2359,N_183,N_1197);
or U2360 (N_2360,N_1688,N_833);
nor U2361 (N_2361,N_804,N_1637);
xnor U2362 (N_2362,N_14,In_4645);
nand U2363 (N_2363,In_4302,N_223);
nand U2364 (N_2364,In_885,N_1244);
or U2365 (N_2365,In_800,N_1034);
nor U2366 (N_2366,N_365,N_1167);
or U2367 (N_2367,In_3939,N_310);
and U2368 (N_2368,In_4545,In_2152);
or U2369 (N_2369,N_1564,N_1177);
and U2370 (N_2370,N_177,In_426);
nor U2371 (N_2371,In_4353,N_62);
or U2372 (N_2372,N_1667,N_447);
or U2373 (N_2373,N_1130,N_799);
nand U2374 (N_2374,N_817,In_2209);
and U2375 (N_2375,N_1445,N_107);
or U2376 (N_2376,N_1647,In_2716);
nand U2377 (N_2377,In_76,N_1571);
xnor U2378 (N_2378,N_406,In_334);
xnor U2379 (N_2379,N_1743,N_1215);
xnor U2380 (N_2380,N_10,N_50);
nand U2381 (N_2381,In_4571,In_2883);
and U2382 (N_2382,In_4662,In_3672);
nor U2383 (N_2383,N_1513,In_2989);
or U2384 (N_2384,In_1088,N_635);
nor U2385 (N_2385,N_613,N_1881);
xnor U2386 (N_2386,N_1522,N_395);
nand U2387 (N_2387,N_1832,N_532);
or U2388 (N_2388,In_4520,N_1280);
xnor U2389 (N_2389,N_391,N_1470);
or U2390 (N_2390,N_1071,In_3180);
nor U2391 (N_2391,N_468,In_3268);
and U2392 (N_2392,In_2115,N_818);
nand U2393 (N_2393,N_1136,N_1908);
nand U2394 (N_2394,N_1860,N_1350);
nor U2395 (N_2395,In_1223,In_2597);
xnor U2396 (N_2396,N_1162,In_2056);
nor U2397 (N_2397,N_1043,N_908);
or U2398 (N_2398,N_1558,In_1568);
nand U2399 (N_2399,In_1655,In_4495);
or U2400 (N_2400,In_1570,N_1840);
xnor U2401 (N_2401,N_1058,N_1347);
nor U2402 (N_2402,N_1112,In_2335);
xnor U2403 (N_2403,In_432,N_1804);
nand U2404 (N_2404,N_544,In_2243);
nor U2405 (N_2405,In_471,N_1150);
or U2406 (N_2406,N_610,N_1521);
and U2407 (N_2407,N_1728,N_501);
and U2408 (N_2408,In_2633,N_1427);
or U2409 (N_2409,In_4385,N_1601);
and U2410 (N_2410,In_4636,N_425);
xnor U2411 (N_2411,In_3628,In_4506);
or U2412 (N_2412,In_2128,N_1020);
xnor U2413 (N_2413,N_1540,N_561);
and U2414 (N_2414,N_40,In_1262);
nand U2415 (N_2415,N_1993,N_1719);
or U2416 (N_2416,In_1282,In_1738);
nor U2417 (N_2417,In_2562,In_1529);
xnor U2418 (N_2418,In_2869,N_1148);
nor U2419 (N_2419,N_175,N_1442);
or U2420 (N_2420,N_1206,N_1623);
nor U2421 (N_2421,N_1090,N_955);
xnor U2422 (N_2422,In_308,N_418);
or U2423 (N_2423,N_845,N_528);
and U2424 (N_2424,In_1948,N_1617);
nor U2425 (N_2425,N_966,In_4125);
nand U2426 (N_2426,In_2204,N_60);
nand U2427 (N_2427,In_1854,In_3177);
or U2428 (N_2428,N_377,In_3745);
xor U2429 (N_2429,In_138,N_555);
nor U2430 (N_2430,N_1164,N_1117);
xor U2431 (N_2431,N_1992,N_793);
or U2432 (N_2432,N_1753,In_2098);
nand U2433 (N_2433,In_2227,N_186);
nand U2434 (N_2434,N_247,N_1578);
nand U2435 (N_2435,N_1534,N_668);
xnor U2436 (N_2436,In_1804,N_611);
or U2437 (N_2437,N_1361,N_258);
nor U2438 (N_2438,N_1441,In_2751);
nand U2439 (N_2439,N_568,N_1911);
and U2440 (N_2440,N_142,N_1920);
nor U2441 (N_2441,N_661,N_1484);
nand U2442 (N_2442,N_749,In_2538);
or U2443 (N_2443,N_362,In_3271);
nand U2444 (N_2444,In_293,N_358);
and U2445 (N_2445,In_3195,N_1984);
or U2446 (N_2446,N_1219,N_234);
xnor U2447 (N_2447,In_602,N_771);
nand U2448 (N_2448,In_3533,In_2388);
or U2449 (N_2449,In_3530,N_1896);
or U2450 (N_2450,In_1240,In_1593);
nand U2451 (N_2451,N_1270,N_1706);
nand U2452 (N_2452,N_557,N_128);
and U2453 (N_2453,In_2258,N_405);
nor U2454 (N_2454,N_1668,In_1534);
nor U2455 (N_2455,N_1025,N_1620);
or U2456 (N_2456,N_1791,N_1650);
nor U2457 (N_2457,In_376,In_4199);
xnor U2458 (N_2458,In_77,N_1771);
and U2459 (N_2459,N_1191,N_1326);
and U2460 (N_2460,N_97,N_1548);
nand U2461 (N_2461,N_1843,In_619);
and U2462 (N_2462,N_290,N_1895);
xor U2463 (N_2463,N_160,N_1391);
xnor U2464 (N_2464,In_74,In_3677);
and U2465 (N_2465,N_1672,N_111);
nand U2466 (N_2466,N_585,N_1665);
or U2467 (N_2467,N_1788,N_504);
and U2468 (N_2468,In_2404,N_7);
xor U2469 (N_2469,N_1581,N_1277);
nand U2470 (N_2470,In_422,N_1406);
nand U2471 (N_2471,N_1366,In_4629);
nor U2472 (N_2472,In_3043,In_3957);
nand U2473 (N_2473,N_629,In_4503);
nor U2474 (N_2474,N_153,N_1781);
or U2475 (N_2475,In_179,In_3920);
and U2476 (N_2476,N_481,N_695);
and U2477 (N_2477,In_1999,N_126);
nand U2478 (N_2478,N_37,N_64);
nand U2479 (N_2479,In_2406,N_138);
and U2480 (N_2480,N_70,N_253);
nor U2481 (N_2481,N_1147,N_1235);
nand U2482 (N_2482,N_1510,In_4540);
and U2483 (N_2483,In_2407,N_1153);
nand U2484 (N_2484,In_4738,N_1568);
or U2485 (N_2485,N_284,In_3345);
nand U2486 (N_2486,N_71,N_538);
xnor U2487 (N_2487,In_2850,In_1386);
xor U2488 (N_2488,In_2827,N_1987);
or U2489 (N_2489,N_359,N_1869);
nand U2490 (N_2490,N_1475,N_475);
nand U2491 (N_2491,N_797,In_3114);
or U2492 (N_2492,In_456,N_1463);
xnor U2493 (N_2493,In_2911,In_3242);
nor U2494 (N_2494,N_944,In_3472);
nand U2495 (N_2495,In_4453,N_374);
and U2496 (N_2496,N_1670,N_201);
nand U2497 (N_2497,N_281,N_1687);
nor U2498 (N_2498,N_1759,N_878);
nor U2499 (N_2499,N_222,In_1487);
nand U2500 (N_2500,In_4305,N_1448);
or U2501 (N_2501,N_717,N_1236);
or U2502 (N_2502,N_24,N_1113);
or U2503 (N_2503,N_1402,N_341);
or U2504 (N_2504,In_450,N_443);
nand U2505 (N_2505,N_243,In_3414);
and U2506 (N_2506,In_3415,N_378);
or U2507 (N_2507,In_930,N_1867);
xnor U2508 (N_2508,N_399,N_79);
nor U2509 (N_2509,N_1431,N_293);
xnor U2510 (N_2510,N_906,N_1311);
xor U2511 (N_2511,N_382,N_1939);
or U2512 (N_2512,In_3201,In_2433);
and U2513 (N_2513,In_4157,N_518);
xor U2514 (N_2514,N_498,N_755);
and U2515 (N_2515,In_4114,N_1943);
and U2516 (N_2516,N_825,N_1999);
nand U2517 (N_2517,N_1806,N_1611);
nor U2518 (N_2518,N_652,N_80);
or U2519 (N_2519,In_259,In_2343);
and U2520 (N_2520,In_2555,In_1402);
nor U2521 (N_2521,In_454,In_4852);
or U2522 (N_2522,N_393,N_45);
xnor U2523 (N_2523,In_2093,N_316);
or U2524 (N_2524,N_1192,N_1704);
xor U2525 (N_2525,In_4232,N_894);
xor U2526 (N_2526,N_1403,N_934);
nor U2527 (N_2527,In_2899,N_408);
nand U2528 (N_2528,N_524,N_477);
and U2529 (N_2529,N_590,N_684);
nand U2530 (N_2530,N_782,In_4497);
xor U2531 (N_2531,In_3832,N_1169);
and U2532 (N_2532,N_905,N_1218);
or U2533 (N_2533,In_1039,N_89);
nor U2534 (N_2534,In_1113,N_240);
nor U2535 (N_2535,N_1174,N_1619);
or U2536 (N_2536,In_192,N_1549);
and U2537 (N_2537,N_1490,In_3229);
nand U2538 (N_2538,N_1525,N_1618);
nor U2539 (N_2539,N_1069,N_380);
xnor U2540 (N_2540,N_904,N_1814);
nand U2541 (N_2541,In_1701,N_885);
xor U2542 (N_2542,N_618,In_1399);
nand U2543 (N_2543,N_1310,N_1551);
nand U2544 (N_2544,In_3480,In_2183);
xor U2545 (N_2545,N_960,In_3387);
nand U2546 (N_2546,In_206,In_1862);
or U2547 (N_2547,In_288,In_630);
or U2548 (N_2548,In_1665,N_1859);
xnor U2549 (N_2549,N_1338,N_907);
nor U2550 (N_2550,N_453,N_29);
nand U2551 (N_2551,N_764,N_1055);
nor U2552 (N_2552,N_1691,N_1377);
xnor U2553 (N_2553,N_1303,In_1172);
xor U2554 (N_2554,N_1271,N_686);
or U2555 (N_2555,N_1194,In_3255);
nand U2556 (N_2556,N_1813,N_441);
and U2557 (N_2557,N_1700,N_1553);
nand U2558 (N_2558,N_884,N_324);
or U2559 (N_2559,In_388,N_1784);
nor U2560 (N_2560,In_4036,N_1418);
and U2561 (N_2561,N_47,N_433);
and U2562 (N_2562,In_173,N_1410);
xor U2563 (N_2563,N_41,In_1640);
or U2564 (N_2564,N_1476,N_768);
xnor U2565 (N_2565,N_1247,N_985);
nor U2566 (N_2566,In_4019,N_75);
and U2567 (N_2567,N_910,In_118);
xor U2568 (N_2568,N_1602,In_3446);
xnor U2569 (N_2569,In_774,In_2094);
nor U2570 (N_2570,N_593,N_1931);
xor U2571 (N_2571,N_1161,In_2102);
or U2572 (N_2572,N_1550,In_684);
nor U2573 (N_2573,N_159,N_891);
nor U2574 (N_2574,In_1349,In_1026);
nor U2575 (N_2575,In_1544,N_25);
or U2576 (N_2576,In_3190,N_17);
xnor U2577 (N_2577,N_941,In_4068);
or U2578 (N_2578,N_1455,N_942);
nand U2579 (N_2579,N_375,N_445);
and U2580 (N_2580,N_571,In_61);
xnor U2581 (N_2581,N_752,N_1775);
or U2582 (N_2582,N_1731,N_1500);
and U2583 (N_2583,In_1495,N_1084);
xnor U2584 (N_2584,N_1154,N_1726);
nand U2585 (N_2585,In_597,N_582);
and U2586 (N_2586,N_1979,In_3314);
xor U2587 (N_2587,N_1569,In_1604);
nor U2588 (N_2588,In_2201,In_4618);
xor U2589 (N_2589,N_303,N_1646);
nor U2590 (N_2590,N_1186,N_607);
and U2591 (N_2591,N_961,In_3679);
nand U2592 (N_2592,N_300,In_2079);
or U2593 (N_2593,In_1142,N_1287);
or U2594 (N_2594,In_4499,N_1629);
nor U2595 (N_2595,N_1969,N_986);
or U2596 (N_2596,N_232,N_1076);
and U2597 (N_2597,N_1890,N_803);
nor U2598 (N_2598,N_1085,N_777);
nor U2599 (N_2599,In_2764,N_335);
and U2600 (N_2600,N_623,N_903);
nor U2601 (N_2601,N_1284,N_603);
xnor U2602 (N_2602,In_3503,In_1646);
nor U2603 (N_2603,In_2512,N_1489);
nor U2604 (N_2604,In_4158,N_82);
nor U2605 (N_2605,N_137,In_2068);
and U2606 (N_2606,N_998,N_1100);
nor U2607 (N_2607,N_1272,N_1561);
nor U2608 (N_2608,In_3551,N_728);
or U2609 (N_2609,In_4972,In_2563);
and U2610 (N_2610,In_397,N_1156);
and U2611 (N_2611,In_4998,In_1841);
and U2612 (N_2612,In_2412,N_1382);
xnor U2613 (N_2613,N_1607,In_3748);
nand U2614 (N_2614,In_1683,N_1899);
or U2615 (N_2615,N_164,In_3729);
nand U2616 (N_2616,N_822,N_542);
nand U2617 (N_2617,N_373,N_982);
and U2618 (N_2618,N_1600,N_1820);
and U2619 (N_2619,N_457,N_1267);
and U2620 (N_2620,N_1738,In_653);
xor U2621 (N_2621,In_4936,In_3913);
nand U2622 (N_2622,N_1152,In_128);
or U2623 (N_2623,N_1892,In_691);
nor U2624 (N_2624,N_1648,N_829);
xnor U2625 (N_2625,In_1541,N_548);
nand U2626 (N_2626,In_966,N_594);
nand U2627 (N_2627,N_808,N_835);
nor U2628 (N_2628,In_3406,N_1198);
or U2629 (N_2629,N_1502,N_245);
nor U2630 (N_2630,N_241,N_463);
xor U2631 (N_2631,In_2180,N_689);
and U2632 (N_2632,In_3191,N_705);
or U2633 (N_2633,N_774,N_1449);
xnor U2634 (N_2634,N_92,In_4006);
xnor U2635 (N_2635,N_1797,In_204);
xnor U2636 (N_2636,N_779,In_3798);
nor U2637 (N_2637,N_1000,N_1885);
nor U2638 (N_2638,N_340,N_605);
xnor U2639 (N_2639,N_662,N_1013);
or U2640 (N_2640,N_608,In_4547);
and U2641 (N_2641,In_1697,N_124);
xor U2642 (N_2642,In_4630,N_1344);
and U2643 (N_2643,N_1745,In_4661);
or U2644 (N_2644,In_3777,In_1607);
nand U2645 (N_2645,N_1603,In_385);
nor U2646 (N_2646,N_1269,N_1009);
and U2647 (N_2647,N_466,N_628);
xor U2648 (N_2648,In_3391,N_1790);
xor U2649 (N_2649,N_1388,In_3822);
and U2650 (N_2650,In_444,In_2279);
or U2651 (N_2651,N_588,In_4343);
nand U2652 (N_2652,In_3618,In_4117);
nand U2653 (N_2653,In_1831,N_263);
and U2654 (N_2654,N_616,N_402);
nand U2655 (N_2655,N_615,N_1826);
xnor U2656 (N_2656,N_1654,N_981);
nand U2657 (N_2657,In_1806,In_4254);
and U2658 (N_2658,N_993,N_1636);
xnor U2659 (N_2659,N_330,In_2288);
and U2660 (N_2660,In_3553,In_3045);
or U2661 (N_2661,In_3318,N_1032);
or U2662 (N_2662,N_182,N_1518);
xor U2663 (N_2663,N_1514,N_1316);
or U2664 (N_2664,In_43,N_1990);
nand U2665 (N_2665,N_889,N_1045);
xnor U2666 (N_2666,In_1268,In_3050);
nand U2667 (N_2667,In_4703,N_1717);
xnor U2668 (N_2668,In_3434,N_682);
and U2669 (N_2669,In_3536,N_1541);
nand U2670 (N_2670,In_3865,N_1794);
and U2671 (N_2671,N_254,N_1276);
xor U2672 (N_2672,N_1836,N_437);
xor U2673 (N_2673,N_1755,N_746);
nor U2674 (N_2674,In_1929,In_4925);
nor U2675 (N_2675,N_1461,N_1047);
xor U2676 (N_2676,In_2895,N_1595);
and U2677 (N_2677,N_516,In_4822);
or U2678 (N_2678,In_3090,N_1373);
or U2679 (N_2679,N_1913,N_1021);
and U2680 (N_2680,N_1737,N_1997);
and U2681 (N_2681,In_2430,In_2200);
and U2682 (N_2682,N_1912,N_1723);
and U2683 (N_2683,N_1963,In_3072);
and U2684 (N_2684,In_1225,N_1875);
nor U2685 (N_2685,N_84,N_703);
and U2686 (N_2686,N_1579,N_1353);
nor U2687 (N_2687,N_1973,N_1872);
xor U2688 (N_2688,N_1308,N_643);
xnor U2689 (N_2689,In_2342,In_2862);
xor U2690 (N_2690,N_1078,N_480);
xnor U2691 (N_2691,N_1309,N_1891);
nand U2692 (N_2692,N_34,N_937);
nor U2693 (N_2693,N_488,N_1002);
xnor U2694 (N_2694,N_828,N_1178);
and U2695 (N_2695,N_637,N_452);
and U2696 (N_2696,N_1846,In_2338);
xor U2697 (N_2697,In_3505,In_2132);
and U2698 (N_2698,N_121,In_2655);
xnor U2699 (N_2699,In_4792,N_840);
nand U2700 (N_2700,N_1799,N_1429);
and U2701 (N_2701,N_388,In_273);
nand U2702 (N_2702,In_3403,In_2526);
nor U2703 (N_2703,In_3888,N_1395);
nor U2704 (N_2704,N_595,N_181);
nor U2705 (N_2705,N_1829,N_412);
or U2706 (N_2706,In_4788,In_2590);
nor U2707 (N_2707,N_1536,In_2669);
nor U2708 (N_2708,N_1428,N_19);
xnor U2709 (N_2709,N_533,N_509);
xor U2710 (N_2710,N_1471,N_1432);
or U2711 (N_2711,In_4918,In_1482);
or U2712 (N_2712,N_461,In_4761);
or U2713 (N_2713,N_556,N_123);
and U2714 (N_2714,In_2328,N_1176);
nand U2715 (N_2715,N_1570,N_503);
and U2716 (N_2716,N_1193,N_879);
xor U2717 (N_2717,N_694,N_1606);
or U2718 (N_2718,N_309,N_1230);
and U2719 (N_2719,N_640,N_1212);
nand U2720 (N_2720,N_383,N_398);
nor U2721 (N_2721,N_744,In_2956);
nor U2722 (N_2722,N_552,N_809);
nand U2723 (N_2723,N_1098,N_558);
and U2724 (N_2724,In_3951,N_1505);
and U2725 (N_2725,N_553,In_3332);
xor U2726 (N_2726,N_922,N_731);
nor U2727 (N_2727,N_954,N_1980);
nor U2728 (N_2728,N_1998,N_1874);
or U2729 (N_2729,N_389,N_105);
or U2730 (N_2730,N_1721,In_748);
nand U2731 (N_2731,In_2635,N_1120);
nor U2732 (N_2732,In_2708,In_1933);
and U2733 (N_2733,In_1900,N_267);
and U2734 (N_2734,N_776,N_923);
and U2735 (N_2735,N_1727,N_860);
xnor U2736 (N_2736,N_118,In_1036);
or U2737 (N_2737,N_969,N_1898);
nor U2738 (N_2738,N_735,N_1616);
and U2739 (N_2739,N_1234,In_154);
and U2740 (N_2740,In_3284,In_4586);
or U2741 (N_2741,N_116,N_530);
nor U2742 (N_2742,N_1261,In_1731);
nor U2743 (N_2743,N_1828,N_251);
or U2744 (N_2744,N_535,N_1925);
nor U2745 (N_2745,N_1904,In_880);
and U2746 (N_2746,In_3259,In_2987);
or U2747 (N_2747,In_3216,In_186);
or U2748 (N_2748,N_332,In_4332);
xor U2749 (N_2749,In_2142,N_1882);
and U2750 (N_2750,N_688,In_1159);
nor U2751 (N_2751,In_1072,N_1756);
nand U2752 (N_2752,In_4334,N_280);
nand U2753 (N_2753,N_1529,In_1493);
nand U2754 (N_2754,N_1004,N_1336);
nor U2755 (N_2755,N_151,N_1533);
and U2756 (N_2756,N_811,In_2443);
nor U2757 (N_2757,N_1811,N_537);
and U2758 (N_2758,N_1389,N_1321);
or U2759 (N_2759,N_1452,N_1592);
or U2760 (N_2760,N_1985,N_1559);
nand U2761 (N_2761,In_2076,N_440);
or U2762 (N_2762,In_1618,N_387);
nand U2763 (N_2763,N_1635,N_1143);
or U2764 (N_2764,N_424,N_208);
nand U2765 (N_2765,N_1083,N_692);
nor U2766 (N_2766,In_603,N_971);
nand U2767 (N_2767,N_701,N_1923);
nor U2768 (N_2768,N_1589,N_366);
and U2769 (N_2769,N_1666,In_4252);
nand U2770 (N_2770,N_837,In_1371);
and U2771 (N_2771,N_1517,N_1394);
xor U2772 (N_2772,In_1699,In_3461);
nor U2773 (N_2773,In_3835,N_890);
xor U2774 (N_2774,N_994,N_298);
and U2775 (N_2775,In_3317,N_1459);
nor U2776 (N_2776,N_1810,In_573);
nand U2777 (N_2777,In_2424,N_56);
nand U2778 (N_2778,In_833,N_104);
nand U2779 (N_2779,N_205,In_3776);
nor U2780 (N_2780,N_439,N_1739);
or U2781 (N_2781,In_2391,In_2131);
nor U2782 (N_2782,N_149,N_868);
nor U2783 (N_2783,N_249,N_285);
and U2784 (N_2784,N_51,N_487);
nor U2785 (N_2785,N_1341,N_1278);
nand U2786 (N_2786,N_1707,In_27);
xnor U2787 (N_2787,N_1906,In_4175);
nand U2788 (N_2788,In_153,In_4315);
xor U2789 (N_2789,In_1833,N_1986);
xor U2790 (N_2790,N_1274,N_133);
nand U2791 (N_2791,In_808,In_3989);
or U2792 (N_2792,N_1188,N_876);
or U2793 (N_2793,In_2768,N_302);
nor U2794 (N_2794,N_1481,N_671);
and U2795 (N_2795,In_1418,N_102);
nand U2796 (N_2796,N_1172,N_66);
nand U2797 (N_2797,In_2516,N_1955);
and U2798 (N_2798,In_3493,N_619);
xnor U2799 (N_2799,In_3276,N_156);
xor U2800 (N_2800,N_979,N_794);
nand U2801 (N_2801,N_796,N_219);
nor U2802 (N_2802,N_1642,N_1961);
xor U2803 (N_2803,N_575,In_3661);
nor U2804 (N_2804,N_384,N_1118);
nand U2805 (N_2805,In_2341,In_1961);
or U2806 (N_2806,In_4711,N_325);
or U2807 (N_2807,N_1848,N_1909);
nor U2808 (N_2808,In_1100,N_1888);
or U2809 (N_2809,N_1134,In_1263);
nand U2810 (N_2810,N_196,In_4709);
xor U2811 (N_2811,N_61,N_675);
nor U2812 (N_2812,In_3799,In_3273);
nor U2813 (N_2813,N_1155,In_3425);
nor U2814 (N_2814,In_245,N_1852);
nand U2815 (N_2815,N_1638,N_125);
nand U2816 (N_2816,N_601,N_586);
nand U2817 (N_2817,N_1695,In_3502);
and U2818 (N_2818,In_4836,In_2025);
nor U2819 (N_2819,In_87,N_1411);
nand U2820 (N_2820,In_4522,N_502);
xnor U2821 (N_2821,N_1300,N_161);
and U2822 (N_2822,N_572,N_1228);
nand U2823 (N_2823,In_2999,In_3065);
or U2824 (N_2824,N_1656,In_2847);
xor U2825 (N_2825,N_1632,In_3143);
nor U2826 (N_2826,N_421,N_154);
nor U2827 (N_2827,In_4638,N_314);
or U2828 (N_2828,N_292,N_162);
nand U2829 (N_2829,In_2222,N_1067);
nand U2830 (N_2830,In_2218,N_44);
nand U2831 (N_2831,N_1102,In_4846);
nand U2832 (N_2832,N_226,N_1472);
or U2833 (N_2833,N_262,N_1757);
nor U2834 (N_2834,In_3905,N_863);
nor U2835 (N_2835,N_1762,In_1217);
nand U2836 (N_2836,In_967,N_1698);
nor U2837 (N_2837,In_139,N_1474);
xor U2838 (N_2838,N_1131,N_235);
nor U2839 (N_2839,In_217,N_1841);
and U2840 (N_2840,N_483,N_1486);
nand U2841 (N_2841,N_428,N_1497);
nand U2842 (N_2842,N_260,N_580);
nand U2843 (N_2843,N_1290,N_1040);
and U2844 (N_2844,In_2084,N_1785);
nor U2845 (N_2845,In_2237,N_816);
nand U2846 (N_2846,N_207,N_983);
and U2847 (N_2847,In_2739,In_4819);
or U2848 (N_2848,N_1531,In_2);
xor U2849 (N_2849,In_2686,N_88);
nor U2850 (N_2850,N_179,N_873);
and U2851 (N_2851,In_4612,N_824);
nor U2852 (N_2852,N_192,In_3181);
or U2853 (N_2853,N_1694,N_881);
and U2854 (N_2854,N_600,N_1231);
nor U2855 (N_2855,In_791,N_959);
and U2856 (N_2856,N_1577,N_1028);
and U2857 (N_2857,N_565,In_4347);
or U2858 (N_2858,In_3167,In_4521);
and U2859 (N_2859,N_193,N_1238);
or U2860 (N_2860,In_2168,N_1296);
xnor U2861 (N_2861,N_1363,N_892);
nand U2862 (N_2862,N_737,In_4569);
nor U2863 (N_2863,In_4421,N_1233);
nor U2864 (N_2864,N_1714,N_988);
nand U2865 (N_2865,N_195,N_1246);
nor U2866 (N_2866,N_1653,In_2472);
xor U2867 (N_2867,N_1044,N_912);
and U2868 (N_2868,In_2336,N_31);
or U2869 (N_2869,N_854,N_925);
or U2870 (N_2870,N_1368,In_3948);
xnor U2871 (N_2871,N_1815,N_1319);
nor U2872 (N_2872,N_28,In_18);
or U2873 (N_2873,N_1735,In_4828);
nand U2874 (N_2874,N_1671,In_681);
and U2875 (N_2875,In_252,In_4224);
xor U2876 (N_2876,N_289,N_203);
nand U2877 (N_2877,N_574,N_827);
xor U2878 (N_2878,N_1805,N_1103);
or U2879 (N_2879,N_1555,N_1950);
nor U2880 (N_2880,In_203,N_1622);
nor U2881 (N_2881,In_2285,N_1408);
or U2882 (N_2882,N_1934,In_1967);
nor U2883 (N_2883,In_935,N_415);
and U2884 (N_2884,N_345,In_4677);
nor U2885 (N_2885,In_2447,N_1501);
nor U2886 (N_2886,N_103,N_1110);
and U2887 (N_2887,N_563,In_4475);
nand U2888 (N_2888,N_1304,N_626);
nand U2889 (N_2889,In_101,N_1574);
or U2890 (N_2890,In_2264,N_1528);
and U2891 (N_2891,N_888,In_2864);
xor U2892 (N_2892,In_4399,In_4339);
xnor U2893 (N_2893,N_396,N_784);
nor U2894 (N_2894,N_482,N_995);
nand U2895 (N_2895,N_1889,N_1038);
nand U2896 (N_2896,N_206,N_1722);
and U2897 (N_2897,N_1732,N_1535);
nand U2898 (N_2898,N_500,N_631);
nand U2899 (N_2899,N_1237,N_78);
or U2900 (N_2900,N_1932,N_1072);
nand U2901 (N_2901,N_745,In_3880);
or U2902 (N_2902,In_1803,N_1293);
nand U2903 (N_2903,N_507,N_1295);
nor U2904 (N_2904,N_1075,In_4930);
or U2905 (N_2905,In_4317,N_625);
or U2906 (N_2906,N_1144,N_1921);
or U2907 (N_2907,N_1202,In_2727);
xnor U2908 (N_2908,N_551,In_929);
or U2909 (N_2909,N_135,N_0);
nand U2910 (N_2910,N_1059,In_4901);
nor U2911 (N_2911,In_132,In_4040);
and U2912 (N_2912,In_3843,N_1342);
nand U2913 (N_2913,N_1544,N_1970);
nand U2914 (N_2914,In_2405,In_3885);
nand U2915 (N_2915,N_620,N_438);
and U2916 (N_2916,N_211,N_1946);
and U2917 (N_2917,In_3923,In_2569);
or U2918 (N_2918,N_560,N_1291);
and U2919 (N_2919,N_921,N_1077);
nor U2920 (N_2920,N_839,N_1444);
xnor U2921 (N_2921,N_1125,N_1097);
xor U2922 (N_2922,In_1670,N_1954);
or U2923 (N_2923,N_1948,N_132);
and U2924 (N_2924,N_999,N_1011);
or U2925 (N_2925,N_591,N_1624);
nor U2926 (N_2926,N_147,In_3418);
nor U2927 (N_2927,In_2652,N_1547);
nor U2928 (N_2928,N_667,N_274);
nor U2929 (N_2929,N_1699,In_1126);
nand U2930 (N_2930,In_1808,N_1114);
xor U2931 (N_2931,N_531,N_987);
xnor U2932 (N_2932,N_992,In_3736);
xor U2933 (N_2933,N_1439,In_1244);
and U2934 (N_2934,N_853,In_1500);
or U2935 (N_2935,N_1823,N_287);
and U2936 (N_2936,N_1029,N_1381);
xor U2937 (N_2937,N_1012,N_1351);
and U2938 (N_2938,N_1584,N_180);
nand U2939 (N_2939,In_2836,N_581);
nor U2940 (N_2940,N_1268,In_2300);
nand U2941 (N_2941,In_3591,N_802);
and U2942 (N_2942,N_1255,N_810);
xor U2943 (N_2943,N_1024,N_1772);
or U2944 (N_2944,N_831,In_4973);
nor U2945 (N_2945,N_624,N_55);
or U2946 (N_2946,N_1119,N_1224);
or U2947 (N_2947,N_1991,In_1209);
and U2948 (N_2948,In_951,N_1750);
or U2949 (N_2949,In_2466,In_650);
nor U2950 (N_2950,In_1463,N_866);
nand U2951 (N_2951,N_1938,In_3183);
nand U2952 (N_2952,N_638,N_691);
nor U2953 (N_2953,N_1673,In_2303);
nor U2954 (N_2954,N_1730,N_353);
and U2955 (N_2955,N_163,N_953);
nand U2956 (N_2956,In_3631,N_318);
and U2957 (N_2957,N_1974,In_671);
xor U2958 (N_2958,N_1214,In_4071);
and U2959 (N_2959,N_724,In_2905);
nand U2960 (N_2960,In_1673,N_120);
nor U2961 (N_2961,In_2848,N_1663);
nand U2962 (N_2962,In_4273,N_1652);
nor U2963 (N_2963,In_789,N_1051);
xnor U2964 (N_2964,N_1868,N_1415);
or U2965 (N_2965,N_1511,N_1260);
nor U2966 (N_2966,N_301,In_2242);
nand U2967 (N_2967,In_2837,N_1286);
or U2968 (N_2968,N_57,In_1473);
nand U2969 (N_2969,N_85,N_1983);
and U2970 (N_2970,N_431,N_1123);
or U2971 (N_2971,In_135,In_1335);
nor U2972 (N_2972,N_1958,N_1933);
nor U2973 (N_2973,In_134,N_1957);
or U2974 (N_2974,In_3687,N_1325);
or U2975 (N_2975,N_1145,In_865);
and U2976 (N_2976,N_32,In_4561);
nor U2977 (N_2977,N_1951,N_704);
and U2978 (N_2978,N_973,N_1496);
nand U2979 (N_2979,N_1400,N_77);
nand U2980 (N_2980,In_1483,N_1655);
xnor U2981 (N_2981,In_1109,In_570);
or U2982 (N_2982,N_1640,N_495);
or U2983 (N_2983,In_764,N_1543);
or U2984 (N_2984,N_1049,N_648);
xnor U2985 (N_2985,In_3408,In_4106);
nor U2986 (N_2986,N_523,In_1914);
or U2987 (N_2987,In_2834,N_3);
nand U2988 (N_2988,N_1035,N_644);
xnor U2989 (N_2989,In_3829,N_806);
xnor U2990 (N_2990,In_1437,N_699);
xor U2991 (N_2991,In_2757,N_872);
nor U2992 (N_2992,N_470,N_351);
and U2993 (N_2993,N_931,N_526);
nor U2994 (N_2994,N_602,In_3915);
nand U2995 (N_2995,N_1248,N_1423);
and U2996 (N_2996,N_1052,N_690);
xor U2997 (N_2997,N_1343,N_842);
or U2998 (N_2998,In_17,N_1710);
nor U2999 (N_2999,In_455,N_1249);
nor U3000 (N_3000,N_1264,N_350);
nand U3001 (N_3001,In_1578,In_2797);
and U3002 (N_3002,N_1916,N_242);
xor U3003 (N_3003,In_100,N_225);
or U3004 (N_3004,In_3753,N_676);
xnor U3005 (N_3005,N_1211,N_210);
xnor U3006 (N_3006,N_1039,In_1145);
nor U3007 (N_3007,In_3509,N_83);
nand U3008 (N_3008,N_1996,N_1108);
or U3009 (N_3009,N_379,N_54);
xor U3010 (N_3010,N_609,In_1973);
nor U3011 (N_3011,N_244,N_1758);
or U3012 (N_3012,N_171,In_4447);
and U3013 (N_3013,N_536,N_525);
nand U3014 (N_3014,In_2897,N_1358);
and U3015 (N_3015,N_199,In_695);
and U3016 (N_3016,N_321,N_404);
and U3017 (N_3017,In_867,N_190);
xnor U3018 (N_3018,In_3021,In_3614);
nor U3019 (N_3019,In_591,N_947);
xor U3020 (N_3020,N_1692,In_2838);
or U3021 (N_3021,N_184,N_911);
or U3022 (N_3022,N_81,N_167);
or U3023 (N_3023,N_1664,N_1480);
and U3024 (N_3024,In_513,N_1822);
nand U3025 (N_3025,N_1426,N_1307);
xnor U3026 (N_3026,N_943,N_508);
nor U3027 (N_3027,N_427,In_4419);
or U3028 (N_3028,In_4556,In_84);
nor U3029 (N_3029,N_972,In_284);
nor U3030 (N_3030,N_1792,In_497);
xor U3031 (N_3031,In_2744,N_522);
nand U3032 (N_3032,N_1657,N_1436);
and U3033 (N_3033,N_397,In_3343);
nor U3034 (N_3034,N_1962,N_1128);
or U3035 (N_3035,In_3146,N_975);
and U3036 (N_3036,N_1397,N_257);
or U3037 (N_3037,In_3003,N_965);
nor U3038 (N_3038,In_4338,In_2557);
nor U3039 (N_3039,N_1598,In_2842);
or U3040 (N_3040,In_4275,N_1749);
xor U3041 (N_3041,N_269,N_1447);
or U3042 (N_3042,In_4456,N_1099);
or U3043 (N_3043,In_162,N_1751);
nor U3044 (N_3044,N_718,N_1747);
or U3045 (N_3045,N_1742,N_1245);
xor U3046 (N_3046,N_1780,N_1807);
or U3047 (N_3047,N_1519,N_464);
nand U3048 (N_3048,N_1205,N_800);
nor U3049 (N_3049,N_547,In_4449);
nand U3050 (N_3050,N_1265,N_569);
nor U3051 (N_3051,N_9,In_2431);
nor U3052 (N_3052,N_1301,N_271);
nor U3053 (N_3053,In_1404,N_1485);
nor U3054 (N_3054,N_1216,N_150);
nor U3055 (N_3055,In_2064,N_423);
or U3056 (N_3056,N_630,N_368);
or U3057 (N_3057,In_2502,N_1643);
and U3058 (N_3058,N_1509,N_1591);
nor U3059 (N_3059,N_1464,N_1335);
and U3060 (N_3060,N_237,N_209);
and U3061 (N_3061,N_1409,N_627);
and U3062 (N_3062,In_4249,N_633);
xor U3063 (N_3063,In_1147,In_3280);
nand U3064 (N_3064,N_1660,In_4696);
or U3065 (N_3065,In_105,In_1546);
and U3066 (N_3066,In_622,N_762);
xnor U3067 (N_3067,N_1947,N_554);
xor U3068 (N_3068,N_753,In_2027);
nor U3069 (N_3069,N_134,In_240);
or U3070 (N_3070,N_1504,N_1056);
xor U3071 (N_3071,In_2252,N_1503);
and U3072 (N_3072,N_887,N_783);
and U3073 (N_3073,N_497,In_1626);
and U3074 (N_3074,N_282,N_1166);
and U3075 (N_3075,In_4034,In_332);
and U3076 (N_3076,In_1162,In_1403);
nand U3077 (N_3077,N_347,N_136);
nor U3078 (N_3078,In_2255,N_1597);
and U3079 (N_3079,N_871,N_436);
nand U3080 (N_3080,In_424,N_36);
nand U3081 (N_3081,N_693,In_21);
nor U3082 (N_3082,N_1132,N_112);
and U3083 (N_3083,N_446,In_2330);
nand U3084 (N_3084,N_410,N_1563);
and U3085 (N_3085,N_579,In_4129);
xor U3086 (N_3086,In_3474,N_933);
or U3087 (N_3087,In_3283,N_798);
or U3088 (N_3088,N_1473,In_4713);
xnor U3089 (N_3089,N_606,N_1421);
nand U3090 (N_3090,In_742,N_945);
nor U3091 (N_3091,In_2823,N_1062);
and U3092 (N_3092,N_1065,N_1001);
xor U3093 (N_3093,N_870,In_1562);
xnor U3094 (N_3094,In_496,N_313);
nand U3095 (N_3095,In_4913,N_1953);
xnor U3096 (N_3096,In_4594,N_1199);
or U3097 (N_3097,In_3164,N_1712);
or U3098 (N_3098,N_1816,N_1088);
xor U3099 (N_3099,In_4898,In_1548);
xnor U3100 (N_3100,N_326,N_451);
xnor U3101 (N_3101,N_1163,N_1645);
nor U3102 (N_3102,N_792,N_805);
nor U3103 (N_3103,N_1405,N_787);
xnor U3104 (N_3104,N_990,N_1346);
and U3105 (N_3105,In_4309,N_176);
nand U3106 (N_3106,In_428,In_2534);
nand U3107 (N_3107,In_4893,N_1944);
or U3108 (N_3108,In_486,N_348);
or U3109 (N_3109,N_559,N_1419);
nor U3110 (N_3110,N_651,N_727);
xnor U3111 (N_3111,N_641,N_272);
nand U3112 (N_3112,In_3532,N_471);
or U3113 (N_3113,N_141,N_1240);
xnor U3114 (N_3114,In_3134,In_1515);
nand U3115 (N_3115,N_1189,In_60);
xor U3116 (N_3116,In_755,N_90);
nor U3117 (N_3117,N_299,In_1598);
nand U3118 (N_3118,N_567,N_1802);
nor U3119 (N_3119,N_1116,In_1486);
nor U3120 (N_3120,In_4637,In_1047);
and U3121 (N_3121,N_407,N_1139);
and U3122 (N_3122,In_533,N_520);
and U3123 (N_3123,In_1127,N_1165);
and U3124 (N_3124,In_4211,N_1357);
or U3125 (N_3125,N_144,N_765);
nand U3126 (N_3126,N_1115,N_390);
nand U3127 (N_3127,In_4011,N_1594);
and U3128 (N_3128,N_1003,In_387);
or U3129 (N_3129,In_3869,N_1995);
or U3130 (N_3130,In_2772,In_4919);
nand U3131 (N_3131,In_3306,N_1006);
xnor U3132 (N_3132,N_1262,N_1708);
xor U3133 (N_3133,In_3716,In_368);
and U3134 (N_3134,N_1711,N_1375);
and U3135 (N_3135,N_145,In_3382);
and U3136 (N_3136,N_1322,In_1937);
nand U3137 (N_3137,In_4996,In_4592);
or U3138 (N_3138,In_1780,N_1734);
and U3139 (N_3139,N_114,N_1430);
and U3140 (N_3140,N_1257,In_4136);
and U3141 (N_3141,N_1935,N_1053);
nor U3142 (N_3142,N_1796,N_1967);
or U3143 (N_3143,N_1917,N_238);
nand U3144 (N_3144,N_1080,N_1289);
nand U3145 (N_3145,In_4572,N_218);
and U3146 (N_3146,N_1818,In_3738);
and U3147 (N_3147,N_1649,N_775);
xor U3148 (N_3148,N_781,N_1614);
or U3149 (N_3149,N_493,N_1539);
nor U3150 (N_3150,N_1488,N_227);
nor U3151 (N_3151,N_950,In_1583);
and U3152 (N_3152,N_1530,In_1433);
nand U3153 (N_3153,In_3863,N_1905);
xnor U3154 (N_3154,In_301,N_12);
nand U3155 (N_3155,N_672,In_4115);
or U3156 (N_3156,N_1438,In_554);
and U3157 (N_3157,N_939,In_3730);
nand U3158 (N_3158,In_3933,N_650);
and U3159 (N_3159,N_1928,In_4633);
nand U3160 (N_3160,N_360,In_4057);
and U3161 (N_3161,N_1479,In_1307);
or U3162 (N_3162,N_1680,N_1227);
nand U3163 (N_3163,N_1399,In_340);
xnor U3164 (N_3164,N_320,In_3615);
and U3165 (N_3165,N_277,N_1225);
and U3166 (N_3166,In_2138,N_527);
and U3167 (N_3167,N_756,In_3312);
or U3168 (N_3168,N_517,In_165);
nand U3169 (N_3169,N_268,N_1170);
xor U3170 (N_3170,In_3248,N_1675);
nand U3171 (N_3171,N_1367,N_1929);
or U3172 (N_3172,N_68,N_1837);
nand U3173 (N_3173,In_247,N_1557);
nand U3174 (N_3174,In_4751,In_406);
nand U3175 (N_3175,N_248,N_1195);
nor U3176 (N_3176,N_1768,N_1064);
and U3177 (N_3177,N_1288,N_678);
nand U3178 (N_3178,In_1747,N_455);
nor U3179 (N_3179,N_1355,In_11);
xor U3180 (N_3180,In_462,N_1106);
or U3181 (N_3181,N_723,N_935);
xor U3182 (N_3182,N_930,N_570);
nor U3183 (N_3183,N_1456,In_3970);
nor U3184 (N_3184,In_4715,In_4810);
nand U3185 (N_3185,N_1516,N_578);
and U3186 (N_3186,N_926,N_1387);
nor U3187 (N_3187,In_914,In_2898);
nor U3188 (N_3188,In_504,N_962);
nand U3189 (N_3189,N_1924,In_2370);
and U3190 (N_3190,N_1175,N_152);
and U3191 (N_3191,N_1879,N_669);
nand U3192 (N_3192,In_1182,N_758);
xor U3193 (N_3193,In_1325,N_319);
nand U3194 (N_3194,In_2931,N_1819);
nand U3195 (N_3195,N_1787,In_1037);
xnor U3196 (N_3196,N_754,In_718);
xor U3197 (N_3197,N_1242,In_3715);
and U3198 (N_3198,N_1371,In_215);
xnor U3199 (N_3199,N_165,N_1015);
nor U3200 (N_3200,N_1588,N_820);
nand U3201 (N_3201,N_204,In_545);
nand U3202 (N_3202,N_371,N_951);
or U3203 (N_3203,N_479,In_4328);
nor U3204 (N_3204,N_1266,N_465);
and U3205 (N_3205,In_3122,In_2226);
xnor U3206 (N_3206,In_2611,N_416);
nand U3207 (N_3207,In_1874,N_2);
nor U3208 (N_3208,In_3692,N_228);
nand U3209 (N_3209,N_751,In_1003);
and U3210 (N_3210,N_1253,In_4720);
nor U3211 (N_3211,N_460,N_1703);
or U3212 (N_3212,In_965,N_967);
xnor U3213 (N_3213,N_212,N_1070);
xor U3214 (N_3214,In_4505,N_949);
nor U3215 (N_3215,N_364,In_112);
and U3216 (N_3216,N_1965,In_323);
xnor U3217 (N_3217,In_1065,N_1086);
nor U3218 (N_3218,N_432,N_1585);
nor U3219 (N_3219,In_185,N_821);
nor U3220 (N_3220,N_1285,N_110);
nor U3221 (N_3221,In_4440,N_1482);
nor U3222 (N_3222,In_799,In_1919);
nand U3223 (N_3223,N_213,N_773);
nor U3224 (N_3224,N_86,N_1808);
and U3225 (N_3225,N_1861,In_595);
xor U3226 (N_3226,In_2065,N_1337);
or U3227 (N_3227,In_3696,N_505);
nand U3228 (N_3228,N_539,N_392);
xor U3229 (N_3229,N_867,In_3057);
or U3230 (N_3230,In_1491,N_733);
nor U3231 (N_3231,N_1789,N_916);
nor U3232 (N_3232,N_869,N_231);
and U3233 (N_3233,In_1066,N_1507);
xor U3234 (N_3234,In_4714,N_1856);
nor U3235 (N_3235,In_2126,In_3401);
or U3236 (N_3236,N_617,N_826);
nand U3237 (N_3237,N_1821,N_312);
or U3238 (N_3238,In_4080,N_448);
or U3239 (N_3239,N_709,N_400);
and U3240 (N_3240,N_233,N_200);
or U3241 (N_3241,N_42,N_924);
xnor U3242 (N_3242,N_1313,N_738);
nor U3243 (N_3243,N_1964,In_4417);
or U3244 (N_3244,N_899,In_3668);
nor U3245 (N_3245,In_51,N_1201);
and U3246 (N_3246,In_256,In_4623);
xnor U3247 (N_3247,N_984,N_874);
and U3248 (N_3248,N_276,In_4140);
xor U3249 (N_3249,N_772,N_766);
xor U3250 (N_3250,In_3398,N_46);
and U3251 (N_3251,N_1446,N_936);
and U3252 (N_3252,In_1971,N_1223);
nor U3253 (N_3253,N_188,In_1134);
or U3254 (N_3254,N_1677,In_655);
nand U3255 (N_3255,In_547,In_235);
and U3256 (N_3256,N_1451,In_3197);
or U3257 (N_3257,In_4917,In_818);
nand U3258 (N_3258,In_4265,In_3858);
or U3259 (N_3259,In_2995,In_4486);
or U3260 (N_3260,N_456,N_647);
xor U3261 (N_3261,N_583,N_413);
nor U3262 (N_3262,In_3719,N_1862);
and U3263 (N_3263,N_372,In_1677);
and U3264 (N_3264,N_976,N_989);
or U3265 (N_3265,N_1434,N_1776);
nand U3266 (N_3266,N_1066,N_91);
nand U3267 (N_3267,N_113,N_1159);
xnor U3268 (N_3268,In_4390,N_900);
and U3269 (N_3269,In_2663,N_173);
xnor U3270 (N_3270,In_4736,N_401);
or U3271 (N_3271,In_4833,In_4851);
xnor U3272 (N_3272,N_1349,N_221);
xnor U3273 (N_3273,In_4746,In_2386);
or U3274 (N_3274,N_1546,In_1897);
xnor U3275 (N_3275,N_1752,N_1417);
nor U3276 (N_3276,N_174,In_1822);
nand U3277 (N_3277,In_4111,In_1357);
nand U3278 (N_3278,N_1041,N_266);
or U3279 (N_3279,In_4279,N_977);
nor U3280 (N_3280,In_2191,In_3135);
nor U3281 (N_3281,N_194,In_2725);
or U3282 (N_3282,N_1870,N_1146);
and U3283 (N_3283,N_1803,N_1180);
or U3284 (N_3284,N_722,N_69);
nand U3285 (N_3285,In_1319,N_467);
nor U3286 (N_3286,N_1037,N_333);
and U3287 (N_3287,N_1683,N_666);
or U3288 (N_3288,N_1741,In_1457);
nor U3289 (N_3289,In_2276,N_685);
and U3290 (N_3290,In_4582,N_813);
nor U3291 (N_3291,N_1241,N_30);
nor U3292 (N_3292,N_1196,N_741);
nand U3293 (N_3293,In_2456,In_231);
or U3294 (N_3294,N_1493,N_1018);
and U3295 (N_3295,In_1320,N_747);
nor U3296 (N_3296,N_711,In_3170);
xor U3297 (N_3297,In_4483,N_716);
nor U3298 (N_3298,N_1779,N_1556);
nand U3299 (N_3299,In_511,N_1689);
nand U3300 (N_3300,In_2275,In_1358);
and U3301 (N_3301,In_1873,N_1748);
nand U3302 (N_3302,N_952,N_614);
or U3303 (N_3303,N_489,N_763);
nand U3304 (N_3304,N_1127,N_712);
or U3305 (N_3305,N_1552,N_1831);
nor U3306 (N_3306,N_736,N_1520);
nor U3307 (N_3307,In_438,In_1882);
xor U3308 (N_3308,N_1720,N_224);
nor U3309 (N_3309,N_72,N_1613);
nor U3310 (N_3310,N_1782,N_169);
nor U3311 (N_3311,N_968,In_212);
or U3312 (N_3312,N_1764,N_830);
xnor U3313 (N_3313,In_1062,N_1952);
nor U3314 (N_3314,In_4294,N_1104);
nor U3315 (N_3315,In_906,N_1770);
nand U3316 (N_3316,N_434,In_311);
xor U3317 (N_3317,In_4139,In_225);
xor U3318 (N_3318,N_1385,N_189);
and U3319 (N_3319,N_343,N_1437);
nor U3320 (N_3320,N_444,N_1217);
nand U3321 (N_3321,N_1095,N_1918);
nand U3322 (N_3322,In_3416,In_407);
nor U3323 (N_3323,In_4744,N_1783);
or U3324 (N_3324,In_1612,N_367);
xor U3325 (N_3325,N_39,In_4133);
nand U3326 (N_3326,N_1101,In_3665);
xnor U3327 (N_3327,N_1661,N_1679);
or U3328 (N_3328,N_1865,N_948);
nand U3329 (N_3329,In_1236,N_1239);
nor U3330 (N_3330,In_4700,N_970);
nand U3331 (N_3331,In_3037,N_843);
nor U3332 (N_3332,In_2414,N_1761);
and U3333 (N_3333,N_1140,In_12);
or U3334 (N_3334,N_8,In_788);
nor U3335 (N_3335,N_18,In_4849);
nor U3336 (N_3336,N_250,N_1725);
and U3337 (N_3337,N_311,N_76);
and U3338 (N_3338,N_815,N_101);
nand U3339 (N_3339,In_3286,In_3497);
and U3340 (N_3340,N_1545,N_1259);
nand U3341 (N_3341,N_789,N_748);
nand U3342 (N_3342,In_2645,N_216);
nand U3343 (N_3343,N_1327,In_3066);
nand U3344 (N_3344,N_1884,N_732);
or U3345 (N_3345,In_3365,N_1709);
nand U3346 (N_3346,In_1279,N_429);
nor U3347 (N_3347,N_278,N_902);
or U3348 (N_3348,N_1498,N_1554);
xnor U3349 (N_3349,In_1315,N_956);
nor U3350 (N_3350,N_1850,N_1082);
nand U3351 (N_3351,N_265,In_1020);
nand U3352 (N_3352,N_680,N_1801);
and U3353 (N_3353,N_1079,N_346);
or U3354 (N_3354,N_597,N_1937);
nand U3355 (N_3355,In_1526,N_1631);
nand U3356 (N_3356,N_1919,N_1333);
xnor U3357 (N_3357,In_2537,In_2193);
nand U3358 (N_3358,N_98,N_1669);
or U3359 (N_3359,N_1537,In_4614);
and U3360 (N_3360,In_525,N_679);
nand U3361 (N_3361,In_2874,In_1524);
xnor U3362 (N_3362,In_4222,In_3766);
xor U3363 (N_3363,N_496,N_1279);
and U3364 (N_3364,N_13,N_1157);
and U3365 (N_3365,In_213,In_2488);
and U3366 (N_3366,N_743,N_1978);
or U3367 (N_3367,In_1297,N_883);
xor U3368 (N_3368,N_1910,In_214);
nand U3369 (N_3369,N_1390,N_1678);
nor U3370 (N_3370,In_3795,N_499);
nand U3371 (N_3371,In_2223,N_1094);
or U3372 (N_3372,N_529,N_996);
or U3373 (N_3373,N_770,In_3089);
xnor U3374 (N_3374,In_3071,N_117);
and U3375 (N_3375,N_604,N_1696);
nor U3376 (N_3376,In_4598,N_336);
nand U3377 (N_3377,In_1055,In_2514);
nand U3378 (N_3378,In_3002,N_914);
xnor U3379 (N_3379,N_1515,N_856);
or U3380 (N_3380,In_1782,N_1701);
xor U3381 (N_3381,In_452,N_1433);
xnor U3382 (N_3382,N_549,N_1864);
or U3383 (N_3383,N_1760,N_875);
or U3384 (N_3384,N_4,N_599);
and U3385 (N_3385,N_929,N_49);
or U3386 (N_3386,N_918,N_229);
xnor U3387 (N_3387,In_3266,In_2794);
or U3388 (N_3388,N_940,N_636);
xnor U3389 (N_3389,In_2401,N_1054);
or U3390 (N_3390,In_2733,N_1184);
nand U3391 (N_3391,In_1447,In_392);
xor U3392 (N_3392,In_453,In_599);
xnor U3393 (N_3393,N_185,N_1729);
nor U3394 (N_3394,N_1587,N_1477);
or U3395 (N_3395,N_564,N_698);
and U3396 (N_3396,N_848,In_4033);
nor U3397 (N_3397,N_857,N_256);
xor U3398 (N_3398,N_259,In_756);
and U3399 (N_3399,N_713,N_469);
or U3400 (N_3400,N_919,In_2124);
nand U3401 (N_3401,N_759,N_1016);
xnor U3402 (N_3402,N_1527,N_486);
xnor U3403 (N_3403,In_3328,N_801);
and U3404 (N_3404,N_761,N_1258);
and U3405 (N_3405,In_1480,N_1630);
nand U3406 (N_3406,N_849,N_1562);
xor U3407 (N_3407,N_1994,N_1364);
xnor U3408 (N_3408,N_1512,N_1684);
nand U3409 (N_3409,N_858,In_3097);
nand U3410 (N_3410,In_2305,N_1424);
or U3411 (N_3411,In_372,In_2580);
nand U3412 (N_3412,N_1036,In_587);
or U3413 (N_3413,N_674,N_1930);
and U3414 (N_3414,N_1275,In_2011);
or U3415 (N_3415,N_1014,N_823);
or U3416 (N_3416,In_2054,N_1033);
or U3417 (N_3417,N_306,In_4452);
and U3418 (N_3418,N_1662,N_119);
and U3419 (N_3419,N_946,N_146);
nor U3420 (N_3420,N_1200,N_1483);
nor U3421 (N_3421,In_246,N_286);
or U3422 (N_3422,In_4410,N_1830);
nand U3423 (N_3423,N_1362,N_920);
nand U3424 (N_3424,In_4812,N_1221);
xnor U3425 (N_3425,N_355,N_834);
xor U3426 (N_3426,In_2123,N_1847);
nand U3427 (N_3427,In_4414,N_510);
xnor U3428 (N_3428,N_814,N_1111);
nor U3429 (N_3429,N_100,N_1866);
nor U3430 (N_3430,N_63,N_1329);
or U3431 (N_3431,In_3054,In_1112);
nor U3432 (N_3432,N_710,N_1126);
nor U3433 (N_3433,In_3793,N_658);
nand U3434 (N_3434,N_1845,N_1767);
nor U3435 (N_3435,N_707,In_1090);
nor U3436 (N_3436,N_665,In_1243);
xor U3437 (N_3437,In_1692,N_1454);
xnor U3438 (N_3438,N_1508,N_1007);
or U3439 (N_3439,In_3595,N_1282);
nor U3440 (N_3440,N_1320,N_1878);
nor U3441 (N_3441,In_1622,N_1765);
and U3442 (N_3442,N_381,In_1060);
nand U3443 (N_3443,N_1407,In_2074);
nand U3444 (N_3444,N_1942,N_1297);
nand U3445 (N_3445,N_1129,N_573);
nand U3446 (N_3446,N_1352,N_202);
xor U3447 (N_3447,N_155,N_576);
nor U3448 (N_3448,In_4056,N_1702);
xor U3449 (N_3449,N_1839,N_719);
or U3450 (N_3450,In_2349,In_4498);
nand U3451 (N_3451,N_1940,N_297);
and U3452 (N_3452,In_3428,In_119);
and U3453 (N_3453,N_1190,N_1774);
xnor U3454 (N_3454,In_3322,N_1305);
nand U3455 (N_3455,In_4658,In_1199);
or U3456 (N_3456,N_356,N_305);
nor U3457 (N_3457,N_275,N_1927);
xor U3458 (N_3458,N_1676,N_1314);
and U3459 (N_3459,In_682,In_523);
and U3460 (N_3460,In_4459,In_3545);
nor U3461 (N_3461,N_122,In_4004);
and U3462 (N_3462,N_1294,N_1506);
xnor U3463 (N_3463,N_317,N_1465);
and U3464 (N_3464,In_3101,In_2734);
nor U3465 (N_3465,N_1605,In_91);
and U3466 (N_3466,N_1093,N_622);
xnor U3467 (N_3467,In_3223,N_478);
and U3468 (N_3468,N_1769,N_323);
nand U3469 (N_3469,In_405,N_1838);
and U3470 (N_3470,N_739,N_791);
nand U3471 (N_3471,N_217,N_577);
nand U3472 (N_3472,N_1853,N_1492);
nand U3473 (N_3473,In_933,N_861);
and U3474 (N_3474,N_170,N_657);
or U3475 (N_3475,N_462,N_1376);
nor U3476 (N_3476,N_706,N_1532);
nor U3477 (N_3477,N_1413,N_1604);
or U3478 (N_3478,N_1229,N_1736);
xnor U3479 (N_3479,N_864,N_1977);
or U3480 (N_3480,N_1468,N_473);
xnor U3481 (N_3481,N_1746,N_729);
nand U3482 (N_3482,N_653,In_1735);
xnor U3483 (N_3483,In_191,N_655);
nor U3484 (N_3484,N_882,N_1331);
nor U3485 (N_3485,In_2272,N_1185);
nor U3486 (N_3486,In_698,In_4797);
nor U3487 (N_3487,N_283,N_1893);
nor U3488 (N_3488,N_1754,In_3683);
or U3489 (N_3489,N_1763,N_187);
nor U3490 (N_3490,N_730,N_1250);
or U3491 (N_3491,N_1491,In_4131);
and U3492 (N_3492,N_1306,In_3751);
xnor U3493 (N_3493,N_38,N_1232);
xor U3494 (N_3494,N_1715,N_157);
nor U3495 (N_3495,N_261,In_1917);
nor U3496 (N_3496,N_6,N_459);
or U3497 (N_3497,In_2289,N_978);
nor U3498 (N_3498,In_1739,N_1374);
nor U3499 (N_3499,N_1487,N_1945);
nor U3500 (N_3500,N_166,In_2727);
and U3501 (N_3501,N_46,In_74);
or U3502 (N_3502,In_3122,N_585);
nor U3503 (N_3503,N_1781,N_1104);
and U3504 (N_3504,N_418,N_1527);
nor U3505 (N_3505,N_1864,In_4453);
or U3506 (N_3506,N_660,In_1402);
xor U3507 (N_3507,N_1695,N_1332);
and U3508 (N_3508,In_4459,N_1018);
or U3509 (N_3509,N_662,In_1548);
or U3510 (N_3510,N_933,In_1262);
and U3511 (N_3511,N_827,In_11);
nor U3512 (N_3512,N_1246,N_1717);
nand U3513 (N_3513,N_422,N_79);
xnor U3514 (N_3514,N_1857,N_1536);
nand U3515 (N_3515,In_100,N_1115);
xnor U3516 (N_3516,In_2330,N_1282);
xnor U3517 (N_3517,N_1740,N_933);
and U3518 (N_3518,N_737,N_404);
nand U3519 (N_3519,N_875,In_3122);
nand U3520 (N_3520,In_589,In_1047);
nand U3521 (N_3521,N_98,N_716);
nor U3522 (N_3522,N_812,N_1046);
nand U3523 (N_3523,N_1100,N_213);
nor U3524 (N_3524,N_356,In_2534);
nor U3525 (N_3525,In_3191,N_1307);
nand U3526 (N_3526,In_2407,N_1334);
nand U3527 (N_3527,N_1063,N_1717);
nand U3528 (N_3528,In_3480,N_1676);
and U3529 (N_3529,N_1310,N_1960);
nor U3530 (N_3530,N_149,N_446);
and U3531 (N_3531,In_84,N_224);
xor U3532 (N_3532,N_195,N_1346);
and U3533 (N_3533,N_247,In_2742);
nand U3534 (N_3534,In_4612,In_1873);
and U3535 (N_3535,N_729,N_1537);
and U3536 (N_3536,In_2684,N_382);
and U3537 (N_3537,In_3461,N_1950);
nor U3538 (N_3538,N_850,N_1373);
and U3539 (N_3539,N_1109,N_107);
xnor U3540 (N_3540,N_649,N_1367);
or U3541 (N_3541,In_2974,N_247);
or U3542 (N_3542,N_594,N_617);
xor U3543 (N_3543,N_503,N_302);
xnor U3544 (N_3544,N_980,N_914);
or U3545 (N_3545,N_1350,N_1492);
nor U3546 (N_3546,N_56,In_486);
nand U3547 (N_3547,N_466,N_93);
xor U3548 (N_3548,In_1548,N_377);
nor U3549 (N_3549,N_1400,N_139);
xor U3550 (N_3550,In_1259,N_776);
or U3551 (N_3551,In_3425,N_1359);
or U3552 (N_3552,N_1509,In_4661);
nor U3553 (N_3553,In_1534,N_1550);
or U3554 (N_3554,N_1451,N_899);
nor U3555 (N_3555,N_472,In_2027);
xnor U3556 (N_3556,N_1224,N_289);
and U3557 (N_3557,N_1907,In_3869);
nor U3558 (N_3558,N_1399,In_3197);
nand U3559 (N_3559,N_88,N_1512);
nor U3560 (N_3560,N_174,In_1803);
and U3561 (N_3561,In_2338,N_1745);
nor U3562 (N_3562,N_1314,N_815);
nand U3563 (N_3563,In_1112,N_1120);
or U3564 (N_3564,N_1520,N_437);
nand U3565 (N_3565,In_1483,N_1369);
and U3566 (N_3566,N_821,In_3276);
nand U3567 (N_3567,N_939,In_162);
nor U3568 (N_3568,In_4788,N_824);
and U3569 (N_3569,N_972,N_1882);
nor U3570 (N_3570,In_493,N_561);
nor U3571 (N_3571,N_715,N_304);
nand U3572 (N_3572,N_1365,N_1747);
xnor U3573 (N_3573,In_4973,N_1454);
nand U3574 (N_3574,N_431,N_363);
and U3575 (N_3575,N_55,In_3677);
and U3576 (N_3576,N_567,N_902);
nand U3577 (N_3577,In_2899,In_2081);
and U3578 (N_3578,N_1078,N_1529);
or U3579 (N_3579,N_11,N_757);
xnor U3580 (N_3580,N_824,In_2488);
or U3581 (N_3581,In_3181,In_3758);
xnor U3582 (N_3582,N_1127,In_1971);
xnor U3583 (N_3583,In_4711,N_1765);
nor U3584 (N_3584,N_1125,In_4034);
nand U3585 (N_3585,N_1912,N_163);
nor U3586 (N_3586,N_45,In_462);
and U3587 (N_3587,N_452,In_599);
or U3588 (N_3588,In_533,In_1937);
and U3589 (N_3589,In_167,N_1770);
nand U3590 (N_3590,In_4955,N_1708);
and U3591 (N_3591,N_969,In_27);
nor U3592 (N_3592,N_1630,In_1822);
nand U3593 (N_3593,N_225,N_598);
or U3594 (N_3594,N_694,In_2716);
nor U3595 (N_3595,N_913,N_521);
xor U3596 (N_3596,In_650,N_1891);
and U3597 (N_3597,N_1270,In_2407);
or U3598 (N_3598,N_335,N_1006);
and U3599 (N_3599,N_1390,N_15);
nor U3600 (N_3600,N_1337,N_1476);
xor U3601 (N_3601,In_2255,N_703);
and U3602 (N_3602,N_1081,N_1602);
and U3603 (N_3603,In_573,N_1697);
xor U3604 (N_3604,N_1860,In_3146);
nand U3605 (N_3605,N_1971,In_3195);
and U3606 (N_3606,N_1124,N_422);
nand U3607 (N_3607,N_538,N_286);
xor U3608 (N_3608,In_1699,N_1982);
and U3609 (N_3609,In_1699,N_261);
nand U3610 (N_3610,In_3502,N_979);
nor U3611 (N_3611,In_4421,In_4582);
or U3612 (N_3612,N_366,N_258);
nand U3613 (N_3613,N_733,N_141);
nor U3614 (N_3614,N_382,N_938);
nor U3615 (N_3615,In_3509,N_1218);
nand U3616 (N_3616,N_1903,In_755);
nor U3617 (N_3617,In_3450,N_1466);
xnor U3618 (N_3618,N_999,N_199);
nand U3619 (N_3619,N_1425,In_17);
nand U3620 (N_3620,N_1250,N_488);
nand U3621 (N_3621,In_408,N_281);
nor U3622 (N_3622,N_876,In_4124);
nand U3623 (N_3623,N_1937,N_692);
nand U3624 (N_3624,N_1950,N_1190);
or U3625 (N_3625,N_225,In_1483);
nand U3626 (N_3626,In_4614,In_684);
and U3627 (N_3627,N_789,N_648);
nor U3628 (N_3628,N_645,In_2961);
nor U3629 (N_3629,N_1002,N_658);
nand U3630 (N_3630,N_1057,N_865);
nand U3631 (N_3631,N_319,N_1242);
and U3632 (N_3632,N_1180,N_1529);
nor U3633 (N_3633,In_2128,N_506);
xnor U3634 (N_3634,N_44,N_1917);
xnor U3635 (N_3635,In_1905,N_1196);
and U3636 (N_3636,In_4040,In_452);
and U3637 (N_3637,In_655,N_1359);
xor U3638 (N_3638,N_20,N_735);
nand U3639 (N_3639,N_873,N_1665);
xnor U3640 (N_3640,In_4305,In_4751);
xnor U3641 (N_3641,In_4036,N_480);
and U3642 (N_3642,N_1265,N_483);
nor U3643 (N_3643,In_4540,N_1460);
or U3644 (N_3644,In_589,N_681);
or U3645 (N_3645,In_3835,N_1223);
nand U3646 (N_3646,N_900,In_4972);
xnor U3647 (N_3647,N_1267,In_4040);
nor U3648 (N_3648,In_135,N_321);
xnor U3649 (N_3649,In_2305,In_3472);
and U3650 (N_3650,N_1490,N_1272);
nor U3651 (N_3651,In_4129,N_1835);
and U3652 (N_3652,In_1780,In_951);
and U3653 (N_3653,N_1595,N_1489);
nor U3654 (N_3654,N_1992,N_17);
and U3655 (N_3655,N_746,N_1551);
nand U3656 (N_3656,In_588,In_4556);
nand U3657 (N_3657,N_690,N_1143);
xnor U3658 (N_3658,N_278,N_1805);
nand U3659 (N_3659,N_1441,In_2742);
nor U3660 (N_3660,N_106,N_1572);
xor U3661 (N_3661,In_2,N_1261);
and U3662 (N_3662,N_124,In_1159);
xnor U3663 (N_3663,In_2893,In_3533);
xor U3664 (N_3664,N_923,N_84);
nor U3665 (N_3665,N_82,In_764);
xnor U3666 (N_3666,N_1721,N_1664);
and U3667 (N_3667,N_747,In_2076);
or U3668 (N_3668,N_953,N_1416);
xor U3669 (N_3669,N_1029,N_1125);
or U3670 (N_3670,N_1504,N_993);
nand U3671 (N_3671,In_1236,N_1274);
xnor U3672 (N_3672,N_339,In_1493);
and U3673 (N_3673,N_961,In_406);
and U3674 (N_3674,In_1780,In_1747);
and U3675 (N_3675,N_367,N_27);
and U3676 (N_3676,N_824,N_203);
or U3677 (N_3677,N_1555,N_1376);
or U3678 (N_3678,In_1758,In_1447);
nor U3679 (N_3679,In_225,In_4475);
or U3680 (N_3680,N_150,In_653);
xnor U3681 (N_3681,N_10,N_112);
or U3682 (N_3682,N_263,N_389);
nor U3683 (N_3683,N_886,N_1491);
or U3684 (N_3684,N_1377,N_651);
or U3685 (N_3685,N_574,In_4385);
or U3686 (N_3686,N_567,N_380);
or U3687 (N_3687,In_697,N_1079);
or U3688 (N_3688,N_1409,N_725);
nor U3689 (N_3689,N_724,N_532);
and U3690 (N_3690,N_1861,In_1961);
and U3691 (N_3691,N_1552,In_3719);
nand U3692 (N_3692,In_3655,N_603);
or U3693 (N_3693,In_288,N_877);
and U3694 (N_3694,N_1891,In_454);
and U3695 (N_3695,N_589,In_1335);
nor U3696 (N_3696,In_4770,N_1900);
nand U3697 (N_3697,N_361,N_1489);
nand U3698 (N_3698,N_1885,N_1849);
nand U3699 (N_3699,In_4503,In_908);
or U3700 (N_3700,In_4936,N_330);
nor U3701 (N_3701,N_874,In_3736);
xnor U3702 (N_3702,In_373,N_67);
or U3703 (N_3703,N_1926,N_1070);
xor U3704 (N_3704,In_1495,In_2911);
nor U3705 (N_3705,N_1875,N_1770);
xor U3706 (N_3706,N_1519,In_424);
or U3707 (N_3707,N_1915,N_1182);
nand U3708 (N_3708,N_1219,In_1036);
or U3709 (N_3709,N_439,N_984);
or U3710 (N_3710,N_1517,N_587);
or U3711 (N_3711,N_1649,N_218);
xnor U3712 (N_3712,N_525,N_1660);
and U3713 (N_3713,In_2764,N_1325);
nor U3714 (N_3714,N_1533,In_2278);
and U3715 (N_3715,N_412,In_4265);
xnor U3716 (N_3716,N_866,N_1752);
nand U3717 (N_3717,N_974,N_1819);
nand U3718 (N_3718,N_1702,N_1969);
nor U3719 (N_3719,In_2869,N_1058);
nor U3720 (N_3720,In_695,In_2242);
xor U3721 (N_3721,In_597,N_1906);
or U3722 (N_3722,N_1090,In_3628);
nand U3723 (N_3723,In_272,In_1090);
and U3724 (N_3724,N_1232,In_3177);
xor U3725 (N_3725,In_1386,N_1339);
nor U3726 (N_3726,N_1928,In_1107);
nor U3727 (N_3727,N_1639,N_494);
nor U3728 (N_3728,In_3156,In_4582);
nand U3729 (N_3729,N_236,In_1403);
nor U3730 (N_3730,N_308,In_3097);
nand U3731 (N_3731,N_214,In_2030);
nand U3732 (N_3732,In_3408,N_1387);
or U3733 (N_3733,N_1117,In_4375);
or U3734 (N_3734,N_1470,N_1387);
and U3735 (N_3735,N_1719,N_1245);
xor U3736 (N_3736,N_292,N_94);
xor U3737 (N_3737,N_452,In_1487);
and U3738 (N_3738,N_866,In_4459);
xor U3739 (N_3739,N_1757,N_406);
or U3740 (N_3740,In_3454,In_2074);
nor U3741 (N_3741,N_1973,N_858);
and U3742 (N_3742,N_1080,N_1720);
nor U3743 (N_3743,N_1518,N_350);
nand U3744 (N_3744,N_1709,N_482);
nand U3745 (N_3745,N_1312,N_1580);
xor U3746 (N_3746,N_23,N_1868);
xnor U3747 (N_3747,N_1288,N_1657);
xor U3748 (N_3748,In_3177,N_1097);
xor U3749 (N_3749,In_4449,N_1012);
nor U3750 (N_3750,N_1702,N_1426);
nor U3751 (N_3751,In_684,N_688);
nor U3752 (N_3752,In_4390,In_4139);
or U3753 (N_3753,N_655,In_1618);
xnor U3754 (N_3754,In_405,In_1066);
nor U3755 (N_3755,N_1697,In_1223);
xor U3756 (N_3756,In_3065,N_1155);
nand U3757 (N_3757,N_147,N_1605);
or U3758 (N_3758,N_103,In_1546);
and U3759 (N_3759,N_1613,In_3558);
xor U3760 (N_3760,N_1557,In_4449);
nor U3761 (N_3761,N_889,N_813);
xor U3762 (N_3762,In_1217,In_4872);
xor U3763 (N_3763,N_921,N_884);
and U3764 (N_3764,In_2562,N_1671);
nor U3765 (N_3765,In_1349,N_1967);
and U3766 (N_3766,N_1931,N_668);
and U3767 (N_3767,N_1293,N_1694);
and U3768 (N_3768,N_621,N_1449);
and U3769 (N_3769,In_4761,In_4232);
or U3770 (N_3770,In_2847,N_1901);
nor U3771 (N_3771,N_1143,N_1530);
or U3772 (N_3772,In_4339,N_1024);
nand U3773 (N_3773,In_4788,N_1814);
or U3774 (N_3774,In_1126,In_1655);
xor U3775 (N_3775,In_1057,In_3201);
nor U3776 (N_3776,N_944,N_871);
xnor U3777 (N_3777,In_2264,N_215);
and U3778 (N_3778,N_1727,N_1835);
or U3779 (N_3779,N_307,N_1164);
xor U3780 (N_3780,N_1361,N_1561);
nand U3781 (N_3781,In_4919,In_4539);
and U3782 (N_3782,N_397,N_1959);
nand U3783 (N_3783,In_3122,N_1854);
nor U3784 (N_3784,In_4849,N_93);
xor U3785 (N_3785,N_394,N_1640);
xnor U3786 (N_3786,In_4859,N_1517);
or U3787 (N_3787,In_452,N_1365);
and U3788 (N_3788,N_1487,In_4071);
and U3789 (N_3789,N_935,N_1698);
xor U3790 (N_3790,In_422,In_2401);
and U3791 (N_3791,N_1063,N_18);
and U3792 (N_3792,N_1262,In_4633);
and U3793 (N_3793,In_3266,N_1891);
or U3794 (N_3794,In_764,N_141);
nor U3795 (N_3795,In_4399,N_571);
nor U3796 (N_3796,N_1164,N_1116);
nor U3797 (N_3797,N_84,N_584);
nand U3798 (N_3798,In_1147,In_2864);
and U3799 (N_3799,N_330,N_545);
xor U3800 (N_3800,N_1431,In_4867);
xor U3801 (N_3801,In_4556,N_1097);
nand U3802 (N_3802,In_3314,N_1353);
or U3803 (N_3803,N_1896,N_1330);
or U3804 (N_3804,N_632,In_3370);
or U3805 (N_3805,N_597,N_34);
xnor U3806 (N_3806,N_1434,In_4700);
and U3807 (N_3807,N_149,N_1704);
nand U3808 (N_3808,N_35,In_1967);
nor U3809 (N_3809,In_2935,N_819);
and U3810 (N_3810,N_726,N_1089);
nand U3811 (N_3811,In_3893,In_671);
nor U3812 (N_3812,N_1535,In_4294);
nand U3813 (N_3813,N_1808,In_1183);
or U3814 (N_3814,In_252,In_3824);
nor U3815 (N_3815,N_1543,In_4131);
nor U3816 (N_3816,In_4522,N_1107);
xor U3817 (N_3817,N_1142,N_530);
or U3818 (N_3818,In_4474,N_205);
xor U3819 (N_3819,N_1009,In_695);
and U3820 (N_3820,N_1475,In_4338);
and U3821 (N_3821,In_101,In_4269);
nand U3822 (N_3822,In_2193,N_591);
and U3823 (N_3823,N_1306,N_1397);
xor U3824 (N_3824,In_339,In_1919);
or U3825 (N_3825,N_1487,In_3844);
and U3826 (N_3826,In_1145,N_1930);
xor U3827 (N_3827,In_2905,In_2401);
or U3828 (N_3828,N_822,In_547);
and U3829 (N_3829,In_3832,N_24);
nand U3830 (N_3830,N_1167,N_1093);
nor U3831 (N_3831,N_1144,N_1940);
or U3832 (N_3832,N_1812,N_1697);
nor U3833 (N_3833,N_1966,N_1492);
or U3834 (N_3834,N_196,In_3480);
or U3835 (N_3835,N_1010,N_1583);
or U3836 (N_3836,In_3736,In_4973);
and U3837 (N_3837,In_3382,In_4136);
xnor U3838 (N_3838,N_364,In_2837);
xnor U3839 (N_3839,N_345,N_805);
and U3840 (N_3840,In_1999,N_1357);
nand U3841 (N_3841,N_1349,N_1860);
or U3842 (N_3842,N_69,N_1315);
nand U3843 (N_3843,N_1221,N_1582);
or U3844 (N_3844,In_2443,In_4505);
xnor U3845 (N_3845,N_568,N_425);
nor U3846 (N_3846,N_725,N_1673);
xnor U3847 (N_3847,N_1653,N_205);
xnor U3848 (N_3848,In_1967,In_4272);
nor U3849 (N_3849,N_1698,N_1074);
nand U3850 (N_3850,N_1208,N_1063);
and U3851 (N_3851,N_1248,N_261);
nand U3852 (N_3852,N_1317,N_941);
nor U3853 (N_3853,N_1061,N_705);
nand U3854 (N_3854,N_684,N_1360);
and U3855 (N_3855,N_699,N_475);
nand U3856 (N_3856,N_1240,In_4746);
or U3857 (N_3857,N_1814,N_1002);
or U3858 (N_3858,N_68,N_239);
xor U3859 (N_3859,N_1003,N_116);
or U3860 (N_3860,In_695,N_491);
nand U3861 (N_3861,In_191,In_2079);
nor U3862 (N_3862,N_1510,In_4036);
and U3863 (N_3863,In_3655,In_1936);
nor U3864 (N_3864,In_3773,N_1336);
and U3865 (N_3865,N_1711,N_14);
or U3866 (N_3866,N_1469,N_1708);
nand U3867 (N_3867,In_3216,N_1679);
xnor U3868 (N_3868,N_1902,N_488);
nor U3869 (N_3869,N_1532,N_704);
and U3870 (N_3870,N_1122,N_1534);
nand U3871 (N_3871,N_1711,N_564);
xor U3872 (N_3872,In_1463,N_1957);
and U3873 (N_3873,In_3951,In_1622);
nand U3874 (N_3874,N_805,N_1168);
xnor U3875 (N_3875,N_1988,N_255);
xnor U3876 (N_3876,N_127,In_3946);
nor U3877 (N_3877,In_1182,N_962);
nor U3878 (N_3878,N_937,In_4122);
xor U3879 (N_3879,N_74,In_4809);
nor U3880 (N_3880,N_540,In_2131);
xor U3881 (N_3881,In_3873,N_1736);
xor U3882 (N_3882,N_1191,N_292);
and U3883 (N_3883,N_1086,In_4605);
nor U3884 (N_3884,N_855,N_341);
nor U3885 (N_3885,N_1752,N_1358);
nor U3886 (N_3886,In_3065,N_1142);
nor U3887 (N_3887,N_1066,N_765);
and U3888 (N_3888,In_966,N_695);
or U3889 (N_3889,N_295,N_1640);
or U3890 (N_3890,In_4598,In_4997);
or U3891 (N_3891,In_4057,N_1073);
nand U3892 (N_3892,In_1060,N_1259);
and U3893 (N_3893,N_506,N_1352);
or U3894 (N_3894,N_235,N_1720);
and U3895 (N_3895,N_977,N_1455);
or U3896 (N_3896,N_1595,In_755);
nand U3897 (N_3897,N_697,N_16);
nand U3898 (N_3898,In_1736,N_202);
and U3899 (N_3899,In_1622,In_3425);
nand U3900 (N_3900,N_286,N_1774);
xor U3901 (N_3901,In_2234,In_3177);
xor U3902 (N_3902,N_435,N_1237);
nand U3903 (N_3903,N_668,In_2725);
or U3904 (N_3904,In_2935,In_1243);
or U3905 (N_3905,N_1934,In_4594);
or U3906 (N_3906,N_1997,N_432);
or U3907 (N_3907,N_806,N_1437);
nand U3908 (N_3908,N_742,In_3614);
and U3909 (N_3909,In_2848,In_1177);
xor U3910 (N_3910,N_1455,In_2200);
nor U3911 (N_3911,In_3913,N_798);
xnor U3912 (N_3912,In_4984,N_1268);
nand U3913 (N_3913,N_1207,In_240);
xnor U3914 (N_3914,N_1857,In_554);
and U3915 (N_3915,In_774,N_938);
nor U3916 (N_3916,N_18,N_1023);
nand U3917 (N_3917,N_1380,N_1894);
nor U3918 (N_3918,In_3497,In_4677);
or U3919 (N_3919,In_4571,N_1168);
xor U3920 (N_3920,N_195,In_4377);
and U3921 (N_3921,N_976,N_1337);
and U3922 (N_3922,N_370,N_1142);
and U3923 (N_3923,N_1838,In_4334);
nand U3924 (N_3924,N_456,N_606);
and U3925 (N_3925,N_955,N_196);
xnor U3926 (N_3926,N_1574,In_2222);
nand U3927 (N_3927,N_540,N_1837);
or U3928 (N_3928,N_1951,N_1544);
xnor U3929 (N_3929,N_693,N_1799);
nor U3930 (N_3930,N_875,In_2580);
xor U3931 (N_3931,N_853,N_1320);
nand U3932 (N_3932,N_1699,N_454);
xor U3933 (N_3933,N_1655,N_1291);
or U3934 (N_3934,N_1013,N_458);
nor U3935 (N_3935,N_1991,N_1158);
and U3936 (N_3936,In_3097,In_3946);
nand U3937 (N_3937,N_74,In_1279);
or U3938 (N_3938,N_1881,In_4714);
or U3939 (N_3939,In_781,In_2590);
nor U3940 (N_3940,N_99,N_41);
or U3941 (N_3941,N_350,N_338);
nor U3942 (N_3942,N_755,N_353);
and U3943 (N_3943,N_1962,N_1658);
nor U3944 (N_3944,In_2243,N_1085);
xnor U3945 (N_3945,N_1,N_876);
nand U3946 (N_3946,N_1447,In_1546);
and U3947 (N_3947,N_1955,In_2995);
nand U3948 (N_3948,In_3748,N_742);
and U3949 (N_3949,In_4571,N_605);
or U3950 (N_3950,In_3844,In_1917);
xnor U3951 (N_3951,In_4254,N_579);
or U3952 (N_3952,N_1902,In_388);
nand U3953 (N_3953,N_1560,N_1563);
and U3954 (N_3954,In_217,N_1820);
and U3955 (N_3955,N_1803,N_1595);
and U3956 (N_3956,N_1292,In_1854);
nor U3957 (N_3957,N_1994,N_1905);
or U3958 (N_3958,N_3,In_2874);
xor U3959 (N_3959,In_4836,In_1319);
nor U3960 (N_3960,N_1376,In_4713);
nand U3961 (N_3961,N_1325,N_1951);
nor U3962 (N_3962,In_965,N_855);
and U3963 (N_3963,N_863,N_1066);
nor U3964 (N_3964,In_2721,N_143);
xor U3965 (N_3965,N_989,N_1402);
xnor U3966 (N_3966,N_745,N_1420);
nor U3967 (N_3967,In_1915,In_2911);
and U3968 (N_3968,N_1753,N_470);
nor U3969 (N_3969,N_958,N_863);
and U3970 (N_3970,N_892,In_2189);
nor U3971 (N_3971,In_3480,N_1205);
nand U3972 (N_3972,N_1560,N_1119);
and U3973 (N_3973,N_1466,N_645);
nand U3974 (N_3974,N_1875,N_317);
nor U3975 (N_3975,In_3692,N_1189);
nand U3976 (N_3976,N_1252,N_1847);
nand U3977 (N_3977,N_236,N_691);
or U3978 (N_3978,In_3169,N_1024);
and U3979 (N_3979,N_133,N_1341);
nand U3980 (N_3980,N_608,N_478);
xnor U3981 (N_3981,N_942,N_797);
or U3982 (N_3982,N_1431,N_1342);
nand U3983 (N_3983,N_310,N_1183);
xor U3984 (N_3984,N_1497,N_1780);
and U3985 (N_3985,In_455,In_4131);
nand U3986 (N_3986,N_1094,N_1051);
nand U3987 (N_3987,N_1766,In_4919);
nor U3988 (N_3988,N_1790,In_3614);
nor U3989 (N_3989,In_3766,N_1495);
xor U3990 (N_3990,N_1870,N_134);
nand U3991 (N_3991,In_748,N_1482);
or U3992 (N_3992,In_2227,N_1276);
and U3993 (N_3993,N_1506,In_2285);
and U3994 (N_3994,In_162,In_4637);
nand U3995 (N_3995,N_91,N_41);
nand U3996 (N_3996,N_1755,N_1129);
or U3997 (N_3997,N_1688,N_1047);
nor U3998 (N_3998,N_1067,In_1804);
or U3999 (N_3999,N_1727,In_1279);
xor U4000 (N_4000,N_2729,N_3948);
and U4001 (N_4001,N_2691,N_2350);
nor U4002 (N_4002,N_2391,N_3640);
nor U4003 (N_4003,N_3944,N_3504);
nor U4004 (N_4004,N_2803,N_2148);
or U4005 (N_4005,N_2302,N_2035);
xor U4006 (N_4006,N_2839,N_2010);
nor U4007 (N_4007,N_3184,N_3069);
nor U4008 (N_4008,N_3838,N_2790);
nand U4009 (N_4009,N_2493,N_2125);
or U4010 (N_4010,N_3606,N_3506);
and U4011 (N_4011,N_3732,N_2914);
nor U4012 (N_4012,N_2544,N_3302);
nor U4013 (N_4013,N_3756,N_3719);
and U4014 (N_4014,N_2249,N_3533);
nand U4015 (N_4015,N_2868,N_2353);
nand U4016 (N_4016,N_3730,N_3201);
and U4017 (N_4017,N_2157,N_2910);
xor U4018 (N_4018,N_2099,N_3537);
nor U4019 (N_4019,N_2956,N_3662);
nand U4020 (N_4020,N_3355,N_2895);
nor U4021 (N_4021,N_3768,N_3113);
nand U4022 (N_4022,N_2921,N_3748);
or U4023 (N_4023,N_2251,N_3656);
xor U4024 (N_4024,N_2813,N_2404);
or U4025 (N_4025,N_2036,N_2153);
or U4026 (N_4026,N_3362,N_3042);
nand U4027 (N_4027,N_2294,N_3356);
xnor U4028 (N_4028,N_3697,N_2114);
and U4029 (N_4029,N_3933,N_2333);
and U4030 (N_4030,N_3546,N_3381);
xor U4031 (N_4031,N_2420,N_3554);
nand U4032 (N_4032,N_3293,N_3314);
nor U4033 (N_4033,N_2082,N_2534);
xnor U4034 (N_4034,N_3815,N_2015);
or U4035 (N_4035,N_2108,N_3325);
xnor U4036 (N_4036,N_2945,N_2808);
or U4037 (N_4037,N_3103,N_2201);
or U4038 (N_4038,N_3307,N_3954);
nand U4039 (N_4039,N_2820,N_2609);
nor U4040 (N_4040,N_2199,N_3187);
xnor U4041 (N_4041,N_3932,N_3185);
nor U4042 (N_4042,N_2998,N_2715);
and U4043 (N_4043,N_3050,N_2115);
xnor U4044 (N_4044,N_2445,N_2573);
xor U4045 (N_4045,N_2190,N_2159);
or U4046 (N_4046,N_3889,N_2365);
or U4047 (N_4047,N_2287,N_3845);
nor U4048 (N_4048,N_2706,N_3995);
and U4049 (N_4049,N_3249,N_2112);
or U4050 (N_4050,N_3903,N_2279);
xnor U4051 (N_4051,N_3475,N_2075);
and U4052 (N_4052,N_2459,N_3658);
or U4053 (N_4053,N_3073,N_2216);
and U4054 (N_4054,N_3476,N_2598);
xor U4055 (N_4055,N_2801,N_3923);
and U4056 (N_4056,N_2139,N_2384);
nor U4057 (N_4057,N_2746,N_3760);
nand U4058 (N_4058,N_3959,N_2781);
xor U4059 (N_4059,N_2622,N_2649);
xor U4060 (N_4060,N_3603,N_2673);
nor U4061 (N_4061,N_2507,N_3028);
or U4062 (N_4062,N_3345,N_2959);
and U4063 (N_4063,N_2854,N_3638);
nand U4064 (N_4064,N_3856,N_3502);
nand U4065 (N_4065,N_3967,N_3007);
or U4066 (N_4066,N_2032,N_3005);
nor U4067 (N_4067,N_3551,N_2906);
nor U4068 (N_4068,N_3762,N_3189);
and U4069 (N_4069,N_2499,N_2227);
nand U4070 (N_4070,N_2861,N_3994);
or U4071 (N_4071,N_3677,N_2393);
or U4072 (N_4072,N_2777,N_2197);
and U4073 (N_4073,N_2555,N_3421);
and U4074 (N_4074,N_2186,N_3904);
or U4075 (N_4075,N_3898,N_3951);
nor U4076 (N_4076,N_2345,N_3444);
xnor U4077 (N_4077,N_2289,N_2497);
and U4078 (N_4078,N_3055,N_2319);
nand U4079 (N_4079,N_2326,N_3065);
or U4080 (N_4080,N_3135,N_3264);
nand U4081 (N_4081,N_2455,N_3150);
nand U4082 (N_4082,N_2750,N_2958);
xor U4083 (N_4083,N_3346,N_2709);
xor U4084 (N_4084,N_3172,N_3012);
xnor U4085 (N_4085,N_3848,N_2274);
xnor U4086 (N_4086,N_3819,N_3206);
nand U4087 (N_4087,N_2933,N_3695);
and U4088 (N_4088,N_2204,N_3383);
xor U4089 (N_4089,N_2177,N_3046);
xor U4090 (N_4090,N_2261,N_3772);
nand U4091 (N_4091,N_2782,N_3975);
or U4092 (N_4092,N_3575,N_3597);
and U4093 (N_4093,N_3268,N_2971);
xnor U4094 (N_4094,N_2331,N_2200);
nand U4095 (N_4095,N_2038,N_3557);
xor U4096 (N_4096,N_3099,N_3990);
nand U4097 (N_4097,N_3952,N_2309);
and U4098 (N_4098,N_2702,N_2191);
nor U4099 (N_4099,N_2654,N_3207);
xnor U4100 (N_4100,N_2775,N_2795);
nor U4101 (N_4101,N_2539,N_3622);
or U4102 (N_4102,N_2024,N_3626);
xor U4103 (N_4103,N_2018,N_2448);
xnor U4104 (N_4104,N_3721,N_3374);
nor U4105 (N_4105,N_2286,N_2442);
nand U4106 (N_4106,N_2124,N_2911);
or U4107 (N_4107,N_3254,N_2441);
nor U4108 (N_4108,N_2903,N_2436);
xor U4109 (N_4109,N_3231,N_2460);
xnor U4110 (N_4110,N_2704,N_3218);
and U4111 (N_4111,N_2554,N_2826);
nand U4112 (N_4112,N_2072,N_2561);
nand U4113 (N_4113,N_3577,N_3870);
nand U4114 (N_4114,N_2871,N_2918);
nand U4115 (N_4115,N_3177,N_2389);
nand U4116 (N_4116,N_2060,N_2402);
and U4117 (N_4117,N_3263,N_3864);
nand U4118 (N_4118,N_2986,N_2532);
xnor U4119 (N_4119,N_3781,N_3270);
nor U4120 (N_4120,N_3223,N_2504);
or U4121 (N_4121,N_2007,N_2821);
and U4122 (N_4122,N_2527,N_2583);
or U4123 (N_4123,N_2901,N_3003);
or U4124 (N_4124,N_3262,N_3633);
or U4125 (N_4125,N_3868,N_2881);
and U4126 (N_4126,N_2011,N_3163);
nor U4127 (N_4127,N_2033,N_2163);
or U4128 (N_4128,N_3623,N_3233);
or U4129 (N_4129,N_3988,N_3497);
xor U4130 (N_4130,N_2482,N_3459);
nand U4131 (N_4131,N_2217,N_3826);
nand U4132 (N_4132,N_3429,N_2266);
xor U4133 (N_4133,N_3029,N_3559);
and U4134 (N_4134,N_3479,N_3717);
xor U4135 (N_4135,N_2117,N_3538);
and U4136 (N_4136,N_3271,N_2156);
nand U4137 (N_4137,N_2833,N_2046);
or U4138 (N_4138,N_3681,N_3043);
or U4139 (N_4139,N_2541,N_2263);
and U4140 (N_4140,N_2693,N_2488);
xnor U4141 (N_4141,N_2714,N_2999);
or U4142 (N_4142,N_3128,N_2961);
xnor U4143 (N_4143,N_2860,N_2167);
and U4144 (N_4144,N_2503,N_2847);
or U4145 (N_4145,N_2663,N_3365);
nand U4146 (N_4146,N_2373,N_3058);
or U4147 (N_4147,N_3326,N_2666);
or U4148 (N_4148,N_3956,N_2919);
or U4149 (N_4149,N_3339,N_2815);
nand U4150 (N_4150,N_3408,N_3914);
nor U4151 (N_4151,N_2763,N_3410);
nand U4152 (N_4152,N_2343,N_2852);
nor U4153 (N_4153,N_3129,N_3417);
xor U4154 (N_4154,N_3066,N_2454);
nand U4155 (N_4155,N_3379,N_2092);
nand U4156 (N_4156,N_2669,N_3261);
nand U4157 (N_4157,N_2981,N_2472);
xor U4158 (N_4158,N_2337,N_3440);
and U4159 (N_4159,N_3322,N_3100);
or U4160 (N_4160,N_2665,N_3616);
or U4161 (N_4161,N_2856,N_2681);
or U4162 (N_4162,N_3996,N_3032);
or U4163 (N_4163,N_2427,N_2796);
and U4164 (N_4164,N_3037,N_2275);
nand U4165 (N_4165,N_3160,N_2152);
nor U4166 (N_4166,N_3666,N_2458);
nor U4167 (N_4167,N_3534,N_3727);
nand U4168 (N_4168,N_2413,N_2676);
or U4169 (N_4169,N_2461,N_3225);
nor U4170 (N_4170,N_2724,N_2996);
xor U4171 (N_4171,N_3652,N_3125);
xnor U4172 (N_4172,N_3074,N_2762);
and U4173 (N_4173,N_2338,N_3624);
xor U4174 (N_4174,N_3503,N_2579);
nor U4175 (N_4175,N_2096,N_2935);
nand U4176 (N_4176,N_3422,N_2738);
xor U4177 (N_4177,N_3494,N_3495);
or U4178 (N_4178,N_3399,N_2645);
nand U4179 (N_4179,N_3902,N_2019);
nor U4180 (N_4180,N_3824,N_3349);
nand U4181 (N_4181,N_2987,N_2926);
or U4182 (N_4182,N_3619,N_3816);
nor U4183 (N_4183,N_2209,N_2969);
and U4184 (N_4184,N_2859,N_3361);
nor U4185 (N_4185,N_3310,N_2941);
and U4186 (N_4186,N_3237,N_2136);
and U4187 (N_4187,N_2451,N_2978);
or U4188 (N_4188,N_2589,N_3894);
nor U4189 (N_4189,N_3700,N_3654);
or U4190 (N_4190,N_3871,N_2749);
and U4191 (N_4191,N_3153,N_3614);
or U4192 (N_4192,N_3663,N_2247);
nor U4193 (N_4193,N_3333,N_3387);
or U4194 (N_4194,N_2180,N_3543);
or U4195 (N_4195,N_3910,N_3794);
nand U4196 (N_4196,N_3330,N_2651);
or U4197 (N_4197,N_2169,N_2515);
nor U4198 (N_4198,N_3085,N_3409);
or U4199 (N_4199,N_2193,N_2980);
nand U4200 (N_4200,N_3696,N_2196);
or U4201 (N_4201,N_2964,N_2601);
nor U4202 (N_4202,N_3507,N_3465);
nand U4203 (N_4203,N_3404,N_3305);
xor U4204 (N_4204,N_2138,N_3735);
nand U4205 (N_4205,N_2817,N_3808);
or U4206 (N_4206,N_3525,N_2265);
nor U4207 (N_4207,N_3803,N_3216);
xor U4208 (N_4208,N_3512,N_3139);
or U4209 (N_4209,N_3392,N_3532);
or U4210 (N_4210,N_2065,N_2627);
nand U4211 (N_4211,N_2122,N_2770);
and U4212 (N_4212,N_3335,N_2017);
or U4213 (N_4213,N_2475,N_3167);
nand U4214 (N_4214,N_2248,N_2178);
and U4215 (N_4215,N_2634,N_3131);
and U4216 (N_4216,N_3805,N_2235);
xor U4217 (N_4217,N_3395,N_2698);
and U4218 (N_4218,N_3832,N_3242);
xor U4219 (N_4219,N_2757,N_3403);
xor U4220 (N_4220,N_3318,N_3490);
and U4221 (N_4221,N_3215,N_2735);
and U4222 (N_4222,N_2085,N_3574);
xnor U4223 (N_4223,N_2540,N_2473);
nor U4224 (N_4224,N_3137,N_3885);
xnor U4225 (N_4225,N_2814,N_3340);
and U4226 (N_4226,N_2581,N_3428);
nor U4227 (N_4227,N_2421,N_2298);
or U4228 (N_4228,N_2510,N_2246);
nor U4229 (N_4229,N_2466,N_2822);
xnor U4230 (N_4230,N_3839,N_2327);
xor U4231 (N_4231,N_2412,N_2536);
xor U4232 (N_4232,N_2121,N_3170);
or U4233 (N_4233,N_2374,N_2483);
nor U4234 (N_4234,N_2359,N_3847);
nor U4235 (N_4235,N_3936,N_3204);
nor U4236 (N_4236,N_2525,N_2074);
nor U4237 (N_4237,N_2551,N_2277);
nor U4238 (N_4238,N_3863,N_2680);
and U4239 (N_4239,N_3929,N_2872);
nor U4240 (N_4240,N_3558,N_2106);
nor U4241 (N_4241,N_3049,N_3369);
or U4242 (N_4242,N_3222,N_3252);
xor U4243 (N_4243,N_3670,N_3935);
or U4244 (N_4244,N_3843,N_2633);
or U4245 (N_4245,N_2849,N_2982);
nor U4246 (N_4246,N_2495,N_3061);
nor U4247 (N_4247,N_3977,N_3306);
nor U4248 (N_4248,N_2638,N_3778);
nor U4249 (N_4249,N_3829,N_2722);
nor U4250 (N_4250,N_3442,N_2269);
nand U4251 (N_4251,N_3517,N_3548);
nand U4252 (N_4252,N_2563,N_2479);
and U4253 (N_4253,N_2809,N_2765);
and U4254 (N_4254,N_3972,N_2097);
nand U4255 (N_4255,N_2165,N_2192);
nand U4256 (N_4256,N_3458,N_2054);
nor U4257 (N_4257,N_2751,N_3436);
nand U4258 (N_4258,N_3704,N_2635);
xnor U4259 (N_4259,N_3774,N_2219);
nor U4260 (N_4260,N_3284,N_2823);
xor U4261 (N_4261,N_2592,N_3942);
and U4262 (N_4262,N_2487,N_2925);
nor U4263 (N_4263,N_2582,N_3934);
xor U4264 (N_4264,N_3985,N_2432);
and U4265 (N_4265,N_2284,N_2357);
or U4266 (N_4266,N_2913,N_2008);
nor U4267 (N_4267,N_3390,N_2417);
xor U4268 (N_4268,N_2344,N_3716);
xnor U4269 (N_4269,N_2937,N_3583);
and U4270 (N_4270,N_3324,N_2968);
and U4271 (N_4271,N_2256,N_3777);
nor U4272 (N_4272,N_2712,N_3641);
nand U4273 (N_4273,N_3315,N_3859);
and U4274 (N_4274,N_3445,N_3023);
xor U4275 (N_4275,N_3414,N_3776);
xnor U4276 (N_4276,N_3097,N_2317);
nor U4277 (N_4277,N_3115,N_2686);
nor U4278 (N_4278,N_2876,N_2789);
xnor U4279 (N_4279,N_2772,N_2137);
nand U4280 (N_4280,N_3499,N_2807);
or U4281 (N_4281,N_2840,N_2250);
nor U4282 (N_4282,N_2595,N_2143);
nand U4283 (N_4283,N_2688,N_2324);
or U4284 (N_4284,N_3680,N_3560);
nor U4285 (N_4285,N_2005,N_2494);
nand U4286 (N_4286,N_2077,N_2875);
or U4287 (N_4287,N_2816,N_3511);
or U4288 (N_4288,N_2089,N_3950);
nor U4289 (N_4289,N_2118,N_3120);
or U4290 (N_4290,N_3474,N_2929);
and U4291 (N_4291,N_3960,N_2175);
or U4292 (N_4292,N_3290,N_3643);
nor U4293 (N_4293,N_2129,N_2321);
nor U4294 (N_4294,N_2398,N_3737);
nand U4295 (N_4295,N_3620,N_3926);
nor U4296 (N_4296,N_2492,N_2119);
nor U4297 (N_4297,N_2194,N_3057);
nand U4298 (N_4298,N_3689,N_2542);
or U4299 (N_4299,N_2245,N_3683);
or U4300 (N_4300,N_3782,N_2073);
xnor U4301 (N_4301,N_3759,N_3287);
nand U4302 (N_4302,N_3797,N_2838);
and U4303 (N_4303,N_3004,N_2362);
and U4304 (N_4304,N_3478,N_2556);
nand U4305 (N_4305,N_3970,N_3412);
nor U4306 (N_4306,N_3068,N_3178);
xnor U4307 (N_4307,N_2127,N_2034);
and U4308 (N_4308,N_2785,N_3541);
nor U4309 (N_4309,N_2526,N_2012);
or U4310 (N_4310,N_3174,N_2113);
xnor U4311 (N_4311,N_3925,N_3449);
or U4312 (N_4312,N_3814,N_2195);
nor U4313 (N_4313,N_2993,N_2835);
nor U4314 (N_4314,N_2737,N_2375);
and U4315 (N_4315,N_2597,N_2845);
xor U4316 (N_4316,N_2335,N_2141);
nand U4317 (N_4317,N_3605,N_3562);
nand U4318 (N_4318,N_3397,N_2985);
and U4319 (N_4319,N_3675,N_3523);
nor U4320 (N_4320,N_3011,N_2890);
nand U4321 (N_4321,N_2316,N_2356);
nor U4322 (N_4322,N_3527,N_3796);
or U4323 (N_4323,N_3489,N_3779);
or U4324 (N_4324,N_2111,N_3687);
or U4325 (N_4325,N_3432,N_2128);
and U4326 (N_4326,N_3292,N_3389);
nor U4327 (N_4327,N_3338,N_3569);
nor U4328 (N_4328,N_3480,N_3878);
nor U4329 (N_4329,N_3198,N_3496);
xor U4330 (N_4330,N_2967,N_3299);
and U4331 (N_4331,N_2867,N_3630);
nand U4332 (N_4332,N_2948,N_3062);
nand U4333 (N_4333,N_3565,N_3539);
nor U4334 (N_4334,N_3118,N_2960);
nand U4335 (N_4335,N_3590,N_3446);
or U4336 (N_4336,N_3133,N_2006);
nor U4337 (N_4337,N_3837,N_2378);
xor U4338 (N_4338,N_3966,N_2748);
or U4339 (N_4339,N_2135,N_2283);
xor U4340 (N_4340,N_3659,N_3621);
nor U4341 (N_4341,N_3400,N_2208);
or U4342 (N_4342,N_2626,N_2218);
and U4343 (N_4343,N_3833,N_2411);
or U4344 (N_4344,N_2798,N_2002);
xor U4345 (N_4345,N_3352,N_2325);
nand U4346 (N_4346,N_3370,N_2829);
and U4347 (N_4347,N_2270,N_2656);
and U4348 (N_4348,N_2334,N_2014);
nor U4349 (N_4349,N_3450,N_3881);
nor U4350 (N_4350,N_2831,N_3513);
xor U4351 (N_4351,N_2304,N_3752);
nand U4352 (N_4352,N_2701,N_3526);
or U4353 (N_4353,N_3462,N_3300);
nand U4354 (N_4354,N_3039,N_2907);
xnor U4355 (N_4355,N_3741,N_3866);
nand U4356 (N_4356,N_3107,N_3679);
and U4357 (N_4357,N_3056,N_2667);
nand U4358 (N_4358,N_2853,N_3976);
nand U4359 (N_4359,N_3745,N_3088);
and U4360 (N_4360,N_2509,N_2733);
xor U4361 (N_4361,N_2290,N_2857);
nor U4362 (N_4362,N_3441,N_3992);
or U4363 (N_4363,N_2502,N_2400);
and U4364 (N_4364,N_3722,N_3612);
xor U4365 (N_4365,N_3544,N_2130);
or U4366 (N_4366,N_2569,N_2004);
or U4367 (N_4367,N_3301,N_3147);
nand U4368 (N_4368,N_3709,N_3867);
and U4369 (N_4369,N_3141,N_2151);
xnor U4370 (N_4370,N_2491,N_2946);
nand U4371 (N_4371,N_2804,N_3281);
nor U4372 (N_4372,N_2930,N_2048);
or U4373 (N_4373,N_2550,N_2576);
and U4374 (N_4374,N_3013,N_3265);
xnor U4375 (N_4375,N_2766,N_2568);
nand U4376 (N_4376,N_3757,N_3649);
nand U4377 (N_4377,N_3158,N_3336);
xnor U4378 (N_4378,N_3010,N_3647);
nor U4379 (N_4379,N_2564,N_3602);
xor U4380 (N_4380,N_3821,N_3059);
and U4381 (N_4381,N_2030,N_3684);
or U4382 (N_4382,N_3105,N_3609);
or U4383 (N_4383,N_3921,N_3175);
nor U4384 (N_4384,N_2767,N_3550);
or U4385 (N_4385,N_2932,N_3214);
nand U4386 (N_4386,N_2366,N_3733);
nor U4387 (N_4387,N_3750,N_2323);
nand U4388 (N_4388,N_3485,N_2668);
and U4389 (N_4389,N_2575,N_3908);
or U4390 (N_4390,N_3718,N_2642);
and U4391 (N_4391,N_2992,N_2897);
nor U4392 (N_4392,N_3580,N_2203);
nor U4393 (N_4393,N_2719,N_2489);
or U4394 (N_4394,N_3121,N_2887);
and U4395 (N_4395,N_3209,N_3382);
nor U4396 (N_4396,N_3702,N_2874);
xnor U4397 (N_4397,N_3317,N_3849);
xnor U4398 (N_4398,N_2098,N_2655);
and U4399 (N_4399,N_3228,N_3134);
and U4400 (N_4400,N_2025,N_2022);
and U4401 (N_4401,N_2718,N_2332);
nand U4402 (N_4402,N_2272,N_2239);
and U4403 (N_4403,N_3452,N_3396);
nand U4404 (N_4404,N_2285,N_3655);
or U4405 (N_4405,N_2027,N_3787);
xnor U4406 (N_4406,N_2705,N_3909);
and U4407 (N_4407,N_2524,N_2320);
nand U4408 (N_4408,N_3501,N_2434);
nor U4409 (N_4409,N_3251,N_3740);
xnor U4410 (N_4410,N_3146,N_3822);
nand U4411 (N_4411,N_3469,N_3993);
nand U4412 (N_4412,N_3457,N_3211);
or U4413 (N_4413,N_2703,N_3785);
or U4414 (N_4414,N_3997,N_3269);
nor U4415 (N_4415,N_3792,N_3706);
xor U4416 (N_4416,N_3599,N_3940);
and U4417 (N_4417,N_2846,N_3094);
nand U4418 (N_4418,N_2549,N_2403);
xnor U4419 (N_4419,N_3522,N_3698);
or U4420 (N_4420,N_3138,N_2444);
nor U4421 (N_4421,N_2023,N_2602);
and U4422 (N_4422,N_2588,N_2259);
or U4423 (N_4423,N_2844,N_3596);
and U4424 (N_4424,N_2039,N_2214);
nor U4425 (N_4425,N_3810,N_2303);
and U4426 (N_4426,N_2614,N_2878);
nor U4427 (N_4427,N_3991,N_2707);
and U4428 (N_4428,N_2425,N_3391);
xnor U4429 (N_4429,N_2963,N_2858);
nor U4430 (N_4430,N_3416,N_3608);
nand U4431 (N_4431,N_2222,N_2570);
and U4432 (N_4432,N_3401,N_2950);
xor U4433 (N_4433,N_2288,N_2580);
and U4434 (N_4434,N_2720,N_2088);
nand U4435 (N_4435,N_2690,N_3931);
or U4436 (N_4436,N_2896,N_3793);
xnor U4437 (N_4437,N_2684,N_2140);
and U4438 (N_4438,N_2947,N_3584);
nand U4439 (N_4439,N_3283,N_3686);
nand U4440 (N_4440,N_3919,N_2828);
nor U4441 (N_4441,N_3887,N_2083);
or U4442 (N_4442,N_3842,N_3825);
and U4443 (N_4443,N_3297,N_2734);
nor U4444 (N_4444,N_3747,N_2340);
nand U4445 (N_4445,N_3430,N_3453);
xnor U4446 (N_4446,N_2979,N_2087);
xor U4447 (N_4447,N_3986,N_3974);
nand U4448 (N_4448,N_2753,N_2870);
nor U4449 (N_4449,N_3203,N_2086);
nor U4450 (N_4450,N_2439,N_3834);
nand U4451 (N_4451,N_3102,N_2485);
or U4452 (N_4452,N_2970,N_3286);
or U4453 (N_4453,N_3811,N_2100);
nor U4454 (N_4454,N_3586,N_3949);
or U4455 (N_4455,N_3364,N_2800);
and U4456 (N_4456,N_3617,N_3720);
or U4457 (N_4457,N_3962,N_3644);
nand U4458 (N_4458,N_3064,N_2126);
nor U4459 (N_4459,N_2604,N_2276);
and U4460 (N_4460,N_3398,N_2805);
and U4461 (N_4461,N_2567,N_3406);
xnor U4462 (N_4462,N_2243,N_2730);
or U4463 (N_4463,N_3818,N_3607);
nand U4464 (N_4464,N_2574,N_3114);
xor U4465 (N_4465,N_3169,N_2314);
xor U4466 (N_4466,N_3197,N_3279);
xor U4467 (N_4467,N_3230,N_2689);
and U4468 (N_4468,N_2519,N_3329);
and U4469 (N_4469,N_3874,N_3259);
xnor U4470 (N_4470,N_2939,N_2144);
nand U4471 (N_4471,N_2414,N_3529);
nand U4472 (N_4472,N_2422,N_2168);
or U4473 (N_4473,N_3423,N_3799);
and U4474 (N_4474,N_3276,N_2799);
xnor U4475 (N_4475,N_2797,N_3765);
or U4476 (N_4476,N_3742,N_2301);
and U4477 (N_4477,N_2557,N_2437);
and U4478 (N_4478,N_3854,N_3196);
nor U4479 (N_4479,N_2424,N_3535);
nand U4480 (N_4480,N_3463,N_2467);
nor U4481 (N_4481,N_2202,N_2062);
and U4482 (N_4482,N_3831,N_2670);
nand U4483 (N_4483,N_2174,N_2043);
nand U4484 (N_4484,N_3298,N_3937);
xor U4485 (N_4485,N_2530,N_3176);
xor U4486 (N_4486,N_3433,N_3989);
xnor U4487 (N_4487,N_2055,N_2132);
or U4488 (N_4488,N_3360,N_3130);
xnor U4489 (N_4489,N_2189,N_2363);
and U4490 (N_4490,N_2486,N_3645);
nor U4491 (N_4491,N_2212,N_2741);
nand U4492 (N_4492,N_3723,N_2812);
and U4493 (N_4493,N_3078,N_2093);
xor U4494 (N_4494,N_2533,N_2708);
xnor U4495 (N_4495,N_3775,N_3587);
nand U4496 (N_4496,N_2342,N_2181);
and U4497 (N_4497,N_3195,N_2824);
nand U4498 (N_4498,N_3555,N_3869);
and U4499 (N_4499,N_2754,N_2677);
nand U4500 (N_4500,N_3895,N_2029);
or U4501 (N_4501,N_2382,N_3860);
nor U4502 (N_4502,N_3347,N_3664);
nor U4503 (N_4503,N_3813,N_2794);
or U4504 (N_4504,N_3090,N_2862);
and U4505 (N_4505,N_2565,N_3783);
or U4506 (N_4506,N_3632,N_2182);
nand U4507 (N_4507,N_3669,N_2990);
and U4508 (N_4508,N_3646,N_3296);
xnor U4509 (N_4509,N_2123,N_2780);
nand U4510 (N_4510,N_2435,N_2058);
or U4511 (N_4511,N_3256,N_3294);
and U4512 (N_4512,N_2401,N_2103);
and U4513 (N_4513,N_2415,N_3155);
xnor U4514 (N_4514,N_2917,N_3123);
nor U4515 (N_4515,N_2657,N_2884);
nor U4516 (N_4516,N_3071,N_3875);
and U4517 (N_4517,N_3229,N_3671);
xor U4518 (N_4518,N_2740,N_2236);
or U4519 (N_4519,N_2966,N_2296);
and U4520 (N_4520,N_2695,N_3427);
xnor U4521 (N_4521,N_2395,N_3613);
nand U4522 (N_4522,N_3806,N_2224);
or U4523 (N_4523,N_2786,N_2571);
xor U4524 (N_4524,N_3239,N_3024);
xor U4525 (N_4525,N_2912,N_3913);
nor U4526 (N_4526,N_3888,N_2464);
xnor U4527 (N_4527,N_2995,N_2056);
nand U4528 (N_4528,N_2905,N_3038);
xor U4529 (N_4529,N_2372,N_3500);
nor U4530 (N_4530,N_3034,N_3701);
and U4531 (N_4531,N_3767,N_3104);
nor U4532 (N_4532,N_2449,N_2512);
or U4533 (N_4533,N_2110,N_3419);
xnor U4534 (N_4534,N_2755,N_3255);
or U4535 (N_4535,N_3938,N_3308);
xnor U4536 (N_4536,N_2776,N_3968);
nor U4537 (N_4537,N_3200,N_3426);
xnor U4538 (N_4538,N_3183,N_2318);
nand U4539 (N_4539,N_2465,N_2888);
or U4540 (N_4540,N_3245,N_3348);
nor U4541 (N_4541,N_3127,N_3828);
nor U4542 (N_4542,N_2347,N_3079);
or U4543 (N_4543,N_2063,N_3212);
and U4544 (N_4544,N_3112,N_3044);
or U4545 (N_4545,N_2976,N_3648);
nor U4546 (N_4546,N_2943,N_2205);
and U4547 (N_4547,N_3905,N_2150);
nand U4548 (N_4548,N_3486,N_3247);
xor U4549 (N_4549,N_2721,N_3093);
nand U4550 (N_4550,N_3162,N_3357);
or U4551 (N_4551,N_3077,N_2773);
xnor U4552 (N_4552,N_3791,N_2067);
and U4553 (N_4553,N_2644,N_3411);
or U4554 (N_4554,N_2674,N_2047);
and U4555 (N_4555,N_2611,N_3418);
xnor U4556 (N_4556,N_3194,N_2084);
nand U4557 (N_4557,N_2390,N_3893);
xor U4558 (N_4558,N_3969,N_3650);
and U4559 (N_4559,N_3520,N_2553);
and U4560 (N_4560,N_2944,N_3610);
xor U4561 (N_4561,N_3576,N_2920);
xor U4562 (N_4562,N_3600,N_3116);
nand U4563 (N_4563,N_2954,N_3764);
or U4564 (N_4564,N_2710,N_2842);
xnor U4565 (N_4565,N_3961,N_3006);
xnor U4566 (N_4566,N_2725,N_2069);
nor U4567 (N_4567,N_2416,N_2953);
or U4568 (N_4568,N_3947,N_2514);
nor U4569 (N_4569,N_3710,N_3876);
or U4570 (N_4570,N_3140,N_2450);
and U4571 (N_4571,N_2505,N_3545);
nor U4572 (N_4572,N_2000,N_3707);
and U4573 (N_4573,N_2234,N_2552);
or U4574 (N_4574,N_2051,N_3691);
nand U4575 (N_4575,N_2768,N_3081);
and U4576 (N_4576,N_2339,N_3257);
or U4577 (N_4577,N_3763,N_3375);
and U4578 (N_4578,N_2535,N_3291);
xnor U4579 (N_4579,N_2972,N_3674);
nor U4580 (N_4580,N_3915,N_3862);
nor U4581 (N_4581,N_2659,N_2806);
nor U4582 (N_4582,N_2779,N_3784);
xnor U4583 (N_4583,N_2231,N_2220);
and U4584 (N_4584,N_3086,N_3505);
and U4585 (N_4585,N_3036,N_2962);
or U4586 (N_4586,N_3823,N_3731);
nand U4587 (N_4587,N_3708,N_2281);
nor U4588 (N_4588,N_3143,N_3958);
and U4589 (N_4589,N_2975,N_3070);
or U4590 (N_4590,N_3568,N_3892);
or U4591 (N_4591,N_3117,N_3728);
nand U4592 (N_4592,N_2613,N_3323);
nor U4593 (N_4593,N_2662,N_2716);
xor U4594 (N_4594,N_3240,N_3564);
nand U4595 (N_4595,N_3015,N_2225);
nor U4596 (N_4596,N_3119,N_3981);
xor U4597 (N_4597,N_2457,N_2723);
or U4598 (N_4598,N_2769,N_2898);
or U4599 (N_4599,N_2057,N_2658);
or U4600 (N_4600,N_3786,N_3561);
nand U4601 (N_4601,N_2699,N_3008);
nor U4602 (N_4602,N_3907,N_2240);
and U4603 (N_4603,N_3841,N_3897);
xnor U4604 (N_4604,N_3598,N_3528);
and U4605 (N_4605,N_2818,N_2299);
xor U4606 (N_4606,N_3266,N_3110);
or U4607 (N_4607,N_3556,N_3435);
nor U4608 (N_4608,N_3373,N_2660);
nand U4609 (N_4609,N_3682,N_2104);
and U4610 (N_4610,N_3589,N_2206);
nor U4611 (N_4611,N_2478,N_2358);
nor U4612 (N_4612,N_3817,N_2452);
nand U4613 (N_4613,N_3998,N_2566);
nor U4614 (N_4614,N_2593,N_3802);
nand U4615 (N_4615,N_3124,N_3482);
nor U4616 (N_4616,N_3920,N_3366);
and U4617 (N_4617,N_2254,N_2059);
nand U4618 (N_4618,N_2409,N_2028);
nor U4619 (N_4619,N_3788,N_2682);
nor U4620 (N_4620,N_2185,N_2031);
nor U4621 (N_4621,N_3122,N_2468);
xor U4622 (N_4622,N_2523,N_2848);
xnor U4623 (N_4623,N_2310,N_2923);
nand U4624 (N_4624,N_2894,N_2650);
xor U4625 (N_4625,N_3547,N_2001);
xnor U4626 (N_4626,N_3186,N_2641);
or U4627 (N_4627,N_2355,N_3592);
and U4628 (N_4628,N_3773,N_2238);
and U4629 (N_4629,N_3101,N_2469);
nor U4630 (N_4630,N_2600,N_2170);
xor U4631 (N_4631,N_2438,N_2880);
and U4632 (N_4632,N_3835,N_2016);
xor U4633 (N_4633,N_2949,N_3924);
nor U4634 (N_4634,N_2778,N_2955);
nor U4635 (N_4635,N_3091,N_2330);
xor U4636 (N_4636,N_3804,N_3639);
xor U4637 (N_4637,N_3258,N_3443);
and U4638 (N_4638,N_2392,N_2076);
nand U4639 (N_4639,N_2511,N_3001);
or U4640 (N_4640,N_3917,N_2596);
nor U4641 (N_4641,N_2242,N_2756);
and U4642 (N_4642,N_3579,N_3083);
nor U4643 (N_4643,N_2470,N_3464);
or U4644 (N_4644,N_2383,N_3999);
nand U4645 (N_4645,N_3363,N_2447);
or U4646 (N_4646,N_2893,N_3578);
and U4647 (N_4647,N_2346,N_3076);
and U4648 (N_4648,N_3328,N_2009);
nor U4649 (N_4649,N_2207,N_3724);
nor U4650 (N_4650,N_3930,N_3234);
nor U4651 (N_4651,N_3221,N_3219);
xor U4652 (N_4652,N_2370,N_3770);
or U4653 (N_4653,N_3883,N_3705);
xnor U4654 (N_4654,N_2278,N_3665);
and U4655 (N_4655,N_3852,N_2648);
xor U4656 (N_4656,N_2639,N_3653);
xor U4657 (N_4657,N_2834,N_2223);
nand U4658 (N_4658,N_2607,N_2500);
and U4659 (N_4659,N_2013,N_3795);
nor U4660 (N_4660,N_3713,N_2496);
or U4661 (N_4661,N_2984,N_3588);
and U4662 (N_4662,N_3041,N_2367);
or U4663 (N_4663,N_2899,N_2810);
or U4664 (N_4664,N_3213,N_2520);
or U4665 (N_4665,N_3567,N_3912);
and U4666 (N_4666,N_2529,N_3132);
or U4667 (N_4667,N_3751,N_3054);
and U4668 (N_4668,N_3725,N_3855);
and U4669 (N_4669,N_3965,N_2610);
and U4670 (N_4670,N_3045,N_2900);
nor U4671 (N_4671,N_3978,N_3844);
xor U4672 (N_4672,N_2991,N_2694);
and U4673 (N_4673,N_3342,N_3405);
nand U4674 (N_4674,N_2989,N_2830);
nand U4675 (N_4675,N_2599,N_3438);
xor U4676 (N_4676,N_3235,N_2743);
and U4677 (N_4677,N_3420,N_2547);
or U4678 (N_4678,N_3983,N_3260);
or U4679 (N_4679,N_3487,N_3629);
nor U4680 (N_4680,N_3943,N_2394);
or U4681 (N_4681,N_2672,N_3715);
nor U4682 (N_4682,N_3359,N_2508);
xor U4683 (N_4683,N_2952,N_2973);
nand U4684 (N_4684,N_3080,N_3385);
nand U4685 (N_4685,N_2026,N_3946);
xor U4686 (N_4686,N_3455,N_2802);
or U4687 (N_4687,N_2692,N_2161);
and U4688 (N_4688,N_2405,N_3549);
nor U4689 (N_4689,N_2187,N_3027);
nand U4690 (N_4690,N_3145,N_2446);
xnor U4691 (N_4691,N_3199,N_2109);
and U4692 (N_4692,N_3246,N_3319);
and U4693 (N_4693,N_3018,N_3492);
xor U4694 (N_4694,N_3384,N_2376);
nand U4695 (N_4695,N_3282,N_2388);
nor U4696 (N_4696,N_2864,N_3769);
nand U4697 (N_4697,N_2041,N_2623);
xnor U4698 (N_4698,N_2481,N_2974);
nor U4699 (N_4699,N_3744,N_3636);
and U4700 (N_4700,N_3415,N_3673);
or U4701 (N_4701,N_2837,N_2850);
nor U4702 (N_4702,N_2841,N_3351);
and U4703 (N_4703,N_2528,N_3278);
nor U4704 (N_4704,N_2377,N_2179);
or U4705 (N_4705,N_3205,N_2071);
or U4706 (N_4706,N_2591,N_3918);
xor U4707 (N_4707,N_2387,N_3467);
nand U4708 (N_4708,N_3635,N_3516);
and U4709 (N_4709,N_2764,N_2090);
xor U4710 (N_4710,N_3571,N_2134);
nor U4711 (N_4711,N_3060,N_2162);
or U4712 (N_4712,N_3454,N_3190);
xnor U4713 (N_4713,N_2428,N_2210);
nor U4714 (N_4714,N_3243,N_3836);
and U4715 (N_4715,N_2371,N_2079);
and U4716 (N_4716,N_2352,N_2360);
or U4717 (N_4717,N_3780,N_3144);
nor U4718 (N_4718,N_2241,N_2827);
nor U4719 (N_4719,N_3304,N_3052);
xnor U4720 (N_4720,N_2661,N_2262);
and U4721 (N_4721,N_3161,N_2305);
or U4722 (N_4722,N_3481,N_3809);
xnor U4723 (N_4723,N_2147,N_2329);
nor U4724 (N_4724,N_3460,N_3530);
or U4725 (N_4725,N_3484,N_3573);
nor U4726 (N_4726,N_2518,N_2700);
nand U4727 (N_4727,N_3009,N_3514);
nor U4728 (N_4728,N_2490,N_2631);
nand U4729 (N_4729,N_3685,N_2183);
xnor U4730 (N_4730,N_3582,N_2101);
nand U4731 (N_4731,N_2758,N_2647);
or U4732 (N_4732,N_2229,N_2760);
xnor U4733 (N_4733,N_2843,N_2883);
xor U4734 (N_4734,N_3964,N_3106);
xnor U4735 (N_4735,N_2784,N_3726);
nor U4736 (N_4736,N_3188,N_2471);
xnor U4737 (N_4737,N_3386,N_3618);
nor U4738 (N_4738,N_2044,N_3274);
and U4739 (N_4739,N_2909,N_3217);
and U4740 (N_4740,N_3168,N_3873);
xnor U4741 (N_4741,N_3693,N_3377);
nand U4742 (N_4742,N_3350,N_2221);
nand U4743 (N_4743,N_3238,N_3232);
nor U4744 (N_4744,N_2940,N_2938);
and U4745 (N_4745,N_3890,N_3156);
nor U4746 (N_4746,N_2537,N_3466);
nor U4747 (N_4747,N_2885,N_3179);
nor U4748 (N_4748,N_2625,N_3634);
nand U4749 (N_4749,N_2257,N_2983);
nor U4750 (N_4750,N_2328,N_3220);
and U4751 (N_4751,N_3971,N_3448);
and U4752 (N_4752,N_3309,N_2928);
nor U4753 (N_4753,N_2892,N_3236);
xor U4754 (N_4754,N_2386,N_2522);
nand U4755 (N_4755,N_2213,N_3850);
nor U4756 (N_4756,N_3688,N_3536);
nor U4757 (N_4757,N_3790,N_3758);
xnor U4758 (N_4758,N_2521,N_3801);
xor U4759 (N_4759,N_3771,N_2173);
xnor U4760 (N_4760,N_3468,N_2252);
and U4761 (N_4761,N_3272,N_2922);
nor U4762 (N_4762,N_3192,N_3882);
xnor U4763 (N_4763,N_3846,N_2443);
or U4764 (N_4764,N_3031,N_2307);
xor U4765 (N_4765,N_2745,N_2717);
nand U4766 (N_4766,N_3729,N_2267);
xor U4767 (N_4767,N_2232,N_3152);
nor U4768 (N_4768,N_2931,N_2731);
or U4769 (N_4769,N_2792,N_3572);
nand U4770 (N_4770,N_2145,N_3380);
nor U4771 (N_4771,N_3289,N_3025);
xor U4772 (N_4772,N_3660,N_3973);
or U4773 (N_4773,N_2994,N_2164);
and U4774 (N_4774,N_3789,N_3524);
or U4775 (N_4775,N_2433,N_2149);
or U4776 (N_4776,N_2936,N_3712);
nand U4777 (N_4777,N_2477,N_2951);
or U4778 (N_4778,N_2788,N_3703);
xnor U4779 (N_4779,N_2253,N_2379);
xnor U4780 (N_4780,N_2440,N_3911);
nand U4781 (N_4781,N_2040,N_3173);
or U4782 (N_4782,N_3072,N_3637);
nor U4783 (N_4783,N_2882,N_3180);
or U4784 (N_4784,N_3367,N_3916);
nor U4785 (N_4785,N_2578,N_3471);
and U4786 (N_4786,N_3585,N_2675);
nand U4787 (N_4787,N_3181,N_2397);
or U4788 (N_4788,N_3303,N_3111);
nor U4789 (N_4789,N_3877,N_2430);
xor U4790 (N_4790,N_2866,N_2258);
nand U4791 (N_4791,N_2476,N_3461);
xnor U4792 (N_4792,N_2619,N_2517);
nor U4793 (N_4793,N_3288,N_3227);
nor U4794 (N_4794,N_2865,N_2211);
and U4795 (N_4795,N_2997,N_3955);
or U4796 (N_4796,N_2685,N_2646);
or U4797 (N_4797,N_3053,N_3157);
xor U4798 (N_4798,N_3595,N_3865);
or U4799 (N_4799,N_3108,N_3566);
or U4800 (N_4800,N_2683,N_3857);
xor U4801 (N_4801,N_2902,N_3320);
or U4802 (N_4802,N_2879,N_2158);
or U4803 (N_4803,N_2618,N_3402);
nor U4804 (N_4804,N_2747,N_3531);
and U4805 (N_4805,N_3941,N_3540);
nor U4806 (N_4806,N_2612,N_3807);
xor U4807 (N_4807,N_2396,N_2759);
nand U4808 (N_4808,N_3332,N_2643);
nor U4809 (N_4809,N_2620,N_3341);
and U4810 (N_4810,N_2484,N_2313);
xnor U4811 (N_4811,N_2977,N_2742);
or U4812 (N_4812,N_2653,N_3749);
or U4813 (N_4813,N_3021,N_3142);
nand U4814 (N_4814,N_2226,N_2908);
xor U4815 (N_4815,N_3711,N_2543);
and U4816 (N_4816,N_2546,N_2431);
nor U4817 (N_4817,N_2761,N_2506);
nor U4818 (N_4818,N_3337,N_2577);
nor U4819 (N_4819,N_3515,N_3316);
nor U4820 (N_4820,N_3491,N_2280);
and U4821 (N_4821,N_3820,N_2783);
nand U4822 (N_4822,N_3668,N_3226);
nor U4823 (N_4823,N_3250,N_3224);
xnor U4824 (N_4824,N_2832,N_3368);
nand U4825 (N_4825,N_3739,N_3891);
or U4826 (N_4826,N_2538,N_3470);
nand U4827 (N_4827,N_3311,N_2516);
and U4828 (N_4828,N_2697,N_2726);
nor U4829 (N_4829,N_3331,N_2559);
or U4830 (N_4830,N_3136,N_3148);
and U4831 (N_4831,N_2050,N_2774);
xnor U4832 (N_4832,N_3019,N_2605);
or U4833 (N_4833,N_2306,N_2419);
nor U4834 (N_4834,N_3182,N_3126);
xnor U4835 (N_4835,N_2652,N_2230);
nand U4836 (N_4836,N_3002,N_3075);
nand U4837 (N_4837,N_2531,N_2244);
nand U4838 (N_4838,N_2904,N_3388);
and U4839 (N_4839,N_3886,N_3812);
nand U4840 (N_4840,N_2988,N_3358);
nand U4841 (N_4841,N_3191,N_3672);
and U4842 (N_4842,N_2819,N_3285);
nor U4843 (N_4843,N_2462,N_3084);
or U4844 (N_4844,N_3743,N_2713);
xor U4845 (N_4845,N_2052,N_3030);
and U4846 (N_4846,N_2615,N_2003);
nand U4847 (N_4847,N_2696,N_3593);
xor U4848 (N_4848,N_2480,N_2545);
or U4849 (N_4849,N_3089,N_2341);
and U4850 (N_4850,N_2070,N_2608);
nor U4851 (N_4851,N_2172,N_3063);
xor U4852 (N_4852,N_3208,N_2322);
xor U4853 (N_4853,N_2916,N_3447);
nand U4854 (N_4854,N_3642,N_2078);
xnor U4855 (N_4855,N_2548,N_2957);
nand U4856 (N_4856,N_3872,N_2188);
xnor U4857 (N_4857,N_3657,N_2664);
nor U4858 (N_4858,N_3040,N_3051);
xor U4859 (N_4859,N_2836,N_3628);
or U4860 (N_4860,N_2348,N_2572);
and U4861 (N_4861,N_3202,N_2297);
xnor U4862 (N_4862,N_2045,N_2671);
or U4863 (N_4863,N_2873,N_2791);
and U4864 (N_4864,N_3880,N_3164);
or U4865 (N_4865,N_2727,N_2630);
nand U4866 (N_4866,N_3945,N_2105);
nand U4867 (N_4867,N_2587,N_2942);
or U4868 (N_4868,N_3858,N_2068);
nand U4869 (N_4869,N_3800,N_3017);
and U4870 (N_4870,N_3754,N_3906);
nand U4871 (N_4871,N_3927,N_3244);
or U4872 (N_4872,N_3425,N_2064);
xnor U4873 (N_4873,N_3151,N_3899);
nand U4874 (N_4874,N_3248,N_3378);
and U4875 (N_4875,N_2886,N_3098);
xor U4876 (N_4876,N_2728,N_2851);
nand U4877 (N_4877,N_3353,N_3980);
nor U4878 (N_4878,N_2228,N_3939);
nand U4879 (N_4879,N_3280,N_3987);
or U4880 (N_4880,N_3407,N_2049);
and U4881 (N_4881,N_2354,N_2590);
xor U4882 (N_4882,N_2368,N_3953);
nand U4883 (N_4883,N_2198,N_2154);
or U4884 (N_4884,N_3313,N_2863);
nand U4885 (N_4885,N_2825,N_3900);
nand U4886 (N_4886,N_2736,N_2636);
xor U4887 (N_4887,N_3879,N_3210);
nand U4888 (N_4888,N_3631,N_3483);
nor U4889 (N_4889,N_3542,N_2131);
nand U4890 (N_4890,N_2927,N_2501);
or U4891 (N_4891,N_2037,N_2042);
nor U4892 (N_4892,N_3334,N_2351);
nor U4893 (N_4893,N_2255,N_2264);
or U4894 (N_4894,N_2380,N_3035);
or U4895 (N_4895,N_3047,N_2640);
nor U4896 (N_4896,N_3521,N_2752);
nor U4897 (N_4897,N_3736,N_2120);
xor U4898 (N_4898,N_2381,N_3149);
xor U4899 (N_4899,N_2877,N_2142);
nand U4900 (N_4900,N_3667,N_2349);
and U4901 (N_4901,N_3661,N_2273);
xnor U4902 (N_4902,N_3552,N_3431);
nand U4903 (N_4903,N_3761,N_2787);
nand U4904 (N_4904,N_3413,N_3581);
and U4905 (N_4905,N_3277,N_2408);
xnor U4906 (N_4906,N_3753,N_3678);
nand U4907 (N_4907,N_2687,N_2293);
or U4908 (N_4908,N_3033,N_3022);
nand U4909 (N_4909,N_3518,N_3928);
or U4910 (N_4910,N_3734,N_2418);
nor U4911 (N_4911,N_2369,N_2053);
nand U4912 (N_4912,N_2410,N_2637);
xor U4913 (N_4913,N_2364,N_3295);
xor U4914 (N_4914,N_2233,N_2463);
and U4915 (N_4915,N_3253,N_2474);
nand U4916 (N_4916,N_2406,N_3692);
nor U4917 (N_4917,N_3884,N_3510);
and U4918 (N_4918,N_3473,N_2771);
and U4919 (N_4919,N_2385,N_2621);
and U4920 (N_4920,N_3594,N_2094);
xor U4921 (N_4921,N_3508,N_2632);
and U4922 (N_4922,N_2292,N_3109);
or U4923 (N_4923,N_2793,N_3193);
nor U4924 (N_4924,N_3343,N_2679);
xnor U4925 (N_4925,N_3171,N_2426);
and U4926 (N_4926,N_3020,N_3861);
nand U4927 (N_4927,N_2617,N_2624);
or U4928 (N_4928,N_2361,N_2215);
and U4929 (N_4929,N_2184,N_3275);
and U4930 (N_4930,N_2260,N_3312);
xor U4931 (N_4931,N_3694,N_3087);
xnor U4932 (N_4932,N_3853,N_3488);
or U4933 (N_4933,N_2744,N_2584);
nand U4934 (N_4934,N_3591,N_3026);
or U4935 (N_4935,N_3627,N_3766);
xnor U4936 (N_4936,N_2606,N_3957);
and U4937 (N_4937,N_2300,N_3493);
nand U4938 (N_4938,N_2160,N_3611);
and U4939 (N_4939,N_2558,N_2429);
nand U4940 (N_4940,N_2095,N_2021);
or U4941 (N_4941,N_3394,N_3273);
or U4942 (N_4942,N_2146,N_3096);
nor U4943 (N_4943,N_2513,N_2080);
xor U4944 (N_4944,N_2061,N_2116);
or U4945 (N_4945,N_3376,N_2171);
xor U4946 (N_4946,N_3601,N_2586);
nand U4947 (N_4947,N_3159,N_2628);
nor U4948 (N_4948,N_3896,N_3354);
nor U4949 (N_4949,N_3344,N_2107);
nand U4950 (N_4950,N_3166,N_3615);
and U4951 (N_4951,N_2291,N_3690);
xnor U4952 (N_4952,N_2407,N_3434);
or U4953 (N_4953,N_3451,N_2811);
and U4954 (N_4954,N_3092,N_3676);
and U4955 (N_4955,N_2066,N_3016);
xor U4956 (N_4956,N_3553,N_2562);
and U4957 (N_4957,N_2456,N_2739);
nor U4958 (N_4958,N_3165,N_3456);
xnor U4959 (N_4959,N_3563,N_2271);
nand U4960 (N_4960,N_3437,N_2237);
and U4961 (N_4961,N_3651,N_2091);
or U4962 (N_4962,N_3321,N_3901);
xor U4963 (N_4963,N_2965,N_2282);
nand U4964 (N_4964,N_3699,N_3851);
or U4965 (N_4965,N_2020,N_3830);
nand U4966 (N_4966,N_3048,N_3714);
xnor U4967 (N_4967,N_3424,N_2711);
and U4968 (N_4968,N_2889,N_2934);
nand U4969 (N_4969,N_2629,N_3746);
xnor U4970 (N_4970,N_3477,N_2594);
and U4971 (N_4971,N_3241,N_2498);
xor U4972 (N_4972,N_2924,N_3267);
and U4973 (N_4973,N_2133,N_3840);
and U4974 (N_4974,N_3000,N_2453);
and U4975 (N_4975,N_3963,N_3498);
or U4976 (N_4976,N_3738,N_2678);
and U4977 (N_4977,N_3095,N_2166);
or U4978 (N_4978,N_2423,N_3922);
and U4979 (N_4979,N_2603,N_3472);
nand U4980 (N_4980,N_2295,N_3067);
xor U4981 (N_4981,N_3154,N_2315);
nor U4982 (N_4982,N_3604,N_3371);
xor U4983 (N_4983,N_2311,N_2869);
nand U4984 (N_4984,N_3519,N_2732);
xor U4985 (N_4985,N_2915,N_2891);
nor U4986 (N_4986,N_3509,N_3982);
nand U4987 (N_4987,N_2176,N_2336);
or U4988 (N_4988,N_2560,N_3372);
nand U4989 (N_4989,N_2308,N_3798);
and U4990 (N_4990,N_3082,N_2616);
nor U4991 (N_4991,N_3984,N_3439);
and U4992 (N_4992,N_2081,N_2155);
xor U4993 (N_4993,N_3570,N_2312);
and U4994 (N_4994,N_2102,N_2268);
xor U4995 (N_4995,N_3755,N_3327);
nor U4996 (N_4996,N_2855,N_3393);
nor U4997 (N_4997,N_3827,N_2399);
nor U4998 (N_4998,N_3979,N_3625);
nand U4999 (N_4999,N_3014,N_2585);
nand U5000 (N_5000,N_3019,N_2501);
and U5001 (N_5001,N_3022,N_3211);
nor U5002 (N_5002,N_2847,N_3561);
nor U5003 (N_5003,N_2261,N_2615);
and U5004 (N_5004,N_2638,N_2092);
or U5005 (N_5005,N_2970,N_2452);
nand U5006 (N_5006,N_3568,N_3849);
and U5007 (N_5007,N_3822,N_2855);
xnor U5008 (N_5008,N_2204,N_2102);
and U5009 (N_5009,N_3959,N_2076);
nand U5010 (N_5010,N_2110,N_3575);
nand U5011 (N_5011,N_3451,N_2068);
and U5012 (N_5012,N_2227,N_3715);
and U5013 (N_5013,N_3162,N_2370);
xnor U5014 (N_5014,N_3766,N_3850);
xor U5015 (N_5015,N_3991,N_3825);
nand U5016 (N_5016,N_3452,N_2411);
or U5017 (N_5017,N_3062,N_3832);
nand U5018 (N_5018,N_2324,N_3583);
xor U5019 (N_5019,N_3578,N_2913);
and U5020 (N_5020,N_3890,N_3472);
nor U5021 (N_5021,N_3599,N_3805);
or U5022 (N_5022,N_3485,N_3546);
and U5023 (N_5023,N_3648,N_3975);
nor U5024 (N_5024,N_3179,N_2594);
nor U5025 (N_5025,N_2926,N_3659);
nor U5026 (N_5026,N_3390,N_2383);
or U5027 (N_5027,N_3178,N_3835);
nand U5028 (N_5028,N_3897,N_2333);
nand U5029 (N_5029,N_3815,N_2703);
xor U5030 (N_5030,N_2122,N_2212);
nor U5031 (N_5031,N_3446,N_2370);
xor U5032 (N_5032,N_3930,N_2484);
nand U5033 (N_5033,N_2119,N_3676);
nor U5034 (N_5034,N_3678,N_3376);
xnor U5035 (N_5035,N_2316,N_3902);
nor U5036 (N_5036,N_2665,N_3975);
nor U5037 (N_5037,N_2141,N_3627);
xnor U5038 (N_5038,N_2733,N_3077);
xor U5039 (N_5039,N_3695,N_3657);
or U5040 (N_5040,N_3796,N_2908);
and U5041 (N_5041,N_2180,N_3033);
or U5042 (N_5042,N_2633,N_3358);
or U5043 (N_5043,N_2810,N_3960);
nor U5044 (N_5044,N_2265,N_3924);
and U5045 (N_5045,N_2993,N_3878);
or U5046 (N_5046,N_2926,N_3575);
or U5047 (N_5047,N_2147,N_2674);
and U5048 (N_5048,N_3138,N_2992);
xor U5049 (N_5049,N_2485,N_3348);
nor U5050 (N_5050,N_3486,N_2227);
nor U5051 (N_5051,N_3324,N_2382);
xnor U5052 (N_5052,N_3387,N_3683);
nor U5053 (N_5053,N_3032,N_2553);
xnor U5054 (N_5054,N_2082,N_2948);
and U5055 (N_5055,N_3545,N_3306);
or U5056 (N_5056,N_2187,N_2092);
nor U5057 (N_5057,N_2819,N_2527);
nor U5058 (N_5058,N_2388,N_2536);
xor U5059 (N_5059,N_3337,N_3001);
nand U5060 (N_5060,N_2410,N_3559);
nor U5061 (N_5061,N_3679,N_2587);
xor U5062 (N_5062,N_3551,N_3450);
or U5063 (N_5063,N_2942,N_2004);
xnor U5064 (N_5064,N_2919,N_3750);
nand U5065 (N_5065,N_3503,N_2098);
nand U5066 (N_5066,N_3331,N_3512);
nor U5067 (N_5067,N_2073,N_3130);
xor U5068 (N_5068,N_3142,N_2960);
nor U5069 (N_5069,N_3273,N_3136);
xor U5070 (N_5070,N_3530,N_2628);
nand U5071 (N_5071,N_3481,N_2413);
and U5072 (N_5072,N_3481,N_2308);
nand U5073 (N_5073,N_2605,N_2264);
nor U5074 (N_5074,N_2573,N_2331);
nor U5075 (N_5075,N_3240,N_3284);
xnor U5076 (N_5076,N_2823,N_3074);
nand U5077 (N_5077,N_2748,N_3193);
nand U5078 (N_5078,N_3390,N_3849);
nand U5079 (N_5079,N_3188,N_2247);
nor U5080 (N_5080,N_3441,N_3392);
and U5081 (N_5081,N_3206,N_2161);
nand U5082 (N_5082,N_3503,N_3831);
nor U5083 (N_5083,N_2973,N_3253);
nor U5084 (N_5084,N_2094,N_2578);
nor U5085 (N_5085,N_3716,N_2096);
xnor U5086 (N_5086,N_3086,N_2061);
or U5087 (N_5087,N_3021,N_2928);
nor U5088 (N_5088,N_2667,N_3671);
xor U5089 (N_5089,N_2028,N_2657);
xor U5090 (N_5090,N_2029,N_2432);
nand U5091 (N_5091,N_2130,N_2815);
and U5092 (N_5092,N_3107,N_2590);
xnor U5093 (N_5093,N_2970,N_3248);
xnor U5094 (N_5094,N_2777,N_3884);
xor U5095 (N_5095,N_2627,N_2805);
nor U5096 (N_5096,N_2698,N_3683);
xnor U5097 (N_5097,N_2952,N_3270);
nand U5098 (N_5098,N_2200,N_3291);
or U5099 (N_5099,N_3212,N_3602);
nor U5100 (N_5100,N_3797,N_3923);
nand U5101 (N_5101,N_3325,N_2322);
or U5102 (N_5102,N_2599,N_2086);
xor U5103 (N_5103,N_2388,N_2526);
or U5104 (N_5104,N_3516,N_2690);
nor U5105 (N_5105,N_2050,N_2522);
or U5106 (N_5106,N_2262,N_3641);
or U5107 (N_5107,N_2924,N_2168);
nor U5108 (N_5108,N_2194,N_3729);
xor U5109 (N_5109,N_2862,N_2633);
xnor U5110 (N_5110,N_2846,N_3233);
xnor U5111 (N_5111,N_2315,N_2398);
or U5112 (N_5112,N_3960,N_3007);
xnor U5113 (N_5113,N_3236,N_3810);
or U5114 (N_5114,N_3692,N_2104);
nand U5115 (N_5115,N_3764,N_2103);
nor U5116 (N_5116,N_2760,N_3699);
xnor U5117 (N_5117,N_2282,N_3565);
xnor U5118 (N_5118,N_2289,N_2787);
nand U5119 (N_5119,N_2727,N_3232);
nand U5120 (N_5120,N_3743,N_3704);
and U5121 (N_5121,N_3420,N_3390);
and U5122 (N_5122,N_2649,N_2662);
and U5123 (N_5123,N_3129,N_3108);
xor U5124 (N_5124,N_3466,N_3340);
or U5125 (N_5125,N_2217,N_3455);
xor U5126 (N_5126,N_2933,N_3934);
and U5127 (N_5127,N_2370,N_3544);
nor U5128 (N_5128,N_3988,N_2808);
or U5129 (N_5129,N_3651,N_2531);
and U5130 (N_5130,N_3782,N_2160);
xor U5131 (N_5131,N_3339,N_3996);
nor U5132 (N_5132,N_3228,N_2306);
nand U5133 (N_5133,N_2165,N_2810);
and U5134 (N_5134,N_2844,N_2291);
nand U5135 (N_5135,N_3657,N_2421);
nand U5136 (N_5136,N_2079,N_3493);
nor U5137 (N_5137,N_3439,N_2740);
nand U5138 (N_5138,N_2467,N_3964);
xor U5139 (N_5139,N_2240,N_3115);
nand U5140 (N_5140,N_3603,N_2471);
and U5141 (N_5141,N_3242,N_2531);
or U5142 (N_5142,N_2924,N_2853);
and U5143 (N_5143,N_2540,N_3284);
nand U5144 (N_5144,N_3013,N_3368);
xnor U5145 (N_5145,N_2392,N_3672);
nand U5146 (N_5146,N_2863,N_2948);
nor U5147 (N_5147,N_2387,N_3617);
nand U5148 (N_5148,N_3153,N_3497);
xnor U5149 (N_5149,N_3895,N_2984);
xnor U5150 (N_5150,N_2760,N_2779);
xnor U5151 (N_5151,N_3901,N_3227);
and U5152 (N_5152,N_3284,N_3740);
xor U5153 (N_5153,N_2091,N_3279);
nor U5154 (N_5154,N_2723,N_3516);
nand U5155 (N_5155,N_3611,N_2334);
nor U5156 (N_5156,N_2565,N_3233);
or U5157 (N_5157,N_3632,N_2304);
nand U5158 (N_5158,N_2125,N_2065);
or U5159 (N_5159,N_3677,N_2436);
or U5160 (N_5160,N_2636,N_3018);
or U5161 (N_5161,N_2898,N_2304);
and U5162 (N_5162,N_3527,N_3931);
xnor U5163 (N_5163,N_3102,N_3900);
nand U5164 (N_5164,N_2900,N_3245);
or U5165 (N_5165,N_2958,N_3775);
xnor U5166 (N_5166,N_2812,N_3625);
and U5167 (N_5167,N_3733,N_3105);
nor U5168 (N_5168,N_2093,N_2631);
and U5169 (N_5169,N_2080,N_3604);
nor U5170 (N_5170,N_2697,N_3105);
xnor U5171 (N_5171,N_3851,N_2810);
xor U5172 (N_5172,N_2028,N_3338);
xnor U5173 (N_5173,N_3462,N_2908);
nand U5174 (N_5174,N_2766,N_2733);
and U5175 (N_5175,N_2484,N_2717);
nand U5176 (N_5176,N_3474,N_2035);
and U5177 (N_5177,N_2131,N_2049);
nor U5178 (N_5178,N_3189,N_2934);
or U5179 (N_5179,N_3402,N_2724);
nand U5180 (N_5180,N_3991,N_2600);
nand U5181 (N_5181,N_3559,N_2879);
nand U5182 (N_5182,N_2890,N_2123);
nand U5183 (N_5183,N_3860,N_2249);
or U5184 (N_5184,N_2117,N_2583);
nand U5185 (N_5185,N_2684,N_3176);
and U5186 (N_5186,N_2675,N_3423);
nor U5187 (N_5187,N_3015,N_3792);
nor U5188 (N_5188,N_3368,N_3634);
xor U5189 (N_5189,N_2950,N_2575);
nor U5190 (N_5190,N_3140,N_2788);
nor U5191 (N_5191,N_3667,N_3062);
or U5192 (N_5192,N_2344,N_2909);
nor U5193 (N_5193,N_2047,N_2113);
nor U5194 (N_5194,N_2220,N_2132);
and U5195 (N_5195,N_3013,N_3383);
or U5196 (N_5196,N_2662,N_3792);
xnor U5197 (N_5197,N_2212,N_3426);
nand U5198 (N_5198,N_2877,N_3119);
xnor U5199 (N_5199,N_2484,N_3348);
xnor U5200 (N_5200,N_2077,N_3656);
nor U5201 (N_5201,N_3026,N_3614);
nand U5202 (N_5202,N_2243,N_2987);
and U5203 (N_5203,N_3961,N_3795);
nand U5204 (N_5204,N_3586,N_3027);
or U5205 (N_5205,N_2821,N_2835);
or U5206 (N_5206,N_2633,N_2807);
xnor U5207 (N_5207,N_2194,N_3911);
nand U5208 (N_5208,N_2127,N_3083);
nand U5209 (N_5209,N_2903,N_3957);
or U5210 (N_5210,N_3012,N_2436);
or U5211 (N_5211,N_2517,N_3866);
xor U5212 (N_5212,N_3839,N_2628);
nor U5213 (N_5213,N_2245,N_3355);
xor U5214 (N_5214,N_2169,N_2683);
nor U5215 (N_5215,N_3287,N_3049);
and U5216 (N_5216,N_2602,N_2561);
xnor U5217 (N_5217,N_3431,N_3144);
nor U5218 (N_5218,N_3567,N_3921);
xnor U5219 (N_5219,N_3979,N_3398);
nor U5220 (N_5220,N_2964,N_2681);
nand U5221 (N_5221,N_2021,N_2730);
and U5222 (N_5222,N_3718,N_2512);
xor U5223 (N_5223,N_3072,N_3356);
nor U5224 (N_5224,N_2547,N_2136);
and U5225 (N_5225,N_3860,N_2034);
nor U5226 (N_5226,N_2270,N_2709);
nor U5227 (N_5227,N_3629,N_3137);
xor U5228 (N_5228,N_2479,N_3135);
and U5229 (N_5229,N_3548,N_2875);
nor U5230 (N_5230,N_3309,N_2102);
and U5231 (N_5231,N_2248,N_2939);
xnor U5232 (N_5232,N_2943,N_2179);
and U5233 (N_5233,N_2767,N_2562);
nand U5234 (N_5234,N_2155,N_2931);
nor U5235 (N_5235,N_2919,N_2110);
xnor U5236 (N_5236,N_2095,N_3028);
xnor U5237 (N_5237,N_3819,N_2691);
xnor U5238 (N_5238,N_2908,N_3718);
and U5239 (N_5239,N_2525,N_3150);
nor U5240 (N_5240,N_3208,N_3083);
and U5241 (N_5241,N_3593,N_3763);
and U5242 (N_5242,N_2122,N_3775);
nor U5243 (N_5243,N_3889,N_2930);
nand U5244 (N_5244,N_3518,N_3320);
nor U5245 (N_5245,N_2479,N_3806);
nand U5246 (N_5246,N_3757,N_3106);
xnor U5247 (N_5247,N_3399,N_2559);
xor U5248 (N_5248,N_3212,N_3245);
or U5249 (N_5249,N_3372,N_2729);
or U5250 (N_5250,N_3981,N_3319);
nor U5251 (N_5251,N_3830,N_2358);
and U5252 (N_5252,N_3442,N_2850);
and U5253 (N_5253,N_3740,N_3812);
or U5254 (N_5254,N_3180,N_2225);
or U5255 (N_5255,N_3928,N_2369);
nand U5256 (N_5256,N_3753,N_2641);
xnor U5257 (N_5257,N_3348,N_3805);
xor U5258 (N_5258,N_3536,N_3257);
nand U5259 (N_5259,N_2649,N_2582);
nor U5260 (N_5260,N_3476,N_3883);
or U5261 (N_5261,N_3398,N_3331);
and U5262 (N_5262,N_2625,N_3490);
and U5263 (N_5263,N_3403,N_3565);
nor U5264 (N_5264,N_2844,N_3615);
xor U5265 (N_5265,N_2739,N_2836);
and U5266 (N_5266,N_2431,N_2012);
or U5267 (N_5267,N_2961,N_3235);
nor U5268 (N_5268,N_3844,N_2022);
or U5269 (N_5269,N_2008,N_3475);
nand U5270 (N_5270,N_3020,N_3285);
nand U5271 (N_5271,N_3972,N_3648);
xnor U5272 (N_5272,N_2511,N_2238);
or U5273 (N_5273,N_2468,N_2941);
and U5274 (N_5274,N_3022,N_3214);
nor U5275 (N_5275,N_3415,N_2058);
nor U5276 (N_5276,N_2056,N_2878);
nand U5277 (N_5277,N_2997,N_2903);
and U5278 (N_5278,N_2509,N_3876);
nor U5279 (N_5279,N_3397,N_2008);
or U5280 (N_5280,N_3784,N_3464);
and U5281 (N_5281,N_2230,N_2464);
and U5282 (N_5282,N_2590,N_2449);
and U5283 (N_5283,N_2892,N_2161);
or U5284 (N_5284,N_2816,N_3240);
nor U5285 (N_5285,N_2295,N_3231);
nor U5286 (N_5286,N_2122,N_2636);
and U5287 (N_5287,N_2040,N_3945);
and U5288 (N_5288,N_3858,N_3186);
nor U5289 (N_5289,N_3554,N_3375);
nand U5290 (N_5290,N_2400,N_2061);
or U5291 (N_5291,N_2118,N_2399);
and U5292 (N_5292,N_2432,N_3828);
nor U5293 (N_5293,N_3557,N_2059);
nor U5294 (N_5294,N_3949,N_2585);
nor U5295 (N_5295,N_2919,N_3863);
nor U5296 (N_5296,N_3200,N_2793);
or U5297 (N_5297,N_2002,N_2937);
or U5298 (N_5298,N_3981,N_3670);
or U5299 (N_5299,N_3666,N_2115);
or U5300 (N_5300,N_2202,N_3883);
nor U5301 (N_5301,N_2871,N_2944);
or U5302 (N_5302,N_3733,N_2550);
xor U5303 (N_5303,N_3049,N_3591);
and U5304 (N_5304,N_2293,N_2511);
and U5305 (N_5305,N_2620,N_2042);
nand U5306 (N_5306,N_2548,N_3028);
nor U5307 (N_5307,N_3880,N_3959);
nand U5308 (N_5308,N_2606,N_2158);
nand U5309 (N_5309,N_3850,N_3893);
or U5310 (N_5310,N_2149,N_2041);
xnor U5311 (N_5311,N_3754,N_3309);
or U5312 (N_5312,N_2266,N_3555);
nand U5313 (N_5313,N_2896,N_3992);
and U5314 (N_5314,N_2537,N_2603);
and U5315 (N_5315,N_3573,N_2958);
xnor U5316 (N_5316,N_2782,N_2444);
xnor U5317 (N_5317,N_3173,N_2577);
xor U5318 (N_5318,N_2346,N_2647);
nand U5319 (N_5319,N_3438,N_3217);
and U5320 (N_5320,N_2440,N_2191);
or U5321 (N_5321,N_3244,N_3209);
nor U5322 (N_5322,N_2392,N_2341);
xnor U5323 (N_5323,N_3492,N_2972);
and U5324 (N_5324,N_3298,N_2609);
nor U5325 (N_5325,N_3910,N_2309);
or U5326 (N_5326,N_3493,N_3511);
and U5327 (N_5327,N_2996,N_3336);
or U5328 (N_5328,N_2821,N_3579);
and U5329 (N_5329,N_3887,N_2957);
and U5330 (N_5330,N_2721,N_2210);
and U5331 (N_5331,N_2309,N_2289);
nand U5332 (N_5332,N_2058,N_2756);
nor U5333 (N_5333,N_3032,N_3380);
nor U5334 (N_5334,N_3891,N_3817);
xor U5335 (N_5335,N_3452,N_3554);
xnor U5336 (N_5336,N_3188,N_3045);
nor U5337 (N_5337,N_3685,N_3299);
and U5338 (N_5338,N_2007,N_2564);
nor U5339 (N_5339,N_2112,N_2783);
and U5340 (N_5340,N_2216,N_2834);
and U5341 (N_5341,N_3062,N_3189);
nor U5342 (N_5342,N_2368,N_2783);
and U5343 (N_5343,N_2510,N_2692);
nor U5344 (N_5344,N_3566,N_3913);
or U5345 (N_5345,N_2372,N_2482);
nor U5346 (N_5346,N_3481,N_3055);
or U5347 (N_5347,N_3249,N_3585);
xnor U5348 (N_5348,N_3122,N_3766);
or U5349 (N_5349,N_2636,N_2851);
and U5350 (N_5350,N_3623,N_3788);
nor U5351 (N_5351,N_2962,N_2512);
or U5352 (N_5352,N_2388,N_2194);
nand U5353 (N_5353,N_2752,N_2444);
and U5354 (N_5354,N_2432,N_2257);
xnor U5355 (N_5355,N_3054,N_3112);
or U5356 (N_5356,N_3171,N_2436);
nor U5357 (N_5357,N_3228,N_2061);
and U5358 (N_5358,N_3292,N_3517);
or U5359 (N_5359,N_2662,N_3659);
nand U5360 (N_5360,N_2767,N_2187);
and U5361 (N_5361,N_3936,N_3816);
xor U5362 (N_5362,N_2580,N_2376);
nand U5363 (N_5363,N_3153,N_3639);
nor U5364 (N_5364,N_2918,N_3668);
or U5365 (N_5365,N_2914,N_3167);
nand U5366 (N_5366,N_2424,N_2847);
nand U5367 (N_5367,N_2205,N_2174);
nor U5368 (N_5368,N_2432,N_2548);
xor U5369 (N_5369,N_2597,N_3516);
nor U5370 (N_5370,N_2991,N_3366);
and U5371 (N_5371,N_2277,N_2572);
and U5372 (N_5372,N_3112,N_3643);
nand U5373 (N_5373,N_2553,N_2192);
or U5374 (N_5374,N_3292,N_2361);
xor U5375 (N_5375,N_3539,N_3642);
nand U5376 (N_5376,N_2626,N_3278);
nand U5377 (N_5377,N_3330,N_2222);
xnor U5378 (N_5378,N_2018,N_3694);
and U5379 (N_5379,N_3076,N_3586);
or U5380 (N_5380,N_2290,N_3315);
and U5381 (N_5381,N_3253,N_3403);
nor U5382 (N_5382,N_3435,N_2623);
nor U5383 (N_5383,N_3587,N_3290);
or U5384 (N_5384,N_2299,N_2272);
or U5385 (N_5385,N_2658,N_2767);
or U5386 (N_5386,N_2788,N_3786);
and U5387 (N_5387,N_2182,N_2213);
and U5388 (N_5388,N_3321,N_3328);
xor U5389 (N_5389,N_3656,N_2768);
xor U5390 (N_5390,N_2320,N_2075);
nand U5391 (N_5391,N_2097,N_3415);
nand U5392 (N_5392,N_2918,N_3624);
nand U5393 (N_5393,N_3713,N_2154);
nor U5394 (N_5394,N_3439,N_3928);
nand U5395 (N_5395,N_2425,N_3664);
and U5396 (N_5396,N_2801,N_2193);
and U5397 (N_5397,N_3828,N_3961);
nand U5398 (N_5398,N_3569,N_2334);
xor U5399 (N_5399,N_2107,N_3232);
or U5400 (N_5400,N_3747,N_3123);
and U5401 (N_5401,N_2026,N_3725);
xnor U5402 (N_5402,N_3541,N_2997);
xnor U5403 (N_5403,N_3222,N_3897);
xor U5404 (N_5404,N_2741,N_3077);
nand U5405 (N_5405,N_3308,N_3973);
xor U5406 (N_5406,N_2020,N_3730);
nand U5407 (N_5407,N_3923,N_2305);
and U5408 (N_5408,N_2653,N_3269);
nor U5409 (N_5409,N_3233,N_3228);
nor U5410 (N_5410,N_3169,N_2550);
nor U5411 (N_5411,N_3230,N_3283);
and U5412 (N_5412,N_2834,N_3111);
nand U5413 (N_5413,N_3034,N_3524);
nor U5414 (N_5414,N_2534,N_3011);
nand U5415 (N_5415,N_3074,N_2850);
nand U5416 (N_5416,N_3523,N_3779);
and U5417 (N_5417,N_3186,N_3879);
xnor U5418 (N_5418,N_3093,N_2528);
or U5419 (N_5419,N_2611,N_3209);
nand U5420 (N_5420,N_3230,N_3379);
xor U5421 (N_5421,N_3521,N_2352);
xnor U5422 (N_5422,N_2688,N_2014);
and U5423 (N_5423,N_2189,N_3510);
and U5424 (N_5424,N_3613,N_3898);
nand U5425 (N_5425,N_2768,N_2183);
and U5426 (N_5426,N_3938,N_3595);
nand U5427 (N_5427,N_2254,N_3609);
and U5428 (N_5428,N_3512,N_3195);
or U5429 (N_5429,N_3668,N_2766);
nand U5430 (N_5430,N_3046,N_2332);
and U5431 (N_5431,N_2207,N_3692);
nand U5432 (N_5432,N_2895,N_3733);
xnor U5433 (N_5433,N_2335,N_2554);
xor U5434 (N_5434,N_2540,N_2326);
nor U5435 (N_5435,N_3933,N_2234);
nand U5436 (N_5436,N_3811,N_2096);
nand U5437 (N_5437,N_3733,N_2319);
or U5438 (N_5438,N_3036,N_3959);
nor U5439 (N_5439,N_2642,N_2179);
xor U5440 (N_5440,N_2869,N_2025);
or U5441 (N_5441,N_2950,N_2824);
nand U5442 (N_5442,N_2848,N_3930);
xnor U5443 (N_5443,N_2788,N_3469);
or U5444 (N_5444,N_2602,N_3630);
nor U5445 (N_5445,N_2831,N_2590);
xnor U5446 (N_5446,N_2499,N_3167);
nand U5447 (N_5447,N_2439,N_3354);
and U5448 (N_5448,N_2684,N_3518);
xnor U5449 (N_5449,N_2047,N_2726);
xor U5450 (N_5450,N_3677,N_3696);
or U5451 (N_5451,N_2438,N_3073);
nor U5452 (N_5452,N_3497,N_2117);
nand U5453 (N_5453,N_3126,N_3990);
xnor U5454 (N_5454,N_2307,N_3381);
or U5455 (N_5455,N_3697,N_3955);
or U5456 (N_5456,N_2633,N_2180);
nor U5457 (N_5457,N_2386,N_2358);
and U5458 (N_5458,N_2847,N_3949);
xor U5459 (N_5459,N_2390,N_3997);
nand U5460 (N_5460,N_2972,N_2866);
and U5461 (N_5461,N_2119,N_2947);
nor U5462 (N_5462,N_2193,N_3284);
nand U5463 (N_5463,N_2991,N_3028);
and U5464 (N_5464,N_2709,N_3169);
and U5465 (N_5465,N_3383,N_2325);
nor U5466 (N_5466,N_3081,N_3993);
and U5467 (N_5467,N_2568,N_2590);
nor U5468 (N_5468,N_3393,N_2904);
or U5469 (N_5469,N_3636,N_2369);
or U5470 (N_5470,N_3347,N_2478);
xnor U5471 (N_5471,N_3038,N_3439);
and U5472 (N_5472,N_2679,N_2778);
nand U5473 (N_5473,N_3054,N_3863);
and U5474 (N_5474,N_2813,N_2532);
xnor U5475 (N_5475,N_2596,N_2705);
xnor U5476 (N_5476,N_2044,N_2638);
xnor U5477 (N_5477,N_2046,N_2545);
or U5478 (N_5478,N_3848,N_3790);
and U5479 (N_5479,N_3243,N_2030);
nand U5480 (N_5480,N_2615,N_3789);
nand U5481 (N_5481,N_3297,N_3370);
nor U5482 (N_5482,N_2215,N_2147);
xnor U5483 (N_5483,N_2819,N_3799);
or U5484 (N_5484,N_2346,N_3531);
and U5485 (N_5485,N_2982,N_3718);
or U5486 (N_5486,N_2150,N_3761);
or U5487 (N_5487,N_3011,N_3741);
nor U5488 (N_5488,N_3383,N_3993);
nand U5489 (N_5489,N_2789,N_3999);
nor U5490 (N_5490,N_2931,N_3201);
and U5491 (N_5491,N_2725,N_2509);
xor U5492 (N_5492,N_2495,N_3745);
nor U5493 (N_5493,N_2169,N_3233);
nand U5494 (N_5494,N_3959,N_3061);
or U5495 (N_5495,N_2161,N_3893);
xnor U5496 (N_5496,N_3248,N_3316);
xnor U5497 (N_5497,N_3899,N_2122);
or U5498 (N_5498,N_3186,N_2620);
nor U5499 (N_5499,N_3698,N_2720);
or U5500 (N_5500,N_3981,N_2720);
nor U5501 (N_5501,N_2025,N_3296);
xnor U5502 (N_5502,N_3675,N_2848);
xnor U5503 (N_5503,N_3143,N_3415);
and U5504 (N_5504,N_3785,N_3205);
nand U5505 (N_5505,N_2613,N_3213);
and U5506 (N_5506,N_3678,N_2646);
nor U5507 (N_5507,N_2730,N_3412);
or U5508 (N_5508,N_2754,N_2138);
nor U5509 (N_5509,N_2840,N_2575);
nor U5510 (N_5510,N_2677,N_3201);
xnor U5511 (N_5511,N_3666,N_2993);
or U5512 (N_5512,N_2622,N_3771);
nor U5513 (N_5513,N_2799,N_2341);
nand U5514 (N_5514,N_3651,N_2533);
xor U5515 (N_5515,N_3054,N_3799);
or U5516 (N_5516,N_3435,N_2423);
xor U5517 (N_5517,N_2530,N_3219);
nand U5518 (N_5518,N_3807,N_3313);
xnor U5519 (N_5519,N_2851,N_2360);
nor U5520 (N_5520,N_2067,N_3966);
or U5521 (N_5521,N_2670,N_2573);
nand U5522 (N_5522,N_3295,N_3298);
nand U5523 (N_5523,N_2160,N_3344);
or U5524 (N_5524,N_3606,N_3791);
nand U5525 (N_5525,N_3917,N_3286);
xor U5526 (N_5526,N_2753,N_3724);
or U5527 (N_5527,N_3180,N_3455);
or U5528 (N_5528,N_2572,N_2379);
nor U5529 (N_5529,N_3523,N_2601);
nor U5530 (N_5530,N_2239,N_2343);
and U5531 (N_5531,N_2169,N_2110);
nor U5532 (N_5532,N_2434,N_2873);
nand U5533 (N_5533,N_3253,N_3740);
nor U5534 (N_5534,N_3965,N_3531);
xnor U5535 (N_5535,N_2423,N_3396);
xnor U5536 (N_5536,N_2115,N_2739);
xnor U5537 (N_5537,N_2734,N_2537);
or U5538 (N_5538,N_3108,N_3190);
xor U5539 (N_5539,N_3613,N_3257);
xor U5540 (N_5540,N_3312,N_2803);
nor U5541 (N_5541,N_2206,N_2290);
nand U5542 (N_5542,N_2334,N_2109);
xor U5543 (N_5543,N_3577,N_3766);
and U5544 (N_5544,N_3490,N_3085);
nand U5545 (N_5545,N_3995,N_3227);
nand U5546 (N_5546,N_3488,N_2438);
xnor U5547 (N_5547,N_3434,N_3988);
nor U5548 (N_5548,N_3627,N_2653);
nor U5549 (N_5549,N_2351,N_2529);
nor U5550 (N_5550,N_3702,N_2508);
and U5551 (N_5551,N_2381,N_3393);
nor U5552 (N_5552,N_3422,N_3403);
and U5553 (N_5553,N_3795,N_3635);
nand U5554 (N_5554,N_2681,N_3714);
nand U5555 (N_5555,N_3353,N_3038);
or U5556 (N_5556,N_2262,N_3581);
nor U5557 (N_5557,N_3184,N_2321);
xnor U5558 (N_5558,N_2748,N_3009);
and U5559 (N_5559,N_3583,N_2560);
xnor U5560 (N_5560,N_2012,N_3333);
nor U5561 (N_5561,N_2839,N_3205);
and U5562 (N_5562,N_3945,N_3408);
and U5563 (N_5563,N_3816,N_3522);
xor U5564 (N_5564,N_3930,N_2500);
and U5565 (N_5565,N_2736,N_2690);
nand U5566 (N_5566,N_3086,N_2469);
nand U5567 (N_5567,N_2974,N_2037);
nand U5568 (N_5568,N_2969,N_2447);
nand U5569 (N_5569,N_3478,N_3752);
xor U5570 (N_5570,N_2731,N_3048);
xnor U5571 (N_5571,N_2154,N_3600);
nor U5572 (N_5572,N_3954,N_3441);
nor U5573 (N_5573,N_3631,N_3952);
xnor U5574 (N_5574,N_2940,N_2728);
and U5575 (N_5575,N_2411,N_3713);
nor U5576 (N_5576,N_2921,N_2219);
xor U5577 (N_5577,N_2638,N_2097);
xor U5578 (N_5578,N_3569,N_3457);
or U5579 (N_5579,N_3071,N_3548);
and U5580 (N_5580,N_3309,N_2198);
and U5581 (N_5581,N_2521,N_3643);
nor U5582 (N_5582,N_3988,N_3474);
or U5583 (N_5583,N_2681,N_2538);
nand U5584 (N_5584,N_2507,N_3517);
and U5585 (N_5585,N_3807,N_3771);
or U5586 (N_5586,N_3429,N_2334);
or U5587 (N_5587,N_3336,N_2051);
or U5588 (N_5588,N_2571,N_3638);
or U5589 (N_5589,N_2968,N_2720);
nand U5590 (N_5590,N_2681,N_3311);
xor U5591 (N_5591,N_2718,N_3534);
xor U5592 (N_5592,N_2923,N_2099);
nor U5593 (N_5593,N_2154,N_3179);
and U5594 (N_5594,N_3239,N_2688);
nor U5595 (N_5595,N_2449,N_3343);
nor U5596 (N_5596,N_2490,N_3242);
nand U5597 (N_5597,N_2515,N_2258);
nand U5598 (N_5598,N_3095,N_2632);
nor U5599 (N_5599,N_3559,N_2383);
nand U5600 (N_5600,N_2336,N_3459);
nand U5601 (N_5601,N_2440,N_3432);
and U5602 (N_5602,N_3415,N_3262);
and U5603 (N_5603,N_2894,N_2053);
xnor U5604 (N_5604,N_3726,N_2420);
xor U5605 (N_5605,N_2195,N_2411);
or U5606 (N_5606,N_3844,N_2864);
nor U5607 (N_5607,N_3770,N_3912);
xnor U5608 (N_5608,N_2899,N_3273);
or U5609 (N_5609,N_3370,N_3000);
and U5610 (N_5610,N_2445,N_3468);
and U5611 (N_5611,N_3569,N_3060);
or U5612 (N_5612,N_2625,N_3725);
nand U5613 (N_5613,N_2606,N_3288);
xor U5614 (N_5614,N_2972,N_2164);
nand U5615 (N_5615,N_3925,N_2099);
nor U5616 (N_5616,N_3739,N_2033);
xnor U5617 (N_5617,N_3447,N_2214);
nor U5618 (N_5618,N_2622,N_3095);
xnor U5619 (N_5619,N_3559,N_2355);
nor U5620 (N_5620,N_2300,N_2529);
xnor U5621 (N_5621,N_2241,N_3387);
nor U5622 (N_5622,N_3173,N_2252);
and U5623 (N_5623,N_3440,N_3197);
or U5624 (N_5624,N_2511,N_3005);
nand U5625 (N_5625,N_2153,N_3946);
and U5626 (N_5626,N_3739,N_2167);
nand U5627 (N_5627,N_3210,N_3308);
nor U5628 (N_5628,N_3883,N_2807);
and U5629 (N_5629,N_2128,N_3507);
and U5630 (N_5630,N_3529,N_3927);
xor U5631 (N_5631,N_3168,N_3267);
or U5632 (N_5632,N_2312,N_3765);
and U5633 (N_5633,N_3788,N_3616);
nand U5634 (N_5634,N_2037,N_3264);
and U5635 (N_5635,N_3491,N_2226);
nor U5636 (N_5636,N_3484,N_2707);
nor U5637 (N_5637,N_2764,N_2303);
or U5638 (N_5638,N_2626,N_3511);
or U5639 (N_5639,N_3557,N_2048);
nand U5640 (N_5640,N_2418,N_2868);
and U5641 (N_5641,N_3808,N_2084);
and U5642 (N_5642,N_3278,N_2977);
nand U5643 (N_5643,N_2296,N_2150);
nand U5644 (N_5644,N_2741,N_2349);
and U5645 (N_5645,N_2828,N_3705);
nor U5646 (N_5646,N_3102,N_2069);
and U5647 (N_5647,N_3958,N_2391);
and U5648 (N_5648,N_3115,N_3735);
nor U5649 (N_5649,N_2897,N_2102);
and U5650 (N_5650,N_3787,N_3242);
or U5651 (N_5651,N_3561,N_2404);
nand U5652 (N_5652,N_3535,N_2436);
nor U5653 (N_5653,N_2555,N_3701);
nand U5654 (N_5654,N_2852,N_3142);
nor U5655 (N_5655,N_3293,N_2817);
xor U5656 (N_5656,N_2971,N_2699);
and U5657 (N_5657,N_3300,N_2898);
nand U5658 (N_5658,N_2448,N_3373);
or U5659 (N_5659,N_2829,N_2194);
and U5660 (N_5660,N_2821,N_3832);
and U5661 (N_5661,N_3991,N_2134);
xnor U5662 (N_5662,N_2200,N_3239);
nand U5663 (N_5663,N_2111,N_3038);
or U5664 (N_5664,N_2981,N_2960);
nor U5665 (N_5665,N_2408,N_2003);
or U5666 (N_5666,N_3063,N_2872);
xnor U5667 (N_5667,N_3477,N_2411);
nand U5668 (N_5668,N_2322,N_2204);
and U5669 (N_5669,N_2334,N_3972);
and U5670 (N_5670,N_2802,N_3870);
xor U5671 (N_5671,N_2682,N_2963);
or U5672 (N_5672,N_3910,N_3005);
nand U5673 (N_5673,N_2183,N_2157);
xor U5674 (N_5674,N_3976,N_3637);
nor U5675 (N_5675,N_3071,N_3046);
nand U5676 (N_5676,N_3803,N_3600);
xnor U5677 (N_5677,N_3329,N_3290);
nand U5678 (N_5678,N_2796,N_2098);
nor U5679 (N_5679,N_2407,N_2247);
xnor U5680 (N_5680,N_2743,N_2352);
nor U5681 (N_5681,N_2610,N_3401);
and U5682 (N_5682,N_3784,N_2442);
nand U5683 (N_5683,N_3185,N_2926);
xnor U5684 (N_5684,N_2602,N_3421);
xor U5685 (N_5685,N_3833,N_2544);
or U5686 (N_5686,N_3635,N_2326);
and U5687 (N_5687,N_2539,N_2875);
and U5688 (N_5688,N_2955,N_3605);
nor U5689 (N_5689,N_2451,N_3572);
xnor U5690 (N_5690,N_2901,N_2067);
or U5691 (N_5691,N_3763,N_3173);
nor U5692 (N_5692,N_3948,N_3074);
xnor U5693 (N_5693,N_3269,N_2102);
and U5694 (N_5694,N_3443,N_2534);
nand U5695 (N_5695,N_3067,N_2273);
nor U5696 (N_5696,N_2136,N_3611);
and U5697 (N_5697,N_2440,N_2662);
nand U5698 (N_5698,N_3778,N_2753);
nand U5699 (N_5699,N_3551,N_3006);
or U5700 (N_5700,N_3373,N_3792);
nand U5701 (N_5701,N_3687,N_2577);
nor U5702 (N_5702,N_2121,N_3149);
or U5703 (N_5703,N_3212,N_3648);
and U5704 (N_5704,N_2881,N_2617);
and U5705 (N_5705,N_3094,N_3689);
nand U5706 (N_5706,N_2393,N_3715);
and U5707 (N_5707,N_3383,N_2504);
xnor U5708 (N_5708,N_3601,N_3696);
nand U5709 (N_5709,N_3271,N_2435);
nor U5710 (N_5710,N_2873,N_2069);
xnor U5711 (N_5711,N_2520,N_2144);
nor U5712 (N_5712,N_3607,N_3602);
nor U5713 (N_5713,N_2784,N_2468);
xnor U5714 (N_5714,N_2875,N_3463);
and U5715 (N_5715,N_2486,N_3377);
and U5716 (N_5716,N_2356,N_2574);
xnor U5717 (N_5717,N_3810,N_3085);
and U5718 (N_5718,N_3490,N_3390);
xnor U5719 (N_5719,N_2415,N_2417);
nor U5720 (N_5720,N_3790,N_2327);
xor U5721 (N_5721,N_2230,N_2393);
or U5722 (N_5722,N_3890,N_2792);
nor U5723 (N_5723,N_3995,N_2558);
nor U5724 (N_5724,N_3104,N_3984);
nor U5725 (N_5725,N_2442,N_2998);
nor U5726 (N_5726,N_3670,N_2649);
xnor U5727 (N_5727,N_2452,N_2814);
or U5728 (N_5728,N_3107,N_3249);
nand U5729 (N_5729,N_2237,N_2093);
or U5730 (N_5730,N_3200,N_2685);
xor U5731 (N_5731,N_3215,N_2566);
or U5732 (N_5732,N_2680,N_2963);
xor U5733 (N_5733,N_2330,N_2984);
and U5734 (N_5734,N_2470,N_2035);
nor U5735 (N_5735,N_3008,N_3312);
nand U5736 (N_5736,N_3297,N_2970);
and U5737 (N_5737,N_3955,N_3713);
or U5738 (N_5738,N_2406,N_2192);
nor U5739 (N_5739,N_3284,N_3768);
or U5740 (N_5740,N_2171,N_2793);
xor U5741 (N_5741,N_2732,N_2756);
or U5742 (N_5742,N_3386,N_2817);
nor U5743 (N_5743,N_3318,N_2908);
nor U5744 (N_5744,N_3430,N_2464);
xor U5745 (N_5745,N_3758,N_3676);
nor U5746 (N_5746,N_3265,N_3580);
and U5747 (N_5747,N_2153,N_2207);
or U5748 (N_5748,N_2741,N_3854);
nand U5749 (N_5749,N_3766,N_3737);
xnor U5750 (N_5750,N_2698,N_2650);
xnor U5751 (N_5751,N_2456,N_2727);
and U5752 (N_5752,N_2534,N_3136);
nor U5753 (N_5753,N_3038,N_3952);
nor U5754 (N_5754,N_2589,N_2406);
nand U5755 (N_5755,N_3523,N_3164);
or U5756 (N_5756,N_3567,N_2267);
and U5757 (N_5757,N_3288,N_3843);
or U5758 (N_5758,N_2437,N_3360);
and U5759 (N_5759,N_3231,N_3015);
nand U5760 (N_5760,N_2366,N_2408);
nor U5761 (N_5761,N_3056,N_2161);
and U5762 (N_5762,N_3850,N_3531);
nor U5763 (N_5763,N_2395,N_3866);
and U5764 (N_5764,N_3003,N_3111);
nand U5765 (N_5765,N_3104,N_2404);
nand U5766 (N_5766,N_2163,N_3873);
and U5767 (N_5767,N_3863,N_2302);
nor U5768 (N_5768,N_3563,N_3989);
xnor U5769 (N_5769,N_3986,N_2568);
nand U5770 (N_5770,N_2451,N_2850);
and U5771 (N_5771,N_2797,N_2279);
and U5772 (N_5772,N_2788,N_2462);
or U5773 (N_5773,N_3362,N_2587);
and U5774 (N_5774,N_3245,N_3981);
and U5775 (N_5775,N_3132,N_2145);
and U5776 (N_5776,N_2713,N_3759);
xnor U5777 (N_5777,N_3217,N_3960);
xor U5778 (N_5778,N_3104,N_2246);
nor U5779 (N_5779,N_3822,N_2101);
xor U5780 (N_5780,N_3574,N_3857);
nor U5781 (N_5781,N_3116,N_3557);
and U5782 (N_5782,N_3986,N_3939);
and U5783 (N_5783,N_3057,N_3665);
nor U5784 (N_5784,N_3859,N_3526);
and U5785 (N_5785,N_3327,N_2446);
nand U5786 (N_5786,N_2078,N_2270);
and U5787 (N_5787,N_2736,N_3271);
nor U5788 (N_5788,N_3804,N_3922);
xor U5789 (N_5789,N_2453,N_3629);
nand U5790 (N_5790,N_2645,N_2241);
nor U5791 (N_5791,N_2710,N_2420);
xnor U5792 (N_5792,N_2473,N_2937);
and U5793 (N_5793,N_3366,N_2988);
nand U5794 (N_5794,N_3902,N_2344);
or U5795 (N_5795,N_2606,N_3135);
nor U5796 (N_5796,N_3007,N_2503);
and U5797 (N_5797,N_2683,N_2981);
nand U5798 (N_5798,N_3151,N_2335);
and U5799 (N_5799,N_2300,N_3549);
or U5800 (N_5800,N_3815,N_3654);
nor U5801 (N_5801,N_2009,N_3615);
xor U5802 (N_5802,N_2847,N_2969);
nor U5803 (N_5803,N_2147,N_2622);
nor U5804 (N_5804,N_2199,N_2858);
and U5805 (N_5805,N_3092,N_2533);
and U5806 (N_5806,N_3001,N_3942);
xor U5807 (N_5807,N_2801,N_2007);
or U5808 (N_5808,N_2889,N_3711);
and U5809 (N_5809,N_3768,N_2452);
nand U5810 (N_5810,N_3861,N_2147);
nand U5811 (N_5811,N_3028,N_2306);
xor U5812 (N_5812,N_3435,N_3882);
nor U5813 (N_5813,N_3123,N_3130);
or U5814 (N_5814,N_3413,N_3052);
xnor U5815 (N_5815,N_2016,N_2715);
and U5816 (N_5816,N_3723,N_3664);
nor U5817 (N_5817,N_3993,N_2195);
xnor U5818 (N_5818,N_2798,N_2132);
nor U5819 (N_5819,N_3301,N_2386);
or U5820 (N_5820,N_3263,N_2380);
xor U5821 (N_5821,N_2499,N_3812);
nand U5822 (N_5822,N_3912,N_3458);
or U5823 (N_5823,N_2783,N_3363);
nor U5824 (N_5824,N_3263,N_3594);
xor U5825 (N_5825,N_3082,N_3462);
nor U5826 (N_5826,N_3883,N_3065);
and U5827 (N_5827,N_3624,N_3245);
or U5828 (N_5828,N_2500,N_3430);
or U5829 (N_5829,N_2664,N_2473);
or U5830 (N_5830,N_2998,N_2392);
and U5831 (N_5831,N_3885,N_2163);
or U5832 (N_5832,N_3474,N_3327);
nand U5833 (N_5833,N_3878,N_3706);
nor U5834 (N_5834,N_2919,N_3290);
xnor U5835 (N_5835,N_2612,N_3967);
xor U5836 (N_5836,N_3023,N_3770);
and U5837 (N_5837,N_3279,N_2129);
nor U5838 (N_5838,N_3411,N_3326);
or U5839 (N_5839,N_3552,N_3612);
or U5840 (N_5840,N_2750,N_3719);
or U5841 (N_5841,N_3038,N_2444);
and U5842 (N_5842,N_2968,N_3970);
xnor U5843 (N_5843,N_2712,N_3392);
nand U5844 (N_5844,N_3433,N_2410);
nand U5845 (N_5845,N_3650,N_3628);
and U5846 (N_5846,N_3914,N_2793);
nor U5847 (N_5847,N_3110,N_2245);
nand U5848 (N_5848,N_2585,N_3496);
nor U5849 (N_5849,N_3606,N_3141);
and U5850 (N_5850,N_3726,N_2222);
and U5851 (N_5851,N_2086,N_3903);
xor U5852 (N_5852,N_3169,N_2765);
and U5853 (N_5853,N_2122,N_3259);
nor U5854 (N_5854,N_3385,N_3969);
or U5855 (N_5855,N_2132,N_3708);
nand U5856 (N_5856,N_3663,N_2478);
nand U5857 (N_5857,N_2401,N_2192);
xnor U5858 (N_5858,N_2594,N_3557);
nor U5859 (N_5859,N_2265,N_3151);
xor U5860 (N_5860,N_2156,N_2376);
xor U5861 (N_5861,N_2802,N_2704);
nand U5862 (N_5862,N_3929,N_3046);
nor U5863 (N_5863,N_2722,N_2480);
xor U5864 (N_5864,N_3886,N_3815);
or U5865 (N_5865,N_3926,N_2239);
nor U5866 (N_5866,N_3770,N_2964);
or U5867 (N_5867,N_3000,N_2702);
xor U5868 (N_5868,N_3766,N_3389);
and U5869 (N_5869,N_2656,N_3300);
or U5870 (N_5870,N_3300,N_3900);
xor U5871 (N_5871,N_3224,N_2715);
or U5872 (N_5872,N_2826,N_3026);
and U5873 (N_5873,N_3504,N_3835);
xor U5874 (N_5874,N_3437,N_3970);
xnor U5875 (N_5875,N_3008,N_3152);
and U5876 (N_5876,N_2076,N_2272);
nor U5877 (N_5877,N_2849,N_2111);
xnor U5878 (N_5878,N_3459,N_2679);
xnor U5879 (N_5879,N_3155,N_2158);
nand U5880 (N_5880,N_3921,N_2015);
xor U5881 (N_5881,N_3159,N_3259);
and U5882 (N_5882,N_2748,N_3062);
or U5883 (N_5883,N_3903,N_2741);
or U5884 (N_5884,N_2334,N_2031);
or U5885 (N_5885,N_3069,N_3170);
nor U5886 (N_5886,N_3333,N_3979);
and U5887 (N_5887,N_3267,N_2782);
nor U5888 (N_5888,N_2241,N_3400);
and U5889 (N_5889,N_3266,N_3917);
xor U5890 (N_5890,N_2404,N_3099);
or U5891 (N_5891,N_3362,N_3588);
xnor U5892 (N_5892,N_2261,N_3666);
nor U5893 (N_5893,N_3838,N_2764);
nor U5894 (N_5894,N_2501,N_3831);
nand U5895 (N_5895,N_2580,N_2373);
or U5896 (N_5896,N_3286,N_3536);
and U5897 (N_5897,N_2755,N_3333);
and U5898 (N_5898,N_3485,N_3157);
xnor U5899 (N_5899,N_2689,N_2772);
nand U5900 (N_5900,N_2748,N_2045);
nand U5901 (N_5901,N_3005,N_2590);
xor U5902 (N_5902,N_3990,N_3574);
or U5903 (N_5903,N_3077,N_2551);
nand U5904 (N_5904,N_2674,N_3083);
nor U5905 (N_5905,N_3850,N_2125);
or U5906 (N_5906,N_3173,N_2362);
nand U5907 (N_5907,N_3009,N_3587);
nor U5908 (N_5908,N_2654,N_2976);
or U5909 (N_5909,N_3485,N_3098);
or U5910 (N_5910,N_3115,N_2867);
nor U5911 (N_5911,N_3951,N_3712);
and U5912 (N_5912,N_3158,N_2442);
nand U5913 (N_5913,N_2763,N_3328);
nor U5914 (N_5914,N_3506,N_3729);
nor U5915 (N_5915,N_3576,N_3488);
or U5916 (N_5916,N_3293,N_2074);
xor U5917 (N_5917,N_2586,N_2921);
nand U5918 (N_5918,N_3414,N_3144);
or U5919 (N_5919,N_3539,N_3444);
xnor U5920 (N_5920,N_2064,N_3868);
nand U5921 (N_5921,N_2014,N_3977);
or U5922 (N_5922,N_3909,N_2286);
xor U5923 (N_5923,N_3050,N_2126);
xor U5924 (N_5924,N_3655,N_3269);
and U5925 (N_5925,N_2860,N_3194);
and U5926 (N_5926,N_3295,N_2437);
and U5927 (N_5927,N_2519,N_3892);
or U5928 (N_5928,N_3834,N_3606);
nand U5929 (N_5929,N_3624,N_3115);
and U5930 (N_5930,N_2479,N_2601);
and U5931 (N_5931,N_2353,N_3299);
or U5932 (N_5932,N_2447,N_2720);
nand U5933 (N_5933,N_3383,N_2817);
nand U5934 (N_5934,N_2936,N_2177);
or U5935 (N_5935,N_2720,N_3467);
and U5936 (N_5936,N_3086,N_3284);
and U5937 (N_5937,N_2920,N_3127);
xor U5938 (N_5938,N_2522,N_2985);
and U5939 (N_5939,N_2350,N_3841);
or U5940 (N_5940,N_2839,N_2175);
or U5941 (N_5941,N_2496,N_2935);
xnor U5942 (N_5942,N_2108,N_3635);
or U5943 (N_5943,N_3710,N_2529);
nor U5944 (N_5944,N_2110,N_3022);
and U5945 (N_5945,N_3544,N_2826);
or U5946 (N_5946,N_3970,N_2650);
nor U5947 (N_5947,N_2941,N_2786);
xor U5948 (N_5948,N_3359,N_3430);
nand U5949 (N_5949,N_2271,N_2354);
xor U5950 (N_5950,N_3852,N_3735);
xor U5951 (N_5951,N_2360,N_2372);
or U5952 (N_5952,N_3810,N_2729);
xor U5953 (N_5953,N_2916,N_2223);
nor U5954 (N_5954,N_3721,N_2499);
or U5955 (N_5955,N_2210,N_3134);
nor U5956 (N_5956,N_3650,N_2192);
nor U5957 (N_5957,N_2535,N_2465);
nor U5958 (N_5958,N_2443,N_2305);
and U5959 (N_5959,N_3371,N_2202);
nand U5960 (N_5960,N_3202,N_3684);
xor U5961 (N_5961,N_3717,N_3816);
and U5962 (N_5962,N_2600,N_3807);
and U5963 (N_5963,N_3740,N_3743);
and U5964 (N_5964,N_2334,N_2146);
nand U5965 (N_5965,N_2778,N_3076);
nand U5966 (N_5966,N_2388,N_3738);
nand U5967 (N_5967,N_2141,N_3747);
or U5968 (N_5968,N_3599,N_3992);
nand U5969 (N_5969,N_3738,N_3980);
nand U5970 (N_5970,N_2435,N_2425);
or U5971 (N_5971,N_3180,N_2084);
and U5972 (N_5972,N_3091,N_2026);
nor U5973 (N_5973,N_2499,N_2178);
and U5974 (N_5974,N_2387,N_3095);
nor U5975 (N_5975,N_2988,N_3671);
nand U5976 (N_5976,N_2282,N_2061);
nor U5977 (N_5977,N_3321,N_2049);
nand U5978 (N_5978,N_2108,N_2834);
nand U5979 (N_5979,N_2518,N_2303);
and U5980 (N_5980,N_2973,N_2635);
xnor U5981 (N_5981,N_2528,N_2786);
nor U5982 (N_5982,N_2845,N_2462);
nor U5983 (N_5983,N_3740,N_2318);
or U5984 (N_5984,N_3319,N_2111);
nor U5985 (N_5985,N_3049,N_3138);
xor U5986 (N_5986,N_2124,N_3407);
nor U5987 (N_5987,N_3578,N_3698);
and U5988 (N_5988,N_2065,N_3444);
nand U5989 (N_5989,N_3084,N_3034);
nand U5990 (N_5990,N_2811,N_2399);
xnor U5991 (N_5991,N_3941,N_2524);
xor U5992 (N_5992,N_3699,N_3455);
xnor U5993 (N_5993,N_3723,N_3569);
xor U5994 (N_5994,N_3416,N_2395);
nor U5995 (N_5995,N_2045,N_3151);
xor U5996 (N_5996,N_3257,N_2896);
nor U5997 (N_5997,N_3000,N_2100);
or U5998 (N_5998,N_2530,N_2111);
nor U5999 (N_5999,N_2732,N_3629);
nand U6000 (N_6000,N_5042,N_5383);
and U6001 (N_6001,N_5266,N_4573);
and U6002 (N_6002,N_4759,N_5679);
and U6003 (N_6003,N_5457,N_4056);
nand U6004 (N_6004,N_4121,N_4371);
and U6005 (N_6005,N_5808,N_5045);
or U6006 (N_6006,N_4649,N_5711);
nand U6007 (N_6007,N_4102,N_4194);
and U6008 (N_6008,N_4541,N_5104);
nor U6009 (N_6009,N_5773,N_5409);
nor U6010 (N_6010,N_5989,N_4819);
xnor U6011 (N_6011,N_4171,N_5064);
xnor U6012 (N_6012,N_4313,N_5872);
or U6013 (N_6013,N_5322,N_4531);
nor U6014 (N_6014,N_5502,N_5215);
or U6015 (N_6015,N_4600,N_4461);
nand U6016 (N_6016,N_5429,N_5174);
xnor U6017 (N_6017,N_4682,N_5867);
nand U6018 (N_6018,N_4504,N_5547);
nor U6019 (N_6019,N_5360,N_4611);
xnor U6020 (N_6020,N_5603,N_5198);
nor U6021 (N_6021,N_4091,N_4775);
and U6022 (N_6022,N_5372,N_5850);
and U6023 (N_6023,N_4314,N_5203);
nor U6024 (N_6024,N_5995,N_4637);
xor U6025 (N_6025,N_5614,N_5173);
nor U6026 (N_6026,N_4807,N_4206);
xor U6027 (N_6027,N_4319,N_5578);
or U6028 (N_6028,N_5983,N_5088);
nand U6029 (N_6029,N_4908,N_4557);
nor U6030 (N_6030,N_4550,N_5021);
xnor U6031 (N_6031,N_5297,N_4279);
nor U6032 (N_6032,N_4652,N_5269);
nand U6033 (N_6033,N_4059,N_5506);
and U6034 (N_6034,N_5859,N_4125);
nor U6035 (N_6035,N_4561,N_4006);
and U6036 (N_6036,N_5272,N_5075);
nor U6037 (N_6037,N_5294,N_5468);
or U6038 (N_6038,N_4638,N_5252);
nor U6039 (N_6039,N_4182,N_4164);
or U6040 (N_6040,N_4812,N_5304);
nand U6041 (N_6041,N_4712,N_4583);
and U6042 (N_6042,N_5564,N_4814);
and U6043 (N_6043,N_4594,N_4835);
or U6044 (N_6044,N_4894,N_4018);
xor U6045 (N_6045,N_4867,N_4554);
and U6046 (N_6046,N_5384,N_4996);
xor U6047 (N_6047,N_4847,N_4792);
xnor U6048 (N_6048,N_5340,N_5149);
nor U6049 (N_6049,N_5566,N_4346);
nand U6050 (N_6050,N_5754,N_5542);
or U6051 (N_6051,N_4196,N_5151);
nand U6052 (N_6052,N_4132,N_4238);
or U6053 (N_6053,N_4403,N_4258);
nand U6054 (N_6054,N_4640,N_5108);
and U6055 (N_6055,N_4767,N_5038);
nor U6056 (N_6056,N_5598,N_5565);
nor U6057 (N_6057,N_4119,N_4278);
xnor U6058 (N_6058,N_5971,N_5703);
or U6059 (N_6059,N_5790,N_4489);
nor U6060 (N_6060,N_4694,N_5433);
xor U6061 (N_6061,N_4919,N_4200);
xor U6062 (N_6062,N_5617,N_4046);
and U6063 (N_6063,N_4273,N_5782);
xnor U6064 (N_6064,N_5054,N_5114);
and U6065 (N_6065,N_4395,N_4872);
and U6066 (N_6066,N_5411,N_5885);
xnor U6067 (N_6067,N_4645,N_4928);
or U6068 (N_6068,N_4739,N_5972);
and U6069 (N_6069,N_5658,N_5262);
or U6070 (N_6070,N_4513,N_4257);
xnor U6071 (N_6071,N_5017,N_5874);
nor U6072 (N_6072,N_5159,N_5955);
or U6073 (N_6073,N_5014,N_5800);
and U6074 (N_6074,N_5192,N_4113);
nand U6075 (N_6075,N_4197,N_4893);
and U6076 (N_6076,N_5690,N_5018);
nor U6077 (N_6077,N_5477,N_5356);
and U6078 (N_6078,N_4223,N_5655);
xnor U6079 (N_6079,N_4551,N_5928);
nand U6080 (N_6080,N_4868,N_5734);
nand U6081 (N_6081,N_4260,N_5556);
nand U6082 (N_6082,N_4444,N_5838);
nand U6083 (N_6083,N_5568,N_4415);
xnor U6084 (N_6084,N_5713,N_5211);
or U6085 (N_6085,N_4624,N_4949);
or U6086 (N_6086,N_5720,N_4857);
nand U6087 (N_6087,N_5438,N_4881);
nand U6088 (N_6088,N_4103,N_4219);
or U6089 (N_6089,N_4410,N_4912);
or U6090 (N_6090,N_4741,N_5237);
xor U6091 (N_6091,N_4272,N_4115);
or U6092 (N_6092,N_5353,N_5856);
and U6093 (N_6093,N_4824,N_5688);
or U6094 (N_6094,N_4790,N_5462);
nand U6095 (N_6095,N_5915,N_5794);
and U6096 (N_6096,N_4470,N_4136);
nand U6097 (N_6097,N_5534,N_5315);
and U6098 (N_6098,N_5579,N_5293);
and U6099 (N_6099,N_5555,N_5373);
and U6100 (N_6100,N_5426,N_5403);
nand U6101 (N_6101,N_4352,N_4799);
xor U6102 (N_6102,N_5076,N_5635);
and U6103 (N_6103,N_5424,N_5685);
nor U6104 (N_6104,N_4560,N_5148);
nor U6105 (N_6105,N_4475,N_5560);
or U6106 (N_6106,N_4337,N_5508);
and U6107 (N_6107,N_5553,N_4175);
and U6108 (N_6108,N_5952,N_5707);
xnor U6109 (N_6109,N_5168,N_4163);
and U6110 (N_6110,N_5227,N_4034);
xor U6111 (N_6111,N_4750,N_5739);
or U6112 (N_6112,N_5153,N_5611);
xor U6113 (N_6113,N_5706,N_5585);
nand U6114 (N_6114,N_4340,N_5851);
xnor U6115 (N_6115,N_5359,N_5319);
and U6116 (N_6116,N_4331,N_4099);
and U6117 (N_6117,N_4031,N_4098);
nor U6118 (N_6118,N_4510,N_5646);
nand U6119 (N_6119,N_5309,N_4703);
nor U6120 (N_6120,N_4935,N_5427);
xor U6121 (N_6121,N_5764,N_5879);
xor U6122 (N_6122,N_4945,N_5898);
xor U6123 (N_6123,N_4083,N_4515);
xor U6124 (N_6124,N_4774,N_4368);
nor U6125 (N_6125,N_4071,N_5759);
xor U6126 (N_6126,N_4044,N_4746);
xor U6127 (N_6127,N_4347,N_5220);
and U6128 (N_6128,N_4616,N_5852);
and U6129 (N_6129,N_4834,N_4570);
or U6130 (N_6130,N_5871,N_4931);
nand U6131 (N_6131,N_5965,N_4051);
or U6132 (N_6132,N_5669,N_5784);
xor U6133 (N_6133,N_5170,N_4229);
and U6134 (N_6134,N_4282,N_4907);
and U6135 (N_6135,N_5999,N_5847);
nand U6136 (N_6136,N_4202,N_5277);
and U6137 (N_6137,N_5721,N_4357);
and U6138 (N_6138,N_5523,N_5901);
or U6139 (N_6139,N_4829,N_4449);
nand U6140 (N_6140,N_4360,N_4298);
nor U6141 (N_6141,N_4998,N_4985);
nor U6142 (N_6142,N_5959,N_5033);
nor U6143 (N_6143,N_5126,N_5815);
nor U6144 (N_6144,N_5280,N_5714);
nor U6145 (N_6145,N_5208,N_4597);
and U6146 (N_6146,N_5939,N_5922);
or U6147 (N_6147,N_4938,N_5730);
nand U6148 (N_6148,N_5748,N_5893);
nor U6149 (N_6149,N_4388,N_5752);
nor U6150 (N_6150,N_5056,N_5327);
xnor U6151 (N_6151,N_5248,N_5591);
or U6152 (N_6152,N_5011,N_5960);
or U6153 (N_6153,N_4086,N_5738);
or U6154 (N_6154,N_4978,N_4979);
and U6155 (N_6155,N_5695,N_5588);
nor U6156 (N_6156,N_4190,N_4075);
or U6157 (N_6157,N_5582,N_4370);
or U6158 (N_6158,N_4224,N_5044);
nor U6159 (N_6159,N_4663,N_4458);
nor U6160 (N_6160,N_5886,N_4361);
nor U6161 (N_6161,N_5094,N_5116);
xor U6162 (N_6162,N_5620,N_4954);
nand U6163 (N_6163,N_5615,N_4653);
xnor U6164 (N_6164,N_4249,N_5821);
nor U6165 (N_6165,N_5767,N_5681);
and U6166 (N_6166,N_4827,N_4971);
nor U6167 (N_6167,N_5795,N_4195);
or U6168 (N_6168,N_4303,N_5736);
or U6169 (N_6169,N_4207,N_5806);
nor U6170 (N_6170,N_4657,N_4902);
nand U6171 (N_6171,N_5843,N_5586);
or U6172 (N_6172,N_4130,N_5762);
nor U6173 (N_6173,N_4491,N_4270);
nand U6174 (N_6174,N_4329,N_4925);
nand U6175 (N_6175,N_5222,N_4536);
or U6176 (N_6176,N_5414,N_4577);
or U6177 (N_6177,N_4112,N_4991);
nor U6178 (N_6178,N_4431,N_4015);
nor U6179 (N_6179,N_5077,N_5670);
or U6180 (N_6180,N_4129,N_4213);
and U6181 (N_6181,N_4064,N_4830);
and U6182 (N_6182,N_5910,N_5692);
xnor U6183 (N_6183,N_4888,N_4910);
nand U6184 (N_6184,N_5569,N_4023);
nor U6185 (N_6185,N_5050,N_5974);
nand U6186 (N_6186,N_5334,N_5543);
and U6187 (N_6187,N_4517,N_4968);
nand U6188 (N_6188,N_5811,N_4050);
or U6189 (N_6189,N_5010,N_5188);
nor U6190 (N_6190,N_4588,N_4225);
or U6191 (N_6191,N_5863,N_5613);
nor U6192 (N_6192,N_5507,N_5870);
nor U6193 (N_6193,N_5497,N_5877);
nand U6194 (N_6194,N_4743,N_4854);
nand U6195 (N_6195,N_5740,N_4151);
nor U6196 (N_6196,N_4719,N_5083);
or U6197 (N_6197,N_5717,N_5944);
and U6198 (N_6198,N_5328,N_5678);
xor U6199 (N_6199,N_4684,N_5123);
or U6200 (N_6200,N_4062,N_5365);
xor U6201 (N_6201,N_5557,N_4176);
nor U6202 (N_6202,N_4078,N_4698);
nor U6203 (N_6203,N_4832,N_5650);
nor U6204 (N_6204,N_4842,N_5936);
xnor U6205 (N_6205,N_5996,N_4443);
xor U6206 (N_6206,N_4535,N_5458);
nand U6207 (N_6207,N_5501,N_4929);
nand U6208 (N_6208,N_4027,N_4951);
nor U6209 (N_6209,N_4798,N_4492);
xor U6210 (N_6210,N_4514,N_4339);
nand U6211 (N_6211,N_4181,N_4628);
or U6212 (N_6212,N_4709,N_4858);
nand U6213 (N_6213,N_4956,N_5826);
or U6214 (N_6214,N_5078,N_4484);
and U6215 (N_6215,N_4528,N_4265);
nor U6216 (N_6216,N_4215,N_4763);
nor U6217 (N_6217,N_4362,N_5481);
xor U6218 (N_6218,N_4483,N_4785);
nor U6219 (N_6219,N_4678,N_5391);
xor U6220 (N_6220,N_4077,N_4903);
nor U6221 (N_6221,N_4363,N_4969);
nor U6222 (N_6222,N_5254,N_5621);
and U6223 (N_6223,N_4669,N_4480);
and U6224 (N_6224,N_5063,N_4315);
or U6225 (N_6225,N_5967,N_5172);
nand U6226 (N_6226,N_5179,N_5141);
nor U6227 (N_6227,N_4578,N_5402);
or U6228 (N_6228,N_4000,N_4731);
and U6229 (N_6229,N_5407,N_4451);
nand U6230 (N_6230,N_5758,N_5776);
and U6231 (N_6231,N_4727,N_4636);
nor U6232 (N_6232,N_5715,N_4376);
xor U6233 (N_6233,N_5610,N_4297);
and U6234 (N_6234,N_5594,N_4639);
or U6235 (N_6235,N_4665,N_5558);
and U6236 (N_6236,N_4381,N_5487);
or U6237 (N_6237,N_4417,N_4596);
or U6238 (N_6238,N_4017,N_5397);
nand U6239 (N_6239,N_5250,N_5401);
and U6240 (N_6240,N_5068,N_5238);
nand U6241 (N_6241,N_4328,N_4335);
or U6242 (N_6242,N_4808,N_4498);
or U6243 (N_6243,N_4664,N_5865);
xnor U6244 (N_6244,N_5793,N_5000);
nand U6245 (N_6245,N_5651,N_4274);
and U6246 (N_6246,N_5786,N_4038);
and U6247 (N_6247,N_4210,N_5226);
and U6248 (N_6248,N_4345,N_5789);
and U6249 (N_6249,N_5367,N_4780);
nand U6250 (N_6250,N_5639,N_4602);
and U6251 (N_6251,N_4654,N_4679);
nor U6252 (N_6252,N_4506,N_4478);
xnor U6253 (N_6253,N_5043,N_5381);
nor U6254 (N_6254,N_5288,N_5259);
xnor U6255 (N_6255,N_5829,N_5702);
or U6256 (N_6256,N_4526,N_4745);
nor U6257 (N_6257,N_4672,N_4326);
and U6258 (N_6258,N_5066,N_5496);
and U6259 (N_6259,N_4146,N_5812);
or U6260 (N_6260,N_5694,N_4592);
nand U6261 (N_6261,N_5583,N_4082);
nand U6262 (N_6262,N_4012,N_4898);
nor U6263 (N_6263,N_4227,N_5317);
nand U6264 (N_6264,N_5988,N_4527);
xnor U6265 (N_6265,N_4024,N_4632);
and U6266 (N_6266,N_5465,N_5004);
xnor U6267 (N_6267,N_4145,N_4423);
xnor U6268 (N_6268,N_5742,N_5062);
xor U6269 (N_6269,N_4646,N_5991);
xnor U6270 (N_6270,N_5029,N_5316);
and U6271 (N_6271,N_4294,N_5780);
nand U6272 (N_6272,N_5976,N_5489);
xnor U6273 (N_6273,N_5131,N_4601);
and U6274 (N_6274,N_5979,N_4633);
nand U6275 (N_6275,N_4953,N_5331);
nand U6276 (N_6276,N_4503,N_4656);
xnor U6277 (N_6277,N_5798,N_4674);
nand U6278 (N_6278,N_4373,N_5107);
nand U6279 (N_6279,N_4725,N_5453);
nor U6280 (N_6280,N_5535,N_5275);
nand U6281 (N_6281,N_5303,N_5561);
xor U6282 (N_6282,N_5846,N_5015);
and U6283 (N_6283,N_5765,N_5526);
nand U6284 (N_6284,N_4932,N_5949);
nand U6285 (N_6285,N_5485,N_5102);
nand U6286 (N_6286,N_4563,N_5330);
and U6287 (N_6287,N_4734,N_4730);
nand U6288 (N_6288,N_5065,N_4614);
nand U6289 (N_6289,N_5619,N_5563);
and U6290 (N_6290,N_4939,N_5325);
nor U6291 (N_6291,N_5530,N_4304);
and U6292 (N_6292,N_5858,N_5417);
nand U6293 (N_6293,N_5122,N_4149);
or U6294 (N_6294,N_4567,N_4866);
xnor U6295 (N_6295,N_4096,N_5421);
and U6296 (N_6296,N_4609,N_4160);
or U6297 (N_6297,N_5051,N_4635);
nand U6298 (N_6298,N_5190,N_4686);
or U6299 (N_6299,N_4972,N_5897);
nand U6300 (N_6300,N_5349,N_4334);
and U6301 (N_6301,N_5095,N_5419);
nor U6302 (N_6302,N_5517,N_4895);
and U6303 (N_6303,N_4961,N_5060);
and U6304 (N_6304,N_5344,N_4066);
nor U6305 (N_6305,N_5169,N_4862);
and U6306 (N_6306,N_4019,N_4037);
and U6307 (N_6307,N_5907,N_5251);
xor U6308 (N_6308,N_4469,N_4965);
or U6309 (N_6309,N_5389,N_5212);
nand U6310 (N_6310,N_4618,N_5638);
and U6311 (N_6311,N_4598,N_4205);
nand U6312 (N_6312,N_5541,N_5467);
or U6313 (N_6313,N_5006,N_4002);
nor U6314 (N_6314,N_4994,N_5495);
nand U6315 (N_6315,N_4687,N_4997);
xnor U6316 (N_6316,N_5625,N_5954);
nor U6317 (N_6317,N_4794,N_5580);
xor U6318 (N_6318,N_5282,N_5306);
and U6319 (N_6319,N_5059,N_5009);
nor U6320 (N_6320,N_5657,N_4380);
xor U6321 (N_6321,N_5341,N_4651);
and U6322 (N_6322,N_4732,N_5022);
xnor U6323 (N_6323,N_4983,N_4539);
and U6324 (N_6324,N_4786,N_5797);
or U6325 (N_6325,N_4524,N_5378);
nand U6326 (N_6326,N_5836,N_4467);
nand U6327 (N_6327,N_4555,N_5781);
and U6328 (N_6328,N_4057,N_5813);
or U6329 (N_6329,N_4354,N_4138);
xor U6330 (N_6330,N_4148,N_5571);
or U6331 (N_6331,N_4833,N_4288);
nor U6332 (N_6332,N_4990,N_5082);
and U6333 (N_6333,N_5396,N_4885);
or U6334 (N_6334,N_4843,N_5086);
nor U6335 (N_6335,N_4400,N_5333);
nor U6336 (N_6336,N_4033,N_5069);
xor U6337 (N_6337,N_5031,N_5117);
nor U6338 (N_6338,N_5181,N_4101);
xnor U6339 (N_6339,N_5070,N_5519);
xnor U6340 (N_6340,N_4424,N_4590);
nand U6341 (N_6341,N_5089,N_5351);
xnor U6342 (N_6342,N_4540,N_5618);
xor U6343 (N_6343,N_5731,N_5005);
nand U6344 (N_6344,N_4574,N_4747);
nor U6345 (N_6345,N_4011,N_5405);
or U6346 (N_6346,N_5112,N_4781);
or U6347 (N_6347,N_5674,N_5106);
or U6348 (N_6348,N_4511,N_4957);
or U6349 (N_6349,N_4166,N_4586);
nor U6350 (N_6350,N_5521,N_4496);
and U6351 (N_6351,N_5223,N_4733);
or U6352 (N_6352,N_5347,N_5778);
nor U6353 (N_6353,N_4967,N_4382);
or U6354 (N_6354,N_5125,N_5525);
nor U6355 (N_6355,N_4448,N_4520);
xnor U6356 (N_6356,N_5937,N_5242);
nand U6357 (N_6357,N_5935,N_5440);
nand U6358 (N_6358,N_4074,N_5616);
and U6359 (N_6359,N_4806,N_4825);
and U6360 (N_6360,N_4509,N_4543);
xnor U6361 (N_6361,N_5137,N_5825);
nand U6362 (N_6362,N_5743,N_5802);
nor U6363 (N_6363,N_5918,N_5777);
xnor U6364 (N_6364,N_5769,N_5354);
and U6365 (N_6365,N_4026,N_5864);
nor U6366 (N_6366,N_4292,N_4058);
xor U6367 (N_6367,N_4622,N_5358);
nor U6368 (N_6368,N_5691,N_4005);
nor U6369 (N_6369,N_5895,N_4061);
nor U6370 (N_6370,N_5435,N_4591);
nor U6371 (N_6371,N_4133,N_4783);
xor U6372 (N_6372,N_4795,N_5719);
or U6373 (N_6373,N_4142,N_5945);
nor U6374 (N_6374,N_5712,N_5861);
or U6375 (N_6375,N_4960,N_4521);
and U6376 (N_6376,N_5039,N_5528);
nand U6377 (N_6377,N_5080,N_5912);
and U6378 (N_6378,N_5196,N_4744);
xor U6379 (N_6379,N_4700,N_5992);
and U6380 (N_6380,N_5474,N_4441);
and U6381 (N_6381,N_5158,N_4135);
xnor U6382 (N_6382,N_5923,N_5040);
nand U6383 (N_6383,N_4845,N_4787);
or U6384 (N_6384,N_5200,N_4547);
and U6385 (N_6385,N_5966,N_5162);
and U6386 (N_6386,N_5410,N_5355);
and U6387 (N_6387,N_5442,N_5377);
nor U6388 (N_6388,N_5732,N_5267);
nand U6389 (N_6389,N_5150,N_5138);
and U6390 (N_6390,N_4120,N_5946);
xor U6391 (N_6391,N_5164,N_5118);
xnor U6392 (N_6392,N_4240,N_4482);
nor U6393 (N_6393,N_4261,N_4416);
or U6394 (N_6394,N_4421,N_4230);
nand U6395 (N_6395,N_5337,N_4239);
nand U6396 (N_6396,N_5264,N_4418);
xor U6397 (N_6397,N_5240,N_5504);
nand U6398 (N_6398,N_4490,N_4926);
or U6399 (N_6399,N_5810,N_5265);
nor U6400 (N_6400,N_5166,N_5536);
xnor U6401 (N_6401,N_4185,N_4826);
xnor U6402 (N_6402,N_4964,N_4715);
nor U6403 (N_6403,N_4359,N_5380);
nand U6404 (N_6404,N_4198,N_4934);
xnor U6405 (N_6405,N_4275,N_4766);
nor U6406 (N_6406,N_5513,N_4253);
or U6407 (N_6407,N_5127,N_5640);
nor U6408 (N_6408,N_4450,N_5156);
and U6409 (N_6409,N_4048,N_4587);
nor U6410 (N_6410,N_4559,N_4068);
or U6411 (N_6411,N_4505,N_5332);
or U6412 (N_6412,N_4378,N_4729);
and U6413 (N_6413,N_4407,N_5163);
nor U6414 (N_6414,N_4810,N_4765);
nand U6415 (N_6415,N_4726,N_5961);
or U6416 (N_6416,N_5592,N_4948);
and U6417 (N_6417,N_5796,N_4406);
xor U6418 (N_6418,N_5013,N_5097);
and U6419 (N_6419,N_5724,N_5318);
or U6420 (N_6420,N_5216,N_5628);
nor U6421 (N_6421,N_5735,N_4621);
xnor U6422 (N_6422,N_4377,N_5788);
or U6423 (N_6423,N_5147,N_4073);
nand U6424 (N_6424,N_4047,N_5835);
or U6425 (N_6425,N_5024,N_4626);
and U6426 (N_6426,N_5270,N_4660);
and U6427 (N_6427,N_5109,N_4105);
or U6428 (N_6428,N_5575,N_4777);
nand U6429 (N_6429,N_4152,N_4013);
nor U6430 (N_6430,N_5363,N_5387);
nand U6431 (N_6431,N_4372,N_5749);
or U6432 (N_6432,N_5883,N_4818);
nand U6433 (N_6433,N_4286,N_5866);
and U6434 (N_6434,N_5230,N_4094);
nor U6435 (N_6435,N_5607,N_5668);
nand U6436 (N_6436,N_5531,N_5087);
xnor U6437 (N_6437,N_4762,N_5143);
nand U6438 (N_6438,N_5336,N_4411);
nand U6439 (N_6439,N_5385,N_4916);
nand U6440 (N_6440,N_4816,N_4771);
nand U6441 (N_6441,N_4309,N_5343);
nor U6442 (N_6442,N_4008,N_5818);
and U6443 (N_6443,N_5152,N_4214);
or U6444 (N_6444,N_4683,N_4049);
xor U6445 (N_6445,N_4671,N_5452);
nand U6446 (N_6446,N_5180,N_5997);
and U6447 (N_6447,N_5182,N_4923);
nand U6448 (N_6448,N_4568,N_5518);
nand U6449 (N_6449,N_5020,N_5185);
or U6450 (N_6450,N_4124,N_5132);
and U6451 (N_6451,N_5984,N_4917);
and U6452 (N_6452,N_4104,N_5311);
or U6453 (N_6453,N_5134,N_5527);
or U6454 (N_6454,N_4473,N_5683);
nor U6455 (N_6455,N_4927,N_4434);
and U6456 (N_6456,N_5008,N_4126);
nor U6457 (N_6457,N_4982,N_4263);
xor U6458 (N_6458,N_4922,N_5284);
and U6459 (N_6459,N_4021,N_5823);
nor U6460 (N_6460,N_4307,N_5718);
or U6461 (N_6461,N_4837,N_5079);
xor U6462 (N_6462,N_4341,N_5231);
nor U6463 (N_6463,N_4529,N_5205);
nand U6464 (N_6464,N_4259,N_4179);
nor U6465 (N_6465,N_4374,N_4385);
or U6466 (N_6466,N_4344,N_5799);
or U6467 (N_6467,N_4070,N_4690);
nand U6468 (N_6468,N_5105,N_5194);
nor U6469 (N_6469,N_4147,N_5964);
nor U6470 (N_6470,N_4255,N_5128);
nand U6471 (N_6471,N_5932,N_5197);
and U6472 (N_6472,N_5689,N_4141);
nor U6473 (N_6473,N_4580,N_4685);
nor U6474 (N_6474,N_5570,N_5933);
xor U6475 (N_6475,N_5993,N_4457);
and U6476 (N_6476,N_5374,N_5436);
or U6477 (N_6477,N_4760,N_5839);
nand U6478 (N_6478,N_5868,N_5854);
xor U6479 (N_6479,N_4268,N_4658);
or U6480 (N_6480,N_5505,N_5225);
or U6481 (N_6481,N_4092,N_5774);
and U6482 (N_6482,N_4604,N_4793);
or U6483 (N_6483,N_4853,N_4875);
or U6484 (N_6484,N_5286,N_5023);
nand U6485 (N_6485,N_5888,N_4123);
nand U6486 (N_6486,N_5445,N_4396);
and U6487 (N_6487,N_5210,N_4134);
nor U6488 (N_6488,N_4822,N_4287);
or U6489 (N_6489,N_5837,N_5834);
nand U6490 (N_6490,N_5028,N_4264);
xnor U6491 (N_6491,N_5486,N_4946);
nand U6492 (N_6492,N_4079,N_5941);
xnor U6493 (N_6493,N_5924,N_5757);
and U6494 (N_6494,N_5310,N_4289);
nor U6495 (N_6495,N_5906,N_5455);
and U6496 (N_6496,N_5103,N_4276);
xor U6497 (N_6497,N_5982,N_5772);
xor U6498 (N_6498,N_5970,N_4324);
nor U6499 (N_6499,N_5684,N_5219);
nor U6500 (N_6500,N_5274,N_5509);
nand U6501 (N_6501,N_4659,N_4004);
and U6502 (N_6502,N_4438,N_5241);
nor U6503 (N_6503,N_4460,N_5551);
nor U6504 (N_6504,N_4488,N_4106);
or U6505 (N_6505,N_4212,N_4800);
nor U6506 (N_6506,N_4533,N_4452);
and U6507 (N_6507,N_5652,N_4617);
nor U6508 (N_6508,N_4128,N_4704);
nor U6509 (N_6509,N_5431,N_5963);
or U6510 (N_6510,N_5887,N_4291);
nor U6511 (N_6511,N_4876,N_4619);
and U6512 (N_6512,N_5538,N_4081);
nand U6513 (N_6513,N_4302,N_5642);
nor U6514 (N_6514,N_4043,N_5199);
nand U6515 (N_6515,N_4670,N_5443);
xnor U6516 (N_6516,N_5144,N_5687);
nor U6517 (N_6517,N_4349,N_4140);
and U6518 (N_6518,N_5710,N_4523);
xor U6519 (N_6519,N_5665,N_4456);
and U6520 (N_6520,N_4369,N_5191);
and U6521 (N_6521,N_5929,N_4992);
xor U6522 (N_6522,N_4797,N_4477);
and U6523 (N_6523,N_5019,N_5801);
and U6524 (N_6524,N_4446,N_5375);
or U6525 (N_6525,N_4365,N_5708);
nand U6526 (N_6526,N_5892,N_4820);
nor U6527 (N_6527,N_4241,N_5037);
nand U6528 (N_6528,N_5361,N_5581);
or U6529 (N_6529,N_5876,N_5473);
nor U6530 (N_6530,N_4072,N_4821);
nand U6531 (N_6531,N_4174,N_5048);
or U6532 (N_6532,N_4001,N_5290);
nor U6533 (N_6533,N_4764,N_4886);
xor U6534 (N_6534,N_4311,N_4327);
and U6535 (N_6535,N_5820,N_5382);
and U6536 (N_6536,N_5430,N_4187);
or U6537 (N_6537,N_5296,N_5942);
and U6538 (N_6538,N_5480,N_4462);
and U6539 (N_6539,N_4052,N_4706);
and U6540 (N_6540,N_5753,N_5756);
nand U6541 (N_6541,N_4981,N_5003);
or U6542 (N_6542,N_4076,N_4963);
nor U6543 (N_6543,N_5574,N_5605);
xnor U6544 (N_6544,N_4413,N_5699);
nor U6545 (N_6545,N_4608,N_5201);
nor U6546 (N_6546,N_4020,N_5140);
nor U6547 (N_6547,N_4728,N_4436);
or U6548 (N_6548,N_4322,N_5161);
nand U6549 (N_6549,N_5940,N_4110);
nand U6550 (N_6550,N_5400,N_5511);
nor U6551 (N_6551,N_5627,N_4010);
nor U6552 (N_6552,N_5479,N_5771);
and U6553 (N_6553,N_5247,N_5499);
nor U6554 (N_6554,N_4242,N_4525);
xor U6555 (N_6555,N_4634,N_4693);
and U6556 (N_6556,N_4883,N_5920);
nor U6557 (N_6557,N_4769,N_4947);
xor U6558 (N_6558,N_5012,N_5600);
xnor U6559 (N_6559,N_4384,N_4802);
or U6560 (N_6560,N_4299,N_4542);
nor U6561 (N_6561,N_5312,N_5157);
nor U6562 (N_6562,N_4231,N_5841);
nand U6563 (N_6563,N_4920,N_5673);
and U6564 (N_6564,N_5572,N_4468);
nand U6565 (N_6565,N_4995,N_5298);
or U6566 (N_6566,N_5943,N_4770);
nand U6567 (N_6567,N_4137,N_5217);
nand U6568 (N_6568,N_4711,N_4882);
nor U6569 (N_6569,N_5110,N_4695);
xnor U6570 (N_6570,N_5894,N_4389);
and U6571 (N_6571,N_4718,N_4673);
and U6572 (N_6572,N_5745,N_4156);
or U6573 (N_6573,N_4713,N_5700);
and U6574 (N_6574,N_4699,N_5962);
and U6575 (N_6575,N_5667,N_5408);
xnor U6576 (N_6576,N_4773,N_4203);
and U6577 (N_6577,N_4154,N_4538);
xnor U6578 (N_6578,N_4356,N_5729);
and U6579 (N_6579,N_4784,N_5493);
xnor U6580 (N_6580,N_5680,N_4863);
xor U6581 (N_6581,N_5649,N_5055);
xnor U6582 (N_6582,N_4911,N_5656);
and U6583 (N_6583,N_4173,N_4519);
xnor U6584 (N_6584,N_5121,N_4691);
nor U6585 (N_6585,N_4753,N_5633);
nand U6586 (N_6586,N_4648,N_5073);
nor U6587 (N_6587,N_4168,N_4880);
nand U6588 (N_6588,N_4724,N_4201);
xor U6589 (N_6589,N_5209,N_4918);
nand U6590 (N_6590,N_4941,N_4962);
xnor U6591 (N_6591,N_4722,N_5368);
nor U6592 (N_6592,N_5348,N_5597);
xnor U6593 (N_6593,N_4111,N_5239);
and U6594 (N_6594,N_4192,N_4401);
nor U6595 (N_6595,N_5034,N_4668);
nand U6596 (N_6596,N_5573,N_5889);
and U6597 (N_6597,N_4285,N_5931);
nor U6598 (N_6598,N_5595,N_5321);
and U6599 (N_6599,N_4317,N_4623);
nor U6600 (N_6600,N_5978,N_4476);
nor U6601 (N_6601,N_4342,N_5914);
or U6602 (N_6602,N_4850,N_5833);
and U6603 (N_6603,N_4650,N_5930);
or U6604 (N_6604,N_4364,N_4831);
or U6605 (N_6605,N_5195,N_4487);
nand U6606 (N_6606,N_5589,N_4404);
xnor U6607 (N_6607,N_4390,N_4507);
nor U6608 (N_6608,N_5300,N_4677);
nor U6609 (N_6609,N_4569,N_4943);
or U6610 (N_6610,N_4855,N_4063);
and U6611 (N_6611,N_5666,N_4815);
nand U6612 (N_6612,N_4899,N_5522);
xnor U6613 (N_6613,N_5916,N_5146);
nor U6614 (N_6614,N_4921,N_4589);
and U6615 (N_6615,N_5785,N_5926);
nand U6616 (N_6616,N_4169,N_4262);
nor U6617 (N_6617,N_4610,N_5994);
and U6618 (N_6618,N_4325,N_4655);
nand U6619 (N_6619,N_4191,N_4778);
xor U6620 (N_6620,N_4445,N_4914);
or U6621 (N_6621,N_4183,N_4705);
or U6622 (N_6622,N_4508,N_4353);
nand U6623 (N_6623,N_4290,N_5258);
nand U6624 (N_6624,N_4720,N_4321);
nand U6625 (N_6625,N_4701,N_4887);
nor U6626 (N_6626,N_4761,N_4900);
xnor U6627 (N_6627,N_4556,N_5726);
nor U6628 (N_6628,N_4114,N_4358);
and U6629 (N_6629,N_5634,N_4131);
or U6630 (N_6630,N_4028,N_4980);
xor U6631 (N_6631,N_5853,N_5295);
or U6632 (N_6632,N_5478,N_5969);
xor U6633 (N_6633,N_5213,N_5289);
and U6634 (N_6634,N_5339,N_5469);
or U6635 (N_6635,N_4466,N_5602);
nor U6636 (N_6636,N_5448,N_4150);
xnor U6637 (N_6637,N_5891,N_5559);
nand U6638 (N_6638,N_4613,N_4742);
and U6639 (N_6639,N_4877,N_5084);
nand U6640 (N_6640,N_5459,N_4065);
nor U6641 (N_6641,N_4454,N_4584);
or U6642 (N_6642,N_4859,N_4465);
and U6643 (N_6643,N_5464,N_4425);
and U6644 (N_6644,N_5263,N_5664);
xor U6645 (N_6645,N_5903,N_5099);
nand U6646 (N_6646,N_4429,N_4776);
or U6647 (N_6647,N_4428,N_4296);
nand U6648 (N_6648,N_5184,N_5204);
xnor U6649 (N_6649,N_4740,N_5661);
or U6650 (N_6650,N_5067,N_5404);
and U6651 (N_6651,N_5737,N_5819);
nor U6652 (N_6652,N_4398,N_4248);
xnor U6653 (N_6653,N_4579,N_4813);
xnor U6654 (N_6654,N_4984,N_4393);
or U6655 (N_6655,N_4714,N_4256);
nand U6656 (N_6656,N_4474,N_5256);
nand U6657 (N_6657,N_5845,N_4355);
nand U6658 (N_6658,N_5395,N_5456);
nand U6659 (N_6659,N_4986,N_4751);
and U6660 (N_6660,N_4823,N_4316);
nor U6661 (N_6661,N_4499,N_4630);
nand U6662 (N_6662,N_4045,N_5362);
or U6663 (N_6663,N_5036,N_5911);
nor U6664 (N_6664,N_4779,N_4915);
xnor U6665 (N_6665,N_5981,N_4804);
xor U6666 (N_6666,N_5193,N_5135);
and U6667 (N_6667,N_4332,N_5545);
or U6668 (N_6668,N_4772,N_5057);
nor U6669 (N_6669,N_5305,N_4305);
nand U6670 (N_6670,N_4471,N_4738);
or U6671 (N_6671,N_4933,N_4338);
nand U6672 (N_6672,N_4088,N_5115);
nand U6673 (N_6673,N_5046,N_5221);
and U6674 (N_6674,N_5938,N_4143);
nor U6675 (N_6675,N_4840,N_4427);
nor U6676 (N_6676,N_4864,N_5760);
and U6677 (N_6677,N_5139,N_4717);
or U6678 (N_6678,N_5549,N_5516);
nor U6679 (N_6679,N_5364,N_4844);
or U6680 (N_6680,N_4952,N_4204);
nand U6681 (N_6681,N_5085,N_5093);
nor U6682 (N_6682,N_4522,N_4530);
nand U6683 (N_6683,N_4716,N_5342);
nor U6684 (N_6684,N_5260,N_5584);
xor U6685 (N_6685,N_5291,N_4737);
xnor U6686 (N_6686,N_4565,N_5727);
nand U6687 (N_6687,N_5675,N_5145);
nand U6688 (N_6688,N_5779,N_4860);
and U6689 (N_6689,N_4817,N_5189);
xor U6690 (N_6690,N_5763,N_4805);
xor U6691 (N_6691,N_4437,N_4629);
or U6692 (N_6692,N_4245,N_4537);
nor U6693 (N_6693,N_5129,N_4892);
and U6694 (N_6694,N_5186,N_5491);
xor U6695 (N_6695,N_5723,N_4226);
xnor U6696 (N_6696,N_4702,N_5980);
xor U6697 (N_6697,N_4494,N_5896);
xnor U6698 (N_6698,N_5278,N_4180);
or U6699 (N_6699,N_5905,N_5552);
nor U6700 (N_6700,N_4025,N_5596);
nand U6701 (N_6701,N_4890,N_4566);
nor U6702 (N_6702,N_5326,N_4768);
nor U6703 (N_6703,N_4252,N_5329);
nor U6704 (N_6704,N_4924,N_5653);
or U6705 (N_6705,N_5268,N_4032);
and U6706 (N_6706,N_5787,N_5968);
nor U6707 (N_6707,N_4426,N_5809);
and U6708 (N_6708,N_4267,N_5142);
and U6709 (N_6709,N_5840,N_4688);
or U6710 (N_6710,N_5623,N_5725);
nor U6711 (N_6711,N_4350,N_4676);
nand U6712 (N_6712,N_4942,N_5925);
xnor U6713 (N_6713,N_4419,N_5855);
or U6714 (N_6714,N_4442,N_5313);
xnor U6715 (N_6715,N_5124,N_5816);
nor U6716 (N_6716,N_5647,N_4606);
and U6717 (N_6717,N_4246,N_5550);
nand U6718 (N_6718,N_5609,N_4796);
xor U6719 (N_6719,N_4901,N_5096);
nor U6720 (N_6720,N_5323,N_5371);
nor U6721 (N_6721,N_5601,N_4117);
xor U6722 (N_6722,N_5366,N_4386);
or U6723 (N_6723,N_5255,N_5308);
nand U6724 (N_6724,N_5958,N_4266);
nor U6725 (N_6725,N_5599,N_4975);
xor U6726 (N_6726,N_5369,N_5947);
nand U6727 (N_6727,N_4184,N_4036);
or U6728 (N_6728,N_5253,N_4803);
xor U6729 (N_6729,N_4736,N_5283);
nor U6730 (N_6730,N_5470,N_5998);
and U6731 (N_6731,N_5900,N_4402);
nor U6732 (N_6732,N_5660,N_5576);
and U6733 (N_6733,N_5704,N_4846);
nand U6734 (N_6734,N_5287,N_5654);
nand U6735 (N_6735,N_5415,N_4562);
and U6736 (N_6736,N_4089,N_4936);
xor U6737 (N_6737,N_4897,N_4891);
or U6738 (N_6738,N_5728,N_5392);
and U6739 (N_6739,N_4828,N_4170);
or U6740 (N_6740,N_5975,N_5320);
nor U6741 (N_6741,N_5081,N_5663);
or U6742 (N_6742,N_5643,N_5881);
nand U6743 (N_6743,N_4615,N_5488);
xor U6744 (N_6744,N_4913,N_4155);
nand U6745 (N_6745,N_5016,N_5091);
nand U6746 (N_6746,N_5622,N_5324);
xor U6747 (N_6747,N_4666,N_4625);
xor U6748 (N_6748,N_4999,N_4607);
xor U6749 (N_6749,N_5335,N_4937);
and U6750 (N_6750,N_5276,N_4035);
xor U6751 (N_6751,N_4055,N_5444);
nor U6752 (N_6752,N_4735,N_5463);
nand U6753 (N_6753,N_5546,N_5744);
and U6754 (N_6754,N_4647,N_4612);
nor U6755 (N_6755,N_4841,N_4383);
xor U6756 (N_6756,N_5314,N_5554);
and U6757 (N_6757,N_4409,N_4177);
nand U6758 (N_6758,N_5987,N_4486);
or U6759 (N_6759,N_5412,N_4084);
nor U6760 (N_6760,N_4399,N_4572);
nand U6761 (N_6761,N_5630,N_5842);
nor U6762 (N_6762,N_5577,N_5136);
nor U6763 (N_6763,N_4433,N_5281);
xor U6764 (N_6764,N_4493,N_4186);
and U6765 (N_6765,N_5857,N_4988);
or U6766 (N_6766,N_5904,N_4247);
nor U6767 (N_6767,N_5399,N_4878);
and U6768 (N_6768,N_4233,N_5167);
and U6769 (N_6769,N_4440,N_4394);
and U6770 (N_6770,N_4930,N_5299);
and U6771 (N_6771,N_4041,N_4464);
or U6772 (N_6772,N_4871,N_4116);
nor U6773 (N_6773,N_4755,N_4479);
and U6774 (N_6774,N_4879,N_4789);
nor U6775 (N_6775,N_5919,N_4723);
or U6776 (N_6776,N_5722,N_4014);
nand U6777 (N_6777,N_4243,N_5733);
or U6778 (N_6778,N_5460,N_5376);
nand U6779 (N_6779,N_5913,N_5672);
nor U6780 (N_6780,N_4167,N_4721);
or U6781 (N_6781,N_4696,N_5370);
nand U6782 (N_6782,N_5827,N_5053);
xor U6783 (N_6783,N_4122,N_4323);
or U6784 (N_6784,N_5814,N_4391);
and U6785 (N_6785,N_4977,N_5593);
xnor U6786 (N_6786,N_4330,N_5951);
xor U6787 (N_6787,N_4042,N_4387);
nand U6788 (N_6788,N_5232,N_5207);
nand U6789 (N_6789,N_4218,N_4809);
nand U6790 (N_6790,N_5027,N_4662);
or U6791 (N_6791,N_4300,N_5187);
nor U6792 (N_6792,N_4144,N_5768);
or U6793 (N_6793,N_4220,N_4518);
xor U6794 (N_6794,N_4667,N_4277);
or U6795 (N_6795,N_4221,N_5510);
and U6796 (N_6796,N_5171,N_5948);
or U6797 (N_6797,N_4016,N_5828);
or U6798 (N_6798,N_5899,N_4549);
or U6799 (N_6799,N_4839,N_5416);
nor U6800 (N_6800,N_5500,N_4958);
nand U6801 (N_6801,N_4710,N_5154);
or U6802 (N_6802,N_4811,N_4343);
xnor U6803 (N_6803,N_5428,N_5302);
or U6804 (N_6804,N_4605,N_4432);
xor U6805 (N_6805,N_5902,N_5608);
or U6806 (N_6806,N_4585,N_5165);
xnor U6807 (N_6807,N_5908,N_5472);
and U6808 (N_6808,N_4375,N_4007);
nor U6809 (N_6809,N_4232,N_5498);
xnor U6810 (N_6810,N_4054,N_4053);
and U6811 (N_6811,N_4085,N_5249);
or U6812 (N_6812,N_5632,N_5606);
xor U6813 (N_6813,N_5648,N_5229);
xor U6814 (N_6814,N_5567,N_4090);
nand U6815 (N_6815,N_5471,N_4269);
or U6816 (N_6816,N_5307,N_4909);
or U6817 (N_6817,N_5246,N_4748);
xnor U6818 (N_6818,N_4420,N_4595);
nand U6819 (N_6819,N_4463,N_4250);
and U6820 (N_6820,N_4564,N_5446);
or U6821 (N_6821,N_5953,N_5637);
or U6822 (N_6822,N_4552,N_5990);
nor U6823 (N_6823,N_4100,N_4139);
nand U6824 (N_6824,N_5035,N_5176);
nor U6825 (N_6825,N_5803,N_5177);
xnor U6826 (N_6826,N_5873,N_5072);
nand U6827 (N_6827,N_4158,N_5529);
nor U6828 (N_6828,N_5475,N_5461);
xnor U6829 (N_6829,N_4283,N_5693);
or U6830 (N_6830,N_5629,N_5860);
and U6831 (N_6831,N_5747,N_5869);
and U6832 (N_6832,N_5388,N_5224);
nand U6833 (N_6833,N_5515,N_5133);
nand U6834 (N_6834,N_5454,N_5659);
and U6835 (N_6835,N_5092,N_5235);
nor U6836 (N_6836,N_4162,N_5450);
or U6837 (N_6837,N_4284,N_4532);
or U6838 (N_6838,N_4333,N_4974);
nor U6839 (N_6839,N_5927,N_5766);
nor U6840 (N_6840,N_5030,N_4366);
xor U6841 (N_6841,N_4087,N_5824);
or U6842 (N_6842,N_5346,N_5466);
or U6843 (N_6843,N_4689,N_5449);
and U6844 (N_6844,N_5032,N_5245);
xor U6845 (N_6845,N_4481,N_5849);
nor U6846 (N_6846,N_4620,N_5878);
nand U6847 (N_6847,N_4500,N_5301);
xor U6848 (N_6848,N_5697,N_4849);
xnor U6849 (N_6849,N_4348,N_4109);
xor U6850 (N_6850,N_5590,N_4955);
or U6851 (N_6851,N_4642,N_5830);
xnor U6852 (N_6852,N_4312,N_4641);
nand U6853 (N_6853,N_4306,N_5671);
nand U6854 (N_6854,N_4217,N_4749);
and U6855 (N_6855,N_5160,N_4495);
or U6856 (N_6856,N_5775,N_4576);
nor U6857 (N_6857,N_4336,N_4318);
xnor U6858 (N_6858,N_4544,N_4675);
nor U6859 (N_6859,N_4692,N_5350);
xor U6860 (N_6860,N_5476,N_5832);
xor U6861 (N_6861,N_5537,N_5386);
and U6862 (N_6862,N_5183,N_5490);
nand U6863 (N_6863,N_5884,N_5909);
or U6864 (N_6864,N_5049,N_4534);
or U6865 (N_6865,N_4869,N_4447);
nand U6866 (N_6866,N_4756,N_5202);
nand U6867 (N_6867,N_4966,N_5398);
or U6868 (N_6868,N_4234,N_4707);
nor U6869 (N_6869,N_4097,N_5761);
nand U6870 (N_6870,N_4905,N_5934);
nand U6871 (N_6871,N_5271,N_5755);
and U6872 (N_6872,N_4067,N_4697);
and U6873 (N_6873,N_5236,N_5432);
xnor U6874 (N_6874,N_4801,N_5425);
or U6875 (N_6875,N_5273,N_5524);
nand U6876 (N_6876,N_5434,N_5804);
nor U6877 (N_6877,N_4422,N_4235);
nand U6878 (N_6878,N_5393,N_5484);
xnor U6879 (N_6879,N_5805,N_5413);
nor U6880 (N_6880,N_5130,N_5041);
xnor U6881 (N_6881,N_5956,N_4865);
or U6882 (N_6882,N_5279,N_4127);
or U6883 (N_6883,N_5113,N_5817);
xnor U6884 (N_6884,N_5822,N_5292);
xor U6885 (N_6885,N_4208,N_4581);
nand U6886 (N_6886,N_4178,N_4153);
or U6887 (N_6887,N_4582,N_5233);
nand U6888 (N_6888,N_4993,N_4310);
or U6889 (N_6889,N_5007,N_4367);
or U6890 (N_6890,N_5716,N_5119);
and U6891 (N_6891,N_4856,N_4884);
xnor U6892 (N_6892,N_4188,N_4603);
and U6893 (N_6893,N_5379,N_4873);
and U6894 (N_6894,N_5514,N_5644);
and U6895 (N_6895,N_4575,N_5100);
nand U6896 (N_6896,N_5026,N_5071);
nand U6897 (N_6897,N_5494,N_5645);
and U6898 (N_6898,N_4681,N_4320);
and U6899 (N_6899,N_5482,N_5701);
or U6900 (N_6900,N_4851,N_5352);
nor U6901 (N_6901,N_5844,N_5741);
nor U6902 (N_6902,N_4959,N_5807);
xor U6903 (N_6903,N_4501,N_5533);
nor U6904 (N_6904,N_4039,N_5977);
or U6905 (N_6905,N_5746,N_4412);
nor U6906 (N_6906,N_5539,N_5612);
or U6907 (N_6907,N_5390,N_5986);
and U6908 (N_6908,N_4453,N_4455);
and U6909 (N_6909,N_5052,N_4165);
nand U6910 (N_6910,N_4022,N_4029);
xnor U6911 (N_6911,N_4571,N_5423);
and U6912 (N_6912,N_5705,N_4643);
and U6913 (N_6913,N_4896,N_4472);
nor U6914 (N_6914,N_5394,N_4870);
nand U6915 (N_6915,N_4251,N_4293);
and U6916 (N_6916,N_5422,N_4599);
or U6917 (N_6917,N_4502,N_5698);
nand U6918 (N_6918,N_5770,N_5676);
nor U6919 (N_6919,N_5406,N_5338);
nand U6920 (N_6920,N_5917,N_5120);
nor U6921 (N_6921,N_4161,N_4782);
xor U6922 (N_6922,N_4280,N_4631);
nor U6923 (N_6923,N_5587,N_5001);
and U6924 (N_6924,N_5985,N_4976);
nor U6925 (N_6925,N_5604,N_4593);
nand U6926 (N_6926,N_4295,N_5257);
and U6927 (N_6927,N_4199,N_4661);
or U6928 (N_6928,N_4172,N_4644);
nor U6929 (N_6929,N_5631,N_4211);
and U6930 (N_6930,N_5512,N_4414);
nor U6931 (N_6931,N_4553,N_5111);
and U6932 (N_6932,N_4003,N_5098);
nand U6933 (N_6933,N_4545,N_5061);
or U6934 (N_6934,N_5101,N_4237);
or U6935 (N_6935,N_4405,N_4430);
and U6936 (N_6936,N_5451,N_5058);
or U6937 (N_6937,N_4209,N_4392);
xnor U6938 (N_6938,N_4351,N_5562);
nor U6939 (N_6939,N_4254,N_4236);
and U6940 (N_6940,N_5751,N_4308);
or U6941 (N_6941,N_5696,N_4788);
nand U6942 (N_6942,N_4861,N_4439);
nand U6943 (N_6943,N_5624,N_5548);
and U6944 (N_6944,N_4379,N_5791);
xor U6945 (N_6945,N_4940,N_5957);
or U6946 (N_6946,N_4497,N_5709);
nor U6947 (N_6947,N_4989,N_4485);
nor U6948 (N_6948,N_5540,N_5437);
or U6949 (N_6949,N_5441,N_5047);
or U6950 (N_6950,N_4157,N_4060);
xnor U6951 (N_6951,N_4108,N_5686);
xor U6952 (N_6952,N_5218,N_4009);
and U6953 (N_6953,N_5677,N_4093);
nor U6954 (N_6954,N_4836,N_5439);
or U6955 (N_6955,N_5544,N_4397);
and U6956 (N_6956,N_4754,N_4040);
and U6957 (N_6957,N_4558,N_4874);
xor U6958 (N_6958,N_5243,N_5002);
and U6959 (N_6959,N_5244,N_5973);
nand U6960 (N_6960,N_4271,N_5261);
xnor U6961 (N_6961,N_5074,N_5178);
nor U6962 (N_6962,N_5025,N_4030);
xor U6963 (N_6963,N_4216,N_5155);
or U6964 (N_6964,N_4516,N_5880);
nor U6965 (N_6965,N_4546,N_4889);
nor U6966 (N_6966,N_5641,N_5750);
nand U6967 (N_6967,N_4838,N_5520);
xor U6968 (N_6968,N_4757,N_5831);
nand U6969 (N_6969,N_5418,N_4228);
nand U6970 (N_6970,N_5503,N_5950);
nor U6971 (N_6971,N_4987,N_4680);
nand U6972 (N_6972,N_5447,N_5848);
nand U6973 (N_6973,N_4193,N_5175);
nor U6974 (N_6974,N_5228,N_5420);
and U6975 (N_6975,N_4944,N_4627);
nand U6976 (N_6976,N_4950,N_5345);
nand U6977 (N_6977,N_4159,N_5862);
nand U6978 (N_6978,N_4973,N_5636);
or U6979 (N_6979,N_4408,N_4080);
xor U6980 (N_6980,N_4069,N_5285);
nor U6981 (N_6981,N_4189,N_4708);
and U6982 (N_6982,N_4301,N_4758);
and U6983 (N_6983,N_5626,N_4970);
or U6984 (N_6984,N_4459,N_5682);
nand U6985 (N_6985,N_5921,N_5234);
nor U6986 (N_6986,N_4107,N_5662);
nor U6987 (N_6987,N_4904,N_4848);
xor U6988 (N_6988,N_4095,N_5532);
and U6989 (N_6989,N_4791,N_5214);
xnor U6990 (N_6990,N_5792,N_5890);
nor U6991 (N_6991,N_5492,N_4906);
and U6992 (N_6992,N_5206,N_5882);
or U6993 (N_6993,N_5783,N_4548);
and U6994 (N_6994,N_4512,N_5875);
nand U6995 (N_6995,N_4852,N_5090);
or U6996 (N_6996,N_5483,N_4281);
or U6997 (N_6997,N_4244,N_4222);
and U6998 (N_6998,N_4118,N_4752);
nand U6999 (N_6999,N_5357,N_4435);
nor U7000 (N_7000,N_4383,N_4945);
nand U7001 (N_7001,N_5676,N_5823);
or U7002 (N_7002,N_5816,N_4813);
nor U7003 (N_7003,N_5587,N_4748);
nand U7004 (N_7004,N_4767,N_4533);
or U7005 (N_7005,N_4252,N_4184);
xor U7006 (N_7006,N_4597,N_4838);
and U7007 (N_7007,N_4208,N_4314);
and U7008 (N_7008,N_4199,N_4295);
and U7009 (N_7009,N_4449,N_4431);
nand U7010 (N_7010,N_5209,N_5896);
and U7011 (N_7011,N_5192,N_4680);
or U7012 (N_7012,N_5316,N_5279);
xor U7013 (N_7013,N_4055,N_4319);
nand U7014 (N_7014,N_5129,N_4004);
and U7015 (N_7015,N_5599,N_5046);
xor U7016 (N_7016,N_4863,N_4633);
xor U7017 (N_7017,N_5545,N_5069);
xnor U7018 (N_7018,N_5725,N_5952);
or U7019 (N_7019,N_4569,N_4460);
nor U7020 (N_7020,N_4246,N_5916);
or U7021 (N_7021,N_4686,N_4791);
or U7022 (N_7022,N_4958,N_5239);
nand U7023 (N_7023,N_4743,N_4238);
nor U7024 (N_7024,N_4560,N_5453);
or U7025 (N_7025,N_5545,N_5814);
nor U7026 (N_7026,N_5454,N_5788);
xnor U7027 (N_7027,N_5560,N_5009);
or U7028 (N_7028,N_5025,N_4548);
nor U7029 (N_7029,N_5197,N_4787);
and U7030 (N_7030,N_5949,N_4771);
nor U7031 (N_7031,N_5826,N_5418);
nand U7032 (N_7032,N_4396,N_5871);
nand U7033 (N_7033,N_4747,N_5442);
nand U7034 (N_7034,N_5546,N_4359);
nand U7035 (N_7035,N_4129,N_4947);
or U7036 (N_7036,N_4165,N_5851);
nor U7037 (N_7037,N_4407,N_5981);
nor U7038 (N_7038,N_5518,N_4831);
nand U7039 (N_7039,N_5425,N_4633);
nor U7040 (N_7040,N_5421,N_4591);
or U7041 (N_7041,N_4778,N_5723);
nand U7042 (N_7042,N_5513,N_5624);
nand U7043 (N_7043,N_5892,N_5813);
or U7044 (N_7044,N_5308,N_4844);
nor U7045 (N_7045,N_4219,N_4960);
and U7046 (N_7046,N_4698,N_5432);
xnor U7047 (N_7047,N_4453,N_5138);
and U7048 (N_7048,N_5107,N_4011);
nand U7049 (N_7049,N_5816,N_4447);
nand U7050 (N_7050,N_4497,N_5685);
and U7051 (N_7051,N_5880,N_4536);
nand U7052 (N_7052,N_4412,N_4853);
and U7053 (N_7053,N_4202,N_4223);
nand U7054 (N_7054,N_5060,N_5984);
and U7055 (N_7055,N_4286,N_5017);
or U7056 (N_7056,N_4365,N_5796);
nor U7057 (N_7057,N_4523,N_4486);
nand U7058 (N_7058,N_4333,N_5224);
or U7059 (N_7059,N_4854,N_4810);
and U7060 (N_7060,N_4307,N_4750);
nor U7061 (N_7061,N_5062,N_4429);
nand U7062 (N_7062,N_5087,N_4465);
xnor U7063 (N_7063,N_4960,N_5827);
or U7064 (N_7064,N_5679,N_5639);
nor U7065 (N_7065,N_5223,N_4990);
nand U7066 (N_7066,N_4495,N_4520);
and U7067 (N_7067,N_5888,N_4959);
and U7068 (N_7068,N_4943,N_5633);
nor U7069 (N_7069,N_5287,N_5416);
nand U7070 (N_7070,N_5807,N_5572);
xor U7071 (N_7071,N_4810,N_4706);
nor U7072 (N_7072,N_5381,N_4029);
xnor U7073 (N_7073,N_5130,N_5871);
nor U7074 (N_7074,N_5095,N_4782);
or U7075 (N_7075,N_5276,N_4281);
xnor U7076 (N_7076,N_5887,N_4668);
or U7077 (N_7077,N_4302,N_4030);
nor U7078 (N_7078,N_5710,N_4275);
and U7079 (N_7079,N_4326,N_4532);
and U7080 (N_7080,N_4402,N_4120);
nand U7081 (N_7081,N_4235,N_4473);
and U7082 (N_7082,N_5589,N_4200);
xnor U7083 (N_7083,N_4191,N_4550);
nand U7084 (N_7084,N_4842,N_5627);
nor U7085 (N_7085,N_4256,N_4116);
and U7086 (N_7086,N_5620,N_5341);
xor U7087 (N_7087,N_5447,N_5783);
nor U7088 (N_7088,N_5205,N_4901);
and U7089 (N_7089,N_4847,N_5302);
xnor U7090 (N_7090,N_4105,N_5313);
and U7091 (N_7091,N_5823,N_5112);
nand U7092 (N_7092,N_4436,N_4891);
xnor U7093 (N_7093,N_4378,N_5007);
xor U7094 (N_7094,N_5323,N_4224);
nor U7095 (N_7095,N_5026,N_4202);
xnor U7096 (N_7096,N_4379,N_5167);
or U7097 (N_7097,N_4918,N_4380);
nor U7098 (N_7098,N_5536,N_5682);
nand U7099 (N_7099,N_4868,N_5705);
or U7100 (N_7100,N_5051,N_5002);
nor U7101 (N_7101,N_5480,N_5558);
nand U7102 (N_7102,N_4260,N_5790);
and U7103 (N_7103,N_5962,N_5025);
xor U7104 (N_7104,N_4085,N_5807);
nand U7105 (N_7105,N_4863,N_5239);
nand U7106 (N_7106,N_4135,N_5827);
or U7107 (N_7107,N_4907,N_4772);
nor U7108 (N_7108,N_4591,N_5698);
xor U7109 (N_7109,N_4095,N_5658);
xnor U7110 (N_7110,N_4290,N_4398);
and U7111 (N_7111,N_4510,N_5822);
or U7112 (N_7112,N_5957,N_5053);
and U7113 (N_7113,N_5172,N_4041);
and U7114 (N_7114,N_4628,N_4077);
nand U7115 (N_7115,N_5197,N_4520);
xnor U7116 (N_7116,N_5546,N_5669);
nand U7117 (N_7117,N_4246,N_4063);
and U7118 (N_7118,N_4205,N_5360);
or U7119 (N_7119,N_4000,N_4732);
or U7120 (N_7120,N_5042,N_4596);
or U7121 (N_7121,N_5637,N_5839);
or U7122 (N_7122,N_5556,N_5633);
xnor U7123 (N_7123,N_4810,N_5252);
xor U7124 (N_7124,N_4410,N_4778);
xor U7125 (N_7125,N_4046,N_4544);
and U7126 (N_7126,N_4347,N_4660);
or U7127 (N_7127,N_4695,N_4804);
and U7128 (N_7128,N_5775,N_5293);
xnor U7129 (N_7129,N_5267,N_4536);
nor U7130 (N_7130,N_4315,N_5475);
nand U7131 (N_7131,N_5387,N_5287);
nand U7132 (N_7132,N_4550,N_5090);
and U7133 (N_7133,N_4581,N_4168);
xnor U7134 (N_7134,N_5531,N_4695);
xnor U7135 (N_7135,N_4579,N_5612);
and U7136 (N_7136,N_4624,N_5173);
or U7137 (N_7137,N_4660,N_4295);
xor U7138 (N_7138,N_5620,N_5121);
or U7139 (N_7139,N_5999,N_4374);
xor U7140 (N_7140,N_5266,N_5686);
nand U7141 (N_7141,N_4591,N_4812);
nor U7142 (N_7142,N_5831,N_5748);
nor U7143 (N_7143,N_5511,N_4043);
nor U7144 (N_7144,N_5597,N_5589);
xor U7145 (N_7145,N_5087,N_5608);
xnor U7146 (N_7146,N_4975,N_5841);
or U7147 (N_7147,N_4088,N_5296);
or U7148 (N_7148,N_4046,N_4859);
nor U7149 (N_7149,N_5323,N_4182);
nor U7150 (N_7150,N_5237,N_4557);
xnor U7151 (N_7151,N_5632,N_5839);
xnor U7152 (N_7152,N_4407,N_4016);
or U7153 (N_7153,N_4433,N_5251);
xnor U7154 (N_7154,N_5564,N_4753);
or U7155 (N_7155,N_4621,N_4245);
or U7156 (N_7156,N_4440,N_5549);
or U7157 (N_7157,N_5308,N_4211);
nor U7158 (N_7158,N_5533,N_5506);
nand U7159 (N_7159,N_5423,N_4354);
nand U7160 (N_7160,N_4063,N_5438);
or U7161 (N_7161,N_4618,N_5000);
nand U7162 (N_7162,N_5038,N_4870);
and U7163 (N_7163,N_5378,N_5723);
nor U7164 (N_7164,N_5176,N_5599);
and U7165 (N_7165,N_5924,N_4349);
nand U7166 (N_7166,N_4223,N_5431);
xnor U7167 (N_7167,N_5376,N_4631);
nand U7168 (N_7168,N_4680,N_4318);
nand U7169 (N_7169,N_4797,N_5938);
or U7170 (N_7170,N_4776,N_4666);
nand U7171 (N_7171,N_4276,N_5524);
nor U7172 (N_7172,N_5427,N_5218);
xor U7173 (N_7173,N_4481,N_5702);
or U7174 (N_7174,N_5453,N_4252);
and U7175 (N_7175,N_4193,N_4169);
or U7176 (N_7176,N_5990,N_4963);
or U7177 (N_7177,N_4932,N_4049);
xnor U7178 (N_7178,N_5027,N_4334);
xor U7179 (N_7179,N_5406,N_5071);
xnor U7180 (N_7180,N_5997,N_5134);
nor U7181 (N_7181,N_4312,N_5599);
nand U7182 (N_7182,N_5122,N_5063);
or U7183 (N_7183,N_5660,N_5273);
and U7184 (N_7184,N_5678,N_5994);
and U7185 (N_7185,N_4404,N_4802);
xor U7186 (N_7186,N_4722,N_4687);
nor U7187 (N_7187,N_5909,N_5344);
or U7188 (N_7188,N_5796,N_4250);
nand U7189 (N_7189,N_5289,N_4908);
and U7190 (N_7190,N_4735,N_5783);
xnor U7191 (N_7191,N_4947,N_5131);
xor U7192 (N_7192,N_4674,N_4121);
xor U7193 (N_7193,N_4228,N_5027);
nand U7194 (N_7194,N_5432,N_5615);
nor U7195 (N_7195,N_5754,N_5232);
nand U7196 (N_7196,N_4996,N_5875);
and U7197 (N_7197,N_4892,N_5301);
nand U7198 (N_7198,N_4784,N_5775);
or U7199 (N_7199,N_4434,N_4757);
nor U7200 (N_7200,N_4461,N_4939);
and U7201 (N_7201,N_5202,N_5847);
xnor U7202 (N_7202,N_5211,N_5301);
nor U7203 (N_7203,N_5220,N_5387);
and U7204 (N_7204,N_4594,N_5350);
xor U7205 (N_7205,N_4800,N_5996);
xnor U7206 (N_7206,N_5795,N_5184);
nand U7207 (N_7207,N_4096,N_5879);
nand U7208 (N_7208,N_4205,N_5862);
and U7209 (N_7209,N_4698,N_5075);
or U7210 (N_7210,N_4506,N_5382);
nand U7211 (N_7211,N_4360,N_4516);
nand U7212 (N_7212,N_4144,N_5691);
nand U7213 (N_7213,N_5084,N_5232);
nor U7214 (N_7214,N_4634,N_5135);
or U7215 (N_7215,N_5097,N_4873);
or U7216 (N_7216,N_5536,N_5904);
or U7217 (N_7217,N_5799,N_5034);
nor U7218 (N_7218,N_5392,N_5101);
nor U7219 (N_7219,N_5492,N_4242);
xnor U7220 (N_7220,N_5773,N_5438);
or U7221 (N_7221,N_5206,N_4961);
xnor U7222 (N_7222,N_5716,N_4179);
nor U7223 (N_7223,N_5079,N_4448);
nor U7224 (N_7224,N_4230,N_5651);
or U7225 (N_7225,N_5675,N_4476);
nand U7226 (N_7226,N_4206,N_4386);
nand U7227 (N_7227,N_5717,N_5255);
or U7228 (N_7228,N_4003,N_5880);
nor U7229 (N_7229,N_4250,N_5571);
or U7230 (N_7230,N_5998,N_4604);
xnor U7231 (N_7231,N_5786,N_4705);
and U7232 (N_7232,N_4690,N_5957);
or U7233 (N_7233,N_5262,N_4108);
xnor U7234 (N_7234,N_4648,N_5527);
nand U7235 (N_7235,N_5190,N_4945);
nand U7236 (N_7236,N_5256,N_4268);
xor U7237 (N_7237,N_4090,N_5879);
nand U7238 (N_7238,N_4092,N_4094);
nand U7239 (N_7239,N_4316,N_4260);
xnor U7240 (N_7240,N_5673,N_4568);
nor U7241 (N_7241,N_4385,N_4815);
and U7242 (N_7242,N_5914,N_4123);
or U7243 (N_7243,N_5729,N_4306);
nor U7244 (N_7244,N_5640,N_5480);
nor U7245 (N_7245,N_5509,N_5204);
nand U7246 (N_7246,N_5927,N_4251);
nand U7247 (N_7247,N_5171,N_4111);
nand U7248 (N_7248,N_4315,N_4472);
xor U7249 (N_7249,N_5887,N_4505);
and U7250 (N_7250,N_5731,N_4322);
xor U7251 (N_7251,N_4608,N_4694);
xnor U7252 (N_7252,N_4172,N_5156);
xnor U7253 (N_7253,N_4847,N_5188);
or U7254 (N_7254,N_4611,N_5600);
and U7255 (N_7255,N_5533,N_5155);
and U7256 (N_7256,N_4067,N_4445);
nor U7257 (N_7257,N_4765,N_4738);
nor U7258 (N_7258,N_4671,N_4154);
xnor U7259 (N_7259,N_5085,N_5490);
nand U7260 (N_7260,N_5105,N_4906);
and U7261 (N_7261,N_4167,N_5244);
nand U7262 (N_7262,N_4511,N_4926);
or U7263 (N_7263,N_5638,N_4852);
or U7264 (N_7264,N_4398,N_4810);
or U7265 (N_7265,N_5246,N_4365);
or U7266 (N_7266,N_5372,N_4529);
nand U7267 (N_7267,N_4155,N_4018);
nand U7268 (N_7268,N_4476,N_5790);
nor U7269 (N_7269,N_4921,N_5194);
and U7270 (N_7270,N_4226,N_5612);
nor U7271 (N_7271,N_4813,N_5606);
xnor U7272 (N_7272,N_4158,N_4898);
or U7273 (N_7273,N_4058,N_4186);
nor U7274 (N_7274,N_5030,N_5590);
nor U7275 (N_7275,N_5041,N_4814);
nor U7276 (N_7276,N_4022,N_4436);
nor U7277 (N_7277,N_5743,N_5836);
nor U7278 (N_7278,N_5757,N_5816);
xnor U7279 (N_7279,N_5631,N_5744);
nand U7280 (N_7280,N_4201,N_5624);
xnor U7281 (N_7281,N_5161,N_4581);
nand U7282 (N_7282,N_4662,N_4296);
and U7283 (N_7283,N_5804,N_5110);
nand U7284 (N_7284,N_4536,N_4516);
and U7285 (N_7285,N_5106,N_4926);
nor U7286 (N_7286,N_4654,N_4856);
and U7287 (N_7287,N_5609,N_5592);
nand U7288 (N_7288,N_5627,N_4943);
or U7289 (N_7289,N_4545,N_5439);
xnor U7290 (N_7290,N_5944,N_5327);
nand U7291 (N_7291,N_4133,N_5406);
and U7292 (N_7292,N_4342,N_5061);
nor U7293 (N_7293,N_5201,N_5884);
nand U7294 (N_7294,N_5398,N_5239);
nand U7295 (N_7295,N_4491,N_5328);
nand U7296 (N_7296,N_5562,N_5044);
nand U7297 (N_7297,N_4161,N_4492);
and U7298 (N_7298,N_5270,N_4824);
and U7299 (N_7299,N_4818,N_5024);
nand U7300 (N_7300,N_5726,N_4230);
and U7301 (N_7301,N_5574,N_5732);
and U7302 (N_7302,N_5712,N_4229);
or U7303 (N_7303,N_4930,N_4254);
xnor U7304 (N_7304,N_4289,N_4458);
xor U7305 (N_7305,N_5982,N_4113);
nand U7306 (N_7306,N_4823,N_5258);
and U7307 (N_7307,N_4318,N_5137);
and U7308 (N_7308,N_4310,N_4623);
and U7309 (N_7309,N_4583,N_4050);
or U7310 (N_7310,N_4760,N_5220);
nand U7311 (N_7311,N_4013,N_5803);
or U7312 (N_7312,N_4955,N_5511);
or U7313 (N_7313,N_5563,N_4904);
and U7314 (N_7314,N_4176,N_5576);
and U7315 (N_7315,N_4541,N_5369);
nand U7316 (N_7316,N_5533,N_4892);
or U7317 (N_7317,N_4879,N_4664);
nor U7318 (N_7318,N_4652,N_4854);
and U7319 (N_7319,N_5154,N_4879);
nand U7320 (N_7320,N_5580,N_5093);
and U7321 (N_7321,N_4968,N_4778);
nor U7322 (N_7322,N_5416,N_4534);
or U7323 (N_7323,N_5654,N_5703);
nand U7324 (N_7324,N_5281,N_4860);
nand U7325 (N_7325,N_5011,N_4994);
nand U7326 (N_7326,N_5033,N_5685);
nand U7327 (N_7327,N_4014,N_5544);
xor U7328 (N_7328,N_4572,N_4285);
nand U7329 (N_7329,N_5201,N_5048);
nor U7330 (N_7330,N_4086,N_5321);
nor U7331 (N_7331,N_4378,N_4219);
and U7332 (N_7332,N_5891,N_4979);
and U7333 (N_7333,N_4113,N_5534);
nor U7334 (N_7334,N_4604,N_4629);
nor U7335 (N_7335,N_5324,N_5406);
or U7336 (N_7336,N_5429,N_4115);
nor U7337 (N_7337,N_5477,N_4524);
nand U7338 (N_7338,N_4493,N_5702);
and U7339 (N_7339,N_5135,N_5005);
and U7340 (N_7340,N_4051,N_4150);
and U7341 (N_7341,N_4743,N_4663);
xor U7342 (N_7342,N_5289,N_5858);
and U7343 (N_7343,N_4514,N_4272);
nand U7344 (N_7344,N_5123,N_5665);
or U7345 (N_7345,N_4148,N_5288);
and U7346 (N_7346,N_5594,N_4895);
xor U7347 (N_7347,N_5287,N_5425);
nand U7348 (N_7348,N_4234,N_5831);
and U7349 (N_7349,N_4515,N_4119);
nor U7350 (N_7350,N_4846,N_4905);
and U7351 (N_7351,N_4747,N_5467);
and U7352 (N_7352,N_5689,N_5931);
or U7353 (N_7353,N_5205,N_4458);
or U7354 (N_7354,N_5994,N_4539);
or U7355 (N_7355,N_4507,N_5647);
and U7356 (N_7356,N_4965,N_5093);
and U7357 (N_7357,N_5626,N_5870);
nor U7358 (N_7358,N_4989,N_5623);
nor U7359 (N_7359,N_5339,N_4546);
nor U7360 (N_7360,N_4239,N_4325);
nor U7361 (N_7361,N_4740,N_4160);
nand U7362 (N_7362,N_5981,N_5610);
nor U7363 (N_7363,N_5317,N_4505);
or U7364 (N_7364,N_4253,N_4897);
and U7365 (N_7365,N_5014,N_4592);
nor U7366 (N_7366,N_5152,N_5902);
xnor U7367 (N_7367,N_4503,N_4110);
nor U7368 (N_7368,N_4723,N_5775);
and U7369 (N_7369,N_5522,N_4287);
nand U7370 (N_7370,N_4820,N_5387);
xor U7371 (N_7371,N_4498,N_5509);
nor U7372 (N_7372,N_4246,N_5423);
nand U7373 (N_7373,N_4390,N_4227);
nor U7374 (N_7374,N_4141,N_5402);
or U7375 (N_7375,N_4400,N_4542);
or U7376 (N_7376,N_5270,N_4223);
nor U7377 (N_7377,N_4308,N_5712);
nand U7378 (N_7378,N_4746,N_4221);
and U7379 (N_7379,N_5188,N_5395);
or U7380 (N_7380,N_4606,N_4556);
or U7381 (N_7381,N_5558,N_4185);
xnor U7382 (N_7382,N_4701,N_5518);
nor U7383 (N_7383,N_4452,N_5651);
xnor U7384 (N_7384,N_5238,N_5130);
nand U7385 (N_7385,N_4410,N_5094);
or U7386 (N_7386,N_4372,N_5525);
and U7387 (N_7387,N_4713,N_5234);
xnor U7388 (N_7388,N_4966,N_5148);
nor U7389 (N_7389,N_5651,N_4384);
and U7390 (N_7390,N_5399,N_4585);
or U7391 (N_7391,N_4158,N_4704);
or U7392 (N_7392,N_5740,N_4056);
xor U7393 (N_7393,N_5509,N_4509);
nand U7394 (N_7394,N_5153,N_4320);
nor U7395 (N_7395,N_4961,N_5687);
and U7396 (N_7396,N_4324,N_5556);
nand U7397 (N_7397,N_4771,N_5295);
xor U7398 (N_7398,N_4712,N_4238);
nor U7399 (N_7399,N_4634,N_5196);
or U7400 (N_7400,N_4511,N_5352);
xor U7401 (N_7401,N_5312,N_4323);
nand U7402 (N_7402,N_4473,N_4421);
nand U7403 (N_7403,N_5803,N_5958);
nor U7404 (N_7404,N_4628,N_4111);
and U7405 (N_7405,N_4858,N_4112);
or U7406 (N_7406,N_5782,N_5662);
or U7407 (N_7407,N_5269,N_5498);
or U7408 (N_7408,N_5801,N_5539);
or U7409 (N_7409,N_5068,N_5835);
nor U7410 (N_7410,N_5654,N_5729);
xor U7411 (N_7411,N_4057,N_4058);
or U7412 (N_7412,N_5734,N_4547);
nor U7413 (N_7413,N_5704,N_4207);
or U7414 (N_7414,N_4396,N_4753);
or U7415 (N_7415,N_5750,N_5838);
nand U7416 (N_7416,N_4454,N_4215);
xor U7417 (N_7417,N_4427,N_4788);
and U7418 (N_7418,N_4612,N_4231);
nor U7419 (N_7419,N_5091,N_5768);
nor U7420 (N_7420,N_5655,N_5548);
nand U7421 (N_7421,N_4718,N_5007);
or U7422 (N_7422,N_4097,N_4279);
xor U7423 (N_7423,N_5459,N_5659);
or U7424 (N_7424,N_5619,N_5587);
nand U7425 (N_7425,N_5577,N_5372);
and U7426 (N_7426,N_5794,N_4560);
xnor U7427 (N_7427,N_5389,N_5218);
xnor U7428 (N_7428,N_4992,N_5139);
nand U7429 (N_7429,N_4939,N_4853);
and U7430 (N_7430,N_4414,N_4025);
and U7431 (N_7431,N_5398,N_5941);
or U7432 (N_7432,N_4103,N_5922);
nor U7433 (N_7433,N_4098,N_4120);
nand U7434 (N_7434,N_5734,N_4071);
nand U7435 (N_7435,N_4460,N_4791);
or U7436 (N_7436,N_4277,N_4106);
nand U7437 (N_7437,N_5752,N_5071);
or U7438 (N_7438,N_5532,N_4138);
or U7439 (N_7439,N_5328,N_5106);
nand U7440 (N_7440,N_4770,N_5307);
and U7441 (N_7441,N_4055,N_4798);
and U7442 (N_7442,N_5510,N_5810);
xnor U7443 (N_7443,N_5337,N_4556);
nand U7444 (N_7444,N_4618,N_5558);
and U7445 (N_7445,N_5276,N_4199);
nand U7446 (N_7446,N_4093,N_5294);
nor U7447 (N_7447,N_4287,N_5660);
nand U7448 (N_7448,N_4183,N_4572);
and U7449 (N_7449,N_4350,N_4839);
nor U7450 (N_7450,N_4569,N_5594);
nor U7451 (N_7451,N_4337,N_5584);
or U7452 (N_7452,N_4393,N_5885);
and U7453 (N_7453,N_5123,N_5505);
and U7454 (N_7454,N_5974,N_4474);
or U7455 (N_7455,N_5543,N_5125);
nand U7456 (N_7456,N_5749,N_5174);
and U7457 (N_7457,N_4429,N_4483);
or U7458 (N_7458,N_5965,N_5087);
or U7459 (N_7459,N_4085,N_4573);
or U7460 (N_7460,N_5894,N_5059);
nor U7461 (N_7461,N_4030,N_4527);
nand U7462 (N_7462,N_4492,N_4766);
and U7463 (N_7463,N_5827,N_4930);
and U7464 (N_7464,N_5496,N_4000);
or U7465 (N_7465,N_4073,N_5446);
or U7466 (N_7466,N_5748,N_5049);
and U7467 (N_7467,N_4389,N_5274);
xor U7468 (N_7468,N_4166,N_4283);
xnor U7469 (N_7469,N_5171,N_4847);
nor U7470 (N_7470,N_4140,N_4835);
or U7471 (N_7471,N_5332,N_4737);
nor U7472 (N_7472,N_4372,N_5962);
xnor U7473 (N_7473,N_4282,N_4877);
and U7474 (N_7474,N_4675,N_4563);
nand U7475 (N_7475,N_4908,N_4862);
and U7476 (N_7476,N_5586,N_4261);
or U7477 (N_7477,N_4647,N_5617);
nor U7478 (N_7478,N_4842,N_5203);
and U7479 (N_7479,N_5075,N_5406);
or U7480 (N_7480,N_5866,N_5156);
nor U7481 (N_7481,N_4843,N_4376);
nor U7482 (N_7482,N_4914,N_5640);
nor U7483 (N_7483,N_5007,N_5825);
xnor U7484 (N_7484,N_5031,N_4347);
xnor U7485 (N_7485,N_5117,N_5441);
nand U7486 (N_7486,N_4296,N_5529);
or U7487 (N_7487,N_5167,N_5451);
xnor U7488 (N_7488,N_4007,N_4926);
nand U7489 (N_7489,N_4342,N_4341);
nor U7490 (N_7490,N_4350,N_4461);
or U7491 (N_7491,N_5300,N_4913);
nor U7492 (N_7492,N_5549,N_4407);
and U7493 (N_7493,N_4966,N_4829);
and U7494 (N_7494,N_4109,N_5147);
or U7495 (N_7495,N_4266,N_5929);
xnor U7496 (N_7496,N_5836,N_5027);
and U7497 (N_7497,N_5042,N_5919);
and U7498 (N_7498,N_4253,N_4184);
nand U7499 (N_7499,N_5573,N_4786);
nand U7500 (N_7500,N_5821,N_5172);
xnor U7501 (N_7501,N_5871,N_5336);
xnor U7502 (N_7502,N_4665,N_5299);
nand U7503 (N_7503,N_4346,N_4172);
nand U7504 (N_7504,N_4182,N_4869);
and U7505 (N_7505,N_5399,N_4626);
and U7506 (N_7506,N_4216,N_4816);
nand U7507 (N_7507,N_5130,N_4309);
and U7508 (N_7508,N_5861,N_5663);
nor U7509 (N_7509,N_5686,N_5822);
xor U7510 (N_7510,N_5305,N_4323);
or U7511 (N_7511,N_4347,N_4442);
xnor U7512 (N_7512,N_5360,N_5733);
xnor U7513 (N_7513,N_4609,N_5779);
nand U7514 (N_7514,N_5171,N_5901);
nand U7515 (N_7515,N_4842,N_5799);
nand U7516 (N_7516,N_5022,N_5405);
or U7517 (N_7517,N_4226,N_4244);
or U7518 (N_7518,N_4296,N_4454);
or U7519 (N_7519,N_5459,N_4127);
nor U7520 (N_7520,N_4816,N_5594);
nor U7521 (N_7521,N_4514,N_4758);
xor U7522 (N_7522,N_5942,N_5831);
or U7523 (N_7523,N_4779,N_4623);
nor U7524 (N_7524,N_4479,N_5461);
and U7525 (N_7525,N_5830,N_4936);
xor U7526 (N_7526,N_5545,N_5072);
nor U7527 (N_7527,N_4149,N_4650);
nor U7528 (N_7528,N_5659,N_4806);
and U7529 (N_7529,N_4297,N_5404);
nand U7530 (N_7530,N_4406,N_4453);
and U7531 (N_7531,N_4720,N_4977);
xnor U7532 (N_7532,N_4077,N_4174);
xnor U7533 (N_7533,N_4227,N_4369);
nor U7534 (N_7534,N_4794,N_4479);
nor U7535 (N_7535,N_4429,N_5856);
xor U7536 (N_7536,N_4367,N_4371);
and U7537 (N_7537,N_4953,N_5519);
and U7538 (N_7538,N_4132,N_4390);
or U7539 (N_7539,N_5914,N_4818);
or U7540 (N_7540,N_4529,N_5019);
nor U7541 (N_7541,N_4969,N_5504);
or U7542 (N_7542,N_4969,N_5552);
xor U7543 (N_7543,N_5003,N_5041);
or U7544 (N_7544,N_4568,N_5450);
and U7545 (N_7545,N_5420,N_4947);
nor U7546 (N_7546,N_4383,N_4828);
nand U7547 (N_7547,N_4341,N_4304);
nor U7548 (N_7548,N_5377,N_4641);
nand U7549 (N_7549,N_4334,N_5656);
or U7550 (N_7550,N_4316,N_5413);
nand U7551 (N_7551,N_5711,N_5777);
nor U7552 (N_7552,N_4602,N_4961);
nand U7553 (N_7553,N_4468,N_4374);
nor U7554 (N_7554,N_5442,N_5525);
nand U7555 (N_7555,N_5547,N_5241);
nand U7556 (N_7556,N_5432,N_5727);
and U7557 (N_7557,N_4397,N_5361);
or U7558 (N_7558,N_4963,N_4529);
nand U7559 (N_7559,N_5710,N_4352);
nor U7560 (N_7560,N_4192,N_5237);
and U7561 (N_7561,N_5085,N_4755);
and U7562 (N_7562,N_4302,N_5186);
nand U7563 (N_7563,N_4943,N_4934);
nand U7564 (N_7564,N_5879,N_4024);
nand U7565 (N_7565,N_5760,N_5985);
nand U7566 (N_7566,N_5486,N_4942);
xnor U7567 (N_7567,N_4119,N_4863);
or U7568 (N_7568,N_4550,N_4047);
nor U7569 (N_7569,N_4717,N_5602);
xor U7570 (N_7570,N_4448,N_4297);
and U7571 (N_7571,N_4270,N_5454);
nand U7572 (N_7572,N_5271,N_5660);
or U7573 (N_7573,N_5078,N_4303);
or U7574 (N_7574,N_5173,N_5995);
or U7575 (N_7575,N_4785,N_4196);
or U7576 (N_7576,N_5447,N_4149);
and U7577 (N_7577,N_5642,N_4774);
nand U7578 (N_7578,N_4426,N_4876);
or U7579 (N_7579,N_4058,N_4232);
nand U7580 (N_7580,N_4327,N_4761);
or U7581 (N_7581,N_5759,N_5168);
and U7582 (N_7582,N_5428,N_4038);
or U7583 (N_7583,N_4409,N_5403);
nand U7584 (N_7584,N_4596,N_5284);
nor U7585 (N_7585,N_4075,N_5395);
nand U7586 (N_7586,N_4912,N_5663);
nand U7587 (N_7587,N_5786,N_4758);
xnor U7588 (N_7588,N_5076,N_4502);
and U7589 (N_7589,N_5280,N_5018);
or U7590 (N_7590,N_4828,N_5191);
xnor U7591 (N_7591,N_5375,N_4244);
nor U7592 (N_7592,N_5614,N_4278);
nand U7593 (N_7593,N_4232,N_5376);
or U7594 (N_7594,N_4255,N_4081);
nand U7595 (N_7595,N_4884,N_5916);
nor U7596 (N_7596,N_5904,N_5038);
and U7597 (N_7597,N_4129,N_5898);
and U7598 (N_7598,N_4468,N_5693);
or U7599 (N_7599,N_4205,N_5697);
or U7600 (N_7600,N_4024,N_4875);
or U7601 (N_7601,N_4367,N_5673);
xor U7602 (N_7602,N_5959,N_5844);
xor U7603 (N_7603,N_5731,N_5494);
xor U7604 (N_7604,N_4382,N_4190);
or U7605 (N_7605,N_4976,N_4362);
or U7606 (N_7606,N_5053,N_4543);
nor U7607 (N_7607,N_5696,N_5123);
or U7608 (N_7608,N_4047,N_4083);
nand U7609 (N_7609,N_5353,N_5741);
xnor U7610 (N_7610,N_5189,N_5046);
and U7611 (N_7611,N_4022,N_5189);
xnor U7612 (N_7612,N_5966,N_4212);
nor U7613 (N_7613,N_5169,N_4653);
nor U7614 (N_7614,N_4855,N_4698);
xnor U7615 (N_7615,N_4433,N_5897);
and U7616 (N_7616,N_4712,N_4182);
nand U7617 (N_7617,N_4705,N_5675);
nand U7618 (N_7618,N_4991,N_4974);
xor U7619 (N_7619,N_5855,N_4326);
nor U7620 (N_7620,N_4650,N_4146);
or U7621 (N_7621,N_4770,N_4213);
or U7622 (N_7622,N_5004,N_5563);
xor U7623 (N_7623,N_4942,N_5737);
nand U7624 (N_7624,N_5423,N_4762);
nor U7625 (N_7625,N_5694,N_5692);
nand U7626 (N_7626,N_4514,N_4699);
and U7627 (N_7627,N_4123,N_5228);
nand U7628 (N_7628,N_4230,N_5634);
or U7629 (N_7629,N_4422,N_5105);
and U7630 (N_7630,N_4849,N_4742);
nor U7631 (N_7631,N_4025,N_5400);
or U7632 (N_7632,N_4117,N_5252);
nand U7633 (N_7633,N_4279,N_4645);
and U7634 (N_7634,N_5852,N_4670);
nor U7635 (N_7635,N_5434,N_5568);
and U7636 (N_7636,N_4911,N_5374);
or U7637 (N_7637,N_4562,N_5892);
or U7638 (N_7638,N_4773,N_5424);
or U7639 (N_7639,N_5597,N_5868);
or U7640 (N_7640,N_4644,N_5510);
or U7641 (N_7641,N_4582,N_4452);
nor U7642 (N_7642,N_4303,N_4263);
nand U7643 (N_7643,N_4636,N_4339);
and U7644 (N_7644,N_4889,N_4710);
nand U7645 (N_7645,N_4668,N_5672);
nor U7646 (N_7646,N_5745,N_4172);
and U7647 (N_7647,N_4824,N_4949);
and U7648 (N_7648,N_5798,N_4150);
xnor U7649 (N_7649,N_5124,N_4645);
xnor U7650 (N_7650,N_4974,N_5532);
nand U7651 (N_7651,N_5748,N_4948);
xnor U7652 (N_7652,N_5403,N_4389);
and U7653 (N_7653,N_5265,N_4064);
or U7654 (N_7654,N_5994,N_5991);
or U7655 (N_7655,N_5619,N_5458);
and U7656 (N_7656,N_5047,N_4501);
xor U7657 (N_7657,N_4209,N_5839);
nand U7658 (N_7658,N_5857,N_4190);
and U7659 (N_7659,N_4267,N_5811);
nor U7660 (N_7660,N_5600,N_4216);
xor U7661 (N_7661,N_4993,N_5568);
or U7662 (N_7662,N_5573,N_5928);
nand U7663 (N_7663,N_4450,N_5067);
or U7664 (N_7664,N_4316,N_4080);
and U7665 (N_7665,N_5953,N_4120);
xnor U7666 (N_7666,N_4235,N_5469);
xor U7667 (N_7667,N_5290,N_4923);
or U7668 (N_7668,N_4273,N_5181);
or U7669 (N_7669,N_4547,N_4653);
nor U7670 (N_7670,N_5476,N_4791);
and U7671 (N_7671,N_4492,N_5172);
or U7672 (N_7672,N_4646,N_4501);
nor U7673 (N_7673,N_5275,N_5001);
xnor U7674 (N_7674,N_5976,N_5362);
xnor U7675 (N_7675,N_4854,N_4261);
xnor U7676 (N_7676,N_5259,N_4175);
nor U7677 (N_7677,N_4332,N_5399);
or U7678 (N_7678,N_4222,N_4359);
nor U7679 (N_7679,N_4153,N_5272);
xnor U7680 (N_7680,N_5510,N_5383);
nand U7681 (N_7681,N_4697,N_4489);
and U7682 (N_7682,N_5670,N_5254);
or U7683 (N_7683,N_4796,N_4079);
or U7684 (N_7684,N_5402,N_4703);
nand U7685 (N_7685,N_4218,N_5966);
and U7686 (N_7686,N_5267,N_5396);
and U7687 (N_7687,N_5555,N_4471);
or U7688 (N_7688,N_4575,N_5614);
nand U7689 (N_7689,N_4063,N_4650);
and U7690 (N_7690,N_5369,N_4291);
nor U7691 (N_7691,N_5274,N_4890);
or U7692 (N_7692,N_5756,N_4308);
nor U7693 (N_7693,N_4353,N_5566);
and U7694 (N_7694,N_5063,N_4179);
and U7695 (N_7695,N_4482,N_5693);
nor U7696 (N_7696,N_4172,N_4877);
nor U7697 (N_7697,N_5496,N_4772);
nand U7698 (N_7698,N_4176,N_4179);
and U7699 (N_7699,N_4787,N_5428);
nor U7700 (N_7700,N_5842,N_4621);
nand U7701 (N_7701,N_4466,N_5845);
nand U7702 (N_7702,N_5420,N_4431);
or U7703 (N_7703,N_5832,N_4197);
or U7704 (N_7704,N_4576,N_4509);
nor U7705 (N_7705,N_4968,N_5838);
nand U7706 (N_7706,N_4808,N_4639);
nand U7707 (N_7707,N_5072,N_5884);
and U7708 (N_7708,N_5288,N_5657);
and U7709 (N_7709,N_5071,N_5185);
and U7710 (N_7710,N_4800,N_5619);
nor U7711 (N_7711,N_4199,N_5822);
nor U7712 (N_7712,N_4060,N_4805);
nor U7713 (N_7713,N_5304,N_4298);
or U7714 (N_7714,N_4774,N_5845);
nor U7715 (N_7715,N_4397,N_5980);
or U7716 (N_7716,N_5236,N_5338);
and U7717 (N_7717,N_5634,N_4679);
nand U7718 (N_7718,N_4355,N_4650);
xor U7719 (N_7719,N_4560,N_4183);
xnor U7720 (N_7720,N_4805,N_4020);
nand U7721 (N_7721,N_4971,N_4175);
nor U7722 (N_7722,N_4788,N_4940);
or U7723 (N_7723,N_4309,N_5804);
nor U7724 (N_7724,N_4556,N_4728);
nand U7725 (N_7725,N_4008,N_5318);
xor U7726 (N_7726,N_5554,N_4893);
xor U7727 (N_7727,N_5603,N_4265);
nor U7728 (N_7728,N_4927,N_5600);
xor U7729 (N_7729,N_5976,N_5406);
and U7730 (N_7730,N_4158,N_5028);
nand U7731 (N_7731,N_5552,N_4035);
nor U7732 (N_7732,N_5551,N_5646);
nand U7733 (N_7733,N_5238,N_4475);
xnor U7734 (N_7734,N_5493,N_5328);
nand U7735 (N_7735,N_5240,N_4623);
nor U7736 (N_7736,N_5644,N_4366);
nor U7737 (N_7737,N_5977,N_5371);
nor U7738 (N_7738,N_5091,N_5121);
or U7739 (N_7739,N_5300,N_5440);
and U7740 (N_7740,N_4574,N_5181);
xnor U7741 (N_7741,N_5581,N_5713);
xor U7742 (N_7742,N_5092,N_4595);
nor U7743 (N_7743,N_5309,N_4753);
nor U7744 (N_7744,N_4345,N_5198);
nand U7745 (N_7745,N_4797,N_5983);
xor U7746 (N_7746,N_5175,N_4941);
or U7747 (N_7747,N_4756,N_5894);
nor U7748 (N_7748,N_5596,N_5884);
xor U7749 (N_7749,N_4716,N_4178);
xnor U7750 (N_7750,N_4748,N_4449);
and U7751 (N_7751,N_5522,N_4726);
and U7752 (N_7752,N_4825,N_5785);
nor U7753 (N_7753,N_5797,N_5801);
or U7754 (N_7754,N_5137,N_4774);
nand U7755 (N_7755,N_4359,N_5452);
or U7756 (N_7756,N_4205,N_5770);
or U7757 (N_7757,N_4694,N_4540);
nor U7758 (N_7758,N_4512,N_5791);
nand U7759 (N_7759,N_4286,N_5909);
nor U7760 (N_7760,N_5052,N_4003);
or U7761 (N_7761,N_5017,N_5670);
and U7762 (N_7762,N_5758,N_4890);
and U7763 (N_7763,N_4388,N_5004);
and U7764 (N_7764,N_4192,N_5943);
nand U7765 (N_7765,N_4361,N_5721);
xnor U7766 (N_7766,N_5366,N_4951);
xnor U7767 (N_7767,N_4350,N_5056);
nand U7768 (N_7768,N_5468,N_4798);
xor U7769 (N_7769,N_5100,N_4351);
and U7770 (N_7770,N_5319,N_4144);
nor U7771 (N_7771,N_5273,N_4946);
or U7772 (N_7772,N_4618,N_4682);
or U7773 (N_7773,N_5700,N_4320);
nand U7774 (N_7774,N_4566,N_5785);
nand U7775 (N_7775,N_5717,N_5544);
nor U7776 (N_7776,N_5790,N_4775);
nand U7777 (N_7777,N_4432,N_5561);
nand U7778 (N_7778,N_5319,N_5920);
or U7779 (N_7779,N_5490,N_4577);
nor U7780 (N_7780,N_4552,N_4294);
or U7781 (N_7781,N_4851,N_4297);
nand U7782 (N_7782,N_5574,N_5595);
and U7783 (N_7783,N_4054,N_5793);
or U7784 (N_7784,N_5882,N_4595);
xnor U7785 (N_7785,N_5261,N_5724);
nor U7786 (N_7786,N_5694,N_5950);
nor U7787 (N_7787,N_4873,N_5316);
nor U7788 (N_7788,N_4477,N_4944);
nand U7789 (N_7789,N_4280,N_5129);
nand U7790 (N_7790,N_5036,N_5601);
nand U7791 (N_7791,N_5235,N_4968);
and U7792 (N_7792,N_5887,N_4267);
xor U7793 (N_7793,N_5113,N_5505);
nand U7794 (N_7794,N_5783,N_4322);
xnor U7795 (N_7795,N_5550,N_5534);
nand U7796 (N_7796,N_5607,N_5345);
or U7797 (N_7797,N_5950,N_5507);
and U7798 (N_7798,N_4031,N_4117);
nand U7799 (N_7799,N_5520,N_4965);
nand U7800 (N_7800,N_4946,N_4335);
nand U7801 (N_7801,N_5528,N_5864);
and U7802 (N_7802,N_5117,N_4119);
and U7803 (N_7803,N_5538,N_5035);
or U7804 (N_7804,N_4295,N_4519);
and U7805 (N_7805,N_4018,N_4236);
nor U7806 (N_7806,N_4380,N_5631);
xnor U7807 (N_7807,N_4054,N_4798);
and U7808 (N_7808,N_4368,N_4763);
or U7809 (N_7809,N_5031,N_4835);
nor U7810 (N_7810,N_5387,N_4292);
nor U7811 (N_7811,N_5901,N_4233);
xnor U7812 (N_7812,N_5446,N_5598);
or U7813 (N_7813,N_5470,N_4189);
xnor U7814 (N_7814,N_4562,N_4981);
nand U7815 (N_7815,N_5019,N_4211);
xor U7816 (N_7816,N_4199,N_5975);
or U7817 (N_7817,N_5862,N_5136);
nand U7818 (N_7818,N_5506,N_4606);
or U7819 (N_7819,N_4657,N_5066);
or U7820 (N_7820,N_5798,N_4099);
xor U7821 (N_7821,N_5117,N_4978);
or U7822 (N_7822,N_5296,N_5997);
and U7823 (N_7823,N_5455,N_5404);
or U7824 (N_7824,N_4833,N_4949);
and U7825 (N_7825,N_4713,N_4809);
and U7826 (N_7826,N_4751,N_5202);
xnor U7827 (N_7827,N_5032,N_4360);
and U7828 (N_7828,N_4781,N_4078);
or U7829 (N_7829,N_5243,N_4373);
and U7830 (N_7830,N_4372,N_4314);
nand U7831 (N_7831,N_5999,N_4416);
or U7832 (N_7832,N_4744,N_5353);
xnor U7833 (N_7833,N_4122,N_4592);
and U7834 (N_7834,N_4468,N_4731);
xnor U7835 (N_7835,N_4445,N_5172);
or U7836 (N_7836,N_4687,N_4198);
and U7837 (N_7837,N_4119,N_5910);
nand U7838 (N_7838,N_4275,N_4257);
nand U7839 (N_7839,N_4759,N_4931);
or U7840 (N_7840,N_4893,N_5452);
and U7841 (N_7841,N_5777,N_4164);
nand U7842 (N_7842,N_5299,N_5985);
nor U7843 (N_7843,N_5152,N_5930);
and U7844 (N_7844,N_4050,N_5307);
nand U7845 (N_7845,N_5666,N_5715);
and U7846 (N_7846,N_4985,N_5631);
nand U7847 (N_7847,N_5298,N_4984);
nand U7848 (N_7848,N_5392,N_4385);
or U7849 (N_7849,N_5305,N_4165);
xor U7850 (N_7850,N_5880,N_5658);
xnor U7851 (N_7851,N_4084,N_4629);
and U7852 (N_7852,N_4736,N_5877);
and U7853 (N_7853,N_4749,N_4704);
xnor U7854 (N_7854,N_4638,N_5935);
nand U7855 (N_7855,N_5906,N_5057);
or U7856 (N_7856,N_5678,N_5130);
nand U7857 (N_7857,N_4558,N_5693);
and U7858 (N_7858,N_5693,N_5596);
or U7859 (N_7859,N_5192,N_5927);
or U7860 (N_7860,N_4852,N_5400);
nor U7861 (N_7861,N_4842,N_4731);
nand U7862 (N_7862,N_4799,N_5961);
and U7863 (N_7863,N_5362,N_4474);
or U7864 (N_7864,N_4251,N_5659);
nand U7865 (N_7865,N_5102,N_5938);
and U7866 (N_7866,N_5014,N_4373);
nand U7867 (N_7867,N_5914,N_5093);
nor U7868 (N_7868,N_4428,N_5947);
nand U7869 (N_7869,N_4085,N_4946);
nand U7870 (N_7870,N_5118,N_4098);
or U7871 (N_7871,N_4436,N_5253);
nor U7872 (N_7872,N_4161,N_4107);
or U7873 (N_7873,N_5465,N_4820);
or U7874 (N_7874,N_5860,N_4616);
xnor U7875 (N_7875,N_5505,N_5960);
nor U7876 (N_7876,N_5229,N_5339);
nand U7877 (N_7877,N_4940,N_4942);
xor U7878 (N_7878,N_4690,N_4887);
nand U7879 (N_7879,N_5354,N_5740);
nand U7880 (N_7880,N_5151,N_5646);
or U7881 (N_7881,N_4826,N_5785);
or U7882 (N_7882,N_5056,N_4676);
nand U7883 (N_7883,N_4333,N_4775);
and U7884 (N_7884,N_5631,N_4102);
nand U7885 (N_7885,N_4611,N_4821);
nand U7886 (N_7886,N_4855,N_4091);
nand U7887 (N_7887,N_5698,N_5761);
nor U7888 (N_7888,N_5579,N_5077);
nor U7889 (N_7889,N_4972,N_5405);
nand U7890 (N_7890,N_5114,N_5758);
and U7891 (N_7891,N_5829,N_5238);
nand U7892 (N_7892,N_4240,N_4581);
nor U7893 (N_7893,N_4723,N_4437);
xor U7894 (N_7894,N_5351,N_5134);
nor U7895 (N_7895,N_5020,N_5249);
xor U7896 (N_7896,N_5461,N_5677);
nand U7897 (N_7897,N_4552,N_5923);
nand U7898 (N_7898,N_5275,N_5733);
xor U7899 (N_7899,N_5708,N_4518);
and U7900 (N_7900,N_5120,N_5690);
or U7901 (N_7901,N_4986,N_5740);
nor U7902 (N_7902,N_4511,N_4682);
and U7903 (N_7903,N_4215,N_4789);
nand U7904 (N_7904,N_4149,N_4789);
xor U7905 (N_7905,N_4283,N_4190);
nand U7906 (N_7906,N_4215,N_4854);
nand U7907 (N_7907,N_5995,N_4718);
nor U7908 (N_7908,N_4108,N_4117);
nand U7909 (N_7909,N_5843,N_4159);
and U7910 (N_7910,N_4963,N_4953);
xnor U7911 (N_7911,N_4520,N_4564);
and U7912 (N_7912,N_5013,N_5912);
and U7913 (N_7913,N_4899,N_4101);
nand U7914 (N_7914,N_5122,N_5612);
nor U7915 (N_7915,N_5029,N_4429);
nand U7916 (N_7916,N_4232,N_5596);
nand U7917 (N_7917,N_5871,N_5785);
or U7918 (N_7918,N_4284,N_4446);
nor U7919 (N_7919,N_5985,N_4411);
nor U7920 (N_7920,N_5160,N_4713);
nand U7921 (N_7921,N_5193,N_4589);
nand U7922 (N_7922,N_5129,N_4946);
or U7923 (N_7923,N_4763,N_5999);
nor U7924 (N_7924,N_5207,N_5552);
nand U7925 (N_7925,N_5671,N_4208);
nand U7926 (N_7926,N_5953,N_4071);
nor U7927 (N_7927,N_4283,N_4062);
nand U7928 (N_7928,N_4486,N_5409);
and U7929 (N_7929,N_5312,N_4953);
or U7930 (N_7930,N_5883,N_4221);
nand U7931 (N_7931,N_5922,N_4971);
and U7932 (N_7932,N_4181,N_5989);
nand U7933 (N_7933,N_4975,N_4275);
xor U7934 (N_7934,N_5807,N_4865);
nor U7935 (N_7935,N_4307,N_5777);
nor U7936 (N_7936,N_5135,N_4123);
or U7937 (N_7937,N_4175,N_4306);
xnor U7938 (N_7938,N_5126,N_5646);
nand U7939 (N_7939,N_4377,N_5819);
or U7940 (N_7940,N_4854,N_4552);
or U7941 (N_7941,N_4600,N_5432);
or U7942 (N_7942,N_5433,N_5393);
xnor U7943 (N_7943,N_4732,N_5612);
nor U7944 (N_7944,N_4220,N_5201);
nand U7945 (N_7945,N_4526,N_4706);
nor U7946 (N_7946,N_5359,N_4042);
or U7947 (N_7947,N_5722,N_4838);
or U7948 (N_7948,N_5541,N_5147);
xor U7949 (N_7949,N_5204,N_4245);
and U7950 (N_7950,N_5889,N_5642);
nor U7951 (N_7951,N_5288,N_4867);
nor U7952 (N_7952,N_4438,N_4805);
nor U7953 (N_7953,N_5627,N_5251);
nor U7954 (N_7954,N_4566,N_5528);
and U7955 (N_7955,N_5819,N_4427);
xor U7956 (N_7956,N_5308,N_4074);
nor U7957 (N_7957,N_4798,N_5225);
nor U7958 (N_7958,N_5290,N_5802);
nor U7959 (N_7959,N_5471,N_5109);
nand U7960 (N_7960,N_4341,N_5848);
xor U7961 (N_7961,N_5278,N_5495);
nand U7962 (N_7962,N_4630,N_5815);
nor U7963 (N_7963,N_4280,N_5492);
xnor U7964 (N_7964,N_4619,N_5650);
nor U7965 (N_7965,N_5423,N_4295);
nand U7966 (N_7966,N_5261,N_5867);
or U7967 (N_7967,N_4588,N_4786);
nand U7968 (N_7968,N_4282,N_5479);
nor U7969 (N_7969,N_4427,N_4350);
nand U7970 (N_7970,N_4804,N_5823);
nor U7971 (N_7971,N_5796,N_4128);
nand U7972 (N_7972,N_4533,N_4342);
nor U7973 (N_7973,N_5793,N_5152);
and U7974 (N_7974,N_5972,N_5616);
and U7975 (N_7975,N_4735,N_5208);
nand U7976 (N_7976,N_5336,N_4956);
or U7977 (N_7977,N_4719,N_4860);
and U7978 (N_7978,N_4873,N_4812);
or U7979 (N_7979,N_5941,N_4282);
nand U7980 (N_7980,N_5272,N_5479);
nor U7981 (N_7981,N_5204,N_4336);
and U7982 (N_7982,N_4645,N_5604);
or U7983 (N_7983,N_5236,N_4727);
xnor U7984 (N_7984,N_4541,N_5531);
and U7985 (N_7985,N_4030,N_5174);
nor U7986 (N_7986,N_5937,N_4570);
nor U7987 (N_7987,N_5143,N_4679);
and U7988 (N_7988,N_5059,N_4837);
and U7989 (N_7989,N_4619,N_4664);
nor U7990 (N_7990,N_5445,N_4352);
or U7991 (N_7991,N_5661,N_4974);
and U7992 (N_7992,N_4461,N_4164);
xnor U7993 (N_7993,N_4797,N_4555);
xor U7994 (N_7994,N_5021,N_4481);
xor U7995 (N_7995,N_4592,N_4560);
and U7996 (N_7996,N_4804,N_5694);
nand U7997 (N_7997,N_5112,N_4107);
and U7998 (N_7998,N_4884,N_4607);
or U7999 (N_7999,N_4561,N_5330);
nand U8000 (N_8000,N_7293,N_7021);
nor U8001 (N_8001,N_6385,N_6696);
xnor U8002 (N_8002,N_6555,N_7841);
and U8003 (N_8003,N_6827,N_7887);
or U8004 (N_8004,N_7644,N_6971);
or U8005 (N_8005,N_6624,N_7588);
nand U8006 (N_8006,N_7777,N_6714);
or U8007 (N_8007,N_7881,N_6300);
nor U8008 (N_8008,N_6351,N_6799);
nor U8009 (N_8009,N_6182,N_6665);
nand U8010 (N_8010,N_7194,N_6749);
nor U8011 (N_8011,N_7773,N_7082);
and U8012 (N_8012,N_7158,N_6109);
or U8013 (N_8013,N_6968,N_7381);
and U8014 (N_8014,N_7006,N_7675);
nand U8015 (N_8015,N_7579,N_6629);
nand U8016 (N_8016,N_6607,N_7778);
nand U8017 (N_8017,N_7134,N_7815);
xor U8018 (N_8018,N_7650,N_7418);
nor U8019 (N_8019,N_7272,N_7053);
nand U8020 (N_8020,N_7851,N_7958);
nor U8021 (N_8021,N_6908,N_7984);
or U8022 (N_8022,N_6259,N_7745);
and U8023 (N_8023,N_7485,N_7502);
nor U8024 (N_8024,N_6635,N_7942);
and U8025 (N_8025,N_6043,N_7700);
or U8026 (N_8026,N_6691,N_6783);
nor U8027 (N_8027,N_7446,N_6806);
nor U8028 (N_8028,N_6614,N_7245);
nor U8029 (N_8029,N_6287,N_6413);
xnor U8030 (N_8030,N_6653,N_7026);
or U8031 (N_8031,N_6595,N_7155);
xnor U8032 (N_8032,N_7742,N_6710);
or U8033 (N_8033,N_7087,N_7596);
or U8034 (N_8034,N_6907,N_6443);
xnor U8035 (N_8035,N_7556,N_7540);
xnor U8036 (N_8036,N_7455,N_6458);
nand U8037 (N_8037,N_6520,N_6857);
and U8038 (N_8038,N_6552,N_7761);
nand U8039 (N_8039,N_7013,N_6808);
xnor U8040 (N_8040,N_6242,N_6723);
nor U8041 (N_8041,N_7270,N_7722);
or U8042 (N_8042,N_6886,N_6567);
and U8043 (N_8043,N_6227,N_6013);
nand U8044 (N_8044,N_6042,N_7498);
nand U8045 (N_8045,N_6522,N_7263);
nor U8046 (N_8046,N_7928,N_6344);
xor U8047 (N_8047,N_7501,N_6140);
xnor U8048 (N_8048,N_7358,N_6817);
nand U8049 (N_8049,N_6918,N_6705);
nand U8050 (N_8050,N_7019,N_7216);
nor U8051 (N_8051,N_7255,N_6816);
nor U8052 (N_8052,N_7766,N_7543);
nand U8053 (N_8053,N_7756,N_7546);
nor U8054 (N_8054,N_6402,N_7506);
xnor U8055 (N_8055,N_6155,N_6851);
xor U8056 (N_8056,N_7944,N_6164);
nand U8057 (N_8057,N_6684,N_6240);
nor U8058 (N_8058,N_6536,N_6391);
nor U8059 (N_8059,N_6432,N_6184);
xnor U8060 (N_8060,N_6766,N_6990);
nor U8061 (N_8061,N_6267,N_7915);
nor U8062 (N_8062,N_7594,N_7156);
or U8063 (N_8063,N_6069,N_6643);
nand U8064 (N_8064,N_6196,N_6394);
and U8065 (N_8065,N_6950,N_6294);
or U8066 (N_8066,N_7201,N_6778);
xnor U8067 (N_8067,N_6644,N_7044);
nand U8068 (N_8068,N_7696,N_6500);
and U8069 (N_8069,N_6145,N_6987);
nand U8070 (N_8070,N_7059,N_7244);
xor U8071 (N_8071,N_6802,N_7380);
nand U8072 (N_8072,N_6764,N_7593);
xnor U8073 (N_8073,N_7517,N_6779);
or U8074 (N_8074,N_7937,N_7065);
nand U8075 (N_8075,N_6153,N_6998);
nor U8076 (N_8076,N_7012,N_7122);
xor U8077 (N_8077,N_6591,N_7187);
nand U8078 (N_8078,N_6492,N_6895);
or U8079 (N_8079,N_6780,N_7600);
and U8080 (N_8080,N_7646,N_6731);
or U8081 (N_8081,N_6833,N_7298);
and U8082 (N_8082,N_7489,N_6899);
nand U8083 (N_8083,N_6221,N_7412);
and U8084 (N_8084,N_6868,N_7772);
or U8085 (N_8085,N_7120,N_6218);
and U8086 (N_8086,N_7787,N_7254);
xnor U8087 (N_8087,N_6323,N_7822);
xnor U8088 (N_8088,N_6251,N_7676);
xor U8089 (N_8089,N_6133,N_7930);
and U8090 (N_8090,N_7541,N_7148);
or U8091 (N_8091,N_7842,N_6979);
nand U8092 (N_8092,N_6960,N_7170);
or U8093 (N_8093,N_7525,N_7709);
and U8094 (N_8094,N_6200,N_7670);
xor U8095 (N_8095,N_7265,N_6129);
xor U8096 (N_8096,N_6436,N_6733);
nor U8097 (N_8097,N_6231,N_6161);
and U8098 (N_8098,N_6455,N_7018);
nand U8099 (N_8099,N_6144,N_6257);
nand U8100 (N_8100,N_7178,N_6842);
xor U8101 (N_8101,N_6469,N_6573);
or U8102 (N_8102,N_7797,N_7622);
nor U8103 (N_8103,N_6172,N_6272);
or U8104 (N_8104,N_6836,N_7220);
nand U8105 (N_8105,N_6570,N_6178);
or U8106 (N_8106,N_7324,N_7616);
and U8107 (N_8107,N_7620,N_7770);
and U8108 (N_8108,N_6265,N_6532);
and U8109 (N_8109,N_6912,N_6266);
nor U8110 (N_8110,N_6224,N_7981);
nand U8111 (N_8111,N_6847,N_7360);
nand U8112 (N_8112,N_6832,N_7430);
xnor U8113 (N_8113,N_6337,N_6716);
nand U8114 (N_8114,N_7292,N_7399);
nor U8115 (N_8115,N_6073,N_7578);
xor U8116 (N_8116,N_6407,N_6309);
xnor U8117 (N_8117,N_6858,N_7138);
nand U8118 (N_8118,N_6188,N_6415);
nand U8119 (N_8119,N_6098,N_7076);
xor U8120 (N_8120,N_7384,N_7189);
or U8121 (N_8121,N_6750,N_6122);
xnor U8122 (N_8122,N_6429,N_7343);
nor U8123 (N_8123,N_6694,N_6598);
or U8124 (N_8124,N_6856,N_6137);
xnor U8125 (N_8125,N_6491,N_7979);
nand U8126 (N_8126,N_6818,N_6546);
or U8127 (N_8127,N_7703,N_6017);
xor U8128 (N_8128,N_7690,N_7479);
or U8129 (N_8129,N_6647,N_7832);
nor U8130 (N_8130,N_6777,N_7728);
nand U8131 (N_8131,N_6316,N_7748);
nand U8132 (N_8132,N_6550,N_6815);
nor U8133 (N_8133,N_7727,N_6295);
or U8134 (N_8134,N_7046,N_7632);
nand U8135 (N_8135,N_7757,N_7075);
and U8136 (N_8136,N_7544,N_7685);
xnor U8137 (N_8137,N_7512,N_6774);
nand U8138 (N_8138,N_6634,N_6232);
and U8139 (N_8139,N_7840,N_7619);
nand U8140 (N_8140,N_6400,N_7654);
and U8141 (N_8141,N_7705,N_6332);
and U8142 (N_8142,N_7320,N_6428);
and U8143 (N_8143,N_7420,N_7718);
and U8144 (N_8144,N_7785,N_7629);
xnor U8145 (N_8145,N_7768,N_7362);
xnor U8146 (N_8146,N_6088,N_6030);
or U8147 (N_8147,N_6601,N_7901);
and U8148 (N_8148,N_7488,N_6092);
or U8149 (N_8149,N_6989,N_7874);
nor U8150 (N_8150,N_7107,N_7406);
xnor U8151 (N_8151,N_6752,N_6449);
or U8152 (N_8152,N_7001,N_6454);
nand U8153 (N_8153,N_6590,N_6540);
xnor U8154 (N_8154,N_6225,N_6810);
and U8155 (N_8155,N_6057,N_7049);
or U8156 (N_8156,N_7597,N_6826);
xnor U8157 (N_8157,N_7157,N_6538);
and U8158 (N_8158,N_7214,N_7369);
nor U8159 (N_8159,N_7505,N_7653);
nand U8160 (N_8160,N_7197,N_7932);
and U8161 (N_8161,N_7023,N_6748);
xnor U8162 (N_8162,N_6105,N_7762);
nor U8163 (N_8163,N_6525,N_7929);
xnor U8164 (N_8164,N_7831,N_7972);
xnor U8165 (N_8165,N_6049,N_6486);
xor U8166 (N_8166,N_7280,N_7467);
nor U8167 (N_8167,N_6789,N_7310);
nor U8168 (N_8168,N_7459,N_7970);
and U8169 (N_8169,N_7868,N_6163);
nand U8170 (N_8170,N_7266,N_7529);
or U8171 (N_8171,N_6015,N_6473);
nor U8172 (N_8172,N_6479,N_6768);
or U8173 (N_8173,N_7865,N_7213);
nand U8174 (N_8174,N_7834,N_6130);
xor U8175 (N_8175,N_6211,N_6565);
nor U8176 (N_8176,N_6509,N_7977);
or U8177 (N_8177,N_6563,N_6319);
or U8178 (N_8178,N_6001,N_7165);
nor U8179 (N_8179,N_7429,N_6303);
nor U8180 (N_8180,N_6341,N_7448);
nor U8181 (N_8181,N_6116,N_6485);
and U8182 (N_8182,N_7303,N_6234);
nor U8183 (N_8183,N_6951,N_6060);
or U8184 (N_8184,N_6809,N_6219);
nand U8185 (N_8185,N_6311,N_6050);
or U8186 (N_8186,N_6837,N_6439);
and U8187 (N_8187,N_7481,N_7334);
nor U8188 (N_8188,N_7346,N_6146);
nor U8189 (N_8189,N_6587,N_6276);
xnor U8190 (N_8190,N_6425,N_6077);
nand U8191 (N_8191,N_7872,N_6167);
or U8192 (N_8192,N_7108,N_6275);
and U8193 (N_8193,N_6361,N_7763);
nor U8194 (N_8194,N_6884,N_7336);
and U8195 (N_8195,N_7047,N_6493);
nand U8196 (N_8196,N_6788,N_6269);
xor U8197 (N_8197,N_7795,N_6727);
xor U8198 (N_8198,N_6956,N_6403);
nor U8199 (N_8199,N_7090,N_6983);
and U8200 (N_8200,N_6835,N_6593);
or U8201 (N_8201,N_7206,N_7827);
nand U8202 (N_8202,N_6961,N_6529);
and U8203 (N_8203,N_6838,N_6729);
and U8204 (N_8204,N_7079,N_6156);
xnor U8205 (N_8205,N_7402,N_7250);
nor U8206 (N_8206,N_7441,N_6505);
nor U8207 (N_8207,N_6585,N_6084);
nand U8208 (N_8208,N_7248,N_7256);
or U8209 (N_8209,N_7449,N_7192);
nor U8210 (N_8210,N_6735,N_6249);
or U8211 (N_8211,N_7613,N_6574);
nor U8212 (N_8212,N_7724,N_6707);
xor U8213 (N_8213,N_6016,N_6296);
nand U8214 (N_8214,N_7036,N_7628);
xnor U8215 (N_8215,N_7764,N_6503);
nor U8216 (N_8216,N_6474,N_6357);
nand U8217 (N_8217,N_6264,N_7311);
xor U8218 (N_8218,N_7663,N_6758);
xor U8219 (N_8219,N_7988,N_7852);
xor U8220 (N_8220,N_7624,N_7518);
xor U8221 (N_8221,N_7424,N_7810);
nand U8222 (N_8222,N_7144,N_7875);
nor U8223 (N_8223,N_6076,N_6701);
nand U8224 (N_8224,N_7199,N_7866);
nand U8225 (N_8225,N_7224,N_6605);
nor U8226 (N_8226,N_7465,N_7561);
nor U8227 (N_8227,N_7045,N_6321);
or U8228 (N_8228,N_7538,N_6081);
nand U8229 (N_8229,N_7603,N_6358);
nor U8230 (N_8230,N_7683,N_7721);
or U8231 (N_8231,N_7209,N_6741);
nor U8232 (N_8232,N_6176,N_6066);
nor U8233 (N_8233,N_6526,N_7736);
nand U8234 (N_8234,N_6663,N_6352);
and U8235 (N_8235,N_6468,N_7273);
and U8236 (N_8236,N_7438,N_7798);
xnor U8237 (N_8237,N_6139,N_7029);
xor U8238 (N_8238,N_7464,N_7800);
and U8239 (N_8239,N_6630,N_7274);
and U8240 (N_8240,N_7442,N_6160);
and U8241 (N_8241,N_7028,N_7050);
or U8242 (N_8242,N_6058,N_7635);
nor U8243 (N_8243,N_6313,N_7747);
nand U8244 (N_8244,N_7377,N_7180);
and U8245 (N_8245,N_7602,N_6995);
nand U8246 (N_8246,N_7363,N_7809);
xnor U8247 (N_8247,N_6909,N_7316);
xnor U8248 (N_8248,N_6112,N_7470);
nor U8249 (N_8249,N_6359,N_7751);
nand U8250 (N_8250,N_6527,N_7553);
or U8251 (N_8251,N_7953,N_6033);
and U8252 (N_8252,N_7184,N_6256);
or U8253 (N_8253,N_7704,N_7060);
or U8254 (N_8254,N_6602,N_7965);
xnor U8255 (N_8255,N_7813,N_7780);
xor U8256 (N_8256,N_7035,N_6233);
or U8257 (N_8257,N_7514,N_6312);
or U8258 (N_8258,N_6878,N_6064);
and U8259 (N_8259,N_7067,N_7308);
nor U8260 (N_8260,N_6367,N_6271);
or U8261 (N_8261,N_7431,N_7627);
and U8262 (N_8262,N_7235,N_6584);
and U8263 (N_8263,N_6094,N_7519);
xnor U8264 (N_8264,N_7701,N_7281);
or U8265 (N_8265,N_7504,N_7612);
xor U8266 (N_8266,N_6984,N_7963);
and U8267 (N_8267,N_7411,N_6834);
xnor U8268 (N_8268,N_6949,N_7400);
and U8269 (N_8269,N_7951,N_7322);
xnor U8270 (N_8270,N_7111,N_6170);
nand U8271 (N_8271,N_7782,N_6162);
or U8272 (N_8272,N_7608,N_7347);
or U8273 (N_8273,N_7856,N_6955);
and U8274 (N_8274,N_6114,N_7174);
and U8275 (N_8275,N_7008,N_6807);
xor U8276 (N_8276,N_6355,N_7914);
nor U8277 (N_8277,N_7423,N_7847);
and U8278 (N_8278,N_7992,N_7261);
xor U8279 (N_8279,N_7185,N_6263);
nand U8280 (N_8280,N_6915,N_6554);
xor U8281 (N_8281,N_6656,N_6688);
nand U8282 (N_8282,N_6769,N_7557);
and U8283 (N_8283,N_7776,N_7935);
xor U8284 (N_8284,N_6293,N_7241);
xor U8285 (N_8285,N_6457,N_6551);
and U8286 (N_8286,N_7038,N_7434);
and U8287 (N_8287,N_6134,N_7807);
and U8288 (N_8288,N_7127,N_6034);
or U8289 (N_8289,N_6037,N_7016);
nor U8290 (N_8290,N_7176,N_6943);
or U8291 (N_8291,N_7652,N_7159);
nor U8292 (N_8292,N_6152,N_7329);
nand U8293 (N_8293,N_6262,N_7539);
or U8294 (N_8294,N_7665,N_6792);
nand U8295 (N_8295,N_6072,N_6947);
nor U8296 (N_8296,N_7548,N_6327);
and U8297 (N_8297,N_7210,N_6260);
and U8298 (N_8298,N_6787,N_6444);
xor U8299 (N_8299,N_6074,N_7295);
xor U8300 (N_8300,N_6543,N_7689);
and U8301 (N_8301,N_6306,N_6250);
xnor U8302 (N_8302,N_7099,N_7925);
or U8303 (N_8303,N_6518,N_6149);
or U8304 (N_8304,N_6702,N_6869);
or U8305 (N_8305,N_7251,N_7480);
nand U8306 (N_8306,N_6075,N_7618);
or U8307 (N_8307,N_7404,N_7169);
nand U8308 (N_8308,N_6596,N_6434);
nand U8309 (N_8309,N_6118,N_6223);
xor U8310 (N_8310,N_6372,N_6369);
and U8311 (N_8311,N_6461,N_7149);
nand U8312 (N_8312,N_7212,N_7861);
and U8313 (N_8313,N_7054,N_7089);
and U8314 (N_8314,N_6592,N_7843);
nor U8315 (N_8315,N_6870,N_7486);
xnor U8316 (N_8316,N_6089,N_6209);
and U8317 (N_8317,N_7153,N_7503);
nor U8318 (N_8318,N_6667,N_7331);
xor U8319 (N_8319,N_6619,N_7335);
nor U8320 (N_8320,N_7458,N_6314);
nor U8321 (N_8321,N_7607,N_6548);
nand U8322 (N_8322,N_7447,N_6099);
or U8323 (N_8323,N_6119,N_6775);
or U8324 (N_8324,N_6241,N_6477);
nand U8325 (N_8325,N_6708,N_7071);
nor U8326 (N_8326,N_6395,N_7080);
or U8327 (N_8327,N_7996,N_7885);
xor U8328 (N_8328,N_7106,N_7905);
xnor U8329 (N_8329,N_7510,N_6463);
nand U8330 (N_8330,N_6333,N_7877);
nor U8331 (N_8331,N_7614,N_6004);
nor U8332 (N_8332,N_6483,N_7625);
xor U8333 (N_8333,N_7077,N_7168);
xnor U8334 (N_8334,N_6903,N_7511);
or U8335 (N_8335,N_6005,N_7826);
or U8336 (N_8336,N_6627,N_7048);
and U8337 (N_8337,N_6946,N_7710);
nand U8338 (N_8338,N_7788,N_6517);
nor U8339 (N_8339,N_7830,N_7121);
nand U8340 (N_8340,N_7695,N_7582);
xnor U8341 (N_8341,N_6639,N_7383);
nand U8342 (N_8342,N_6572,N_7898);
and U8343 (N_8343,N_7806,N_6419);
nand U8344 (N_8344,N_6141,N_6801);
and U8345 (N_8345,N_7348,N_7355);
and U8346 (N_8346,N_7417,N_7811);
xnor U8347 (N_8347,N_6589,N_6180);
or U8348 (N_8348,N_7037,N_6322);
xor U8349 (N_8349,N_7978,N_7032);
nor U8350 (N_8350,N_7799,N_6438);
xnor U8351 (N_8351,N_6675,N_6524);
xnor U8352 (N_8352,N_6892,N_6481);
and U8353 (N_8353,N_7714,N_6487);
and U8354 (N_8354,N_7774,N_6340);
nor U8355 (N_8355,N_6952,N_6658);
nand U8356 (N_8356,N_6864,N_6380);
nor U8357 (N_8357,N_7203,N_7139);
or U8358 (N_8358,N_7143,N_6922);
nand U8359 (N_8359,N_6091,N_7740);
nand U8360 (N_8360,N_7387,N_6362);
nand U8361 (N_8361,N_7102,N_6508);
nand U8362 (N_8362,N_6097,N_7271);
or U8363 (N_8363,N_7660,N_7982);
nand U8364 (N_8364,N_6096,N_7081);
or U8365 (N_8365,N_6896,N_7516);
or U8366 (N_8366,N_6687,N_6757);
xor U8367 (N_8367,N_7796,N_7252);
and U8368 (N_8368,N_7581,N_7783);
nand U8369 (N_8369,N_7083,N_6677);
nand U8370 (N_8370,N_7668,N_6044);
or U8371 (N_8371,N_7836,N_7960);
or U8372 (N_8372,N_7679,N_7737);
or U8373 (N_8373,N_6499,N_7655);
nor U8374 (N_8374,N_7850,N_6212);
nor U8375 (N_8375,N_6239,N_7222);
and U8376 (N_8376,N_6746,N_7306);
xor U8377 (N_8377,N_7661,N_6165);
and U8378 (N_8378,N_6193,N_6237);
or U8379 (N_8379,N_6978,N_6823);
nor U8380 (N_8380,N_6482,N_6038);
and U8381 (N_8381,N_7995,N_7426);
nand U8382 (N_8382,N_7072,N_6738);
nor U8383 (N_8383,N_6699,N_7994);
nand U8384 (N_8384,N_6274,N_6804);
nor U8385 (N_8385,N_7916,N_6795);
xor U8386 (N_8386,N_7940,N_7911);
xor U8387 (N_8387,N_6288,N_7805);
nor U8388 (N_8388,N_7061,N_7883);
nand U8389 (N_8389,N_6625,N_6925);
xor U8390 (N_8390,N_7171,N_7969);
xnor U8391 (N_8391,N_6537,N_7971);
nand U8392 (N_8392,N_6255,N_7591);
nand U8393 (N_8393,N_7136,N_7894);
or U8394 (N_8394,N_6932,N_7299);
xnor U8395 (N_8395,N_6437,N_7857);
nand U8396 (N_8396,N_6530,N_6539);
and U8397 (N_8397,N_6852,N_7326);
or U8398 (N_8398,N_7116,N_7056);
nand U8399 (N_8399,N_7662,N_7279);
and U8400 (N_8400,N_6618,N_6582);
and U8401 (N_8401,N_7871,N_7422);
or U8402 (N_8402,N_6668,N_6011);
or U8403 (N_8403,N_6514,N_7824);
nor U8404 (N_8404,N_6353,N_7225);
or U8405 (N_8405,N_7386,N_6756);
nand U8406 (N_8406,N_6916,N_6025);
xor U8407 (N_8407,N_6280,N_7900);
nor U8408 (N_8408,N_6652,N_6045);
and U8409 (N_8409,N_6003,N_6125);
or U8410 (N_8410,N_6247,N_6082);
or U8411 (N_8411,N_6945,N_6685);
xnor U8412 (N_8412,N_7317,N_6143);
and U8413 (N_8413,N_7964,N_7078);
and U8414 (N_8414,N_7005,N_7321);
nand U8415 (N_8415,N_7207,N_7651);
nor U8416 (N_8416,N_6666,N_6431);
nor U8417 (N_8417,N_6298,N_7140);
and U8418 (N_8418,N_6475,N_7477);
nand U8419 (N_8419,N_6065,N_6270);
xnor U8420 (N_8420,N_7941,N_7730);
nor U8421 (N_8421,N_7182,N_6975);
xnor U8422 (N_8422,N_7816,N_7440);
and U8423 (N_8423,N_6648,N_7070);
xor U8424 (N_8424,N_7698,N_6174);
xor U8425 (N_8425,N_6336,N_7133);
and U8426 (N_8426,N_7095,N_7907);
or U8427 (N_8427,N_7642,N_6024);
xnor U8428 (N_8428,N_6036,N_6051);
or U8429 (N_8429,N_7712,N_6035);
nand U8430 (N_8430,N_7388,N_6791);
nor U8431 (N_8431,N_7577,N_7200);
nor U8432 (N_8432,N_7571,N_7247);
or U8433 (N_8433,N_7638,N_6459);
and U8434 (N_8434,N_6008,N_6906);
nand U8435 (N_8435,N_6236,N_7946);
nand U8436 (N_8436,N_7876,N_6661);
nand U8437 (N_8437,N_6558,N_7068);
xor U8438 (N_8438,N_6376,N_7333);
xor U8439 (N_8439,N_7733,N_7338);
or U8440 (N_8440,N_7599,N_6334);
or U8441 (N_8441,N_7961,N_7376);
nor U8442 (N_8442,N_6124,N_7862);
nor U8443 (N_8443,N_7484,N_7909);
xnor U8444 (N_8444,N_7015,N_6770);
nor U8445 (N_8445,N_6087,N_7482);
nand U8446 (N_8446,N_7318,N_6566);
nor U8447 (N_8447,N_6282,N_6278);
xor U8448 (N_8448,N_6637,N_6890);
and U8449 (N_8449,N_7967,N_6732);
nor U8450 (N_8450,N_6612,N_6887);
or U8451 (N_8451,N_7419,N_6579);
nor U8452 (N_8452,N_6371,N_7781);
and U8453 (N_8453,N_6564,N_7496);
nor U8454 (N_8454,N_7104,N_6384);
xnor U8455 (N_8455,N_7345,N_7472);
nand U8456 (N_8456,N_6150,N_7957);
xor U8457 (N_8457,N_7461,N_7835);
or U8458 (N_8458,N_7154,N_6451);
xor U8459 (N_8459,N_7490,N_7893);
or U8460 (N_8460,N_6187,N_7566);
or U8461 (N_8461,N_6797,N_7833);
and U8462 (N_8462,N_7713,N_7466);
nor U8463 (N_8463,N_6660,N_6767);
nand U8464 (N_8464,N_6919,N_7439);
and U8465 (N_8465,N_7390,N_7753);
or U8466 (N_8466,N_7064,N_7277);
nor U8467 (N_8467,N_6157,N_7626);
and U8468 (N_8468,N_7110,N_6244);
or U8469 (N_8469,N_6626,N_6190);
nand U8470 (N_8470,N_6202,N_6268);
xnor U8471 (N_8471,N_6997,N_7164);
nor U8472 (N_8472,N_6389,N_6678);
or U8473 (N_8473,N_6938,N_7792);
or U8474 (N_8474,N_6720,N_6325);
or U8475 (N_8475,N_7723,N_6902);
nand U8476 (N_8476,N_6616,N_6910);
xnor U8477 (N_8477,N_6805,N_7687);
xnor U8478 (N_8478,N_7167,N_6308);
xnor U8479 (N_8479,N_7999,N_7196);
xor U8480 (N_8480,N_6029,N_6742);
nand U8481 (N_8481,N_7414,N_7589);
xor U8482 (N_8482,N_6460,N_7902);
xor U8483 (N_8483,N_6388,N_7084);
xnor U8484 (N_8484,N_7873,N_6695);
xnor U8485 (N_8485,N_6205,N_7658);
nand U8486 (N_8486,N_6430,N_7983);
xnor U8487 (N_8487,N_7249,N_6230);
xor U8488 (N_8488,N_7804,N_6893);
and U8489 (N_8489,N_7339,N_6450);
nand U8490 (N_8490,N_7463,N_7294);
or U8491 (N_8491,N_7405,N_6417);
nor U8492 (N_8492,N_6183,N_7112);
xor U8493 (N_8493,N_6095,N_6867);
nand U8494 (N_8494,N_6194,N_7135);
nand U8495 (N_8495,N_7791,N_6026);
and U8496 (N_8496,N_6781,N_6422);
and U8497 (N_8497,N_6628,N_6027);
and U8498 (N_8498,N_7694,N_6923);
nand U8499 (N_8499,N_7137,N_6354);
and U8500 (N_8500,N_6722,N_7846);
or U8501 (N_8501,N_6498,N_7610);
nor U8502 (N_8502,N_7462,N_6970);
or U8503 (N_8503,N_7927,N_6286);
xor U8504 (N_8504,N_6914,N_7499);
and U8505 (N_8505,N_6397,N_6401);
xnor U8506 (N_8506,N_6220,N_6640);
nor U8507 (N_8507,N_7234,N_6819);
nor U8508 (N_8508,N_6261,N_7002);
xnor U8509 (N_8509,N_6674,N_7014);
or U8510 (N_8510,N_6410,N_7814);
nor U8511 (N_8511,N_6138,N_6273);
nor U8512 (N_8512,N_6706,N_6166);
nand U8513 (N_8513,N_6690,N_6228);
or U8514 (N_8514,N_7373,N_6398);
nand U8515 (N_8515,N_7895,N_7731);
and U8516 (N_8516,N_7172,N_6649);
xor U8517 (N_8517,N_6504,N_7073);
or U8518 (N_8518,N_6703,N_6755);
and U8519 (N_8519,N_7606,N_7395);
or U8520 (N_8520,N_7580,N_6488);
xnor U8521 (N_8521,N_6243,N_7948);
nand U8522 (N_8522,N_7604,N_7146);
and U8523 (N_8523,N_7240,N_7243);
and U8524 (N_8524,N_6659,N_7296);
or U8525 (N_8525,N_6046,N_6147);
xor U8526 (N_8526,N_7575,N_7945);
nor U8527 (N_8527,N_6031,N_7558);
xnor U8528 (N_8528,N_7474,N_6448);
or U8529 (N_8529,N_6641,N_6364);
nor U8530 (N_8530,N_6631,N_6542);
or U8531 (N_8531,N_7794,N_6854);
xnor U8532 (N_8532,N_7198,N_7849);
or U8533 (N_8533,N_6506,N_6830);
xnor U8534 (N_8534,N_7681,N_7344);
nor U8535 (N_8535,N_7052,N_7669);
nand U8536 (N_8536,N_7125,N_7202);
xor U8537 (N_8537,N_7547,N_7260);
nand U8538 (N_8538,N_7990,N_7565);
nor U8539 (N_8539,N_6023,N_7283);
and U8540 (N_8540,N_7688,N_7232);
and U8541 (N_8541,N_7542,N_6850);
or U8542 (N_8542,N_7789,N_7743);
and U8543 (N_8543,N_6053,N_6453);
nand U8544 (N_8544,N_6071,N_6424);
nand U8545 (N_8545,N_7601,N_6516);
nor U8546 (N_8546,N_6396,N_7101);
nor U8547 (N_8547,N_7531,N_7314);
nand U8548 (N_8548,N_6339,N_7738);
or U8549 (N_8549,N_6657,N_6418);
nor U8550 (N_8550,N_7410,N_7545);
nor U8551 (N_8551,N_6597,N_6447);
or U8552 (N_8552,N_6820,N_6622);
and U8553 (N_8553,N_7150,N_6588);
and U8554 (N_8554,N_7215,N_6894);
and U8555 (N_8555,N_7803,N_6063);
or U8556 (N_8556,N_6958,N_6055);
xnor U8557 (N_8557,N_7332,N_6101);
nand U8558 (N_8558,N_7991,N_6365);
or U8559 (N_8559,N_6222,N_7350);
nor U8560 (N_8560,N_6603,N_7163);
or U8561 (N_8561,N_7926,N_6967);
nand U8562 (N_8562,N_7643,N_6203);
or U8563 (N_8563,N_7784,N_7986);
nor U8564 (N_8564,N_7903,N_6210);
xor U8565 (N_8565,N_7408,N_7943);
nor U8566 (N_8566,N_6412,N_7204);
nand U8567 (N_8567,N_7889,N_7923);
xnor U8568 (N_8568,N_7487,N_7105);
nor U8569 (N_8569,N_7349,N_7177);
xor U8570 (N_8570,N_7123,N_6994);
nand U8571 (N_8571,N_6600,N_6136);
nand U8572 (N_8572,N_6683,N_6502);
or U8573 (N_8573,N_6317,N_7309);
or U8574 (N_8574,N_7401,N_7523);
xnor U8575 (N_8575,N_6476,N_7631);
nand U8576 (N_8576,N_6191,N_7246);
nand U8577 (N_8577,N_6800,N_7515);
nand U8578 (N_8578,N_6168,N_6700);
or U8579 (N_8579,N_7147,N_7890);
and U8580 (N_8580,N_7371,N_7181);
and U8581 (N_8581,N_6704,N_6040);
and U8582 (N_8582,N_7397,N_6299);
or U8583 (N_8583,N_6414,N_6470);
nor U8584 (N_8584,N_6888,N_6845);
nor U8585 (N_8585,N_7741,N_7912);
nor U8586 (N_8586,N_7374,N_6284);
xnor U8587 (N_8587,N_6093,N_7567);
nor U8588 (N_8588,N_7574,N_7884);
xor U8589 (N_8589,N_7759,N_7492);
nand U8590 (N_8590,N_7573,N_6480);
nor U8591 (N_8591,N_7173,N_7708);
xor U8592 (N_8592,N_7664,N_7648);
xnor U8593 (N_8593,N_6747,N_7230);
nor U8594 (N_8594,N_7183,N_7987);
xnor U8595 (N_8595,N_6872,N_7069);
and U8596 (N_8596,N_6773,N_6734);
nand U8597 (N_8597,N_7495,N_7920);
nand U8598 (N_8598,N_6079,N_7208);
nor U8599 (N_8599,N_6996,N_7673);
and U8600 (N_8600,N_6420,N_7478);
xnor U8601 (N_8601,N_7340,N_7735);
nand U8602 (N_8602,N_6954,N_6957);
xnor U8603 (N_8603,N_6494,N_6304);
or U8604 (N_8604,N_7611,N_6466);
xor U8605 (N_8605,N_6512,N_7236);
or U8606 (N_8606,N_7304,N_6171);
and U8607 (N_8607,N_6335,N_6252);
nor U8608 (N_8608,N_7537,N_6936);
or U8609 (N_8609,N_6966,N_7678);
xor U8610 (N_8610,N_7886,N_7359);
or U8611 (N_8611,N_7218,N_7880);
or U8612 (N_8612,N_6848,N_6427);
and U8613 (N_8613,N_6724,N_7568);
nor U8614 (N_8614,N_6192,N_6028);
and U8615 (N_8615,N_6839,N_7924);
xor U8616 (N_8616,N_6988,N_6599);
nand U8617 (N_8617,N_7456,N_6158);
nor U8618 (N_8618,N_7584,N_7952);
xor U8619 (N_8619,N_7509,N_7973);
or U8620 (N_8620,N_6697,N_6762);
and U8621 (N_8621,N_6464,N_7564);
or U8622 (N_8622,N_6416,N_7726);
nand U8623 (N_8623,N_6324,N_6289);
nor U8624 (N_8624,N_6928,N_7956);
nor U8625 (N_8625,N_6841,N_6490);
xnor U8626 (N_8626,N_7302,N_7837);
or U8627 (N_8627,N_6179,N_7715);
nor U8628 (N_8628,N_6373,N_7022);
and U8629 (N_8629,N_7985,N_6577);
nor U8630 (N_8630,N_6404,N_6014);
and U8631 (N_8631,N_6726,N_7767);
nor U8632 (N_8632,N_6285,N_7285);
xor U8633 (N_8633,N_6173,N_7922);
xor U8634 (N_8634,N_7917,N_7585);
nand U8635 (N_8635,N_6803,N_7253);
nor U8636 (N_8636,N_7838,N_6204);
nor U8637 (N_8637,N_6462,N_7892);
nor U8638 (N_8638,N_6128,N_7086);
xor U8639 (N_8639,N_7382,N_7931);
or U8640 (N_8640,N_7193,N_7904);
nand U8641 (N_8641,N_6226,N_6692);
nor U8642 (N_8642,N_7020,N_6484);
nor U8643 (N_8643,N_6880,N_6739);
and U8644 (N_8644,N_7520,N_7141);
nand U8645 (N_8645,N_7755,N_6513);
nand U8646 (N_8646,N_7968,N_7950);
and U8647 (N_8647,N_6980,N_7719);
nor U8648 (N_8648,N_6553,N_7030);
nand U8649 (N_8649,N_6794,N_7451);
and U8650 (N_8650,N_6070,N_6636);
and U8651 (N_8651,N_7550,N_6531);
nand U8652 (N_8652,N_6195,N_7055);
xor U8653 (N_8653,N_6693,N_6213);
xnor U8654 (N_8654,N_7717,N_6189);
nor U8655 (N_8655,N_6297,N_6972);
nor U8656 (N_8656,N_6510,N_7491);
or U8657 (N_8657,N_7552,N_7711);
and U8658 (N_8658,N_6655,N_6840);
nand U8659 (N_8659,N_6258,N_7375);
and U8660 (N_8660,N_7469,N_7732);
nor U8661 (N_8661,N_7818,N_7330);
and U8662 (N_8662,N_7497,N_7454);
and U8663 (N_8663,N_7063,N_7559);
nor U8664 (N_8664,N_6246,N_6776);
or U8665 (N_8665,N_7290,N_6982);
nor U8666 (N_8666,N_7131,N_7284);
and U8667 (N_8667,N_6712,N_7191);
and U8668 (N_8668,N_7563,N_7186);
nor U8669 (N_8669,N_7353,N_6370);
nand U8670 (N_8670,N_6604,N_7033);
nand U8671 (N_8671,N_7680,N_7808);
nor U8672 (N_8672,N_6467,N_6117);
nand U8673 (N_8673,N_6159,N_6085);
and U8674 (N_8674,N_7088,N_7074);
nor U8675 (N_8675,N_7356,N_7468);
xor U8676 (N_8676,N_6654,N_6366);
and U8677 (N_8677,N_6889,N_6523);
or U8678 (N_8678,N_6993,N_6594);
xor U8679 (N_8679,N_7307,N_7166);
and U8680 (N_8680,N_7769,N_7749);
nor U8681 (N_8681,N_6557,N_7098);
or U8682 (N_8682,N_7117,N_6843);
or U8683 (N_8683,N_6547,N_6151);
or U8684 (N_8684,N_7219,N_7899);
and U8685 (N_8685,N_7119,N_6745);
and U8686 (N_8686,N_7853,N_6719);
nand U8687 (N_8687,N_7342,N_7839);
and U8688 (N_8688,N_7354,N_6920);
nand U8689 (N_8689,N_6127,N_6754);
nand U8690 (N_8690,N_7162,N_6865);
or U8691 (N_8691,N_7569,N_6435);
or U8692 (N_8692,N_7771,N_6559);
and U8693 (N_8693,N_6328,N_7507);
or U8694 (N_8694,N_6786,N_6944);
or U8695 (N_8695,N_7621,N_7421);
nor U8696 (N_8696,N_6214,N_6904);
and U8697 (N_8697,N_7551,N_6866);
nor U8698 (N_8698,N_6534,N_6349);
and U8699 (N_8699,N_7017,N_6609);
nand U8700 (N_8700,N_6964,N_7231);
or U8701 (N_8701,N_6671,N_6763);
nand U8702 (N_8702,N_6495,N_6853);
nor U8703 (N_8703,N_7779,N_6078);
nor U8704 (N_8704,N_7793,N_6933);
nor U8705 (N_8705,N_6154,N_6569);
or U8706 (N_8706,N_6342,N_6446);
xor U8707 (N_8707,N_6381,N_6891);
nand U8708 (N_8708,N_7027,N_6849);
or U8709 (N_8709,N_7416,N_6507);
nand U8710 (N_8710,N_7473,N_6560);
and U8711 (N_8711,N_7450,N_6897);
and U8712 (N_8712,N_7175,N_6528);
nor U8713 (N_8713,N_7684,N_6248);
nor U8714 (N_8714,N_6790,N_7933);
xnor U8715 (N_8715,N_7639,N_7433);
nor U8716 (N_8716,N_6662,N_6544);
xor U8717 (N_8717,N_7124,N_7093);
nor U8718 (N_8718,N_6377,N_7527);
or U8719 (N_8719,N_6650,N_6201);
nand U8720 (N_8720,N_6562,N_6929);
or U8721 (N_8721,N_6059,N_7640);
nor U8722 (N_8722,N_7337,N_6215);
and U8723 (N_8723,N_6318,N_6501);
nand U8724 (N_8724,N_6580,N_6440);
and U8725 (N_8725,N_6277,N_7398);
and U8726 (N_8726,N_7828,N_7586);
xnor U8727 (N_8727,N_6103,N_7259);
and U8728 (N_8728,N_7888,N_6709);
nand U8729 (N_8729,N_7372,N_6669);
or U8730 (N_8730,N_6633,N_6730);
nor U8731 (N_8731,N_6814,N_6375);
nand U8732 (N_8732,N_7691,N_7993);
and U8733 (N_8733,N_6301,N_6113);
or U8734 (N_8734,N_6061,N_7536);
nand U8735 (N_8735,N_6782,N_6632);
nand U8736 (N_8736,N_6969,N_7634);
or U8737 (N_8737,N_6759,N_7003);
xor U8738 (N_8738,N_6292,N_7867);
xor U8739 (N_8739,N_7291,N_6305);
and U8740 (N_8740,N_7094,N_7041);
or U8741 (N_8741,N_7409,N_6822);
or U8742 (N_8742,N_6725,N_6613);
nand U8743 (N_8743,N_7966,N_6921);
nand U8744 (N_8744,N_6924,N_6876);
or U8745 (N_8745,N_7361,N_6208);
nand U8746 (N_8746,N_7351,N_7436);
nand U8747 (N_8747,N_6421,N_6392);
and U8748 (N_8748,N_7858,N_6737);
nand U8749 (N_8749,N_6338,N_7393);
and U8750 (N_8750,N_6829,N_6177);
or U8751 (N_8751,N_6090,N_6310);
xor U8752 (N_8752,N_7671,N_6383);
and U8753 (N_8753,N_7300,N_6885);
or U8754 (N_8754,N_7118,N_7921);
nor U8755 (N_8755,N_6939,N_6861);
and U8756 (N_8756,N_7513,N_6433);
xnor U8757 (N_8757,N_7508,N_6253);
xnor U8758 (N_8758,N_6002,N_6356);
xor U8759 (N_8759,N_6423,N_6608);
nand U8760 (N_8760,N_7534,N_6107);
and U8761 (N_8761,N_6348,N_7211);
nor U8762 (N_8762,N_6541,N_7394);
or U8763 (N_8763,N_7042,N_7297);
nor U8764 (N_8764,N_7583,N_6199);
xor U8765 (N_8765,N_6813,N_6682);
nor U8766 (N_8766,N_6115,N_6022);
nand U8767 (N_8767,N_7605,N_6824);
xor U8768 (N_8768,N_7453,N_6142);
or U8769 (N_8769,N_6390,N_7570);
nand U8770 (N_8770,N_6010,N_7649);
xnor U8771 (N_8771,N_7934,N_7011);
xnor U8772 (N_8772,N_7863,N_7949);
xor U8773 (N_8773,N_6855,N_7007);
or U8774 (N_8774,N_6883,N_7313);
xnor U8775 (N_8775,N_7365,N_6796);
xor U8776 (N_8776,N_6761,N_6465);
and U8777 (N_8777,N_7939,N_6676);
nand U8778 (N_8778,N_6307,N_7962);
or U8779 (N_8779,N_7910,N_7460);
nor U8780 (N_8780,N_7975,N_7976);
nand U8781 (N_8781,N_6426,N_7829);
nor U8782 (N_8782,N_6645,N_6931);
nor U8783 (N_8783,N_7328,N_7392);
xnor U8784 (N_8784,N_7659,N_6175);
xor U8785 (N_8785,N_6583,N_7366);
nor U8786 (N_8786,N_7615,N_6497);
or U8787 (N_8787,N_6545,N_6568);
and U8788 (N_8788,N_7897,N_6811);
nand U8789 (N_8789,N_7657,N_6977);
nand U8790 (N_8790,N_6646,N_7617);
and U8791 (N_8791,N_7752,N_7860);
xor U8792 (N_8792,N_7151,N_7085);
nand U8793 (N_8793,N_6120,N_6571);
nor U8794 (N_8794,N_7364,N_7264);
or U8795 (N_8795,N_6679,N_7609);
nor U8796 (N_8796,N_6360,N_7413);
nor U8797 (N_8797,N_7672,N_7744);
xor U8798 (N_8798,N_7989,N_6406);
and U8799 (N_8799,N_6717,N_6409);
nor U8800 (N_8800,N_6041,N_6111);
nand U8801 (N_8801,N_6689,N_7034);
or U8802 (N_8802,N_6935,N_6986);
and U8803 (N_8803,N_7352,N_7997);
nor U8804 (N_8804,N_7819,N_7775);
or U8805 (N_8805,N_6108,N_6672);
and U8806 (N_8806,N_6575,N_6386);
xor U8807 (N_8807,N_7286,N_7370);
or U8808 (N_8808,N_6680,N_6753);
xor U8809 (N_8809,N_6981,N_6456);
xor U8810 (N_8810,N_6863,N_7327);
nor U8811 (N_8811,N_7521,N_7103);
and U8812 (N_8812,N_6728,N_6515);
and U8813 (N_8813,N_7457,N_7974);
or U8814 (N_8814,N_6721,N_6772);
or U8815 (N_8815,N_7734,N_6623);
or U8816 (N_8816,N_6875,N_6131);
and U8817 (N_8817,N_6744,N_7633);
or U8818 (N_8818,N_7385,N_7720);
nand U8819 (N_8819,N_6080,N_7312);
nand U8820 (N_8820,N_6611,N_6331);
xor U8821 (N_8821,N_7476,N_6452);
nand U8822 (N_8822,N_7555,N_7403);
nand U8823 (N_8823,N_7267,N_6771);
xor U8824 (N_8824,N_7445,N_7301);
xor U8825 (N_8825,N_6039,N_6326);
nand U8826 (N_8826,N_6793,N_7623);
nand U8827 (N_8827,N_7576,N_6006);
nand U8828 (N_8828,N_7287,N_7666);
nor U8829 (N_8829,N_6673,N_6106);
nor U8830 (N_8830,N_7522,N_6104);
and U8831 (N_8831,N_6186,N_7535);
nand U8832 (N_8832,N_7739,N_7786);
nor U8833 (N_8833,N_7257,N_6681);
nor U8834 (N_8834,N_6181,N_6216);
and U8835 (N_8835,N_6974,N_6068);
nand U8836 (N_8836,N_6472,N_6664);
and U8837 (N_8837,N_7595,N_7262);
nor U8838 (N_8838,N_7870,N_7239);
nor U8839 (N_8839,N_6067,N_6638);
xnor U8840 (N_8840,N_7554,N_7217);
or U8841 (N_8841,N_7323,N_6581);
xor U8842 (N_8842,N_6535,N_6126);
or U8843 (N_8843,N_6062,N_7697);
xnor U8844 (N_8844,N_6279,N_6927);
and U8845 (N_8845,N_7844,N_7592);
and U8846 (N_8846,N_6048,N_7238);
nor U8847 (N_8847,N_6020,N_7702);
or U8848 (N_8848,N_6110,N_7378);
xnor U8849 (N_8849,N_7908,N_6290);
or U8850 (N_8850,N_6363,N_6411);
and U8851 (N_8851,N_6021,N_7746);
nand U8852 (N_8852,N_6291,N_6054);
nand U8853 (N_8853,N_6881,N_6940);
or U8854 (N_8854,N_7319,N_6642);
nor U8855 (N_8855,N_6408,N_6715);
nand U8856 (N_8856,N_7500,N_7528);
nor U8857 (N_8857,N_6521,N_6281);
nor U8858 (N_8858,N_7275,N_7161);
nor U8859 (N_8859,N_6478,N_6825);
xnor U8860 (N_8860,N_7237,N_7590);
xor U8861 (N_8861,N_6471,N_6962);
and U8862 (N_8862,N_6877,N_6012);
or U8863 (N_8863,N_6345,N_6941);
and U8864 (N_8864,N_7142,N_7706);
and U8865 (N_8865,N_7674,N_6405);
nor U8866 (N_8866,N_6718,N_6238);
and U8867 (N_8867,N_7998,N_7437);
nor U8868 (N_8868,N_7882,N_6670);
nor U8869 (N_8869,N_7699,N_6686);
nor U8870 (N_8870,N_7641,N_6874);
or U8871 (N_8871,N_7647,N_7896);
nand U8872 (N_8872,N_7205,N_7258);
and U8873 (N_8873,N_7954,N_6330);
nand U8874 (N_8874,N_7725,N_7919);
nand U8875 (N_8875,N_6346,N_6991);
or U8876 (N_8876,N_6217,N_7379);
and U8877 (N_8877,N_7288,N_7452);
xnor U8878 (N_8878,N_6901,N_7980);
and U8879 (N_8879,N_6379,N_7572);
xnor U8880 (N_8880,N_7869,N_7475);
nor U8881 (N_8881,N_7959,N_6930);
xnor U8882 (N_8882,N_7471,N_6828);
nor U8883 (N_8883,N_7878,N_6254);
nor U8884 (N_8884,N_6821,N_7637);
or U8885 (N_8885,N_7765,N_6019);
xor U8886 (N_8886,N_6937,N_7109);
and U8887 (N_8887,N_7160,N_7845);
xnor U8888 (N_8888,N_7010,N_7057);
nand U8889 (N_8889,N_7000,N_7855);
or U8890 (N_8890,N_7686,N_6846);
and U8891 (N_8891,N_7750,N_7821);
or U8892 (N_8892,N_6871,N_6329);
nor U8893 (N_8893,N_7587,N_6760);
or U8894 (N_8894,N_6948,N_7918);
xor U8895 (N_8895,N_7004,N_6812);
nor U8896 (N_8896,N_6913,N_6844);
nand U8897 (N_8897,N_6953,N_6132);
nor U8898 (N_8898,N_6047,N_7113);
xnor U8899 (N_8899,N_7645,N_6713);
xor U8900 (N_8900,N_6610,N_7656);
nor U8901 (N_8901,N_6148,N_6973);
xnor U8902 (N_8902,N_6556,N_6032);
or U8903 (N_8903,N_6882,N_7936);
or U8904 (N_8904,N_7062,N_6320);
or U8905 (N_8905,N_6135,N_7812);
nor U8906 (N_8906,N_7391,N_6965);
or U8907 (N_8907,N_6765,N_7825);
and U8908 (N_8908,N_7278,N_6121);
or U8909 (N_8909,N_6736,N_7693);
and U8910 (N_8910,N_7229,N_7692);
or U8911 (N_8911,N_7848,N_6229);
and U8912 (N_8912,N_6086,N_6533);
xnor U8913 (N_8913,N_6831,N_6123);
and U8914 (N_8914,N_7115,N_7524);
xnor U8915 (N_8915,N_6315,N_6496);
and U8916 (N_8916,N_6100,N_6976);
nor U8917 (N_8917,N_6586,N_7227);
nor U8918 (N_8918,N_7040,N_7667);
or U8919 (N_8919,N_7707,N_7341);
nand U8920 (N_8920,N_7801,N_7879);
xnor U8921 (N_8921,N_7066,N_7289);
nor U8922 (N_8922,N_6198,N_6235);
and U8923 (N_8923,N_7802,N_7425);
nand U8924 (N_8924,N_6615,N_7276);
xor U8925 (N_8925,N_7415,N_7758);
or U8926 (N_8926,N_7682,N_6445);
xor U8927 (N_8927,N_7483,N_6617);
and U8928 (N_8928,N_7228,N_6651);
and U8929 (N_8929,N_6784,N_7129);
nor U8930 (N_8930,N_7043,N_6007);
and U8931 (N_8931,N_7190,N_7096);
or U8932 (N_8932,N_7427,N_7494);
and U8933 (N_8933,N_7636,N_7242);
nor U8934 (N_8934,N_6959,N_6009);
xnor U8935 (N_8935,N_6740,N_7092);
or U8936 (N_8936,N_6859,N_7357);
and U8937 (N_8937,N_7039,N_7233);
and U8938 (N_8938,N_7091,N_6862);
and U8939 (N_8939,N_7562,N_7526);
or U8940 (N_8940,N_7223,N_6343);
nor U8941 (N_8941,N_6621,N_7396);
and U8942 (N_8942,N_7195,N_7817);
or U8943 (N_8943,N_7854,N_6056);
xnor U8944 (N_8944,N_7268,N_6999);
nand U8945 (N_8945,N_7630,N_7859);
nand U8946 (N_8946,N_7790,N_7754);
xnor U8947 (N_8947,N_6185,N_6083);
nor U8948 (N_8948,N_6519,N_6387);
and U8949 (N_8949,N_7443,N_6963);
nor U8950 (N_8950,N_6711,N_6382);
nand U8951 (N_8951,N_6000,N_7282);
and U8952 (N_8952,N_6900,N_6441);
nor U8953 (N_8953,N_7221,N_7864);
or U8954 (N_8954,N_7114,N_7906);
xor U8955 (N_8955,N_7560,N_7145);
or U8956 (N_8956,N_6350,N_6169);
or U8957 (N_8957,N_7226,N_7009);
or U8958 (N_8958,N_6873,N_7428);
nand U8959 (N_8959,N_7823,N_7269);
nor U8960 (N_8960,N_6911,N_6751);
or U8961 (N_8961,N_6374,N_7368);
and U8962 (N_8962,N_7152,N_6378);
or U8963 (N_8963,N_6442,N_7530);
nor U8964 (N_8964,N_6879,N_6052);
nor U8965 (N_8965,N_7305,N_7716);
and U8966 (N_8966,N_6245,N_7913);
nor U8967 (N_8967,N_7820,N_7891);
and U8968 (N_8968,N_7389,N_7493);
nor U8969 (N_8969,N_7025,N_6926);
or U8970 (N_8970,N_7432,N_6785);
and U8971 (N_8971,N_6368,N_6743);
and U8972 (N_8972,N_7024,N_6549);
or U8973 (N_8973,N_7760,N_6917);
xor U8974 (N_8974,N_7533,N_6798);
nand U8975 (N_8975,N_7677,N_6302);
xnor U8976 (N_8976,N_6860,N_7955);
xor U8977 (N_8977,N_7532,N_6578);
nand U8978 (N_8978,N_6905,N_7315);
nor U8979 (N_8979,N_6576,N_6511);
nand U8980 (N_8980,N_7100,N_7130);
xnor U8981 (N_8981,N_6985,N_6393);
and U8982 (N_8982,N_6207,N_6018);
nor U8983 (N_8983,N_7598,N_6399);
and U8984 (N_8984,N_7325,N_7031);
nor U8985 (N_8985,N_6283,N_7132);
xnor U8986 (N_8986,N_7097,N_7367);
nand U8987 (N_8987,N_6934,N_7549);
nand U8988 (N_8988,N_6197,N_7435);
or U8989 (N_8989,N_6898,N_7051);
xor U8990 (N_8990,N_7179,N_6347);
nand U8991 (N_8991,N_6698,N_7188);
or U8992 (N_8992,N_6606,N_6489);
or U8993 (N_8993,N_7947,N_7729);
nor U8994 (N_8994,N_7407,N_7126);
nand U8995 (N_8995,N_6992,N_7128);
nor U8996 (N_8996,N_7058,N_6206);
nor U8997 (N_8997,N_6561,N_6620);
and U8998 (N_8998,N_7444,N_6942);
and U8999 (N_8999,N_6102,N_7938);
xor U9000 (N_9000,N_7670,N_7259);
xor U9001 (N_9001,N_6671,N_7225);
or U9002 (N_9002,N_7387,N_6253);
or U9003 (N_9003,N_6387,N_7523);
nand U9004 (N_9004,N_6350,N_6010);
or U9005 (N_9005,N_7333,N_7768);
and U9006 (N_9006,N_6000,N_6465);
nand U9007 (N_9007,N_6525,N_6982);
xor U9008 (N_9008,N_6622,N_6700);
and U9009 (N_9009,N_7603,N_7649);
nand U9010 (N_9010,N_7207,N_6935);
nor U9011 (N_9011,N_7112,N_6002);
nor U9012 (N_9012,N_6614,N_7221);
xor U9013 (N_9013,N_7358,N_6007);
and U9014 (N_9014,N_7073,N_7487);
and U9015 (N_9015,N_7452,N_6398);
nor U9016 (N_9016,N_6216,N_7523);
nor U9017 (N_9017,N_6546,N_7481);
nand U9018 (N_9018,N_7809,N_6909);
nand U9019 (N_9019,N_6498,N_6735);
nor U9020 (N_9020,N_6284,N_6337);
and U9021 (N_9021,N_6396,N_6787);
or U9022 (N_9022,N_7752,N_7966);
nor U9023 (N_9023,N_7404,N_6270);
or U9024 (N_9024,N_6254,N_7937);
nand U9025 (N_9025,N_7078,N_6370);
and U9026 (N_9026,N_6271,N_7069);
nor U9027 (N_9027,N_7219,N_6945);
nand U9028 (N_9028,N_6152,N_7609);
nand U9029 (N_9029,N_6679,N_6757);
xor U9030 (N_9030,N_6049,N_6870);
xnor U9031 (N_9031,N_7575,N_7310);
or U9032 (N_9032,N_7978,N_6237);
and U9033 (N_9033,N_6511,N_6114);
or U9034 (N_9034,N_6617,N_7128);
nand U9035 (N_9035,N_6859,N_6832);
or U9036 (N_9036,N_7247,N_6847);
or U9037 (N_9037,N_7819,N_7389);
and U9038 (N_9038,N_6388,N_7749);
or U9039 (N_9039,N_7927,N_7111);
nand U9040 (N_9040,N_6926,N_7929);
or U9041 (N_9041,N_6304,N_7329);
nand U9042 (N_9042,N_6211,N_7009);
nand U9043 (N_9043,N_6500,N_7853);
or U9044 (N_9044,N_7548,N_7392);
xor U9045 (N_9045,N_7903,N_6433);
nor U9046 (N_9046,N_7255,N_7473);
xor U9047 (N_9047,N_7215,N_6337);
xnor U9048 (N_9048,N_6009,N_6913);
or U9049 (N_9049,N_6517,N_7667);
or U9050 (N_9050,N_6823,N_7055);
nor U9051 (N_9051,N_7558,N_6849);
nand U9052 (N_9052,N_7459,N_7371);
nand U9053 (N_9053,N_7176,N_7853);
and U9054 (N_9054,N_7519,N_6697);
or U9055 (N_9055,N_6956,N_7222);
xnor U9056 (N_9056,N_7126,N_7755);
nand U9057 (N_9057,N_7358,N_7558);
xor U9058 (N_9058,N_6646,N_7973);
xnor U9059 (N_9059,N_6048,N_7014);
and U9060 (N_9060,N_7625,N_6778);
nor U9061 (N_9061,N_6283,N_7462);
and U9062 (N_9062,N_7303,N_6223);
or U9063 (N_9063,N_6289,N_7080);
or U9064 (N_9064,N_6221,N_6240);
or U9065 (N_9065,N_7891,N_7981);
xnor U9066 (N_9066,N_7961,N_6769);
nor U9067 (N_9067,N_6468,N_6198);
nand U9068 (N_9068,N_7809,N_6277);
nor U9069 (N_9069,N_6246,N_7053);
and U9070 (N_9070,N_6197,N_6685);
nand U9071 (N_9071,N_7918,N_6716);
or U9072 (N_9072,N_7108,N_7864);
nor U9073 (N_9073,N_6026,N_7238);
nor U9074 (N_9074,N_6236,N_7346);
or U9075 (N_9075,N_7954,N_7422);
or U9076 (N_9076,N_7102,N_7841);
or U9077 (N_9077,N_7636,N_6040);
nor U9078 (N_9078,N_7510,N_6875);
xnor U9079 (N_9079,N_7455,N_6133);
nand U9080 (N_9080,N_6352,N_7565);
xnor U9081 (N_9081,N_7448,N_7254);
or U9082 (N_9082,N_7900,N_6685);
nand U9083 (N_9083,N_6189,N_6365);
and U9084 (N_9084,N_6217,N_6004);
or U9085 (N_9085,N_6951,N_6562);
and U9086 (N_9086,N_6694,N_6015);
and U9087 (N_9087,N_6926,N_7665);
nand U9088 (N_9088,N_7541,N_6251);
and U9089 (N_9089,N_6625,N_7096);
and U9090 (N_9090,N_6326,N_6143);
nand U9091 (N_9091,N_6609,N_7407);
and U9092 (N_9092,N_7942,N_7593);
xor U9093 (N_9093,N_6208,N_6127);
nor U9094 (N_9094,N_7682,N_6463);
xnor U9095 (N_9095,N_7400,N_6442);
xor U9096 (N_9096,N_7656,N_7645);
xnor U9097 (N_9097,N_6299,N_6970);
nand U9098 (N_9098,N_7153,N_7336);
and U9099 (N_9099,N_7578,N_7550);
and U9100 (N_9100,N_7372,N_7781);
nor U9101 (N_9101,N_6527,N_7812);
or U9102 (N_9102,N_7892,N_7511);
nand U9103 (N_9103,N_6597,N_7650);
nand U9104 (N_9104,N_6957,N_7937);
or U9105 (N_9105,N_6601,N_7211);
nor U9106 (N_9106,N_6802,N_7408);
or U9107 (N_9107,N_6601,N_6156);
or U9108 (N_9108,N_7186,N_6542);
nand U9109 (N_9109,N_7448,N_7335);
xor U9110 (N_9110,N_7208,N_7910);
nor U9111 (N_9111,N_6911,N_6641);
nor U9112 (N_9112,N_6466,N_6380);
or U9113 (N_9113,N_6069,N_7008);
or U9114 (N_9114,N_6555,N_6200);
or U9115 (N_9115,N_6293,N_7189);
and U9116 (N_9116,N_6143,N_6461);
and U9117 (N_9117,N_7956,N_7767);
nand U9118 (N_9118,N_7713,N_6705);
nand U9119 (N_9119,N_7627,N_6593);
or U9120 (N_9120,N_6114,N_6396);
or U9121 (N_9121,N_6479,N_7139);
nor U9122 (N_9122,N_6560,N_7390);
and U9123 (N_9123,N_6578,N_7573);
or U9124 (N_9124,N_6845,N_6307);
nor U9125 (N_9125,N_6384,N_7304);
nand U9126 (N_9126,N_6697,N_6771);
xnor U9127 (N_9127,N_6662,N_7529);
or U9128 (N_9128,N_7639,N_6124);
nor U9129 (N_9129,N_7860,N_7180);
xor U9130 (N_9130,N_7049,N_6528);
or U9131 (N_9131,N_6484,N_6475);
or U9132 (N_9132,N_6510,N_7101);
and U9133 (N_9133,N_7387,N_6762);
and U9134 (N_9134,N_6928,N_7419);
nand U9135 (N_9135,N_7870,N_7007);
and U9136 (N_9136,N_7196,N_6695);
nand U9137 (N_9137,N_7807,N_7257);
or U9138 (N_9138,N_7834,N_6751);
nand U9139 (N_9139,N_6276,N_6777);
nand U9140 (N_9140,N_6965,N_6992);
nor U9141 (N_9141,N_7865,N_7638);
nor U9142 (N_9142,N_7919,N_7530);
xnor U9143 (N_9143,N_7783,N_6265);
or U9144 (N_9144,N_6273,N_6946);
or U9145 (N_9145,N_6216,N_7765);
or U9146 (N_9146,N_6662,N_7419);
and U9147 (N_9147,N_7128,N_7226);
or U9148 (N_9148,N_7129,N_7030);
or U9149 (N_9149,N_6771,N_6534);
or U9150 (N_9150,N_7073,N_6664);
xnor U9151 (N_9151,N_7412,N_7953);
nand U9152 (N_9152,N_6881,N_6849);
nor U9153 (N_9153,N_7707,N_7646);
xor U9154 (N_9154,N_7952,N_6908);
or U9155 (N_9155,N_7788,N_7391);
nand U9156 (N_9156,N_7718,N_7963);
xor U9157 (N_9157,N_6666,N_6387);
and U9158 (N_9158,N_7214,N_7808);
xor U9159 (N_9159,N_7012,N_6017);
nor U9160 (N_9160,N_7289,N_7365);
or U9161 (N_9161,N_6065,N_7589);
or U9162 (N_9162,N_6803,N_6139);
nor U9163 (N_9163,N_6560,N_6441);
or U9164 (N_9164,N_7769,N_6638);
xnor U9165 (N_9165,N_7670,N_7242);
nand U9166 (N_9166,N_7459,N_6369);
or U9167 (N_9167,N_6107,N_7148);
xor U9168 (N_9168,N_7558,N_7767);
and U9169 (N_9169,N_6919,N_6261);
and U9170 (N_9170,N_6772,N_6518);
or U9171 (N_9171,N_7101,N_6487);
xor U9172 (N_9172,N_6702,N_7989);
nand U9173 (N_9173,N_6923,N_7616);
or U9174 (N_9174,N_7239,N_6568);
xnor U9175 (N_9175,N_6001,N_6154);
and U9176 (N_9176,N_6866,N_7859);
nand U9177 (N_9177,N_7208,N_7754);
or U9178 (N_9178,N_7823,N_6939);
or U9179 (N_9179,N_7323,N_6845);
and U9180 (N_9180,N_6646,N_6989);
nand U9181 (N_9181,N_7724,N_6031);
xor U9182 (N_9182,N_7447,N_7987);
and U9183 (N_9183,N_6352,N_7109);
nor U9184 (N_9184,N_6593,N_6506);
or U9185 (N_9185,N_6009,N_6795);
nor U9186 (N_9186,N_6936,N_7798);
or U9187 (N_9187,N_7949,N_7586);
xor U9188 (N_9188,N_7397,N_7432);
nand U9189 (N_9189,N_7573,N_7130);
and U9190 (N_9190,N_7489,N_7269);
nand U9191 (N_9191,N_7601,N_6222);
and U9192 (N_9192,N_7020,N_7784);
nand U9193 (N_9193,N_7309,N_6368);
nand U9194 (N_9194,N_7883,N_7644);
or U9195 (N_9195,N_7002,N_7217);
nand U9196 (N_9196,N_7813,N_7639);
nand U9197 (N_9197,N_6090,N_7010);
xnor U9198 (N_9198,N_7836,N_7609);
nor U9199 (N_9199,N_6912,N_7507);
xor U9200 (N_9200,N_7294,N_6279);
or U9201 (N_9201,N_7211,N_7671);
xnor U9202 (N_9202,N_7610,N_7227);
nor U9203 (N_9203,N_7223,N_7522);
or U9204 (N_9204,N_6954,N_6014);
nor U9205 (N_9205,N_6789,N_7598);
nor U9206 (N_9206,N_7069,N_6208);
nor U9207 (N_9207,N_6242,N_6810);
xor U9208 (N_9208,N_7695,N_7914);
nor U9209 (N_9209,N_6709,N_6784);
and U9210 (N_9210,N_6641,N_6834);
xor U9211 (N_9211,N_7944,N_6803);
nand U9212 (N_9212,N_6820,N_6318);
or U9213 (N_9213,N_7424,N_6731);
xnor U9214 (N_9214,N_7317,N_6372);
nor U9215 (N_9215,N_6832,N_7799);
or U9216 (N_9216,N_7125,N_7285);
and U9217 (N_9217,N_7243,N_6919);
nand U9218 (N_9218,N_6032,N_7292);
and U9219 (N_9219,N_6593,N_7177);
xor U9220 (N_9220,N_6172,N_6534);
and U9221 (N_9221,N_6554,N_7727);
xor U9222 (N_9222,N_6375,N_7487);
xnor U9223 (N_9223,N_7130,N_7076);
nor U9224 (N_9224,N_7553,N_7885);
or U9225 (N_9225,N_7925,N_6894);
nor U9226 (N_9226,N_7410,N_6589);
or U9227 (N_9227,N_6192,N_7841);
nand U9228 (N_9228,N_7988,N_7685);
and U9229 (N_9229,N_6100,N_6000);
nor U9230 (N_9230,N_7972,N_6925);
nor U9231 (N_9231,N_6924,N_6727);
and U9232 (N_9232,N_7479,N_7226);
or U9233 (N_9233,N_7328,N_6773);
or U9234 (N_9234,N_6652,N_7693);
or U9235 (N_9235,N_6029,N_7291);
and U9236 (N_9236,N_6432,N_6348);
nand U9237 (N_9237,N_6089,N_7247);
nor U9238 (N_9238,N_6307,N_6830);
or U9239 (N_9239,N_7633,N_7332);
nor U9240 (N_9240,N_6715,N_7751);
nor U9241 (N_9241,N_7707,N_7032);
and U9242 (N_9242,N_6116,N_7240);
or U9243 (N_9243,N_7663,N_7099);
xor U9244 (N_9244,N_6249,N_6158);
nand U9245 (N_9245,N_6495,N_6696);
nand U9246 (N_9246,N_7850,N_6234);
nor U9247 (N_9247,N_7793,N_6162);
nand U9248 (N_9248,N_6408,N_7587);
xor U9249 (N_9249,N_6575,N_7208);
xnor U9250 (N_9250,N_6808,N_6036);
and U9251 (N_9251,N_6455,N_6407);
nor U9252 (N_9252,N_7589,N_7961);
xor U9253 (N_9253,N_6746,N_6519);
nor U9254 (N_9254,N_6608,N_7181);
nor U9255 (N_9255,N_6501,N_7491);
xnor U9256 (N_9256,N_6356,N_7834);
and U9257 (N_9257,N_7411,N_6494);
nand U9258 (N_9258,N_6861,N_6000);
nor U9259 (N_9259,N_7065,N_7693);
nor U9260 (N_9260,N_6790,N_6954);
xnor U9261 (N_9261,N_6829,N_7330);
xnor U9262 (N_9262,N_7507,N_6682);
nand U9263 (N_9263,N_7125,N_6694);
or U9264 (N_9264,N_6638,N_6182);
xnor U9265 (N_9265,N_7970,N_6987);
or U9266 (N_9266,N_6396,N_6043);
xnor U9267 (N_9267,N_7941,N_7323);
nand U9268 (N_9268,N_6027,N_7810);
and U9269 (N_9269,N_7753,N_7290);
xor U9270 (N_9270,N_7442,N_6977);
xor U9271 (N_9271,N_7725,N_7534);
and U9272 (N_9272,N_6078,N_7606);
xor U9273 (N_9273,N_6016,N_7036);
or U9274 (N_9274,N_7098,N_7174);
or U9275 (N_9275,N_6075,N_7095);
and U9276 (N_9276,N_7233,N_6241);
nor U9277 (N_9277,N_6071,N_6062);
nor U9278 (N_9278,N_6629,N_6635);
or U9279 (N_9279,N_7720,N_7694);
or U9280 (N_9280,N_6495,N_7059);
nand U9281 (N_9281,N_6258,N_6768);
nand U9282 (N_9282,N_7240,N_7734);
xnor U9283 (N_9283,N_6049,N_7220);
and U9284 (N_9284,N_7304,N_6253);
or U9285 (N_9285,N_7615,N_7007);
nor U9286 (N_9286,N_6012,N_6155);
and U9287 (N_9287,N_6989,N_7939);
nor U9288 (N_9288,N_6908,N_7783);
nor U9289 (N_9289,N_6171,N_6205);
nor U9290 (N_9290,N_7300,N_7123);
nand U9291 (N_9291,N_6081,N_7717);
nand U9292 (N_9292,N_7751,N_7283);
and U9293 (N_9293,N_6478,N_7132);
and U9294 (N_9294,N_7513,N_7889);
or U9295 (N_9295,N_7827,N_6843);
nor U9296 (N_9296,N_7291,N_7367);
xor U9297 (N_9297,N_6362,N_6597);
or U9298 (N_9298,N_7083,N_6213);
or U9299 (N_9299,N_6216,N_6230);
nor U9300 (N_9300,N_6513,N_7680);
nand U9301 (N_9301,N_7100,N_6158);
or U9302 (N_9302,N_7626,N_6143);
or U9303 (N_9303,N_6765,N_6468);
and U9304 (N_9304,N_7306,N_6862);
or U9305 (N_9305,N_7231,N_6101);
xnor U9306 (N_9306,N_6125,N_7371);
and U9307 (N_9307,N_6801,N_7718);
nand U9308 (N_9308,N_6140,N_7672);
nand U9309 (N_9309,N_6948,N_7749);
and U9310 (N_9310,N_7663,N_7723);
xor U9311 (N_9311,N_6161,N_7245);
and U9312 (N_9312,N_7277,N_6066);
and U9313 (N_9313,N_6876,N_7087);
nand U9314 (N_9314,N_7831,N_7277);
and U9315 (N_9315,N_7347,N_7826);
and U9316 (N_9316,N_7760,N_7004);
nor U9317 (N_9317,N_6431,N_7062);
nand U9318 (N_9318,N_6042,N_6571);
and U9319 (N_9319,N_6969,N_7733);
and U9320 (N_9320,N_7822,N_7018);
xor U9321 (N_9321,N_7598,N_6947);
xnor U9322 (N_9322,N_6061,N_6990);
or U9323 (N_9323,N_7359,N_7748);
and U9324 (N_9324,N_7114,N_6738);
nand U9325 (N_9325,N_7424,N_6373);
xor U9326 (N_9326,N_7476,N_7126);
and U9327 (N_9327,N_6117,N_6692);
xnor U9328 (N_9328,N_6789,N_6539);
nand U9329 (N_9329,N_6892,N_6498);
nand U9330 (N_9330,N_6850,N_7101);
nand U9331 (N_9331,N_6456,N_7347);
nand U9332 (N_9332,N_7374,N_7396);
xnor U9333 (N_9333,N_6230,N_7004);
or U9334 (N_9334,N_6822,N_6730);
or U9335 (N_9335,N_7564,N_6552);
and U9336 (N_9336,N_6520,N_6174);
and U9337 (N_9337,N_7636,N_7396);
nor U9338 (N_9338,N_7679,N_6508);
or U9339 (N_9339,N_6959,N_6261);
or U9340 (N_9340,N_7452,N_6924);
xor U9341 (N_9341,N_6081,N_6417);
or U9342 (N_9342,N_7021,N_6261);
xor U9343 (N_9343,N_7321,N_6824);
or U9344 (N_9344,N_6627,N_7249);
and U9345 (N_9345,N_6335,N_6281);
and U9346 (N_9346,N_7929,N_6432);
nor U9347 (N_9347,N_6437,N_7721);
nand U9348 (N_9348,N_7884,N_6658);
nor U9349 (N_9349,N_7607,N_7574);
nand U9350 (N_9350,N_6404,N_7590);
nor U9351 (N_9351,N_6833,N_7459);
nand U9352 (N_9352,N_6447,N_7451);
or U9353 (N_9353,N_6762,N_6745);
nand U9354 (N_9354,N_6631,N_6088);
nand U9355 (N_9355,N_7716,N_7336);
nand U9356 (N_9356,N_7820,N_7918);
and U9357 (N_9357,N_6894,N_7467);
or U9358 (N_9358,N_6693,N_7814);
nand U9359 (N_9359,N_6048,N_7411);
and U9360 (N_9360,N_6288,N_7944);
xor U9361 (N_9361,N_7624,N_6665);
xor U9362 (N_9362,N_7747,N_7343);
nor U9363 (N_9363,N_6453,N_6090);
nand U9364 (N_9364,N_6957,N_7204);
and U9365 (N_9365,N_6589,N_6779);
xor U9366 (N_9366,N_6229,N_6843);
or U9367 (N_9367,N_6794,N_7108);
and U9368 (N_9368,N_6591,N_6467);
xor U9369 (N_9369,N_6672,N_6895);
nor U9370 (N_9370,N_7867,N_7789);
or U9371 (N_9371,N_7238,N_7672);
or U9372 (N_9372,N_6541,N_6377);
nor U9373 (N_9373,N_6285,N_6701);
xor U9374 (N_9374,N_7803,N_7866);
or U9375 (N_9375,N_6873,N_6260);
nand U9376 (N_9376,N_6054,N_7671);
nor U9377 (N_9377,N_7596,N_7412);
xor U9378 (N_9378,N_6465,N_6498);
nor U9379 (N_9379,N_7128,N_7270);
nor U9380 (N_9380,N_7012,N_6823);
and U9381 (N_9381,N_6466,N_7692);
nor U9382 (N_9382,N_7178,N_7901);
xnor U9383 (N_9383,N_6370,N_7677);
and U9384 (N_9384,N_7989,N_7255);
nand U9385 (N_9385,N_7683,N_6216);
nor U9386 (N_9386,N_7052,N_6685);
nand U9387 (N_9387,N_7209,N_7661);
xnor U9388 (N_9388,N_6079,N_6563);
and U9389 (N_9389,N_6680,N_7545);
nor U9390 (N_9390,N_7046,N_7695);
or U9391 (N_9391,N_7050,N_7371);
xor U9392 (N_9392,N_6593,N_7360);
or U9393 (N_9393,N_6881,N_7755);
xnor U9394 (N_9394,N_7728,N_6934);
nand U9395 (N_9395,N_6263,N_6767);
and U9396 (N_9396,N_7625,N_7936);
nor U9397 (N_9397,N_7563,N_6485);
nand U9398 (N_9398,N_7580,N_7025);
nand U9399 (N_9399,N_6173,N_7470);
nor U9400 (N_9400,N_6553,N_6404);
nor U9401 (N_9401,N_6384,N_6618);
xnor U9402 (N_9402,N_6458,N_6626);
nor U9403 (N_9403,N_6268,N_7573);
or U9404 (N_9404,N_6230,N_6592);
nor U9405 (N_9405,N_7157,N_7086);
and U9406 (N_9406,N_6600,N_6846);
nor U9407 (N_9407,N_6957,N_7855);
nand U9408 (N_9408,N_6794,N_7854);
xor U9409 (N_9409,N_6355,N_6076);
nor U9410 (N_9410,N_6482,N_6192);
and U9411 (N_9411,N_7009,N_6771);
nor U9412 (N_9412,N_7639,N_7143);
nor U9413 (N_9413,N_6083,N_7990);
and U9414 (N_9414,N_6046,N_7997);
nand U9415 (N_9415,N_6175,N_7730);
and U9416 (N_9416,N_7295,N_6085);
nor U9417 (N_9417,N_7439,N_6012);
or U9418 (N_9418,N_7365,N_7489);
nand U9419 (N_9419,N_6245,N_7367);
nor U9420 (N_9420,N_7958,N_6634);
and U9421 (N_9421,N_7958,N_7754);
xnor U9422 (N_9422,N_7311,N_7387);
nand U9423 (N_9423,N_7224,N_6167);
nand U9424 (N_9424,N_6844,N_6753);
nand U9425 (N_9425,N_6369,N_7693);
and U9426 (N_9426,N_6819,N_7985);
nor U9427 (N_9427,N_7422,N_6480);
nor U9428 (N_9428,N_6537,N_7913);
or U9429 (N_9429,N_7368,N_6478);
xor U9430 (N_9430,N_6564,N_6405);
or U9431 (N_9431,N_7598,N_6410);
and U9432 (N_9432,N_6938,N_6617);
and U9433 (N_9433,N_7100,N_7065);
or U9434 (N_9434,N_6952,N_6248);
nor U9435 (N_9435,N_7417,N_7413);
nand U9436 (N_9436,N_7299,N_6317);
xor U9437 (N_9437,N_7260,N_7574);
nand U9438 (N_9438,N_6371,N_7102);
nor U9439 (N_9439,N_6670,N_7370);
and U9440 (N_9440,N_7407,N_6427);
and U9441 (N_9441,N_7455,N_7623);
xor U9442 (N_9442,N_7159,N_7207);
or U9443 (N_9443,N_7727,N_7842);
xnor U9444 (N_9444,N_7963,N_7444);
and U9445 (N_9445,N_7043,N_7164);
nand U9446 (N_9446,N_6156,N_6298);
nand U9447 (N_9447,N_6268,N_6925);
and U9448 (N_9448,N_7216,N_6399);
nor U9449 (N_9449,N_6737,N_6496);
or U9450 (N_9450,N_7221,N_6205);
and U9451 (N_9451,N_6356,N_6771);
and U9452 (N_9452,N_7181,N_7578);
and U9453 (N_9453,N_7403,N_7591);
or U9454 (N_9454,N_7410,N_6927);
nor U9455 (N_9455,N_6348,N_6296);
nand U9456 (N_9456,N_6962,N_7104);
and U9457 (N_9457,N_6943,N_6873);
or U9458 (N_9458,N_7255,N_7798);
or U9459 (N_9459,N_6160,N_7577);
or U9460 (N_9460,N_6804,N_6400);
and U9461 (N_9461,N_6114,N_7775);
xor U9462 (N_9462,N_7233,N_6152);
nand U9463 (N_9463,N_7967,N_7115);
xor U9464 (N_9464,N_7304,N_7558);
xor U9465 (N_9465,N_7976,N_6402);
xnor U9466 (N_9466,N_7281,N_7140);
xor U9467 (N_9467,N_7971,N_6056);
nand U9468 (N_9468,N_7053,N_6358);
and U9469 (N_9469,N_7042,N_7352);
and U9470 (N_9470,N_7890,N_6145);
or U9471 (N_9471,N_6981,N_6466);
and U9472 (N_9472,N_6378,N_7027);
or U9473 (N_9473,N_6533,N_7087);
nand U9474 (N_9474,N_6499,N_6066);
nand U9475 (N_9475,N_6416,N_7414);
nand U9476 (N_9476,N_6089,N_7917);
nand U9477 (N_9477,N_7390,N_7917);
or U9478 (N_9478,N_6752,N_7826);
and U9479 (N_9479,N_6106,N_7896);
nand U9480 (N_9480,N_6262,N_7481);
or U9481 (N_9481,N_6021,N_6420);
nor U9482 (N_9482,N_7471,N_7942);
nand U9483 (N_9483,N_7905,N_6008);
nand U9484 (N_9484,N_6952,N_6068);
xor U9485 (N_9485,N_7153,N_7144);
nor U9486 (N_9486,N_7330,N_7814);
xnor U9487 (N_9487,N_7468,N_7443);
nor U9488 (N_9488,N_7309,N_7927);
and U9489 (N_9489,N_6676,N_7699);
nand U9490 (N_9490,N_7381,N_7201);
nor U9491 (N_9491,N_7586,N_6365);
nand U9492 (N_9492,N_7296,N_6786);
nand U9493 (N_9493,N_7589,N_7467);
nand U9494 (N_9494,N_6954,N_6214);
nand U9495 (N_9495,N_7013,N_7394);
xnor U9496 (N_9496,N_6028,N_6298);
or U9497 (N_9497,N_7970,N_6312);
nor U9498 (N_9498,N_6617,N_7526);
and U9499 (N_9499,N_7408,N_7125);
nor U9500 (N_9500,N_6078,N_7021);
nor U9501 (N_9501,N_6276,N_7350);
and U9502 (N_9502,N_7574,N_6905);
and U9503 (N_9503,N_7078,N_7988);
nand U9504 (N_9504,N_6692,N_6671);
nor U9505 (N_9505,N_7409,N_6377);
and U9506 (N_9506,N_7404,N_7005);
nand U9507 (N_9507,N_6281,N_6313);
and U9508 (N_9508,N_7840,N_7293);
or U9509 (N_9509,N_6513,N_7310);
nor U9510 (N_9510,N_6745,N_6424);
and U9511 (N_9511,N_7582,N_6440);
xor U9512 (N_9512,N_6766,N_7746);
or U9513 (N_9513,N_7097,N_7483);
nor U9514 (N_9514,N_6186,N_7041);
and U9515 (N_9515,N_6655,N_7972);
or U9516 (N_9516,N_7093,N_7380);
nand U9517 (N_9517,N_6974,N_6397);
nor U9518 (N_9518,N_6848,N_7650);
or U9519 (N_9519,N_6005,N_6407);
xnor U9520 (N_9520,N_6802,N_7192);
xnor U9521 (N_9521,N_7969,N_6419);
or U9522 (N_9522,N_7445,N_7593);
xor U9523 (N_9523,N_7424,N_7568);
xnor U9524 (N_9524,N_7636,N_6269);
xor U9525 (N_9525,N_6564,N_6987);
nand U9526 (N_9526,N_6350,N_6422);
nor U9527 (N_9527,N_6001,N_7695);
nand U9528 (N_9528,N_6909,N_7384);
and U9529 (N_9529,N_6183,N_6096);
and U9530 (N_9530,N_7873,N_7979);
nand U9531 (N_9531,N_6547,N_7525);
and U9532 (N_9532,N_7975,N_6486);
or U9533 (N_9533,N_6918,N_7398);
xnor U9534 (N_9534,N_7381,N_6839);
xor U9535 (N_9535,N_6328,N_7869);
xnor U9536 (N_9536,N_7259,N_7830);
and U9537 (N_9537,N_7242,N_6588);
nor U9538 (N_9538,N_7399,N_6840);
and U9539 (N_9539,N_6474,N_7807);
nand U9540 (N_9540,N_7840,N_7429);
xor U9541 (N_9541,N_7296,N_7202);
nor U9542 (N_9542,N_7106,N_6142);
xor U9543 (N_9543,N_6738,N_6019);
and U9544 (N_9544,N_6706,N_6471);
or U9545 (N_9545,N_7595,N_6096);
or U9546 (N_9546,N_6552,N_6049);
or U9547 (N_9547,N_6530,N_6445);
xor U9548 (N_9548,N_7903,N_6462);
nand U9549 (N_9549,N_7330,N_6082);
nor U9550 (N_9550,N_6106,N_7606);
or U9551 (N_9551,N_7211,N_7122);
and U9552 (N_9552,N_7406,N_7664);
nor U9553 (N_9553,N_7607,N_7603);
and U9554 (N_9554,N_6122,N_7765);
and U9555 (N_9555,N_6711,N_7317);
or U9556 (N_9556,N_7093,N_7426);
or U9557 (N_9557,N_7207,N_7768);
or U9558 (N_9558,N_7966,N_6987);
xor U9559 (N_9559,N_6528,N_6511);
xor U9560 (N_9560,N_6219,N_7425);
nor U9561 (N_9561,N_7736,N_7835);
nand U9562 (N_9562,N_7390,N_6591);
nor U9563 (N_9563,N_6821,N_6740);
nor U9564 (N_9564,N_7295,N_7384);
nand U9565 (N_9565,N_6470,N_7725);
and U9566 (N_9566,N_7245,N_6252);
nand U9567 (N_9567,N_6589,N_7628);
nor U9568 (N_9568,N_7963,N_6115);
nor U9569 (N_9569,N_6976,N_6978);
or U9570 (N_9570,N_7063,N_6934);
nand U9571 (N_9571,N_7460,N_7878);
nand U9572 (N_9572,N_6701,N_7016);
and U9573 (N_9573,N_7239,N_6328);
nand U9574 (N_9574,N_6914,N_7008);
and U9575 (N_9575,N_6921,N_6356);
or U9576 (N_9576,N_7834,N_6429);
xor U9577 (N_9577,N_6338,N_6472);
nor U9578 (N_9578,N_7040,N_6793);
and U9579 (N_9579,N_6934,N_6802);
nand U9580 (N_9580,N_7352,N_7538);
nand U9581 (N_9581,N_6375,N_7861);
nand U9582 (N_9582,N_6917,N_7530);
nand U9583 (N_9583,N_7191,N_6955);
or U9584 (N_9584,N_7938,N_7591);
and U9585 (N_9585,N_7832,N_7596);
xnor U9586 (N_9586,N_7623,N_6286);
and U9587 (N_9587,N_6587,N_7080);
nor U9588 (N_9588,N_7663,N_6570);
and U9589 (N_9589,N_6412,N_7580);
nor U9590 (N_9590,N_7977,N_7032);
or U9591 (N_9591,N_6872,N_7410);
or U9592 (N_9592,N_6255,N_7140);
nand U9593 (N_9593,N_6521,N_6458);
nand U9594 (N_9594,N_6951,N_6322);
and U9595 (N_9595,N_6307,N_6821);
xor U9596 (N_9596,N_7549,N_6819);
or U9597 (N_9597,N_7975,N_7585);
nor U9598 (N_9598,N_6339,N_6511);
and U9599 (N_9599,N_7705,N_7824);
xor U9600 (N_9600,N_7179,N_7155);
or U9601 (N_9601,N_7475,N_7053);
nor U9602 (N_9602,N_6860,N_6119);
nand U9603 (N_9603,N_7469,N_6007);
and U9604 (N_9604,N_7781,N_6384);
nor U9605 (N_9605,N_7211,N_7975);
and U9606 (N_9606,N_6570,N_6256);
nor U9607 (N_9607,N_7472,N_7262);
nand U9608 (N_9608,N_6360,N_7060);
and U9609 (N_9609,N_7436,N_6223);
or U9610 (N_9610,N_6176,N_6078);
or U9611 (N_9611,N_7604,N_6416);
xnor U9612 (N_9612,N_7397,N_7971);
xnor U9613 (N_9613,N_7867,N_7148);
nor U9614 (N_9614,N_6084,N_6884);
xor U9615 (N_9615,N_7472,N_6432);
nand U9616 (N_9616,N_6594,N_6321);
nand U9617 (N_9617,N_6108,N_6914);
nand U9618 (N_9618,N_7911,N_6117);
and U9619 (N_9619,N_6163,N_6965);
xor U9620 (N_9620,N_6027,N_6138);
nor U9621 (N_9621,N_6595,N_7128);
nand U9622 (N_9622,N_6687,N_6064);
xor U9623 (N_9623,N_6952,N_6445);
nor U9624 (N_9624,N_7620,N_6816);
or U9625 (N_9625,N_7989,N_6810);
xor U9626 (N_9626,N_6471,N_7959);
and U9627 (N_9627,N_7130,N_7796);
xnor U9628 (N_9628,N_6773,N_7414);
or U9629 (N_9629,N_7791,N_6419);
nor U9630 (N_9630,N_7466,N_6197);
or U9631 (N_9631,N_6967,N_7907);
nand U9632 (N_9632,N_7426,N_6865);
nand U9633 (N_9633,N_7411,N_7231);
or U9634 (N_9634,N_6669,N_7794);
or U9635 (N_9635,N_6274,N_6339);
and U9636 (N_9636,N_6149,N_7240);
xnor U9637 (N_9637,N_6616,N_6782);
nand U9638 (N_9638,N_7030,N_6801);
nor U9639 (N_9639,N_6900,N_7252);
or U9640 (N_9640,N_6968,N_6499);
nand U9641 (N_9641,N_6917,N_6556);
and U9642 (N_9642,N_6645,N_6427);
xnor U9643 (N_9643,N_7078,N_7469);
nor U9644 (N_9644,N_7839,N_6557);
or U9645 (N_9645,N_6016,N_6840);
nand U9646 (N_9646,N_7992,N_7262);
or U9647 (N_9647,N_6994,N_7080);
or U9648 (N_9648,N_7029,N_6890);
or U9649 (N_9649,N_7166,N_6481);
and U9650 (N_9650,N_7427,N_7109);
nor U9651 (N_9651,N_6193,N_6199);
xor U9652 (N_9652,N_6998,N_7576);
xor U9653 (N_9653,N_6060,N_6467);
nand U9654 (N_9654,N_7967,N_6419);
or U9655 (N_9655,N_6721,N_7351);
xnor U9656 (N_9656,N_6398,N_6194);
xnor U9657 (N_9657,N_7487,N_6311);
xnor U9658 (N_9658,N_7648,N_7971);
nor U9659 (N_9659,N_6522,N_7305);
xor U9660 (N_9660,N_7767,N_6628);
nand U9661 (N_9661,N_7817,N_7997);
nand U9662 (N_9662,N_7751,N_6205);
and U9663 (N_9663,N_6886,N_6591);
or U9664 (N_9664,N_6475,N_7563);
nor U9665 (N_9665,N_6063,N_6718);
or U9666 (N_9666,N_7394,N_6651);
xnor U9667 (N_9667,N_6880,N_7872);
xor U9668 (N_9668,N_7608,N_6271);
nand U9669 (N_9669,N_7008,N_7958);
nor U9670 (N_9670,N_7995,N_6097);
nand U9671 (N_9671,N_6593,N_6641);
nor U9672 (N_9672,N_6679,N_6660);
nand U9673 (N_9673,N_7973,N_7944);
or U9674 (N_9674,N_6439,N_7147);
and U9675 (N_9675,N_6722,N_7813);
nand U9676 (N_9676,N_6306,N_7311);
and U9677 (N_9677,N_7009,N_7396);
or U9678 (N_9678,N_6133,N_7704);
or U9679 (N_9679,N_6207,N_6550);
nor U9680 (N_9680,N_6804,N_7209);
xnor U9681 (N_9681,N_6747,N_7131);
nand U9682 (N_9682,N_6703,N_7387);
or U9683 (N_9683,N_7306,N_7491);
nand U9684 (N_9684,N_7767,N_6536);
xor U9685 (N_9685,N_6709,N_7137);
xor U9686 (N_9686,N_6940,N_7566);
or U9687 (N_9687,N_6397,N_6205);
xor U9688 (N_9688,N_7990,N_6748);
or U9689 (N_9689,N_6457,N_6365);
nand U9690 (N_9690,N_7343,N_7281);
and U9691 (N_9691,N_6144,N_7413);
nor U9692 (N_9692,N_6040,N_7579);
xor U9693 (N_9693,N_6460,N_6612);
or U9694 (N_9694,N_7172,N_7025);
or U9695 (N_9695,N_7161,N_7811);
nand U9696 (N_9696,N_7220,N_6192);
and U9697 (N_9697,N_6614,N_7835);
xor U9698 (N_9698,N_6690,N_7046);
nor U9699 (N_9699,N_6669,N_7346);
xnor U9700 (N_9700,N_6148,N_6428);
xor U9701 (N_9701,N_6370,N_6838);
nor U9702 (N_9702,N_6152,N_7846);
or U9703 (N_9703,N_6560,N_6740);
nor U9704 (N_9704,N_7210,N_6453);
nor U9705 (N_9705,N_6168,N_6418);
nand U9706 (N_9706,N_6814,N_6350);
and U9707 (N_9707,N_6288,N_7597);
xor U9708 (N_9708,N_6980,N_6333);
or U9709 (N_9709,N_7938,N_6998);
nand U9710 (N_9710,N_6136,N_7667);
and U9711 (N_9711,N_6530,N_7940);
xor U9712 (N_9712,N_6541,N_6291);
nand U9713 (N_9713,N_6783,N_7949);
or U9714 (N_9714,N_6834,N_6178);
nand U9715 (N_9715,N_6862,N_6363);
xor U9716 (N_9716,N_6521,N_6202);
or U9717 (N_9717,N_7760,N_6803);
nor U9718 (N_9718,N_7605,N_7796);
or U9719 (N_9719,N_6801,N_7407);
or U9720 (N_9720,N_7118,N_7160);
xnor U9721 (N_9721,N_7001,N_6662);
and U9722 (N_9722,N_6841,N_7948);
nor U9723 (N_9723,N_6307,N_6083);
xor U9724 (N_9724,N_6812,N_6446);
xor U9725 (N_9725,N_6314,N_7024);
or U9726 (N_9726,N_7220,N_6313);
nor U9727 (N_9727,N_6178,N_6612);
xor U9728 (N_9728,N_7265,N_7503);
or U9729 (N_9729,N_7367,N_6393);
nand U9730 (N_9730,N_7012,N_6361);
xnor U9731 (N_9731,N_7335,N_7034);
nand U9732 (N_9732,N_7060,N_7502);
nand U9733 (N_9733,N_7501,N_6656);
xor U9734 (N_9734,N_6465,N_6500);
and U9735 (N_9735,N_6709,N_7724);
or U9736 (N_9736,N_6762,N_7498);
and U9737 (N_9737,N_6922,N_7586);
nor U9738 (N_9738,N_6377,N_7107);
nand U9739 (N_9739,N_7013,N_6987);
or U9740 (N_9740,N_6510,N_6830);
nor U9741 (N_9741,N_7465,N_7025);
or U9742 (N_9742,N_6005,N_6309);
xnor U9743 (N_9743,N_7391,N_7876);
xnor U9744 (N_9744,N_6170,N_7883);
or U9745 (N_9745,N_6668,N_6107);
and U9746 (N_9746,N_6487,N_6402);
or U9747 (N_9747,N_7558,N_6264);
nor U9748 (N_9748,N_6266,N_6023);
nor U9749 (N_9749,N_7214,N_6259);
nand U9750 (N_9750,N_7520,N_6414);
and U9751 (N_9751,N_7425,N_7047);
or U9752 (N_9752,N_7618,N_6733);
or U9753 (N_9753,N_6408,N_7019);
xor U9754 (N_9754,N_6742,N_6915);
and U9755 (N_9755,N_7609,N_7995);
nand U9756 (N_9756,N_7893,N_7513);
nand U9757 (N_9757,N_7819,N_6634);
xnor U9758 (N_9758,N_6749,N_6408);
and U9759 (N_9759,N_7038,N_7585);
or U9760 (N_9760,N_6299,N_7196);
nand U9761 (N_9761,N_6241,N_7599);
xnor U9762 (N_9762,N_6238,N_6427);
nor U9763 (N_9763,N_7232,N_6453);
nor U9764 (N_9764,N_7978,N_7856);
and U9765 (N_9765,N_6196,N_6873);
nand U9766 (N_9766,N_7586,N_7182);
nand U9767 (N_9767,N_6029,N_7630);
nor U9768 (N_9768,N_6096,N_7627);
xnor U9769 (N_9769,N_6258,N_7876);
or U9770 (N_9770,N_6299,N_7655);
or U9771 (N_9771,N_7888,N_6734);
nor U9772 (N_9772,N_6122,N_7960);
and U9773 (N_9773,N_6487,N_7299);
or U9774 (N_9774,N_7829,N_7139);
and U9775 (N_9775,N_7464,N_7778);
or U9776 (N_9776,N_7011,N_6473);
nand U9777 (N_9777,N_7159,N_7161);
nor U9778 (N_9778,N_7700,N_6985);
xnor U9779 (N_9779,N_7919,N_6624);
and U9780 (N_9780,N_6510,N_6072);
or U9781 (N_9781,N_6229,N_7234);
nand U9782 (N_9782,N_7939,N_7582);
nor U9783 (N_9783,N_6883,N_7161);
xor U9784 (N_9784,N_6132,N_6006);
and U9785 (N_9785,N_6563,N_6859);
nor U9786 (N_9786,N_6684,N_6872);
xor U9787 (N_9787,N_6181,N_7549);
or U9788 (N_9788,N_7672,N_7221);
xor U9789 (N_9789,N_7120,N_7230);
nand U9790 (N_9790,N_7604,N_7590);
and U9791 (N_9791,N_7647,N_7183);
nor U9792 (N_9792,N_7426,N_7699);
nor U9793 (N_9793,N_7012,N_6714);
or U9794 (N_9794,N_6770,N_6630);
nor U9795 (N_9795,N_7236,N_6832);
and U9796 (N_9796,N_6144,N_6649);
xnor U9797 (N_9797,N_6056,N_6720);
or U9798 (N_9798,N_7242,N_7266);
and U9799 (N_9799,N_6262,N_6325);
nand U9800 (N_9800,N_7520,N_7506);
nand U9801 (N_9801,N_6450,N_6233);
and U9802 (N_9802,N_7210,N_6072);
nor U9803 (N_9803,N_7658,N_6536);
xor U9804 (N_9804,N_6875,N_6101);
nand U9805 (N_9805,N_7427,N_6861);
nor U9806 (N_9806,N_6523,N_6794);
or U9807 (N_9807,N_6648,N_7202);
nand U9808 (N_9808,N_6765,N_7306);
or U9809 (N_9809,N_6082,N_6737);
nor U9810 (N_9810,N_6891,N_6216);
nor U9811 (N_9811,N_7380,N_7081);
or U9812 (N_9812,N_6405,N_7369);
and U9813 (N_9813,N_6298,N_6727);
or U9814 (N_9814,N_7029,N_6207);
or U9815 (N_9815,N_6284,N_7171);
and U9816 (N_9816,N_7046,N_7762);
nor U9817 (N_9817,N_7836,N_6867);
xor U9818 (N_9818,N_6164,N_6918);
nand U9819 (N_9819,N_6932,N_7094);
nor U9820 (N_9820,N_7786,N_6398);
xor U9821 (N_9821,N_7857,N_6585);
nor U9822 (N_9822,N_6111,N_6820);
and U9823 (N_9823,N_7008,N_6330);
and U9824 (N_9824,N_7842,N_7529);
xnor U9825 (N_9825,N_6997,N_6355);
nor U9826 (N_9826,N_6551,N_6208);
and U9827 (N_9827,N_7894,N_7530);
xor U9828 (N_9828,N_6909,N_6772);
or U9829 (N_9829,N_6299,N_6942);
nand U9830 (N_9830,N_6075,N_6797);
nand U9831 (N_9831,N_7585,N_7709);
and U9832 (N_9832,N_7011,N_7955);
and U9833 (N_9833,N_7312,N_7176);
nand U9834 (N_9834,N_7915,N_7447);
nor U9835 (N_9835,N_6836,N_6011);
and U9836 (N_9836,N_7068,N_6841);
or U9837 (N_9837,N_6230,N_7303);
and U9838 (N_9838,N_7638,N_6252);
and U9839 (N_9839,N_6123,N_7653);
or U9840 (N_9840,N_7312,N_7505);
and U9841 (N_9841,N_7204,N_7905);
and U9842 (N_9842,N_6132,N_6634);
and U9843 (N_9843,N_7177,N_6789);
nor U9844 (N_9844,N_7910,N_6486);
xor U9845 (N_9845,N_6469,N_6282);
xor U9846 (N_9846,N_6330,N_7075);
xnor U9847 (N_9847,N_7261,N_7380);
and U9848 (N_9848,N_7452,N_6059);
and U9849 (N_9849,N_7579,N_7954);
xnor U9850 (N_9850,N_7017,N_7014);
and U9851 (N_9851,N_7917,N_6423);
and U9852 (N_9852,N_7789,N_6585);
or U9853 (N_9853,N_6434,N_6167);
nor U9854 (N_9854,N_6006,N_7651);
or U9855 (N_9855,N_7007,N_6741);
nand U9856 (N_9856,N_6393,N_7184);
xnor U9857 (N_9857,N_6837,N_7700);
nor U9858 (N_9858,N_6279,N_6317);
nand U9859 (N_9859,N_7430,N_6728);
and U9860 (N_9860,N_6904,N_7756);
xnor U9861 (N_9861,N_6110,N_6140);
or U9862 (N_9862,N_7364,N_6863);
nor U9863 (N_9863,N_6887,N_7679);
xnor U9864 (N_9864,N_6520,N_7692);
nand U9865 (N_9865,N_6479,N_6778);
and U9866 (N_9866,N_6225,N_7199);
and U9867 (N_9867,N_7780,N_7303);
nor U9868 (N_9868,N_7930,N_6803);
and U9869 (N_9869,N_7407,N_6183);
and U9870 (N_9870,N_7118,N_6756);
nand U9871 (N_9871,N_6958,N_6220);
nand U9872 (N_9872,N_7094,N_7864);
and U9873 (N_9873,N_7994,N_7326);
nand U9874 (N_9874,N_6635,N_6687);
nand U9875 (N_9875,N_7963,N_6310);
nand U9876 (N_9876,N_7514,N_6731);
nand U9877 (N_9877,N_7081,N_6374);
nor U9878 (N_9878,N_6850,N_7564);
xnor U9879 (N_9879,N_7742,N_6287);
or U9880 (N_9880,N_6696,N_6155);
and U9881 (N_9881,N_6734,N_7626);
nor U9882 (N_9882,N_7788,N_7719);
nor U9883 (N_9883,N_7615,N_6155);
nand U9884 (N_9884,N_7778,N_7609);
nor U9885 (N_9885,N_6109,N_7937);
nand U9886 (N_9886,N_7583,N_7123);
or U9887 (N_9887,N_7891,N_7194);
nand U9888 (N_9888,N_7795,N_6697);
or U9889 (N_9889,N_6066,N_6873);
nor U9890 (N_9890,N_7762,N_6864);
nand U9891 (N_9891,N_7723,N_6733);
nand U9892 (N_9892,N_7017,N_6323);
nor U9893 (N_9893,N_6386,N_6742);
nor U9894 (N_9894,N_6479,N_7922);
nand U9895 (N_9895,N_7173,N_7015);
nand U9896 (N_9896,N_7355,N_6268);
xor U9897 (N_9897,N_7873,N_7899);
or U9898 (N_9898,N_6299,N_7741);
nor U9899 (N_9899,N_6820,N_7157);
xnor U9900 (N_9900,N_6901,N_7330);
xor U9901 (N_9901,N_7552,N_6433);
and U9902 (N_9902,N_7742,N_6341);
nand U9903 (N_9903,N_6242,N_7540);
or U9904 (N_9904,N_6836,N_7685);
or U9905 (N_9905,N_7927,N_7212);
xor U9906 (N_9906,N_6052,N_7984);
or U9907 (N_9907,N_6108,N_7278);
nor U9908 (N_9908,N_6751,N_7922);
xor U9909 (N_9909,N_6201,N_7355);
nand U9910 (N_9910,N_6609,N_6664);
and U9911 (N_9911,N_6380,N_6573);
nand U9912 (N_9912,N_7896,N_6129);
or U9913 (N_9913,N_7762,N_7071);
nor U9914 (N_9914,N_7848,N_6066);
and U9915 (N_9915,N_6629,N_7340);
xnor U9916 (N_9916,N_6663,N_6262);
nor U9917 (N_9917,N_6334,N_6619);
or U9918 (N_9918,N_6700,N_7503);
nor U9919 (N_9919,N_6480,N_6472);
and U9920 (N_9920,N_6943,N_6881);
nor U9921 (N_9921,N_7036,N_7388);
nor U9922 (N_9922,N_6127,N_6583);
nand U9923 (N_9923,N_7652,N_7011);
nor U9924 (N_9924,N_7576,N_6387);
or U9925 (N_9925,N_7935,N_6041);
or U9926 (N_9926,N_6642,N_7070);
nor U9927 (N_9927,N_7961,N_6468);
xor U9928 (N_9928,N_7016,N_6247);
xor U9929 (N_9929,N_7279,N_6263);
and U9930 (N_9930,N_7270,N_7798);
or U9931 (N_9931,N_6562,N_6793);
xnor U9932 (N_9932,N_7566,N_6240);
nor U9933 (N_9933,N_7856,N_7776);
and U9934 (N_9934,N_7935,N_6704);
nor U9935 (N_9935,N_7965,N_7405);
nor U9936 (N_9936,N_7620,N_6145);
nor U9937 (N_9937,N_7301,N_7461);
nand U9938 (N_9938,N_7752,N_7991);
or U9939 (N_9939,N_6165,N_7298);
nand U9940 (N_9940,N_6718,N_6908);
xor U9941 (N_9941,N_6568,N_7073);
xnor U9942 (N_9942,N_6345,N_6765);
and U9943 (N_9943,N_6406,N_6829);
nor U9944 (N_9944,N_6307,N_7312);
xor U9945 (N_9945,N_6579,N_6409);
xnor U9946 (N_9946,N_7527,N_6711);
and U9947 (N_9947,N_6835,N_6241);
or U9948 (N_9948,N_6668,N_6302);
xor U9949 (N_9949,N_6957,N_6234);
nor U9950 (N_9950,N_7397,N_6547);
xor U9951 (N_9951,N_6667,N_6955);
nand U9952 (N_9952,N_6005,N_7071);
nor U9953 (N_9953,N_7048,N_6589);
and U9954 (N_9954,N_6691,N_7601);
and U9955 (N_9955,N_7484,N_7170);
and U9956 (N_9956,N_6547,N_7829);
nand U9957 (N_9957,N_6396,N_7324);
and U9958 (N_9958,N_6159,N_7941);
nand U9959 (N_9959,N_7793,N_6984);
nor U9960 (N_9960,N_6635,N_6652);
nand U9961 (N_9961,N_6611,N_6814);
or U9962 (N_9962,N_6446,N_6950);
nor U9963 (N_9963,N_6053,N_6059);
nor U9964 (N_9964,N_6788,N_7882);
and U9965 (N_9965,N_6430,N_6100);
xnor U9966 (N_9966,N_6056,N_6510);
xor U9967 (N_9967,N_6324,N_7804);
nand U9968 (N_9968,N_6350,N_7504);
xor U9969 (N_9969,N_6523,N_6140);
xnor U9970 (N_9970,N_6510,N_7206);
nand U9971 (N_9971,N_6256,N_6344);
xor U9972 (N_9972,N_6915,N_6968);
xor U9973 (N_9973,N_7563,N_6348);
and U9974 (N_9974,N_7906,N_7381);
or U9975 (N_9975,N_6999,N_6473);
or U9976 (N_9976,N_6099,N_7938);
or U9977 (N_9977,N_7324,N_7787);
or U9978 (N_9978,N_7404,N_7962);
or U9979 (N_9979,N_7083,N_7178);
nand U9980 (N_9980,N_6821,N_7087);
nor U9981 (N_9981,N_6944,N_7066);
nand U9982 (N_9982,N_6927,N_6801);
and U9983 (N_9983,N_7653,N_6058);
and U9984 (N_9984,N_7815,N_7664);
nor U9985 (N_9985,N_6984,N_6334);
nand U9986 (N_9986,N_6651,N_6384);
xnor U9987 (N_9987,N_7659,N_7638);
nor U9988 (N_9988,N_6035,N_6862);
or U9989 (N_9989,N_6055,N_7890);
and U9990 (N_9990,N_6873,N_7507);
nor U9991 (N_9991,N_6228,N_7893);
or U9992 (N_9992,N_6355,N_6194);
nand U9993 (N_9993,N_6558,N_7431);
or U9994 (N_9994,N_7231,N_7461);
nor U9995 (N_9995,N_6627,N_6877);
nand U9996 (N_9996,N_7354,N_6682);
and U9997 (N_9997,N_6527,N_7708);
nand U9998 (N_9998,N_7982,N_6305);
and U9999 (N_9999,N_6939,N_6051);
or U10000 (N_10000,N_8969,N_9375);
xor U10001 (N_10001,N_9923,N_8937);
nand U10002 (N_10002,N_9719,N_9631);
and U10003 (N_10003,N_8290,N_8305);
and U10004 (N_10004,N_8180,N_9304);
or U10005 (N_10005,N_8995,N_8485);
or U10006 (N_10006,N_9232,N_9668);
nand U10007 (N_10007,N_9676,N_8943);
xor U10008 (N_10008,N_8516,N_8585);
xor U10009 (N_10009,N_9750,N_8751);
xnor U10010 (N_10010,N_8131,N_8138);
and U10011 (N_10011,N_9553,N_8438);
or U10012 (N_10012,N_9595,N_8467);
nor U10013 (N_10013,N_9885,N_9773);
nor U10014 (N_10014,N_8491,N_9052);
nand U10015 (N_10015,N_9729,N_8448);
or U10016 (N_10016,N_9662,N_8096);
and U10017 (N_10017,N_8837,N_8222);
xnor U10018 (N_10018,N_9563,N_9366);
and U10019 (N_10019,N_8980,N_8699);
nor U10020 (N_10020,N_8115,N_9382);
nor U10021 (N_10021,N_9428,N_9368);
nor U10022 (N_10022,N_9878,N_9852);
or U10023 (N_10023,N_9578,N_8089);
or U10024 (N_10024,N_9126,N_8850);
nand U10025 (N_10025,N_9021,N_8679);
xnor U10026 (N_10026,N_9141,N_8987);
or U10027 (N_10027,N_8554,N_8122);
nor U10028 (N_10028,N_8879,N_9624);
nor U10029 (N_10029,N_8403,N_9127);
nor U10030 (N_10030,N_9854,N_9308);
xor U10031 (N_10031,N_9910,N_9935);
nor U10032 (N_10032,N_9986,N_8855);
xnor U10033 (N_10033,N_9797,N_8731);
xor U10034 (N_10034,N_9765,N_8001);
or U10035 (N_10035,N_9206,N_9476);
nor U10036 (N_10036,N_8050,N_9350);
or U10037 (N_10037,N_8375,N_9969);
nand U10038 (N_10038,N_9786,N_9282);
nor U10039 (N_10039,N_9680,N_8301);
and U10040 (N_10040,N_8727,N_8159);
nand U10041 (N_10041,N_8744,N_9734);
and U10042 (N_10042,N_8640,N_8259);
xor U10043 (N_10043,N_9877,N_9023);
xor U10044 (N_10044,N_8875,N_9748);
or U10045 (N_10045,N_9086,N_8674);
nor U10046 (N_10046,N_9186,N_8016);
or U10047 (N_10047,N_8595,N_8144);
xor U10048 (N_10048,N_9900,N_9699);
or U10049 (N_10049,N_8657,N_9795);
nor U10050 (N_10050,N_8346,N_8120);
and U10051 (N_10051,N_9567,N_9669);
xnor U10052 (N_10052,N_8619,N_9293);
xor U10053 (N_10053,N_9303,N_8005);
nand U10054 (N_10054,N_9770,N_9889);
nor U10055 (N_10055,N_9895,N_8726);
nand U10056 (N_10056,N_9180,N_9971);
xor U10057 (N_10057,N_9510,N_8009);
nor U10058 (N_10058,N_9035,N_9159);
nand U10059 (N_10059,N_8368,N_9735);
and U10060 (N_10060,N_9262,N_8559);
or U10061 (N_10061,N_8062,N_9164);
xor U10062 (N_10062,N_9808,N_9656);
and U10063 (N_10063,N_8832,N_9416);
nor U10064 (N_10064,N_9178,N_9201);
nor U10065 (N_10065,N_8454,N_8464);
or U10066 (N_10066,N_8961,N_9477);
xnor U10067 (N_10067,N_9810,N_8757);
nand U10068 (N_10068,N_9414,N_8999);
nand U10069 (N_10069,N_8521,N_8265);
or U10070 (N_10070,N_8897,N_8064);
and U10071 (N_10071,N_8538,N_8019);
or U10072 (N_10072,N_8351,N_8091);
or U10073 (N_10073,N_9242,N_9427);
nand U10074 (N_10074,N_8246,N_9523);
nand U10075 (N_10075,N_8769,N_9988);
nor U10076 (N_10076,N_8851,N_9783);
and U10077 (N_10077,N_8904,N_8917);
or U10078 (N_10078,N_8208,N_9198);
and U10079 (N_10079,N_8866,N_9799);
nor U10080 (N_10080,N_8379,N_8313);
or U10081 (N_10081,N_8027,N_9079);
nand U10082 (N_10082,N_9049,N_8892);
or U10083 (N_10083,N_9949,N_9845);
xor U10084 (N_10084,N_9913,N_8022);
nor U10085 (N_10085,N_9564,N_9939);
xor U10086 (N_10086,N_9492,N_8788);
nand U10087 (N_10087,N_9485,N_8548);
xnor U10088 (N_10088,N_9957,N_9015);
nor U10089 (N_10089,N_9468,N_9214);
or U10090 (N_10090,N_8603,N_8911);
nand U10091 (N_10091,N_8841,N_8630);
nand U10092 (N_10092,N_8692,N_9531);
or U10093 (N_10093,N_9431,N_9752);
and U10094 (N_10094,N_8371,N_9310);
xor U10095 (N_10095,N_9334,N_8030);
nor U10096 (N_10096,N_8746,N_9784);
nor U10097 (N_10097,N_9276,N_9705);
xnor U10098 (N_10098,N_8785,N_8730);
xor U10099 (N_10099,N_9514,N_9486);
nand U10100 (N_10100,N_9311,N_9634);
nand U10101 (N_10101,N_9886,N_9220);
and U10102 (N_10102,N_8354,N_8452);
or U10103 (N_10103,N_8444,N_8772);
and U10104 (N_10104,N_8971,N_9400);
and U10105 (N_10105,N_8581,N_8325);
and U10106 (N_10106,N_8948,N_9767);
or U10107 (N_10107,N_9073,N_9793);
nand U10108 (N_10108,N_8473,N_8939);
nor U10109 (N_10109,N_8577,N_9391);
nand U10110 (N_10110,N_8938,N_8658);
nor U10111 (N_10111,N_9029,N_9619);
nand U10112 (N_10112,N_8076,N_9365);
and U10113 (N_10113,N_9273,N_9299);
or U10114 (N_10114,N_8041,N_9807);
and U10115 (N_10115,N_8528,N_8736);
or U10116 (N_10116,N_8154,N_9608);
xor U10117 (N_10117,N_9157,N_9881);
and U10118 (N_10118,N_8712,N_8389);
xor U10119 (N_10119,N_9363,N_9353);
or U10120 (N_10120,N_8953,N_8037);
nor U10121 (N_10121,N_8517,N_9067);
and U10122 (N_10122,N_8298,N_9134);
or U10123 (N_10123,N_8654,N_8197);
or U10124 (N_10124,N_9392,N_8890);
and U10125 (N_10125,N_9947,N_8775);
or U10126 (N_10126,N_9140,N_9535);
nor U10127 (N_10127,N_8113,N_8213);
and U10128 (N_10128,N_8275,N_9016);
nor U10129 (N_10129,N_9494,N_8251);
and U10130 (N_10130,N_9051,N_9243);
nand U10131 (N_10131,N_9686,N_8916);
nor U10132 (N_10132,N_8578,N_9867);
xor U10133 (N_10133,N_8139,N_8795);
nor U10134 (N_10134,N_9459,N_9280);
xor U10135 (N_10135,N_9199,N_9862);
xor U10136 (N_10136,N_8622,N_8912);
and U10137 (N_10137,N_8359,N_9707);
nor U10138 (N_10138,N_8253,N_8596);
or U10139 (N_10139,N_8886,N_9866);
nor U10140 (N_10140,N_8592,N_9483);
nand U10141 (N_10141,N_9339,N_8484);
nand U10142 (N_10142,N_8922,N_8176);
or U10143 (N_10143,N_8803,N_8461);
nor U10144 (N_10144,N_8449,N_9641);
nor U10145 (N_10145,N_8898,N_9039);
nand U10146 (N_10146,N_9708,N_9458);
and U10147 (N_10147,N_9925,N_8966);
and U10148 (N_10148,N_8196,N_8593);
nor U10149 (N_10149,N_9471,N_9008);
or U10150 (N_10150,N_9905,N_9462);
or U10151 (N_10151,N_9024,N_8807);
nor U10152 (N_10152,N_8299,N_9060);
or U10153 (N_10153,N_8386,N_8935);
or U10154 (N_10154,N_9106,N_8084);
xnor U10155 (N_10155,N_9628,N_9706);
nand U10156 (N_10156,N_8771,N_8340);
and U10157 (N_10157,N_9283,N_9150);
or U10158 (N_10158,N_8157,N_8686);
nand U10159 (N_10159,N_9192,N_8993);
or U10160 (N_10160,N_9075,N_9521);
nand U10161 (N_10161,N_9110,N_8681);
xnor U10162 (N_10162,N_9166,N_8295);
or U10163 (N_10163,N_8069,N_9644);
nand U10164 (N_10164,N_8814,N_9948);
xor U10165 (N_10165,N_8535,N_8306);
or U10166 (N_10166,N_8576,N_9170);
nor U10167 (N_10167,N_9507,N_8921);
xor U10168 (N_10168,N_8008,N_9014);
xnor U10169 (N_10169,N_9167,N_8732);
or U10170 (N_10170,N_9020,N_9371);
or U10171 (N_10171,N_8219,N_9518);
nand U10172 (N_10172,N_9831,N_9978);
nor U10173 (N_10173,N_8924,N_9983);
nor U10174 (N_10174,N_9010,N_8767);
xor U10175 (N_10175,N_9244,N_8840);
nand U10176 (N_10176,N_9519,N_8025);
nand U10177 (N_10177,N_9102,N_9697);
nor U10178 (N_10178,N_9314,N_9464);
nor U10179 (N_10179,N_8844,N_8988);
xnor U10180 (N_10180,N_9187,N_8315);
or U10181 (N_10181,N_9078,N_9745);
or U10182 (N_10182,N_8737,N_9069);
or U10183 (N_10183,N_9824,N_8136);
nor U10184 (N_10184,N_8616,N_8662);
nand U10185 (N_10185,N_9162,N_9747);
nor U10186 (N_10186,N_8205,N_8796);
or U10187 (N_10187,N_8017,N_8615);
xnor U10188 (N_10188,N_8335,N_9076);
xor U10189 (N_10189,N_9355,N_8942);
xnor U10190 (N_10190,N_8905,N_8116);
nand U10191 (N_10191,N_9144,N_9582);
or U10192 (N_10192,N_9099,N_9149);
nand U10193 (N_10193,N_9530,N_9466);
or U10194 (N_10194,N_8468,N_8831);
xor U10195 (N_10195,N_8469,N_8446);
nor U10196 (N_10196,N_8040,N_8542);
or U10197 (N_10197,N_9426,N_8989);
nand U10198 (N_10198,N_8230,N_8811);
nand U10199 (N_10199,N_9250,N_8445);
nand U10200 (N_10200,N_8045,N_9586);
xnor U10201 (N_10201,N_9440,N_8612);
nor U10202 (N_10202,N_8264,N_9216);
or U10203 (N_10203,N_8678,N_9671);
nand U10204 (N_10204,N_9826,N_8475);
nand U10205 (N_10205,N_9114,N_9038);
nor U10206 (N_10206,N_9924,N_9288);
and U10207 (N_10207,N_8617,N_8863);
and U10208 (N_10208,N_8967,N_9843);
nand U10209 (N_10209,N_9876,N_8682);
or U10210 (N_10210,N_8433,N_9221);
nand U10211 (N_10211,N_9962,N_9522);
nand U10212 (N_10212,N_8323,N_9543);
and U10213 (N_10213,N_8716,N_9028);
xor U10214 (N_10214,N_9160,N_8195);
nor U10215 (N_10215,N_8053,N_8412);
nor U10216 (N_10216,N_9871,N_9329);
xnor U10217 (N_10217,N_9196,N_8470);
nor U10218 (N_10218,N_9951,N_8293);
nand U10219 (N_10219,N_8199,N_8909);
nor U10220 (N_10220,N_8319,N_8366);
nor U10221 (N_10221,N_9835,N_9987);
or U10222 (N_10222,N_9480,N_8234);
and U10223 (N_10223,N_9724,N_8228);
and U10224 (N_10224,N_9657,N_9224);
xnor U10225 (N_10225,N_9761,N_9456);
xor U10226 (N_10226,N_8297,N_8914);
and U10227 (N_10227,N_9812,N_8443);
and U10228 (N_10228,N_8407,N_8128);
and U10229 (N_10229,N_8854,N_9333);
xor U10230 (N_10230,N_9238,N_8164);
and U10231 (N_10231,N_9135,N_9819);
and U10232 (N_10232,N_9768,N_8170);
nand U10233 (N_10233,N_9723,N_9335);
or U10234 (N_10234,N_9960,N_9025);
nor U10235 (N_10235,N_9241,N_9615);
and U10236 (N_10236,N_9357,N_9146);
nand U10237 (N_10237,N_8507,N_9848);
nand U10238 (N_10238,N_8573,N_8479);
and U10239 (N_10239,N_8247,N_8110);
or U10240 (N_10240,N_8787,N_8970);
or U10241 (N_10241,N_8959,N_9248);
and U10242 (N_10242,N_8294,N_8758);
nor U10243 (N_10243,N_9091,N_9124);
and U10244 (N_10244,N_8387,N_8608);
nor U10245 (N_10245,N_9551,N_9785);
nor U10246 (N_10246,N_9129,N_8415);
or U10247 (N_10247,N_8777,N_8474);
nand U10248 (N_10248,N_9070,N_9133);
and U10249 (N_10249,N_8644,N_9901);
nor U10250 (N_10250,N_8931,N_9554);
xor U10251 (N_10251,N_9270,N_8376);
and U10252 (N_10252,N_8702,N_8129);
nand U10253 (N_10253,N_8423,N_9300);
or U10254 (N_10254,N_8843,N_8722);
or U10255 (N_10255,N_9568,N_8348);
nor U10256 (N_10256,N_9573,N_9019);
or U10257 (N_10257,N_8383,N_9090);
xor U10258 (N_10258,N_8893,N_9571);
xnor U10259 (N_10259,N_9092,N_9614);
and U10260 (N_10260,N_8172,N_8639);
nor U10261 (N_10261,N_8127,N_9976);
nor U10262 (N_10262,N_9269,N_8400);
nor U10263 (N_10263,N_8891,N_9229);
nor U10264 (N_10264,N_9666,N_9764);
nand U10265 (N_10265,N_8026,N_8123);
or U10266 (N_10266,N_9646,N_9756);
nand U10267 (N_10267,N_9207,N_8887);
and U10268 (N_10268,N_8508,N_9804);
nand U10269 (N_10269,N_8108,N_9181);
nand U10270 (N_10270,N_9902,N_8677);
xor U10271 (N_10271,N_9089,N_9922);
nor U10272 (N_10272,N_9694,N_9147);
or U10273 (N_10273,N_8838,N_9683);
nand U10274 (N_10274,N_8033,N_9423);
and U10275 (N_10275,N_9246,N_9968);
nor U10276 (N_10276,N_9593,N_8761);
or U10277 (N_10277,N_8856,N_8109);
and U10278 (N_10278,N_8688,N_9513);
nor U10279 (N_10279,N_8867,N_9673);
nor U10280 (N_10280,N_8309,N_8582);
xor U10281 (N_10281,N_9284,N_9585);
nor U10282 (N_10282,N_9237,N_9703);
nor U10283 (N_10283,N_9690,N_8384);
or U10284 (N_10284,N_8551,N_9364);
and U10285 (N_10285,N_9481,N_9006);
nand U10286 (N_10286,N_9626,N_8362);
xnor U10287 (N_10287,N_8604,N_8557);
nand U10288 (N_10288,N_9063,N_8532);
and U10289 (N_10289,N_8072,N_9447);
nor U10290 (N_10290,N_8784,N_9378);
xnor U10291 (N_10291,N_9583,N_8958);
or U10292 (N_10292,N_8566,N_9463);
or U10293 (N_10293,N_8206,N_9687);
xnor U10294 (N_10294,N_8598,N_9528);
or U10295 (N_10295,N_9704,N_8952);
and U10296 (N_10296,N_8248,N_9744);
or U10297 (N_10297,N_8738,N_8003);
or U10298 (N_10298,N_9544,N_8283);
or U10299 (N_10299,N_9562,N_9825);
or U10300 (N_10300,N_8882,N_9332);
xnor U10301 (N_10301,N_9974,N_9251);
xor U10302 (N_10302,N_8870,N_8960);
xnor U10303 (N_10303,N_8156,N_9491);
nor U10304 (N_10304,N_8816,N_8515);
nor U10305 (N_10305,N_9596,N_9658);
xor U10306 (N_10306,N_8261,N_8365);
and U10307 (N_10307,N_8105,N_8990);
or U10308 (N_10308,N_9610,N_8719);
nand U10309 (N_10309,N_8029,N_9377);
xor U10310 (N_10310,N_8575,N_9636);
nor U10311 (N_10311,N_9194,N_8011);
and U10312 (N_10312,N_8160,N_8162);
nand U10313 (N_10313,N_9053,N_9839);
or U10314 (N_10314,N_8895,N_9853);
nor U10315 (N_10315,N_8530,N_9439);
nor U10316 (N_10316,N_9442,N_9574);
or U10317 (N_10317,N_8104,N_8018);
or U10318 (N_10318,N_9601,N_9632);
and U10319 (N_10319,N_8168,N_9286);
or U10320 (N_10320,N_9849,N_8951);
nor U10321 (N_10321,N_9322,N_9712);
or U10322 (N_10322,N_8773,N_8986);
nand U10323 (N_10323,N_9236,N_9200);
and U10324 (N_10324,N_8286,N_8865);
nor U10325 (N_10325,N_9163,N_8057);
xor U10326 (N_10326,N_8133,N_8497);
or U10327 (N_10327,N_9370,N_9331);
nor U10328 (N_10328,N_8547,N_9139);
and U10329 (N_10329,N_8896,N_9208);
nor U10330 (N_10330,N_8266,N_9277);
xor U10331 (N_10331,N_8087,N_8546);
nor U10332 (N_10332,N_8745,N_9591);
nand U10333 (N_10333,N_9112,N_9555);
and U10334 (N_10334,N_8881,N_9077);
nor U10335 (N_10335,N_8178,N_8556);
or U10336 (N_10336,N_8839,N_8928);
and U10337 (N_10337,N_8137,N_8095);
and U10338 (N_10338,N_9105,N_9472);
xnor U10339 (N_10339,N_9572,N_9319);
nor U10340 (N_10340,N_8974,N_9418);
xor U10341 (N_10341,N_8793,N_9190);
or U10342 (N_10342,N_9235,N_9561);
nor U10343 (N_10343,N_8304,N_9965);
nor U10344 (N_10344,N_9757,N_9343);
or U10345 (N_10345,N_9725,N_8397);
nand U10346 (N_10346,N_9711,N_9088);
xnor U10347 (N_10347,N_8963,N_9302);
nand U10348 (N_10348,N_8460,N_8262);
nand U10349 (N_10349,N_8915,N_9045);
nand U10350 (N_10350,N_8106,N_9295);
nor U10351 (N_10351,N_9788,N_9637);
nand U10352 (N_10352,N_8859,N_8550);
xor U10353 (N_10353,N_8425,N_8392);
or U10354 (N_10354,N_9640,N_8975);
xor U10355 (N_10355,N_8908,N_8250);
xor U10356 (N_10356,N_8028,N_8427);
and U10357 (N_10357,N_8277,N_9228);
nor U10358 (N_10358,N_8358,N_9087);
xor U10359 (N_10359,N_8725,N_8889);
nand U10360 (N_10360,N_8192,N_8165);
or U10361 (N_10361,N_9718,N_8077);
or U10362 (N_10362,N_8142,N_9130);
nand U10363 (N_10363,N_9000,N_8501);
or U10364 (N_10364,N_8601,N_9672);
nand U10365 (N_10365,N_8606,N_9432);
or U10366 (N_10366,N_8329,N_9281);
xnor U10367 (N_10367,N_8512,N_9171);
xor U10368 (N_10368,N_8442,N_9037);
and U10369 (N_10369,N_8241,N_9057);
or U10370 (N_10370,N_9546,N_9920);
nor U10371 (N_10371,N_8821,N_9805);
and U10372 (N_10372,N_8780,N_9222);
xnor U10373 (N_10373,N_9473,N_9663);
and U10374 (N_10374,N_9611,N_8571);
xnor U10375 (N_10375,N_9465,N_9980);
nand U10376 (N_10376,N_9800,N_8272);
nand U10377 (N_10377,N_8631,N_9880);
and U10378 (N_10378,N_8620,N_9356);
or U10379 (N_10379,N_8079,N_8390);
and U10380 (N_10380,N_8704,N_8363);
or U10381 (N_10381,N_8169,N_9675);
and U10382 (N_10382,N_8059,N_9966);
nand U10383 (N_10383,N_9802,N_8884);
xor U10384 (N_10384,N_9113,N_9959);
xor U10385 (N_10385,N_9909,N_8307);
nor U10386 (N_10386,N_8352,N_9501);
nand U10387 (N_10387,N_9137,N_8391);
and U10388 (N_10388,N_8536,N_8268);
xnor U10389 (N_10389,N_8878,N_8919);
nand U10390 (N_10390,N_9929,N_8827);
or U10391 (N_10391,N_9142,N_8225);
xnor U10392 (N_10392,N_9500,N_9009);
or U10393 (N_10393,N_8393,N_8718);
and U10394 (N_10394,N_9257,N_8260);
and U10395 (N_10395,N_8683,N_8698);
nand U10396 (N_10396,N_8539,N_8429);
and U10397 (N_10397,N_9738,N_8976);
nand U10398 (N_10398,N_8524,N_8308);
or U10399 (N_10399,N_9556,N_8060);
or U10400 (N_10400,N_8355,N_9858);
nor U10401 (N_10401,N_9384,N_9434);
nor U10402 (N_10402,N_8944,N_9047);
nand U10403 (N_10403,N_9916,N_8957);
or U10404 (N_10404,N_8885,N_8347);
nand U10405 (N_10405,N_9525,N_9495);
and U10406 (N_10406,N_9478,N_9512);
xor U10407 (N_10407,N_8013,N_8242);
and U10408 (N_10408,N_9892,N_8276);
nand U10409 (N_10409,N_8665,N_9374);
or U10410 (N_10410,N_9497,N_9504);
nand U10411 (N_10411,N_9685,N_8861);
and U10412 (N_10412,N_9975,N_8078);
nand U10413 (N_10413,N_8666,N_8950);
or U10414 (N_10414,N_8254,N_8171);
nor U10415 (N_10415,N_8941,N_9155);
xnor U10416 (N_10416,N_8140,N_9681);
and U10417 (N_10417,N_8669,N_9763);
and U10418 (N_10418,N_8372,N_9732);
nand U10419 (N_10419,N_8428,N_9717);
or U10420 (N_10420,N_8086,N_8006);
xor U10421 (N_10421,N_9515,N_8012);
xnor U10422 (N_10422,N_8395,N_8070);
or U10423 (N_10423,N_9891,N_8519);
and U10424 (N_10424,N_8637,N_9787);
and U10425 (N_10425,N_9508,N_9074);
nor U10426 (N_10426,N_8167,N_8094);
and U10427 (N_10427,N_8733,N_8152);
and U10428 (N_10428,N_9505,N_9271);
and U10429 (N_10429,N_8804,N_8215);
nand U10430 (N_10430,N_8054,N_8404);
nor U10431 (N_10431,N_8965,N_8002);
nand U10432 (N_10432,N_9930,N_9204);
nor U10433 (N_10433,N_8690,N_8709);
or U10434 (N_10434,N_9823,N_9780);
and U10435 (N_10435,N_8798,N_9347);
xor U10436 (N_10436,N_8742,N_9827);
and U10437 (N_10437,N_8321,N_9046);
nor U10438 (N_10438,N_9443,N_9817);
nor U10439 (N_10439,N_9760,N_9639);
nor U10440 (N_10440,N_9390,N_9234);
nand U10441 (N_10441,N_8609,N_8098);
nor U10442 (N_10442,N_9449,N_9684);
nor U10443 (N_10443,N_9055,N_8910);
or U10444 (N_10444,N_9818,N_9184);
and U10445 (N_10445,N_8764,N_9996);
and U10446 (N_10446,N_8752,N_9813);
or U10447 (N_10447,N_9677,N_9660);
xnor U10448 (N_10448,N_9450,N_8800);
and U10449 (N_10449,N_9851,N_8143);
xor U10450 (N_10450,N_8531,N_8421);
and U10451 (N_10451,N_9942,N_8177);
nand U10452 (N_10452,N_9205,N_9383);
and U10453 (N_10453,N_9231,N_8982);
nand U10454 (N_10454,N_9175,N_9145);
nand U10455 (N_10455,N_9991,N_9433);
xnor U10456 (N_10456,N_9064,N_8860);
or U10457 (N_10457,N_9517,N_9781);
and U10458 (N_10458,N_9584,N_8587);
and U10459 (N_10459,N_8877,N_8147);
nor U10460 (N_10460,N_9549,N_8034);
and U10461 (N_10461,N_9590,N_8332);
and U10462 (N_10462,N_8229,N_9954);
nor U10463 (N_10463,N_8211,N_9602);
nand U10464 (N_10464,N_8201,N_8361);
or U10465 (N_10465,N_9926,N_9225);
nand U10466 (N_10466,N_9451,N_9183);
or U10467 (N_10467,N_9402,N_9606);
and U10468 (N_10468,N_8711,N_9362);
xnor U10469 (N_10469,N_8755,N_8422);
or U10470 (N_10470,N_8563,N_9301);
and U10471 (N_10471,N_8488,N_9887);
or U10472 (N_10472,N_8472,N_9566);
nor U10473 (N_10473,N_8327,N_8207);
and U10474 (N_10474,N_8426,N_9188);
or U10475 (N_10475,N_9217,N_8097);
or U10476 (N_10476,N_8155,N_8405);
and U10477 (N_10477,N_8061,N_8588);
or U10478 (N_10478,N_8820,N_9550);
or U10479 (N_10479,N_9796,N_8537);
nor U10480 (N_10480,N_8161,N_9017);
nor U10481 (N_10481,N_8249,N_8151);
or U10482 (N_10482,N_8694,N_8697);
and U10483 (N_10483,N_9457,N_9545);
nand U10484 (N_10484,N_9430,N_9645);
nand U10485 (N_10485,N_9307,N_8858);
and U10486 (N_10486,N_8118,N_9227);
or U10487 (N_10487,N_8936,N_8983);
and U10488 (N_10488,N_9026,N_8656);
or U10489 (N_10489,N_8985,N_8710);
nand U10490 (N_10490,N_9503,N_8728);
and U10491 (N_10491,N_8907,N_9801);
nand U10492 (N_10492,N_8130,N_8845);
nor U10493 (N_10493,N_9318,N_9218);
or U10494 (N_10494,N_9226,N_8090);
nor U10495 (N_10495,N_9811,N_8480);
nand U10496 (N_10496,N_8614,N_9899);
nor U10497 (N_10497,N_9309,N_9758);
xor U10498 (N_10498,N_9109,N_9674);
or U10499 (N_10499,N_8634,N_8994);
nand U10500 (N_10500,N_8673,N_9202);
nand U10501 (N_10501,N_9984,N_9897);
nand U10502 (N_10502,N_9529,N_8227);
or U10503 (N_10503,N_9179,N_9570);
nand U10504 (N_10504,N_9828,N_9575);
nor U10505 (N_10505,N_8280,N_9148);
nor U10506 (N_10506,N_9132,N_8065);
and U10507 (N_10507,N_8316,N_9789);
and U10508 (N_10508,N_9937,N_9328);
nand U10509 (N_10509,N_8432,N_9952);
nor U10510 (N_10510,N_8545,N_9420);
and U10511 (N_10511,N_8646,N_8552);
or U10512 (N_10512,N_8570,N_9185);
or U10513 (N_10513,N_9569,N_8453);
xor U10514 (N_10514,N_9361,N_8713);
nor U10515 (N_10515,N_9098,N_9290);
xnor U10516 (N_10516,N_9031,N_8659);
xor U10517 (N_10517,N_8774,N_9613);
and U10518 (N_10518,N_8900,N_9888);
xor U10519 (N_10519,N_8344,N_8287);
nand U10520 (N_10520,N_8408,N_9095);
and U10521 (N_10521,N_8493,N_8633);
xnor U10522 (N_10522,N_9413,N_9741);
or U10523 (N_10523,N_8797,N_9419);
or U10524 (N_10524,N_9174,N_8973);
and U10525 (N_10525,N_8871,N_9082);
and U10526 (N_10526,N_8600,N_9903);
nor U10527 (N_10527,N_8223,N_9598);
and U10528 (N_10528,N_8714,N_8613);
nand U10529 (N_10529,N_9169,N_9771);
nor U10530 (N_10530,N_9928,N_9516);
and U10531 (N_10531,N_8166,N_9855);
xor U10532 (N_10532,N_9772,N_8490);
nand U10533 (N_10533,N_9272,N_8124);
nand U10534 (N_10534,N_8342,N_9345);
nand U10535 (N_10535,N_8465,N_9890);
xnor U10536 (N_10536,N_9609,N_8221);
or U10537 (N_10537,N_9981,N_9832);
and U10538 (N_10538,N_8930,N_9742);
nand U10539 (N_10539,N_8288,N_9746);
and U10540 (N_10540,N_8257,N_9769);
and U10541 (N_10541,N_8753,N_9018);
nor U10542 (N_10542,N_8792,N_8781);
nor U10543 (N_10543,N_8252,N_8477);
or U10544 (N_10544,N_8607,N_8946);
nand U10545 (N_10545,N_9873,N_9482);
nand U10546 (N_10546,N_8406,N_9212);
nor U10547 (N_10547,N_8014,N_9943);
nor U10548 (N_10548,N_9104,N_9197);
xnor U10549 (N_10549,N_8085,N_8701);
or U10550 (N_10550,N_8135,N_8954);
nand U10551 (N_10551,N_8083,N_8852);
xor U10552 (N_10552,N_9189,N_8194);
or U10553 (N_10553,N_9223,N_9404);
and U10554 (N_10554,N_9806,N_9868);
or U10555 (N_10555,N_9211,N_8876);
and U10556 (N_10556,N_9123,N_9274);
xor U10557 (N_10557,N_9870,N_9306);
nor U10558 (N_10558,N_9651,N_9992);
xnor U10559 (N_10559,N_8883,N_9933);
nand U10560 (N_10560,N_8112,N_9193);
or U10561 (N_10561,N_8451,N_8068);
or U10562 (N_10562,N_8273,N_9395);
or U10563 (N_10563,N_8345,N_8431);
nand U10564 (N_10564,N_8463,N_8093);
or U10565 (N_10565,N_8430,N_9094);
xor U10566 (N_10566,N_9315,N_8652);
nor U10567 (N_10567,N_8968,N_9253);
or U10568 (N_10568,N_9511,N_9898);
xor U10569 (N_10569,N_8927,N_9397);
nand U10570 (N_10570,N_9814,N_9403);
nand U10571 (N_10571,N_9444,N_9240);
nand U10572 (N_10572,N_8747,N_9857);
or U10573 (N_10573,N_8239,N_9066);
nand U10574 (N_10574,N_9093,N_9438);
nor U10575 (N_10575,N_8783,N_8148);
nand U10576 (N_10576,N_9999,N_8218);
nand U10577 (N_10577,N_9998,N_9592);
or U10578 (N_10578,N_9325,N_9979);
and U10579 (N_10579,N_9625,N_9861);
nor U10580 (N_10580,N_8399,N_9172);
xor U10581 (N_10581,N_8868,N_9537);
xnor U10582 (N_10582,N_8672,N_9260);
or U10583 (N_10583,N_8163,N_9594);
nand U10584 (N_10584,N_8232,N_8434);
nand U10585 (N_10585,N_8826,N_9557);
and U10586 (N_10586,N_8956,N_9847);
xnor U10587 (N_10587,N_8805,N_8322);
and U10588 (N_10588,N_9386,N_9359);
nor U10589 (N_10589,N_8216,N_8992);
nand U10590 (N_10590,N_8047,N_9844);
and U10591 (N_10591,N_8689,N_9617);
nor U10592 (N_10592,N_9219,N_9062);
and U10593 (N_10593,N_9421,N_8526);
or U10594 (N_10594,N_9798,N_8696);
xnor U10595 (N_10595,N_9003,N_9349);
nand U10596 (N_10596,N_8739,N_9883);
nor U10597 (N_10597,N_8506,N_8661);
nor U10598 (N_10598,N_9896,N_8031);
nor U10599 (N_10599,N_8561,N_8303);
or U10600 (N_10600,N_9713,N_8934);
and U10601 (N_10601,N_8720,N_8190);
and U10602 (N_10602,N_8735,N_9372);
nand U10603 (N_10603,N_9279,N_8754);
or U10604 (N_10604,N_8641,N_8502);
or U10605 (N_10605,N_9007,N_9520);
nor U10606 (N_10606,N_9577,N_9875);
xnor U10607 (N_10607,N_9605,N_8409);
nand U10608 (N_10608,N_8191,N_8184);
xor U10609 (N_10609,N_8117,N_9401);
and U10610 (N_10610,N_8705,N_8768);
and U10611 (N_10611,N_8349,N_9581);
nor U10612 (N_10612,N_9941,N_8602);
nor U10613 (N_10613,N_8707,N_9351);
or U10614 (N_10614,N_8700,N_9822);
nor U10615 (N_10615,N_8459,N_8869);
nor U10616 (N_10616,N_9532,N_8183);
and U10617 (N_10617,N_8763,N_9004);
xnor U10618 (N_10618,N_9940,N_9589);
xor U10619 (N_10619,N_8623,N_9932);
xor U10620 (N_10620,N_9213,N_8906);
nor U10621 (N_10621,N_9816,N_8802);
nor U10622 (N_10622,N_8036,N_8779);
or U10623 (N_10623,N_9970,N_9158);
and U10624 (N_10624,N_8353,N_9499);
nand U10625 (N_10625,N_8255,N_8830);
or U10626 (N_10626,N_8828,N_9101);
xnor U10627 (N_10627,N_9367,N_8092);
xor U10628 (N_10628,N_9714,N_8567);
xnor U10629 (N_10629,N_8534,N_8317);
or U10630 (N_10630,N_9252,N_8075);
and U10631 (N_10631,N_9864,N_9638);
xnor U10632 (N_10632,N_9406,N_9346);
and U10633 (N_10633,N_8145,N_8413);
nor U10634 (N_10634,N_8670,N_9080);
nor U10635 (N_10635,N_8023,N_8498);
xnor U10636 (N_10636,N_9002,N_9267);
or U10637 (N_10637,N_9239,N_9005);
nand U10638 (N_10638,N_8328,N_8649);
xor U10639 (N_10639,N_8173,N_8334);
nand U10640 (N_10640,N_8455,N_8284);
and U10641 (N_10641,N_8790,N_8274);
nand U10642 (N_10642,N_8642,N_8326);
and U10643 (N_10643,N_9548,N_9389);
nand U10644 (N_10644,N_9679,N_8541);
nor U10645 (N_10645,N_9326,N_8680);
xor U10646 (N_10646,N_8048,N_8586);
xor U10647 (N_10647,N_9107,N_8121);
xor U10648 (N_10648,N_9030,N_8505);
nor U10649 (N_10649,N_9460,N_8185);
or U10650 (N_10650,N_8558,N_8217);
nor U10651 (N_10651,N_9268,N_8175);
nand U10652 (N_10652,N_9261,N_8369);
xnor U10653 (N_10653,N_8436,N_9749);
and U10654 (N_10654,N_8715,N_8063);
and U10655 (N_10655,N_8564,N_8972);
xor U10656 (N_10656,N_9751,N_8482);
xor U10657 (N_10657,N_9915,N_9558);
nor U10658 (N_10658,N_9730,N_9872);
xor U10659 (N_10659,N_8650,N_8849);
nor U10660 (N_10660,N_9540,N_8074);
or U10661 (N_10661,N_9678,N_8627);
nor U10662 (N_10662,N_8964,N_8226);
or U10663 (N_10663,N_8333,N_9341);
nor U10664 (N_10664,N_8336,N_8132);
nand U10665 (N_10665,N_9792,N_9790);
or U10666 (N_10666,N_9168,N_8638);
and U10667 (N_10667,N_9461,N_9759);
nand U10668 (N_10668,N_9893,N_8671);
nand U10669 (N_10669,N_9316,N_8141);
or U10670 (N_10670,N_8381,N_8233);
xnor U10671 (N_10671,N_8000,N_9600);
xnor U10672 (N_10672,N_9266,N_9931);
nand U10673 (N_10673,N_9664,N_8815);
xor U10674 (N_10674,N_8370,N_9647);
xnor U10675 (N_10675,N_9407,N_8504);
or U10676 (N_10676,N_9882,N_8741);
nand U10677 (N_10677,N_8923,N_8402);
or U10678 (N_10678,N_8724,N_9559);
xor U10679 (N_10679,N_9209,N_9245);
nand U10680 (N_10680,N_8782,N_9360);
and U10681 (N_10681,N_8778,N_8150);
and U10682 (N_10682,N_8476,N_8597);
and U10683 (N_10683,N_9081,N_9040);
and U10684 (N_10684,N_9487,N_9436);
xnor U10685 (N_10685,N_9736,N_8801);
xnor U10686 (N_10686,N_8997,N_8337);
xor U10687 (N_10687,N_8888,N_9833);
xor U10688 (N_10688,N_8338,N_9399);
and U10689 (N_10689,N_9542,N_8533);
and U10690 (N_10690,N_9452,N_9136);
and U10691 (N_10691,N_9665,N_9289);
and U10692 (N_10692,N_9352,N_9115);
nand U10693 (N_10693,N_9342,N_8495);
nand U10694 (N_10694,N_8894,N_8902);
nor U10695 (N_10695,N_9779,N_9344);
nor U10696 (N_10696,N_8913,N_8420);
or U10697 (N_10697,N_8099,N_9753);
nor U10698 (N_10698,N_8046,N_8605);
xnor U10699 (N_10699,N_8812,N_8624);
and U10700 (N_10700,N_9138,N_8569);
xnor U10701 (N_10701,N_8962,N_9936);
nand U10702 (N_10702,N_9312,N_9254);
nor U10703 (N_10703,N_8621,N_9448);
nand U10704 (N_10704,N_9776,N_8292);
or U10705 (N_10705,N_9337,N_9393);
or U10706 (N_10706,N_9695,N_8655);
and U10707 (N_10707,N_9398,N_8158);
nor U10708 (N_10708,N_8320,N_8626);
or U10709 (N_10709,N_9117,N_9036);
nand U10710 (N_10710,N_9726,N_9263);
nor U10711 (N_10711,N_8487,N_8373);
or U10712 (N_10712,N_8610,N_8693);
nor U10713 (N_10713,N_8945,N_9408);
xor U10714 (N_10714,N_9484,N_9305);
nor U10715 (N_10715,N_9958,N_9041);
or U10716 (N_10716,N_8748,N_8510);
nor U10717 (N_10717,N_9195,N_9469);
and U10718 (N_10718,N_9264,N_9338);
xnor U10719 (N_10719,N_9424,N_9526);
xnor U10720 (N_10720,N_9298,N_8478);
or U10721 (N_10721,N_9454,N_8981);
nor U10722 (N_10722,N_9938,N_9176);
and U10723 (N_10723,N_8010,N_8457);
and U10724 (N_10724,N_9043,N_8410);
or U10725 (N_10725,N_9230,N_9821);
or U10726 (N_10726,N_8071,N_8873);
or U10727 (N_10727,N_9165,N_8651);
nand U10728 (N_10728,N_8198,N_9652);
xor U10729 (N_10729,N_9737,N_8676);
and U10730 (N_10730,N_9777,N_9841);
or U10731 (N_10731,N_9728,N_9358);
nand U10732 (N_10732,N_9033,N_9097);
nor U10733 (N_10733,N_9667,N_8125);
nand U10734 (N_10734,N_9379,N_8204);
xor U10735 (N_10735,N_9904,N_8044);
xor U10736 (N_10736,N_8675,N_9489);
or U10737 (N_10737,N_8189,N_9654);
xnor U10738 (N_10738,N_8687,N_9912);
or U10739 (N_10739,N_9579,N_8664);
xnor U10740 (N_10740,N_8529,N_8214);
nor U10741 (N_10741,N_8269,N_9838);
xnor U10742 (N_10742,N_8004,N_9068);
nor U10743 (N_10743,N_8932,N_9946);
nand U10744 (N_10744,N_9733,N_8367);
xor U10745 (N_10745,N_8357,N_8511);
or U10746 (N_10746,N_9203,N_9417);
or U10747 (N_10747,N_8401,N_9953);
nor U10748 (N_10748,N_8996,N_8481);
or U10749 (N_10749,N_9405,N_8419);
nor U10750 (N_10750,N_8822,N_8523);
xor U10751 (N_10751,N_9956,N_8817);
or U10752 (N_10752,N_9474,N_8695);
or U10753 (N_10753,N_8149,N_8833);
nand U10754 (N_10754,N_9710,N_9616);
or U10755 (N_10755,N_8991,N_9815);
or U10756 (N_10756,N_8267,N_9034);
and U10757 (N_10757,N_9533,N_8584);
nor U10758 (N_10758,N_9445,N_9580);
xor U10759 (N_10759,N_9552,N_8296);
xnor U10760 (N_10760,N_8289,N_9177);
nor U10761 (N_10761,N_9688,N_8291);
nand U10762 (N_10762,N_9154,N_9967);
nand U10763 (N_10763,N_8636,N_8067);
xnor U10764 (N_10764,N_8360,N_9620);
nor U10765 (N_10765,N_8925,N_8052);
nand U10766 (N_10766,N_9982,N_9294);
or U10767 (N_10767,N_9387,N_8717);
nor U10768 (N_10768,N_9643,N_8663);
nand U10769 (N_10769,N_9103,N_9536);
nand U10770 (N_10770,N_8107,N_8188);
or U10771 (N_10771,N_8660,N_9455);
or U10772 (N_10772,N_9964,N_8824);
and U10773 (N_10773,N_9860,N_9354);
or U10774 (N_10774,N_9285,N_9215);
or U10775 (N_10775,N_9441,N_8500);
or U10776 (N_10776,N_9032,N_9323);
or U10777 (N_10777,N_8020,N_9650);
or U10778 (N_10778,N_9373,N_8813);
nor U10779 (N_10779,N_9409,N_9945);
xor U10780 (N_10780,N_8186,N_8789);
nor U10781 (N_10781,N_8134,N_8015);
nand U10782 (N_10782,N_8278,N_8643);
xor U10783 (N_10783,N_8377,N_9065);
or U10784 (N_10784,N_8209,N_8414);
or U10785 (N_10785,N_9990,N_9291);
xor U10786 (N_10786,N_8589,N_8632);
or U10787 (N_10787,N_9085,N_8102);
xor U10788 (N_10788,N_8231,N_9722);
nand U10789 (N_10789,N_8200,N_8021);
nand U10790 (N_10790,N_9108,N_8418);
nor U10791 (N_10791,N_8721,N_8126);
xnor U10792 (N_10792,N_9258,N_8339);
nor U10793 (N_10793,N_8520,N_9330);
or U10794 (N_10794,N_9934,N_8765);
nor U10795 (N_10795,N_8647,N_9698);
nand U10796 (N_10796,N_8509,N_9918);
or U10797 (N_10797,N_9013,N_8979);
and U10798 (N_10798,N_9775,N_9412);
and U10799 (N_10799,N_9121,N_9727);
nand U10800 (N_10800,N_8494,N_8549);
xnor U10801 (N_10801,N_8101,N_8684);
nor U10802 (N_10802,N_9803,N_9894);
or U10803 (N_10803,N_8416,N_8263);
or U10804 (N_10804,N_9836,N_8635);
and U10805 (N_10805,N_9490,N_8645);
xnor U10806 (N_10806,N_8312,N_9119);
xor U10807 (N_10807,N_8836,N_8901);
and U10808 (N_10808,N_9396,N_8918);
xor U10809 (N_10809,N_8629,N_9794);
nand U10810 (N_10810,N_8411,N_8580);
xnor U10811 (N_10811,N_8734,N_8503);
nor U10812 (N_10812,N_9829,N_8947);
or U10813 (N_10813,N_8594,N_8311);
nor U10814 (N_10814,N_9324,N_9865);
nor U10815 (N_10815,N_8760,N_9116);
nor U10816 (N_10816,N_8591,N_9642);
xor U10817 (N_10817,N_8857,N_9755);
xnor U10818 (N_10818,N_9287,N_9275);
nand U10819 (N_10819,N_8628,N_9618);
or U10820 (N_10820,N_9716,N_8691);
xor U10821 (N_10821,N_9731,N_9720);
nand U10822 (N_10822,N_9597,N_9778);
and U10823 (N_10823,N_8489,N_9842);
or U10824 (N_10824,N_9599,N_9256);
nand U10825 (N_10825,N_8435,N_8574);
or U10826 (N_10826,N_8111,N_9622);
or U10827 (N_10827,N_9696,N_8146);
nand U10828 (N_10828,N_8210,N_9649);
and U10829 (N_10829,N_9629,N_9118);
xor U10830 (N_10830,N_8055,N_9059);
nand U10831 (N_10831,N_9425,N_8038);
nor U10832 (N_10832,N_8625,N_9612);
or U10833 (N_10833,N_8080,N_9173);
nor U10834 (N_10834,N_9233,N_9340);
nand U10835 (N_10835,N_9538,N_8224);
and U10836 (N_10836,N_9648,N_9963);
xor U10837 (N_10837,N_8842,N_8486);
or U10838 (N_10838,N_8527,N_9422);
xnor U10839 (N_10839,N_8039,N_8864);
nand U10840 (N_10840,N_9056,N_9385);
or U10841 (N_10841,N_8553,N_8978);
or U10842 (N_10842,N_9131,N_9488);
nor U10843 (N_10843,N_8560,N_9576);
and U10844 (N_10844,N_9313,N_8685);
nand U10845 (N_10845,N_8073,N_9633);
and U10846 (N_10846,N_9689,N_8417);
xnor U10847 (N_10847,N_8220,N_9700);
xor U10848 (N_10848,N_9498,N_9655);
xnor U10849 (N_10849,N_8281,N_8555);
xnor U10850 (N_10850,N_9411,N_9061);
nand U10851 (N_10851,N_9739,N_8007);
xor U10852 (N_10852,N_8762,N_9791);
nand U10853 (N_10853,N_9496,N_8471);
nand U10854 (N_10854,N_8174,N_8100);
nand U10855 (N_10855,N_9921,N_8378);
nand U10856 (N_10856,N_9911,N_8808);
nor U10857 (N_10857,N_8703,N_8977);
xnor U10858 (N_10858,N_9429,N_8032);
and U10859 (N_10859,N_8544,N_9547);
and U10860 (N_10860,N_9388,N_9604);
xor U10861 (N_10861,N_9410,N_8848);
nand U10862 (N_10862,N_9348,N_8853);
or U10863 (N_10863,N_8153,N_9919);
nor U10864 (N_10864,N_9627,N_8374);
xnor U10865 (N_10865,N_8270,N_8042);
nor U10866 (N_10866,N_9944,N_9914);
nand U10867 (N_10867,N_8794,N_9415);
nand U10868 (N_10868,N_8302,N_9467);
and U10869 (N_10869,N_8310,N_9782);
nand U10870 (N_10870,N_8579,N_8648);
xnor U10871 (N_10871,N_8653,N_9565);
xor U10872 (N_10872,N_9743,N_9623);
and U10873 (N_10873,N_8998,N_8258);
nand U10874 (N_10874,N_8447,N_8513);
and U10875 (N_10875,N_8066,N_8024);
nor U10876 (N_10876,N_9721,N_8282);
nor U10877 (N_10877,N_9995,N_8382);
nand U10878 (N_10878,N_9058,N_8492);
and U10879 (N_10879,N_9977,N_8238);
and U10880 (N_10880,N_8929,N_8437);
nand U10881 (N_10881,N_8388,N_8872);
and U10882 (N_10882,N_8456,N_9506);
nor U10883 (N_10883,N_8880,N_9297);
or U10884 (N_10884,N_8766,N_8818);
and U10885 (N_10885,N_9740,N_8236);
nand U10886 (N_10886,N_8203,N_9670);
nor U10887 (N_10887,N_8193,N_9376);
and U10888 (N_10888,N_8182,N_9152);
and U10889 (N_10889,N_8244,N_8082);
and U10890 (N_10890,N_9044,N_9446);
and U10891 (N_10891,N_9054,N_8318);
xnor U10892 (N_10892,N_9100,N_8847);
and U10893 (N_10893,N_9840,N_9682);
nor U10894 (N_10894,N_9156,N_9691);
and U10895 (N_10895,N_8043,N_9762);
xnor U10896 (N_10896,N_9908,N_9182);
nor U10897 (N_10897,N_9027,N_8396);
or U10898 (N_10898,N_8750,N_8862);
nand U10899 (N_10899,N_9321,N_8819);
nor U10900 (N_10900,N_9320,N_8187);
nor U10901 (N_10901,N_9394,N_8179);
and U10902 (N_10902,N_8245,N_9278);
nor U10903 (N_10903,N_8572,N_8394);
and U10904 (N_10904,N_9249,N_8364);
nor U10905 (N_10905,N_9042,N_8599);
and U10906 (N_10906,N_9859,N_8770);
and U10907 (N_10907,N_9072,N_8240);
nand U10908 (N_10908,N_8759,N_8940);
and U10909 (N_10909,N_8743,N_9317);
and U10910 (N_10910,N_8212,N_9603);
nor U10911 (N_10911,N_9048,N_9292);
nor U10912 (N_10912,N_9071,N_9527);
and U10913 (N_10913,N_8522,N_8279);
nand U10914 (N_10914,N_9524,N_8499);
xor U10915 (N_10915,N_9693,N_9381);
nand U10916 (N_10916,N_9435,N_8835);
nand U10917 (N_10917,N_8450,N_8829);
nor U10918 (N_10918,N_8341,N_9011);
and U10919 (N_10919,N_9453,N_9884);
xnor U10920 (N_10920,N_9820,N_8119);
or U10921 (N_10921,N_8568,N_9973);
or U10922 (N_10922,N_9927,N_9111);
xnor U10923 (N_10923,N_8324,N_9709);
nor U10924 (N_10924,N_9153,N_8899);
or U10925 (N_10925,N_8518,N_8256);
or U10926 (N_10926,N_9143,N_9470);
or U10927 (N_10927,N_9012,N_9327);
or U10928 (N_10928,N_9994,N_8776);
nor U10929 (N_10929,N_9259,N_8668);
nand U10930 (N_10930,N_8458,N_9874);
nand U10931 (N_10931,N_9834,N_8756);
or U10932 (N_10932,N_8496,N_8398);
nor U10933 (N_10933,N_9001,N_9879);
nand U10934 (N_10934,N_8202,N_9630);
or U10935 (N_10935,N_8525,N_9509);
nor U10936 (N_10936,N_9702,N_9869);
nand U10937 (N_10937,N_8103,N_8424);
nand U10938 (N_10938,N_8058,N_8285);
nor U10939 (N_10939,N_9961,N_8949);
xor U10940 (N_10940,N_9766,N_9661);
or U10941 (N_10941,N_8874,N_8806);
nand U10942 (N_10942,N_8809,N_8271);
nor U10943 (N_10943,N_9128,N_9022);
xnor U10944 (N_10944,N_9950,N_9161);
nand U10945 (N_10945,N_9050,N_9659);
or U10946 (N_10946,N_8729,N_8955);
nor U10947 (N_10947,N_8514,N_8611);
nand U10948 (N_10948,N_9539,N_9856);
or U10949 (N_10949,N_9493,N_9541);
nor U10950 (N_10950,N_8343,N_8823);
or U10951 (N_10951,N_8466,N_9380);
or U10952 (N_10952,N_8051,N_8181);
or U10953 (N_10953,N_9475,N_8708);
nor U10954 (N_10954,N_8543,N_8810);
xor U10955 (N_10955,N_8565,N_8237);
nor U10956 (N_10956,N_9621,N_8562);
xnor U10957 (N_10957,N_8590,N_9296);
and U10958 (N_10958,N_8088,N_9369);
and U10959 (N_10959,N_9502,N_8799);
nand U10960 (N_10960,N_8331,N_8618);
nand U10961 (N_10961,N_9122,N_8314);
nor U10962 (N_10962,N_9588,N_9906);
or U10963 (N_10963,N_8984,N_9096);
nor U10964 (N_10964,N_8056,N_8440);
nand U10965 (N_10965,N_8926,N_9265);
or U10966 (N_10966,N_9336,N_9534);
nand U10967 (N_10967,N_9993,N_8049);
and U10968 (N_10968,N_9151,N_8356);
nor U10969 (N_10969,N_9125,N_9850);
or U10970 (N_10970,N_8540,N_8114);
xnor U10971 (N_10971,N_9653,N_8825);
nor U10972 (N_10972,N_9255,N_9437);
and U10973 (N_10973,N_9809,N_9635);
xor U10974 (N_10974,N_8791,N_9083);
or U10975 (N_10975,N_9084,N_8667);
or U10976 (N_10976,N_8350,N_9247);
and U10977 (N_10977,N_9863,N_9917);
or U10978 (N_10978,N_8786,N_9715);
nor U10979 (N_10979,N_8035,N_9210);
nand U10980 (N_10980,N_9907,N_8385);
xnor U10981 (N_10981,N_9972,N_8462);
nand U10982 (N_10982,N_9774,N_9479);
nand U10983 (N_10983,N_8740,N_8441);
xnor U10984 (N_10984,N_8081,N_8834);
xnor U10985 (N_10985,N_8483,N_8933);
nor U10986 (N_10986,N_8380,N_9607);
and U10987 (N_10987,N_9560,N_9997);
xor U10988 (N_10988,N_8706,N_8583);
nor U10989 (N_10989,N_8846,N_8235);
nor U10990 (N_10990,N_9692,N_8903);
nor U10991 (N_10991,N_9837,N_8920);
nand U10992 (N_10992,N_9701,N_8330);
nand U10993 (N_10993,N_8243,N_8749);
xor U10994 (N_10994,N_9985,N_9587);
xnor U10995 (N_10995,N_9120,N_8300);
xnor U10996 (N_10996,N_9830,N_9846);
xor U10997 (N_10997,N_9989,N_8723);
nor U10998 (N_10998,N_9754,N_9955);
and U10999 (N_10999,N_8439,N_9191);
xor U11000 (N_11000,N_9186,N_9431);
xor U11001 (N_11001,N_9405,N_9571);
nand U11002 (N_11002,N_9307,N_9824);
xor U11003 (N_11003,N_9895,N_9463);
nand U11004 (N_11004,N_9725,N_8755);
and U11005 (N_11005,N_8121,N_8639);
nor U11006 (N_11006,N_8317,N_9825);
nand U11007 (N_11007,N_8717,N_9343);
nor U11008 (N_11008,N_8677,N_9125);
nand U11009 (N_11009,N_8682,N_8951);
xor U11010 (N_11010,N_8895,N_8328);
nand U11011 (N_11011,N_9121,N_8384);
nand U11012 (N_11012,N_8463,N_9548);
nand U11013 (N_11013,N_8123,N_8032);
and U11014 (N_11014,N_9927,N_9035);
xor U11015 (N_11015,N_8939,N_8308);
xnor U11016 (N_11016,N_9989,N_8768);
or U11017 (N_11017,N_8679,N_8178);
or U11018 (N_11018,N_8287,N_9202);
xnor U11019 (N_11019,N_8452,N_8051);
or U11020 (N_11020,N_8398,N_8631);
xor U11021 (N_11021,N_9309,N_9536);
and U11022 (N_11022,N_8123,N_8241);
nand U11023 (N_11023,N_8888,N_9627);
nand U11024 (N_11024,N_8687,N_9466);
xnor U11025 (N_11025,N_9928,N_9541);
and U11026 (N_11026,N_9730,N_9114);
or U11027 (N_11027,N_9963,N_8664);
or U11028 (N_11028,N_9236,N_9131);
nor U11029 (N_11029,N_8203,N_9709);
nand U11030 (N_11030,N_8963,N_8373);
xnor U11031 (N_11031,N_8871,N_8809);
or U11032 (N_11032,N_9978,N_8129);
nand U11033 (N_11033,N_8514,N_8344);
and U11034 (N_11034,N_9100,N_8351);
nand U11035 (N_11035,N_8263,N_8288);
or U11036 (N_11036,N_8305,N_8711);
xor U11037 (N_11037,N_9750,N_8465);
nand U11038 (N_11038,N_9505,N_8518);
nand U11039 (N_11039,N_9101,N_9447);
nand U11040 (N_11040,N_8699,N_9723);
nand U11041 (N_11041,N_8216,N_8716);
nand U11042 (N_11042,N_8355,N_8164);
nor U11043 (N_11043,N_8170,N_8793);
or U11044 (N_11044,N_9316,N_9149);
nand U11045 (N_11045,N_8443,N_8414);
or U11046 (N_11046,N_9260,N_8822);
or U11047 (N_11047,N_8461,N_8107);
and U11048 (N_11048,N_9003,N_8549);
xnor U11049 (N_11049,N_9935,N_9937);
or U11050 (N_11050,N_9097,N_9579);
nand U11051 (N_11051,N_9384,N_9227);
and U11052 (N_11052,N_8127,N_9232);
xor U11053 (N_11053,N_8405,N_8705);
nand U11054 (N_11054,N_8267,N_9816);
nor U11055 (N_11055,N_9656,N_8935);
or U11056 (N_11056,N_8108,N_9246);
or U11057 (N_11057,N_9875,N_9155);
nor U11058 (N_11058,N_9447,N_8210);
or U11059 (N_11059,N_9910,N_9114);
and U11060 (N_11060,N_8128,N_9046);
xnor U11061 (N_11061,N_9645,N_9273);
and U11062 (N_11062,N_9915,N_8395);
xnor U11063 (N_11063,N_9196,N_8443);
and U11064 (N_11064,N_8327,N_9501);
and U11065 (N_11065,N_9881,N_8548);
nor U11066 (N_11066,N_9749,N_8713);
nor U11067 (N_11067,N_9914,N_8313);
nand U11068 (N_11068,N_8380,N_8180);
xor U11069 (N_11069,N_9827,N_9322);
xnor U11070 (N_11070,N_8410,N_9278);
xnor U11071 (N_11071,N_9773,N_9994);
nor U11072 (N_11072,N_9997,N_9656);
nand U11073 (N_11073,N_8399,N_9382);
or U11074 (N_11074,N_9209,N_9105);
and U11075 (N_11075,N_9772,N_8883);
and U11076 (N_11076,N_9399,N_8816);
nor U11077 (N_11077,N_9412,N_9720);
nor U11078 (N_11078,N_9176,N_9866);
or U11079 (N_11079,N_8172,N_8009);
or U11080 (N_11080,N_9898,N_9222);
nand U11081 (N_11081,N_8842,N_9639);
or U11082 (N_11082,N_9744,N_9838);
nand U11083 (N_11083,N_8459,N_9031);
xnor U11084 (N_11084,N_9257,N_8170);
nor U11085 (N_11085,N_9726,N_9955);
nor U11086 (N_11086,N_9383,N_8398);
and U11087 (N_11087,N_8061,N_8043);
and U11088 (N_11088,N_8271,N_8780);
xnor U11089 (N_11089,N_9589,N_9711);
or U11090 (N_11090,N_8047,N_9604);
and U11091 (N_11091,N_8896,N_9019);
or U11092 (N_11092,N_8501,N_9219);
nand U11093 (N_11093,N_9385,N_9561);
nand U11094 (N_11094,N_9329,N_8083);
xor U11095 (N_11095,N_9913,N_8431);
nand U11096 (N_11096,N_8994,N_9894);
or U11097 (N_11097,N_8639,N_9033);
and U11098 (N_11098,N_9175,N_9240);
and U11099 (N_11099,N_9038,N_9339);
or U11100 (N_11100,N_8572,N_8733);
xnor U11101 (N_11101,N_9865,N_8608);
or U11102 (N_11102,N_9072,N_8896);
nor U11103 (N_11103,N_8407,N_8517);
or U11104 (N_11104,N_9002,N_8044);
xor U11105 (N_11105,N_8599,N_9321);
or U11106 (N_11106,N_9420,N_9286);
or U11107 (N_11107,N_9120,N_9986);
nor U11108 (N_11108,N_9506,N_9371);
nand U11109 (N_11109,N_8218,N_9261);
or U11110 (N_11110,N_9226,N_9260);
nor U11111 (N_11111,N_9766,N_8252);
nand U11112 (N_11112,N_8205,N_8738);
nand U11113 (N_11113,N_8459,N_9860);
and U11114 (N_11114,N_9535,N_8060);
nor U11115 (N_11115,N_8175,N_8728);
nor U11116 (N_11116,N_9367,N_9715);
xnor U11117 (N_11117,N_8086,N_8999);
nand U11118 (N_11118,N_8635,N_9521);
xnor U11119 (N_11119,N_8544,N_9934);
or U11120 (N_11120,N_8264,N_8696);
or U11121 (N_11121,N_9294,N_9231);
nand U11122 (N_11122,N_8306,N_8033);
xnor U11123 (N_11123,N_8863,N_8210);
nor U11124 (N_11124,N_8480,N_8890);
nand U11125 (N_11125,N_9992,N_9981);
nor U11126 (N_11126,N_9913,N_9400);
nand U11127 (N_11127,N_9947,N_8427);
or U11128 (N_11128,N_9637,N_9043);
nor U11129 (N_11129,N_8134,N_8527);
and U11130 (N_11130,N_8618,N_8697);
nand U11131 (N_11131,N_9449,N_8970);
nor U11132 (N_11132,N_8060,N_8151);
xnor U11133 (N_11133,N_9836,N_8619);
xor U11134 (N_11134,N_9119,N_8578);
nor U11135 (N_11135,N_9244,N_8008);
or U11136 (N_11136,N_9415,N_9999);
nand U11137 (N_11137,N_8650,N_9298);
and U11138 (N_11138,N_8473,N_9756);
or U11139 (N_11139,N_8713,N_8652);
nand U11140 (N_11140,N_9707,N_8342);
nor U11141 (N_11141,N_8558,N_8481);
and U11142 (N_11142,N_9482,N_8945);
or U11143 (N_11143,N_8931,N_9439);
or U11144 (N_11144,N_8608,N_8129);
xor U11145 (N_11145,N_9062,N_9359);
nand U11146 (N_11146,N_8282,N_9964);
or U11147 (N_11147,N_8165,N_8443);
or U11148 (N_11148,N_9127,N_8203);
nand U11149 (N_11149,N_8435,N_9766);
xnor U11150 (N_11150,N_8256,N_9382);
nand U11151 (N_11151,N_9447,N_9634);
nor U11152 (N_11152,N_8675,N_8184);
or U11153 (N_11153,N_9538,N_9636);
and U11154 (N_11154,N_8653,N_8503);
and U11155 (N_11155,N_8111,N_9874);
or U11156 (N_11156,N_8691,N_9057);
nor U11157 (N_11157,N_9949,N_8272);
or U11158 (N_11158,N_8224,N_9905);
xnor U11159 (N_11159,N_8422,N_9451);
and U11160 (N_11160,N_8122,N_8422);
or U11161 (N_11161,N_8762,N_9377);
xor U11162 (N_11162,N_9990,N_9845);
nand U11163 (N_11163,N_8172,N_8557);
and U11164 (N_11164,N_8251,N_8693);
nor U11165 (N_11165,N_8362,N_8517);
xor U11166 (N_11166,N_8054,N_8375);
nand U11167 (N_11167,N_8592,N_8959);
and U11168 (N_11168,N_8579,N_9724);
or U11169 (N_11169,N_8767,N_8136);
nand U11170 (N_11170,N_8172,N_9955);
nor U11171 (N_11171,N_9063,N_9457);
nand U11172 (N_11172,N_9392,N_9578);
xor U11173 (N_11173,N_9969,N_9760);
nor U11174 (N_11174,N_9343,N_8223);
nand U11175 (N_11175,N_8808,N_9087);
nor U11176 (N_11176,N_8310,N_9314);
nor U11177 (N_11177,N_9432,N_9059);
nand U11178 (N_11178,N_8540,N_9740);
or U11179 (N_11179,N_9709,N_8299);
or U11180 (N_11180,N_8468,N_8583);
and U11181 (N_11181,N_9736,N_8066);
xnor U11182 (N_11182,N_8750,N_8487);
and U11183 (N_11183,N_9177,N_9946);
nand U11184 (N_11184,N_9587,N_9497);
or U11185 (N_11185,N_8230,N_9354);
nor U11186 (N_11186,N_8892,N_9161);
nor U11187 (N_11187,N_9239,N_9705);
nand U11188 (N_11188,N_9397,N_9287);
or U11189 (N_11189,N_9348,N_8851);
or U11190 (N_11190,N_9284,N_8467);
xnor U11191 (N_11191,N_9308,N_8047);
xor U11192 (N_11192,N_8218,N_9455);
or U11193 (N_11193,N_9697,N_9372);
nand U11194 (N_11194,N_9510,N_9004);
and U11195 (N_11195,N_9510,N_8143);
nor U11196 (N_11196,N_9250,N_8083);
nand U11197 (N_11197,N_9849,N_8829);
nand U11198 (N_11198,N_9877,N_9823);
xnor U11199 (N_11199,N_8556,N_9168);
and U11200 (N_11200,N_9105,N_8660);
xnor U11201 (N_11201,N_8486,N_9310);
and U11202 (N_11202,N_9041,N_8678);
nor U11203 (N_11203,N_9467,N_9724);
or U11204 (N_11204,N_9675,N_9253);
or U11205 (N_11205,N_8752,N_9417);
nor U11206 (N_11206,N_9900,N_8560);
or U11207 (N_11207,N_8866,N_9015);
xor U11208 (N_11208,N_9525,N_8219);
xor U11209 (N_11209,N_8355,N_8529);
and U11210 (N_11210,N_9258,N_8553);
nand U11211 (N_11211,N_9481,N_9334);
xor U11212 (N_11212,N_9237,N_9305);
nor U11213 (N_11213,N_9986,N_8551);
and U11214 (N_11214,N_9238,N_8792);
and U11215 (N_11215,N_9134,N_8628);
and U11216 (N_11216,N_8347,N_9932);
and U11217 (N_11217,N_8995,N_8108);
nand U11218 (N_11218,N_8664,N_9595);
nand U11219 (N_11219,N_9324,N_9913);
nand U11220 (N_11220,N_8806,N_8020);
xnor U11221 (N_11221,N_8172,N_9560);
nor U11222 (N_11222,N_9609,N_8290);
nor U11223 (N_11223,N_8219,N_8856);
nor U11224 (N_11224,N_8447,N_9139);
nand U11225 (N_11225,N_9574,N_8474);
and U11226 (N_11226,N_8962,N_8718);
or U11227 (N_11227,N_8876,N_8980);
and U11228 (N_11228,N_9465,N_8911);
nor U11229 (N_11229,N_9091,N_8401);
and U11230 (N_11230,N_8037,N_9519);
and U11231 (N_11231,N_9019,N_8021);
and U11232 (N_11232,N_8719,N_9987);
xnor U11233 (N_11233,N_8792,N_9614);
nor U11234 (N_11234,N_8476,N_8966);
and U11235 (N_11235,N_9416,N_9844);
nand U11236 (N_11236,N_9824,N_8770);
nor U11237 (N_11237,N_9820,N_9051);
xnor U11238 (N_11238,N_8951,N_9687);
nand U11239 (N_11239,N_9985,N_9357);
and U11240 (N_11240,N_9907,N_8169);
xor U11241 (N_11241,N_9713,N_9618);
and U11242 (N_11242,N_9903,N_8679);
or U11243 (N_11243,N_8198,N_9782);
or U11244 (N_11244,N_9835,N_9884);
nor U11245 (N_11245,N_9338,N_8412);
nand U11246 (N_11246,N_9600,N_8737);
nand U11247 (N_11247,N_8103,N_8429);
and U11248 (N_11248,N_9116,N_9046);
and U11249 (N_11249,N_9676,N_8985);
xnor U11250 (N_11250,N_9573,N_8784);
nand U11251 (N_11251,N_9172,N_9900);
nor U11252 (N_11252,N_8729,N_9257);
nor U11253 (N_11253,N_8310,N_9138);
xnor U11254 (N_11254,N_9516,N_9943);
nor U11255 (N_11255,N_8804,N_8089);
nor U11256 (N_11256,N_8454,N_9393);
and U11257 (N_11257,N_8803,N_9773);
xnor U11258 (N_11258,N_8473,N_8708);
or U11259 (N_11259,N_9167,N_8146);
or U11260 (N_11260,N_8502,N_9473);
nor U11261 (N_11261,N_9765,N_8609);
xnor U11262 (N_11262,N_8925,N_8320);
xor U11263 (N_11263,N_9623,N_8481);
nand U11264 (N_11264,N_8307,N_9291);
and U11265 (N_11265,N_9362,N_9589);
nand U11266 (N_11266,N_8423,N_9080);
nor U11267 (N_11267,N_9039,N_8614);
xor U11268 (N_11268,N_9438,N_9256);
and U11269 (N_11269,N_9634,N_9769);
nand U11270 (N_11270,N_8783,N_8595);
or U11271 (N_11271,N_8688,N_8764);
xor U11272 (N_11272,N_8254,N_8170);
nand U11273 (N_11273,N_9391,N_8075);
or U11274 (N_11274,N_9867,N_8443);
nand U11275 (N_11275,N_9716,N_9060);
xnor U11276 (N_11276,N_9542,N_8943);
nor U11277 (N_11277,N_8482,N_8979);
xor U11278 (N_11278,N_8370,N_8591);
or U11279 (N_11279,N_8289,N_9000);
nand U11280 (N_11280,N_8145,N_9621);
nand U11281 (N_11281,N_9976,N_9362);
or U11282 (N_11282,N_8123,N_9975);
or U11283 (N_11283,N_9914,N_8008);
xor U11284 (N_11284,N_9595,N_9052);
or U11285 (N_11285,N_9148,N_9429);
nand U11286 (N_11286,N_8432,N_9469);
or U11287 (N_11287,N_9398,N_8165);
nand U11288 (N_11288,N_9214,N_9001);
nor U11289 (N_11289,N_9458,N_9586);
nand U11290 (N_11290,N_9027,N_9487);
nand U11291 (N_11291,N_9960,N_9918);
and U11292 (N_11292,N_9617,N_8160);
and U11293 (N_11293,N_8278,N_8822);
nand U11294 (N_11294,N_8874,N_8152);
nand U11295 (N_11295,N_8992,N_8456);
nor U11296 (N_11296,N_8096,N_8074);
nor U11297 (N_11297,N_8990,N_8247);
nor U11298 (N_11298,N_8791,N_8189);
nand U11299 (N_11299,N_9743,N_8981);
or U11300 (N_11300,N_8935,N_9536);
nor U11301 (N_11301,N_8689,N_8367);
xor U11302 (N_11302,N_9292,N_8913);
xor U11303 (N_11303,N_9630,N_9645);
or U11304 (N_11304,N_9439,N_8290);
xor U11305 (N_11305,N_8364,N_9422);
nor U11306 (N_11306,N_9416,N_9900);
or U11307 (N_11307,N_8770,N_9469);
nor U11308 (N_11308,N_9868,N_9963);
xor U11309 (N_11309,N_8081,N_9390);
or U11310 (N_11310,N_9761,N_8323);
nor U11311 (N_11311,N_8774,N_8955);
xor U11312 (N_11312,N_8944,N_8238);
xnor U11313 (N_11313,N_9140,N_9646);
and U11314 (N_11314,N_9132,N_8298);
nor U11315 (N_11315,N_8644,N_9614);
nand U11316 (N_11316,N_9077,N_8030);
nor U11317 (N_11317,N_9591,N_8898);
nor U11318 (N_11318,N_8805,N_8167);
and U11319 (N_11319,N_9962,N_8984);
and U11320 (N_11320,N_9495,N_8259);
or U11321 (N_11321,N_9253,N_9047);
nand U11322 (N_11322,N_8980,N_8047);
nand U11323 (N_11323,N_8191,N_9343);
xnor U11324 (N_11324,N_9293,N_9796);
or U11325 (N_11325,N_9480,N_8324);
nor U11326 (N_11326,N_8900,N_9508);
nor U11327 (N_11327,N_9965,N_8859);
xnor U11328 (N_11328,N_9601,N_9949);
nor U11329 (N_11329,N_8686,N_8758);
nand U11330 (N_11330,N_9144,N_9788);
nand U11331 (N_11331,N_9040,N_8475);
xnor U11332 (N_11332,N_8708,N_8418);
nor U11333 (N_11333,N_8919,N_9873);
xnor U11334 (N_11334,N_8354,N_8447);
or U11335 (N_11335,N_9268,N_8104);
or U11336 (N_11336,N_9543,N_8087);
nor U11337 (N_11337,N_9506,N_9760);
nand U11338 (N_11338,N_9951,N_8760);
nor U11339 (N_11339,N_9269,N_8724);
nand U11340 (N_11340,N_9706,N_8306);
nor U11341 (N_11341,N_8235,N_9674);
nor U11342 (N_11342,N_8148,N_9947);
nand U11343 (N_11343,N_8911,N_9687);
and U11344 (N_11344,N_9749,N_8399);
nor U11345 (N_11345,N_8933,N_8371);
xor U11346 (N_11346,N_9501,N_9854);
nand U11347 (N_11347,N_9662,N_8555);
xor U11348 (N_11348,N_9820,N_9093);
xnor U11349 (N_11349,N_9047,N_8065);
nand U11350 (N_11350,N_8587,N_8214);
nand U11351 (N_11351,N_8641,N_8692);
xnor U11352 (N_11352,N_8385,N_9885);
nor U11353 (N_11353,N_8836,N_9712);
nor U11354 (N_11354,N_9018,N_9752);
nor U11355 (N_11355,N_8187,N_9705);
xnor U11356 (N_11356,N_9125,N_8286);
nand U11357 (N_11357,N_9843,N_8749);
nand U11358 (N_11358,N_9997,N_8129);
xor U11359 (N_11359,N_9114,N_9277);
nor U11360 (N_11360,N_9681,N_8763);
nor U11361 (N_11361,N_9944,N_9274);
xnor U11362 (N_11362,N_9764,N_8311);
nand U11363 (N_11363,N_8213,N_8803);
xnor U11364 (N_11364,N_9008,N_9145);
or U11365 (N_11365,N_9425,N_8948);
and U11366 (N_11366,N_8668,N_8756);
xnor U11367 (N_11367,N_9609,N_9453);
or U11368 (N_11368,N_9224,N_8231);
or U11369 (N_11369,N_8335,N_8421);
nand U11370 (N_11370,N_9794,N_8124);
nor U11371 (N_11371,N_9456,N_9383);
or U11372 (N_11372,N_9906,N_8339);
and U11373 (N_11373,N_8801,N_9303);
nor U11374 (N_11374,N_8171,N_8153);
or U11375 (N_11375,N_8517,N_8066);
and U11376 (N_11376,N_8154,N_9371);
nand U11377 (N_11377,N_9755,N_8540);
or U11378 (N_11378,N_9587,N_9789);
xnor U11379 (N_11379,N_8639,N_9498);
nor U11380 (N_11380,N_9789,N_9365);
xnor U11381 (N_11381,N_9498,N_9601);
or U11382 (N_11382,N_8637,N_9185);
or U11383 (N_11383,N_9960,N_8294);
xor U11384 (N_11384,N_8321,N_8009);
nand U11385 (N_11385,N_9028,N_9132);
xor U11386 (N_11386,N_8992,N_8752);
or U11387 (N_11387,N_8520,N_9474);
and U11388 (N_11388,N_8962,N_8434);
and U11389 (N_11389,N_8064,N_9891);
or U11390 (N_11390,N_9662,N_8758);
xor U11391 (N_11391,N_9561,N_8489);
nor U11392 (N_11392,N_8661,N_8388);
or U11393 (N_11393,N_8500,N_9778);
xnor U11394 (N_11394,N_8437,N_8858);
xor U11395 (N_11395,N_8267,N_9432);
nor U11396 (N_11396,N_8276,N_9688);
and U11397 (N_11397,N_8690,N_9910);
nand U11398 (N_11398,N_8390,N_9218);
and U11399 (N_11399,N_8409,N_9308);
nand U11400 (N_11400,N_9212,N_9563);
and U11401 (N_11401,N_8375,N_8022);
nor U11402 (N_11402,N_8221,N_8016);
and U11403 (N_11403,N_9160,N_9577);
or U11404 (N_11404,N_8761,N_9370);
nor U11405 (N_11405,N_8481,N_9789);
nand U11406 (N_11406,N_9037,N_9276);
xnor U11407 (N_11407,N_9241,N_8562);
nand U11408 (N_11408,N_9124,N_8515);
and U11409 (N_11409,N_9998,N_8438);
xnor U11410 (N_11410,N_8034,N_8090);
xor U11411 (N_11411,N_9319,N_8082);
and U11412 (N_11412,N_9048,N_8196);
or U11413 (N_11413,N_8236,N_9359);
nand U11414 (N_11414,N_9463,N_9960);
nor U11415 (N_11415,N_8777,N_8034);
or U11416 (N_11416,N_8748,N_9076);
or U11417 (N_11417,N_9748,N_8795);
nand U11418 (N_11418,N_9240,N_8982);
nand U11419 (N_11419,N_9950,N_9724);
and U11420 (N_11420,N_9398,N_9093);
xnor U11421 (N_11421,N_9694,N_8863);
nand U11422 (N_11422,N_8399,N_8060);
nor U11423 (N_11423,N_9030,N_8240);
and U11424 (N_11424,N_8579,N_8554);
nand U11425 (N_11425,N_8345,N_8115);
or U11426 (N_11426,N_8738,N_8511);
nand U11427 (N_11427,N_8273,N_9739);
and U11428 (N_11428,N_8255,N_9172);
and U11429 (N_11429,N_9125,N_9370);
nand U11430 (N_11430,N_8301,N_8053);
and U11431 (N_11431,N_8492,N_8133);
nor U11432 (N_11432,N_8466,N_9226);
nand U11433 (N_11433,N_8789,N_9674);
nor U11434 (N_11434,N_8182,N_9951);
nand U11435 (N_11435,N_8896,N_8784);
nand U11436 (N_11436,N_8662,N_8119);
xnor U11437 (N_11437,N_8540,N_9142);
or U11438 (N_11438,N_8522,N_9827);
and U11439 (N_11439,N_9671,N_9224);
xor U11440 (N_11440,N_8197,N_9679);
or U11441 (N_11441,N_8158,N_9919);
nand U11442 (N_11442,N_8454,N_8825);
xnor U11443 (N_11443,N_8427,N_9889);
xnor U11444 (N_11444,N_8721,N_8482);
nor U11445 (N_11445,N_8098,N_9635);
and U11446 (N_11446,N_9137,N_8263);
and U11447 (N_11447,N_8144,N_8516);
or U11448 (N_11448,N_8262,N_9906);
nand U11449 (N_11449,N_9832,N_8031);
nor U11450 (N_11450,N_8191,N_8720);
and U11451 (N_11451,N_8732,N_8686);
or U11452 (N_11452,N_8685,N_8762);
nor U11453 (N_11453,N_8858,N_8726);
nor U11454 (N_11454,N_8357,N_9670);
or U11455 (N_11455,N_8325,N_8150);
and U11456 (N_11456,N_8345,N_9742);
nand U11457 (N_11457,N_8229,N_9806);
and U11458 (N_11458,N_8652,N_9144);
nand U11459 (N_11459,N_9313,N_9548);
nand U11460 (N_11460,N_8021,N_9525);
and U11461 (N_11461,N_8031,N_9091);
nor U11462 (N_11462,N_8469,N_9135);
xnor U11463 (N_11463,N_9636,N_9630);
nor U11464 (N_11464,N_8984,N_8370);
xnor U11465 (N_11465,N_9163,N_8711);
and U11466 (N_11466,N_8368,N_9432);
or U11467 (N_11467,N_8151,N_9565);
or U11468 (N_11468,N_8530,N_8065);
nor U11469 (N_11469,N_8602,N_9234);
nor U11470 (N_11470,N_9915,N_9266);
nand U11471 (N_11471,N_8315,N_8190);
nor U11472 (N_11472,N_9798,N_9452);
or U11473 (N_11473,N_9269,N_8234);
nand U11474 (N_11474,N_8905,N_9823);
nor U11475 (N_11475,N_8199,N_8105);
nor U11476 (N_11476,N_8150,N_9560);
nor U11477 (N_11477,N_9755,N_9503);
or U11478 (N_11478,N_8375,N_8087);
nand U11479 (N_11479,N_9220,N_8425);
or U11480 (N_11480,N_8483,N_8580);
and U11481 (N_11481,N_8161,N_9546);
xnor U11482 (N_11482,N_8314,N_9014);
and U11483 (N_11483,N_8221,N_9789);
nand U11484 (N_11484,N_9797,N_8941);
xnor U11485 (N_11485,N_9050,N_9666);
nand U11486 (N_11486,N_9119,N_9209);
nand U11487 (N_11487,N_9963,N_9216);
xnor U11488 (N_11488,N_9769,N_8841);
nor U11489 (N_11489,N_8788,N_9026);
xnor U11490 (N_11490,N_9982,N_9675);
or U11491 (N_11491,N_8843,N_9556);
xor U11492 (N_11492,N_9000,N_8529);
xnor U11493 (N_11493,N_9029,N_8420);
or U11494 (N_11494,N_9749,N_8183);
nand U11495 (N_11495,N_8522,N_9861);
nand U11496 (N_11496,N_8152,N_9977);
and U11497 (N_11497,N_9083,N_8146);
and U11498 (N_11498,N_9104,N_8066);
nor U11499 (N_11499,N_8999,N_8071);
xnor U11500 (N_11500,N_9709,N_8689);
and U11501 (N_11501,N_9633,N_8592);
nand U11502 (N_11502,N_9252,N_9095);
nand U11503 (N_11503,N_8580,N_9971);
nand U11504 (N_11504,N_9732,N_9968);
and U11505 (N_11505,N_8648,N_8652);
xor U11506 (N_11506,N_8066,N_9343);
xor U11507 (N_11507,N_8725,N_8885);
and U11508 (N_11508,N_9913,N_8478);
nor U11509 (N_11509,N_9311,N_9640);
or U11510 (N_11510,N_9040,N_9725);
and U11511 (N_11511,N_8442,N_9595);
nor U11512 (N_11512,N_8991,N_9701);
and U11513 (N_11513,N_9580,N_8326);
nand U11514 (N_11514,N_9732,N_9759);
xor U11515 (N_11515,N_9095,N_9136);
nor U11516 (N_11516,N_8117,N_8938);
xor U11517 (N_11517,N_9053,N_8937);
and U11518 (N_11518,N_8347,N_9128);
and U11519 (N_11519,N_8221,N_9962);
nand U11520 (N_11520,N_8994,N_8892);
and U11521 (N_11521,N_9628,N_9119);
xor U11522 (N_11522,N_8222,N_9464);
xnor U11523 (N_11523,N_9359,N_8078);
and U11524 (N_11524,N_8756,N_9727);
or U11525 (N_11525,N_8931,N_8080);
or U11526 (N_11526,N_8111,N_9828);
or U11527 (N_11527,N_9352,N_9921);
nor U11528 (N_11528,N_8994,N_8478);
nor U11529 (N_11529,N_9008,N_9933);
xor U11530 (N_11530,N_9216,N_9625);
xor U11531 (N_11531,N_9964,N_8570);
nand U11532 (N_11532,N_9641,N_9078);
nor U11533 (N_11533,N_9411,N_8181);
nor U11534 (N_11534,N_8637,N_8935);
nand U11535 (N_11535,N_9567,N_8443);
xor U11536 (N_11536,N_8434,N_8852);
and U11537 (N_11537,N_8115,N_8733);
nor U11538 (N_11538,N_9372,N_8904);
xor U11539 (N_11539,N_9586,N_9786);
and U11540 (N_11540,N_8902,N_8965);
nor U11541 (N_11541,N_9114,N_8411);
nor U11542 (N_11542,N_8622,N_9715);
xor U11543 (N_11543,N_9543,N_9046);
nor U11544 (N_11544,N_8700,N_9439);
or U11545 (N_11545,N_8271,N_8247);
nor U11546 (N_11546,N_9027,N_9815);
nand U11547 (N_11547,N_9461,N_8692);
and U11548 (N_11548,N_8229,N_8570);
nand U11549 (N_11549,N_8216,N_9655);
or U11550 (N_11550,N_8701,N_9127);
xor U11551 (N_11551,N_9877,N_8624);
and U11552 (N_11552,N_9404,N_9231);
or U11553 (N_11553,N_8713,N_8741);
or U11554 (N_11554,N_8242,N_8967);
nor U11555 (N_11555,N_9189,N_9300);
nand U11556 (N_11556,N_8686,N_8699);
nor U11557 (N_11557,N_8574,N_8537);
nor U11558 (N_11558,N_9368,N_9874);
nor U11559 (N_11559,N_9349,N_8364);
or U11560 (N_11560,N_8453,N_9511);
or U11561 (N_11561,N_8701,N_8307);
and U11562 (N_11562,N_8070,N_8614);
xnor U11563 (N_11563,N_8842,N_9262);
and U11564 (N_11564,N_9655,N_8188);
nand U11565 (N_11565,N_9314,N_8734);
or U11566 (N_11566,N_9212,N_9243);
nor U11567 (N_11567,N_9784,N_8196);
nor U11568 (N_11568,N_9450,N_8649);
nor U11569 (N_11569,N_9109,N_9652);
or U11570 (N_11570,N_9804,N_8976);
and U11571 (N_11571,N_9236,N_8628);
nor U11572 (N_11572,N_8614,N_9944);
nor U11573 (N_11573,N_8852,N_8339);
nor U11574 (N_11574,N_9639,N_9661);
xnor U11575 (N_11575,N_8054,N_9620);
nor U11576 (N_11576,N_9813,N_8664);
and U11577 (N_11577,N_8697,N_8982);
or U11578 (N_11578,N_9320,N_8001);
or U11579 (N_11579,N_9560,N_9584);
or U11580 (N_11580,N_9483,N_8245);
nand U11581 (N_11581,N_9892,N_8795);
or U11582 (N_11582,N_8152,N_9782);
nor U11583 (N_11583,N_9390,N_8481);
xor U11584 (N_11584,N_8841,N_8482);
xnor U11585 (N_11585,N_8769,N_9848);
xor U11586 (N_11586,N_9432,N_8976);
xor U11587 (N_11587,N_9796,N_8566);
nand U11588 (N_11588,N_8816,N_9989);
nand U11589 (N_11589,N_8837,N_8892);
or U11590 (N_11590,N_8275,N_8544);
xor U11591 (N_11591,N_9550,N_8398);
xnor U11592 (N_11592,N_9564,N_8616);
nand U11593 (N_11593,N_9735,N_8182);
or U11594 (N_11594,N_9080,N_8665);
xor U11595 (N_11595,N_9634,N_9706);
or U11596 (N_11596,N_8225,N_8246);
xnor U11597 (N_11597,N_9638,N_8685);
and U11598 (N_11598,N_9215,N_9276);
or U11599 (N_11599,N_9484,N_9628);
nand U11600 (N_11600,N_9832,N_9860);
nor U11601 (N_11601,N_9326,N_8983);
and U11602 (N_11602,N_8507,N_9430);
nor U11603 (N_11603,N_9969,N_8376);
or U11604 (N_11604,N_8956,N_8117);
and U11605 (N_11605,N_9947,N_9143);
or U11606 (N_11606,N_8809,N_8601);
nand U11607 (N_11607,N_8222,N_8112);
nand U11608 (N_11608,N_9681,N_9730);
and U11609 (N_11609,N_9204,N_8256);
nor U11610 (N_11610,N_8914,N_8466);
and U11611 (N_11611,N_9407,N_9229);
or U11612 (N_11612,N_8270,N_8817);
nor U11613 (N_11613,N_9912,N_9894);
xor U11614 (N_11614,N_9192,N_8143);
and U11615 (N_11615,N_8659,N_9124);
and U11616 (N_11616,N_9598,N_9409);
nor U11617 (N_11617,N_9609,N_8503);
and U11618 (N_11618,N_8632,N_9223);
nand U11619 (N_11619,N_8080,N_9184);
nand U11620 (N_11620,N_8812,N_9340);
xor U11621 (N_11621,N_8522,N_8166);
nand U11622 (N_11622,N_9775,N_9572);
nand U11623 (N_11623,N_9480,N_9373);
and U11624 (N_11624,N_8015,N_8025);
xor U11625 (N_11625,N_9934,N_9546);
xnor U11626 (N_11626,N_9825,N_8109);
nand U11627 (N_11627,N_9127,N_9453);
or U11628 (N_11628,N_9669,N_9131);
nor U11629 (N_11629,N_8394,N_9196);
and U11630 (N_11630,N_8685,N_9531);
nor U11631 (N_11631,N_9522,N_8453);
or U11632 (N_11632,N_8675,N_9006);
nand U11633 (N_11633,N_8274,N_8864);
xor U11634 (N_11634,N_9720,N_8793);
nor U11635 (N_11635,N_8029,N_9204);
nor U11636 (N_11636,N_9766,N_9122);
nor U11637 (N_11637,N_9043,N_9157);
and U11638 (N_11638,N_9084,N_8918);
nor U11639 (N_11639,N_9593,N_9870);
and U11640 (N_11640,N_8984,N_9972);
nand U11641 (N_11641,N_8564,N_9024);
xnor U11642 (N_11642,N_9122,N_8284);
nor U11643 (N_11643,N_8051,N_8577);
xor U11644 (N_11644,N_8782,N_9761);
nor U11645 (N_11645,N_8674,N_9419);
xor U11646 (N_11646,N_9927,N_9077);
and U11647 (N_11647,N_9123,N_8035);
nand U11648 (N_11648,N_9828,N_9099);
or U11649 (N_11649,N_8454,N_8065);
xnor U11650 (N_11650,N_8235,N_8035);
xnor U11651 (N_11651,N_9411,N_9320);
nor U11652 (N_11652,N_9664,N_9316);
and U11653 (N_11653,N_8390,N_9675);
or U11654 (N_11654,N_8310,N_8889);
nor U11655 (N_11655,N_9063,N_9466);
or U11656 (N_11656,N_8886,N_9940);
xnor U11657 (N_11657,N_9598,N_8374);
xnor U11658 (N_11658,N_8286,N_8593);
nand U11659 (N_11659,N_9614,N_8675);
nor U11660 (N_11660,N_8307,N_8903);
xor U11661 (N_11661,N_8941,N_9702);
xnor U11662 (N_11662,N_8883,N_9361);
xnor U11663 (N_11663,N_8289,N_9656);
nand U11664 (N_11664,N_8070,N_9006);
nor U11665 (N_11665,N_8498,N_8841);
and U11666 (N_11666,N_9902,N_8499);
or U11667 (N_11667,N_8991,N_9720);
nand U11668 (N_11668,N_9973,N_9614);
or U11669 (N_11669,N_9749,N_8098);
or U11670 (N_11670,N_9926,N_9476);
xnor U11671 (N_11671,N_8461,N_8053);
xor U11672 (N_11672,N_9525,N_9282);
nand U11673 (N_11673,N_8656,N_9410);
nor U11674 (N_11674,N_8001,N_9723);
nand U11675 (N_11675,N_9979,N_8509);
nand U11676 (N_11676,N_9538,N_8146);
or U11677 (N_11677,N_8012,N_8557);
and U11678 (N_11678,N_8117,N_8806);
nand U11679 (N_11679,N_9191,N_9335);
nand U11680 (N_11680,N_9190,N_8862);
and U11681 (N_11681,N_9520,N_9341);
nor U11682 (N_11682,N_8071,N_8118);
xor U11683 (N_11683,N_9596,N_8358);
nor U11684 (N_11684,N_9442,N_9100);
and U11685 (N_11685,N_8857,N_8044);
nor U11686 (N_11686,N_8871,N_9584);
nor U11687 (N_11687,N_8120,N_8736);
or U11688 (N_11688,N_9295,N_8367);
xor U11689 (N_11689,N_8574,N_9417);
xnor U11690 (N_11690,N_9487,N_9141);
nor U11691 (N_11691,N_9696,N_9366);
nand U11692 (N_11692,N_8575,N_8489);
and U11693 (N_11693,N_9882,N_8276);
xor U11694 (N_11694,N_8589,N_9789);
nor U11695 (N_11695,N_9228,N_9287);
or U11696 (N_11696,N_9895,N_8553);
nand U11697 (N_11697,N_9977,N_9387);
nor U11698 (N_11698,N_8691,N_9234);
or U11699 (N_11699,N_8853,N_9699);
and U11700 (N_11700,N_9011,N_8389);
nand U11701 (N_11701,N_8672,N_9223);
or U11702 (N_11702,N_9511,N_9610);
or U11703 (N_11703,N_8913,N_8305);
nor U11704 (N_11704,N_9004,N_8214);
xnor U11705 (N_11705,N_8139,N_8428);
nor U11706 (N_11706,N_8081,N_9553);
nor U11707 (N_11707,N_9108,N_9424);
xnor U11708 (N_11708,N_9933,N_9676);
nand U11709 (N_11709,N_8593,N_8176);
nand U11710 (N_11710,N_9537,N_9343);
xor U11711 (N_11711,N_9154,N_8128);
nor U11712 (N_11712,N_8171,N_8628);
xnor U11713 (N_11713,N_9819,N_8948);
nor U11714 (N_11714,N_9029,N_8016);
nand U11715 (N_11715,N_9218,N_8927);
xor U11716 (N_11716,N_8038,N_8723);
nor U11717 (N_11717,N_9018,N_8416);
and U11718 (N_11718,N_9690,N_9216);
nand U11719 (N_11719,N_8152,N_8424);
or U11720 (N_11720,N_9353,N_8521);
and U11721 (N_11721,N_8864,N_9614);
xor U11722 (N_11722,N_9143,N_9755);
nor U11723 (N_11723,N_9469,N_9542);
or U11724 (N_11724,N_9310,N_8293);
nor U11725 (N_11725,N_8639,N_8201);
nand U11726 (N_11726,N_9482,N_8079);
xor U11727 (N_11727,N_9597,N_8700);
or U11728 (N_11728,N_9161,N_9123);
and U11729 (N_11729,N_8073,N_9698);
or U11730 (N_11730,N_9543,N_8277);
xor U11731 (N_11731,N_9760,N_8295);
or U11732 (N_11732,N_9986,N_8018);
or U11733 (N_11733,N_9705,N_8692);
xnor U11734 (N_11734,N_9036,N_8326);
or U11735 (N_11735,N_9373,N_9857);
or U11736 (N_11736,N_9858,N_8822);
nand U11737 (N_11737,N_8676,N_8798);
xor U11738 (N_11738,N_9008,N_8576);
nand U11739 (N_11739,N_8809,N_9055);
and U11740 (N_11740,N_8524,N_9233);
xor U11741 (N_11741,N_8050,N_8802);
nor U11742 (N_11742,N_9403,N_8241);
nand U11743 (N_11743,N_8958,N_9035);
xnor U11744 (N_11744,N_9587,N_9698);
and U11745 (N_11745,N_9471,N_8663);
xor U11746 (N_11746,N_9786,N_8568);
or U11747 (N_11747,N_8238,N_9862);
nor U11748 (N_11748,N_8536,N_9572);
or U11749 (N_11749,N_8726,N_8715);
and U11750 (N_11750,N_9353,N_8077);
nor U11751 (N_11751,N_8845,N_9471);
or U11752 (N_11752,N_8644,N_8018);
nand U11753 (N_11753,N_8893,N_9297);
xor U11754 (N_11754,N_9754,N_9099);
xor U11755 (N_11755,N_9335,N_8930);
xnor U11756 (N_11756,N_8818,N_9259);
or U11757 (N_11757,N_8922,N_9807);
or U11758 (N_11758,N_9684,N_8914);
nor U11759 (N_11759,N_8988,N_8708);
or U11760 (N_11760,N_8312,N_8097);
or U11761 (N_11761,N_8988,N_9335);
and U11762 (N_11762,N_9146,N_9945);
or U11763 (N_11763,N_8157,N_9115);
or U11764 (N_11764,N_8201,N_9507);
or U11765 (N_11765,N_8162,N_9034);
or U11766 (N_11766,N_9507,N_9317);
or U11767 (N_11767,N_9215,N_8062);
and U11768 (N_11768,N_8889,N_8518);
nand U11769 (N_11769,N_9588,N_8460);
or U11770 (N_11770,N_9517,N_9467);
or U11771 (N_11771,N_9068,N_9655);
xnor U11772 (N_11772,N_9074,N_9338);
nor U11773 (N_11773,N_9365,N_8412);
xnor U11774 (N_11774,N_8107,N_9870);
nor U11775 (N_11775,N_8796,N_9162);
nor U11776 (N_11776,N_9963,N_8991);
nand U11777 (N_11777,N_9819,N_8333);
nor U11778 (N_11778,N_8820,N_8487);
or U11779 (N_11779,N_8288,N_8772);
nor U11780 (N_11780,N_9438,N_8717);
xor U11781 (N_11781,N_9102,N_9521);
nor U11782 (N_11782,N_9296,N_8050);
nor U11783 (N_11783,N_8757,N_9540);
or U11784 (N_11784,N_9908,N_8313);
or U11785 (N_11785,N_9264,N_8172);
or U11786 (N_11786,N_8022,N_9331);
nand U11787 (N_11787,N_8210,N_9788);
nand U11788 (N_11788,N_9604,N_8087);
and U11789 (N_11789,N_8233,N_8439);
nand U11790 (N_11790,N_8792,N_9698);
nor U11791 (N_11791,N_9450,N_9845);
nor U11792 (N_11792,N_8106,N_8959);
or U11793 (N_11793,N_8487,N_8916);
or U11794 (N_11794,N_8695,N_9499);
xnor U11795 (N_11795,N_9330,N_9718);
nor U11796 (N_11796,N_8876,N_8931);
xnor U11797 (N_11797,N_8750,N_8199);
xnor U11798 (N_11798,N_9291,N_9777);
nor U11799 (N_11799,N_9050,N_8454);
nand U11800 (N_11800,N_8107,N_9931);
or U11801 (N_11801,N_8101,N_9167);
nor U11802 (N_11802,N_9945,N_8237);
and U11803 (N_11803,N_9005,N_9796);
nand U11804 (N_11804,N_9615,N_9024);
and U11805 (N_11805,N_9220,N_9835);
and U11806 (N_11806,N_9954,N_8312);
nand U11807 (N_11807,N_8099,N_9149);
xor U11808 (N_11808,N_8096,N_9733);
or U11809 (N_11809,N_8655,N_8012);
xnor U11810 (N_11810,N_9149,N_8105);
xnor U11811 (N_11811,N_9249,N_9435);
xnor U11812 (N_11812,N_8885,N_9678);
and U11813 (N_11813,N_9533,N_9961);
xnor U11814 (N_11814,N_9649,N_9225);
xor U11815 (N_11815,N_9338,N_8444);
or U11816 (N_11816,N_8865,N_8909);
nand U11817 (N_11817,N_8557,N_9425);
xnor U11818 (N_11818,N_8455,N_8629);
nand U11819 (N_11819,N_9980,N_9453);
nor U11820 (N_11820,N_9951,N_8171);
xnor U11821 (N_11821,N_8668,N_9492);
and U11822 (N_11822,N_9296,N_8799);
and U11823 (N_11823,N_9281,N_9697);
nand U11824 (N_11824,N_9630,N_8031);
nor U11825 (N_11825,N_9205,N_8766);
nor U11826 (N_11826,N_8958,N_9890);
nand U11827 (N_11827,N_9094,N_9655);
and U11828 (N_11828,N_9475,N_8355);
nor U11829 (N_11829,N_8573,N_8788);
or U11830 (N_11830,N_9562,N_8632);
nor U11831 (N_11831,N_8944,N_9217);
and U11832 (N_11832,N_9179,N_9238);
and U11833 (N_11833,N_9226,N_8357);
nor U11834 (N_11834,N_8454,N_8888);
nor U11835 (N_11835,N_8424,N_9267);
or U11836 (N_11836,N_9625,N_8727);
xor U11837 (N_11837,N_8233,N_8096);
nand U11838 (N_11838,N_9855,N_9735);
and U11839 (N_11839,N_9185,N_9563);
nor U11840 (N_11840,N_9816,N_9603);
and U11841 (N_11841,N_9580,N_8916);
or U11842 (N_11842,N_8414,N_8648);
nor U11843 (N_11843,N_8884,N_9277);
or U11844 (N_11844,N_8634,N_9283);
xnor U11845 (N_11845,N_9300,N_8305);
and U11846 (N_11846,N_9735,N_9986);
and U11847 (N_11847,N_9045,N_9071);
nand U11848 (N_11848,N_9526,N_9719);
or U11849 (N_11849,N_8792,N_8427);
nor U11850 (N_11850,N_8355,N_9175);
nand U11851 (N_11851,N_8977,N_9451);
xnor U11852 (N_11852,N_8061,N_9198);
nor U11853 (N_11853,N_8470,N_8409);
nand U11854 (N_11854,N_9291,N_9018);
nand U11855 (N_11855,N_9376,N_9672);
xor U11856 (N_11856,N_9072,N_8657);
nor U11857 (N_11857,N_9147,N_9052);
xor U11858 (N_11858,N_8219,N_8824);
and U11859 (N_11859,N_9755,N_8838);
and U11860 (N_11860,N_9474,N_8717);
nor U11861 (N_11861,N_8623,N_9279);
nand U11862 (N_11862,N_8570,N_8051);
xnor U11863 (N_11863,N_8239,N_9357);
and U11864 (N_11864,N_8814,N_8955);
xor U11865 (N_11865,N_9741,N_8308);
or U11866 (N_11866,N_9940,N_8258);
and U11867 (N_11867,N_9145,N_8229);
xnor U11868 (N_11868,N_8409,N_8310);
nor U11869 (N_11869,N_9183,N_8635);
nor U11870 (N_11870,N_9518,N_8976);
nor U11871 (N_11871,N_9830,N_9377);
and U11872 (N_11872,N_8118,N_8872);
or U11873 (N_11873,N_9036,N_9482);
or U11874 (N_11874,N_8677,N_8193);
xnor U11875 (N_11875,N_8837,N_8338);
nand U11876 (N_11876,N_8762,N_9917);
nor U11877 (N_11877,N_9876,N_9230);
xnor U11878 (N_11878,N_9274,N_9332);
xor U11879 (N_11879,N_9062,N_9714);
xnor U11880 (N_11880,N_9047,N_8778);
and U11881 (N_11881,N_9395,N_8219);
or U11882 (N_11882,N_8975,N_9292);
or U11883 (N_11883,N_9226,N_8383);
xnor U11884 (N_11884,N_9006,N_9692);
xnor U11885 (N_11885,N_9971,N_9446);
nor U11886 (N_11886,N_8521,N_9020);
or U11887 (N_11887,N_8328,N_8904);
nand U11888 (N_11888,N_8926,N_8974);
nor U11889 (N_11889,N_8849,N_8024);
nand U11890 (N_11890,N_9949,N_9458);
nand U11891 (N_11891,N_9139,N_9921);
and U11892 (N_11892,N_8290,N_9858);
and U11893 (N_11893,N_8449,N_9289);
or U11894 (N_11894,N_8795,N_9701);
xnor U11895 (N_11895,N_8498,N_8658);
xor U11896 (N_11896,N_8577,N_9421);
xnor U11897 (N_11897,N_9331,N_8190);
xnor U11898 (N_11898,N_8125,N_8812);
nor U11899 (N_11899,N_8475,N_8409);
and U11900 (N_11900,N_9551,N_8833);
xnor U11901 (N_11901,N_8845,N_9145);
nand U11902 (N_11902,N_9506,N_8954);
xnor U11903 (N_11903,N_8798,N_8459);
nor U11904 (N_11904,N_8518,N_8814);
or U11905 (N_11905,N_8913,N_9066);
nor U11906 (N_11906,N_9809,N_8043);
and U11907 (N_11907,N_8714,N_9963);
nand U11908 (N_11908,N_9358,N_9505);
nor U11909 (N_11909,N_9860,N_8769);
nand U11910 (N_11910,N_8614,N_8324);
xor U11911 (N_11911,N_8562,N_9981);
xor U11912 (N_11912,N_8598,N_9367);
xor U11913 (N_11913,N_8830,N_8975);
nor U11914 (N_11914,N_8298,N_9113);
xnor U11915 (N_11915,N_8693,N_8880);
or U11916 (N_11916,N_9328,N_9695);
nor U11917 (N_11917,N_8353,N_8498);
or U11918 (N_11918,N_9975,N_9764);
xor U11919 (N_11919,N_8439,N_9358);
xor U11920 (N_11920,N_8770,N_8810);
and U11921 (N_11921,N_8764,N_8787);
or U11922 (N_11922,N_9724,N_9966);
nor U11923 (N_11923,N_8357,N_8614);
nor U11924 (N_11924,N_8819,N_9077);
or U11925 (N_11925,N_8495,N_9291);
nand U11926 (N_11926,N_8642,N_8167);
nand U11927 (N_11927,N_8615,N_8628);
and U11928 (N_11928,N_8397,N_8145);
and U11929 (N_11929,N_9092,N_8416);
nand U11930 (N_11930,N_8326,N_8585);
and U11931 (N_11931,N_8082,N_8861);
and U11932 (N_11932,N_8173,N_9062);
xnor U11933 (N_11933,N_9676,N_8903);
xor U11934 (N_11934,N_8215,N_9157);
or U11935 (N_11935,N_8517,N_9689);
and U11936 (N_11936,N_8773,N_9745);
nand U11937 (N_11937,N_8060,N_8067);
or U11938 (N_11938,N_8379,N_8091);
or U11939 (N_11939,N_9671,N_8817);
or U11940 (N_11940,N_8633,N_8755);
and U11941 (N_11941,N_9067,N_8357);
nand U11942 (N_11942,N_8117,N_8032);
nor U11943 (N_11943,N_9239,N_9336);
and U11944 (N_11944,N_8375,N_8527);
and U11945 (N_11945,N_8470,N_8061);
xnor U11946 (N_11946,N_8796,N_8091);
nor U11947 (N_11947,N_8532,N_8261);
or U11948 (N_11948,N_9340,N_8758);
nand U11949 (N_11949,N_8740,N_9796);
nand U11950 (N_11950,N_8912,N_8846);
or U11951 (N_11951,N_9931,N_9696);
xnor U11952 (N_11952,N_8797,N_8071);
or U11953 (N_11953,N_8865,N_9426);
nand U11954 (N_11954,N_8034,N_8089);
or U11955 (N_11955,N_9143,N_8051);
and U11956 (N_11956,N_9438,N_8387);
nand U11957 (N_11957,N_9963,N_9970);
xor U11958 (N_11958,N_8556,N_9162);
xnor U11959 (N_11959,N_8522,N_8630);
and U11960 (N_11960,N_9433,N_9493);
nor U11961 (N_11961,N_8459,N_8639);
and U11962 (N_11962,N_8806,N_9078);
or U11963 (N_11963,N_8463,N_8832);
nor U11964 (N_11964,N_9977,N_9018);
nand U11965 (N_11965,N_8084,N_9061);
nor U11966 (N_11966,N_9990,N_8147);
and U11967 (N_11967,N_9492,N_8871);
xnor U11968 (N_11968,N_8423,N_9488);
nor U11969 (N_11969,N_8919,N_9608);
or U11970 (N_11970,N_9833,N_8910);
and U11971 (N_11971,N_8491,N_9663);
and U11972 (N_11972,N_8198,N_8867);
nor U11973 (N_11973,N_8394,N_9718);
and U11974 (N_11974,N_8785,N_9739);
nor U11975 (N_11975,N_8923,N_9552);
nand U11976 (N_11976,N_8972,N_9626);
and U11977 (N_11977,N_8833,N_9508);
nand U11978 (N_11978,N_8761,N_8033);
xnor U11979 (N_11979,N_8150,N_9931);
or U11980 (N_11980,N_8811,N_8404);
xor U11981 (N_11981,N_8276,N_8577);
or U11982 (N_11982,N_9313,N_9044);
nand U11983 (N_11983,N_8035,N_8281);
nor U11984 (N_11984,N_9409,N_9445);
xor U11985 (N_11985,N_8068,N_9366);
or U11986 (N_11986,N_9367,N_8684);
nor U11987 (N_11987,N_8233,N_8310);
xor U11988 (N_11988,N_9613,N_8648);
xor U11989 (N_11989,N_9111,N_9029);
xor U11990 (N_11990,N_9015,N_8630);
nor U11991 (N_11991,N_8971,N_9784);
or U11992 (N_11992,N_8884,N_9246);
and U11993 (N_11993,N_9145,N_8973);
nor U11994 (N_11994,N_8394,N_8763);
nand U11995 (N_11995,N_9689,N_8264);
xnor U11996 (N_11996,N_9129,N_9048);
nand U11997 (N_11997,N_8474,N_8986);
nand U11998 (N_11998,N_9990,N_9044);
xor U11999 (N_11999,N_9091,N_8360);
nor U12000 (N_12000,N_11182,N_10090);
and U12001 (N_12001,N_11804,N_10313);
nand U12002 (N_12002,N_11516,N_10155);
nor U12003 (N_12003,N_11877,N_10949);
or U12004 (N_12004,N_11460,N_10542);
nor U12005 (N_12005,N_11979,N_10909);
and U12006 (N_12006,N_10958,N_11030);
or U12007 (N_12007,N_10430,N_11492);
xnor U12008 (N_12008,N_11255,N_10849);
and U12009 (N_12009,N_10582,N_11955);
nor U12010 (N_12010,N_10736,N_11686);
or U12011 (N_12011,N_10629,N_11679);
and U12012 (N_12012,N_11896,N_10088);
nand U12013 (N_12013,N_10150,N_10656);
nor U12014 (N_12014,N_10821,N_11588);
and U12015 (N_12015,N_11494,N_11809);
or U12016 (N_12016,N_10559,N_10563);
and U12017 (N_12017,N_11023,N_10390);
and U12018 (N_12018,N_11172,N_11421);
nor U12019 (N_12019,N_10400,N_10641);
nor U12020 (N_12020,N_10707,N_11487);
xnor U12021 (N_12021,N_10189,N_11943);
xor U12022 (N_12022,N_11483,N_10265);
or U12023 (N_12023,N_11858,N_10982);
or U12024 (N_12024,N_10075,N_10588);
xnor U12025 (N_12025,N_10531,N_11723);
and U12026 (N_12026,N_10491,N_11562);
or U12027 (N_12027,N_10851,N_10085);
and U12028 (N_12028,N_10411,N_10346);
or U12029 (N_12029,N_11749,N_11190);
nand U12030 (N_12030,N_10478,N_10252);
xnor U12031 (N_12031,N_11286,N_11260);
and U12032 (N_12032,N_11589,N_10620);
nor U12033 (N_12033,N_10053,N_11549);
or U12034 (N_12034,N_10771,N_10143);
or U12035 (N_12035,N_11221,N_10939);
or U12036 (N_12036,N_10558,N_11083);
nand U12037 (N_12037,N_11504,N_11718);
or U12038 (N_12038,N_11196,N_11513);
nand U12039 (N_12039,N_11142,N_11807);
or U12040 (N_12040,N_10115,N_11954);
nor U12041 (N_12041,N_10870,N_11108);
nand U12042 (N_12042,N_10255,N_10481);
nor U12043 (N_12043,N_10726,N_10826);
and U12044 (N_12044,N_10731,N_10144);
xor U12045 (N_12045,N_10057,N_11508);
nor U12046 (N_12046,N_10112,N_10283);
nand U12047 (N_12047,N_10197,N_11987);
and U12048 (N_12048,N_11825,N_11621);
nor U12049 (N_12049,N_11606,N_11148);
xor U12050 (N_12050,N_11009,N_11453);
and U12051 (N_12051,N_11697,N_11365);
nor U12052 (N_12052,N_11950,N_11355);
nand U12053 (N_12053,N_10887,N_10300);
xnor U12054 (N_12054,N_11730,N_11931);
or U12055 (N_12055,N_10750,N_10258);
nand U12056 (N_12056,N_10066,N_11257);
and U12057 (N_12057,N_10050,N_10788);
or U12058 (N_12058,N_11726,N_10698);
xor U12059 (N_12059,N_10477,N_10480);
and U12060 (N_12060,N_10604,N_10800);
or U12061 (N_12061,N_10298,N_11473);
and U12062 (N_12062,N_10233,N_11493);
or U12063 (N_12063,N_11881,N_11534);
and U12064 (N_12064,N_10162,N_10408);
nand U12065 (N_12065,N_11234,N_11966);
nor U12066 (N_12066,N_10371,N_10482);
or U12067 (N_12067,N_11946,N_11694);
nand U12068 (N_12068,N_10178,N_11829);
nor U12069 (N_12069,N_10876,N_10494);
nor U12070 (N_12070,N_11282,N_11795);
and U12071 (N_12071,N_11957,N_10734);
nor U12072 (N_12072,N_10513,N_11331);
or U12073 (N_12073,N_11969,N_10626);
nand U12074 (N_12074,N_11747,N_11936);
nor U12075 (N_12075,N_10625,N_11635);
and U12076 (N_12076,N_10099,N_10303);
nand U12077 (N_12077,N_10093,N_11646);
nor U12078 (N_12078,N_11060,N_11610);
nand U12079 (N_12079,N_10510,N_11456);
nor U12080 (N_12080,N_10406,N_10211);
nand U12081 (N_12081,N_11432,N_11146);
or U12082 (N_12082,N_10727,N_11386);
nor U12083 (N_12083,N_11075,N_10264);
or U12084 (N_12084,N_10945,N_11011);
nand U12085 (N_12085,N_10879,N_10368);
nor U12086 (N_12086,N_10244,N_11485);
and U12087 (N_12087,N_10074,N_11174);
or U12088 (N_12088,N_10677,N_11596);
nor U12089 (N_12089,N_11971,N_11164);
and U12090 (N_12090,N_11656,N_11711);
and U12091 (N_12091,N_10769,N_11844);
nand U12092 (N_12092,N_10512,N_11239);
or U12093 (N_12093,N_11873,N_11007);
nand U12094 (N_12094,N_10374,N_10918);
xor U12095 (N_12095,N_10350,N_10511);
and U12096 (N_12096,N_11527,N_10796);
or U12097 (N_12097,N_11441,N_10396);
nand U12098 (N_12098,N_11219,N_10662);
and U12099 (N_12099,N_10543,N_10683);
nor U12100 (N_12100,N_10185,N_10603);
nand U12101 (N_12101,N_11826,N_10779);
nand U12102 (N_12102,N_10139,N_10899);
xor U12103 (N_12103,N_11842,N_10541);
nor U12104 (N_12104,N_11690,N_10856);
xor U12105 (N_12105,N_11019,N_10450);
and U12106 (N_12106,N_11773,N_11663);
nand U12107 (N_12107,N_11056,N_11698);
or U12108 (N_12108,N_11488,N_11783);
or U12109 (N_12109,N_10621,N_10397);
xnor U12110 (N_12110,N_11367,N_10888);
nand U12111 (N_12111,N_10087,N_11294);
and U12112 (N_12112,N_11029,N_10154);
or U12113 (N_12113,N_11292,N_10033);
nand U12114 (N_12114,N_10292,N_11478);
xor U12115 (N_12115,N_10159,N_10871);
or U12116 (N_12116,N_10591,N_10366);
and U12117 (N_12117,N_10960,N_11303);
xor U12118 (N_12118,N_10343,N_10135);
nor U12119 (N_12119,N_11543,N_11528);
or U12120 (N_12120,N_10897,N_10984);
or U12121 (N_12121,N_11592,N_11402);
nor U12122 (N_12122,N_11268,N_11569);
xnor U12123 (N_12123,N_11976,N_11535);
xor U12124 (N_12124,N_11249,N_10152);
nand U12125 (N_12125,N_10381,N_11093);
nand U12126 (N_12126,N_10000,N_10331);
and U12127 (N_12127,N_11890,N_10966);
xor U12128 (N_12128,N_11160,N_10476);
xnor U12129 (N_12129,N_10978,N_11820);
nand U12130 (N_12130,N_10184,N_10086);
or U12131 (N_12131,N_10901,N_11886);
nor U12132 (N_12132,N_11774,N_11607);
and U12133 (N_12133,N_10117,N_11824);
xnor U12134 (N_12134,N_10239,N_11152);
and U12135 (N_12135,N_10113,N_11150);
nor U12136 (N_12136,N_11887,N_11379);
nor U12137 (N_12137,N_11756,N_10606);
and U12138 (N_12138,N_10109,N_11736);
or U12139 (N_12139,N_10742,N_10860);
nor U12140 (N_12140,N_11251,N_10457);
or U12141 (N_12141,N_10027,N_11900);
nand U12142 (N_12142,N_10003,N_10379);
or U12143 (N_12143,N_11638,N_10056);
xnor U12144 (N_12144,N_10607,N_11136);
nor U12145 (N_12145,N_10496,N_10845);
nand U12146 (N_12146,N_11129,N_11475);
and U12147 (N_12147,N_11835,N_11857);
xor U12148 (N_12148,N_10593,N_10597);
or U12149 (N_12149,N_11574,N_11158);
xnor U12150 (N_12150,N_11440,N_10728);
xor U12151 (N_12151,N_10391,N_11306);
nor U12152 (N_12152,N_10425,N_10441);
nor U12153 (N_12153,N_10141,N_11999);
xor U12154 (N_12154,N_11984,N_10904);
nand U12155 (N_12155,N_11841,N_10746);
or U12156 (N_12156,N_11356,N_11206);
nor U12157 (N_12157,N_10883,N_10912);
or U12158 (N_12158,N_10474,N_10323);
nand U12159 (N_12159,N_11350,N_10289);
or U12160 (N_12160,N_10008,N_10961);
nor U12161 (N_12161,N_11275,N_10758);
nand U12162 (N_12162,N_11342,N_10589);
nor U12163 (N_12163,N_11173,N_10610);
nand U12164 (N_12164,N_11015,N_10175);
and U12165 (N_12165,N_11049,N_10617);
nand U12166 (N_12166,N_10191,N_10213);
nor U12167 (N_12167,N_10473,N_11851);
nand U12168 (N_12168,N_11098,N_11031);
or U12169 (N_12169,N_11256,N_11565);
nand U12170 (N_12170,N_11405,N_11328);
nand U12171 (N_12171,N_11143,N_11016);
and U12172 (N_12172,N_11057,N_11772);
nor U12173 (N_12173,N_11313,N_10520);
or U12174 (N_12174,N_11415,N_10544);
and U12175 (N_12175,N_11464,N_10747);
nand U12176 (N_12176,N_10171,N_10719);
or U12177 (N_12177,N_11994,N_11265);
and U12178 (N_12178,N_10007,N_10556);
or U12179 (N_12179,N_11557,N_10377);
xnor U12180 (N_12180,N_11325,N_10266);
nand U12181 (N_12181,N_11186,N_10598);
xor U12182 (N_12182,N_10420,N_11054);
nor U12183 (N_12183,N_11799,N_11733);
and U12184 (N_12184,N_10678,N_11899);
xor U12185 (N_12185,N_11169,N_10032);
nor U12186 (N_12186,N_11546,N_11720);
nor U12187 (N_12187,N_11207,N_11981);
and U12188 (N_12188,N_11162,N_11629);
nor U12189 (N_12189,N_10291,N_10015);
nand U12190 (N_12190,N_11340,N_10124);
nand U12191 (N_12191,N_10739,N_10226);
xor U12192 (N_12192,N_10757,N_10262);
or U12193 (N_12193,N_10819,N_11768);
xnor U12194 (N_12194,N_10118,N_11601);
and U12195 (N_12195,N_10704,N_11700);
xnor U12196 (N_12196,N_11530,N_10241);
nor U12197 (N_12197,N_11932,N_10082);
nand U12198 (N_12198,N_11259,N_11539);
nand U12199 (N_12199,N_10401,N_11935);
nor U12200 (N_12200,N_10855,N_10920);
nand U12201 (N_12201,N_11753,N_10680);
and U12202 (N_12202,N_10304,N_11874);
or U12203 (N_12203,N_11041,N_11912);
xor U12204 (N_12204,N_10272,N_10914);
nor U12205 (N_12205,N_10947,N_11620);
nand U12206 (N_12206,N_11184,N_11094);
nand U12207 (N_12207,N_11625,N_10455);
xor U12208 (N_12208,N_11645,N_10985);
nor U12209 (N_12209,N_10181,N_10247);
or U12210 (N_12210,N_10072,N_10690);
or U12211 (N_12211,N_11354,N_11231);
xnor U12212 (N_12212,N_11412,N_11246);
xor U12213 (N_12213,N_11691,N_10515);
nor U12214 (N_12214,N_10850,N_11420);
xor U12215 (N_12215,N_10301,N_11069);
nand U12216 (N_12216,N_10808,N_10105);
nand U12217 (N_12217,N_10633,N_10073);
xor U12218 (N_12218,N_10164,N_10968);
or U12219 (N_12219,N_11904,N_10638);
xor U12220 (N_12220,N_10485,N_10717);
or U12221 (N_12221,N_10426,N_10900);
and U12222 (N_12222,N_11208,N_11731);
nand U12223 (N_12223,N_10219,N_11166);
or U12224 (N_12224,N_10334,N_10970);
xor U12225 (N_12225,N_11649,N_11653);
and U12226 (N_12226,N_11805,N_10789);
xnor U12227 (N_12227,N_11659,N_11225);
and U12228 (N_12228,N_11838,N_10890);
and U12229 (N_12229,N_11876,N_10893);
nand U12230 (N_12230,N_11764,N_11024);
xor U12231 (N_12231,N_10695,N_10770);
nor U12232 (N_12232,N_11223,N_11312);
nor U12233 (N_12233,N_11704,N_10803);
nand U12234 (N_12234,N_10632,N_10243);
and U12235 (N_12235,N_10134,N_10248);
xnor U12236 (N_12236,N_10460,N_10205);
nand U12237 (N_12237,N_11837,N_11407);
and U12238 (N_12238,N_11895,N_11665);
and U12239 (N_12239,N_10995,N_11297);
nor U12240 (N_12240,N_11237,N_10299);
nor U12241 (N_12241,N_10596,N_11972);
and U12242 (N_12242,N_11671,N_11018);
xnor U12243 (N_12243,N_11875,N_11830);
and U12244 (N_12244,N_10378,N_10005);
and U12245 (N_12245,N_10220,N_11314);
and U12246 (N_12246,N_10784,N_11337);
nor U12247 (N_12247,N_10691,N_11622);
nor U12248 (N_12248,N_10357,N_11202);
nand U12249 (N_12249,N_10120,N_10980);
nand U12250 (N_12250,N_11428,N_10140);
or U12251 (N_12251,N_11819,N_10853);
nand U12252 (N_12252,N_11640,N_10906);
nor U12253 (N_12253,N_10230,N_10974);
xnor U12254 (N_12254,N_11116,N_11933);
and U12255 (N_12255,N_11956,N_11360);
or U12256 (N_12256,N_10358,N_10294);
xnor U12257 (N_12257,N_11263,N_11803);
or U12258 (N_12258,N_10635,N_10212);
or U12259 (N_12259,N_11616,N_11572);
nor U12260 (N_12260,N_11866,N_11266);
nand U12261 (N_12261,N_11595,N_11279);
nor U12262 (N_12262,N_10297,N_10147);
and U12263 (N_12263,N_10857,N_10242);
xnor U12264 (N_12264,N_11394,N_10192);
nand U12265 (N_12265,N_11114,N_11644);
nor U12266 (N_12266,N_11037,N_11205);
nor U12267 (N_12267,N_10196,N_11179);
xor U12268 (N_12268,N_11519,N_11717);
or U12269 (N_12269,N_10972,N_11135);
xor U12270 (N_12270,N_10993,N_10844);
and U12271 (N_12271,N_11520,N_10538);
or U12272 (N_12272,N_10574,N_11909);
or U12273 (N_12273,N_11132,N_11982);
nand U12274 (N_12274,N_10356,N_10654);
nand U12275 (N_12275,N_10173,N_11657);
and U12276 (N_12276,N_10684,N_11005);
or U12277 (N_12277,N_10138,N_11967);
nand U12278 (N_12278,N_11538,N_11423);
xor U12279 (N_12279,N_10605,N_11105);
xor U12280 (N_12280,N_10250,N_10981);
nand U12281 (N_12281,N_11288,N_11668);
xnor U12282 (N_12282,N_10667,N_11849);
and U12283 (N_12283,N_11194,N_11776);
nand U12284 (N_12284,N_11085,N_10555);
and U12285 (N_12285,N_11099,N_11871);
nor U12286 (N_12286,N_11759,N_11253);
xnor U12287 (N_12287,N_11082,N_11167);
xnor U12288 (N_12288,N_11670,N_11469);
or U12289 (N_12289,N_11087,N_11079);
nor U12290 (N_12290,N_11214,N_11370);
nor U12291 (N_12291,N_10714,N_11917);
or U12292 (N_12292,N_10565,N_10353);
nor U12293 (N_12293,N_10754,N_11706);
xnor U12294 (N_12294,N_11518,N_10218);
and U12295 (N_12295,N_10094,N_10837);
or U12296 (N_12296,N_10385,N_11524);
or U12297 (N_12297,N_10882,N_10711);
nand U12298 (N_12298,N_11074,N_10471);
xor U12299 (N_12299,N_11419,N_11058);
and U12300 (N_12300,N_10669,N_10025);
and U12301 (N_12301,N_11088,N_11168);
nand U12302 (N_12302,N_10658,N_11341);
nand U12303 (N_12303,N_10752,N_11293);
nand U12304 (N_12304,N_11163,N_11398);
xnor U12305 (N_12305,N_10534,N_10487);
nor U12306 (N_12306,N_11865,N_11983);
nor U12307 (N_12307,N_11159,N_11787);
xor U12308 (N_12308,N_10278,N_11335);
nand U12309 (N_12309,N_11115,N_11126);
nand U12310 (N_12310,N_11978,N_10738);
and U12311 (N_12311,N_10125,N_11920);
xor U12312 (N_12312,N_11351,N_10873);
nor U12313 (N_12313,N_10791,N_10994);
nand U12314 (N_12314,N_10618,N_11846);
or U12315 (N_12315,N_11553,N_11675);
nand U12316 (N_12316,N_11725,N_11210);
nor U12317 (N_12317,N_10345,N_10838);
nand U12318 (N_12318,N_10193,N_11063);
xnor U12319 (N_12319,N_10666,N_10664);
or U12320 (N_12320,N_11199,N_10035);
and U12321 (N_12321,N_11848,N_11677);
xor U12322 (N_12322,N_11183,N_10089);
and U12323 (N_12323,N_10720,N_10790);
and U12324 (N_12324,N_11727,N_10330);
or U12325 (N_12325,N_11302,N_11450);
and U12326 (N_12326,N_11012,N_10933);
xnor U12327 (N_12327,N_10528,N_10163);
nand U12328 (N_12328,N_10327,N_10979);
or U12329 (N_12329,N_10448,N_11233);
xor U12330 (N_12330,N_11119,N_11307);
xnor U12331 (N_12331,N_10898,N_10499);
or U12332 (N_12332,N_11793,N_11821);
or U12333 (N_12333,N_11921,N_11661);
xor U12334 (N_12334,N_10367,N_11106);
nand U12335 (N_12335,N_10240,N_11792);
or U12336 (N_12336,N_10546,N_10232);
nor U12337 (N_12337,N_10081,N_10762);
or U12338 (N_12338,N_11790,N_10288);
and U12339 (N_12339,N_10760,N_10409);
nor U12340 (N_12340,N_10608,N_10560);
xor U12341 (N_12341,N_11436,N_10602);
and U12342 (N_12342,N_11339,N_11027);
or U12343 (N_12343,N_10277,N_10279);
xor U12344 (N_12344,N_10780,N_10364);
nand U12345 (N_12345,N_11375,N_10001);
nand U12346 (N_12346,N_10864,N_10946);
and U12347 (N_12347,N_11178,N_10428);
nand U12348 (N_12348,N_10312,N_10149);
nor U12349 (N_12349,N_10948,N_11544);
and U12350 (N_12350,N_11879,N_10701);
nand U12351 (N_12351,N_11669,N_11579);
xnor U12352 (N_12352,N_10263,N_11376);
nor U12353 (N_12353,N_11346,N_11468);
or U12354 (N_12354,N_11811,N_10136);
nor U12355 (N_12355,N_11859,N_10040);
nand U12356 (N_12356,N_10624,N_11134);
and U12357 (N_12357,N_10369,N_11861);
nand U12358 (N_12358,N_10158,N_11446);
xor U12359 (N_12359,N_10080,N_10523);
nor U12360 (N_12360,N_11997,N_10335);
xor U12361 (N_12361,N_11109,N_11385);
and U12362 (N_12362,N_10648,N_11388);
nand U12363 (N_12363,N_10786,N_10270);
nor U12364 (N_12364,N_11433,N_11600);
and U12365 (N_12365,N_10681,N_10071);
xnor U12366 (N_12366,N_10675,N_10551);
nor U12367 (N_12367,N_11964,N_10387);
nand U12368 (N_12368,N_11988,N_10340);
nor U12369 (N_12369,N_10924,N_11794);
xor U12370 (N_12370,N_11953,N_10527);
nor U12371 (N_12371,N_10502,N_10862);
or U12372 (N_12372,N_10505,N_10581);
and U12373 (N_12373,N_11195,N_11028);
or U12374 (N_12374,N_10011,N_11867);
or U12375 (N_12375,N_10932,N_10922);
or U12376 (N_12376,N_10157,N_10380);
and U12377 (N_12377,N_10650,N_11431);
xor U12378 (N_12378,N_11796,N_10835);
xnor U12379 (N_12379,N_10503,N_10399);
and U12380 (N_12380,N_11853,N_10891);
nor U12381 (N_12381,N_11280,N_11816);
xor U12382 (N_12382,N_10584,N_11380);
nor U12383 (N_12383,N_10273,N_11715);
xnor U12384 (N_12384,N_11914,N_11585);
nand U12385 (N_12385,N_10464,N_11065);
xor U12386 (N_12386,N_10537,N_10095);
nand U12387 (N_12387,N_11533,N_11636);
or U12388 (N_12388,N_11020,N_11227);
xnor U12389 (N_12389,N_10319,N_11501);
nand U12390 (N_12390,N_10059,N_10063);
xnor U12391 (N_12391,N_10238,N_10889);
and U12392 (N_12392,N_11322,N_10166);
or U12393 (N_12393,N_11685,N_11652);
nand U12394 (N_12394,N_10023,N_10365);
nand U12395 (N_12395,N_10514,N_10236);
nand U12396 (N_12396,N_11140,N_10637);
or U12397 (N_12397,N_11482,N_11854);
nor U12398 (N_12398,N_11362,N_11568);
nor U12399 (N_12399,N_10058,N_11597);
nand U12400 (N_12400,N_11403,N_10868);
and U12401 (N_12401,N_11800,N_11091);
or U12402 (N_12402,N_11623,N_10322);
xor U12403 (N_12403,N_10841,N_11959);
nand U12404 (N_12404,N_10030,N_10259);
nor U12405 (N_12405,N_10601,N_10116);
nand U12406 (N_12406,N_10179,N_10102);
xnor U12407 (N_12407,N_10685,N_10067);
xnor U12408 (N_12408,N_10045,N_10999);
and U12409 (N_12409,N_11919,N_11590);
or U12410 (N_12410,N_11758,N_10100);
nor U12411 (N_12411,N_11358,N_10828);
nor U12412 (N_12412,N_10165,N_11090);
or U12413 (N_12413,N_10014,N_10987);
and U12414 (N_12414,N_11422,N_11683);
and U12415 (N_12415,N_11701,N_10311);
nand U12416 (N_12416,N_10938,N_10903);
nand U12417 (N_12417,N_11244,N_10051);
nand U12418 (N_12418,N_11141,N_10772);
and U12419 (N_12419,N_10347,N_11515);
nand U12420 (N_12420,N_10777,N_11902);
or U12421 (N_12421,N_11770,N_10160);
and U12422 (N_12422,N_10452,N_10037);
xnor U12423 (N_12423,N_11133,N_10579);
nand U12424 (N_12424,N_10921,N_10847);
and U12425 (N_12425,N_11343,N_11203);
xor U12426 (N_12426,N_10091,N_10983);
xor U12427 (N_12427,N_10807,N_11489);
nor U12428 (N_12428,N_11371,N_11383);
nand U12429 (N_12429,N_11408,N_11414);
nor U12430 (N_12430,N_11329,N_11710);
nand U12431 (N_12431,N_10561,N_11850);
or U12432 (N_12432,N_11102,N_11930);
and U12433 (N_12433,N_11444,N_10630);
xnor U12434 (N_12434,N_10451,N_11377);
or U12435 (N_12435,N_11502,N_11901);
nor U12436 (N_12436,N_10442,N_11532);
or U12437 (N_12437,N_10416,N_10148);
xnor U12438 (N_12438,N_11941,N_10043);
nand U12439 (N_12439,N_11748,N_11801);
nand U12440 (N_12440,N_10054,N_11630);
nand U12441 (N_12441,N_10493,N_11171);
xnor U12442 (N_12442,N_10700,N_11180);
or U12443 (N_12443,N_11406,N_11689);
and U12444 (N_12444,N_11952,N_10077);
xor U12445 (N_12445,N_10950,N_11537);
or U12446 (N_12446,N_10740,N_11192);
or U12447 (N_12447,N_11334,N_11884);
xor U12448 (N_12448,N_10815,N_11637);
nor U12449 (N_12449,N_11110,N_11061);
and U12450 (N_12450,N_10169,N_11215);
and U12451 (N_12451,N_11870,N_11791);
or U12452 (N_12452,N_11359,N_11942);
or U12453 (N_12453,N_11430,N_10142);
and U12454 (N_12454,N_11033,N_10098);
or U12455 (N_12455,N_10216,N_11076);
or U12456 (N_12456,N_10127,N_11789);
nand U12457 (N_12457,N_11240,N_11443);
nand U12458 (N_12458,N_10461,N_11261);
or U12459 (N_12459,N_11584,N_10229);
nand U12460 (N_12460,N_10062,N_11176);
and U12461 (N_12461,N_10595,N_10955);
nand U12462 (N_12462,N_11366,N_11754);
nor U12463 (N_12463,N_11357,N_10393);
nor U12464 (N_12464,N_10097,N_11071);
nand U12465 (N_12465,N_11566,N_11304);
nor U12466 (N_12466,N_11352,N_10768);
and U12467 (N_12467,N_10552,N_10506);
or U12468 (N_12468,N_11096,N_11961);
nand U12469 (N_12469,N_10321,N_10956);
nand U12470 (N_12470,N_11555,N_10553);
or U12471 (N_12471,N_10529,N_10612);
nor U12472 (N_12472,N_10910,N_10295);
xor U12473 (N_12473,N_10281,N_10101);
and U12474 (N_12474,N_10307,N_10475);
nand U12475 (N_12475,N_11291,N_11051);
nor U12476 (N_12476,N_10820,N_11285);
nand U12477 (N_12477,N_10942,N_10863);
or U12478 (N_12478,N_10592,N_10465);
nor U12479 (N_12479,N_11017,N_11642);
or U12480 (N_12480,N_10619,N_10470);
nor U12481 (N_12481,N_10881,N_11561);
and U12482 (N_12482,N_11705,N_11613);
or U12483 (N_12483,N_10383,N_10781);
and U12484 (N_12484,N_10314,N_11521);
or U12485 (N_12485,N_10806,N_11712);
nand U12486 (N_12486,N_11591,N_10965);
xor U12487 (N_12487,N_11880,N_10645);
nor U12488 (N_12488,N_10123,N_11369);
and U12489 (N_12489,N_10251,N_10586);
or U12490 (N_12490,N_10692,N_10111);
xor U12491 (N_12491,N_10352,N_11300);
and U12492 (N_12492,N_10814,N_11393);
nand U12493 (N_12493,N_10957,N_11187);
xnor U12494 (N_12494,N_10745,N_10469);
nor U12495 (N_12495,N_11235,N_10308);
or U12496 (N_12496,N_11573,N_11138);
or U12497 (N_12497,N_10729,N_10895);
and U12498 (N_12498,N_11062,N_10539);
and U12499 (N_12499,N_10268,N_11211);
nand U12500 (N_12500,N_11678,N_11048);
and U12501 (N_12501,N_11722,N_11684);
or U12502 (N_12502,N_10068,N_11626);
and U12503 (N_12503,N_10296,N_10200);
and U12504 (N_12504,N_11778,N_10570);
and U12505 (N_12505,N_11614,N_10713);
xnor U12506 (N_12506,N_10699,N_10599);
or U12507 (N_12507,N_11752,N_10959);
nor U12508 (N_12508,N_11739,N_10341);
xnor U12509 (N_12509,N_11654,N_10817);
and U12510 (N_12510,N_11201,N_10569);
and U12511 (N_12511,N_11818,N_11270);
and U12512 (N_12512,N_11741,N_11598);
xor U12513 (N_12513,N_11633,N_10203);
nand U12514 (N_12514,N_10526,N_10830);
and U12515 (N_12515,N_11860,N_10907);
and U12516 (N_12516,N_10280,N_10207);
and U12517 (N_12517,N_11651,N_10083);
and U12518 (N_12518,N_11021,N_11949);
nand U12519 (N_12519,N_11289,N_10519);
and U12520 (N_12520,N_10886,N_11298);
and U12521 (N_12521,N_10484,N_11276);
or U12522 (N_12522,N_10293,N_11046);
nor U12523 (N_12523,N_10962,N_11911);
xnor U12524 (N_12524,N_10878,N_10517);
nand U12525 (N_12525,N_11193,N_11882);
nand U12526 (N_12526,N_11052,N_10609);
and U12527 (N_12527,N_11695,N_11862);
xor U12528 (N_12528,N_10445,N_11026);
or U12529 (N_12529,N_11274,N_10816);
or U12530 (N_12530,N_11278,N_11389);
xor U12531 (N_12531,N_11245,N_11960);
nor U12532 (N_12532,N_10682,N_11578);
nor U12533 (N_12533,N_10227,N_11889);
nor U12534 (N_12534,N_11438,N_11181);
nand U12535 (N_12535,N_11391,N_10217);
or U12536 (N_12536,N_11459,N_10804);
nand U12537 (N_12537,N_11232,N_10778);
and U12538 (N_12538,N_10285,N_11089);
xnor U12539 (N_12539,N_10577,N_11632);
xor U12540 (N_12540,N_10204,N_11897);
or U12541 (N_12541,N_10706,N_10351);
xnor U12542 (N_12542,N_11531,N_11053);
and U12543 (N_12543,N_11913,N_11229);
nor U12544 (N_12544,N_11022,N_10201);
nand U12545 (N_12545,N_10730,N_10104);
or U12546 (N_12546,N_10753,N_10359);
or U12547 (N_12547,N_11575,N_10657);
xor U12548 (N_12548,N_10320,N_11055);
nand U12549 (N_12549,N_10765,N_10774);
nor U12550 (N_12550,N_10813,N_10575);
and U12551 (N_12551,N_10671,N_11353);
nor U12552 (N_12552,N_10687,N_11499);
nand U12553 (N_12553,N_10508,N_10468);
or U12554 (N_12554,N_11338,N_10718);
and U12555 (N_12555,N_11814,N_10550);
nor U12556 (N_12556,N_11248,N_11937);
nor U12557 (N_12557,N_10249,N_10854);
xor U12558 (N_12558,N_11287,N_11097);
nand U12559 (N_12559,N_11893,N_11505);
and U12560 (N_12560,N_10600,N_11409);
nor U12561 (N_12561,N_10696,N_11107);
xnor U12562 (N_12562,N_11465,N_11583);
and U12563 (N_12563,N_10064,N_10723);
xnor U12564 (N_12564,N_10483,N_11608);
nor U12565 (N_12565,N_10636,N_10302);
and U12566 (N_12566,N_11666,N_10659);
nand U12567 (N_12567,N_11156,N_10188);
nor U12568 (N_12568,N_10818,N_11230);
nand U12569 (N_12569,N_11451,N_11247);
xnor U12570 (N_12570,N_10079,N_10458);
nor U12571 (N_12571,N_11891,N_10829);
nand U12572 (N_12572,N_11045,N_11777);
xnor U12573 (N_12573,N_10348,N_11693);
and U12574 (N_12574,N_11550,N_11477);
or U12575 (N_12575,N_11922,N_10501);
nand U12576 (N_12576,N_10132,N_11604);
and U12577 (N_12577,N_10869,N_11449);
and U12578 (N_12578,N_10256,N_10545);
or U12579 (N_12579,N_10686,N_11615);
nor U12580 (N_12580,N_11498,N_11760);
xor U12581 (N_12581,N_10284,N_11781);
nor U12582 (N_12582,N_11599,N_11382);
and U12583 (N_12583,N_11836,N_10875);
nand U12584 (N_12584,N_10724,N_11204);
and U12585 (N_12585,N_11486,N_10916);
nor U12586 (N_12586,N_11915,N_11560);
or U12587 (N_12587,N_10186,N_11556);
and U12588 (N_12588,N_11373,N_10896);
and U12589 (N_12589,N_11296,N_11918);
and U12590 (N_12590,N_10114,N_11241);
nand U12591 (N_12591,N_11004,N_10590);
nand U12592 (N_12592,N_10253,N_11827);
nand U12593 (N_12593,N_10454,N_11479);
and U12594 (N_12594,N_10509,N_10151);
nand U12595 (N_12595,N_10766,N_10824);
nor U12596 (N_12596,N_11008,N_10246);
or U12597 (N_12597,N_10344,N_11905);
and U12598 (N_12598,N_10438,N_10052);
or U12599 (N_12599,N_10874,N_10013);
and U12600 (N_12600,N_10422,N_11864);
nand U12601 (N_12601,N_11746,N_10764);
or U12602 (N_12602,N_10661,N_11514);
nand U12603 (N_12603,N_10616,N_11080);
nor U12604 (N_12604,N_11552,N_10649);
and U12605 (N_12605,N_10846,N_10905);
or U12606 (N_12606,N_11529,N_10414);
nor U12607 (N_12607,N_11766,N_11605);
and U12608 (N_12608,N_11729,N_10783);
or U12609 (N_12609,N_11197,N_10653);
nand U12610 (N_12610,N_11564,N_11878);
and U12611 (N_12611,N_10180,N_10915);
nor U12612 (N_12612,N_10640,N_11908);
xor U12613 (N_12613,N_11462,N_11650);
nor U12614 (N_12614,N_10756,N_11283);
xor U12615 (N_12615,N_10798,N_11927);
or U12616 (N_12616,N_10221,N_10261);
nand U12617 (N_12617,N_11744,N_10012);
nand U12618 (N_12618,N_11680,N_11970);
or U12619 (N_12619,N_11923,N_10413);
and U12620 (N_12620,N_11467,N_10562);
or U12621 (N_12621,N_11145,N_10833);
xnor U12622 (N_12622,N_11869,N_11582);
nand U12623 (N_12623,N_10540,N_11001);
nor U12624 (N_12624,N_10872,N_11418);
and U12625 (N_12625,N_11673,N_10467);
nor U12626 (N_12626,N_10429,N_11929);
nor U12627 (N_12627,N_10009,N_11013);
or U12628 (N_12628,N_11782,N_10398);
and U12629 (N_12629,N_10504,N_11332);
or U12630 (N_12630,N_11570,N_10363);
nand U12631 (N_12631,N_10388,N_10930);
and U12632 (N_12632,N_11660,N_10997);
nand U12633 (N_12633,N_10190,N_11429);
nand U12634 (N_12634,N_10827,N_10708);
nor U12635 (N_12635,N_11852,N_11831);
nand U12636 (N_12636,N_10885,N_11628);
nor U12637 (N_12637,N_11035,N_11522);
nand U12638 (N_12638,N_11305,N_11284);
nor U12639 (N_12639,N_10926,N_10567);
nor U12640 (N_12640,N_10759,N_11810);
nand U12641 (N_12641,N_11577,N_11993);
nor U12642 (N_12642,N_10549,N_10392);
nor U12643 (N_12643,N_10977,N_10432);
nor U12644 (N_12644,N_11548,N_11154);
or U12645 (N_12645,N_11426,N_11986);
or U12646 (N_12646,N_10183,N_10048);
xor U12647 (N_12647,N_10022,N_11563);
or U12648 (N_12648,N_11345,N_10389);
xor U12649 (N_12649,N_10732,N_10443);
or U12650 (N_12650,N_10020,N_10848);
or U12651 (N_12651,N_11424,N_11551);
nand U12652 (N_12652,N_10038,N_11481);
or U12653 (N_12653,N_11973,N_10967);
nand U12654 (N_12654,N_11243,N_10177);
and U12655 (N_12655,N_10194,N_11363);
and U12656 (N_12656,N_11643,N_10709);
nor U12657 (N_12657,N_10583,N_11315);
xor U12658 (N_12658,N_11618,N_11939);
xnor U12659 (N_12659,N_11798,N_11272);
nand U12660 (N_12660,N_11855,N_11903);
and U12661 (N_12661,N_11813,N_11751);
or U12662 (N_12662,N_10395,N_10336);
nor U12663 (N_12663,N_11702,N_10842);
nor U12664 (N_12664,N_10462,N_10614);
or U12665 (N_12665,N_11258,N_10755);
nand U12666 (N_12666,N_11425,N_10525);
nor U12667 (N_12667,N_11639,N_11101);
nor U12668 (N_12668,N_11699,N_10834);
nand U12669 (N_12669,N_11455,N_11496);
nand U12670 (N_12670,N_10222,N_11536);
xor U12671 (N_12671,N_11435,N_11916);
nor U12672 (N_12672,N_11907,N_11025);
nand U12673 (N_12673,N_11427,N_10403);
nand U12674 (N_12674,N_11822,N_10908);
xnor U12675 (N_12675,N_11655,N_10710);
nor U12676 (N_12676,N_10006,N_11139);
and U12677 (N_12677,N_10195,N_10224);
xor U12678 (N_12678,N_11463,N_10858);
and U12679 (N_12679,N_11311,N_10145);
nand U12680 (N_12680,N_10799,N_11617);
and U12681 (N_12681,N_10447,N_11308);
and U12682 (N_12682,N_11144,N_11175);
nand U12683 (N_12683,N_10975,N_11319);
or U12684 (N_12684,N_10568,N_11439);
nor U12685 (N_12685,N_10024,N_10354);
nor U12686 (N_12686,N_10042,N_11507);
and U12687 (N_12687,N_11112,N_11581);
xnor U12688 (N_12688,N_10639,N_11330);
and U12689 (N_12689,N_11226,N_11732);
xnor U12690 (N_12690,N_11924,N_10436);
and U12691 (N_12691,N_11032,N_10953);
nor U12692 (N_12692,N_10785,N_10679);
nand U12693 (N_12693,N_11775,N_10070);
and U12694 (N_12694,N_10276,N_11349);
nand U12695 (N_12695,N_11762,N_10613);
nor U12696 (N_12696,N_10290,N_10931);
and U12697 (N_12697,N_10773,N_10415);
and U12698 (N_12698,N_10310,N_11399);
or U12699 (N_12699,N_11761,N_10326);
nor U12700 (N_12700,N_11863,N_10174);
xnor U12701 (N_12701,N_11958,N_11068);
or U12702 (N_12702,N_10329,N_11442);
nor U12703 (N_12703,N_10069,N_11050);
nand U12704 (N_12704,N_10940,N_10309);
xnor U12705 (N_12705,N_11868,N_11321);
nand U12706 (N_12706,N_10107,N_10986);
nor U12707 (N_12707,N_10373,N_11189);
nand U12708 (N_12708,N_11200,N_11217);
or U12709 (N_12709,N_11002,N_10971);
or U12710 (N_12710,N_11157,N_10787);
nor U12711 (N_12711,N_11735,N_11832);
nor U12712 (N_12712,N_10376,N_11968);
nor U12713 (N_12713,N_10061,N_11963);
or U12714 (N_12714,N_10126,N_10668);
xor U12715 (N_12715,N_10305,N_11072);
or U12716 (N_12716,N_10802,N_10651);
and U12717 (N_12717,N_11540,N_10424);
and U12718 (N_12718,N_11128,N_11326);
xor U12719 (N_12719,N_11454,N_11262);
or U12720 (N_12720,N_10129,N_10969);
and U12721 (N_12721,N_11372,N_10028);
nand U12722 (N_12722,N_10548,N_10935);
nand U12723 (N_12723,N_11269,N_11962);
xnor U12724 (N_12724,N_10623,N_10122);
and U12725 (N_12725,N_11165,N_11737);
nand U12726 (N_12726,N_11944,N_10029);
and U12727 (N_12727,N_10121,N_11437);
xnor U12728 (N_12728,N_11703,N_11780);
or U12729 (N_12729,N_10911,N_10674);
nor U12730 (N_12730,N_10712,N_10741);
or U12731 (N_12731,N_10693,N_10489);
nand U12732 (N_12732,N_10761,N_10417);
and U12733 (N_12733,N_10486,N_11252);
or U12734 (N_12734,N_11320,N_11721);
or U12735 (N_12735,N_11127,N_10615);
nand U12736 (N_12736,N_10018,N_10716);
xnor U12737 (N_12737,N_10919,N_11317);
or U12738 (N_12738,N_10767,N_11985);
nand U12739 (N_12739,N_10861,N_10076);
and U12740 (N_12740,N_10831,N_11558);
and U12741 (N_12741,N_11070,N_10439);
or U12742 (N_12742,N_10156,N_11324);
xor U12743 (N_12743,N_10325,N_10866);
and U12744 (N_12744,N_11797,N_11198);
and U12745 (N_12745,N_10763,N_11095);
xor U12746 (N_12746,N_11170,N_10421);
or U12747 (N_12747,N_11092,N_11310);
nand U12748 (N_12748,N_10384,N_10973);
nand U12749 (N_12749,N_11510,N_10382);
nor U12750 (N_12750,N_11843,N_10676);
nand U12751 (N_12751,N_10775,N_10776);
or U12752 (N_12752,N_10996,N_11839);
nor U12753 (N_12753,N_10034,N_10809);
xnor U12754 (N_12754,N_10128,N_11059);
nand U12755 (N_12755,N_11624,N_10375);
and U12756 (N_12756,N_11281,N_11808);
nand U12757 (N_12757,N_11396,N_11381);
and U12758 (N_12758,N_10002,N_10315);
nor U12759 (N_12759,N_11709,N_11713);
nor U12760 (N_12760,N_10627,N_11039);
or U12761 (N_12761,N_10260,N_10418);
or U12762 (N_12762,N_11038,N_11611);
xor U12763 (N_12763,N_10643,N_10405);
or U12764 (N_12764,N_11042,N_11743);
nor U12765 (N_12765,N_10198,N_10046);
nor U12766 (N_12766,N_11238,N_10498);
or U12767 (N_12767,N_11526,N_10444);
xnor U12768 (N_12768,N_11368,N_11554);
and U12769 (N_12769,N_11559,N_10078);
nor U12770 (N_12770,N_11416,N_11220);
or U12771 (N_12771,N_11594,N_11224);
xor U12772 (N_12772,N_10702,N_11191);
and U12773 (N_12773,N_11662,N_10187);
nor U12774 (N_12774,N_11763,N_10867);
or U12775 (N_12775,N_11401,N_10286);
xor U12776 (N_12776,N_11845,N_11567);
nor U12777 (N_12777,N_10990,N_10642);
nor U12778 (N_12778,N_10751,N_10594);
nor U12779 (N_12779,N_10694,N_10587);
xor U12780 (N_12780,N_11014,N_10998);
nor U12781 (N_12781,N_11185,N_11461);
xnor U12782 (N_12782,N_11147,N_10355);
xor U12783 (N_12783,N_11472,N_10488);
or U12784 (N_12784,N_10361,N_11254);
or U12785 (N_12785,N_11411,N_10254);
and U12786 (N_12786,N_11696,N_11840);
xnor U12787 (N_12787,N_11000,N_11817);
or U12788 (N_12788,N_10349,N_11177);
nor U12789 (N_12789,N_10507,N_11151);
xor U12790 (N_12790,N_10168,N_11216);
and U12791 (N_12791,N_11047,N_10412);
nor U12792 (N_12792,N_11378,N_11542);
or U12793 (N_12793,N_11682,N_11413);
nand U12794 (N_12794,N_11888,N_10823);
nor U12795 (N_12795,N_11277,N_11500);
or U12796 (N_12796,N_11299,N_10433);
and U12797 (N_12797,N_10782,N_10103);
nand U12798 (N_12798,N_10106,N_11344);
nand U12799 (N_12799,N_11466,N_11410);
xnor U12800 (N_12800,N_10267,N_11619);
xor U12801 (N_12801,N_10884,N_11828);
nor U12802 (N_12802,N_11612,N_10110);
nor U12803 (N_12803,N_10557,N_11404);
or U12804 (N_12804,N_11316,N_10410);
nor U12805 (N_12805,N_10735,N_11417);
nand U12806 (N_12806,N_11397,N_11130);
nand U12807 (N_12807,N_10917,N_11998);
nor U12808 (N_12808,N_10274,N_11086);
xor U12809 (N_12809,N_10176,N_10721);
and U12810 (N_12810,N_11815,N_10328);
or U12811 (N_12811,N_11040,N_10119);
or U12812 (N_12812,N_10670,N_10795);
or U12813 (N_12813,N_10578,N_11137);
xor U12814 (N_12814,N_11833,N_11084);
xnor U12815 (N_12815,N_11892,N_11273);
and U12816 (N_12816,N_10992,N_10342);
and U12817 (N_12817,N_11445,N_10801);
or U12818 (N_12818,N_10036,N_10209);
nand U12819 (N_12819,N_11327,N_11400);
xnor U12820 (N_12820,N_10337,N_10021);
xnor U12821 (N_12821,N_11323,N_10234);
and U12822 (N_12822,N_10275,N_10585);
or U12823 (N_12823,N_10652,N_10832);
xor U12824 (N_12824,N_11627,N_10031);
nand U12825 (N_12825,N_10673,N_10989);
nor U12826 (N_12826,N_10936,N_11131);
and U12827 (N_12827,N_10941,N_11545);
nor U12828 (N_12828,N_11161,N_11188);
nand U12829 (N_12829,N_11883,N_10859);
nand U12830 (N_12830,N_11361,N_10492);
nor U12831 (N_12831,N_11926,N_11676);
nor U12832 (N_12832,N_10665,N_10317);
xor U12833 (N_12833,N_11586,N_10812);
or U12834 (N_12834,N_11672,N_10017);
or U12835 (N_12835,N_11209,N_11708);
nor U12836 (N_12836,N_10839,N_10518);
nor U12837 (N_12837,N_11765,N_10991);
xor U12838 (N_12838,N_10362,N_10840);
and U12839 (N_12839,N_10725,N_10108);
xor U12840 (N_12840,N_10793,N_11100);
and U12841 (N_12841,N_10822,N_11003);
nand U12842 (N_12842,N_10689,N_11996);
nand U12843 (N_12843,N_10456,N_10576);
nand U12844 (N_12844,N_10170,N_10370);
and U12845 (N_12845,N_11898,N_10402);
or U12846 (N_12846,N_10663,N_10237);
or U12847 (N_12847,N_11295,N_11571);
xnor U12848 (N_12848,N_10655,N_10865);
xnor U12849 (N_12849,N_10153,N_11991);
or U12850 (N_12850,N_11318,N_11541);
and U12851 (N_12851,N_11647,N_10805);
and U12852 (N_12852,N_10257,N_10130);
xnor U12853 (N_12853,N_10047,N_10925);
nand U12854 (N_12854,N_11512,N_10928);
xor U12855 (N_12855,N_10161,N_10522);
or U12856 (N_12856,N_11745,N_11847);
and U12857 (N_12857,N_10880,N_11495);
nand U12858 (N_12858,N_10797,N_10810);
and U12859 (N_12859,N_10703,N_11036);
nand U12860 (N_12860,N_10269,N_10877);
or U12861 (N_12861,N_11267,N_10096);
nor U12862 (N_12862,N_10535,N_11497);
xor U12863 (N_12863,N_11448,N_10894);
and U12864 (N_12864,N_10737,N_11785);
or U12865 (N_12865,N_11123,N_10944);
xor U12866 (N_12866,N_11767,N_10228);
and U12867 (N_12867,N_10235,N_11103);
nand U12868 (N_12868,N_10963,N_10811);
or U12869 (N_12869,N_10479,N_10533);
xor U12870 (N_12870,N_11925,N_11806);
nor U12871 (N_12871,N_11738,N_11250);
nor U12872 (N_12872,N_11447,N_11392);
xnor U12873 (N_12873,N_11740,N_11212);
and U12874 (N_12874,N_10937,N_11290);
or U12875 (N_12875,N_11044,N_10434);
xor U12876 (N_12876,N_11491,N_11474);
nor U12877 (N_12877,N_10332,N_11384);
xnor U12878 (N_12878,N_11664,N_10628);
and U12879 (N_12879,N_11336,N_11153);
xnor U12880 (N_12880,N_11771,N_11122);
nand U12881 (N_12881,N_11965,N_10934);
xnor U12882 (N_12882,N_11728,N_11779);
nor U12883 (N_12883,N_10131,N_10449);
nor U12884 (N_12884,N_10573,N_11788);
and U12885 (N_12885,N_10041,N_10927);
nand U12886 (N_12886,N_11587,N_10825);
nor U12887 (N_12887,N_11509,N_11995);
or U12888 (N_12888,N_10146,N_10287);
or U12889 (N_12889,N_11716,N_10532);
nor U12890 (N_12890,N_10902,N_11471);
nand U12891 (N_12891,N_10386,N_11769);
nand U12892 (N_12892,N_11113,N_11517);
xor U12893 (N_12893,N_11149,N_11658);
nand U12894 (N_12894,N_11687,N_10245);
nand U12895 (N_12895,N_11948,N_11511);
xor U12896 (N_12896,N_11506,N_10644);
nand U12897 (N_12897,N_10495,N_11458);
nor U12898 (N_12898,N_11910,N_11714);
nor U12899 (N_12899,N_10459,N_10490);
nor U12900 (N_12900,N_11111,N_10852);
or U12901 (N_12901,N_10055,N_11609);
or U12902 (N_12902,N_10743,N_11348);
and U12903 (N_12903,N_10318,N_10988);
nand U12904 (N_12904,N_10306,N_10133);
or U12905 (N_12905,N_10524,N_11213);
xor U12906 (N_12906,N_11580,N_10748);
xor U12907 (N_12907,N_11593,N_10929);
nand U12908 (N_12908,N_11006,N_10547);
xor U12909 (N_12909,N_10404,N_10010);
xor U12910 (N_12910,N_10733,N_10647);
or U12911 (N_12911,N_11674,N_10019);
nor U12912 (N_12912,N_10206,N_10516);
nor U12913 (N_12913,N_10437,N_10976);
nand U12914 (N_12914,N_11872,N_10049);
or U12915 (N_12915,N_11309,N_11707);
nand U12916 (N_12916,N_10572,N_10208);
nand U12917 (N_12917,N_11755,N_10660);
nor U12918 (N_12918,N_10199,N_11992);
nand U12919 (N_12919,N_10182,N_11364);
nand U12920 (N_12920,N_10044,N_11947);
nand U12921 (N_12921,N_10324,N_10951);
nand U12922 (N_12922,N_11784,N_11347);
nand U12923 (N_12923,N_11742,N_10923);
nand U12924 (N_12924,N_10580,N_10466);
and U12925 (N_12925,N_11975,N_10836);
and U12926 (N_12926,N_10372,N_10215);
and U12927 (N_12927,N_11631,N_11719);
nor U12928 (N_12928,N_10943,N_10394);
nor U12929 (N_12929,N_11938,N_11218);
and U12930 (N_12930,N_11104,N_11242);
nand U12931 (N_12931,N_10497,N_10427);
nor U12932 (N_12932,N_11750,N_11688);
nand U12933 (N_12933,N_11602,N_11980);
xor U12934 (N_12934,N_11066,N_10521);
and U12935 (N_12935,N_10715,N_10202);
or U12936 (N_12936,N_10338,N_11523);
nand U12937 (N_12937,N_11387,N_11945);
or U12938 (N_12938,N_11081,N_10039);
nor U12939 (N_12939,N_11434,N_11476);
or U12940 (N_12940,N_11034,N_10446);
and U12941 (N_12941,N_10564,N_11064);
or U12942 (N_12942,N_10705,N_10360);
nor U12943 (N_12943,N_11906,N_10571);
xnor U12944 (N_12944,N_11480,N_10634);
or U12945 (N_12945,N_10611,N_10271);
and U12946 (N_12946,N_11125,N_10092);
or U12947 (N_12947,N_10954,N_11301);
xnor U12948 (N_12948,N_11155,N_11490);
nor U12949 (N_12949,N_11067,N_11118);
or U12950 (N_12950,N_10004,N_10536);
xor U12951 (N_12951,N_11977,N_10463);
xor U12952 (N_12952,N_11547,N_11457);
xor U12953 (N_12953,N_10913,N_10282);
or U12954 (N_12954,N_10472,N_11934);
nand U12955 (N_12955,N_10407,N_11525);
nor U12956 (N_12956,N_10566,N_10697);
or U12957 (N_12957,N_11940,N_11885);
nor U12958 (N_12958,N_10339,N_10843);
xor U12959 (N_12959,N_11043,N_11990);
nor U12960 (N_12960,N_10316,N_11951);
nor U12961 (N_12961,N_11374,N_11222);
xor U12962 (N_12962,N_10137,N_10744);
xor U12963 (N_12963,N_10084,N_10453);
and U12964 (N_12964,N_11073,N_11928);
or U12965 (N_12965,N_10167,N_11634);
or U12966 (N_12966,N_11856,N_10431);
and U12967 (N_12967,N_10060,N_11974);
nor U12968 (N_12968,N_10435,N_10026);
and U12969 (N_12969,N_11989,N_11603);
and U12970 (N_12970,N_10223,N_10500);
and U12971 (N_12971,N_11010,N_10792);
nor U12972 (N_12972,N_10722,N_11894);
or U12973 (N_12973,N_10622,N_11724);
xor U12974 (N_12974,N_10646,N_10530);
nand U12975 (N_12975,N_11692,N_10688);
xnor U12976 (N_12976,N_11117,N_10225);
and U12977 (N_12977,N_10419,N_11452);
nor U12978 (N_12978,N_10554,N_10952);
nand U12979 (N_12979,N_11648,N_11124);
nor U12980 (N_12980,N_11395,N_11757);
nand U12981 (N_12981,N_11484,N_11667);
and U12982 (N_12982,N_10333,N_11121);
nand U12983 (N_12983,N_11120,N_11823);
nand U12984 (N_12984,N_11390,N_10892);
xnor U12985 (N_12985,N_11470,N_11641);
nand U12986 (N_12986,N_11078,N_11576);
nor U12987 (N_12987,N_10672,N_11802);
or U12988 (N_12988,N_10065,N_11734);
or U12989 (N_12989,N_11812,N_10794);
and U12990 (N_12990,N_11264,N_11786);
or U12991 (N_12991,N_10423,N_10214);
nand U12992 (N_12992,N_11236,N_10016);
nor U12993 (N_12993,N_11834,N_11681);
nand U12994 (N_12994,N_10231,N_11077);
nor U12995 (N_12995,N_10631,N_10172);
xor U12996 (N_12996,N_11228,N_10210);
and U12997 (N_12997,N_10964,N_10749);
nand U12998 (N_12998,N_11503,N_11271);
xor U12999 (N_12999,N_11333,N_10440);
and U13000 (N_13000,N_10420,N_10147);
or U13001 (N_13001,N_11717,N_10636);
xor U13002 (N_13002,N_10928,N_11112);
nor U13003 (N_13003,N_10170,N_10107);
nor U13004 (N_13004,N_10056,N_11889);
or U13005 (N_13005,N_10636,N_10262);
nor U13006 (N_13006,N_10444,N_10010);
and U13007 (N_13007,N_11802,N_10588);
nor U13008 (N_13008,N_10720,N_10194);
and U13009 (N_13009,N_11443,N_10329);
or U13010 (N_13010,N_11408,N_10820);
and U13011 (N_13011,N_10992,N_11143);
and U13012 (N_13012,N_11690,N_11647);
nand U13013 (N_13013,N_11495,N_11863);
or U13014 (N_13014,N_11595,N_10425);
and U13015 (N_13015,N_11165,N_11118);
nand U13016 (N_13016,N_10193,N_10404);
and U13017 (N_13017,N_11489,N_11805);
xnor U13018 (N_13018,N_11178,N_11097);
nor U13019 (N_13019,N_11358,N_10305);
nor U13020 (N_13020,N_11956,N_11547);
xor U13021 (N_13021,N_10204,N_11913);
nor U13022 (N_13022,N_11800,N_10150);
xor U13023 (N_13023,N_10366,N_11263);
xnor U13024 (N_13024,N_10579,N_10299);
nand U13025 (N_13025,N_11329,N_11358);
xnor U13026 (N_13026,N_11947,N_10506);
nor U13027 (N_13027,N_11325,N_11561);
or U13028 (N_13028,N_10941,N_10133);
nand U13029 (N_13029,N_10137,N_10471);
xor U13030 (N_13030,N_11663,N_11977);
nand U13031 (N_13031,N_11119,N_11604);
nand U13032 (N_13032,N_11976,N_10782);
nand U13033 (N_13033,N_10645,N_11989);
nor U13034 (N_13034,N_11224,N_11113);
or U13035 (N_13035,N_10197,N_10668);
nand U13036 (N_13036,N_10068,N_11083);
xor U13037 (N_13037,N_10385,N_11167);
and U13038 (N_13038,N_10939,N_10208);
nor U13039 (N_13039,N_11782,N_11238);
nand U13040 (N_13040,N_11797,N_11749);
nor U13041 (N_13041,N_10474,N_11472);
nor U13042 (N_13042,N_10535,N_11901);
and U13043 (N_13043,N_10059,N_10394);
or U13044 (N_13044,N_10258,N_10869);
nand U13045 (N_13045,N_11797,N_10216);
nand U13046 (N_13046,N_11236,N_11634);
nand U13047 (N_13047,N_10133,N_11335);
nor U13048 (N_13048,N_11614,N_10448);
and U13049 (N_13049,N_11235,N_10616);
nor U13050 (N_13050,N_10268,N_10398);
nor U13051 (N_13051,N_10657,N_10630);
or U13052 (N_13052,N_10196,N_11038);
or U13053 (N_13053,N_11123,N_11550);
xnor U13054 (N_13054,N_10733,N_11381);
xnor U13055 (N_13055,N_11949,N_10920);
or U13056 (N_13056,N_11475,N_10506);
nand U13057 (N_13057,N_10408,N_11634);
and U13058 (N_13058,N_10916,N_10468);
and U13059 (N_13059,N_10082,N_11155);
nor U13060 (N_13060,N_10808,N_11136);
nor U13061 (N_13061,N_11416,N_10637);
nand U13062 (N_13062,N_10267,N_10336);
nand U13063 (N_13063,N_10325,N_10742);
xnor U13064 (N_13064,N_10344,N_11237);
and U13065 (N_13065,N_11973,N_11877);
nor U13066 (N_13066,N_11392,N_10476);
or U13067 (N_13067,N_11863,N_10677);
xor U13068 (N_13068,N_11194,N_11498);
nor U13069 (N_13069,N_11517,N_11697);
or U13070 (N_13070,N_10553,N_10618);
nor U13071 (N_13071,N_10046,N_11359);
and U13072 (N_13072,N_11869,N_10542);
nand U13073 (N_13073,N_10324,N_10050);
nor U13074 (N_13074,N_11724,N_11509);
or U13075 (N_13075,N_10015,N_11226);
nand U13076 (N_13076,N_10039,N_10265);
xor U13077 (N_13077,N_11616,N_10298);
nand U13078 (N_13078,N_11620,N_10675);
nor U13079 (N_13079,N_10529,N_11076);
nand U13080 (N_13080,N_11370,N_10600);
nor U13081 (N_13081,N_10690,N_11191);
or U13082 (N_13082,N_10356,N_10603);
nor U13083 (N_13083,N_10312,N_11487);
or U13084 (N_13084,N_10093,N_11765);
and U13085 (N_13085,N_10083,N_10252);
or U13086 (N_13086,N_10108,N_11429);
or U13087 (N_13087,N_10305,N_10793);
xnor U13088 (N_13088,N_10218,N_10590);
or U13089 (N_13089,N_10862,N_11918);
nand U13090 (N_13090,N_10856,N_11796);
and U13091 (N_13091,N_10202,N_10637);
nand U13092 (N_13092,N_10803,N_10497);
nand U13093 (N_13093,N_10592,N_10967);
nor U13094 (N_13094,N_11034,N_10680);
nor U13095 (N_13095,N_10892,N_10552);
xor U13096 (N_13096,N_10452,N_10491);
nand U13097 (N_13097,N_10440,N_10558);
xor U13098 (N_13098,N_11335,N_11971);
or U13099 (N_13099,N_10589,N_11152);
or U13100 (N_13100,N_10530,N_10754);
and U13101 (N_13101,N_10695,N_10243);
or U13102 (N_13102,N_11697,N_11658);
nor U13103 (N_13103,N_10644,N_10007);
xor U13104 (N_13104,N_10699,N_11517);
or U13105 (N_13105,N_10859,N_10619);
xor U13106 (N_13106,N_10386,N_10425);
nor U13107 (N_13107,N_11195,N_11930);
xor U13108 (N_13108,N_11093,N_10630);
xor U13109 (N_13109,N_10476,N_11492);
xnor U13110 (N_13110,N_11283,N_10815);
xor U13111 (N_13111,N_11833,N_11118);
xor U13112 (N_13112,N_11141,N_10416);
nor U13113 (N_13113,N_10504,N_10118);
and U13114 (N_13114,N_10713,N_10513);
nor U13115 (N_13115,N_10483,N_11367);
nor U13116 (N_13116,N_10947,N_11982);
xor U13117 (N_13117,N_10095,N_10037);
or U13118 (N_13118,N_10947,N_10558);
nor U13119 (N_13119,N_11455,N_10057);
or U13120 (N_13120,N_10863,N_10039);
nand U13121 (N_13121,N_10081,N_10970);
nor U13122 (N_13122,N_11787,N_10543);
xor U13123 (N_13123,N_10959,N_10691);
and U13124 (N_13124,N_10325,N_10404);
and U13125 (N_13125,N_11744,N_11524);
nor U13126 (N_13126,N_11967,N_11890);
xor U13127 (N_13127,N_10856,N_10231);
nand U13128 (N_13128,N_10227,N_11345);
and U13129 (N_13129,N_11041,N_10958);
nand U13130 (N_13130,N_11054,N_11262);
and U13131 (N_13131,N_11056,N_10340);
xor U13132 (N_13132,N_10543,N_10808);
xor U13133 (N_13133,N_10436,N_11306);
or U13134 (N_13134,N_10405,N_10568);
and U13135 (N_13135,N_10366,N_10909);
nand U13136 (N_13136,N_11980,N_10596);
and U13137 (N_13137,N_11172,N_11213);
nand U13138 (N_13138,N_10309,N_11839);
xnor U13139 (N_13139,N_11984,N_10559);
xnor U13140 (N_13140,N_11977,N_10457);
xor U13141 (N_13141,N_11602,N_10742);
xnor U13142 (N_13142,N_10309,N_11567);
nand U13143 (N_13143,N_11661,N_10408);
nand U13144 (N_13144,N_10086,N_11245);
and U13145 (N_13145,N_10950,N_11832);
xor U13146 (N_13146,N_11346,N_11482);
nor U13147 (N_13147,N_10902,N_11672);
or U13148 (N_13148,N_11593,N_11079);
or U13149 (N_13149,N_11728,N_11191);
xnor U13150 (N_13150,N_10588,N_11912);
xor U13151 (N_13151,N_11724,N_11204);
nand U13152 (N_13152,N_11427,N_10231);
xor U13153 (N_13153,N_10429,N_10603);
xnor U13154 (N_13154,N_10308,N_10694);
xnor U13155 (N_13155,N_11951,N_11631);
or U13156 (N_13156,N_10944,N_10346);
nand U13157 (N_13157,N_10415,N_10273);
or U13158 (N_13158,N_10193,N_10811);
and U13159 (N_13159,N_10584,N_10807);
or U13160 (N_13160,N_10702,N_10328);
xor U13161 (N_13161,N_10290,N_10142);
nor U13162 (N_13162,N_10736,N_10745);
and U13163 (N_13163,N_10718,N_11474);
and U13164 (N_13164,N_10014,N_10357);
nor U13165 (N_13165,N_10362,N_10796);
nand U13166 (N_13166,N_10071,N_11029);
nand U13167 (N_13167,N_11148,N_11156);
nand U13168 (N_13168,N_10464,N_10723);
or U13169 (N_13169,N_10001,N_10854);
or U13170 (N_13170,N_11591,N_10055);
nand U13171 (N_13171,N_10967,N_11680);
nand U13172 (N_13172,N_11422,N_10021);
or U13173 (N_13173,N_11211,N_11431);
nor U13174 (N_13174,N_10883,N_11821);
or U13175 (N_13175,N_11006,N_11983);
or U13176 (N_13176,N_11578,N_10086);
or U13177 (N_13177,N_10064,N_11551);
nor U13178 (N_13178,N_10761,N_10730);
nand U13179 (N_13179,N_10719,N_10523);
xnor U13180 (N_13180,N_10334,N_10305);
xnor U13181 (N_13181,N_11192,N_10085);
nand U13182 (N_13182,N_11564,N_11512);
nor U13183 (N_13183,N_10823,N_10296);
nor U13184 (N_13184,N_11993,N_11236);
or U13185 (N_13185,N_11220,N_10349);
and U13186 (N_13186,N_10758,N_11051);
and U13187 (N_13187,N_11171,N_10496);
nor U13188 (N_13188,N_10267,N_11452);
nor U13189 (N_13189,N_11373,N_11097);
xnor U13190 (N_13190,N_10052,N_10537);
nand U13191 (N_13191,N_11906,N_11239);
or U13192 (N_13192,N_11266,N_11764);
nand U13193 (N_13193,N_10305,N_10605);
or U13194 (N_13194,N_11218,N_11926);
and U13195 (N_13195,N_11470,N_10001);
xor U13196 (N_13196,N_11232,N_10407);
or U13197 (N_13197,N_11982,N_11411);
nand U13198 (N_13198,N_11160,N_10570);
and U13199 (N_13199,N_10899,N_10633);
or U13200 (N_13200,N_10739,N_11117);
and U13201 (N_13201,N_10820,N_11633);
nand U13202 (N_13202,N_11182,N_10718);
nand U13203 (N_13203,N_11324,N_11115);
nand U13204 (N_13204,N_11328,N_11172);
nor U13205 (N_13205,N_10212,N_10286);
nand U13206 (N_13206,N_10035,N_10070);
and U13207 (N_13207,N_11740,N_10101);
nand U13208 (N_13208,N_11544,N_10463);
or U13209 (N_13209,N_11860,N_10299);
xor U13210 (N_13210,N_11804,N_11199);
xnor U13211 (N_13211,N_11940,N_11723);
nand U13212 (N_13212,N_11263,N_11176);
nor U13213 (N_13213,N_11327,N_10140);
nor U13214 (N_13214,N_11765,N_10844);
nand U13215 (N_13215,N_10122,N_10718);
or U13216 (N_13216,N_10079,N_10312);
nor U13217 (N_13217,N_11264,N_10091);
nor U13218 (N_13218,N_11737,N_10893);
nand U13219 (N_13219,N_10648,N_10718);
xnor U13220 (N_13220,N_10964,N_11311);
xor U13221 (N_13221,N_10282,N_11666);
or U13222 (N_13222,N_10704,N_11210);
or U13223 (N_13223,N_10507,N_11416);
and U13224 (N_13224,N_10132,N_10221);
or U13225 (N_13225,N_10693,N_10868);
nand U13226 (N_13226,N_10773,N_10252);
and U13227 (N_13227,N_11357,N_10031);
or U13228 (N_13228,N_11192,N_10473);
nor U13229 (N_13229,N_10580,N_10977);
xnor U13230 (N_13230,N_10973,N_10894);
or U13231 (N_13231,N_11554,N_10314);
and U13232 (N_13232,N_11265,N_11311);
or U13233 (N_13233,N_10084,N_10975);
nor U13234 (N_13234,N_11862,N_10458);
and U13235 (N_13235,N_10331,N_11084);
nand U13236 (N_13236,N_11374,N_11408);
nor U13237 (N_13237,N_11294,N_10569);
xnor U13238 (N_13238,N_10940,N_10126);
xor U13239 (N_13239,N_10594,N_10981);
nand U13240 (N_13240,N_10460,N_11597);
or U13241 (N_13241,N_10374,N_11036);
nor U13242 (N_13242,N_11071,N_10239);
or U13243 (N_13243,N_11494,N_11948);
or U13244 (N_13244,N_10402,N_10603);
nand U13245 (N_13245,N_10100,N_11958);
and U13246 (N_13246,N_10131,N_11231);
and U13247 (N_13247,N_10144,N_11746);
and U13248 (N_13248,N_11207,N_11003);
and U13249 (N_13249,N_11437,N_10593);
and U13250 (N_13250,N_11423,N_11085);
and U13251 (N_13251,N_11181,N_11732);
nand U13252 (N_13252,N_10116,N_11937);
or U13253 (N_13253,N_11388,N_11714);
nor U13254 (N_13254,N_10004,N_10960);
nor U13255 (N_13255,N_11703,N_10686);
xnor U13256 (N_13256,N_10100,N_11963);
xor U13257 (N_13257,N_11244,N_11718);
and U13258 (N_13258,N_11705,N_11315);
nor U13259 (N_13259,N_10190,N_11129);
nand U13260 (N_13260,N_10649,N_11455);
or U13261 (N_13261,N_10342,N_10418);
and U13262 (N_13262,N_10527,N_11812);
nor U13263 (N_13263,N_11957,N_10424);
nor U13264 (N_13264,N_11933,N_10243);
or U13265 (N_13265,N_10766,N_11323);
and U13266 (N_13266,N_11618,N_10350);
xor U13267 (N_13267,N_11255,N_11926);
or U13268 (N_13268,N_10236,N_10334);
nor U13269 (N_13269,N_11396,N_11780);
and U13270 (N_13270,N_10315,N_11128);
nor U13271 (N_13271,N_10416,N_10543);
nand U13272 (N_13272,N_10718,N_11327);
or U13273 (N_13273,N_11480,N_11102);
or U13274 (N_13274,N_11270,N_11471);
xor U13275 (N_13275,N_10996,N_10365);
nor U13276 (N_13276,N_11977,N_11178);
xnor U13277 (N_13277,N_11595,N_10069);
or U13278 (N_13278,N_10099,N_10010);
xor U13279 (N_13279,N_11711,N_10075);
or U13280 (N_13280,N_10717,N_11215);
nor U13281 (N_13281,N_10598,N_10603);
nand U13282 (N_13282,N_10158,N_11614);
xor U13283 (N_13283,N_11586,N_10457);
and U13284 (N_13284,N_10333,N_11247);
nand U13285 (N_13285,N_11392,N_10938);
or U13286 (N_13286,N_11009,N_11033);
or U13287 (N_13287,N_10407,N_11548);
nand U13288 (N_13288,N_10331,N_11076);
or U13289 (N_13289,N_11276,N_10629);
and U13290 (N_13290,N_10904,N_11583);
xnor U13291 (N_13291,N_11036,N_10948);
xnor U13292 (N_13292,N_11215,N_10136);
xnor U13293 (N_13293,N_10302,N_11552);
and U13294 (N_13294,N_11046,N_11601);
nor U13295 (N_13295,N_11872,N_11211);
nand U13296 (N_13296,N_10844,N_10412);
or U13297 (N_13297,N_10434,N_10626);
xor U13298 (N_13298,N_10658,N_10156);
and U13299 (N_13299,N_11953,N_10165);
and U13300 (N_13300,N_10091,N_10466);
nand U13301 (N_13301,N_11135,N_11480);
xor U13302 (N_13302,N_11106,N_10161);
nand U13303 (N_13303,N_11492,N_11633);
xor U13304 (N_13304,N_10090,N_10234);
and U13305 (N_13305,N_10630,N_10146);
nor U13306 (N_13306,N_11926,N_11064);
xor U13307 (N_13307,N_10297,N_10773);
nor U13308 (N_13308,N_11847,N_10665);
and U13309 (N_13309,N_11070,N_10259);
nor U13310 (N_13310,N_10032,N_10080);
nor U13311 (N_13311,N_10166,N_10197);
and U13312 (N_13312,N_10469,N_10359);
and U13313 (N_13313,N_11213,N_10579);
and U13314 (N_13314,N_11514,N_11086);
xor U13315 (N_13315,N_10243,N_11078);
or U13316 (N_13316,N_10899,N_10542);
nand U13317 (N_13317,N_10009,N_10984);
xnor U13318 (N_13318,N_10100,N_11778);
nand U13319 (N_13319,N_11753,N_11452);
and U13320 (N_13320,N_11391,N_11759);
nand U13321 (N_13321,N_10087,N_10927);
nand U13322 (N_13322,N_11150,N_11737);
or U13323 (N_13323,N_11988,N_10508);
xnor U13324 (N_13324,N_11318,N_10801);
xor U13325 (N_13325,N_11450,N_11299);
xor U13326 (N_13326,N_11372,N_11716);
nand U13327 (N_13327,N_11809,N_11049);
xnor U13328 (N_13328,N_11046,N_11945);
and U13329 (N_13329,N_11820,N_11062);
and U13330 (N_13330,N_11813,N_10582);
xor U13331 (N_13331,N_11766,N_11394);
nand U13332 (N_13332,N_11301,N_11052);
nand U13333 (N_13333,N_11939,N_10365);
and U13334 (N_13334,N_10898,N_11417);
nor U13335 (N_13335,N_10935,N_11064);
or U13336 (N_13336,N_10241,N_11198);
or U13337 (N_13337,N_11900,N_10047);
and U13338 (N_13338,N_10404,N_10308);
nor U13339 (N_13339,N_11127,N_11373);
or U13340 (N_13340,N_10847,N_11971);
and U13341 (N_13341,N_11820,N_11835);
xnor U13342 (N_13342,N_11502,N_10242);
nor U13343 (N_13343,N_11679,N_11243);
nor U13344 (N_13344,N_11711,N_10292);
and U13345 (N_13345,N_10117,N_11011);
xor U13346 (N_13346,N_10336,N_10695);
or U13347 (N_13347,N_11724,N_11808);
xor U13348 (N_13348,N_11032,N_10254);
nand U13349 (N_13349,N_10927,N_11230);
or U13350 (N_13350,N_11940,N_10835);
or U13351 (N_13351,N_10834,N_11396);
or U13352 (N_13352,N_10091,N_11016);
nor U13353 (N_13353,N_11220,N_11030);
or U13354 (N_13354,N_11255,N_11424);
nand U13355 (N_13355,N_11813,N_11322);
nor U13356 (N_13356,N_10223,N_11163);
and U13357 (N_13357,N_10445,N_10462);
nor U13358 (N_13358,N_11245,N_10963);
or U13359 (N_13359,N_10320,N_11718);
nand U13360 (N_13360,N_11131,N_11643);
and U13361 (N_13361,N_11483,N_11469);
xnor U13362 (N_13362,N_11173,N_10883);
nor U13363 (N_13363,N_11257,N_11080);
and U13364 (N_13364,N_10100,N_10017);
or U13365 (N_13365,N_10430,N_11762);
and U13366 (N_13366,N_11501,N_10091);
nor U13367 (N_13367,N_11418,N_10170);
xor U13368 (N_13368,N_10183,N_10353);
nor U13369 (N_13369,N_10674,N_11676);
or U13370 (N_13370,N_11336,N_11663);
or U13371 (N_13371,N_10717,N_10658);
nand U13372 (N_13372,N_10504,N_11939);
nand U13373 (N_13373,N_10719,N_11566);
nor U13374 (N_13374,N_10078,N_11353);
or U13375 (N_13375,N_10342,N_10907);
and U13376 (N_13376,N_10527,N_11406);
nor U13377 (N_13377,N_10299,N_10692);
nor U13378 (N_13378,N_10889,N_11043);
nor U13379 (N_13379,N_11453,N_11790);
nor U13380 (N_13380,N_11264,N_11580);
xnor U13381 (N_13381,N_11204,N_10297);
and U13382 (N_13382,N_10702,N_10106);
or U13383 (N_13383,N_10805,N_10538);
and U13384 (N_13384,N_10394,N_11030);
nand U13385 (N_13385,N_10385,N_11750);
and U13386 (N_13386,N_10515,N_10001);
xnor U13387 (N_13387,N_11103,N_10605);
nand U13388 (N_13388,N_10828,N_11708);
nor U13389 (N_13389,N_11001,N_10172);
or U13390 (N_13390,N_11330,N_11640);
xor U13391 (N_13391,N_10270,N_11505);
and U13392 (N_13392,N_11572,N_11381);
and U13393 (N_13393,N_10801,N_11268);
xnor U13394 (N_13394,N_11074,N_11527);
nand U13395 (N_13395,N_10951,N_10407);
xor U13396 (N_13396,N_10437,N_11584);
and U13397 (N_13397,N_10159,N_10548);
nand U13398 (N_13398,N_11353,N_11721);
nand U13399 (N_13399,N_11380,N_11120);
or U13400 (N_13400,N_11012,N_11951);
and U13401 (N_13401,N_11825,N_10504);
xor U13402 (N_13402,N_11143,N_11494);
nand U13403 (N_13403,N_10261,N_10237);
and U13404 (N_13404,N_10875,N_11083);
nor U13405 (N_13405,N_10996,N_11920);
or U13406 (N_13406,N_10804,N_11492);
or U13407 (N_13407,N_10920,N_10342);
or U13408 (N_13408,N_11122,N_11195);
nand U13409 (N_13409,N_10624,N_11843);
or U13410 (N_13410,N_11945,N_10225);
or U13411 (N_13411,N_10869,N_11095);
or U13412 (N_13412,N_10127,N_10707);
nand U13413 (N_13413,N_11970,N_10869);
nor U13414 (N_13414,N_10244,N_10346);
or U13415 (N_13415,N_11112,N_11374);
nor U13416 (N_13416,N_10539,N_11537);
and U13417 (N_13417,N_11413,N_11403);
or U13418 (N_13418,N_10145,N_10938);
xnor U13419 (N_13419,N_11567,N_10164);
nor U13420 (N_13420,N_11593,N_10735);
nor U13421 (N_13421,N_11225,N_11069);
nor U13422 (N_13422,N_11948,N_11128);
and U13423 (N_13423,N_10217,N_11738);
or U13424 (N_13424,N_10058,N_11564);
or U13425 (N_13425,N_10318,N_11266);
nor U13426 (N_13426,N_11462,N_11081);
nand U13427 (N_13427,N_10538,N_10833);
nor U13428 (N_13428,N_10970,N_11572);
nor U13429 (N_13429,N_11579,N_11967);
and U13430 (N_13430,N_10730,N_11191);
xor U13431 (N_13431,N_10154,N_10253);
or U13432 (N_13432,N_10392,N_10651);
nand U13433 (N_13433,N_11908,N_11552);
and U13434 (N_13434,N_10090,N_10656);
and U13435 (N_13435,N_10117,N_11606);
nor U13436 (N_13436,N_10825,N_10421);
and U13437 (N_13437,N_11753,N_10814);
xor U13438 (N_13438,N_10031,N_10486);
and U13439 (N_13439,N_10142,N_11145);
or U13440 (N_13440,N_11032,N_11447);
or U13441 (N_13441,N_11417,N_10119);
or U13442 (N_13442,N_10359,N_11378);
nand U13443 (N_13443,N_11647,N_10397);
or U13444 (N_13444,N_11859,N_10965);
nor U13445 (N_13445,N_10211,N_10478);
xnor U13446 (N_13446,N_10872,N_11057);
nor U13447 (N_13447,N_11683,N_10876);
and U13448 (N_13448,N_10796,N_10655);
nor U13449 (N_13449,N_10357,N_11773);
nor U13450 (N_13450,N_10968,N_10357);
and U13451 (N_13451,N_11478,N_10596);
or U13452 (N_13452,N_10750,N_10943);
xor U13453 (N_13453,N_11727,N_11264);
nor U13454 (N_13454,N_10325,N_10966);
xnor U13455 (N_13455,N_10715,N_10188);
nor U13456 (N_13456,N_11405,N_10306);
and U13457 (N_13457,N_10102,N_11603);
and U13458 (N_13458,N_11790,N_10411);
or U13459 (N_13459,N_11109,N_11661);
and U13460 (N_13460,N_10044,N_10473);
or U13461 (N_13461,N_10830,N_10107);
xnor U13462 (N_13462,N_11703,N_10907);
xor U13463 (N_13463,N_10127,N_11535);
and U13464 (N_13464,N_11722,N_11367);
and U13465 (N_13465,N_11199,N_11113);
and U13466 (N_13466,N_11962,N_10678);
xor U13467 (N_13467,N_10596,N_11535);
nand U13468 (N_13468,N_10386,N_11152);
xnor U13469 (N_13469,N_11321,N_10517);
xor U13470 (N_13470,N_10551,N_10070);
or U13471 (N_13471,N_11312,N_11435);
xnor U13472 (N_13472,N_11110,N_11619);
nand U13473 (N_13473,N_10369,N_11968);
nand U13474 (N_13474,N_11717,N_10428);
and U13475 (N_13475,N_11155,N_10279);
or U13476 (N_13476,N_10481,N_10986);
nor U13477 (N_13477,N_11827,N_11394);
xor U13478 (N_13478,N_10942,N_11889);
or U13479 (N_13479,N_11866,N_11487);
or U13480 (N_13480,N_10028,N_11639);
nor U13481 (N_13481,N_10615,N_10358);
and U13482 (N_13482,N_11888,N_10265);
nor U13483 (N_13483,N_11918,N_10650);
or U13484 (N_13484,N_11582,N_11307);
nand U13485 (N_13485,N_11885,N_10391);
and U13486 (N_13486,N_10733,N_11945);
nand U13487 (N_13487,N_10061,N_10445);
nand U13488 (N_13488,N_10551,N_11448);
and U13489 (N_13489,N_11373,N_11140);
xor U13490 (N_13490,N_11282,N_10701);
and U13491 (N_13491,N_11900,N_11229);
or U13492 (N_13492,N_10576,N_10478);
nand U13493 (N_13493,N_11510,N_10087);
and U13494 (N_13494,N_11977,N_11180);
nor U13495 (N_13495,N_10072,N_11479);
and U13496 (N_13496,N_11251,N_11208);
and U13497 (N_13497,N_11141,N_10349);
nand U13498 (N_13498,N_11130,N_11975);
nor U13499 (N_13499,N_11187,N_10353);
and U13500 (N_13500,N_11163,N_11457);
xor U13501 (N_13501,N_11626,N_11987);
xnor U13502 (N_13502,N_11338,N_10221);
and U13503 (N_13503,N_10248,N_10103);
nor U13504 (N_13504,N_11875,N_10410);
and U13505 (N_13505,N_11988,N_11439);
nand U13506 (N_13506,N_10084,N_11730);
or U13507 (N_13507,N_10314,N_11391);
and U13508 (N_13508,N_10632,N_11314);
or U13509 (N_13509,N_10532,N_10979);
nor U13510 (N_13510,N_10897,N_10294);
xnor U13511 (N_13511,N_11093,N_10311);
and U13512 (N_13512,N_10453,N_11714);
or U13513 (N_13513,N_10271,N_11324);
and U13514 (N_13514,N_11449,N_11807);
xnor U13515 (N_13515,N_11675,N_10115);
or U13516 (N_13516,N_11934,N_11346);
or U13517 (N_13517,N_11229,N_11297);
xnor U13518 (N_13518,N_10705,N_10322);
nand U13519 (N_13519,N_10672,N_10818);
xor U13520 (N_13520,N_11289,N_10496);
xnor U13521 (N_13521,N_11727,N_11596);
nand U13522 (N_13522,N_10816,N_10824);
or U13523 (N_13523,N_10127,N_10202);
xor U13524 (N_13524,N_11717,N_10544);
nand U13525 (N_13525,N_10351,N_10157);
or U13526 (N_13526,N_11405,N_10424);
nand U13527 (N_13527,N_11808,N_10646);
nand U13528 (N_13528,N_11000,N_11737);
and U13529 (N_13529,N_11215,N_11213);
and U13530 (N_13530,N_11919,N_11163);
xnor U13531 (N_13531,N_10934,N_10102);
nand U13532 (N_13532,N_11080,N_10733);
xnor U13533 (N_13533,N_10235,N_10299);
nand U13534 (N_13534,N_11812,N_10863);
nor U13535 (N_13535,N_11651,N_11048);
or U13536 (N_13536,N_10515,N_11769);
xor U13537 (N_13537,N_11628,N_11532);
nand U13538 (N_13538,N_11780,N_11531);
nand U13539 (N_13539,N_11101,N_10200);
xor U13540 (N_13540,N_10008,N_10767);
and U13541 (N_13541,N_10467,N_11099);
and U13542 (N_13542,N_10414,N_10102);
xnor U13543 (N_13543,N_10902,N_10796);
xnor U13544 (N_13544,N_11855,N_11494);
or U13545 (N_13545,N_11445,N_10758);
or U13546 (N_13546,N_10902,N_10020);
or U13547 (N_13547,N_10089,N_11720);
xor U13548 (N_13548,N_10786,N_10469);
and U13549 (N_13549,N_10719,N_11048);
nor U13550 (N_13550,N_11882,N_10512);
or U13551 (N_13551,N_10693,N_10441);
nand U13552 (N_13552,N_10225,N_11529);
or U13553 (N_13553,N_10607,N_11371);
nand U13554 (N_13554,N_11728,N_10992);
nand U13555 (N_13555,N_10946,N_11567);
nand U13556 (N_13556,N_11828,N_10495);
nor U13557 (N_13557,N_11608,N_11996);
nand U13558 (N_13558,N_10167,N_10807);
nor U13559 (N_13559,N_11745,N_10305);
nand U13560 (N_13560,N_10358,N_10186);
or U13561 (N_13561,N_10487,N_11860);
xnor U13562 (N_13562,N_11548,N_10628);
xnor U13563 (N_13563,N_11656,N_10096);
or U13564 (N_13564,N_10566,N_10852);
and U13565 (N_13565,N_10117,N_11350);
or U13566 (N_13566,N_11251,N_11996);
or U13567 (N_13567,N_10506,N_10048);
nor U13568 (N_13568,N_11709,N_10494);
xor U13569 (N_13569,N_10120,N_10725);
and U13570 (N_13570,N_10894,N_10954);
xor U13571 (N_13571,N_11177,N_11350);
xor U13572 (N_13572,N_11083,N_10158);
and U13573 (N_13573,N_10364,N_10103);
and U13574 (N_13574,N_11176,N_11853);
nand U13575 (N_13575,N_10572,N_11012);
or U13576 (N_13576,N_11818,N_11860);
and U13577 (N_13577,N_11177,N_11447);
or U13578 (N_13578,N_10757,N_11516);
and U13579 (N_13579,N_11782,N_10763);
nand U13580 (N_13580,N_10082,N_10430);
nand U13581 (N_13581,N_11592,N_11835);
nand U13582 (N_13582,N_11384,N_11778);
and U13583 (N_13583,N_10685,N_11254);
nor U13584 (N_13584,N_10281,N_10640);
nand U13585 (N_13585,N_11078,N_11449);
and U13586 (N_13586,N_10743,N_10967);
nand U13587 (N_13587,N_11245,N_11913);
xnor U13588 (N_13588,N_11621,N_11217);
nand U13589 (N_13589,N_11178,N_10012);
and U13590 (N_13590,N_10332,N_10474);
nor U13591 (N_13591,N_11397,N_11005);
nand U13592 (N_13592,N_10630,N_10430);
nor U13593 (N_13593,N_10831,N_10858);
and U13594 (N_13594,N_10329,N_11264);
nor U13595 (N_13595,N_10310,N_10018);
and U13596 (N_13596,N_10066,N_10059);
and U13597 (N_13597,N_10914,N_10198);
and U13598 (N_13598,N_10096,N_11529);
xnor U13599 (N_13599,N_11355,N_10942);
nor U13600 (N_13600,N_10563,N_10054);
nor U13601 (N_13601,N_10781,N_10995);
and U13602 (N_13602,N_10237,N_10785);
or U13603 (N_13603,N_11336,N_10677);
nor U13604 (N_13604,N_10997,N_10612);
xnor U13605 (N_13605,N_11666,N_10538);
and U13606 (N_13606,N_10539,N_10411);
nor U13607 (N_13607,N_11170,N_11678);
or U13608 (N_13608,N_10090,N_11307);
nor U13609 (N_13609,N_11266,N_10565);
or U13610 (N_13610,N_11849,N_10918);
xor U13611 (N_13611,N_11787,N_11061);
and U13612 (N_13612,N_10830,N_11155);
xor U13613 (N_13613,N_11918,N_10462);
and U13614 (N_13614,N_11727,N_10791);
nand U13615 (N_13615,N_11791,N_10277);
xor U13616 (N_13616,N_11004,N_11714);
and U13617 (N_13617,N_10736,N_11007);
nand U13618 (N_13618,N_11777,N_10707);
nor U13619 (N_13619,N_11841,N_10398);
nand U13620 (N_13620,N_10265,N_10235);
or U13621 (N_13621,N_10267,N_11626);
nor U13622 (N_13622,N_11974,N_11383);
nand U13623 (N_13623,N_10779,N_10419);
nor U13624 (N_13624,N_11674,N_10688);
xor U13625 (N_13625,N_10421,N_10666);
nand U13626 (N_13626,N_11747,N_11935);
nor U13627 (N_13627,N_10016,N_11231);
and U13628 (N_13628,N_10312,N_10409);
and U13629 (N_13629,N_11478,N_10270);
nor U13630 (N_13630,N_10226,N_11862);
xnor U13631 (N_13631,N_11286,N_11050);
and U13632 (N_13632,N_11218,N_10150);
xnor U13633 (N_13633,N_11637,N_10162);
nand U13634 (N_13634,N_10494,N_10610);
or U13635 (N_13635,N_10627,N_10340);
nor U13636 (N_13636,N_11559,N_10331);
or U13637 (N_13637,N_10370,N_11082);
nand U13638 (N_13638,N_10253,N_10992);
nand U13639 (N_13639,N_11728,N_11538);
xor U13640 (N_13640,N_10924,N_10207);
nor U13641 (N_13641,N_11762,N_11869);
nor U13642 (N_13642,N_10275,N_10323);
and U13643 (N_13643,N_10596,N_10224);
and U13644 (N_13644,N_10166,N_11704);
and U13645 (N_13645,N_11883,N_11038);
or U13646 (N_13646,N_10059,N_11856);
xnor U13647 (N_13647,N_10066,N_10524);
nand U13648 (N_13648,N_11344,N_11220);
xor U13649 (N_13649,N_10534,N_10997);
nor U13650 (N_13650,N_10439,N_10480);
nor U13651 (N_13651,N_11718,N_10021);
xor U13652 (N_13652,N_11190,N_11954);
or U13653 (N_13653,N_11533,N_11334);
nor U13654 (N_13654,N_10022,N_10450);
nand U13655 (N_13655,N_11024,N_10849);
or U13656 (N_13656,N_10023,N_11598);
nand U13657 (N_13657,N_11127,N_11183);
nand U13658 (N_13658,N_11453,N_11645);
and U13659 (N_13659,N_10964,N_11959);
xor U13660 (N_13660,N_10919,N_10921);
xor U13661 (N_13661,N_11697,N_10383);
nand U13662 (N_13662,N_11815,N_11727);
nor U13663 (N_13663,N_10535,N_11114);
xor U13664 (N_13664,N_11790,N_10677);
or U13665 (N_13665,N_11354,N_10814);
nand U13666 (N_13666,N_11034,N_10095);
xnor U13667 (N_13667,N_11171,N_10637);
nor U13668 (N_13668,N_11279,N_11240);
nor U13669 (N_13669,N_11623,N_10286);
nor U13670 (N_13670,N_11882,N_11519);
or U13671 (N_13671,N_10037,N_10083);
and U13672 (N_13672,N_10233,N_10800);
xnor U13673 (N_13673,N_10997,N_11598);
xor U13674 (N_13674,N_11695,N_10615);
and U13675 (N_13675,N_11678,N_10222);
and U13676 (N_13676,N_10997,N_11137);
xnor U13677 (N_13677,N_10165,N_10413);
and U13678 (N_13678,N_10247,N_10730);
nand U13679 (N_13679,N_10752,N_10146);
nor U13680 (N_13680,N_11451,N_11605);
and U13681 (N_13681,N_11179,N_10965);
nor U13682 (N_13682,N_10896,N_11811);
and U13683 (N_13683,N_11312,N_10656);
and U13684 (N_13684,N_11600,N_11517);
nand U13685 (N_13685,N_11535,N_11708);
and U13686 (N_13686,N_10039,N_10966);
and U13687 (N_13687,N_11090,N_10670);
nor U13688 (N_13688,N_11380,N_11125);
nand U13689 (N_13689,N_11296,N_11056);
and U13690 (N_13690,N_10870,N_10511);
and U13691 (N_13691,N_10170,N_10994);
or U13692 (N_13692,N_11343,N_11194);
nor U13693 (N_13693,N_10478,N_10257);
nand U13694 (N_13694,N_11196,N_11132);
or U13695 (N_13695,N_11151,N_10691);
or U13696 (N_13696,N_10023,N_10149);
xnor U13697 (N_13697,N_11167,N_10706);
nand U13698 (N_13698,N_10097,N_11447);
xnor U13699 (N_13699,N_10287,N_10512);
xnor U13700 (N_13700,N_10436,N_10037);
xor U13701 (N_13701,N_10655,N_10097);
nor U13702 (N_13702,N_10208,N_10729);
nand U13703 (N_13703,N_10073,N_11383);
or U13704 (N_13704,N_11339,N_11624);
xor U13705 (N_13705,N_11514,N_11573);
or U13706 (N_13706,N_11298,N_11138);
or U13707 (N_13707,N_10566,N_10161);
nor U13708 (N_13708,N_11334,N_10097);
xor U13709 (N_13709,N_10878,N_11124);
nand U13710 (N_13710,N_11140,N_10019);
and U13711 (N_13711,N_11724,N_10604);
and U13712 (N_13712,N_10874,N_11051);
and U13713 (N_13713,N_11391,N_10757);
nand U13714 (N_13714,N_10149,N_10221);
and U13715 (N_13715,N_11052,N_10975);
and U13716 (N_13716,N_10082,N_11351);
or U13717 (N_13717,N_10330,N_10482);
nor U13718 (N_13718,N_11482,N_10165);
nor U13719 (N_13719,N_11993,N_10997);
or U13720 (N_13720,N_11998,N_11405);
and U13721 (N_13721,N_11026,N_11580);
or U13722 (N_13722,N_11206,N_10030);
nand U13723 (N_13723,N_10161,N_10153);
or U13724 (N_13724,N_10491,N_10912);
and U13725 (N_13725,N_10402,N_10087);
nor U13726 (N_13726,N_11848,N_10472);
and U13727 (N_13727,N_10614,N_10748);
nand U13728 (N_13728,N_10299,N_10553);
nor U13729 (N_13729,N_10540,N_10226);
nor U13730 (N_13730,N_11561,N_10258);
xnor U13731 (N_13731,N_11162,N_11178);
nand U13732 (N_13732,N_10322,N_10034);
nand U13733 (N_13733,N_10635,N_10237);
or U13734 (N_13734,N_10407,N_10250);
nor U13735 (N_13735,N_11037,N_10233);
nor U13736 (N_13736,N_10358,N_11731);
nand U13737 (N_13737,N_10937,N_10619);
nor U13738 (N_13738,N_10066,N_10298);
nand U13739 (N_13739,N_10382,N_10776);
nor U13740 (N_13740,N_10407,N_11198);
or U13741 (N_13741,N_11269,N_11352);
or U13742 (N_13742,N_11962,N_10640);
nor U13743 (N_13743,N_10990,N_10954);
or U13744 (N_13744,N_11444,N_11204);
nand U13745 (N_13745,N_11863,N_11963);
and U13746 (N_13746,N_10821,N_10065);
and U13747 (N_13747,N_11023,N_11477);
nand U13748 (N_13748,N_11045,N_10143);
and U13749 (N_13749,N_10247,N_11054);
nor U13750 (N_13750,N_11623,N_10974);
nor U13751 (N_13751,N_10300,N_11828);
and U13752 (N_13752,N_11068,N_11228);
nor U13753 (N_13753,N_11920,N_11218);
and U13754 (N_13754,N_11239,N_11889);
nor U13755 (N_13755,N_10443,N_10398);
xnor U13756 (N_13756,N_10242,N_11501);
nor U13757 (N_13757,N_10329,N_11382);
and U13758 (N_13758,N_11022,N_10479);
nor U13759 (N_13759,N_11507,N_11683);
nor U13760 (N_13760,N_11162,N_10352);
or U13761 (N_13761,N_11077,N_11986);
nor U13762 (N_13762,N_10762,N_10103);
nor U13763 (N_13763,N_11853,N_11754);
and U13764 (N_13764,N_11189,N_11928);
nand U13765 (N_13765,N_11610,N_10745);
xor U13766 (N_13766,N_11731,N_11559);
and U13767 (N_13767,N_11180,N_11225);
xor U13768 (N_13768,N_10927,N_11761);
xor U13769 (N_13769,N_11235,N_10544);
xnor U13770 (N_13770,N_10637,N_10447);
nor U13771 (N_13771,N_10864,N_10789);
nand U13772 (N_13772,N_10786,N_11918);
nor U13773 (N_13773,N_11919,N_11224);
nand U13774 (N_13774,N_10366,N_11785);
and U13775 (N_13775,N_10704,N_11842);
or U13776 (N_13776,N_10384,N_11543);
nor U13777 (N_13777,N_11376,N_11949);
nand U13778 (N_13778,N_10924,N_11289);
xor U13779 (N_13779,N_11117,N_10951);
and U13780 (N_13780,N_10193,N_10914);
xor U13781 (N_13781,N_10941,N_11630);
xnor U13782 (N_13782,N_10387,N_10669);
nor U13783 (N_13783,N_11743,N_10838);
nor U13784 (N_13784,N_10097,N_10704);
xor U13785 (N_13785,N_11072,N_11195);
nor U13786 (N_13786,N_11464,N_10966);
nand U13787 (N_13787,N_11637,N_10667);
and U13788 (N_13788,N_10239,N_11582);
xnor U13789 (N_13789,N_11323,N_11924);
nand U13790 (N_13790,N_11012,N_11584);
or U13791 (N_13791,N_11764,N_10525);
and U13792 (N_13792,N_11003,N_11934);
and U13793 (N_13793,N_11638,N_11899);
nor U13794 (N_13794,N_11713,N_10241);
nor U13795 (N_13795,N_10435,N_10064);
nand U13796 (N_13796,N_11093,N_10820);
xor U13797 (N_13797,N_11385,N_11456);
xor U13798 (N_13798,N_10754,N_10509);
and U13799 (N_13799,N_11859,N_11236);
nand U13800 (N_13800,N_11721,N_10682);
nor U13801 (N_13801,N_11860,N_10603);
xnor U13802 (N_13802,N_10225,N_11227);
xor U13803 (N_13803,N_11736,N_10273);
and U13804 (N_13804,N_10800,N_10278);
nor U13805 (N_13805,N_10714,N_10756);
nor U13806 (N_13806,N_10659,N_11624);
and U13807 (N_13807,N_11476,N_11711);
and U13808 (N_13808,N_10295,N_11829);
xor U13809 (N_13809,N_11549,N_11125);
nor U13810 (N_13810,N_11005,N_11741);
or U13811 (N_13811,N_10018,N_10009);
nand U13812 (N_13812,N_10147,N_10579);
or U13813 (N_13813,N_11622,N_11869);
nor U13814 (N_13814,N_11293,N_11530);
xor U13815 (N_13815,N_10014,N_11839);
nor U13816 (N_13816,N_10459,N_11494);
nand U13817 (N_13817,N_10393,N_11791);
nand U13818 (N_13818,N_11485,N_11893);
nand U13819 (N_13819,N_11417,N_11641);
xor U13820 (N_13820,N_11800,N_10661);
or U13821 (N_13821,N_11255,N_11646);
or U13822 (N_13822,N_11099,N_10486);
or U13823 (N_13823,N_10123,N_10989);
nor U13824 (N_13824,N_11124,N_11774);
nor U13825 (N_13825,N_10220,N_11254);
nor U13826 (N_13826,N_10002,N_11273);
xnor U13827 (N_13827,N_11766,N_11995);
and U13828 (N_13828,N_11832,N_11823);
nand U13829 (N_13829,N_11958,N_11744);
or U13830 (N_13830,N_11337,N_11789);
or U13831 (N_13831,N_11861,N_10003);
nor U13832 (N_13832,N_10654,N_11224);
xnor U13833 (N_13833,N_10526,N_10217);
and U13834 (N_13834,N_11131,N_11733);
xnor U13835 (N_13835,N_10135,N_10878);
xor U13836 (N_13836,N_10405,N_11002);
nand U13837 (N_13837,N_10485,N_10052);
nor U13838 (N_13838,N_11517,N_11002);
nor U13839 (N_13839,N_10164,N_10840);
xnor U13840 (N_13840,N_10800,N_10656);
xnor U13841 (N_13841,N_10687,N_11895);
nor U13842 (N_13842,N_11063,N_11309);
xor U13843 (N_13843,N_10535,N_11950);
nor U13844 (N_13844,N_10470,N_10908);
or U13845 (N_13845,N_10060,N_10042);
or U13846 (N_13846,N_11433,N_11037);
or U13847 (N_13847,N_11002,N_11170);
and U13848 (N_13848,N_10022,N_10253);
nand U13849 (N_13849,N_10974,N_10300);
xnor U13850 (N_13850,N_11604,N_10764);
nand U13851 (N_13851,N_10189,N_11253);
nand U13852 (N_13852,N_11125,N_10837);
or U13853 (N_13853,N_10231,N_10659);
nand U13854 (N_13854,N_11682,N_11616);
nor U13855 (N_13855,N_10519,N_11290);
or U13856 (N_13856,N_10253,N_10725);
xnor U13857 (N_13857,N_10424,N_11267);
xnor U13858 (N_13858,N_11437,N_11801);
xnor U13859 (N_13859,N_11153,N_10141);
xnor U13860 (N_13860,N_10776,N_11861);
and U13861 (N_13861,N_11843,N_10835);
nand U13862 (N_13862,N_11991,N_10125);
nand U13863 (N_13863,N_11739,N_11665);
xnor U13864 (N_13864,N_10337,N_10016);
and U13865 (N_13865,N_10457,N_10015);
xnor U13866 (N_13866,N_11730,N_10101);
nor U13867 (N_13867,N_10479,N_10600);
xnor U13868 (N_13868,N_11578,N_10539);
nand U13869 (N_13869,N_11081,N_10238);
and U13870 (N_13870,N_10090,N_11979);
nand U13871 (N_13871,N_11637,N_10393);
xnor U13872 (N_13872,N_10117,N_11670);
xor U13873 (N_13873,N_11541,N_10333);
xor U13874 (N_13874,N_10420,N_11965);
and U13875 (N_13875,N_11958,N_10087);
xnor U13876 (N_13876,N_11013,N_10403);
or U13877 (N_13877,N_11298,N_11013);
xnor U13878 (N_13878,N_11700,N_10814);
or U13879 (N_13879,N_11030,N_10579);
or U13880 (N_13880,N_11333,N_11321);
xnor U13881 (N_13881,N_10555,N_11454);
nor U13882 (N_13882,N_11255,N_11949);
or U13883 (N_13883,N_11885,N_10444);
and U13884 (N_13884,N_10786,N_11550);
nor U13885 (N_13885,N_11877,N_11609);
xnor U13886 (N_13886,N_10596,N_10589);
nand U13887 (N_13887,N_10909,N_10129);
nand U13888 (N_13888,N_10894,N_11545);
or U13889 (N_13889,N_11694,N_10878);
or U13890 (N_13890,N_11761,N_10271);
nand U13891 (N_13891,N_11230,N_11484);
or U13892 (N_13892,N_11027,N_10394);
or U13893 (N_13893,N_10772,N_10446);
and U13894 (N_13894,N_10348,N_11223);
xor U13895 (N_13895,N_10863,N_11520);
or U13896 (N_13896,N_10953,N_10667);
or U13897 (N_13897,N_11809,N_11466);
and U13898 (N_13898,N_10954,N_11794);
nand U13899 (N_13899,N_10606,N_11872);
xor U13900 (N_13900,N_10838,N_10846);
and U13901 (N_13901,N_10556,N_11058);
nand U13902 (N_13902,N_10238,N_10992);
and U13903 (N_13903,N_11865,N_11495);
nor U13904 (N_13904,N_10647,N_11715);
nand U13905 (N_13905,N_11079,N_10891);
nand U13906 (N_13906,N_10978,N_10269);
nand U13907 (N_13907,N_11314,N_11629);
or U13908 (N_13908,N_11232,N_10093);
xor U13909 (N_13909,N_10619,N_10560);
and U13910 (N_13910,N_10425,N_10619);
and U13911 (N_13911,N_11919,N_10904);
xor U13912 (N_13912,N_10040,N_11456);
or U13913 (N_13913,N_10712,N_10343);
or U13914 (N_13914,N_10629,N_10883);
or U13915 (N_13915,N_10470,N_10900);
xor U13916 (N_13916,N_10433,N_10237);
and U13917 (N_13917,N_11845,N_11469);
or U13918 (N_13918,N_10192,N_10244);
and U13919 (N_13919,N_10466,N_11235);
or U13920 (N_13920,N_10185,N_11881);
nand U13921 (N_13921,N_10369,N_10273);
or U13922 (N_13922,N_10210,N_11509);
nand U13923 (N_13923,N_10485,N_11546);
nor U13924 (N_13924,N_11403,N_11221);
and U13925 (N_13925,N_11118,N_11687);
or U13926 (N_13926,N_11503,N_10317);
nand U13927 (N_13927,N_10405,N_11162);
nand U13928 (N_13928,N_10642,N_11085);
nor U13929 (N_13929,N_10916,N_11995);
nor U13930 (N_13930,N_11003,N_10528);
nor U13931 (N_13931,N_11785,N_10476);
and U13932 (N_13932,N_10115,N_10986);
nand U13933 (N_13933,N_10053,N_10792);
and U13934 (N_13934,N_11142,N_11657);
nand U13935 (N_13935,N_11820,N_10440);
or U13936 (N_13936,N_11714,N_10355);
and U13937 (N_13937,N_10982,N_10882);
nand U13938 (N_13938,N_11186,N_10294);
or U13939 (N_13939,N_10900,N_11605);
nand U13940 (N_13940,N_11429,N_11430);
nand U13941 (N_13941,N_10210,N_11091);
or U13942 (N_13942,N_11482,N_11349);
or U13943 (N_13943,N_10227,N_10981);
and U13944 (N_13944,N_11806,N_11281);
nor U13945 (N_13945,N_10085,N_10398);
nor U13946 (N_13946,N_10465,N_10493);
xor U13947 (N_13947,N_11986,N_10957);
nor U13948 (N_13948,N_11402,N_10462);
and U13949 (N_13949,N_11212,N_10233);
or U13950 (N_13950,N_10890,N_10574);
xnor U13951 (N_13951,N_10997,N_11478);
or U13952 (N_13952,N_11175,N_11174);
xnor U13953 (N_13953,N_11294,N_11687);
or U13954 (N_13954,N_10997,N_10777);
xnor U13955 (N_13955,N_10210,N_11063);
xor U13956 (N_13956,N_11753,N_10555);
nand U13957 (N_13957,N_11612,N_10977);
and U13958 (N_13958,N_11097,N_11144);
xor U13959 (N_13959,N_11594,N_11278);
nand U13960 (N_13960,N_11041,N_11736);
nor U13961 (N_13961,N_11609,N_10015);
nand U13962 (N_13962,N_10741,N_11014);
or U13963 (N_13963,N_11767,N_11525);
and U13964 (N_13964,N_10182,N_11691);
and U13965 (N_13965,N_10838,N_10354);
nor U13966 (N_13966,N_10753,N_10149);
xnor U13967 (N_13967,N_10019,N_11884);
nand U13968 (N_13968,N_10898,N_10623);
nand U13969 (N_13969,N_10962,N_11324);
and U13970 (N_13970,N_11096,N_10947);
and U13971 (N_13971,N_10930,N_11265);
or U13972 (N_13972,N_10644,N_11067);
and U13973 (N_13973,N_11009,N_10882);
xnor U13974 (N_13974,N_10567,N_11956);
or U13975 (N_13975,N_11818,N_11111);
nand U13976 (N_13976,N_11307,N_11085);
nand U13977 (N_13977,N_10214,N_11671);
or U13978 (N_13978,N_10965,N_10527);
or U13979 (N_13979,N_11432,N_11405);
nand U13980 (N_13980,N_10291,N_11898);
nand U13981 (N_13981,N_11364,N_10674);
and U13982 (N_13982,N_11180,N_11769);
or U13983 (N_13983,N_11674,N_10612);
or U13984 (N_13984,N_10878,N_11654);
nand U13985 (N_13985,N_11827,N_10249);
nand U13986 (N_13986,N_10495,N_10801);
nor U13987 (N_13987,N_10782,N_10650);
and U13988 (N_13988,N_11481,N_10614);
and U13989 (N_13989,N_11330,N_10760);
nand U13990 (N_13990,N_10369,N_11394);
nor U13991 (N_13991,N_10738,N_11576);
xnor U13992 (N_13992,N_11416,N_11004);
or U13993 (N_13993,N_10101,N_10330);
and U13994 (N_13994,N_11666,N_11282);
nor U13995 (N_13995,N_11367,N_10181);
nor U13996 (N_13996,N_10741,N_10956);
nor U13997 (N_13997,N_10070,N_10349);
or U13998 (N_13998,N_10776,N_10634);
or U13999 (N_13999,N_11096,N_11112);
nor U14000 (N_14000,N_12467,N_12227);
nor U14001 (N_14001,N_13772,N_13611);
nand U14002 (N_14002,N_13850,N_13006);
nand U14003 (N_14003,N_13536,N_13515);
nor U14004 (N_14004,N_12368,N_13618);
xnor U14005 (N_14005,N_13632,N_12226);
nor U14006 (N_14006,N_12303,N_13789);
nand U14007 (N_14007,N_12459,N_13034);
nor U14008 (N_14008,N_13253,N_12049);
nor U14009 (N_14009,N_13828,N_12559);
or U14010 (N_14010,N_12911,N_13941);
and U14011 (N_14011,N_12040,N_13599);
and U14012 (N_14012,N_13638,N_12074);
and U14013 (N_14013,N_12811,N_13017);
nor U14014 (N_14014,N_12645,N_13930);
or U14015 (N_14015,N_12357,N_13794);
nand U14016 (N_14016,N_12988,N_13606);
or U14017 (N_14017,N_12504,N_12153);
nand U14018 (N_14018,N_12061,N_13561);
nor U14019 (N_14019,N_12594,N_13112);
xor U14020 (N_14020,N_13128,N_12314);
xor U14021 (N_14021,N_12713,N_12742);
nor U14022 (N_14022,N_12428,N_12627);
nor U14023 (N_14023,N_12012,N_13778);
nand U14024 (N_14024,N_13082,N_13304);
nor U14025 (N_14025,N_12066,N_13982);
xnor U14026 (N_14026,N_13922,N_12806);
nor U14027 (N_14027,N_12095,N_12420);
nor U14028 (N_14028,N_12771,N_13373);
nand U14029 (N_14029,N_12112,N_12773);
xnor U14030 (N_14030,N_12525,N_12278);
xor U14031 (N_14031,N_12511,N_13090);
xor U14032 (N_14032,N_13270,N_13799);
nand U14033 (N_14033,N_12633,N_13550);
nor U14034 (N_14034,N_13177,N_13863);
nor U14035 (N_14035,N_13755,N_13061);
nor U14036 (N_14036,N_12608,N_12327);
and U14037 (N_14037,N_12087,N_13258);
nand U14038 (N_14038,N_13595,N_12922);
nor U14039 (N_14039,N_12872,N_12025);
nand U14040 (N_14040,N_12334,N_12978);
or U14041 (N_14041,N_13833,N_13159);
nor U14042 (N_14042,N_12104,N_13329);
and U14043 (N_14043,N_13967,N_13519);
and U14044 (N_14044,N_13609,N_13903);
or U14045 (N_14045,N_12008,N_12807);
and U14046 (N_14046,N_12435,N_13878);
and U14047 (N_14047,N_13736,N_12022);
nand U14048 (N_14048,N_13150,N_13808);
nor U14049 (N_14049,N_12571,N_12223);
xnor U14050 (N_14050,N_13729,N_12609);
or U14051 (N_14051,N_13059,N_12558);
and U14052 (N_14052,N_13044,N_12330);
or U14053 (N_14053,N_12832,N_13847);
nor U14054 (N_14054,N_13840,N_13917);
nand U14055 (N_14055,N_12199,N_12000);
and U14056 (N_14056,N_12100,N_13195);
nand U14057 (N_14057,N_12668,N_13613);
or U14058 (N_14058,N_12004,N_12803);
xor U14059 (N_14059,N_12660,N_13420);
nor U14060 (N_14060,N_12933,N_12494);
nor U14061 (N_14061,N_13610,N_13173);
and U14062 (N_14062,N_12818,N_13877);
nand U14063 (N_14063,N_13607,N_12257);
nor U14064 (N_14064,N_13769,N_13131);
or U14065 (N_14065,N_12768,N_13512);
or U14066 (N_14066,N_13347,N_12109);
xor U14067 (N_14067,N_13156,N_12723);
nor U14068 (N_14068,N_13644,N_12089);
or U14069 (N_14069,N_13255,N_12146);
nor U14070 (N_14070,N_13980,N_12540);
nand U14071 (N_14071,N_13003,N_13055);
nor U14072 (N_14072,N_13331,N_13357);
nand U14073 (N_14073,N_13886,N_12837);
nand U14074 (N_14074,N_12852,N_12834);
nand U14075 (N_14075,N_12062,N_13225);
nand U14076 (N_14076,N_13733,N_12699);
and U14077 (N_14077,N_12746,N_13297);
nor U14078 (N_14078,N_12648,N_13210);
and U14079 (N_14079,N_13603,N_12775);
nor U14080 (N_14080,N_12506,N_12204);
or U14081 (N_14081,N_12508,N_13093);
xnor U14082 (N_14082,N_12077,N_13950);
or U14083 (N_14083,N_12247,N_12736);
and U14084 (N_14084,N_12866,N_13094);
nand U14085 (N_14085,N_12085,N_12339);
nand U14086 (N_14086,N_13287,N_12372);
xnor U14087 (N_14087,N_12934,N_12889);
nand U14088 (N_14088,N_12588,N_12870);
nor U14089 (N_14089,N_13722,N_13309);
xnor U14090 (N_14090,N_12980,N_13237);
nor U14091 (N_14091,N_13263,N_13896);
nor U14092 (N_14092,N_13020,N_13608);
nand U14093 (N_14093,N_13499,N_12280);
and U14094 (N_14094,N_13779,N_13320);
nand U14095 (N_14095,N_12300,N_13506);
nor U14096 (N_14096,N_13694,N_12618);
xor U14097 (N_14097,N_13548,N_13174);
and U14098 (N_14098,N_12892,N_13516);
nor U14099 (N_14099,N_12086,N_13882);
and U14100 (N_14100,N_12875,N_12097);
nor U14101 (N_14101,N_12485,N_12195);
nand U14102 (N_14102,N_13276,N_13222);
nand U14103 (N_14103,N_12333,N_12356);
and U14104 (N_14104,N_12105,N_13569);
and U14105 (N_14105,N_13932,N_12361);
nand U14106 (N_14106,N_12441,N_13440);
nor U14107 (N_14107,N_12293,N_12054);
and U14108 (N_14108,N_13683,N_13666);
xor U14109 (N_14109,N_12938,N_12786);
and U14110 (N_14110,N_13415,N_12555);
or U14111 (N_14111,N_13453,N_12294);
xnor U14112 (N_14112,N_12737,N_12058);
and U14113 (N_14113,N_13949,N_12917);
or U14114 (N_14114,N_13365,N_12297);
or U14115 (N_14115,N_13360,N_12232);
or U14116 (N_14116,N_12250,N_12408);
nor U14117 (N_14117,N_12170,N_13624);
nor U14118 (N_14118,N_13084,N_13057);
and U14119 (N_14119,N_12589,N_13025);
nand U14120 (N_14120,N_12733,N_13243);
and U14121 (N_14121,N_12113,N_13634);
nand U14122 (N_14122,N_13235,N_13612);
or U14123 (N_14123,N_13731,N_13835);
or U14124 (N_14124,N_13909,N_13122);
and U14125 (N_14125,N_12143,N_13132);
nor U14126 (N_14126,N_13598,N_12501);
nor U14127 (N_14127,N_12614,N_12041);
xnor U14128 (N_14128,N_13919,N_13018);
nor U14129 (N_14129,N_12568,N_13629);
nand U14130 (N_14130,N_12584,N_13597);
nand U14131 (N_14131,N_12789,N_12517);
xor U14132 (N_14132,N_13213,N_12045);
nand U14133 (N_14133,N_13208,N_12631);
nor U14134 (N_14134,N_13169,N_13724);
nand U14135 (N_14135,N_13230,N_13231);
or U14136 (N_14136,N_13585,N_12521);
nor U14137 (N_14137,N_12815,N_13868);
xnor U14138 (N_14138,N_13591,N_13524);
nor U14139 (N_14139,N_13446,N_13911);
nor U14140 (N_14140,N_12343,N_13185);
xor U14141 (N_14141,N_12284,N_12901);
nor U14142 (N_14142,N_13383,N_12847);
and U14143 (N_14143,N_12065,N_12299);
and U14144 (N_14144,N_13551,N_13771);
nand U14145 (N_14145,N_12546,N_12003);
or U14146 (N_14146,N_13823,N_12320);
nor U14147 (N_14147,N_12399,N_13509);
nand U14148 (N_14148,N_12890,N_12242);
nor U14149 (N_14149,N_13553,N_12384);
and U14150 (N_14150,N_12636,N_13510);
or U14151 (N_14151,N_12474,N_12784);
nor U14152 (N_14152,N_12562,N_13926);
xor U14153 (N_14153,N_13182,N_12903);
xnor U14154 (N_14154,N_12676,N_13458);
nor U14155 (N_14155,N_13668,N_12311);
xnor U14156 (N_14156,N_13764,N_12125);
xnor U14157 (N_14157,N_12793,N_12183);
nor U14158 (N_14158,N_12478,N_13121);
nand U14159 (N_14159,N_12887,N_13408);
or U14160 (N_14160,N_13049,N_13385);
and U14161 (N_14161,N_13582,N_12079);
nand U14162 (N_14162,N_13368,N_13032);
nor U14163 (N_14163,N_12677,N_12430);
xnor U14164 (N_14164,N_13405,N_12068);
and U14165 (N_14165,N_12581,N_12740);
and U14166 (N_14166,N_12071,N_12440);
nand U14167 (N_14167,N_13052,N_12702);
xor U14168 (N_14168,N_12745,N_12629);
nor U14169 (N_14169,N_13616,N_12635);
xor U14170 (N_14170,N_12126,N_12804);
xnor U14171 (N_14171,N_12265,N_12172);
nand U14172 (N_14172,N_13189,N_13783);
nand U14173 (N_14173,N_13791,N_13924);
nor U14174 (N_14174,N_13389,N_13708);
nand U14175 (N_14175,N_12014,N_12873);
nand U14176 (N_14176,N_13285,N_13647);
nor U14177 (N_14177,N_12292,N_13776);
or U14178 (N_14178,N_12347,N_12448);
or U14179 (N_14179,N_12395,N_13352);
nor U14180 (N_14180,N_12624,N_13832);
nor U14181 (N_14181,N_13223,N_13552);
nand U14182 (N_14182,N_12744,N_12874);
nand U14183 (N_14183,N_13797,N_13397);
nor U14184 (N_14184,N_12490,N_12850);
nor U14185 (N_14185,N_12638,N_12124);
or U14186 (N_14186,N_13404,N_12835);
nand U14187 (N_14187,N_13460,N_13978);
xnor U14188 (N_14188,N_12350,N_12221);
nor U14189 (N_14189,N_12241,N_13447);
nor U14190 (N_14190,N_12527,N_13406);
xor U14191 (N_14191,N_12405,N_12725);
or U14192 (N_14192,N_12586,N_13554);
and U14193 (N_14193,N_12020,N_12164);
nand U14194 (N_14194,N_12050,N_13815);
nor U14195 (N_14195,N_12628,N_13426);
nand U14196 (N_14196,N_13388,N_12947);
xnor U14197 (N_14197,N_12205,N_13951);
nand U14198 (N_14198,N_13105,N_12279);
nor U14199 (N_14199,N_13859,N_13016);
nor U14200 (N_14200,N_13702,N_13410);
nor U14201 (N_14201,N_13417,N_12497);
nor U14202 (N_14202,N_13330,N_12643);
and U14203 (N_14203,N_13313,N_13448);
nand U14204 (N_14204,N_12415,N_12968);
nor U14205 (N_14205,N_13812,N_13190);
or U14206 (N_14206,N_12048,N_12094);
nor U14207 (N_14207,N_12817,N_13322);
xnor U14208 (N_14208,N_13178,N_13146);
nor U14209 (N_14209,N_12138,N_12021);
nand U14210 (N_14210,N_12748,N_12215);
and U14211 (N_14211,N_13572,N_13386);
nor U14212 (N_14212,N_12912,N_12083);
nand U14213 (N_14213,N_13861,N_13176);
nand U14214 (N_14214,N_12503,N_13699);
and U14215 (N_14215,N_13531,N_12871);
nor U14216 (N_14216,N_13450,N_13673);
and U14217 (N_14217,N_13050,N_13845);
and U14218 (N_14218,N_13517,N_12433);
xor U14219 (N_14219,N_13490,N_13558);
xor U14220 (N_14220,N_12619,N_12523);
and U14221 (N_14221,N_12990,N_13805);
nand U14222 (N_14222,N_13328,N_12304);
or U14223 (N_14223,N_12749,N_13803);
nor U14224 (N_14224,N_13894,N_13849);
and U14225 (N_14225,N_12839,N_13854);
nand U14226 (N_14226,N_13179,N_13818);
and U14227 (N_14227,N_13549,N_12262);
nand U14228 (N_14228,N_13977,N_13296);
nor U14229 (N_14229,N_13513,N_13525);
and U14230 (N_14230,N_12877,N_12507);
nor U14231 (N_14231,N_12722,N_13391);
nor U14232 (N_14232,N_13379,N_12222);
nand U14233 (N_14233,N_12683,N_13481);
and U14234 (N_14234,N_13312,N_13398);
nor U14235 (N_14235,N_13002,N_13393);
or U14236 (N_14236,N_13482,N_13895);
xor U14237 (N_14237,N_12403,N_13814);
nand U14238 (N_14238,N_13622,N_13944);
nand U14239 (N_14239,N_12731,N_12704);
nor U14240 (N_14240,N_13143,N_12667);
xor U14241 (N_14241,N_12084,N_13212);
nand U14242 (N_14242,N_13975,N_13884);
or U14243 (N_14243,N_13893,N_12264);
nor U14244 (N_14244,N_12259,N_12753);
xor U14245 (N_14245,N_12998,N_12228);
nand U14246 (N_14246,N_12759,N_13291);
xnor U14247 (N_14247,N_13826,N_12092);
nor U14248 (N_14248,N_12565,N_13505);
nand U14249 (N_14249,N_12034,N_12069);
nor U14250 (N_14250,N_13495,N_12601);
nand U14251 (N_14251,N_13438,N_13269);
nand U14252 (N_14252,N_12857,N_13630);
xnor U14253 (N_14253,N_13675,N_12370);
nand U14254 (N_14254,N_12761,N_13154);
or U14255 (N_14255,N_12772,N_12392);
nand U14256 (N_14256,N_13913,N_13841);
or U14257 (N_14257,N_13838,N_13377);
or U14258 (N_14258,N_13204,N_13245);
nand U14259 (N_14259,N_13374,N_13651);
nand U14260 (N_14260,N_13257,N_12574);
or U14261 (N_14261,N_12822,N_12686);
nor U14262 (N_14262,N_12287,N_12267);
xor U14263 (N_14263,N_12920,N_12452);
or U14264 (N_14264,N_13614,N_13087);
nor U14265 (N_14265,N_13445,N_13750);
nand U14266 (N_14266,N_12055,N_12487);
nor U14267 (N_14267,N_12017,N_13316);
xor U14268 (N_14268,N_13546,N_12332);
and U14269 (N_14269,N_12838,N_12767);
or U14270 (N_14270,N_12578,N_12449);
and U14271 (N_14271,N_12701,N_13014);
or U14272 (N_14272,N_12269,N_13567);
xnor U14273 (N_14273,N_12785,N_13075);
or U14274 (N_14274,N_13311,N_12039);
nand U14275 (N_14275,N_13160,N_12121);
and U14276 (N_14276,N_12496,N_13457);
and U14277 (N_14277,N_13538,N_13083);
nor U14278 (N_14278,N_12982,N_12187);
nand U14279 (N_14279,N_12769,N_13541);
or U14280 (N_14280,N_13762,N_13422);
nand U14281 (N_14281,N_12401,N_13141);
nand U14282 (N_14282,N_12621,N_13749);
and U14283 (N_14283,N_12853,N_13959);
xor U14284 (N_14284,N_12218,N_12475);
xor U14285 (N_14285,N_13931,N_13916);
nand U14286 (N_14286,N_13820,N_12463);
nand U14287 (N_14287,N_12833,N_13110);
nor U14288 (N_14288,N_12549,N_12979);
nor U14289 (N_14289,N_12970,N_13645);
nor U14290 (N_14290,N_12792,N_12605);
nand U14291 (N_14291,N_13649,N_13314);
xnor U14292 (N_14292,N_13487,N_12579);
or U14293 (N_14293,N_12424,N_13214);
nor U14294 (N_14294,N_12886,N_13573);
xor U14295 (N_14295,N_13232,N_13753);
and U14296 (N_14296,N_12386,N_12466);
or U14297 (N_14297,N_13793,N_13958);
xor U14298 (N_14298,N_12144,N_13081);
and U14299 (N_14299,N_13431,N_13413);
nor U14300 (N_14300,N_12567,N_13592);
or U14301 (N_14301,N_13837,N_12539);
and U14302 (N_14302,N_13888,N_13107);
or U14303 (N_14303,N_13286,N_13674);
nor U14304 (N_14304,N_13349,N_13777);
nand U14305 (N_14305,N_13175,N_12597);
xnor U14306 (N_14306,N_12596,N_13339);
nor U14307 (N_14307,N_13273,N_13461);
or U14308 (N_14308,N_12116,N_12305);
nand U14309 (N_14309,N_12093,N_13817);
or U14310 (N_14310,N_13705,N_13477);
or U14311 (N_14311,N_12908,N_12708);
or U14312 (N_14312,N_13716,N_13593);
nor U14313 (N_14313,N_12445,N_12700);
xor U14314 (N_14314,N_12896,N_13117);
or U14315 (N_14315,N_13165,N_13875);
and U14316 (N_14316,N_12393,N_13635);
and U14317 (N_14317,N_13892,N_12741);
or U14318 (N_14318,N_13576,N_13211);
and U14319 (N_14319,N_12688,N_13976);
nor U14320 (N_14320,N_12669,N_13631);
and U14321 (N_14321,N_13046,N_13429);
nor U14322 (N_14322,N_13047,N_13704);
nor U14323 (N_14323,N_13707,N_13155);
xor U14324 (N_14324,N_12245,N_12253);
or U14325 (N_14325,N_12375,N_12770);
nor U14326 (N_14326,N_13943,N_13464);
or U14327 (N_14327,N_12394,N_13292);
and U14328 (N_14328,N_12431,N_12483);
xor U14329 (N_14329,N_13129,N_12937);
xnor U14330 (N_14330,N_13130,N_13470);
nor U14331 (N_14331,N_12024,N_12047);
nand U14332 (N_14332,N_13305,N_12033);
and U14333 (N_14333,N_13378,N_12727);
xnor U14334 (N_14334,N_13372,N_12916);
and U14335 (N_14335,N_13358,N_13168);
nor U14336 (N_14336,N_12028,N_13170);
nor U14337 (N_14337,N_13994,N_13993);
or U14338 (N_14338,N_12159,N_13955);
nor U14339 (N_14339,N_12096,N_13452);
or U14340 (N_14340,N_13663,N_12224);
and U14341 (N_14341,N_12977,N_12321);
and U14342 (N_14342,N_13307,N_13727);
nand U14343 (N_14343,N_13682,N_13118);
and U14344 (N_14344,N_12653,N_13617);
nand U14345 (N_14345,N_13089,N_12328);
nor U14346 (N_14346,N_13157,N_13241);
nor U14347 (N_14347,N_12417,N_13885);
and U14348 (N_14348,N_13187,N_13010);
xnor U14349 (N_14349,N_13425,N_13233);
or U14350 (N_14350,N_13074,N_12208);
nor U14351 (N_14351,N_13180,N_13206);
or U14352 (N_14352,N_12036,N_12705);
nand U14353 (N_14353,N_12575,N_12714);
xnor U14354 (N_14354,N_12359,N_13637);
nor U14355 (N_14355,N_12031,N_12695);
nand U14356 (N_14356,N_13684,N_13923);
xor U14357 (N_14357,N_13427,N_13038);
and U14358 (N_14358,N_12529,N_13945);
nand U14359 (N_14359,N_13865,N_13321);
nor U14360 (N_14360,N_13434,N_12082);
or U14361 (N_14361,N_12698,N_13031);
nand U14362 (N_14362,N_12925,N_13954);
xor U14363 (N_14363,N_13876,N_13532);
or U14364 (N_14364,N_12165,N_12824);
and U14365 (N_14365,N_13503,N_12362);
or U14366 (N_14366,N_13758,N_12882);
nand U14367 (N_14367,N_12078,N_13441);
xor U14368 (N_14368,N_12591,N_12111);
nand U14369 (N_14369,N_12880,N_12632);
nand U14370 (N_14370,N_13897,N_13765);
nor U14371 (N_14371,N_13138,N_12548);
nor U14372 (N_14372,N_12717,N_13571);
and U14373 (N_14373,N_13676,N_12531);
and U14374 (N_14374,N_13900,N_13376);
xor U14375 (N_14375,N_12661,N_12651);
or U14376 (N_14376,N_13315,N_12456);
or U14377 (N_14377,N_12639,N_12842);
xor U14378 (N_14378,N_12751,N_12056);
nand U14379 (N_14379,N_12155,N_12171);
xor U14380 (N_14380,N_12367,N_13407);
xnor U14381 (N_14381,N_13578,N_13891);
nand U14382 (N_14382,N_13703,N_13934);
or U14383 (N_14383,N_13889,N_12486);
nor U14384 (N_14384,N_13801,N_12390);
and U14385 (N_14385,N_13166,N_13589);
nand U14386 (N_14386,N_12997,N_13744);
nand U14387 (N_14387,N_12801,N_12220);
nand U14388 (N_14388,N_12928,N_12239);
nor U14389 (N_14389,N_12290,N_12743);
nor U14390 (N_14390,N_13290,N_13338);
nor U14391 (N_14391,N_12642,N_13730);
and U14392 (N_14392,N_13077,N_12551);
nor U14393 (N_14393,N_13471,N_12935);
and U14394 (N_14394,N_13601,N_13437);
xnor U14395 (N_14395,N_13565,N_12726);
and U14396 (N_14396,N_12943,N_12285);
xnor U14397 (N_14397,N_13192,N_13918);
and U14398 (N_14398,N_12157,N_13557);
xnor U14399 (N_14399,N_13323,N_13660);
nand U14400 (N_14400,N_13158,N_13822);
nor U14401 (N_14401,N_12971,N_12681);
and U14402 (N_14402,N_13834,N_12373);
and U14403 (N_14403,N_12984,N_12240);
nor U14404 (N_14404,N_12388,N_13709);
xor U14405 (N_14405,N_12752,N_12354);
nand U14406 (N_14406,N_13181,N_12592);
xor U14407 (N_14407,N_12337,N_12396);
nand U14408 (N_14408,N_12989,N_13714);
or U14409 (N_14409,N_13665,N_13033);
nand U14410 (N_14410,N_12098,N_13164);
nand U14411 (N_14411,N_12355,N_12493);
and U14412 (N_14412,N_13742,N_12843);
nor U14413 (N_14413,N_12719,N_13428);
nor U14414 (N_14414,N_13927,N_12364);
xnor U14415 (N_14415,N_12295,N_13399);
xor U14416 (N_14416,N_13098,N_13504);
xnor U14417 (N_14417,N_12696,N_12136);
and U14418 (N_14418,N_13964,N_13342);
or U14419 (N_14419,N_13656,N_13806);
and U14420 (N_14420,N_12072,N_12881);
nand U14421 (N_14421,N_13396,N_12132);
and U14422 (N_14422,N_12961,N_12762);
xor U14423 (N_14423,N_13334,N_13853);
nand U14424 (N_14424,N_13879,N_12057);
nand U14425 (N_14425,N_13872,N_12489);
and U14426 (N_14426,N_13186,N_13124);
nand U14427 (N_14427,N_12007,N_13069);
nor U14428 (N_14428,N_12458,N_12940);
nand U14429 (N_14429,N_12996,N_13667);
nand U14430 (N_14430,N_13902,N_13449);
or U14431 (N_14431,N_12663,N_13153);
nand U14432 (N_14432,N_13627,N_13172);
xor U14433 (N_14433,N_12035,N_13343);
nor U14434 (N_14434,N_13364,N_13641);
xor U14435 (N_14435,N_13183,N_12826);
and U14436 (N_14436,N_13721,N_13906);
and U14437 (N_14437,N_12657,N_12999);
nor U14438 (N_14438,N_12500,N_12867);
nor U14439 (N_14439,N_12819,N_13278);
and U14440 (N_14440,N_12595,N_13654);
and U14441 (N_14441,N_12213,N_12409);
xnor U14442 (N_14442,N_12081,N_12813);
or U14443 (N_14443,N_13527,N_12156);
or U14444 (N_14444,N_12992,N_13813);
and U14445 (N_14445,N_12439,N_12387);
nor U14446 (N_14446,N_12831,N_13700);
nand U14447 (N_14447,N_13294,N_12344);
or U14448 (N_14448,N_12029,N_13851);
or U14449 (N_14449,N_13488,N_12108);
and U14450 (N_14450,N_12110,N_13619);
and U14451 (N_14451,N_13662,N_13101);
nand U14452 (N_14452,N_13384,N_12616);
nand U14453 (N_14453,N_12856,N_12502);
xnor U14454 (N_14454,N_13000,N_13479);
nor U14455 (N_14455,N_13325,N_12461);
and U14456 (N_14456,N_12697,N_13957);
xnor U14457 (N_14457,N_12391,N_13860);
and U14458 (N_14458,N_12101,N_13809);
or U14459 (N_14459,N_12322,N_13259);
xnor U14460 (N_14460,N_13562,N_12471);
or U14461 (N_14461,N_13302,N_12271);
nor U14462 (N_14462,N_12052,N_13113);
and U14463 (N_14463,N_13356,N_12583);
and U14464 (N_14464,N_12782,N_13459);
nor U14465 (N_14465,N_13672,N_12821);
or U14466 (N_14466,N_13123,N_13962);
and U14467 (N_14467,N_13247,N_13590);
xnor U14468 (N_14468,N_12134,N_13933);
xnor U14469 (N_14469,N_12230,N_13987);
and U14470 (N_14470,N_12203,N_13827);
nor U14471 (N_14471,N_12902,N_12277);
and U14472 (N_14472,N_13856,N_13560);
or U14473 (N_14473,N_13394,N_13830);
and U14474 (N_14474,N_13579,N_13348);
nor U14475 (N_14475,N_13946,N_13824);
nor U14476 (N_14476,N_13831,N_13870);
nand U14477 (N_14477,N_13528,N_12406);
xnor U14478 (N_14478,N_13811,N_12192);
nor U14479 (N_14479,N_13937,N_13463);
nor U14480 (N_14480,N_13734,N_12965);
nor U14481 (N_14481,N_12664,N_13864);
xnor U14482 (N_14482,N_12122,N_12225);
and U14483 (N_14483,N_12505,N_12480);
and U14484 (N_14484,N_12210,N_12479);
and U14485 (N_14485,N_13474,N_12673);
xnor U14486 (N_14486,N_12691,N_12042);
xnor U14487 (N_14487,N_13855,N_12703);
and U14488 (N_14488,N_12897,N_13989);
or U14489 (N_14489,N_13367,N_12115);
xor U14490 (N_14490,N_12672,N_13690);
and U14491 (N_14491,N_12120,N_13604);
and U14492 (N_14492,N_12185,N_12534);
and U14493 (N_14493,N_13821,N_13792);
nor U14494 (N_14494,N_13686,N_12604);
or U14495 (N_14495,N_13152,N_12810);
nand U14496 (N_14496,N_12532,N_13203);
or U14497 (N_14497,N_13483,N_13220);
or U14498 (N_14498,N_13430,N_12318);
or U14499 (N_14499,N_13713,N_13333);
and U14500 (N_14500,N_13335,N_12900);
nor U14501 (N_14501,N_12561,N_12932);
nand U14502 (N_14502,N_12182,N_13298);
nor U14503 (N_14503,N_12640,N_13785);
xnor U14504 (N_14504,N_13628,N_13738);
nand U14505 (N_14505,N_13843,N_13361);
or U14506 (N_14506,N_12678,N_13277);
xnor U14507 (N_14507,N_12477,N_13256);
and U14508 (N_14508,N_12885,N_13680);
and U14509 (N_14509,N_13380,N_12385);
nand U14510 (N_14510,N_12346,N_13639);
nor U14511 (N_14511,N_12553,N_12335);
xnor U14512 (N_14512,N_13904,N_12926);
or U14513 (N_14513,N_13478,N_12948);
nand U14514 (N_14514,N_13011,N_13184);
xor U14515 (N_14515,N_12805,N_12693);
xnor U14516 (N_14516,N_13621,N_13401);
or U14517 (N_14517,N_13804,N_12070);
and U14518 (N_14518,N_13416,N_12249);
xnor U14519 (N_14519,N_13209,N_12515);
nor U14520 (N_14520,N_12016,N_13246);
and U14521 (N_14521,N_13022,N_13359);
and U14522 (N_14522,N_12312,N_13787);
xnor U14523 (N_14523,N_13088,N_12206);
nand U14524 (N_14524,N_13692,N_13844);
or U14525 (N_14525,N_12718,N_12543);
and U14526 (N_14526,N_13655,N_13414);
xnor U14527 (N_14527,N_13745,N_13048);
nor U14528 (N_14528,N_13111,N_12924);
and U14529 (N_14529,N_12282,N_12296);
and U14530 (N_14530,N_13681,N_12552);
or U14531 (N_14531,N_12956,N_12231);
nor U14532 (N_14532,N_12738,N_12827);
xor U14533 (N_14533,N_13197,N_13371);
nand U14534 (N_14534,N_13332,N_13908);
or U14535 (N_14535,N_13226,N_12283);
and U14536 (N_14536,N_13508,N_13574);
nand U14537 (N_14537,N_13581,N_13915);
or U14538 (N_14538,N_12791,N_12302);
nand U14539 (N_14539,N_12410,N_13036);
and U14540 (N_14540,N_12426,N_13191);
nand U14541 (N_14541,N_13701,N_12235);
nand U14542 (N_14542,N_12603,N_13754);
and U14543 (N_14543,N_13747,N_13486);
nand U14544 (N_14544,N_13171,N_12654);
or U14545 (N_14545,N_12139,N_13969);
and U14546 (N_14546,N_13340,N_13042);
nand U14547 (N_14547,N_12413,N_13988);
and U14548 (N_14548,N_12895,N_13695);
nor U14549 (N_14549,N_13956,N_12706);
nand U14550 (N_14550,N_12455,N_12254);
nor U14551 (N_14551,N_13898,N_13299);
or U14552 (N_14552,N_13147,N_13646);
and U14553 (N_14553,N_12128,N_13545);
or U14554 (N_14554,N_12106,N_13542);
and U14555 (N_14555,N_13491,N_12537);
nand U14556 (N_14556,N_13162,N_13108);
xor U14557 (N_14557,N_12644,N_12141);
nor U14558 (N_14558,N_12038,N_12566);
or U14559 (N_14559,N_13436,N_13858);
xnor U14560 (N_14560,N_12217,N_12888);
or U14561 (N_14561,N_12946,N_12904);
and U14562 (N_14562,N_13984,N_12569);
and U14563 (N_14563,N_13462,N_12338);
nor U14564 (N_14564,N_12258,N_13009);
or U14565 (N_14565,N_12309,N_13697);
or U14566 (N_14566,N_13970,N_12200);
and U14567 (N_14567,N_12600,N_13514);
nand U14568 (N_14568,N_13421,N_13035);
and U14569 (N_14569,N_12602,N_13511);
nand U14570 (N_14570,N_13685,N_13717);
or U14571 (N_14571,N_12091,N_13466);
and U14572 (N_14572,N_12064,N_12286);
and U14573 (N_14573,N_13496,N_12266);
xnor U14574 (N_14574,N_12613,N_12809);
xnor U14575 (N_14575,N_13706,N_13403);
xnor U14576 (N_14576,N_13983,N_13319);
or U14577 (N_14577,N_13045,N_13196);
and U14578 (N_14578,N_12854,N_12363);
nand U14579 (N_14579,N_12959,N_12950);
or U14580 (N_14580,N_12976,N_12914);
xnor U14581 (N_14581,N_13207,N_13099);
or U14582 (N_14582,N_13106,N_12634);
xnor U14583 (N_14583,N_12829,N_12342);
xnor U14584 (N_14584,N_13272,N_13200);
or U14585 (N_14585,N_13788,N_12707);
or U14586 (N_14586,N_12797,N_13874);
or U14587 (N_14587,N_12869,N_12689);
nor U14588 (N_14588,N_13501,N_13746);
or U14589 (N_14589,N_12374,N_12963);
and U14590 (N_14590,N_13523,N_13974);
and U14591 (N_14591,N_12764,N_12812);
nor U14592 (N_14592,N_13234,N_13766);
and U14593 (N_14593,N_13659,N_12724);
nor U14594 (N_14594,N_12353,N_13752);
nor U14595 (N_14595,N_12617,N_12983);
or U14596 (N_14596,N_12099,N_13953);
nand U14597 (N_14597,N_12319,N_12324);
nand U14598 (N_14598,N_13412,N_13972);
xnor U14599 (N_14599,N_13995,N_12734);
nor U14600 (N_14600,N_13715,N_12244);
and U14601 (N_14601,N_13767,N_12536);
xnor U14602 (N_14602,N_13650,N_12891);
nor U14603 (N_14603,N_12180,N_12637);
nand U14604 (N_14604,N_13761,N_13836);
or U14605 (N_14605,N_13940,N_13719);
or U14606 (N_14606,N_12954,N_12044);
xnor U14607 (N_14607,N_12377,N_13202);
nor U14608 (N_14608,N_12468,N_12379);
xor U14609 (N_14609,N_12790,N_12760);
xor U14610 (N_14610,N_12450,N_13219);
and U14611 (N_14611,N_13381,N_12783);
or U14612 (N_14612,N_12991,N_13366);
or U14613 (N_14613,N_12484,N_13288);
nor U14614 (N_14614,N_13116,N_12993);
and U14615 (N_14615,N_12434,N_12747);
xor U14616 (N_14616,N_13043,N_13149);
or U14617 (N_14617,N_13539,N_13345);
xnor U14618 (N_14618,N_13947,N_12646);
or U14619 (N_14619,N_13228,N_12865);
or U14620 (N_14620,N_12414,N_13781);
nand U14621 (N_14621,N_13839,N_12163);
nor U14622 (N_14622,N_13575,N_13188);
and U14623 (N_14623,N_12735,N_12154);
and U14624 (N_14624,N_12929,N_13625);
xor U14625 (N_14625,N_12730,N_12482);
nand U14626 (N_14626,N_12013,N_13104);
and U14627 (N_14627,N_13529,N_12469);
and U14628 (N_14628,N_12272,N_13559);
nand U14629 (N_14629,N_12795,N_13015);
nor U14630 (N_14630,N_13555,N_12006);
or U14631 (N_14631,N_12472,N_13281);
nand U14632 (N_14632,N_12184,N_12102);
nand U14633 (N_14633,N_13530,N_12179);
nand U14634 (N_14634,N_12067,N_13248);
xnor U14635 (N_14635,N_12438,N_12758);
nor U14636 (N_14636,N_13005,N_12899);
nand U14637 (N_14637,N_12957,N_12625);
and U14638 (N_14638,N_12560,N_13040);
xor U14639 (N_14639,N_12127,N_12216);
nand U14640 (N_14640,N_12512,N_13326);
xor U14641 (N_14641,N_13004,N_13938);
and U14642 (N_14642,N_12939,N_13939);
and U14643 (N_14643,N_12690,N_12470);
or U14644 (N_14644,N_13300,N_12298);
and U14645 (N_14645,N_12964,N_12766);
and U14646 (N_14646,N_12550,N_13881);
or U14647 (N_14647,N_13925,N_13802);
nor U14648 (N_14648,N_13521,N_13085);
xor U14649 (N_14649,N_12234,N_12130);
nor U14650 (N_14650,N_12114,N_13748);
or U14651 (N_14651,N_12615,N_12315);
nor U14652 (N_14652,N_12323,N_12142);
nor U14653 (N_14653,N_13687,N_13664);
nor U14654 (N_14654,N_12107,N_12306);
or U14655 (N_14655,N_12263,N_12656);
nand U14656 (N_14656,N_13454,N_13520);
or U14657 (N_14657,N_12329,N_13027);
nand U14658 (N_14658,N_12160,N_13126);
and U14659 (N_14659,N_13914,N_12510);
xor U14660 (N_14660,N_12129,N_12670);
or U14661 (N_14661,N_12577,N_13756);
and U14662 (N_14662,N_12576,N_13873);
and U14663 (N_14663,N_13244,N_13456);
nor U14664 (N_14664,N_12910,N_13021);
nand U14665 (N_14665,N_13301,N_13936);
or U14666 (N_14666,N_13533,N_12945);
or U14667 (N_14667,N_13535,N_12454);
and U14668 (N_14668,N_12599,N_12437);
xnor U14669 (N_14669,N_12196,N_13167);
nor U14670 (N_14670,N_12671,N_13268);
nand U14671 (N_14671,N_12816,N_13540);
nor U14672 (N_14672,N_13807,N_13563);
nor U14673 (N_14673,N_13587,N_12229);
or U14674 (N_14674,N_12799,N_12610);
xor U14675 (N_14675,N_13899,N_13484);
nor U14676 (N_14676,N_13432,N_13921);
nor U14677 (N_14677,N_12080,N_12879);
nand U14678 (N_14678,N_13318,N_13080);
xnor U14679 (N_14679,N_12237,N_12352);
and U14680 (N_14680,N_12756,N_12518);
or U14681 (N_14681,N_12573,N_12612);
nor U14682 (N_14682,N_12491,N_13710);
nor U14683 (N_14683,N_13480,N_12960);
nor U14684 (N_14684,N_12909,N_12582);
or U14685 (N_14685,N_13267,N_12345);
and U14686 (N_14686,N_12191,N_12010);
nand U14687 (N_14687,N_12453,N_12942);
nand U14688 (N_14688,N_13400,N_12710);
nand U14689 (N_14689,N_12754,N_12572);
or U14690 (N_14690,N_13402,N_13007);
xor U14691 (N_14691,N_12623,N_12005);
or U14692 (N_14692,N_12898,N_13566);
nand U14693 (N_14693,N_13056,N_13303);
nor U14694 (N_14694,N_12802,N_13370);
and U14695 (N_14695,N_13240,N_12958);
nor U14696 (N_14696,N_13770,N_12137);
nor U14697 (N_14697,N_12972,N_13133);
xnor U14698 (N_14698,N_12168,N_12019);
xor U14699 (N_14699,N_13584,N_13965);
and U14700 (N_14700,N_13008,N_13774);
nand U14701 (N_14701,N_12611,N_12341);
or U14702 (N_14702,N_12514,N_12348);
and U14703 (N_14703,N_13568,N_12451);
nor U14704 (N_14704,N_12840,N_13489);
nor U14705 (N_14705,N_13757,N_12519);
nor U14706 (N_14706,N_12447,N_12243);
xor U14707 (N_14707,N_13289,N_13825);
or U14708 (N_14708,N_13023,N_12117);
or U14709 (N_14709,N_12161,N_13829);
nor U14710 (N_14710,N_13910,N_12538);
nand U14711 (N_14711,N_13648,N_13229);
nor U14712 (N_14712,N_13051,N_13691);
xor U14713 (N_14713,N_12027,N_12765);
nor U14714 (N_14714,N_12798,N_13282);
or U14715 (N_14715,N_13265,N_13720);
nand U14716 (N_14716,N_12444,N_13079);
or U14717 (N_14717,N_12544,N_13280);
and U14718 (N_14718,N_12481,N_13498);
xor U14719 (N_14719,N_12652,N_12255);
and U14720 (N_14720,N_12140,N_12252);
or U14721 (N_14721,N_12181,N_12397);
or U14722 (N_14722,N_13775,N_13097);
nand U14723 (N_14723,N_13418,N_13693);
or U14724 (N_14724,N_12011,N_13261);
and U14725 (N_14725,N_12135,N_13390);
and U14726 (N_14726,N_12499,N_12694);
and U14727 (N_14727,N_13145,N_13981);
and U14728 (N_14728,N_12953,N_13078);
xnor U14729 (N_14729,N_13966,N_13985);
nor U14730 (N_14730,N_12830,N_12246);
xnor U14731 (N_14731,N_12564,N_13136);
xor U14732 (N_14732,N_13986,N_13115);
and U14733 (N_14733,N_12201,N_13395);
xnor U14734 (N_14734,N_13819,N_13473);
and U14735 (N_14735,N_12404,N_13594);
nor U14736 (N_14736,N_13577,N_13901);
xnor U14737 (N_14737,N_12851,N_12018);
and U14738 (N_14738,N_13869,N_13127);
nand U14739 (N_14739,N_13640,N_13283);
and U14740 (N_14740,N_12655,N_13866);
nand U14741 (N_14741,N_13996,N_12520);
nor U14742 (N_14742,N_13564,N_13657);
xor U14743 (N_14743,N_13522,N_13125);
xor U14744 (N_14744,N_13060,N_12777);
and U14745 (N_14745,N_13295,N_13476);
and U14746 (N_14746,N_12779,N_12412);
nor U14747 (N_14747,N_13239,N_13852);
and U14748 (N_14748,N_12530,N_13526);
and U14749 (N_14749,N_12422,N_13012);
nor U14750 (N_14750,N_12238,N_13274);
and U14751 (N_14751,N_13997,N_12794);
nor U14752 (N_14752,N_12233,N_12340);
nor U14753 (N_14753,N_13275,N_12666);
xor U14754 (N_14754,N_12158,N_13193);
and U14755 (N_14755,N_13790,N_13952);
nand U14756 (N_14756,N_12416,N_13880);
and U14757 (N_14757,N_12236,N_12194);
and U14758 (N_14758,N_12460,N_12598);
and U14759 (N_14759,N_13485,N_13670);
nand U14760 (N_14760,N_13605,N_13643);
or U14761 (N_14761,N_12868,N_12930);
nand U14762 (N_14762,N_12944,N_12214);
nor U14763 (N_14763,N_12418,N_12647);
nor U14764 (N_14764,N_12001,N_12131);
xor U14765 (N_14765,N_12814,N_13163);
or U14766 (N_14766,N_12380,N_12967);
and U14767 (N_14767,N_13652,N_12202);
xor U14768 (N_14768,N_13497,N_12398);
xor U14769 (N_14769,N_12516,N_13194);
xor U14770 (N_14770,N_13768,N_13387);
xnor U14771 (N_14771,N_12622,N_13026);
xor U14772 (N_14772,N_13796,N_12859);
nand U14773 (N_14773,N_13782,N_13935);
and U14774 (N_14774,N_12248,N_13920);
nand U14775 (N_14775,N_12465,N_13580);
or U14776 (N_14776,N_12002,N_13798);
nand U14777 (N_14777,N_12150,N_13369);
nand U14778 (N_14778,N_12585,N_12442);
and U14779 (N_14779,N_12986,N_12973);
nor U14780 (N_14780,N_12209,N_13883);
or U14781 (N_14781,N_13596,N_12995);
nor U14782 (N_14782,N_13725,N_12763);
nor U14783 (N_14783,N_12662,N_12462);
and U14784 (N_14784,N_12739,N_12796);
or U14785 (N_14785,N_12836,N_13216);
or U14786 (N_14786,N_12186,N_13739);
or U14787 (N_14787,N_12729,N_12966);
nor U14788 (N_14788,N_13201,N_13842);
or U14789 (N_14789,N_13534,N_12382);
nor U14790 (N_14790,N_13140,N_12778);
nand U14791 (N_14791,N_12533,N_13236);
and U14792 (N_14792,N_13905,N_12846);
and U14793 (N_14793,N_13161,N_13723);
or U14794 (N_14794,N_12580,N_12861);
or U14795 (N_14795,N_12389,N_12251);
nor U14796 (N_14796,N_13096,N_13423);
and U14797 (N_14797,N_13024,N_12685);
or U14798 (N_14798,N_13998,N_13001);
nor U14799 (N_14799,N_12921,N_12711);
and U14800 (N_14800,N_13443,N_12425);
nor U14801 (N_14801,N_13698,N_12175);
xnor U14802 (N_14802,N_12276,N_12275);
or U14803 (N_14803,N_13929,N_13942);
xnor U14804 (N_14804,N_13784,N_13306);
nand U14805 (N_14805,N_12845,N_12757);
and U14806 (N_14806,N_12090,N_12951);
or U14807 (N_14807,N_13260,N_12169);
xor U14808 (N_14808,N_13679,N_12665);
or U14809 (N_14809,N_12123,N_13867);
and U14810 (N_14810,N_13751,N_12498);
nor U14811 (N_14811,N_12358,N_13633);
xor U14812 (N_14812,N_13636,N_12407);
and U14813 (N_14813,N_13583,N_12193);
and U14814 (N_14814,N_12152,N_13409);
or U14815 (N_14815,N_12755,N_12941);
and U14816 (N_14816,N_13144,N_13350);
nand U14817 (N_14817,N_13215,N_12528);
or U14818 (N_14818,N_12273,N_13028);
nand U14819 (N_14819,N_12288,N_12308);
xnor U14820 (N_14820,N_13846,N_12212);
or U14821 (N_14821,N_13139,N_12674);
xor U14822 (N_14822,N_12905,N_12692);
or U14823 (N_14823,N_13507,N_12059);
nor U14824 (N_14824,N_13472,N_12679);
xor U14825 (N_14825,N_12848,N_12936);
nand U14826 (N_14826,N_12715,N_13948);
nor U14827 (N_14827,N_13251,N_12915);
xnor U14828 (N_14828,N_12524,N_12541);
nand U14829 (N_14829,N_12419,N_12684);
nor U14830 (N_14830,N_12149,N_12884);
nor U14831 (N_14831,N_12682,N_13037);
xor U14832 (N_14832,N_13979,N_13271);
nor U14833 (N_14833,N_13019,N_12488);
or U14834 (N_14834,N_13109,N_13264);
nor U14835 (N_14835,N_12046,N_13973);
nor U14836 (N_14836,N_12307,N_12369);
and U14837 (N_14837,N_12473,N_12860);
xor U14838 (N_14838,N_13076,N_12878);
nor U14839 (N_14839,N_13737,N_13442);
nand U14840 (N_14840,N_12975,N_12148);
nand U14841 (N_14841,N_13677,N_12063);
and U14842 (N_14842,N_12800,N_13279);
xnor U14843 (N_14843,N_12728,N_13543);
nor U14844 (N_14844,N_12509,N_12365);
nor U14845 (N_14845,N_12876,N_13070);
xnor U14846 (N_14846,N_13063,N_12301);
xnor U14847 (N_14847,N_12913,N_13816);
or U14848 (N_14848,N_12687,N_12918);
nand U14849 (N_14849,N_13588,N_12862);
xor U14850 (N_14850,N_12556,N_12554);
nor U14851 (N_14851,N_13671,N_13615);
nand U14852 (N_14852,N_12188,N_12118);
nand U14853 (N_14853,N_13151,N_12985);
and U14854 (N_14854,N_13786,N_12823);
xnor U14855 (N_14855,N_13586,N_12103);
and U14856 (N_14856,N_12787,N_12994);
xnor U14857 (N_14857,N_12371,N_12043);
xor U14858 (N_14858,N_12411,N_12446);
or U14859 (N_14859,N_12981,N_12855);
xor U14860 (N_14860,N_12931,N_12325);
xor U14861 (N_14861,N_12658,N_12844);
or U14862 (N_14862,N_13262,N_12073);
nand U14863 (N_14863,N_13119,N_13327);
xor U14864 (N_14864,N_12015,N_13711);
nor U14865 (N_14865,N_13308,N_12492);
nand U14866 (N_14866,N_13254,N_12590);
nor U14867 (N_14867,N_13455,N_13968);
or U14868 (N_14868,N_13928,N_13242);
nand U14869 (N_14869,N_12781,N_13726);
and U14870 (N_14870,N_12620,N_13759);
or U14871 (N_14871,N_12402,N_12893);
and U14872 (N_14872,N_12820,N_12376);
nor U14873 (N_14873,N_13086,N_12310);
xor U14874 (N_14874,N_13556,N_13991);
nand U14875 (N_14875,N_13857,N_12331);
nor U14876 (N_14876,N_12030,N_13317);
nand U14877 (N_14877,N_12788,N_12421);
and U14878 (N_14878,N_13741,N_13990);
xor U14879 (N_14879,N_12145,N_13871);
or U14880 (N_14880,N_12177,N_13433);
xor U14881 (N_14881,N_12522,N_12513);
nor U14882 (N_14882,N_13134,N_12630);
or U14883 (N_14883,N_12626,N_13284);
nand U14884 (N_14884,N_13067,N_13500);
xor U14885 (N_14885,N_12720,N_13336);
or U14886 (N_14886,N_12053,N_12423);
nor U14887 (N_14887,N_13502,N_13992);
nor U14888 (N_14888,N_13800,N_12432);
and U14889 (N_14889,N_13375,N_13544);
and U14890 (N_14890,N_12774,N_13249);
and U14891 (N_14891,N_13013,N_12808);
or U14892 (N_14892,N_12927,N_13735);
and U14893 (N_14893,N_13669,N_12261);
and U14894 (N_14894,N_13102,N_13064);
xnor U14895 (N_14895,N_13250,N_13626);
or U14896 (N_14896,N_12317,N_13227);
or U14897 (N_14897,N_12955,N_13054);
and U14898 (N_14898,N_12291,N_13848);
xnor U14899 (N_14899,N_12351,N_13354);
nor U14900 (N_14900,N_12952,N_12366);
nor U14901 (N_14901,N_12476,N_12641);
xor U14902 (N_14902,N_12443,N_12167);
nand U14903 (N_14903,N_12547,N_13205);
nor U14904 (N_14904,N_13602,N_13142);
nand U14905 (N_14905,N_12606,N_13073);
xor U14906 (N_14906,N_12464,N_13411);
nand U14907 (N_14907,N_13760,N_12281);
xor U14908 (N_14908,N_13344,N_12457);
nand U14909 (N_14909,N_12949,N_13912);
nor U14910 (N_14910,N_12360,N_12780);
xnor U14911 (N_14911,N_13100,N_13862);
or U14912 (N_14912,N_13221,N_13961);
xor U14913 (N_14913,N_13362,N_13743);
nand U14914 (N_14914,N_13623,N_13780);
nand U14915 (N_14915,N_13065,N_13661);
xnor U14916 (N_14916,N_13658,N_13468);
xor U14917 (N_14917,N_12906,N_13469);
nor U14918 (N_14918,N_12207,N_12197);
nand U14919 (N_14919,N_13058,N_12060);
xnor U14920 (N_14920,N_12119,N_13218);
xnor U14921 (N_14921,N_13890,N_13392);
xor U14922 (N_14922,N_12849,N_12189);
and U14923 (N_14923,N_13537,N_12219);
and U14924 (N_14924,N_12969,N_12032);
xor U14925 (N_14925,N_12716,N_13570);
nor U14926 (N_14926,N_13030,N_12675);
nand U14927 (N_14927,N_13341,N_12858);
nand U14928 (N_14928,N_13310,N_12987);
xnor U14929 (N_14929,N_13696,N_12919);
nor U14930 (N_14930,N_12907,N_12535);
and U14931 (N_14931,N_13114,N_13728);
or U14932 (N_14932,N_13293,N_12289);
or U14933 (N_14933,N_13092,N_12349);
and U14934 (N_14934,N_12166,N_13600);
nor U14935 (N_14935,N_13252,N_13451);
nor U14936 (N_14936,N_12260,N_13091);
or U14937 (N_14937,N_13199,N_13492);
or U14938 (N_14938,N_13039,N_13971);
or U14939 (N_14939,N_13718,N_12570);
nand U14940 (N_14940,N_13999,N_12542);
and U14941 (N_14941,N_13062,N_12680);
and U14942 (N_14942,N_13066,N_13148);
xnor U14943 (N_14943,N_12383,N_13475);
nor U14944 (N_14944,N_12162,N_13135);
or U14945 (N_14945,N_12400,N_12750);
xnor U14946 (N_14946,N_13419,N_12962);
xnor U14947 (N_14947,N_13324,N_12974);
or U14948 (N_14948,N_13266,N_13907);
nand U14949 (N_14949,N_13071,N_12313);
nor U14950 (N_14950,N_12650,N_13493);
nand U14951 (N_14951,N_13355,N_12841);
nand U14952 (N_14952,N_12526,N_12923);
or U14953 (N_14953,N_13620,N_13763);
and U14954 (N_14954,N_12051,N_13642);
and U14955 (N_14955,N_13137,N_12270);
nor U14956 (N_14956,N_12147,N_13224);
xor U14957 (N_14957,N_12009,N_13740);
nand U14958 (N_14958,N_12336,N_12076);
nor U14959 (N_14959,N_12037,N_13095);
or U14960 (N_14960,N_12429,N_12176);
xor U14961 (N_14961,N_13053,N_12274);
nor U14962 (N_14962,N_13494,N_12721);
nand U14963 (N_14963,N_12378,N_13465);
nand U14964 (N_14964,N_13712,N_12863);
nand U14965 (N_14965,N_12709,N_13653);
xor U14966 (N_14966,N_12075,N_13120);
and U14967 (N_14967,N_12256,N_13688);
nor U14968 (N_14968,N_13439,N_13363);
nand U14969 (N_14969,N_12326,N_12557);
nand U14970 (N_14970,N_13353,N_13072);
and U14971 (N_14971,N_12894,N_13518);
nor U14972 (N_14972,N_13678,N_12173);
xnor U14973 (N_14973,N_12732,N_12545);
nand U14974 (N_14974,N_13337,N_13547);
and U14975 (N_14975,N_13103,N_12088);
xnor U14976 (N_14976,N_12427,N_12151);
and U14977 (N_14977,N_12211,N_13887);
nor U14978 (N_14978,N_12776,N_12381);
or U14979 (N_14979,N_12607,N_12174);
nor U14980 (N_14980,N_12563,N_12190);
and U14981 (N_14981,N_13382,N_13732);
or U14982 (N_14982,N_13435,N_12593);
and U14983 (N_14983,N_13810,N_13351);
xnor U14984 (N_14984,N_12828,N_12198);
xor U14985 (N_14985,N_13238,N_13041);
or U14986 (N_14986,N_12436,N_12864);
and U14987 (N_14987,N_13029,N_12649);
nor U14988 (N_14988,N_13795,N_12495);
and U14989 (N_14989,N_13467,N_12178);
nor U14990 (N_14990,N_13068,N_12316);
xnor U14991 (N_14991,N_13773,N_12026);
nand U14992 (N_14992,N_12023,N_12825);
and U14993 (N_14993,N_12712,N_12268);
nor U14994 (N_14994,N_13346,N_13424);
and U14995 (N_14995,N_12587,N_13198);
xor U14996 (N_14996,N_12133,N_13960);
and U14997 (N_14997,N_12883,N_12659);
and U14998 (N_14998,N_13689,N_13444);
nor U14999 (N_14999,N_13217,N_13963);
or U15000 (N_15000,N_12965,N_12524);
nor U15001 (N_15001,N_13492,N_12412);
and U15002 (N_15002,N_12384,N_13750);
nor U15003 (N_15003,N_12092,N_12908);
xnor U15004 (N_15004,N_12914,N_12618);
nor U15005 (N_15005,N_12930,N_13212);
and U15006 (N_15006,N_12987,N_13340);
xnor U15007 (N_15007,N_12637,N_12208);
xnor U15008 (N_15008,N_12821,N_13202);
nand U15009 (N_15009,N_13027,N_12605);
nor U15010 (N_15010,N_12289,N_12985);
nand U15011 (N_15011,N_12561,N_12773);
and U15012 (N_15012,N_12283,N_13764);
and U15013 (N_15013,N_12973,N_12609);
nand U15014 (N_15014,N_13403,N_12832);
or U15015 (N_15015,N_13733,N_13086);
and U15016 (N_15016,N_12161,N_12137);
and U15017 (N_15017,N_12550,N_13637);
nand U15018 (N_15018,N_13858,N_12444);
nand U15019 (N_15019,N_13002,N_12744);
nand U15020 (N_15020,N_12046,N_12576);
nand U15021 (N_15021,N_12016,N_13353);
nor U15022 (N_15022,N_12468,N_13689);
and U15023 (N_15023,N_12169,N_12826);
nand U15024 (N_15024,N_12341,N_13543);
or U15025 (N_15025,N_13358,N_12428);
nor U15026 (N_15026,N_12708,N_13117);
nand U15027 (N_15027,N_12654,N_13400);
xor U15028 (N_15028,N_13930,N_13015);
xnor U15029 (N_15029,N_12783,N_12230);
or U15030 (N_15030,N_12460,N_13730);
and U15031 (N_15031,N_13584,N_13933);
nand U15032 (N_15032,N_12007,N_13918);
and U15033 (N_15033,N_13573,N_13071);
nand U15034 (N_15034,N_13686,N_13571);
nor U15035 (N_15035,N_13423,N_13983);
or U15036 (N_15036,N_12597,N_12591);
or U15037 (N_15037,N_12036,N_13287);
xnor U15038 (N_15038,N_12017,N_12895);
xnor U15039 (N_15039,N_13631,N_13427);
nor U15040 (N_15040,N_12048,N_12482);
nand U15041 (N_15041,N_13557,N_12530);
nor U15042 (N_15042,N_13306,N_13168);
nand U15043 (N_15043,N_13484,N_12732);
nand U15044 (N_15044,N_12617,N_12908);
nor U15045 (N_15045,N_13846,N_13954);
and U15046 (N_15046,N_13694,N_13464);
and U15047 (N_15047,N_12122,N_13984);
or U15048 (N_15048,N_13664,N_13237);
nand U15049 (N_15049,N_13258,N_13644);
nor U15050 (N_15050,N_13341,N_12628);
nand U15051 (N_15051,N_13863,N_12634);
xor U15052 (N_15052,N_13431,N_12525);
or U15053 (N_15053,N_13448,N_13105);
nor U15054 (N_15054,N_12812,N_12340);
and U15055 (N_15055,N_12602,N_12783);
or U15056 (N_15056,N_12524,N_12741);
or U15057 (N_15057,N_12635,N_12983);
nand U15058 (N_15058,N_13295,N_12440);
nand U15059 (N_15059,N_13527,N_12213);
xor U15060 (N_15060,N_13568,N_13468);
xor U15061 (N_15061,N_12267,N_13917);
nand U15062 (N_15062,N_12663,N_12581);
and U15063 (N_15063,N_13080,N_12400);
and U15064 (N_15064,N_13746,N_12828);
nor U15065 (N_15065,N_13134,N_13903);
nor U15066 (N_15066,N_13435,N_13709);
and U15067 (N_15067,N_12570,N_12372);
xnor U15068 (N_15068,N_12236,N_13123);
and U15069 (N_15069,N_13653,N_13650);
and U15070 (N_15070,N_13038,N_13004);
and U15071 (N_15071,N_12757,N_12032);
and U15072 (N_15072,N_12975,N_13197);
nor U15073 (N_15073,N_12990,N_12812);
nor U15074 (N_15074,N_13911,N_13274);
nor U15075 (N_15075,N_12261,N_12880);
xor U15076 (N_15076,N_13266,N_13695);
nand U15077 (N_15077,N_13806,N_12876);
and U15078 (N_15078,N_13862,N_12231);
nor U15079 (N_15079,N_13878,N_12330);
xnor U15080 (N_15080,N_13429,N_13695);
xnor U15081 (N_15081,N_12365,N_12403);
xnor U15082 (N_15082,N_13690,N_12598);
nand U15083 (N_15083,N_12979,N_13154);
and U15084 (N_15084,N_12280,N_13300);
nor U15085 (N_15085,N_13847,N_13481);
nor U15086 (N_15086,N_13384,N_12799);
xor U15087 (N_15087,N_13268,N_13137);
or U15088 (N_15088,N_13688,N_12503);
and U15089 (N_15089,N_13287,N_13028);
xor U15090 (N_15090,N_13317,N_13845);
and U15091 (N_15091,N_13154,N_13889);
and U15092 (N_15092,N_13872,N_13533);
nor U15093 (N_15093,N_12392,N_13202);
xor U15094 (N_15094,N_12514,N_12138);
xor U15095 (N_15095,N_12880,N_13452);
or U15096 (N_15096,N_13897,N_13612);
nand U15097 (N_15097,N_13263,N_13054);
and U15098 (N_15098,N_12871,N_13553);
nor U15099 (N_15099,N_13913,N_12023);
and U15100 (N_15100,N_13355,N_13878);
nand U15101 (N_15101,N_12174,N_13488);
or U15102 (N_15102,N_13076,N_12052);
or U15103 (N_15103,N_13534,N_13330);
xnor U15104 (N_15104,N_13949,N_12378);
nand U15105 (N_15105,N_12140,N_12575);
xnor U15106 (N_15106,N_13022,N_13626);
xnor U15107 (N_15107,N_13164,N_12965);
or U15108 (N_15108,N_13580,N_13220);
nand U15109 (N_15109,N_12771,N_13779);
and U15110 (N_15110,N_13540,N_13530);
nor U15111 (N_15111,N_12084,N_12663);
nor U15112 (N_15112,N_13971,N_13205);
nand U15113 (N_15113,N_13630,N_13930);
nand U15114 (N_15114,N_12103,N_13529);
nor U15115 (N_15115,N_12623,N_12169);
nor U15116 (N_15116,N_12361,N_13467);
or U15117 (N_15117,N_13921,N_12241);
nand U15118 (N_15118,N_13769,N_12760);
xnor U15119 (N_15119,N_13349,N_13633);
xnor U15120 (N_15120,N_13029,N_12297);
or U15121 (N_15121,N_12384,N_12207);
nor U15122 (N_15122,N_13635,N_13454);
nor U15123 (N_15123,N_12357,N_13641);
and U15124 (N_15124,N_13471,N_12439);
nand U15125 (N_15125,N_13255,N_12883);
nand U15126 (N_15126,N_13522,N_13000);
nor U15127 (N_15127,N_12348,N_13122);
nand U15128 (N_15128,N_13940,N_13558);
or U15129 (N_15129,N_13826,N_13567);
nor U15130 (N_15130,N_13981,N_13408);
nand U15131 (N_15131,N_13631,N_13063);
nor U15132 (N_15132,N_13015,N_12657);
and U15133 (N_15133,N_12899,N_12225);
xor U15134 (N_15134,N_13120,N_12682);
nor U15135 (N_15135,N_13652,N_13749);
xor U15136 (N_15136,N_13824,N_13121);
xor U15137 (N_15137,N_12028,N_12291);
or U15138 (N_15138,N_13584,N_12736);
or U15139 (N_15139,N_12903,N_12478);
xor U15140 (N_15140,N_12562,N_12325);
or U15141 (N_15141,N_13368,N_12721);
xnor U15142 (N_15142,N_12009,N_13256);
nand U15143 (N_15143,N_13458,N_13492);
xor U15144 (N_15144,N_13433,N_13355);
and U15145 (N_15145,N_12828,N_12631);
nand U15146 (N_15146,N_12016,N_13160);
nor U15147 (N_15147,N_12262,N_13000);
nor U15148 (N_15148,N_13550,N_12007);
or U15149 (N_15149,N_12437,N_12286);
nand U15150 (N_15150,N_13688,N_12187);
or U15151 (N_15151,N_12250,N_12821);
nand U15152 (N_15152,N_13036,N_12244);
nor U15153 (N_15153,N_13037,N_12430);
or U15154 (N_15154,N_12820,N_12160);
and U15155 (N_15155,N_13795,N_13576);
xor U15156 (N_15156,N_12055,N_12490);
nor U15157 (N_15157,N_12934,N_13283);
or U15158 (N_15158,N_13111,N_12630);
nand U15159 (N_15159,N_13826,N_12761);
or U15160 (N_15160,N_12016,N_12221);
nor U15161 (N_15161,N_13559,N_12829);
nor U15162 (N_15162,N_13035,N_12746);
nand U15163 (N_15163,N_12170,N_12010);
nand U15164 (N_15164,N_12376,N_13035);
nand U15165 (N_15165,N_13652,N_12824);
xnor U15166 (N_15166,N_13846,N_12777);
and U15167 (N_15167,N_13332,N_13821);
and U15168 (N_15168,N_13077,N_13483);
or U15169 (N_15169,N_13804,N_12328);
nor U15170 (N_15170,N_12521,N_12177);
xnor U15171 (N_15171,N_12828,N_12097);
or U15172 (N_15172,N_12941,N_12092);
nand U15173 (N_15173,N_13006,N_13911);
xor U15174 (N_15174,N_13961,N_13663);
nor U15175 (N_15175,N_12003,N_13552);
nand U15176 (N_15176,N_13321,N_13120);
nand U15177 (N_15177,N_12153,N_12448);
nand U15178 (N_15178,N_12647,N_12986);
or U15179 (N_15179,N_13595,N_13329);
nor U15180 (N_15180,N_13249,N_12773);
and U15181 (N_15181,N_12736,N_12720);
nor U15182 (N_15182,N_13845,N_12163);
or U15183 (N_15183,N_13202,N_12005);
nor U15184 (N_15184,N_12845,N_13491);
xor U15185 (N_15185,N_13886,N_12897);
xnor U15186 (N_15186,N_12644,N_12046);
xor U15187 (N_15187,N_12419,N_13000);
xor U15188 (N_15188,N_13107,N_13273);
or U15189 (N_15189,N_13111,N_13317);
and U15190 (N_15190,N_13897,N_13381);
or U15191 (N_15191,N_13882,N_12589);
and U15192 (N_15192,N_13854,N_13075);
nand U15193 (N_15193,N_12810,N_12853);
nand U15194 (N_15194,N_12176,N_12922);
and U15195 (N_15195,N_12078,N_12005);
xnor U15196 (N_15196,N_12797,N_13199);
nand U15197 (N_15197,N_12283,N_13454);
and U15198 (N_15198,N_12797,N_12988);
or U15199 (N_15199,N_13808,N_13741);
and U15200 (N_15200,N_12218,N_13936);
xnor U15201 (N_15201,N_12970,N_12348);
nand U15202 (N_15202,N_12997,N_12014);
or U15203 (N_15203,N_12221,N_13464);
nor U15204 (N_15204,N_12684,N_12298);
xor U15205 (N_15205,N_12490,N_12255);
nor U15206 (N_15206,N_13794,N_12541);
or U15207 (N_15207,N_12948,N_13981);
nor U15208 (N_15208,N_12550,N_13269);
nand U15209 (N_15209,N_13093,N_13725);
or U15210 (N_15210,N_13749,N_13866);
and U15211 (N_15211,N_13319,N_13090);
or U15212 (N_15212,N_12653,N_13569);
and U15213 (N_15213,N_12756,N_12883);
nor U15214 (N_15214,N_13010,N_13257);
and U15215 (N_15215,N_12588,N_13701);
nand U15216 (N_15216,N_12110,N_12048);
or U15217 (N_15217,N_13320,N_13631);
and U15218 (N_15218,N_13315,N_12115);
and U15219 (N_15219,N_13605,N_13629);
nand U15220 (N_15220,N_13866,N_13313);
and U15221 (N_15221,N_13724,N_12639);
nor U15222 (N_15222,N_13598,N_13942);
nand U15223 (N_15223,N_12273,N_12928);
or U15224 (N_15224,N_13795,N_13547);
nor U15225 (N_15225,N_12368,N_13111);
nand U15226 (N_15226,N_13825,N_12190);
nand U15227 (N_15227,N_13685,N_13004);
and U15228 (N_15228,N_13699,N_13177);
and U15229 (N_15229,N_13313,N_13021);
or U15230 (N_15230,N_13398,N_12125);
xor U15231 (N_15231,N_12508,N_13673);
nand U15232 (N_15232,N_12893,N_13971);
nor U15233 (N_15233,N_13556,N_12354);
and U15234 (N_15234,N_13253,N_13237);
xor U15235 (N_15235,N_12485,N_12026);
or U15236 (N_15236,N_13367,N_12322);
and U15237 (N_15237,N_13175,N_12552);
xor U15238 (N_15238,N_13323,N_12175);
nand U15239 (N_15239,N_13494,N_13008);
nand U15240 (N_15240,N_12157,N_12239);
or U15241 (N_15241,N_12096,N_13470);
nand U15242 (N_15242,N_12910,N_12170);
or U15243 (N_15243,N_12239,N_12864);
or U15244 (N_15244,N_12485,N_12908);
nand U15245 (N_15245,N_12076,N_13077);
xor U15246 (N_15246,N_13945,N_12777);
and U15247 (N_15247,N_13947,N_13115);
or U15248 (N_15248,N_13494,N_12666);
and U15249 (N_15249,N_13759,N_12244);
nand U15250 (N_15250,N_12245,N_12612);
nor U15251 (N_15251,N_13688,N_13493);
xnor U15252 (N_15252,N_12803,N_12969);
and U15253 (N_15253,N_13888,N_12317);
nor U15254 (N_15254,N_12091,N_13181);
nand U15255 (N_15255,N_13227,N_13126);
nor U15256 (N_15256,N_13711,N_13762);
nand U15257 (N_15257,N_13994,N_12579);
or U15258 (N_15258,N_13672,N_13684);
and U15259 (N_15259,N_12990,N_12013);
or U15260 (N_15260,N_12006,N_13834);
nand U15261 (N_15261,N_13988,N_13254);
or U15262 (N_15262,N_13834,N_13061);
nor U15263 (N_15263,N_13426,N_12929);
and U15264 (N_15264,N_13258,N_12370);
or U15265 (N_15265,N_12731,N_12358);
xnor U15266 (N_15266,N_12441,N_12118);
xor U15267 (N_15267,N_13729,N_12602);
xor U15268 (N_15268,N_13956,N_13142);
nor U15269 (N_15269,N_13127,N_12806);
nand U15270 (N_15270,N_13404,N_13670);
and U15271 (N_15271,N_12795,N_13734);
or U15272 (N_15272,N_13236,N_12579);
nand U15273 (N_15273,N_12963,N_12829);
and U15274 (N_15274,N_12800,N_13268);
nor U15275 (N_15275,N_13749,N_13357);
nand U15276 (N_15276,N_12166,N_13492);
nor U15277 (N_15277,N_13520,N_13507);
or U15278 (N_15278,N_13178,N_12556);
nor U15279 (N_15279,N_12941,N_13348);
and U15280 (N_15280,N_12078,N_13319);
or U15281 (N_15281,N_13900,N_12144);
nand U15282 (N_15282,N_13046,N_13952);
xnor U15283 (N_15283,N_12719,N_13172);
xor U15284 (N_15284,N_13096,N_13051);
xor U15285 (N_15285,N_12982,N_12986);
xor U15286 (N_15286,N_12113,N_12518);
and U15287 (N_15287,N_13544,N_12809);
xnor U15288 (N_15288,N_12776,N_13595);
and U15289 (N_15289,N_12773,N_12052);
nor U15290 (N_15290,N_13955,N_13672);
or U15291 (N_15291,N_13879,N_13926);
nand U15292 (N_15292,N_12572,N_13260);
and U15293 (N_15293,N_12461,N_13859);
xor U15294 (N_15294,N_12675,N_13722);
and U15295 (N_15295,N_13418,N_12936);
or U15296 (N_15296,N_13355,N_13294);
and U15297 (N_15297,N_13967,N_13162);
nor U15298 (N_15298,N_12855,N_12493);
xnor U15299 (N_15299,N_12080,N_13996);
xor U15300 (N_15300,N_13106,N_13119);
nand U15301 (N_15301,N_12672,N_13734);
xor U15302 (N_15302,N_13339,N_12831);
or U15303 (N_15303,N_13367,N_13104);
or U15304 (N_15304,N_12272,N_12765);
nand U15305 (N_15305,N_12023,N_12701);
and U15306 (N_15306,N_13707,N_12622);
nor U15307 (N_15307,N_12900,N_12970);
nor U15308 (N_15308,N_13438,N_12417);
nor U15309 (N_15309,N_12467,N_12634);
or U15310 (N_15310,N_13746,N_12201);
xor U15311 (N_15311,N_12217,N_13866);
xor U15312 (N_15312,N_13434,N_12550);
nand U15313 (N_15313,N_13687,N_12231);
nor U15314 (N_15314,N_12365,N_13786);
and U15315 (N_15315,N_12228,N_13226);
nor U15316 (N_15316,N_12353,N_13492);
nand U15317 (N_15317,N_12130,N_13994);
or U15318 (N_15318,N_12461,N_12671);
nor U15319 (N_15319,N_12098,N_12180);
nand U15320 (N_15320,N_13692,N_13773);
and U15321 (N_15321,N_13333,N_13201);
nor U15322 (N_15322,N_12383,N_12353);
and U15323 (N_15323,N_12377,N_13981);
nor U15324 (N_15324,N_12723,N_13885);
or U15325 (N_15325,N_12986,N_12974);
or U15326 (N_15326,N_12442,N_12757);
and U15327 (N_15327,N_13921,N_12191);
and U15328 (N_15328,N_12596,N_12263);
and U15329 (N_15329,N_12005,N_12956);
nor U15330 (N_15330,N_13012,N_12548);
or U15331 (N_15331,N_12433,N_13528);
nand U15332 (N_15332,N_13157,N_12366);
nand U15333 (N_15333,N_12891,N_13711);
xnor U15334 (N_15334,N_12828,N_13444);
or U15335 (N_15335,N_13320,N_13703);
nand U15336 (N_15336,N_13666,N_13188);
nand U15337 (N_15337,N_13485,N_13539);
nor U15338 (N_15338,N_13394,N_12396);
nand U15339 (N_15339,N_13572,N_12878);
xor U15340 (N_15340,N_13866,N_13542);
nor U15341 (N_15341,N_12189,N_13790);
and U15342 (N_15342,N_12903,N_13708);
xor U15343 (N_15343,N_13568,N_13310);
nand U15344 (N_15344,N_12474,N_12385);
nor U15345 (N_15345,N_12384,N_12513);
xor U15346 (N_15346,N_13793,N_13431);
nor U15347 (N_15347,N_13196,N_13834);
or U15348 (N_15348,N_12799,N_13336);
xnor U15349 (N_15349,N_13470,N_13702);
xor U15350 (N_15350,N_12792,N_12919);
nand U15351 (N_15351,N_12299,N_13451);
nand U15352 (N_15352,N_12072,N_13075);
and U15353 (N_15353,N_13291,N_13298);
xor U15354 (N_15354,N_13271,N_13105);
nand U15355 (N_15355,N_13879,N_12564);
nand U15356 (N_15356,N_12518,N_13419);
xor U15357 (N_15357,N_12199,N_13295);
nor U15358 (N_15358,N_12047,N_12718);
nand U15359 (N_15359,N_13103,N_13328);
and U15360 (N_15360,N_12317,N_12632);
and U15361 (N_15361,N_13172,N_12974);
xor U15362 (N_15362,N_13770,N_13371);
or U15363 (N_15363,N_13681,N_12539);
nand U15364 (N_15364,N_13554,N_12640);
nand U15365 (N_15365,N_13975,N_13300);
and U15366 (N_15366,N_13388,N_12383);
nand U15367 (N_15367,N_12395,N_13263);
xor U15368 (N_15368,N_13107,N_12845);
and U15369 (N_15369,N_12824,N_13223);
or U15370 (N_15370,N_13329,N_13260);
or U15371 (N_15371,N_13516,N_12413);
or U15372 (N_15372,N_13407,N_13578);
nand U15373 (N_15373,N_13038,N_12696);
or U15374 (N_15374,N_12157,N_13579);
or U15375 (N_15375,N_13032,N_13804);
nand U15376 (N_15376,N_12365,N_13799);
and U15377 (N_15377,N_13846,N_13360);
or U15378 (N_15378,N_12012,N_13448);
nor U15379 (N_15379,N_13749,N_12296);
xor U15380 (N_15380,N_12137,N_13279);
nand U15381 (N_15381,N_12398,N_12322);
nand U15382 (N_15382,N_12880,N_12745);
xor U15383 (N_15383,N_12654,N_13291);
and U15384 (N_15384,N_13639,N_12562);
nor U15385 (N_15385,N_13994,N_13428);
nor U15386 (N_15386,N_13057,N_13085);
nor U15387 (N_15387,N_12667,N_12392);
xnor U15388 (N_15388,N_12983,N_12719);
and U15389 (N_15389,N_12601,N_13988);
nor U15390 (N_15390,N_12679,N_13002);
nand U15391 (N_15391,N_12648,N_12654);
nand U15392 (N_15392,N_13048,N_12626);
nand U15393 (N_15393,N_13893,N_13516);
and U15394 (N_15394,N_13812,N_12438);
or U15395 (N_15395,N_12727,N_13234);
or U15396 (N_15396,N_13298,N_12919);
and U15397 (N_15397,N_13273,N_13762);
xnor U15398 (N_15398,N_12770,N_12072);
and U15399 (N_15399,N_13878,N_12278);
nor U15400 (N_15400,N_12498,N_13616);
xor U15401 (N_15401,N_13540,N_13085);
nor U15402 (N_15402,N_13704,N_12558);
xnor U15403 (N_15403,N_13049,N_12045);
nor U15404 (N_15404,N_13230,N_12223);
nand U15405 (N_15405,N_12655,N_12104);
nor U15406 (N_15406,N_13226,N_12763);
nand U15407 (N_15407,N_12147,N_13913);
nor U15408 (N_15408,N_12502,N_12480);
xor U15409 (N_15409,N_12336,N_13496);
xor U15410 (N_15410,N_13956,N_13106);
or U15411 (N_15411,N_13891,N_13976);
nand U15412 (N_15412,N_13883,N_13980);
nor U15413 (N_15413,N_12545,N_13027);
or U15414 (N_15414,N_13928,N_12136);
or U15415 (N_15415,N_13285,N_12160);
xnor U15416 (N_15416,N_12443,N_12123);
nor U15417 (N_15417,N_13408,N_12888);
nor U15418 (N_15418,N_12646,N_12366);
nor U15419 (N_15419,N_13545,N_13376);
and U15420 (N_15420,N_13517,N_13796);
and U15421 (N_15421,N_13939,N_12185);
and U15422 (N_15422,N_13139,N_12503);
or U15423 (N_15423,N_13367,N_12461);
or U15424 (N_15424,N_13680,N_12167);
xnor U15425 (N_15425,N_13356,N_12244);
or U15426 (N_15426,N_13951,N_13875);
or U15427 (N_15427,N_13119,N_12759);
and U15428 (N_15428,N_12371,N_13005);
or U15429 (N_15429,N_13030,N_12797);
and U15430 (N_15430,N_13441,N_13580);
xor U15431 (N_15431,N_12938,N_12249);
xor U15432 (N_15432,N_12432,N_12398);
and U15433 (N_15433,N_13236,N_13381);
and U15434 (N_15434,N_13144,N_12759);
nor U15435 (N_15435,N_13096,N_12435);
xnor U15436 (N_15436,N_12218,N_12361);
nand U15437 (N_15437,N_12166,N_13704);
nor U15438 (N_15438,N_13021,N_12381);
xor U15439 (N_15439,N_13282,N_13450);
xnor U15440 (N_15440,N_12487,N_12243);
xor U15441 (N_15441,N_12569,N_12779);
and U15442 (N_15442,N_13900,N_13876);
or U15443 (N_15443,N_13337,N_13328);
or U15444 (N_15444,N_12492,N_12587);
xor U15445 (N_15445,N_12175,N_13082);
xor U15446 (N_15446,N_13959,N_12289);
nor U15447 (N_15447,N_12605,N_13454);
xor U15448 (N_15448,N_13898,N_13097);
or U15449 (N_15449,N_12961,N_12211);
nand U15450 (N_15450,N_13609,N_13025);
nand U15451 (N_15451,N_12341,N_12210);
nand U15452 (N_15452,N_12436,N_13983);
or U15453 (N_15453,N_12617,N_12570);
xor U15454 (N_15454,N_13081,N_12476);
nor U15455 (N_15455,N_12451,N_12784);
nand U15456 (N_15456,N_12780,N_13136);
or U15457 (N_15457,N_13532,N_12422);
nor U15458 (N_15458,N_12068,N_12528);
nand U15459 (N_15459,N_13280,N_13505);
or U15460 (N_15460,N_13523,N_13206);
xor U15461 (N_15461,N_12958,N_13131);
or U15462 (N_15462,N_13722,N_12923);
and U15463 (N_15463,N_13183,N_13836);
xor U15464 (N_15464,N_12999,N_12144);
nor U15465 (N_15465,N_12571,N_13673);
or U15466 (N_15466,N_13334,N_13346);
or U15467 (N_15467,N_13378,N_12927);
and U15468 (N_15468,N_12992,N_13117);
and U15469 (N_15469,N_12243,N_13429);
nor U15470 (N_15470,N_12827,N_13329);
or U15471 (N_15471,N_12506,N_13687);
or U15472 (N_15472,N_12610,N_13131);
or U15473 (N_15473,N_12849,N_13705);
nor U15474 (N_15474,N_13272,N_12491);
xnor U15475 (N_15475,N_13036,N_13755);
xor U15476 (N_15476,N_13919,N_12259);
or U15477 (N_15477,N_13150,N_13764);
xor U15478 (N_15478,N_13143,N_13240);
or U15479 (N_15479,N_12304,N_13325);
and U15480 (N_15480,N_12158,N_13666);
nand U15481 (N_15481,N_13449,N_12822);
nor U15482 (N_15482,N_13349,N_12137);
xor U15483 (N_15483,N_13237,N_12498);
or U15484 (N_15484,N_13060,N_13826);
and U15485 (N_15485,N_12876,N_12403);
nor U15486 (N_15486,N_12102,N_13607);
nand U15487 (N_15487,N_13571,N_12034);
nand U15488 (N_15488,N_13436,N_12935);
nand U15489 (N_15489,N_12335,N_13570);
xor U15490 (N_15490,N_12008,N_13156);
nand U15491 (N_15491,N_13869,N_12007);
or U15492 (N_15492,N_12817,N_13683);
nand U15493 (N_15493,N_12046,N_12579);
nor U15494 (N_15494,N_12688,N_13844);
nor U15495 (N_15495,N_13588,N_13687);
nor U15496 (N_15496,N_12449,N_13892);
and U15497 (N_15497,N_12696,N_13820);
and U15498 (N_15498,N_13919,N_13358);
and U15499 (N_15499,N_13826,N_12126);
nand U15500 (N_15500,N_12468,N_12347);
nor U15501 (N_15501,N_13456,N_12767);
xnor U15502 (N_15502,N_13094,N_13916);
nor U15503 (N_15503,N_13788,N_12378);
nor U15504 (N_15504,N_12036,N_13451);
xor U15505 (N_15505,N_12917,N_13218);
nor U15506 (N_15506,N_13380,N_13022);
xnor U15507 (N_15507,N_13604,N_13086);
and U15508 (N_15508,N_12091,N_13785);
xor U15509 (N_15509,N_12789,N_12571);
nor U15510 (N_15510,N_13688,N_12701);
nor U15511 (N_15511,N_12283,N_12994);
xor U15512 (N_15512,N_12592,N_12691);
and U15513 (N_15513,N_12626,N_12052);
nor U15514 (N_15514,N_12041,N_12064);
nor U15515 (N_15515,N_12256,N_13032);
and U15516 (N_15516,N_12004,N_13074);
xor U15517 (N_15517,N_12565,N_12101);
nor U15518 (N_15518,N_12131,N_13389);
or U15519 (N_15519,N_13116,N_13435);
xnor U15520 (N_15520,N_12296,N_13199);
nor U15521 (N_15521,N_13616,N_12046);
nand U15522 (N_15522,N_12892,N_13773);
nand U15523 (N_15523,N_12884,N_12848);
or U15524 (N_15524,N_12857,N_13503);
xnor U15525 (N_15525,N_13401,N_13302);
nor U15526 (N_15526,N_13735,N_12679);
xor U15527 (N_15527,N_13534,N_12316);
nand U15528 (N_15528,N_12197,N_13155);
nor U15529 (N_15529,N_13809,N_13281);
nand U15530 (N_15530,N_13810,N_13896);
xor U15531 (N_15531,N_13944,N_12079);
xor U15532 (N_15532,N_13430,N_13753);
xnor U15533 (N_15533,N_13350,N_12949);
nor U15534 (N_15534,N_12047,N_13971);
or U15535 (N_15535,N_12082,N_12427);
nor U15536 (N_15536,N_12774,N_12832);
or U15537 (N_15537,N_12380,N_12371);
nand U15538 (N_15538,N_13792,N_12492);
xor U15539 (N_15539,N_13523,N_13622);
nor U15540 (N_15540,N_12966,N_12557);
xor U15541 (N_15541,N_13211,N_13806);
or U15542 (N_15542,N_12450,N_13647);
or U15543 (N_15543,N_13693,N_13454);
nor U15544 (N_15544,N_13461,N_12780);
nand U15545 (N_15545,N_12311,N_13682);
and U15546 (N_15546,N_12825,N_13213);
nor U15547 (N_15547,N_13177,N_12434);
nand U15548 (N_15548,N_13869,N_13072);
xnor U15549 (N_15549,N_12418,N_13814);
or U15550 (N_15550,N_12585,N_12751);
xnor U15551 (N_15551,N_12476,N_12701);
nor U15552 (N_15552,N_13906,N_13578);
nor U15553 (N_15553,N_12239,N_13390);
nor U15554 (N_15554,N_12842,N_12856);
nor U15555 (N_15555,N_12504,N_12119);
and U15556 (N_15556,N_13063,N_13987);
or U15557 (N_15557,N_12649,N_12103);
or U15558 (N_15558,N_13032,N_13130);
nand U15559 (N_15559,N_12900,N_12808);
nand U15560 (N_15560,N_12066,N_13389);
nor U15561 (N_15561,N_13342,N_12313);
and U15562 (N_15562,N_13647,N_12599);
xor U15563 (N_15563,N_13643,N_13823);
or U15564 (N_15564,N_13273,N_12425);
or U15565 (N_15565,N_13288,N_12612);
xor U15566 (N_15566,N_12393,N_12798);
nand U15567 (N_15567,N_13914,N_12396);
and U15568 (N_15568,N_12314,N_13771);
xnor U15569 (N_15569,N_12577,N_12346);
and U15570 (N_15570,N_13650,N_12210);
nand U15571 (N_15571,N_13360,N_13359);
or U15572 (N_15572,N_13537,N_12838);
and U15573 (N_15573,N_12067,N_12983);
nand U15574 (N_15574,N_12838,N_13354);
xnor U15575 (N_15575,N_13882,N_12327);
xnor U15576 (N_15576,N_12910,N_12852);
and U15577 (N_15577,N_13689,N_12007);
xor U15578 (N_15578,N_12956,N_12157);
nor U15579 (N_15579,N_12102,N_13268);
and U15580 (N_15580,N_12887,N_12529);
and U15581 (N_15581,N_13374,N_12083);
xnor U15582 (N_15582,N_13909,N_13458);
nor U15583 (N_15583,N_12979,N_12161);
nor U15584 (N_15584,N_12275,N_13837);
nand U15585 (N_15585,N_13641,N_12878);
nand U15586 (N_15586,N_13290,N_12200);
and U15587 (N_15587,N_13840,N_13414);
nor U15588 (N_15588,N_12965,N_13839);
nor U15589 (N_15589,N_12366,N_13734);
xnor U15590 (N_15590,N_13440,N_12320);
or U15591 (N_15591,N_12184,N_13128);
nand U15592 (N_15592,N_13996,N_12851);
and U15593 (N_15593,N_12813,N_13934);
and U15594 (N_15594,N_12396,N_13483);
and U15595 (N_15595,N_12866,N_12625);
and U15596 (N_15596,N_12774,N_13403);
and U15597 (N_15597,N_13042,N_12864);
xnor U15598 (N_15598,N_13572,N_13500);
or U15599 (N_15599,N_12898,N_12328);
nand U15600 (N_15600,N_12146,N_13524);
or U15601 (N_15601,N_12174,N_12500);
and U15602 (N_15602,N_13895,N_13105);
and U15603 (N_15603,N_12261,N_13414);
or U15604 (N_15604,N_13819,N_12015);
xnor U15605 (N_15605,N_13609,N_12220);
nand U15606 (N_15606,N_13498,N_12341);
xor U15607 (N_15607,N_12704,N_12352);
xnor U15608 (N_15608,N_12359,N_12156);
or U15609 (N_15609,N_13847,N_13795);
nor U15610 (N_15610,N_13009,N_13119);
nor U15611 (N_15611,N_12466,N_12318);
xor U15612 (N_15612,N_12321,N_13699);
nor U15613 (N_15613,N_13846,N_12760);
nand U15614 (N_15614,N_13500,N_13362);
xor U15615 (N_15615,N_13614,N_13895);
and U15616 (N_15616,N_12800,N_12420);
xor U15617 (N_15617,N_12085,N_13639);
and U15618 (N_15618,N_13500,N_13832);
nand U15619 (N_15619,N_13830,N_13994);
nor U15620 (N_15620,N_13937,N_13098);
xnor U15621 (N_15621,N_12054,N_13820);
nor U15622 (N_15622,N_13562,N_12868);
and U15623 (N_15623,N_13968,N_12630);
or U15624 (N_15624,N_13523,N_12216);
xor U15625 (N_15625,N_13235,N_13512);
or U15626 (N_15626,N_13509,N_12814);
and U15627 (N_15627,N_13622,N_12349);
nor U15628 (N_15628,N_13956,N_12348);
or U15629 (N_15629,N_12331,N_12667);
nand U15630 (N_15630,N_12432,N_12185);
and U15631 (N_15631,N_12117,N_13817);
and U15632 (N_15632,N_13104,N_12442);
xor U15633 (N_15633,N_12451,N_12755);
nand U15634 (N_15634,N_13164,N_12934);
or U15635 (N_15635,N_12900,N_13036);
nand U15636 (N_15636,N_13075,N_13946);
nand U15637 (N_15637,N_12837,N_13728);
xor U15638 (N_15638,N_12762,N_12268);
and U15639 (N_15639,N_12898,N_13401);
and U15640 (N_15640,N_12916,N_13778);
xor U15641 (N_15641,N_12886,N_13973);
and U15642 (N_15642,N_13537,N_13958);
nand U15643 (N_15643,N_13732,N_12257);
and U15644 (N_15644,N_12277,N_12538);
and U15645 (N_15645,N_12773,N_12221);
and U15646 (N_15646,N_13179,N_12653);
nor U15647 (N_15647,N_12151,N_13796);
nor U15648 (N_15648,N_12616,N_12214);
nor U15649 (N_15649,N_13851,N_12363);
or U15650 (N_15650,N_13986,N_13884);
nor U15651 (N_15651,N_13146,N_13557);
nor U15652 (N_15652,N_12154,N_13459);
nor U15653 (N_15653,N_13881,N_13622);
xor U15654 (N_15654,N_12858,N_13367);
or U15655 (N_15655,N_12862,N_12601);
and U15656 (N_15656,N_13820,N_13789);
nand U15657 (N_15657,N_12370,N_13211);
nand U15658 (N_15658,N_12147,N_12954);
and U15659 (N_15659,N_12485,N_13907);
or U15660 (N_15660,N_13464,N_12001);
nand U15661 (N_15661,N_12704,N_12633);
nor U15662 (N_15662,N_13063,N_13296);
nand U15663 (N_15663,N_13301,N_12032);
nor U15664 (N_15664,N_12386,N_13728);
nor U15665 (N_15665,N_12422,N_13672);
or U15666 (N_15666,N_12761,N_13249);
nand U15667 (N_15667,N_13510,N_13465);
or U15668 (N_15668,N_12416,N_12823);
and U15669 (N_15669,N_13521,N_12084);
or U15670 (N_15670,N_13170,N_13847);
nor U15671 (N_15671,N_13898,N_12717);
and U15672 (N_15672,N_12552,N_13701);
or U15673 (N_15673,N_12449,N_12295);
xnor U15674 (N_15674,N_12106,N_13073);
nand U15675 (N_15675,N_12859,N_13513);
xor U15676 (N_15676,N_12903,N_12735);
or U15677 (N_15677,N_12240,N_13359);
nor U15678 (N_15678,N_13089,N_13583);
nor U15679 (N_15679,N_13284,N_13068);
and U15680 (N_15680,N_12552,N_13037);
and U15681 (N_15681,N_13672,N_12370);
and U15682 (N_15682,N_12994,N_13698);
nor U15683 (N_15683,N_12468,N_13438);
nand U15684 (N_15684,N_13024,N_12529);
nor U15685 (N_15685,N_12790,N_12640);
xor U15686 (N_15686,N_13560,N_12599);
nand U15687 (N_15687,N_12696,N_13756);
nor U15688 (N_15688,N_13510,N_12930);
nand U15689 (N_15689,N_13516,N_12785);
xor U15690 (N_15690,N_12653,N_13906);
nor U15691 (N_15691,N_12989,N_12997);
or U15692 (N_15692,N_13867,N_12106);
xor U15693 (N_15693,N_12422,N_13669);
nor U15694 (N_15694,N_12382,N_13367);
xor U15695 (N_15695,N_13169,N_12447);
xnor U15696 (N_15696,N_12399,N_12290);
nand U15697 (N_15697,N_13964,N_13561);
nand U15698 (N_15698,N_12878,N_13347);
and U15699 (N_15699,N_12334,N_13183);
and U15700 (N_15700,N_13255,N_12788);
or U15701 (N_15701,N_12474,N_13407);
xor U15702 (N_15702,N_12668,N_13591);
xor U15703 (N_15703,N_13634,N_13492);
nor U15704 (N_15704,N_12870,N_12368);
nand U15705 (N_15705,N_13498,N_12024);
or U15706 (N_15706,N_13185,N_13778);
nand U15707 (N_15707,N_13344,N_12646);
nand U15708 (N_15708,N_13768,N_13682);
nand U15709 (N_15709,N_13759,N_12032);
xnor U15710 (N_15710,N_12840,N_12371);
or U15711 (N_15711,N_13244,N_12760);
nor U15712 (N_15712,N_13535,N_12747);
nand U15713 (N_15713,N_12088,N_13784);
nand U15714 (N_15714,N_13772,N_13927);
nand U15715 (N_15715,N_13032,N_12821);
nor U15716 (N_15716,N_13811,N_12860);
nand U15717 (N_15717,N_13219,N_13875);
nand U15718 (N_15718,N_13458,N_13548);
or U15719 (N_15719,N_12434,N_12549);
nor U15720 (N_15720,N_13611,N_13900);
nand U15721 (N_15721,N_12858,N_13695);
and U15722 (N_15722,N_13409,N_13847);
or U15723 (N_15723,N_12642,N_13092);
and U15724 (N_15724,N_12032,N_12336);
xnor U15725 (N_15725,N_13059,N_12724);
or U15726 (N_15726,N_12770,N_12256);
nor U15727 (N_15727,N_13186,N_12307);
nand U15728 (N_15728,N_12436,N_13271);
nor U15729 (N_15729,N_13583,N_13069);
or U15730 (N_15730,N_12186,N_13163);
nand U15731 (N_15731,N_13051,N_13311);
nand U15732 (N_15732,N_12380,N_12028);
xor U15733 (N_15733,N_12032,N_13657);
xor U15734 (N_15734,N_12403,N_13302);
nand U15735 (N_15735,N_12527,N_13175);
nor U15736 (N_15736,N_13072,N_13663);
nor U15737 (N_15737,N_12353,N_13233);
or U15738 (N_15738,N_13975,N_13586);
and U15739 (N_15739,N_13049,N_13468);
nand U15740 (N_15740,N_12189,N_13209);
and U15741 (N_15741,N_13167,N_12799);
nand U15742 (N_15742,N_13622,N_12646);
nand U15743 (N_15743,N_13695,N_13955);
and U15744 (N_15744,N_13180,N_12152);
and U15745 (N_15745,N_13532,N_12206);
nand U15746 (N_15746,N_12515,N_13977);
nand U15747 (N_15747,N_12740,N_13661);
and U15748 (N_15748,N_13466,N_12969);
xnor U15749 (N_15749,N_13081,N_12501);
nand U15750 (N_15750,N_12856,N_13210);
or U15751 (N_15751,N_12007,N_12925);
nand U15752 (N_15752,N_12865,N_12024);
nand U15753 (N_15753,N_12420,N_12958);
nand U15754 (N_15754,N_13130,N_12705);
and U15755 (N_15755,N_12058,N_13168);
nor U15756 (N_15756,N_13984,N_13843);
nand U15757 (N_15757,N_13691,N_12638);
nor U15758 (N_15758,N_12292,N_13472);
and U15759 (N_15759,N_12072,N_13725);
nand U15760 (N_15760,N_12767,N_13090);
nor U15761 (N_15761,N_13076,N_13682);
nand U15762 (N_15762,N_12485,N_12944);
nand U15763 (N_15763,N_12855,N_12783);
and U15764 (N_15764,N_12782,N_13242);
and U15765 (N_15765,N_12615,N_13449);
nor U15766 (N_15766,N_12904,N_12319);
and U15767 (N_15767,N_13135,N_12464);
nor U15768 (N_15768,N_12815,N_13313);
and U15769 (N_15769,N_12959,N_12661);
xnor U15770 (N_15770,N_13037,N_13658);
or U15771 (N_15771,N_13729,N_13495);
or U15772 (N_15772,N_13963,N_12941);
or U15773 (N_15773,N_13334,N_13223);
nand U15774 (N_15774,N_12257,N_12573);
nand U15775 (N_15775,N_12088,N_12470);
nand U15776 (N_15776,N_12533,N_13008);
xnor U15777 (N_15777,N_13552,N_13219);
nand U15778 (N_15778,N_13684,N_13489);
or U15779 (N_15779,N_13303,N_12436);
xnor U15780 (N_15780,N_12460,N_13107);
or U15781 (N_15781,N_13662,N_12296);
nand U15782 (N_15782,N_12111,N_12451);
or U15783 (N_15783,N_13837,N_13553);
or U15784 (N_15784,N_12425,N_12464);
or U15785 (N_15785,N_13664,N_13865);
xor U15786 (N_15786,N_12032,N_13823);
or U15787 (N_15787,N_12555,N_12384);
xnor U15788 (N_15788,N_13073,N_13015);
nand U15789 (N_15789,N_13620,N_12867);
nor U15790 (N_15790,N_13656,N_13060);
nor U15791 (N_15791,N_13705,N_13932);
and U15792 (N_15792,N_12919,N_13051);
or U15793 (N_15793,N_12925,N_12104);
nor U15794 (N_15794,N_13730,N_13493);
nor U15795 (N_15795,N_12751,N_12618);
nand U15796 (N_15796,N_12548,N_12969);
nor U15797 (N_15797,N_13964,N_13564);
nor U15798 (N_15798,N_12598,N_12531);
and U15799 (N_15799,N_13632,N_13918);
xnor U15800 (N_15800,N_13271,N_13477);
xor U15801 (N_15801,N_12829,N_12318);
and U15802 (N_15802,N_13562,N_12405);
or U15803 (N_15803,N_13300,N_13710);
xnor U15804 (N_15804,N_12388,N_12113);
and U15805 (N_15805,N_13492,N_13959);
nand U15806 (N_15806,N_12027,N_13105);
nor U15807 (N_15807,N_13778,N_12381);
nor U15808 (N_15808,N_12320,N_12478);
nor U15809 (N_15809,N_13604,N_13192);
nor U15810 (N_15810,N_13642,N_12602);
nand U15811 (N_15811,N_13121,N_13688);
xnor U15812 (N_15812,N_13548,N_13310);
nand U15813 (N_15813,N_13053,N_13277);
nand U15814 (N_15814,N_13609,N_13298);
nor U15815 (N_15815,N_12284,N_12063);
nand U15816 (N_15816,N_12331,N_13109);
nor U15817 (N_15817,N_13125,N_13042);
nand U15818 (N_15818,N_13677,N_13561);
and U15819 (N_15819,N_13148,N_12967);
xnor U15820 (N_15820,N_13992,N_13614);
or U15821 (N_15821,N_12718,N_13962);
nand U15822 (N_15822,N_13312,N_13145);
nand U15823 (N_15823,N_12594,N_13865);
and U15824 (N_15824,N_12413,N_12857);
or U15825 (N_15825,N_12769,N_12276);
xnor U15826 (N_15826,N_13041,N_12470);
or U15827 (N_15827,N_13307,N_13320);
or U15828 (N_15828,N_13629,N_13497);
nor U15829 (N_15829,N_13918,N_13098);
nand U15830 (N_15830,N_12120,N_13465);
nor U15831 (N_15831,N_13541,N_12281);
nand U15832 (N_15832,N_13587,N_12548);
and U15833 (N_15833,N_12750,N_13603);
nand U15834 (N_15834,N_12792,N_12061);
nand U15835 (N_15835,N_13581,N_13820);
or U15836 (N_15836,N_12316,N_12948);
nor U15837 (N_15837,N_12680,N_12810);
and U15838 (N_15838,N_12385,N_12792);
nor U15839 (N_15839,N_13654,N_13902);
xnor U15840 (N_15840,N_12004,N_12109);
or U15841 (N_15841,N_13269,N_12062);
xor U15842 (N_15842,N_12817,N_12070);
nor U15843 (N_15843,N_12754,N_12530);
or U15844 (N_15844,N_12577,N_12472);
and U15845 (N_15845,N_12566,N_12774);
and U15846 (N_15846,N_13885,N_13808);
nor U15847 (N_15847,N_13269,N_13207);
xnor U15848 (N_15848,N_13554,N_13406);
and U15849 (N_15849,N_13394,N_13599);
xor U15850 (N_15850,N_12927,N_13891);
or U15851 (N_15851,N_13269,N_13971);
nand U15852 (N_15852,N_12255,N_13629);
or U15853 (N_15853,N_13115,N_13654);
nand U15854 (N_15854,N_12808,N_12479);
nand U15855 (N_15855,N_12139,N_13166);
nand U15856 (N_15856,N_12996,N_12480);
xor U15857 (N_15857,N_12752,N_12039);
or U15858 (N_15858,N_12055,N_12634);
or U15859 (N_15859,N_12212,N_12972);
or U15860 (N_15860,N_12119,N_13040);
and U15861 (N_15861,N_13107,N_12612);
nor U15862 (N_15862,N_13014,N_12073);
or U15863 (N_15863,N_12351,N_13457);
xor U15864 (N_15864,N_12576,N_13967);
xnor U15865 (N_15865,N_12536,N_12808);
xnor U15866 (N_15866,N_12149,N_13082);
nor U15867 (N_15867,N_13659,N_13396);
nor U15868 (N_15868,N_13532,N_12964);
xor U15869 (N_15869,N_12495,N_13986);
nand U15870 (N_15870,N_13247,N_13894);
and U15871 (N_15871,N_12140,N_12772);
nand U15872 (N_15872,N_13137,N_12056);
and U15873 (N_15873,N_12023,N_12106);
and U15874 (N_15874,N_12671,N_13999);
nand U15875 (N_15875,N_12905,N_12272);
nor U15876 (N_15876,N_13121,N_13333);
nand U15877 (N_15877,N_12276,N_13667);
xnor U15878 (N_15878,N_12988,N_12745);
nor U15879 (N_15879,N_13569,N_12839);
nand U15880 (N_15880,N_13053,N_13535);
nand U15881 (N_15881,N_12965,N_13190);
nand U15882 (N_15882,N_12075,N_13615);
nor U15883 (N_15883,N_12662,N_12369);
and U15884 (N_15884,N_13745,N_12992);
and U15885 (N_15885,N_13524,N_12188);
nor U15886 (N_15886,N_13533,N_13791);
xor U15887 (N_15887,N_12022,N_13243);
nand U15888 (N_15888,N_13538,N_12634);
and U15889 (N_15889,N_13061,N_12572);
nand U15890 (N_15890,N_13048,N_12348);
and U15891 (N_15891,N_12586,N_12192);
nor U15892 (N_15892,N_12701,N_13564);
and U15893 (N_15893,N_12473,N_13378);
xor U15894 (N_15894,N_13298,N_12637);
xnor U15895 (N_15895,N_13674,N_13673);
or U15896 (N_15896,N_12240,N_13783);
or U15897 (N_15897,N_13967,N_12256);
xnor U15898 (N_15898,N_12924,N_13405);
xor U15899 (N_15899,N_12590,N_12057);
and U15900 (N_15900,N_12849,N_12194);
nor U15901 (N_15901,N_12130,N_13852);
nand U15902 (N_15902,N_13783,N_13890);
or U15903 (N_15903,N_13586,N_12648);
and U15904 (N_15904,N_13946,N_12613);
xor U15905 (N_15905,N_13323,N_12872);
xor U15906 (N_15906,N_13153,N_12640);
and U15907 (N_15907,N_12256,N_13243);
and U15908 (N_15908,N_12745,N_13623);
or U15909 (N_15909,N_12358,N_13942);
and U15910 (N_15910,N_13768,N_12395);
nand U15911 (N_15911,N_12080,N_13282);
or U15912 (N_15912,N_12324,N_13029);
and U15913 (N_15913,N_12635,N_13884);
nand U15914 (N_15914,N_12012,N_12932);
or U15915 (N_15915,N_12283,N_12479);
nor U15916 (N_15916,N_13050,N_13676);
nand U15917 (N_15917,N_12236,N_13895);
and U15918 (N_15918,N_13762,N_12915);
or U15919 (N_15919,N_12858,N_12327);
nand U15920 (N_15920,N_13123,N_13596);
xor U15921 (N_15921,N_13184,N_13284);
nor U15922 (N_15922,N_13478,N_12442);
or U15923 (N_15923,N_13467,N_13042);
xnor U15924 (N_15924,N_12622,N_12201);
and U15925 (N_15925,N_12868,N_12398);
or U15926 (N_15926,N_12265,N_13630);
nand U15927 (N_15927,N_13088,N_12753);
nor U15928 (N_15928,N_13597,N_13824);
and U15929 (N_15929,N_13619,N_12120);
nand U15930 (N_15930,N_13037,N_12792);
and U15931 (N_15931,N_12645,N_13736);
nor U15932 (N_15932,N_13905,N_12907);
xor U15933 (N_15933,N_12900,N_13214);
or U15934 (N_15934,N_13400,N_12521);
nand U15935 (N_15935,N_13914,N_12697);
nand U15936 (N_15936,N_13022,N_12484);
xnor U15937 (N_15937,N_12050,N_13560);
and U15938 (N_15938,N_13469,N_13200);
and U15939 (N_15939,N_13687,N_13457);
nor U15940 (N_15940,N_13362,N_13735);
nand U15941 (N_15941,N_13850,N_12275);
nor U15942 (N_15942,N_12285,N_12101);
xnor U15943 (N_15943,N_12515,N_12173);
nor U15944 (N_15944,N_13811,N_13907);
nor U15945 (N_15945,N_13248,N_13137);
or U15946 (N_15946,N_12605,N_12086);
nor U15947 (N_15947,N_12106,N_12984);
or U15948 (N_15948,N_12208,N_13121);
or U15949 (N_15949,N_12652,N_12628);
nand U15950 (N_15950,N_13104,N_12180);
or U15951 (N_15951,N_13708,N_13381);
nor U15952 (N_15952,N_12860,N_12788);
nor U15953 (N_15953,N_12527,N_12276);
or U15954 (N_15954,N_12253,N_13987);
and U15955 (N_15955,N_13657,N_12169);
or U15956 (N_15956,N_12923,N_12552);
or U15957 (N_15957,N_12448,N_13367);
nor U15958 (N_15958,N_13133,N_13519);
nor U15959 (N_15959,N_12818,N_12516);
nor U15960 (N_15960,N_12110,N_13847);
xnor U15961 (N_15961,N_13225,N_13073);
and U15962 (N_15962,N_12492,N_12330);
or U15963 (N_15963,N_13001,N_13425);
or U15964 (N_15964,N_13294,N_12099);
xor U15965 (N_15965,N_13912,N_13066);
nand U15966 (N_15966,N_13594,N_13944);
nand U15967 (N_15967,N_12022,N_12768);
and U15968 (N_15968,N_13697,N_12411);
nand U15969 (N_15969,N_12002,N_13091);
xnor U15970 (N_15970,N_13822,N_12747);
nor U15971 (N_15971,N_12396,N_12465);
nand U15972 (N_15972,N_12522,N_13034);
nor U15973 (N_15973,N_13921,N_12054);
or U15974 (N_15974,N_13716,N_13918);
or U15975 (N_15975,N_12053,N_13883);
nand U15976 (N_15976,N_13299,N_12760);
nor U15977 (N_15977,N_13858,N_13244);
and U15978 (N_15978,N_12347,N_12924);
and U15979 (N_15979,N_12627,N_13989);
xnor U15980 (N_15980,N_13503,N_13571);
nand U15981 (N_15981,N_12072,N_12477);
nor U15982 (N_15982,N_13290,N_12429);
and U15983 (N_15983,N_12578,N_12705);
or U15984 (N_15984,N_13101,N_12017);
nand U15985 (N_15985,N_13199,N_13855);
nor U15986 (N_15986,N_13629,N_12033);
and U15987 (N_15987,N_13431,N_12881);
or U15988 (N_15988,N_13354,N_12353);
nand U15989 (N_15989,N_12738,N_13144);
nor U15990 (N_15990,N_12083,N_12207);
nand U15991 (N_15991,N_12078,N_13130);
and U15992 (N_15992,N_13470,N_13821);
and U15993 (N_15993,N_12387,N_12577);
and U15994 (N_15994,N_13164,N_13511);
nor U15995 (N_15995,N_12478,N_13211);
nand U15996 (N_15996,N_13823,N_13648);
or U15997 (N_15997,N_12397,N_13447);
xor U15998 (N_15998,N_12973,N_12427);
and U15999 (N_15999,N_12809,N_13251);
and U16000 (N_16000,N_15842,N_14835);
xnor U16001 (N_16001,N_15482,N_15269);
nor U16002 (N_16002,N_15179,N_14176);
or U16003 (N_16003,N_14230,N_15418);
nand U16004 (N_16004,N_14483,N_15350);
and U16005 (N_16005,N_14903,N_14722);
nand U16006 (N_16006,N_14984,N_15756);
nor U16007 (N_16007,N_15515,N_14885);
nand U16008 (N_16008,N_15557,N_14647);
and U16009 (N_16009,N_14394,N_15845);
xnor U16010 (N_16010,N_14619,N_15433);
and U16011 (N_16011,N_15621,N_15454);
or U16012 (N_16012,N_15365,N_14865);
or U16013 (N_16013,N_15170,N_14950);
nor U16014 (N_16014,N_14448,N_15381);
xnor U16015 (N_16015,N_15695,N_14734);
nor U16016 (N_16016,N_14987,N_15735);
or U16017 (N_16017,N_15834,N_14714);
and U16018 (N_16018,N_14046,N_15382);
and U16019 (N_16019,N_14508,N_14995);
xnor U16020 (N_16020,N_14609,N_15214);
nor U16021 (N_16021,N_15188,N_14257);
nand U16022 (N_16022,N_14260,N_14998);
and U16023 (N_16023,N_15945,N_14075);
and U16024 (N_16024,N_14087,N_14828);
and U16025 (N_16025,N_14419,N_14705);
xnor U16026 (N_16026,N_14313,N_15058);
xor U16027 (N_16027,N_14564,N_15244);
xnor U16028 (N_16028,N_15473,N_15994);
and U16029 (N_16029,N_14654,N_14220);
or U16030 (N_16030,N_15070,N_14738);
nor U16031 (N_16031,N_15161,N_15000);
nor U16032 (N_16032,N_14655,N_14287);
nor U16033 (N_16033,N_14898,N_15658);
nand U16034 (N_16034,N_14510,N_15563);
xnor U16035 (N_16035,N_14862,N_15646);
nand U16036 (N_16036,N_14121,N_14604);
nand U16037 (N_16037,N_15668,N_14053);
nand U16038 (N_16038,N_15762,N_14871);
and U16039 (N_16039,N_15728,N_15539);
or U16040 (N_16040,N_15523,N_15870);
nand U16041 (N_16041,N_14954,N_14746);
or U16042 (N_16042,N_15556,N_14852);
nor U16043 (N_16043,N_14826,N_14966);
or U16044 (N_16044,N_15797,N_14308);
xor U16045 (N_16045,N_14331,N_15786);
nand U16046 (N_16046,N_15326,N_14918);
nand U16047 (N_16047,N_15319,N_14468);
xor U16048 (N_16048,N_14110,N_15738);
or U16049 (N_16049,N_15043,N_14690);
nor U16050 (N_16050,N_14893,N_15575);
xnor U16051 (N_16051,N_15030,N_15437);
xnor U16052 (N_16052,N_15074,N_15112);
and U16053 (N_16053,N_14507,N_15248);
or U16054 (N_16054,N_14820,N_15935);
or U16055 (N_16055,N_14550,N_14159);
nand U16056 (N_16056,N_15195,N_15477);
or U16057 (N_16057,N_15184,N_15475);
and U16058 (N_16058,N_15865,N_14493);
nand U16059 (N_16059,N_15354,N_14902);
nor U16060 (N_16060,N_15443,N_14977);
and U16061 (N_16061,N_14624,N_14250);
xor U16062 (N_16062,N_14014,N_15297);
nor U16063 (N_16063,N_14881,N_14780);
nand U16064 (N_16064,N_14704,N_14588);
nand U16065 (N_16065,N_14059,N_15198);
or U16066 (N_16066,N_14910,N_15608);
nand U16067 (N_16067,N_14109,N_15399);
nor U16068 (N_16068,N_14436,N_14727);
and U16069 (N_16069,N_15794,N_15014);
nand U16070 (N_16070,N_15837,N_15872);
or U16071 (N_16071,N_15597,N_14457);
nand U16072 (N_16072,N_15929,N_15614);
or U16073 (N_16073,N_15034,N_15961);
nor U16074 (N_16074,N_15628,N_15122);
nor U16075 (N_16075,N_14720,N_15124);
or U16076 (N_16076,N_14120,N_15585);
nor U16077 (N_16077,N_15751,N_14529);
or U16078 (N_16078,N_14427,N_15873);
nor U16079 (N_16079,N_15877,N_14043);
nor U16080 (N_16080,N_15129,N_15252);
or U16081 (N_16081,N_15208,N_14854);
xor U16082 (N_16082,N_14165,N_15850);
or U16083 (N_16083,N_15143,N_14806);
nand U16084 (N_16084,N_14606,N_14586);
xnor U16085 (N_16085,N_15888,N_15978);
and U16086 (N_16086,N_15398,N_14324);
and U16087 (N_16087,N_15111,N_14982);
or U16088 (N_16088,N_15601,N_14599);
nor U16089 (N_16089,N_14334,N_14636);
xor U16090 (N_16090,N_15419,N_15220);
or U16091 (N_16091,N_14482,N_14288);
or U16092 (N_16092,N_14719,N_15932);
or U16093 (N_16093,N_14639,N_15446);
nor U16094 (N_16094,N_15590,N_15465);
or U16095 (N_16095,N_15414,N_15469);
nor U16096 (N_16096,N_15555,N_15603);
xnor U16097 (N_16097,N_15548,N_14924);
xor U16098 (N_16098,N_15145,N_15496);
xnor U16099 (N_16099,N_14499,N_15956);
nand U16100 (N_16100,N_14375,N_15960);
nor U16101 (N_16101,N_14201,N_14996);
nand U16102 (N_16102,N_14280,N_14878);
nor U16103 (N_16103,N_15595,N_15880);
and U16104 (N_16104,N_15106,N_15624);
nand U16105 (N_16105,N_15222,N_15085);
and U16106 (N_16106,N_15807,N_15329);
xor U16107 (N_16107,N_14859,N_14861);
and U16108 (N_16108,N_14026,N_15080);
xnor U16109 (N_16109,N_14699,N_15981);
nor U16110 (N_16110,N_15627,N_15051);
nor U16111 (N_16111,N_14019,N_14356);
nor U16112 (N_16112,N_14414,N_15013);
and U16113 (N_16113,N_14739,N_15023);
nor U16114 (N_16114,N_15938,N_14904);
nand U16115 (N_16115,N_15755,N_14556);
xor U16116 (N_16116,N_15242,N_15980);
nor U16117 (N_16117,N_14565,N_15238);
or U16118 (N_16118,N_15001,N_15654);
nand U16119 (N_16119,N_15830,N_14174);
xor U16120 (N_16120,N_14882,N_15202);
and U16121 (N_16121,N_14845,N_14147);
or U16122 (N_16122,N_14923,N_14429);
nor U16123 (N_16123,N_14064,N_14160);
and U16124 (N_16124,N_14782,N_15749);
nor U16125 (N_16125,N_15921,N_15788);
or U16126 (N_16126,N_14481,N_14976);
and U16127 (N_16127,N_14042,N_15089);
and U16128 (N_16128,N_14842,N_15512);
xnor U16129 (N_16129,N_14567,N_14101);
xor U16130 (N_16130,N_15985,N_14563);
or U16131 (N_16131,N_15653,N_14351);
or U16132 (N_16132,N_15869,N_14285);
nor U16133 (N_16133,N_15953,N_14616);
xnor U16134 (N_16134,N_14920,N_14623);
xnor U16135 (N_16135,N_14143,N_15160);
xnor U16136 (N_16136,N_14873,N_14384);
nor U16137 (N_16137,N_14184,N_14768);
nand U16138 (N_16138,N_14681,N_15906);
nand U16139 (N_16139,N_15918,N_15661);
or U16140 (N_16140,N_14315,N_14416);
nor U16141 (N_16141,N_15146,N_15140);
nand U16142 (N_16142,N_14518,N_15974);
or U16143 (N_16143,N_14151,N_15169);
and U16144 (N_16144,N_15271,N_14540);
or U16145 (N_16145,N_14115,N_15931);
nand U16146 (N_16146,N_14761,N_14600);
and U16147 (N_16147,N_14291,N_14975);
and U16148 (N_16148,N_14008,N_15341);
nand U16149 (N_16149,N_14072,N_15311);
nand U16150 (N_16150,N_15284,N_14018);
nor U16151 (N_16151,N_15853,N_14863);
xnor U16152 (N_16152,N_15348,N_14325);
or U16153 (N_16153,N_14669,N_14829);
xnor U16154 (N_16154,N_15858,N_14047);
and U16155 (N_16155,N_15340,N_15229);
or U16156 (N_16156,N_14361,N_15417);
nor U16157 (N_16157,N_15404,N_14497);
and U16158 (N_16158,N_14853,N_15474);
or U16159 (N_16159,N_15721,N_14404);
or U16160 (N_16160,N_14601,N_15724);
or U16161 (N_16161,N_15024,N_14985);
nand U16162 (N_16162,N_15879,N_15237);
nor U16163 (N_16163,N_15042,N_15403);
or U16164 (N_16164,N_15141,N_15412);
xnor U16165 (N_16165,N_15163,N_14067);
nor U16166 (N_16166,N_15538,N_15650);
xnor U16167 (N_16167,N_14970,N_15854);
and U16168 (N_16168,N_15368,N_14353);
nand U16169 (N_16169,N_14298,N_14818);
nor U16170 (N_16170,N_15312,N_14801);
xor U16171 (N_16171,N_14908,N_14846);
or U16172 (N_16172,N_15483,N_14848);
nor U16173 (N_16173,N_15409,N_14010);
xnor U16174 (N_16174,N_14281,N_15103);
xor U16175 (N_16175,N_15460,N_14225);
and U16176 (N_16176,N_15611,N_15272);
nor U16177 (N_16177,N_15395,N_14799);
and U16178 (N_16178,N_15839,N_15690);
and U16179 (N_16179,N_14748,N_15200);
or U16180 (N_16180,N_15820,N_15691);
nand U16181 (N_16181,N_15207,N_14857);
nand U16182 (N_16182,N_14232,N_15002);
nor U16183 (N_16183,N_15549,N_14352);
and U16184 (N_16184,N_15359,N_14038);
and U16185 (N_16185,N_15498,N_14033);
nor U16186 (N_16186,N_15586,N_15753);
or U16187 (N_16187,N_14822,N_14055);
nand U16188 (N_16188,N_14126,N_15525);
or U16189 (N_16189,N_14226,N_15508);
xnor U16190 (N_16190,N_14104,N_15031);
or U16191 (N_16191,N_15126,N_15670);
xor U16192 (N_16192,N_15317,N_15645);
nand U16193 (N_16193,N_14093,N_14082);
xnor U16194 (N_16194,N_14145,N_15565);
xnor U16195 (N_16195,N_15809,N_14716);
nor U16196 (N_16196,N_14181,N_14349);
xor U16197 (N_16197,N_14166,N_15912);
nor U16198 (N_16198,N_14643,N_15532);
nor U16199 (N_16199,N_15424,N_15388);
xor U16200 (N_16200,N_14050,N_15727);
and U16201 (N_16201,N_15743,N_15702);
or U16202 (N_16202,N_14138,N_14136);
nor U16203 (N_16203,N_14237,N_14744);
and U16204 (N_16204,N_14022,N_15147);
xor U16205 (N_16205,N_15971,N_15968);
and U16206 (N_16206,N_15801,N_14900);
nor U16207 (N_16207,N_15770,N_15197);
nor U16208 (N_16208,N_15710,N_14407);
and U16209 (N_16209,N_15719,N_15101);
or U16210 (N_16210,N_15400,N_14498);
and U16211 (N_16211,N_14304,N_15159);
nor U16212 (N_16212,N_15174,N_15617);
or U16213 (N_16213,N_14422,N_14812);
or U16214 (N_16214,N_15493,N_14466);
nand U16215 (N_16215,N_15249,N_15201);
or U16216 (N_16216,N_14322,N_15576);
and U16217 (N_16217,N_14317,N_14687);
and U16218 (N_16218,N_14139,N_14559);
and U16219 (N_16219,N_15785,N_15666);
or U16220 (N_16220,N_15472,N_15886);
nand U16221 (N_16221,N_15600,N_15268);
nand U16222 (N_16222,N_14929,N_14302);
xnor U16223 (N_16223,N_15619,N_15745);
nor U16224 (N_16224,N_14376,N_15782);
and U16225 (N_16225,N_15803,N_14763);
and U16226 (N_16226,N_15635,N_15922);
or U16227 (N_16227,N_15102,N_14301);
or U16228 (N_16228,N_15307,N_15892);
xnor U16229 (N_16229,N_14073,N_15992);
and U16230 (N_16230,N_14449,N_14032);
or U16231 (N_16231,N_15573,N_14048);
or U16232 (N_16232,N_14027,N_14157);
nor U16233 (N_16233,N_15954,N_14651);
nand U16234 (N_16234,N_15266,N_15276);
nand U16235 (N_16235,N_15442,N_15587);
nor U16236 (N_16236,N_15527,N_15541);
and U16237 (N_16237,N_14386,N_15881);
xnor U16238 (N_16238,N_15584,N_14735);
xor U16239 (N_16239,N_15625,N_15006);
and U16240 (N_16240,N_15822,N_15187);
xor U16241 (N_16241,N_14702,N_14413);
nand U16242 (N_16242,N_15314,N_14063);
nand U16243 (N_16243,N_15115,N_15393);
nor U16244 (N_16244,N_14580,N_14937);
nor U16245 (N_16245,N_15049,N_14876);
or U16246 (N_16246,N_14869,N_14547);
or U16247 (N_16247,N_14723,N_14103);
or U16248 (N_16248,N_14752,N_14330);
or U16249 (N_16249,N_15748,N_15947);
nand U16250 (N_16250,N_15923,N_15718);
xnor U16251 (N_16251,N_15376,N_15659);
or U16252 (N_16252,N_15939,N_15480);
nand U16253 (N_16253,N_14113,N_14633);
nor U16254 (N_16254,N_15279,N_15866);
xor U16255 (N_16255,N_15760,N_14798);
nand U16256 (N_16256,N_14554,N_15704);
or U16257 (N_16257,N_14221,N_15694);
or U16258 (N_16258,N_14303,N_15946);
nor U16259 (N_16259,N_14571,N_15522);
nor U16260 (N_16260,N_14941,N_14896);
xor U16261 (N_16261,N_15852,N_15097);
or U16262 (N_16262,N_15335,N_15581);
and U16263 (N_16263,N_15909,N_14395);
xnor U16264 (N_16264,N_15720,N_14380);
and U16265 (N_16265,N_14986,N_15543);
nand U16266 (N_16266,N_14775,N_14057);
or U16267 (N_16267,N_15206,N_15204);
and U16268 (N_16268,N_15009,N_15151);
nand U16269 (N_16269,N_15840,N_14792);
nand U16270 (N_16270,N_15976,N_15062);
nand U16271 (N_16271,N_15210,N_15677);
and U16272 (N_16272,N_14204,N_15732);
nand U16273 (N_16273,N_15233,N_14691);
nor U16274 (N_16274,N_14328,N_15185);
nor U16275 (N_16275,N_14167,N_14688);
xnor U16276 (N_16276,N_14194,N_15746);
or U16277 (N_16277,N_14480,N_14238);
and U16278 (N_16278,N_14530,N_15007);
xnor U16279 (N_16279,N_14455,N_14939);
xor U16280 (N_16280,N_14321,N_14843);
nor U16281 (N_16281,N_14659,N_14953);
xnor U16282 (N_16282,N_14294,N_14860);
and U16283 (N_16283,N_15505,N_15158);
or U16284 (N_16284,N_15019,N_14839);
and U16285 (N_16285,N_14085,N_14132);
nand U16286 (N_16286,N_15485,N_15041);
or U16287 (N_16287,N_14195,N_15025);
or U16288 (N_16288,N_15243,N_15674);
and U16289 (N_16289,N_14625,N_15387);
or U16290 (N_16290,N_15048,N_14730);
nand U16291 (N_16291,N_15965,N_15090);
xor U16292 (N_16292,N_15882,N_15864);
xor U16293 (N_16293,N_15351,N_14615);
nand U16294 (N_16294,N_15177,N_14146);
xor U16295 (N_16295,N_14389,N_15529);
nand U16296 (N_16296,N_14751,N_14090);
xnor U16297 (N_16297,N_14830,N_14310);
nand U16298 (N_16298,N_14742,N_15737);
nor U16299 (N_16299,N_14097,N_15245);
or U16300 (N_16300,N_15826,N_14819);
and U16301 (N_16301,N_14094,N_14533);
nor U16302 (N_16302,N_15339,N_14519);
xor U16303 (N_16303,N_14005,N_14016);
and U16304 (N_16304,N_14337,N_14737);
or U16305 (N_16305,N_15664,N_14524);
nor U16306 (N_16306,N_14474,N_15936);
nand U16307 (N_16307,N_14229,N_14522);
and U16308 (N_16308,N_15180,N_14177);
and U16309 (N_16309,N_15959,N_15503);
nor U16310 (N_16310,N_15526,N_14827);
xnor U16311 (N_16311,N_15638,N_14892);
nor U16312 (N_16312,N_14894,N_14442);
nor U16313 (N_16313,N_15769,N_15069);
or U16314 (N_16314,N_15355,N_14015);
nor U16315 (N_16315,N_15752,N_15490);
or U16316 (N_16316,N_14668,N_14078);
and U16317 (N_16317,N_14037,N_15712);
nor U16318 (N_16318,N_14759,N_14172);
and U16319 (N_16319,N_14595,N_14333);
xnor U16320 (N_16320,N_14765,N_15800);
and U16321 (N_16321,N_14607,N_15277);
and U16322 (N_16322,N_14127,N_14756);
xnor U16323 (N_16323,N_15799,N_14758);
xnor U16324 (N_16324,N_14076,N_15846);
and U16325 (N_16325,N_15459,N_15157);
or U16326 (N_16326,N_15464,N_14437);
nor U16327 (N_16327,N_14058,N_14909);
nor U16328 (N_16328,N_15436,N_15036);
and U16329 (N_16329,N_15819,N_14783);
nor U16330 (N_16330,N_14329,N_14771);
nand U16331 (N_16331,N_14593,N_15022);
and U16332 (N_16332,N_14135,N_14823);
xnor U16333 (N_16333,N_14709,N_15969);
and U16334 (N_16334,N_15633,N_14747);
xnor U16335 (N_16335,N_14079,N_15410);
nand U16336 (N_16336,N_15836,N_14045);
and U16337 (N_16337,N_15796,N_14289);
xor U16338 (N_16338,N_14447,N_14585);
or U16339 (N_16339,N_14628,N_15521);
nand U16340 (N_16340,N_15885,N_14488);
and U16341 (N_16341,N_14091,N_15793);
nor U16342 (N_16342,N_14239,N_15430);
nand U16343 (N_16343,N_15189,N_15520);
nand U16344 (N_16344,N_15037,N_14469);
nor U16345 (N_16345,N_14300,N_14698);
nand U16346 (N_16346,N_14980,N_15518);
nand U16347 (N_16347,N_14411,N_14342);
nand U16348 (N_16348,N_15767,N_15280);
xor U16349 (N_16349,N_14895,N_14989);
nor U16350 (N_16350,N_15270,N_15697);
or U16351 (N_16351,N_15369,N_15154);
and U16352 (N_16352,N_14368,N_14247);
nand U16353 (N_16353,N_15703,N_15121);
xnor U16354 (N_16354,N_15110,N_15173);
nor U16355 (N_16355,N_14156,N_14102);
nand U16356 (N_16356,N_14189,N_14506);
nor U16357 (N_16357,N_14131,N_15342);
nor U16358 (N_16358,N_14212,N_14140);
nor U16359 (N_16359,N_15681,N_14921);
nor U16360 (N_16360,N_14244,N_14007);
or U16361 (N_16361,N_14856,N_14814);
xor U16362 (N_16362,N_14453,N_15364);
nand U16363 (N_16363,N_14080,N_14657);
xnor U16364 (N_16364,N_14800,N_14545);
or U16365 (N_16365,N_15715,N_14362);
nand U16366 (N_16366,N_14789,N_15620);
and U16367 (N_16367,N_14978,N_14745);
nor U16368 (N_16368,N_15594,N_15773);
nand U16369 (N_16369,N_14435,N_14273);
xnor U16370 (N_16370,N_15811,N_15156);
or U16371 (N_16371,N_15315,N_14790);
xor U16372 (N_16372,N_14052,N_15942);
nor U16373 (N_16373,N_14809,N_15373);
nand U16374 (N_16374,N_14295,N_14666);
nand U16375 (N_16375,N_15570,N_14383);
nand U16376 (N_16376,N_15887,N_15634);
xnor U16377 (N_16377,N_14182,N_15005);
nor U16378 (N_16378,N_15894,N_15116);
and U16379 (N_16379,N_14387,N_14670);
nand U16380 (N_16380,N_14781,N_14439);
or U16381 (N_16381,N_15630,N_14088);
and U16382 (N_16382,N_14576,N_14675);
or U16383 (N_16383,N_14877,N_14797);
and U16384 (N_16384,N_14426,N_14256);
xor U16385 (N_16385,N_14946,N_15344);
nor U16386 (N_16386,N_15391,N_15679);
nor U16387 (N_16387,N_14804,N_14880);
or U16388 (N_16388,N_15780,N_14926);
nand U16389 (N_16389,N_15120,N_15662);
or U16390 (N_16390,N_14749,N_15078);
xnor U16391 (N_16391,N_15907,N_15723);
xnor U16392 (N_16392,N_14111,N_14107);
nor U16393 (N_16393,N_14645,N_15343);
nand U16394 (N_16394,N_15441,N_15567);
or U16395 (N_16395,N_15528,N_14441);
or U16396 (N_16396,N_15699,N_15913);
xnor U16397 (N_16397,N_15682,N_14712);
or U16398 (N_16398,N_14679,N_15313);
nand U16399 (N_16399,N_14660,N_14613);
xor U16400 (N_16400,N_14897,N_15902);
and U16401 (N_16401,N_15602,N_14150);
and U16402 (N_16402,N_14796,N_15813);
or U16403 (N_16403,N_14803,N_15384);
xnor U16404 (N_16404,N_15133,N_15861);
or U16405 (N_16405,N_14963,N_15775);
nor U16406 (N_16406,N_14543,N_14392);
and U16407 (N_16407,N_14382,N_14390);
or U16408 (N_16408,N_14805,N_14013);
or U16409 (N_16409,N_15814,N_15591);
nor U16410 (N_16410,N_14959,N_14456);
and U16411 (N_16411,N_15226,N_15053);
nand U16412 (N_16412,N_14786,N_14183);
or U16413 (N_16413,N_15429,N_15792);
or U16414 (N_16414,N_15499,N_15998);
and U16415 (N_16415,N_14477,N_14602);
or U16416 (N_16416,N_14290,N_14444);
xnor U16417 (N_16417,N_15278,N_14913);
and U16418 (N_16418,N_14663,N_15017);
nor U16419 (N_16419,N_15516,N_15450);
or U16420 (N_16420,N_15401,N_15919);
nor U16421 (N_16421,N_14401,N_15302);
nand U16422 (N_16422,N_14965,N_14408);
and U16423 (N_16423,N_14542,N_15930);
nand U16424 (N_16424,N_14557,N_15517);
nand U16425 (N_16425,N_14454,N_15578);
xor U16426 (N_16426,N_14207,N_15943);
and U16427 (N_16427,N_14808,N_15808);
nor U16428 (N_16428,N_15725,N_14489);
nand U16429 (N_16429,N_14462,N_14598);
and U16430 (N_16430,N_14574,N_14040);
xor U16431 (N_16431,N_15878,N_14658);
xnor U16432 (N_16432,N_14590,N_14750);
and U16433 (N_16433,N_14592,N_14359);
xnor U16434 (N_16434,N_15232,N_15261);
xnor U16435 (N_16435,N_14060,N_15554);
nand U16436 (N_16436,N_15741,N_15378);
xor U16437 (N_16437,N_15993,N_15445);
and U16438 (N_16438,N_14731,N_14286);
and U16439 (N_16439,N_14224,N_15068);
and U16440 (N_16440,N_14114,N_14089);
xnor U16441 (N_16441,N_14934,N_14695);
nand U16442 (N_16442,N_14193,N_14824);
nor U16443 (N_16443,N_15492,N_14077);
and U16444 (N_16444,N_14662,N_15291);
xor U16445 (N_16445,N_15899,N_14791);
nor U16446 (N_16446,N_14326,N_15322);
xor U16447 (N_16447,N_14400,N_15950);
xnor U16448 (N_16448,N_14555,N_15997);
nor U16449 (N_16449,N_15065,N_15531);
nor U16450 (N_16450,N_14350,N_15641);
xnor U16451 (N_16451,N_15263,N_14642);
and U16452 (N_16452,N_14638,N_15091);
and U16453 (N_16453,N_15763,N_15636);
nand U16454 (N_16454,N_15047,N_15431);
nor U16455 (N_16455,N_15833,N_15372);
and U16456 (N_16456,N_15076,N_14552);
nand U16457 (N_16457,N_14689,N_14673);
xnor U16458 (N_16458,N_14478,N_14402);
and U16459 (N_16459,N_15044,N_14944);
xor U16460 (N_16460,N_14268,N_15972);
xor U16461 (N_16461,N_15218,N_15606);
nor U16462 (N_16462,N_15910,N_15035);
or U16463 (N_16463,N_15008,N_15561);
xor U16464 (N_16464,N_14922,N_14766);
and U16465 (N_16465,N_15394,N_15651);
xor U16466 (N_16466,N_15108,N_15420);
or U16467 (N_16467,N_15687,N_15692);
nor U16468 (N_16468,N_15003,N_15228);
nor U16469 (N_16469,N_15254,N_15977);
xnor U16470 (N_16470,N_15332,N_15761);
or U16471 (N_16471,N_14128,N_15476);
nand U16472 (N_16472,N_14931,N_15716);
and U16473 (N_16473,N_14884,N_14569);
and U16474 (N_16474,N_15361,N_14795);
nor U16475 (N_16475,N_15347,N_15012);
nand U16476 (N_16476,N_14509,N_14274);
nand U16477 (N_16477,N_15027,N_14891);
xor U16478 (N_16478,N_15685,N_15273);
or U16479 (N_16479,N_15487,N_15693);
and U16480 (N_16480,N_14502,N_15572);
nor U16481 (N_16481,N_14205,N_14646);
xnor U16482 (N_16482,N_15300,N_14603);
or U16483 (N_16483,N_14208,N_15577);
nor U16484 (N_16484,N_14886,N_14347);
xnor U16485 (N_16485,N_15029,N_14117);
nor U16486 (N_16486,N_14011,N_14084);
nand U16487 (N_16487,N_15209,N_15453);
nand U16488 (N_16488,N_14335,N_14568);
xnor U16489 (N_16489,N_15324,N_14890);
and U16490 (N_16490,N_15544,N_14206);
nand U16491 (N_16491,N_14832,N_15260);
or U16492 (N_16492,N_15629,N_15655);
and U16493 (N_16493,N_15583,N_15489);
or U16494 (N_16494,N_14762,N_14279);
nand U16495 (N_16495,N_14632,N_15667);
nor U16496 (N_16496,N_15897,N_14610);
and U16497 (N_16497,N_14558,N_15908);
or U16498 (N_16498,N_15726,N_15711);
nand U16499 (N_16499,N_14171,N_14443);
nor U16500 (N_16500,N_15566,N_14770);
and U16501 (N_16501,N_15251,N_14676);
xor U16502 (N_16502,N_15730,N_14717);
or U16503 (N_16503,N_15867,N_14332);
and U16504 (N_16504,N_15432,N_14570);
nand U16505 (N_16505,N_14648,N_15967);
xnor U16506 (N_16506,N_14056,N_15914);
xnor U16507 (N_16507,N_15416,N_15569);
nand U16508 (N_16508,N_15675,N_14141);
xnor U16509 (N_16509,N_15148,N_15898);
nor U16510 (N_16510,N_14945,N_14041);
or U16511 (N_16511,N_14450,N_15966);
xnor U16512 (N_16512,N_15491,N_15904);
xnor U16513 (N_16513,N_14774,N_14405);
xor U16514 (N_16514,N_14988,N_15299);
xor U16515 (N_16515,N_14316,N_14733);
xor U16516 (N_16516,N_15379,N_14083);
xor U16517 (N_16517,N_15114,N_15996);
nand U16518 (N_16518,N_14071,N_14017);
xnor U16519 (N_16519,N_15298,N_15289);
and U16520 (N_16520,N_15783,N_15439);
xnor U16521 (N_16521,N_15766,N_14269);
nor U16522 (N_16522,N_15083,N_15831);
nor U16523 (N_16523,N_14144,N_14433);
and U16524 (N_16524,N_15933,N_15405);
and U16525 (N_16525,N_14787,N_14867);
xnor U16526 (N_16526,N_14283,N_14815);
nand U16527 (N_16527,N_14125,N_14485);
or U16528 (N_16528,N_15402,N_15806);
or U16529 (N_16529,N_14622,N_14451);
or U16530 (N_16530,N_14234,N_15310);
and U16531 (N_16531,N_14684,N_14035);
nand U16532 (N_16532,N_15125,N_15191);
nand U16533 (N_16533,N_14215,N_15764);
nand U16534 (N_16534,N_15057,N_14981);
and U16535 (N_16535,N_14706,N_15562);
nor U16536 (N_16536,N_15479,N_15318);
or U16537 (N_16537,N_15039,N_14844);
nand U16538 (N_16538,N_14729,N_15021);
nand U16539 (N_16539,N_15571,N_14341);
nor U16540 (N_16540,N_15596,N_15790);
or U16541 (N_16541,N_15952,N_14108);
and U16542 (N_16542,N_14412,N_15805);
nand U16543 (N_16543,N_15765,N_14887);
nor U16544 (N_16544,N_15497,N_14534);
xnor U16545 (N_16545,N_14385,N_14248);
and U16546 (N_16546,N_15895,N_14777);
nor U16547 (N_16547,N_15707,N_15413);
or U16548 (N_16548,N_15045,N_15138);
nand U16549 (N_16549,N_15234,N_14947);
nand U16550 (N_16550,N_14118,N_14112);
or U16551 (N_16551,N_14242,N_15925);
and U16552 (N_16552,N_15186,N_14682);
and U16553 (N_16553,N_15537,N_15287);
xor U16554 (N_16554,N_14767,N_15462);
nand U16555 (N_16555,N_14432,N_14068);
and U16556 (N_16556,N_14618,N_14925);
or U16557 (N_16557,N_15285,N_15099);
nand U16558 (N_16558,N_15709,N_15109);
nand U16559 (N_16559,N_14621,N_14521);
and U16560 (N_16560,N_14740,N_15920);
xnor U16561 (N_16561,N_15818,N_15274);
and U16562 (N_16562,N_14840,N_14993);
and U16563 (N_16563,N_14116,N_14784);
or U16564 (N_16564,N_14711,N_15337);
or U16565 (N_16565,N_15964,N_14938);
xor U16566 (N_16566,N_14958,N_14464);
xnor U16567 (N_16567,N_14907,N_14000);
nor U16568 (N_16568,N_15371,N_15192);
xor U16569 (N_16569,N_15194,N_15838);
nor U16570 (N_16570,N_15683,N_15731);
nand U16571 (N_16571,N_14270,N_15451);
or U16572 (N_16572,N_15408,N_14905);
xnor U16573 (N_16573,N_15863,N_15744);
xor U16574 (N_16574,N_14584,N_15357);
nor U16575 (N_16575,N_14227,N_14755);
xnor U16576 (N_16576,N_14410,N_15075);
or U16577 (N_16577,N_15631,N_15995);
xor U16578 (N_16578,N_14213,N_14346);
nor U16579 (N_16579,N_14252,N_14180);
nor U16580 (N_16580,N_15844,N_14323);
and U16581 (N_16581,N_15758,N_14974);
or U16582 (N_16582,N_14933,N_15467);
nor U16583 (N_16583,N_14741,N_14381);
xor U16584 (N_16584,N_15536,N_14211);
nand U16585 (N_16585,N_15828,N_15618);
or U16586 (N_16586,N_15092,N_15081);
or U16587 (N_16587,N_14841,N_14369);
xor U16588 (N_16588,N_14906,N_14501);
or U16589 (N_16589,N_15804,N_15328);
nor U16590 (N_16590,N_15701,N_15481);
xnor U16591 (N_16591,N_14245,N_14198);
and U16592 (N_16592,N_15771,N_15671);
or U16593 (N_16593,N_14235,N_15982);
or U16594 (N_16594,N_14363,N_15678);
nor U16595 (N_16595,N_15363,N_15086);
xnor U16596 (N_16596,N_14575,N_14340);
xor U16597 (N_16597,N_15104,N_15334);
nor U16598 (N_16598,N_14306,N_15463);
nand U16599 (N_16599,N_15338,N_15524);
nand U16600 (N_16600,N_14345,N_15020);
or U16601 (N_16601,N_14992,N_14293);
nand U16602 (N_16602,N_14631,N_14099);
and U16603 (N_16603,N_14495,N_14935);
xnor U16604 (N_16604,N_15055,N_15240);
or U16605 (N_16605,N_15304,N_15589);
xnor U16606 (N_16606,N_14707,N_15167);
and U16607 (N_16607,N_15843,N_14955);
xor U16608 (N_16608,N_14597,N_15987);
nor U16609 (N_16609,N_15470,N_15422);
xnor U16610 (N_16610,N_14092,N_14732);
nand U16611 (N_16611,N_14677,N_15714);
xnor U16612 (N_16612,N_15455,N_14943);
xor U16613 (N_16613,N_15927,N_14743);
and U16614 (N_16614,N_14641,N_15136);
and U16615 (N_16615,N_14142,N_14664);
and U16616 (N_16616,N_14240,N_14972);
nor U16617 (N_16617,N_14962,N_14188);
xor U16618 (N_16618,N_14222,N_15427);
nand U16619 (N_16619,N_15622,N_14173);
nor U16620 (N_16620,N_15336,N_14223);
xor U16621 (N_16621,N_14553,N_14081);
nand U16622 (N_16622,N_14255,N_15305);
or U16623 (N_16623,N_15155,N_14217);
or U16624 (N_16624,N_14149,N_14692);
nand U16625 (N_16625,N_15366,N_14473);
and U16626 (N_16626,N_15303,N_14028);
nand U16627 (N_16627,N_14802,N_15507);
and U16628 (N_16628,N_15327,N_14154);
xnor U16629 (N_16629,N_15759,N_15937);
xnor U16630 (N_16630,N_14579,N_14566);
or U16631 (N_16631,N_14990,N_15088);
nor U16632 (N_16632,N_15066,N_14541);
nand U16633 (N_16633,N_14736,N_15321);
xnor U16634 (N_16634,N_14106,N_15757);
nor U16635 (N_16635,N_15916,N_15264);
xnor U16636 (N_16636,N_14914,N_15944);
and U16637 (N_16637,N_15397,N_15448);
nand U16638 (N_16638,N_15504,N_15514);
xor U16639 (N_16639,N_15903,N_15857);
nand U16640 (N_16640,N_14393,N_15425);
or U16641 (N_16641,N_14561,N_15868);
or U16642 (N_16642,N_15407,N_14834);
or U16643 (N_16643,N_15750,N_14491);
xnor U16644 (N_16644,N_14494,N_14536);
nand U16645 (N_16645,N_14724,N_15456);
nor U16646 (N_16646,N_15468,N_15386);
and U16647 (N_16647,N_15211,N_14314);
nor U16648 (N_16648,N_14233,N_15217);
and U16649 (N_16649,N_14398,N_14152);
or U16650 (N_16650,N_14581,N_15791);
xnor U16651 (N_16651,N_15494,N_15893);
nor U16652 (N_16652,N_14875,N_14810);
nor U16653 (N_16653,N_14098,N_15139);
and U16654 (N_16654,N_15890,N_14973);
and U16655 (N_16655,N_15991,N_15100);
nor U16656 (N_16656,N_14231,N_15362);
nand U16657 (N_16657,N_15308,N_14209);
xor U16658 (N_16658,N_14760,N_14825);
xor U16659 (N_16659,N_14849,N_15706);
nor U16660 (N_16660,N_15135,N_14562);
xnor U16661 (N_16661,N_15293,N_15011);
and U16662 (N_16662,N_14674,N_15325);
nand U16663 (N_16663,N_14504,N_15774);
xor U16664 (N_16664,N_14397,N_15196);
nor U16665 (N_16665,N_14776,N_15059);
and U16666 (N_16666,N_14487,N_15915);
and U16667 (N_16667,N_15449,N_15983);
or U16668 (N_16668,N_15190,N_14275);
and U16669 (N_16669,N_14630,N_15352);
or U16670 (N_16670,N_14589,N_15860);
or U16671 (N_16671,N_14246,N_15900);
xnor U16672 (N_16672,N_14192,N_14339);
or U16673 (N_16673,N_14956,N_14531);
nor U16674 (N_16674,N_15292,N_14137);
and U16675 (N_16675,N_14608,N_14178);
nand U16676 (N_16676,N_15323,N_14034);
nor U16677 (N_16677,N_14187,N_15616);
xnor U16678 (N_16678,N_14197,N_15411);
and U16679 (N_16679,N_15501,N_14374);
xor U16680 (N_16680,N_15823,N_14261);
nor U16681 (N_16681,N_15461,N_15333);
or U16682 (N_16682,N_15152,N_14278);
and U16683 (N_16683,N_15607,N_15729);
or U16684 (N_16684,N_15673,N_15973);
nor U16685 (N_16685,N_15884,N_14200);
nor U16686 (N_16686,N_14277,N_15282);
or U16687 (N_16687,N_14199,N_14214);
nor U16688 (N_16688,N_14003,N_14343);
and U16689 (N_16689,N_15358,N_14888);
nor U16690 (N_16690,N_15579,N_14421);
or U16691 (N_16691,N_15290,N_14100);
xnor U16692 (N_16692,N_14162,N_15789);
nor U16693 (N_16693,N_15406,N_14311);
or U16694 (N_16694,N_15040,N_15193);
nor U16695 (N_16695,N_15948,N_15984);
and U16696 (N_16696,N_14153,N_14715);
or U16697 (N_16697,N_15063,N_14463);
nor U16698 (N_16698,N_15071,N_15989);
nand U16699 (N_16699,N_14292,N_15684);
nand U16700 (N_16700,N_15294,N_15513);
nand U16701 (N_16701,N_14170,N_15440);
and U16702 (N_16702,N_14866,N_15999);
xnor U16703 (N_16703,N_14196,N_14309);
or U16704 (N_16704,N_15374,N_15484);
and U16705 (N_16705,N_14503,N_14870);
and U16706 (N_16706,N_15199,N_14512);
or U16707 (N_16707,N_15847,N_15905);
and U16708 (N_16708,N_14418,N_14122);
nor U16709 (N_16709,N_15640,N_15478);
and U16710 (N_16710,N_15320,N_14572);
xor U16711 (N_16711,N_15262,N_15530);
xnor U16712 (N_16712,N_15660,N_15306);
nor U16713 (N_16713,N_15742,N_14161);
and U16714 (N_16714,N_15739,N_14757);
and U16715 (N_16715,N_14697,N_14587);
nand U16716 (N_16716,N_15656,N_14021);
or U16717 (N_16717,N_15452,N_15010);
nor U16718 (N_16718,N_14940,N_15545);
or U16719 (N_16719,N_14210,N_14336);
nand U16720 (N_16720,N_14864,N_15435);
xor U16721 (N_16721,N_14578,N_14605);
xnor U16722 (N_16722,N_14009,N_14431);
and U16723 (N_16723,N_15500,N_14999);
nor U16724 (N_16724,N_14527,N_14366);
nor U16725 (N_16725,N_15488,N_14773);
nand U16726 (N_16726,N_15415,N_15067);
and U16727 (N_16727,N_14284,N_14415);
nor U16728 (N_16728,N_15547,N_15812);
xor U16729 (N_16729,N_15426,N_14051);
nand U16730 (N_16730,N_15434,N_14831);
xnor U16731 (N_16731,N_15235,N_14219);
and U16732 (N_16732,N_15816,N_14297);
nand U16733 (N_16733,N_15598,N_15768);
xor U16734 (N_16734,N_15649,N_15385);
and U16735 (N_16735,N_14637,N_14190);
xnor U16736 (N_16736,N_15288,N_14917);
xnor U16737 (N_16737,N_15258,N_14764);
nand U16738 (N_16738,N_15802,N_14836);
nor U16739 (N_16739,N_14030,N_14364);
xnor U16740 (N_16740,N_15891,N_14520);
or U16741 (N_16741,N_15613,N_14004);
nor U16742 (N_16742,N_14728,N_15605);
or U16743 (N_16743,N_14259,N_14307);
nor U16744 (N_16744,N_14514,N_15734);
and U16745 (N_16745,N_14879,N_14054);
nand U16746 (N_16746,N_15095,N_14577);
nor U16747 (N_16747,N_14951,N_15652);
and U16748 (N_16748,N_14458,N_14203);
nor U16749 (N_16749,N_15615,N_14927);
nand U16750 (N_16750,N_14484,N_15050);
or U16751 (N_16751,N_14186,N_14296);
nor U16752 (N_16752,N_14693,N_15772);
or U16753 (N_16753,N_15740,N_15079);
nor U16754 (N_16754,N_15444,N_14915);
nor U16755 (N_16755,N_15377,N_15175);
xnor U16756 (N_16756,N_14155,N_14971);
nand U16757 (N_16757,N_14548,N_15582);
and U16758 (N_16758,N_14338,N_15118);
and U16759 (N_16759,N_15219,N_14515);
and U16760 (N_16760,N_14299,N_15623);
or U16761 (N_16761,N_15113,N_15975);
xor U16762 (N_16762,N_15588,N_15941);
or U16763 (N_16763,N_14365,N_14396);
nand U16764 (N_16764,N_14123,N_15182);
xor U16765 (N_16765,N_15849,N_14932);
xor U16766 (N_16766,N_14305,N_14961);
nor U16767 (N_16767,N_14612,N_14778);
nand U16768 (N_16768,N_15301,N_14148);
nor U16769 (N_16769,N_15688,N_14718);
or U16770 (N_16770,N_14276,N_15924);
xnor U16771 (N_16771,N_15223,N_14833);
nand U16772 (N_16772,N_15672,N_14710);
xnor U16773 (N_16773,N_15224,N_15680);
or U16774 (N_16774,N_14357,N_14460);
nor U16775 (N_16775,N_14889,N_14061);
nand U16776 (N_16776,N_15648,N_15553);
nor U16777 (N_16777,N_14133,N_15072);
nor U16778 (N_16778,N_15457,N_15970);
and U16779 (N_16779,N_14528,N_15705);
or U16780 (N_16780,N_14700,N_14459);
or U16781 (N_16781,N_15028,N_14164);
nand U16782 (N_16782,N_15360,N_14969);
and U16783 (N_16783,N_15632,N_15535);
or U16784 (N_16784,N_14957,N_15643);
or U16785 (N_16785,N_14635,N_15986);
and U16786 (N_16786,N_15962,N_15096);
and U16787 (N_16787,N_14228,N_15778);
nor U16788 (N_16788,N_15506,N_15421);
or U16789 (N_16789,N_14838,N_14851);
xor U16790 (N_16790,N_14163,N_15639);
nor U16791 (N_16791,N_14948,N_14899);
or U16792 (N_16792,N_15098,N_15560);
and U16793 (N_16793,N_15957,N_14312);
or U16794 (N_16794,N_15353,N_15370);
nor U16795 (N_16795,N_14678,N_14241);
nor U16796 (N_16796,N_14511,N_15747);
and U16797 (N_16797,N_15215,N_14850);
nand U16798 (N_16798,N_14960,N_15951);
nand U16799 (N_16799,N_14391,N_14236);
or U16800 (N_16800,N_14243,N_14855);
xnor U16801 (N_16801,N_14726,N_14379);
and U16802 (N_16802,N_15940,N_14472);
xor U16803 (N_16803,N_15979,N_14979);
xor U16804 (N_16804,N_15164,N_14430);
xor U16805 (N_16805,N_14769,N_14997);
or U16806 (N_16806,N_15592,N_14202);
nor U16807 (N_16807,N_14360,N_15168);
nor U16808 (N_16808,N_14370,N_15038);
or U16809 (N_16809,N_15779,N_15546);
and U16810 (N_16810,N_14911,N_14964);
nor U16811 (N_16811,N_14377,N_14168);
and U16812 (N_16812,N_15073,N_14445);
and U16813 (N_16813,N_14403,N_14216);
or U16814 (N_16814,N_15094,N_14788);
nor U16815 (N_16815,N_14785,N_15064);
and U16816 (N_16816,N_15669,N_15054);
xnor U16817 (N_16817,N_14912,N_15949);
xnor U16818 (N_16818,N_14617,N_15593);
xnor U16819 (N_16819,N_14271,N_15286);
xor U16820 (N_16820,N_14105,N_14258);
and U16821 (N_16821,N_15926,N_15130);
and U16822 (N_16822,N_14916,N_14611);
nand U16823 (N_16823,N_14344,N_14779);
or U16824 (N_16824,N_15283,N_15330);
nor U16825 (N_16825,N_15511,N_14253);
and U16826 (N_16826,N_15574,N_15955);
or U16827 (N_16827,N_14794,N_14516);
nor U16828 (N_16828,N_14254,N_15247);
nand U16829 (N_16829,N_14614,N_15663);
nand U16830 (N_16830,N_14652,N_15509);
nand U16831 (N_16831,N_14656,N_15295);
or U16832 (N_16832,N_15901,N_14471);
or U16833 (N_16833,N_15137,N_15810);
xor U16834 (N_16834,N_15015,N_14399);
xnor U16835 (N_16835,N_14129,N_14967);
nor U16836 (N_16836,N_15346,N_15534);
nor U16837 (N_16837,N_15230,N_15736);
and U16838 (N_16838,N_14465,N_14650);
or U16839 (N_16839,N_15832,N_14847);
nand U16840 (N_16840,N_14634,N_15060);
nor U16841 (N_16841,N_15231,N_15471);
or U16842 (N_16842,N_14318,N_14367);
nand U16843 (N_16843,N_15821,N_15032);
nand U16844 (N_16844,N_14513,N_14649);
nor U16845 (N_16845,N_15117,N_14428);
and U16846 (N_16846,N_15815,N_15236);
and U16847 (N_16847,N_15851,N_15316);
nand U16848 (N_16848,N_15380,N_14282);
and U16849 (N_16849,N_14983,N_15533);
nand U16850 (N_16850,N_14266,N_14002);
xor U16851 (N_16851,N_15911,N_15383);
or U16852 (N_16852,N_14179,N_14968);
or U16853 (N_16853,N_15061,N_15551);
and U16854 (N_16854,N_14263,N_15787);
xor U16855 (N_16855,N_15795,N_15599);
and U16856 (N_16856,N_15166,N_14538);
nor U16857 (N_16857,N_15874,N_15708);
xnor U16858 (N_16858,N_15150,N_15221);
xor U16859 (N_16859,N_15552,N_14627);
and U16860 (N_16860,N_14119,N_14696);
or U16861 (N_16861,N_15056,N_15128);
nor U16862 (N_16862,N_15657,N_15052);
nand U16863 (N_16863,N_14793,N_15817);
nor U16864 (N_16864,N_14490,N_15246);
nor U16865 (N_16865,N_14095,N_15963);
nor U16866 (N_16866,N_15713,N_14517);
nand U16867 (N_16867,N_14424,N_15637);
nand U16868 (N_16868,N_15722,N_14883);
and U16869 (N_16869,N_14049,N_15580);
nor U16870 (N_16870,N_15754,N_14526);
xor U16871 (N_16871,N_15396,N_15917);
nor U16872 (N_16872,N_15392,N_14476);
xor U16873 (N_16873,N_14858,N_14001);
xnor U16874 (N_16874,N_15349,N_15777);
nand U16875 (N_16875,N_15990,N_14582);
xor U16876 (N_16876,N_15610,N_15700);
nor U16877 (N_16877,N_14546,N_14440);
nor U16878 (N_16878,N_15542,N_14671);
and U16879 (N_16879,N_15213,N_15004);
or U16880 (N_16880,N_14694,N_15458);
xor U16881 (N_16881,N_15356,N_14470);
xor U16882 (N_16882,N_15928,N_15559);
nand U16883 (N_16883,N_14701,N_14523);
or U16884 (N_16884,N_14544,N_15502);
nor U16885 (N_16885,N_14813,N_14754);
nand U16886 (N_16886,N_14874,N_15958);
nor U16887 (N_16887,N_15428,N_15077);
and U16888 (N_16888,N_15093,N_14551);
or U16889 (N_16889,N_15540,N_15871);
xor U16890 (N_16890,N_14423,N_14373);
nor U16891 (N_16891,N_15331,N_14532);
xor U16892 (N_16892,N_14409,N_14272);
and U16893 (N_16893,N_15267,N_15698);
and U16894 (N_16894,N_15896,N_15889);
and U16895 (N_16895,N_14372,N_15642);
or U16896 (N_16896,N_15717,N_14591);
nor U16897 (N_16897,N_14500,N_15558);
nand U16898 (N_16898,N_14417,N_15612);
or U16899 (N_16899,N_14175,N_15689);
xor U16900 (N_16900,N_15026,N_15183);
nor U16901 (N_16901,N_15862,N_14644);
nand U16902 (N_16902,N_15257,N_14492);
and U16903 (N_16903,N_15784,N_15253);
and U16904 (N_16904,N_15176,N_14388);
and U16905 (N_16905,N_14438,N_15134);
xor U16906 (N_16906,N_14006,N_15255);
xor U16907 (N_16907,N_14952,N_14169);
nand U16908 (N_16908,N_14074,N_15016);
xor U16909 (N_16909,N_15519,N_15841);
or U16910 (N_16910,N_14573,N_15875);
and U16911 (N_16911,N_14479,N_14629);
or U16912 (N_16912,N_14348,N_15876);
nor U16913 (N_16913,N_15550,N_15309);
or U16914 (N_16914,N_14525,N_14713);
nor U16915 (N_16915,N_15564,N_15281);
nand U16916 (N_16916,N_14434,N_15676);
and U16917 (N_16917,N_14044,N_14124);
nand U16918 (N_16918,N_15495,N_15239);
or U16919 (N_16919,N_14919,N_15216);
xor U16920 (N_16920,N_14355,N_14596);
and U16921 (N_16921,N_14029,N_14486);
or U16922 (N_16922,N_14065,N_15153);
and U16923 (N_16923,N_15827,N_14837);
or U16924 (N_16924,N_14505,N_15205);
and U16925 (N_16925,N_14708,N_14685);
nand U16926 (N_16926,N_14265,N_15389);
nor U16927 (N_16927,N_15181,N_14158);
or U16928 (N_16928,N_14086,N_14036);
xor U16929 (N_16929,N_14134,N_14930);
xnor U16930 (N_16930,N_15934,N_14446);
nand U16931 (N_16931,N_14406,N_14725);
or U16932 (N_16932,N_14251,N_15466);
nor U16933 (N_16933,N_15647,N_14721);
nor U16934 (N_16934,N_15172,N_15275);
nor U16935 (N_16935,N_14537,N_14020);
xor U16936 (N_16936,N_14901,N_14070);
and U16937 (N_16937,N_14218,N_14096);
nand U16938 (N_16938,N_15241,N_15856);
nand U16939 (N_16939,N_14928,N_14425);
and U16940 (N_16940,N_14539,N_15018);
or U16941 (N_16941,N_14358,N_15256);
nand U16942 (N_16942,N_14031,N_14772);
xnor U16943 (N_16943,N_14371,N_15568);
or U16944 (N_16944,N_15883,N_14264);
or U16945 (N_16945,N_15486,N_14672);
xor U16946 (N_16946,N_14683,N_14991);
nor U16947 (N_16947,N_14475,N_15345);
and U16948 (N_16948,N_14327,N_14942);
and U16949 (N_16949,N_15178,N_15265);
xnor U16950 (N_16950,N_15686,N_14753);
and U16951 (N_16951,N_14594,N_15859);
or U16952 (N_16952,N_15733,N_14023);
or U16953 (N_16953,N_15626,N_15107);
or U16954 (N_16954,N_14069,N_14452);
and U16955 (N_16955,N_15696,N_15250);
or U16956 (N_16956,N_15367,N_14817);
and U16957 (N_16957,N_15119,N_14872);
nand U16958 (N_16958,N_15259,N_15087);
nor U16959 (N_16959,N_15848,N_14354);
nand U16960 (N_16960,N_14461,N_15798);
nand U16961 (N_16961,N_15447,N_14936);
or U16962 (N_16962,N_14549,N_14320);
xor U16963 (N_16963,N_14420,N_15781);
xor U16964 (N_16964,N_15438,N_14821);
nor U16965 (N_16965,N_15165,N_14868);
and U16966 (N_16966,N_14560,N_15227);
nor U16967 (N_16967,N_15296,N_14535);
nor U16968 (N_16968,N_15988,N_14262);
nand U16969 (N_16969,N_15423,N_14012);
or U16970 (N_16970,N_15510,N_14249);
nand U16971 (N_16971,N_15131,N_15825);
or U16972 (N_16972,N_15123,N_14680);
or U16973 (N_16973,N_14130,N_14066);
nand U16974 (N_16974,N_15829,N_14267);
or U16975 (N_16975,N_14378,N_15033);
nor U16976 (N_16976,N_14816,N_14025);
nor U16977 (N_16977,N_14039,N_14024);
nand U16978 (N_16978,N_14949,N_14620);
or U16979 (N_16979,N_15149,N_14062);
xor U16980 (N_16980,N_15390,N_15127);
nor U16981 (N_16981,N_14811,N_14191);
and U16982 (N_16982,N_15835,N_15132);
or U16983 (N_16983,N_14994,N_14807);
xnor U16984 (N_16984,N_15144,N_14185);
nand U16985 (N_16985,N_15084,N_15162);
and U16986 (N_16986,N_15604,N_15375);
and U16987 (N_16987,N_15082,N_15203);
nor U16988 (N_16988,N_15609,N_14626);
or U16989 (N_16989,N_14583,N_14665);
nor U16990 (N_16990,N_14467,N_14667);
nand U16991 (N_16991,N_15171,N_15644);
and U16992 (N_16992,N_15855,N_15212);
nor U16993 (N_16993,N_14703,N_14319);
or U16994 (N_16994,N_15142,N_15225);
or U16995 (N_16995,N_15824,N_15046);
or U16996 (N_16996,N_14496,N_14686);
xor U16997 (N_16997,N_15665,N_14640);
nand U16998 (N_16998,N_15776,N_14661);
and U16999 (N_16999,N_14653,N_15105);
and U17000 (N_17000,N_14901,N_15478);
xnor U17001 (N_17001,N_15709,N_15277);
nor U17002 (N_17002,N_14057,N_14751);
xnor U17003 (N_17003,N_15531,N_14704);
nand U17004 (N_17004,N_15455,N_14956);
and U17005 (N_17005,N_15612,N_14823);
or U17006 (N_17006,N_14155,N_14375);
xor U17007 (N_17007,N_15334,N_15006);
and U17008 (N_17008,N_14650,N_15683);
and U17009 (N_17009,N_15505,N_14458);
nor U17010 (N_17010,N_14381,N_14628);
xnor U17011 (N_17011,N_14869,N_15505);
or U17012 (N_17012,N_15515,N_15877);
nand U17013 (N_17013,N_15930,N_14914);
or U17014 (N_17014,N_15659,N_14077);
nor U17015 (N_17015,N_14690,N_14825);
and U17016 (N_17016,N_15513,N_14203);
and U17017 (N_17017,N_15849,N_15321);
nor U17018 (N_17018,N_15839,N_15407);
nor U17019 (N_17019,N_14619,N_15500);
or U17020 (N_17020,N_14013,N_14135);
xnor U17021 (N_17021,N_14258,N_14423);
nand U17022 (N_17022,N_14233,N_14063);
xor U17023 (N_17023,N_14769,N_15617);
and U17024 (N_17024,N_15895,N_15857);
nand U17025 (N_17025,N_14070,N_15296);
nor U17026 (N_17026,N_14678,N_15395);
or U17027 (N_17027,N_14473,N_14942);
xor U17028 (N_17028,N_15754,N_14334);
nor U17029 (N_17029,N_15032,N_14185);
and U17030 (N_17030,N_15626,N_14453);
nand U17031 (N_17031,N_14873,N_14280);
or U17032 (N_17032,N_15827,N_14139);
xor U17033 (N_17033,N_14266,N_15967);
nand U17034 (N_17034,N_15509,N_14376);
or U17035 (N_17035,N_15692,N_15978);
nor U17036 (N_17036,N_14398,N_15561);
nand U17037 (N_17037,N_14217,N_15319);
nand U17038 (N_17038,N_15720,N_14903);
nand U17039 (N_17039,N_15629,N_15894);
and U17040 (N_17040,N_15620,N_14663);
nor U17041 (N_17041,N_15826,N_15002);
nor U17042 (N_17042,N_15745,N_15743);
nor U17043 (N_17043,N_14098,N_15522);
nand U17044 (N_17044,N_14554,N_14325);
xnor U17045 (N_17045,N_15741,N_15801);
xor U17046 (N_17046,N_15417,N_14533);
nand U17047 (N_17047,N_14335,N_15639);
and U17048 (N_17048,N_14022,N_15251);
xnor U17049 (N_17049,N_15297,N_15349);
nor U17050 (N_17050,N_14195,N_14960);
nand U17051 (N_17051,N_15321,N_15467);
and U17052 (N_17052,N_14273,N_14945);
or U17053 (N_17053,N_15164,N_14106);
or U17054 (N_17054,N_14951,N_15982);
and U17055 (N_17055,N_14787,N_15296);
xnor U17056 (N_17056,N_15425,N_14995);
nand U17057 (N_17057,N_14227,N_14644);
xor U17058 (N_17058,N_15446,N_14137);
xor U17059 (N_17059,N_15409,N_15736);
and U17060 (N_17060,N_14477,N_14564);
nor U17061 (N_17061,N_15607,N_14814);
xnor U17062 (N_17062,N_14072,N_14195);
nand U17063 (N_17063,N_14681,N_15540);
xor U17064 (N_17064,N_14686,N_14046);
and U17065 (N_17065,N_14217,N_15310);
or U17066 (N_17066,N_14123,N_15530);
nand U17067 (N_17067,N_14227,N_15686);
and U17068 (N_17068,N_15875,N_15027);
and U17069 (N_17069,N_14336,N_14728);
or U17070 (N_17070,N_15688,N_15726);
nor U17071 (N_17071,N_15423,N_15245);
and U17072 (N_17072,N_15276,N_14488);
nand U17073 (N_17073,N_15904,N_15830);
nand U17074 (N_17074,N_14406,N_15640);
xor U17075 (N_17075,N_15295,N_14710);
nand U17076 (N_17076,N_14259,N_15760);
nand U17077 (N_17077,N_14127,N_14672);
xnor U17078 (N_17078,N_14892,N_14375);
or U17079 (N_17079,N_14023,N_14455);
nor U17080 (N_17080,N_14394,N_15037);
xor U17081 (N_17081,N_15231,N_14045);
and U17082 (N_17082,N_15562,N_14769);
and U17083 (N_17083,N_15247,N_15822);
or U17084 (N_17084,N_14707,N_14714);
xnor U17085 (N_17085,N_14703,N_14859);
and U17086 (N_17086,N_15219,N_14554);
and U17087 (N_17087,N_14301,N_15643);
nand U17088 (N_17088,N_14457,N_15670);
nand U17089 (N_17089,N_15189,N_14036);
nand U17090 (N_17090,N_14235,N_15500);
or U17091 (N_17091,N_15442,N_15906);
nand U17092 (N_17092,N_14280,N_15891);
xor U17093 (N_17093,N_15355,N_15536);
xnor U17094 (N_17094,N_15289,N_15213);
nand U17095 (N_17095,N_15003,N_15750);
xor U17096 (N_17096,N_14378,N_14231);
nand U17097 (N_17097,N_15930,N_14976);
xor U17098 (N_17098,N_14985,N_15929);
nor U17099 (N_17099,N_14752,N_15348);
and U17100 (N_17100,N_14707,N_14700);
xor U17101 (N_17101,N_14633,N_14393);
xor U17102 (N_17102,N_14705,N_15375);
nor U17103 (N_17103,N_14684,N_14605);
and U17104 (N_17104,N_14530,N_15964);
and U17105 (N_17105,N_14089,N_15867);
and U17106 (N_17106,N_14445,N_14218);
xnor U17107 (N_17107,N_14598,N_14395);
or U17108 (N_17108,N_15251,N_15618);
xnor U17109 (N_17109,N_15641,N_15775);
nand U17110 (N_17110,N_14474,N_14833);
nand U17111 (N_17111,N_14274,N_14276);
nor U17112 (N_17112,N_14988,N_14418);
and U17113 (N_17113,N_14286,N_14955);
xor U17114 (N_17114,N_14459,N_14642);
nand U17115 (N_17115,N_14863,N_15357);
xnor U17116 (N_17116,N_15894,N_14394);
xor U17117 (N_17117,N_15900,N_15047);
and U17118 (N_17118,N_14662,N_15934);
nor U17119 (N_17119,N_14083,N_15084);
and U17120 (N_17120,N_15903,N_14332);
or U17121 (N_17121,N_15095,N_14936);
nor U17122 (N_17122,N_15564,N_14608);
nand U17123 (N_17123,N_14747,N_14617);
xor U17124 (N_17124,N_14664,N_15032);
nand U17125 (N_17125,N_14655,N_14943);
xor U17126 (N_17126,N_14921,N_14637);
nor U17127 (N_17127,N_14561,N_14348);
or U17128 (N_17128,N_14161,N_14003);
and U17129 (N_17129,N_14509,N_14619);
nand U17130 (N_17130,N_14611,N_15597);
nor U17131 (N_17131,N_14546,N_14010);
nor U17132 (N_17132,N_14763,N_15473);
nand U17133 (N_17133,N_14564,N_15458);
xnor U17134 (N_17134,N_14231,N_14202);
nor U17135 (N_17135,N_15005,N_14005);
or U17136 (N_17136,N_14679,N_14216);
xnor U17137 (N_17137,N_14042,N_15279);
nor U17138 (N_17138,N_14842,N_15753);
nand U17139 (N_17139,N_14529,N_14283);
nor U17140 (N_17140,N_15748,N_15494);
xor U17141 (N_17141,N_15575,N_15191);
and U17142 (N_17142,N_14982,N_14716);
xnor U17143 (N_17143,N_15308,N_14417);
nand U17144 (N_17144,N_14409,N_14639);
nand U17145 (N_17145,N_14899,N_14859);
xnor U17146 (N_17146,N_14475,N_15207);
nand U17147 (N_17147,N_14275,N_14521);
nand U17148 (N_17148,N_15379,N_15225);
or U17149 (N_17149,N_14207,N_14897);
nand U17150 (N_17150,N_14312,N_14529);
nor U17151 (N_17151,N_15807,N_15571);
and U17152 (N_17152,N_14240,N_15557);
and U17153 (N_17153,N_15111,N_15179);
nand U17154 (N_17154,N_15281,N_15159);
nand U17155 (N_17155,N_15698,N_14609);
or U17156 (N_17156,N_14754,N_15079);
and U17157 (N_17157,N_15305,N_15455);
nor U17158 (N_17158,N_14595,N_15179);
or U17159 (N_17159,N_14683,N_14941);
and U17160 (N_17160,N_15684,N_14841);
xnor U17161 (N_17161,N_15673,N_15433);
xnor U17162 (N_17162,N_15113,N_15299);
or U17163 (N_17163,N_15747,N_15459);
nor U17164 (N_17164,N_14713,N_15289);
or U17165 (N_17165,N_15941,N_14227);
or U17166 (N_17166,N_15512,N_15822);
xor U17167 (N_17167,N_15413,N_15020);
xor U17168 (N_17168,N_15024,N_14410);
or U17169 (N_17169,N_14214,N_14377);
nor U17170 (N_17170,N_15391,N_15769);
or U17171 (N_17171,N_15381,N_14529);
nand U17172 (N_17172,N_15325,N_15936);
nand U17173 (N_17173,N_14234,N_15577);
xnor U17174 (N_17174,N_14755,N_14587);
nand U17175 (N_17175,N_15775,N_14030);
and U17176 (N_17176,N_15156,N_15769);
and U17177 (N_17177,N_14526,N_14401);
and U17178 (N_17178,N_14763,N_15532);
nand U17179 (N_17179,N_15648,N_15798);
and U17180 (N_17180,N_15276,N_15949);
and U17181 (N_17181,N_15202,N_14481);
nor U17182 (N_17182,N_15365,N_15492);
or U17183 (N_17183,N_14104,N_15407);
xor U17184 (N_17184,N_14274,N_15683);
or U17185 (N_17185,N_15180,N_15498);
nor U17186 (N_17186,N_15968,N_14104);
or U17187 (N_17187,N_15743,N_14622);
or U17188 (N_17188,N_14508,N_14672);
xor U17189 (N_17189,N_15744,N_15895);
xnor U17190 (N_17190,N_15490,N_14873);
or U17191 (N_17191,N_15180,N_15309);
and U17192 (N_17192,N_14280,N_15620);
nor U17193 (N_17193,N_15355,N_15121);
nor U17194 (N_17194,N_15688,N_14728);
nand U17195 (N_17195,N_14634,N_14981);
or U17196 (N_17196,N_15663,N_14273);
or U17197 (N_17197,N_14412,N_14397);
and U17198 (N_17198,N_14357,N_14641);
and U17199 (N_17199,N_14292,N_14353);
nor U17200 (N_17200,N_14607,N_15916);
or U17201 (N_17201,N_14555,N_14345);
xor U17202 (N_17202,N_14440,N_15162);
or U17203 (N_17203,N_15262,N_14485);
and U17204 (N_17204,N_14490,N_15600);
or U17205 (N_17205,N_15791,N_15627);
nor U17206 (N_17206,N_15550,N_14971);
or U17207 (N_17207,N_15224,N_14858);
nand U17208 (N_17208,N_14132,N_15143);
xnor U17209 (N_17209,N_15819,N_14858);
nor U17210 (N_17210,N_15979,N_14735);
or U17211 (N_17211,N_15177,N_14937);
or U17212 (N_17212,N_15794,N_14720);
xor U17213 (N_17213,N_14805,N_15945);
xor U17214 (N_17214,N_15430,N_15314);
xor U17215 (N_17215,N_15186,N_14281);
or U17216 (N_17216,N_14827,N_14561);
xor U17217 (N_17217,N_14063,N_14935);
or U17218 (N_17218,N_14654,N_15272);
and U17219 (N_17219,N_15887,N_15545);
xor U17220 (N_17220,N_15688,N_15213);
or U17221 (N_17221,N_15201,N_15472);
xnor U17222 (N_17222,N_14098,N_15744);
nand U17223 (N_17223,N_15227,N_15990);
or U17224 (N_17224,N_14032,N_15950);
nand U17225 (N_17225,N_15437,N_14290);
or U17226 (N_17226,N_15118,N_14245);
or U17227 (N_17227,N_14217,N_15378);
nand U17228 (N_17228,N_14687,N_14589);
or U17229 (N_17229,N_15596,N_14615);
or U17230 (N_17230,N_14552,N_15515);
nor U17231 (N_17231,N_14235,N_14232);
nor U17232 (N_17232,N_15069,N_15201);
or U17233 (N_17233,N_14282,N_14920);
nor U17234 (N_17234,N_14800,N_14809);
and U17235 (N_17235,N_15317,N_14433);
or U17236 (N_17236,N_15027,N_14796);
nand U17237 (N_17237,N_15883,N_14005);
xnor U17238 (N_17238,N_14960,N_14040);
and U17239 (N_17239,N_15182,N_14172);
nand U17240 (N_17240,N_14538,N_15926);
and U17241 (N_17241,N_14989,N_15542);
nor U17242 (N_17242,N_14932,N_14216);
xor U17243 (N_17243,N_15628,N_14334);
xnor U17244 (N_17244,N_15691,N_14570);
nand U17245 (N_17245,N_14676,N_15553);
nand U17246 (N_17246,N_15503,N_15081);
nand U17247 (N_17247,N_15532,N_15013);
or U17248 (N_17248,N_14973,N_14592);
nor U17249 (N_17249,N_14952,N_14886);
and U17250 (N_17250,N_15951,N_14572);
xnor U17251 (N_17251,N_15045,N_14036);
xnor U17252 (N_17252,N_14425,N_14850);
xor U17253 (N_17253,N_14614,N_15459);
and U17254 (N_17254,N_14234,N_15322);
nor U17255 (N_17255,N_15965,N_15295);
or U17256 (N_17256,N_14862,N_15618);
xnor U17257 (N_17257,N_15870,N_14343);
and U17258 (N_17258,N_14260,N_14591);
nand U17259 (N_17259,N_15469,N_15098);
and U17260 (N_17260,N_14150,N_15036);
or U17261 (N_17261,N_15536,N_15213);
nand U17262 (N_17262,N_14722,N_14429);
nor U17263 (N_17263,N_15621,N_15676);
xor U17264 (N_17264,N_15334,N_14355);
nand U17265 (N_17265,N_14309,N_15532);
or U17266 (N_17266,N_15958,N_14110);
nand U17267 (N_17267,N_14922,N_14144);
and U17268 (N_17268,N_15275,N_14642);
or U17269 (N_17269,N_14469,N_15394);
or U17270 (N_17270,N_14599,N_15169);
and U17271 (N_17271,N_14049,N_14776);
nand U17272 (N_17272,N_15813,N_14464);
xor U17273 (N_17273,N_15512,N_14744);
nor U17274 (N_17274,N_14503,N_14099);
and U17275 (N_17275,N_15036,N_14202);
nor U17276 (N_17276,N_15406,N_15676);
xor U17277 (N_17277,N_14296,N_15886);
nand U17278 (N_17278,N_14084,N_14168);
xnor U17279 (N_17279,N_14954,N_14924);
nand U17280 (N_17280,N_14909,N_15568);
xnor U17281 (N_17281,N_15572,N_15960);
xor U17282 (N_17282,N_15210,N_14896);
xor U17283 (N_17283,N_15276,N_14813);
nand U17284 (N_17284,N_15474,N_14818);
xor U17285 (N_17285,N_14026,N_15884);
nand U17286 (N_17286,N_15560,N_15296);
and U17287 (N_17287,N_14059,N_15439);
xor U17288 (N_17288,N_15508,N_15121);
and U17289 (N_17289,N_15698,N_15591);
and U17290 (N_17290,N_14532,N_15707);
and U17291 (N_17291,N_14919,N_14034);
and U17292 (N_17292,N_15211,N_15630);
and U17293 (N_17293,N_14961,N_15246);
or U17294 (N_17294,N_14193,N_15411);
nand U17295 (N_17295,N_14004,N_15051);
nand U17296 (N_17296,N_14099,N_14170);
nand U17297 (N_17297,N_14179,N_14524);
or U17298 (N_17298,N_14803,N_14236);
and U17299 (N_17299,N_14900,N_15645);
and U17300 (N_17300,N_14501,N_15726);
or U17301 (N_17301,N_15612,N_14904);
nor U17302 (N_17302,N_15240,N_14946);
or U17303 (N_17303,N_14313,N_14715);
and U17304 (N_17304,N_14572,N_15480);
nand U17305 (N_17305,N_14538,N_14887);
nor U17306 (N_17306,N_15354,N_15238);
and U17307 (N_17307,N_15235,N_15272);
xor U17308 (N_17308,N_15781,N_14203);
and U17309 (N_17309,N_15647,N_15029);
and U17310 (N_17310,N_14485,N_14805);
xor U17311 (N_17311,N_14487,N_15150);
or U17312 (N_17312,N_14731,N_14200);
and U17313 (N_17313,N_15119,N_14387);
nor U17314 (N_17314,N_14757,N_15607);
and U17315 (N_17315,N_14397,N_14011);
nor U17316 (N_17316,N_15147,N_15774);
nand U17317 (N_17317,N_14524,N_14531);
nor U17318 (N_17318,N_14497,N_14113);
nor U17319 (N_17319,N_14159,N_14955);
nor U17320 (N_17320,N_15655,N_15093);
and U17321 (N_17321,N_14125,N_15770);
nand U17322 (N_17322,N_14432,N_15258);
nor U17323 (N_17323,N_15067,N_15756);
and U17324 (N_17324,N_14918,N_14960);
nand U17325 (N_17325,N_14328,N_15806);
or U17326 (N_17326,N_14316,N_15591);
or U17327 (N_17327,N_14003,N_14968);
nor U17328 (N_17328,N_14621,N_15943);
nand U17329 (N_17329,N_14243,N_15242);
xor U17330 (N_17330,N_14783,N_14183);
or U17331 (N_17331,N_15884,N_14015);
or U17332 (N_17332,N_14801,N_14718);
nand U17333 (N_17333,N_14910,N_14080);
nand U17334 (N_17334,N_15145,N_14585);
or U17335 (N_17335,N_15297,N_14683);
and U17336 (N_17336,N_15348,N_15770);
xor U17337 (N_17337,N_15604,N_15968);
or U17338 (N_17338,N_14575,N_15020);
or U17339 (N_17339,N_15520,N_15969);
nor U17340 (N_17340,N_15505,N_15832);
and U17341 (N_17341,N_15399,N_15808);
and U17342 (N_17342,N_14147,N_15079);
or U17343 (N_17343,N_15143,N_15369);
nand U17344 (N_17344,N_14757,N_15640);
nand U17345 (N_17345,N_15366,N_14555);
or U17346 (N_17346,N_14358,N_14120);
xnor U17347 (N_17347,N_15774,N_15863);
nor U17348 (N_17348,N_14308,N_15434);
or U17349 (N_17349,N_14734,N_14126);
nor U17350 (N_17350,N_15701,N_14446);
or U17351 (N_17351,N_14127,N_14776);
nor U17352 (N_17352,N_14091,N_15975);
xor U17353 (N_17353,N_15336,N_15134);
or U17354 (N_17354,N_14735,N_15779);
or U17355 (N_17355,N_15476,N_14027);
nor U17356 (N_17356,N_15755,N_15633);
nand U17357 (N_17357,N_15977,N_15999);
nor U17358 (N_17358,N_14442,N_14304);
and U17359 (N_17359,N_14859,N_14973);
nand U17360 (N_17360,N_14600,N_15026);
xor U17361 (N_17361,N_15316,N_14334);
xnor U17362 (N_17362,N_15345,N_14776);
nor U17363 (N_17363,N_15204,N_15914);
nand U17364 (N_17364,N_15490,N_15530);
or U17365 (N_17365,N_14887,N_14597);
xnor U17366 (N_17366,N_15537,N_15302);
nor U17367 (N_17367,N_14989,N_14165);
and U17368 (N_17368,N_15931,N_14672);
nor U17369 (N_17369,N_15447,N_15925);
and U17370 (N_17370,N_15893,N_15094);
nand U17371 (N_17371,N_15533,N_15173);
and U17372 (N_17372,N_15888,N_15445);
nor U17373 (N_17373,N_14262,N_15551);
xnor U17374 (N_17374,N_14150,N_14879);
and U17375 (N_17375,N_15955,N_14888);
xor U17376 (N_17376,N_14553,N_15609);
nor U17377 (N_17377,N_14226,N_15954);
xor U17378 (N_17378,N_14054,N_14177);
nor U17379 (N_17379,N_15574,N_14461);
and U17380 (N_17380,N_15800,N_15053);
and U17381 (N_17381,N_14846,N_15065);
nor U17382 (N_17382,N_15646,N_15525);
nor U17383 (N_17383,N_14619,N_14603);
or U17384 (N_17384,N_14174,N_14366);
nand U17385 (N_17385,N_14854,N_14436);
nand U17386 (N_17386,N_14108,N_15032);
and U17387 (N_17387,N_14247,N_15248);
nor U17388 (N_17388,N_14756,N_15395);
or U17389 (N_17389,N_15751,N_15354);
or U17390 (N_17390,N_14380,N_14648);
and U17391 (N_17391,N_14427,N_15342);
nor U17392 (N_17392,N_15760,N_14561);
or U17393 (N_17393,N_14798,N_14493);
and U17394 (N_17394,N_14178,N_14785);
or U17395 (N_17395,N_15736,N_15826);
nand U17396 (N_17396,N_15689,N_14774);
xor U17397 (N_17397,N_15451,N_14724);
nor U17398 (N_17398,N_14879,N_15910);
xnor U17399 (N_17399,N_14929,N_15525);
xnor U17400 (N_17400,N_14178,N_14441);
nand U17401 (N_17401,N_14862,N_14910);
nor U17402 (N_17402,N_15628,N_14051);
and U17403 (N_17403,N_14927,N_15286);
or U17404 (N_17404,N_15542,N_15958);
or U17405 (N_17405,N_15148,N_14246);
and U17406 (N_17406,N_15671,N_14581);
nand U17407 (N_17407,N_15063,N_14234);
xnor U17408 (N_17408,N_15560,N_15725);
nor U17409 (N_17409,N_15303,N_14592);
nor U17410 (N_17410,N_15963,N_14926);
xor U17411 (N_17411,N_14609,N_14399);
or U17412 (N_17412,N_15971,N_14829);
and U17413 (N_17413,N_14690,N_15661);
nand U17414 (N_17414,N_14786,N_15153);
and U17415 (N_17415,N_15164,N_15229);
and U17416 (N_17416,N_15139,N_15264);
xnor U17417 (N_17417,N_15299,N_14355);
xor U17418 (N_17418,N_14602,N_15858);
nand U17419 (N_17419,N_15728,N_14575);
xnor U17420 (N_17420,N_14466,N_14051);
and U17421 (N_17421,N_14251,N_14787);
nor U17422 (N_17422,N_14994,N_15164);
nor U17423 (N_17423,N_15113,N_15554);
nor U17424 (N_17424,N_14593,N_15113);
nor U17425 (N_17425,N_14158,N_15564);
nand U17426 (N_17426,N_14632,N_14600);
nand U17427 (N_17427,N_15128,N_14352);
xor U17428 (N_17428,N_15654,N_14140);
and U17429 (N_17429,N_14549,N_15653);
nor U17430 (N_17430,N_14317,N_15346);
or U17431 (N_17431,N_14201,N_15108);
or U17432 (N_17432,N_15513,N_14765);
nand U17433 (N_17433,N_15243,N_14659);
xor U17434 (N_17434,N_15749,N_14598);
or U17435 (N_17435,N_14902,N_14713);
xnor U17436 (N_17436,N_15966,N_14491);
and U17437 (N_17437,N_14293,N_15107);
nor U17438 (N_17438,N_14654,N_14149);
nand U17439 (N_17439,N_15722,N_15190);
and U17440 (N_17440,N_15598,N_15463);
nand U17441 (N_17441,N_15664,N_15591);
nor U17442 (N_17442,N_14809,N_14741);
nor U17443 (N_17443,N_15587,N_14341);
nand U17444 (N_17444,N_15074,N_14311);
xor U17445 (N_17445,N_14468,N_15320);
nand U17446 (N_17446,N_14534,N_14805);
nand U17447 (N_17447,N_15470,N_14877);
and U17448 (N_17448,N_15656,N_14747);
nand U17449 (N_17449,N_14346,N_15997);
xnor U17450 (N_17450,N_14892,N_14096);
nor U17451 (N_17451,N_15183,N_14418);
nor U17452 (N_17452,N_15429,N_15126);
nor U17453 (N_17453,N_14365,N_14370);
and U17454 (N_17454,N_15344,N_15871);
nor U17455 (N_17455,N_14871,N_15477);
nand U17456 (N_17456,N_15072,N_15521);
nand U17457 (N_17457,N_14093,N_14027);
or U17458 (N_17458,N_15932,N_14228);
nor U17459 (N_17459,N_14255,N_14566);
and U17460 (N_17460,N_15516,N_15295);
or U17461 (N_17461,N_15616,N_15424);
xor U17462 (N_17462,N_14613,N_15744);
and U17463 (N_17463,N_15597,N_14509);
nor U17464 (N_17464,N_15281,N_15395);
nand U17465 (N_17465,N_14508,N_15760);
nor U17466 (N_17466,N_15936,N_14078);
nor U17467 (N_17467,N_15428,N_15067);
and U17468 (N_17468,N_14872,N_15635);
nand U17469 (N_17469,N_14432,N_15337);
and U17470 (N_17470,N_15487,N_14308);
and U17471 (N_17471,N_15260,N_14125);
nand U17472 (N_17472,N_15974,N_14823);
or U17473 (N_17473,N_14641,N_15806);
xnor U17474 (N_17474,N_15189,N_15956);
xor U17475 (N_17475,N_15205,N_15242);
and U17476 (N_17476,N_14456,N_14544);
nand U17477 (N_17477,N_15708,N_14600);
nor U17478 (N_17478,N_15574,N_15998);
nor U17479 (N_17479,N_14908,N_14545);
xnor U17480 (N_17480,N_14722,N_14519);
and U17481 (N_17481,N_14735,N_15013);
or U17482 (N_17482,N_15441,N_14530);
nand U17483 (N_17483,N_15920,N_14067);
or U17484 (N_17484,N_14053,N_14158);
or U17485 (N_17485,N_15395,N_14565);
nor U17486 (N_17486,N_14184,N_15269);
xor U17487 (N_17487,N_15058,N_14355);
xnor U17488 (N_17488,N_15206,N_14120);
or U17489 (N_17489,N_14746,N_15042);
nor U17490 (N_17490,N_15318,N_15252);
xnor U17491 (N_17491,N_14763,N_15220);
nor U17492 (N_17492,N_15306,N_15360);
nand U17493 (N_17493,N_15031,N_15945);
nand U17494 (N_17494,N_14274,N_15750);
nand U17495 (N_17495,N_15008,N_15927);
xnor U17496 (N_17496,N_14906,N_14187);
or U17497 (N_17497,N_14379,N_14378);
xnor U17498 (N_17498,N_14063,N_15925);
or U17499 (N_17499,N_14158,N_15780);
and U17500 (N_17500,N_14856,N_14316);
nand U17501 (N_17501,N_14873,N_14299);
xor U17502 (N_17502,N_15759,N_14025);
and U17503 (N_17503,N_14205,N_15530);
and U17504 (N_17504,N_15844,N_15505);
or U17505 (N_17505,N_15560,N_14890);
xor U17506 (N_17506,N_14009,N_14076);
nand U17507 (N_17507,N_14674,N_15081);
and U17508 (N_17508,N_15235,N_14689);
or U17509 (N_17509,N_15768,N_14277);
and U17510 (N_17510,N_15314,N_15548);
nand U17511 (N_17511,N_15905,N_14966);
nor U17512 (N_17512,N_14835,N_15878);
or U17513 (N_17513,N_14818,N_15669);
nor U17514 (N_17514,N_14762,N_14586);
nor U17515 (N_17515,N_14591,N_14292);
nand U17516 (N_17516,N_15686,N_14983);
and U17517 (N_17517,N_15216,N_14057);
and U17518 (N_17518,N_14062,N_15270);
nand U17519 (N_17519,N_15827,N_15122);
xnor U17520 (N_17520,N_15303,N_14288);
or U17521 (N_17521,N_14555,N_15370);
xnor U17522 (N_17522,N_15148,N_14495);
and U17523 (N_17523,N_15708,N_15510);
and U17524 (N_17524,N_15350,N_14808);
and U17525 (N_17525,N_14647,N_15517);
nand U17526 (N_17526,N_15189,N_14950);
nor U17527 (N_17527,N_14392,N_15521);
or U17528 (N_17528,N_15909,N_14042);
and U17529 (N_17529,N_14173,N_14144);
xnor U17530 (N_17530,N_14531,N_15384);
nor U17531 (N_17531,N_14694,N_15380);
or U17532 (N_17532,N_15895,N_15643);
nand U17533 (N_17533,N_14664,N_15905);
nand U17534 (N_17534,N_14494,N_15744);
xor U17535 (N_17535,N_15671,N_15767);
nand U17536 (N_17536,N_14412,N_15045);
xnor U17537 (N_17537,N_15873,N_14396);
xor U17538 (N_17538,N_14915,N_15139);
xnor U17539 (N_17539,N_14699,N_15865);
or U17540 (N_17540,N_15934,N_14331);
nor U17541 (N_17541,N_14180,N_14299);
nand U17542 (N_17542,N_15675,N_14053);
nor U17543 (N_17543,N_15783,N_15435);
xor U17544 (N_17544,N_14526,N_14274);
or U17545 (N_17545,N_14351,N_14465);
xnor U17546 (N_17546,N_14601,N_14972);
xor U17547 (N_17547,N_15181,N_14775);
or U17548 (N_17548,N_15079,N_15634);
xor U17549 (N_17549,N_15744,N_15013);
and U17550 (N_17550,N_14479,N_15230);
xor U17551 (N_17551,N_15600,N_14803);
xnor U17552 (N_17552,N_14058,N_15477);
nor U17553 (N_17553,N_15585,N_15624);
or U17554 (N_17554,N_15767,N_14109);
nor U17555 (N_17555,N_15222,N_14526);
nand U17556 (N_17556,N_14950,N_14211);
xnor U17557 (N_17557,N_14707,N_15255);
nor U17558 (N_17558,N_15970,N_15645);
and U17559 (N_17559,N_15764,N_14204);
xnor U17560 (N_17560,N_14282,N_15070);
xor U17561 (N_17561,N_14474,N_14384);
nor U17562 (N_17562,N_14536,N_14723);
nand U17563 (N_17563,N_14092,N_15066);
xor U17564 (N_17564,N_14554,N_14321);
or U17565 (N_17565,N_14789,N_15541);
or U17566 (N_17566,N_15597,N_14784);
or U17567 (N_17567,N_15096,N_15594);
xor U17568 (N_17568,N_15242,N_14519);
xor U17569 (N_17569,N_14760,N_14221);
xnor U17570 (N_17570,N_14917,N_14597);
nand U17571 (N_17571,N_14954,N_14392);
nor U17572 (N_17572,N_14328,N_15423);
nand U17573 (N_17573,N_14547,N_15087);
nand U17574 (N_17574,N_14701,N_15958);
and U17575 (N_17575,N_14478,N_15137);
nor U17576 (N_17576,N_14036,N_15260);
or U17577 (N_17577,N_14486,N_15143);
nand U17578 (N_17578,N_15787,N_14295);
xor U17579 (N_17579,N_15139,N_14198);
and U17580 (N_17580,N_15143,N_15652);
nor U17581 (N_17581,N_14549,N_15934);
nand U17582 (N_17582,N_15407,N_14742);
or U17583 (N_17583,N_14754,N_14116);
or U17584 (N_17584,N_14905,N_15753);
and U17585 (N_17585,N_14325,N_14843);
xnor U17586 (N_17586,N_15975,N_15696);
xnor U17587 (N_17587,N_14167,N_15450);
and U17588 (N_17588,N_14227,N_15217);
xor U17589 (N_17589,N_14220,N_15479);
nor U17590 (N_17590,N_15260,N_15021);
xor U17591 (N_17591,N_15571,N_15955);
nor U17592 (N_17592,N_14430,N_14782);
nor U17593 (N_17593,N_15032,N_14593);
and U17594 (N_17594,N_14446,N_14500);
xnor U17595 (N_17595,N_14390,N_15153);
nor U17596 (N_17596,N_15371,N_14732);
or U17597 (N_17597,N_14085,N_15365);
xnor U17598 (N_17598,N_14119,N_15352);
and U17599 (N_17599,N_14708,N_14491);
xnor U17600 (N_17600,N_14394,N_14425);
nand U17601 (N_17601,N_15565,N_14647);
and U17602 (N_17602,N_14480,N_15377);
nor U17603 (N_17603,N_14423,N_14989);
and U17604 (N_17604,N_14003,N_15204);
or U17605 (N_17605,N_14662,N_15756);
or U17606 (N_17606,N_14954,N_15709);
nand U17607 (N_17607,N_15401,N_15583);
xor U17608 (N_17608,N_15334,N_14409);
or U17609 (N_17609,N_15680,N_14641);
and U17610 (N_17610,N_15399,N_14224);
nand U17611 (N_17611,N_15402,N_14666);
or U17612 (N_17612,N_14129,N_14959);
nor U17613 (N_17613,N_14785,N_15451);
and U17614 (N_17614,N_14736,N_14862);
nor U17615 (N_17615,N_15221,N_15710);
nor U17616 (N_17616,N_15052,N_15916);
xor U17617 (N_17617,N_14460,N_15536);
nand U17618 (N_17618,N_15069,N_14007);
and U17619 (N_17619,N_14842,N_15335);
and U17620 (N_17620,N_15516,N_14298);
nand U17621 (N_17621,N_14291,N_15993);
nand U17622 (N_17622,N_14472,N_15549);
nand U17623 (N_17623,N_15067,N_15863);
or U17624 (N_17624,N_15706,N_14518);
nor U17625 (N_17625,N_14288,N_14364);
nor U17626 (N_17626,N_15836,N_14495);
nor U17627 (N_17627,N_15648,N_14303);
xor U17628 (N_17628,N_15076,N_14942);
nand U17629 (N_17629,N_14042,N_15986);
and U17630 (N_17630,N_14378,N_14127);
xor U17631 (N_17631,N_15320,N_14991);
xor U17632 (N_17632,N_14762,N_14165);
xnor U17633 (N_17633,N_15777,N_15915);
and U17634 (N_17634,N_15261,N_14425);
nand U17635 (N_17635,N_14934,N_14598);
xnor U17636 (N_17636,N_15094,N_15504);
nor U17637 (N_17637,N_15571,N_15809);
xnor U17638 (N_17638,N_15853,N_15783);
xor U17639 (N_17639,N_14807,N_14295);
nand U17640 (N_17640,N_14003,N_14916);
nor U17641 (N_17641,N_15131,N_15798);
xor U17642 (N_17642,N_15913,N_15959);
nand U17643 (N_17643,N_15762,N_15793);
and U17644 (N_17644,N_14035,N_14843);
nor U17645 (N_17645,N_15937,N_15786);
nand U17646 (N_17646,N_14847,N_15535);
nor U17647 (N_17647,N_15007,N_15422);
xor U17648 (N_17648,N_14491,N_15052);
nand U17649 (N_17649,N_14041,N_15437);
or U17650 (N_17650,N_15152,N_14032);
xor U17651 (N_17651,N_14036,N_15739);
or U17652 (N_17652,N_14585,N_15292);
xnor U17653 (N_17653,N_14985,N_14191);
nor U17654 (N_17654,N_15675,N_15253);
nand U17655 (N_17655,N_14914,N_15393);
xnor U17656 (N_17656,N_15041,N_15034);
xor U17657 (N_17657,N_14272,N_15950);
or U17658 (N_17658,N_15381,N_15544);
xor U17659 (N_17659,N_15210,N_14599);
or U17660 (N_17660,N_14379,N_15716);
and U17661 (N_17661,N_15626,N_14360);
or U17662 (N_17662,N_14656,N_14417);
and U17663 (N_17663,N_15995,N_15211);
xnor U17664 (N_17664,N_14474,N_14408);
nand U17665 (N_17665,N_14782,N_15355);
or U17666 (N_17666,N_14349,N_14805);
nand U17667 (N_17667,N_14704,N_14290);
and U17668 (N_17668,N_14529,N_14463);
xor U17669 (N_17669,N_14449,N_14982);
nand U17670 (N_17670,N_14201,N_14566);
nor U17671 (N_17671,N_15877,N_15725);
nor U17672 (N_17672,N_15368,N_15512);
xor U17673 (N_17673,N_15513,N_15608);
nor U17674 (N_17674,N_14095,N_15374);
and U17675 (N_17675,N_14023,N_15666);
nor U17676 (N_17676,N_14213,N_15752);
xor U17677 (N_17677,N_15718,N_14126);
or U17678 (N_17678,N_14880,N_15327);
nand U17679 (N_17679,N_14817,N_14301);
nand U17680 (N_17680,N_15049,N_14121);
or U17681 (N_17681,N_15559,N_14477);
and U17682 (N_17682,N_15397,N_14112);
nor U17683 (N_17683,N_14080,N_14536);
xnor U17684 (N_17684,N_15443,N_14452);
nor U17685 (N_17685,N_15786,N_15233);
and U17686 (N_17686,N_15734,N_15374);
nand U17687 (N_17687,N_15390,N_14452);
nand U17688 (N_17688,N_15936,N_14435);
xnor U17689 (N_17689,N_14492,N_14306);
nand U17690 (N_17690,N_15334,N_15974);
nor U17691 (N_17691,N_15339,N_14748);
or U17692 (N_17692,N_15049,N_14022);
nand U17693 (N_17693,N_15101,N_15218);
nor U17694 (N_17694,N_14461,N_14459);
nor U17695 (N_17695,N_14379,N_15486);
xnor U17696 (N_17696,N_15631,N_14913);
nor U17697 (N_17697,N_14744,N_15811);
xor U17698 (N_17698,N_15449,N_14265);
nor U17699 (N_17699,N_15576,N_14310);
nand U17700 (N_17700,N_14633,N_14421);
nand U17701 (N_17701,N_15140,N_14924);
or U17702 (N_17702,N_14988,N_14017);
xor U17703 (N_17703,N_15971,N_14908);
nor U17704 (N_17704,N_15360,N_15334);
nand U17705 (N_17705,N_14290,N_14732);
or U17706 (N_17706,N_15243,N_14914);
nand U17707 (N_17707,N_15905,N_15918);
and U17708 (N_17708,N_14006,N_15148);
nand U17709 (N_17709,N_14224,N_15383);
nand U17710 (N_17710,N_15132,N_14839);
xnor U17711 (N_17711,N_14300,N_15528);
nand U17712 (N_17712,N_15630,N_15442);
nor U17713 (N_17713,N_15602,N_14489);
and U17714 (N_17714,N_15622,N_14172);
or U17715 (N_17715,N_15544,N_14593);
nor U17716 (N_17716,N_15744,N_15112);
xnor U17717 (N_17717,N_14354,N_14674);
or U17718 (N_17718,N_14629,N_15520);
nor U17719 (N_17719,N_15586,N_15309);
xor U17720 (N_17720,N_15162,N_15816);
xor U17721 (N_17721,N_14093,N_14418);
nand U17722 (N_17722,N_15179,N_15998);
or U17723 (N_17723,N_14582,N_15537);
nor U17724 (N_17724,N_14944,N_14588);
and U17725 (N_17725,N_14014,N_15319);
or U17726 (N_17726,N_15027,N_15295);
and U17727 (N_17727,N_15774,N_15587);
or U17728 (N_17728,N_14894,N_14360);
nand U17729 (N_17729,N_15085,N_15730);
nor U17730 (N_17730,N_14648,N_14435);
xnor U17731 (N_17731,N_15258,N_15246);
nand U17732 (N_17732,N_14776,N_14208);
xor U17733 (N_17733,N_14438,N_15187);
xnor U17734 (N_17734,N_14291,N_15165);
xnor U17735 (N_17735,N_15465,N_14922);
nor U17736 (N_17736,N_14443,N_15026);
xor U17737 (N_17737,N_15318,N_15534);
xor U17738 (N_17738,N_15631,N_14255);
and U17739 (N_17739,N_15772,N_15662);
nand U17740 (N_17740,N_15733,N_14079);
or U17741 (N_17741,N_14831,N_14576);
xnor U17742 (N_17742,N_15698,N_15790);
or U17743 (N_17743,N_14904,N_14968);
and U17744 (N_17744,N_15434,N_14672);
and U17745 (N_17745,N_15116,N_14737);
or U17746 (N_17746,N_14634,N_14707);
nor U17747 (N_17747,N_14224,N_15420);
and U17748 (N_17748,N_15904,N_15502);
and U17749 (N_17749,N_15607,N_15814);
nor U17750 (N_17750,N_15881,N_14311);
nor U17751 (N_17751,N_15042,N_14464);
xnor U17752 (N_17752,N_14144,N_15669);
or U17753 (N_17753,N_14420,N_15634);
nand U17754 (N_17754,N_15755,N_14158);
and U17755 (N_17755,N_15461,N_14622);
nand U17756 (N_17756,N_15671,N_15864);
nor U17757 (N_17757,N_15118,N_15781);
nor U17758 (N_17758,N_15587,N_14259);
nor U17759 (N_17759,N_14088,N_14344);
or U17760 (N_17760,N_14173,N_14829);
xor U17761 (N_17761,N_15289,N_15803);
nor U17762 (N_17762,N_15151,N_15580);
or U17763 (N_17763,N_14582,N_14815);
nand U17764 (N_17764,N_15775,N_15554);
xor U17765 (N_17765,N_15095,N_14106);
and U17766 (N_17766,N_15894,N_14038);
or U17767 (N_17767,N_14365,N_15655);
xnor U17768 (N_17768,N_15490,N_14359);
and U17769 (N_17769,N_14983,N_14159);
or U17770 (N_17770,N_14282,N_14271);
or U17771 (N_17771,N_14107,N_14175);
nand U17772 (N_17772,N_15600,N_14106);
and U17773 (N_17773,N_15479,N_14816);
xnor U17774 (N_17774,N_14498,N_14148);
nor U17775 (N_17775,N_14204,N_15624);
or U17776 (N_17776,N_14787,N_14178);
nor U17777 (N_17777,N_14253,N_15583);
xor U17778 (N_17778,N_15270,N_14086);
nand U17779 (N_17779,N_15785,N_15478);
nor U17780 (N_17780,N_15777,N_14623);
and U17781 (N_17781,N_14511,N_15822);
xor U17782 (N_17782,N_15414,N_14869);
nand U17783 (N_17783,N_15180,N_14692);
nand U17784 (N_17784,N_14023,N_15488);
and U17785 (N_17785,N_15955,N_14316);
xnor U17786 (N_17786,N_15307,N_15559);
xor U17787 (N_17787,N_14966,N_14443);
xor U17788 (N_17788,N_14164,N_14193);
nand U17789 (N_17789,N_15406,N_15423);
and U17790 (N_17790,N_15945,N_15158);
xor U17791 (N_17791,N_14634,N_14868);
nor U17792 (N_17792,N_14946,N_14330);
xnor U17793 (N_17793,N_14995,N_15073);
nand U17794 (N_17794,N_15804,N_15743);
nand U17795 (N_17795,N_15457,N_15511);
nor U17796 (N_17796,N_14678,N_15934);
xnor U17797 (N_17797,N_15272,N_15832);
and U17798 (N_17798,N_14693,N_14657);
xnor U17799 (N_17799,N_14962,N_15273);
nor U17800 (N_17800,N_14834,N_15583);
and U17801 (N_17801,N_14980,N_15153);
or U17802 (N_17802,N_15907,N_15275);
nor U17803 (N_17803,N_15855,N_14244);
nor U17804 (N_17804,N_14607,N_14204);
and U17805 (N_17805,N_15272,N_14603);
and U17806 (N_17806,N_15344,N_15877);
or U17807 (N_17807,N_15457,N_14091);
or U17808 (N_17808,N_15770,N_15325);
xor U17809 (N_17809,N_14365,N_15651);
or U17810 (N_17810,N_15297,N_15937);
and U17811 (N_17811,N_14436,N_15889);
xor U17812 (N_17812,N_15756,N_15814);
and U17813 (N_17813,N_15563,N_15601);
and U17814 (N_17814,N_15853,N_15584);
nor U17815 (N_17815,N_14426,N_15782);
nand U17816 (N_17816,N_15098,N_14993);
nand U17817 (N_17817,N_14040,N_14305);
nor U17818 (N_17818,N_14052,N_14606);
nand U17819 (N_17819,N_15771,N_14434);
and U17820 (N_17820,N_14732,N_14788);
nor U17821 (N_17821,N_14717,N_14735);
xor U17822 (N_17822,N_15770,N_14383);
xnor U17823 (N_17823,N_14395,N_14693);
nand U17824 (N_17824,N_14738,N_14660);
and U17825 (N_17825,N_14662,N_15119);
or U17826 (N_17826,N_15366,N_14336);
nand U17827 (N_17827,N_15877,N_14996);
xor U17828 (N_17828,N_15581,N_14408);
xnor U17829 (N_17829,N_15341,N_15781);
and U17830 (N_17830,N_14071,N_15045);
nand U17831 (N_17831,N_14221,N_15622);
nand U17832 (N_17832,N_15054,N_15353);
and U17833 (N_17833,N_15361,N_15521);
or U17834 (N_17834,N_14793,N_14109);
or U17835 (N_17835,N_15593,N_15133);
xor U17836 (N_17836,N_14318,N_14312);
xnor U17837 (N_17837,N_15947,N_15028);
xor U17838 (N_17838,N_14046,N_15188);
or U17839 (N_17839,N_15836,N_14994);
and U17840 (N_17840,N_15680,N_15886);
xnor U17841 (N_17841,N_15673,N_15646);
or U17842 (N_17842,N_14547,N_14073);
nor U17843 (N_17843,N_14921,N_15369);
and U17844 (N_17844,N_15829,N_15941);
xnor U17845 (N_17845,N_14652,N_14681);
xor U17846 (N_17846,N_15496,N_14465);
nand U17847 (N_17847,N_15993,N_14283);
or U17848 (N_17848,N_15979,N_14690);
xor U17849 (N_17849,N_14173,N_15881);
nor U17850 (N_17850,N_14081,N_15218);
xor U17851 (N_17851,N_14841,N_15129);
and U17852 (N_17852,N_14162,N_15376);
nor U17853 (N_17853,N_15166,N_15777);
and U17854 (N_17854,N_14144,N_14365);
nand U17855 (N_17855,N_14406,N_15961);
and U17856 (N_17856,N_14120,N_15686);
nor U17857 (N_17857,N_15752,N_14182);
nand U17858 (N_17858,N_15731,N_15693);
xnor U17859 (N_17859,N_14568,N_14909);
xnor U17860 (N_17860,N_15959,N_15113);
or U17861 (N_17861,N_14053,N_14038);
or U17862 (N_17862,N_14967,N_15878);
or U17863 (N_17863,N_14764,N_15823);
xnor U17864 (N_17864,N_15132,N_15254);
nand U17865 (N_17865,N_15755,N_15462);
nand U17866 (N_17866,N_15155,N_14734);
xnor U17867 (N_17867,N_14524,N_15063);
nor U17868 (N_17868,N_15962,N_14923);
nand U17869 (N_17869,N_14637,N_14071);
xor U17870 (N_17870,N_15075,N_15658);
and U17871 (N_17871,N_15314,N_15407);
or U17872 (N_17872,N_15587,N_14631);
nor U17873 (N_17873,N_15989,N_15596);
nor U17874 (N_17874,N_15144,N_15618);
or U17875 (N_17875,N_14910,N_15979);
nor U17876 (N_17876,N_14759,N_15292);
or U17877 (N_17877,N_15041,N_15602);
xnor U17878 (N_17878,N_14393,N_14922);
or U17879 (N_17879,N_14125,N_15234);
xor U17880 (N_17880,N_14990,N_14296);
xnor U17881 (N_17881,N_15550,N_14499);
or U17882 (N_17882,N_14195,N_15728);
or U17883 (N_17883,N_14334,N_15738);
and U17884 (N_17884,N_14091,N_14610);
and U17885 (N_17885,N_14557,N_15911);
nor U17886 (N_17886,N_14574,N_15916);
nor U17887 (N_17887,N_15055,N_14589);
nor U17888 (N_17888,N_14548,N_14495);
nor U17889 (N_17889,N_14475,N_14883);
or U17890 (N_17890,N_15445,N_14042);
xor U17891 (N_17891,N_15052,N_15691);
nor U17892 (N_17892,N_15843,N_14404);
and U17893 (N_17893,N_15633,N_15908);
and U17894 (N_17894,N_14698,N_15711);
or U17895 (N_17895,N_14344,N_14747);
nand U17896 (N_17896,N_14474,N_15080);
nand U17897 (N_17897,N_15048,N_15282);
or U17898 (N_17898,N_15483,N_14054);
or U17899 (N_17899,N_14151,N_15266);
nand U17900 (N_17900,N_14162,N_15990);
nor U17901 (N_17901,N_14829,N_15372);
nand U17902 (N_17902,N_14675,N_15997);
nand U17903 (N_17903,N_14350,N_14962);
nand U17904 (N_17904,N_14565,N_14712);
and U17905 (N_17905,N_14819,N_14570);
or U17906 (N_17906,N_14597,N_14799);
nand U17907 (N_17907,N_14251,N_15966);
nor U17908 (N_17908,N_14609,N_15275);
or U17909 (N_17909,N_14145,N_14536);
nor U17910 (N_17910,N_15402,N_14796);
xnor U17911 (N_17911,N_14978,N_14451);
and U17912 (N_17912,N_14364,N_15845);
and U17913 (N_17913,N_14214,N_14122);
nor U17914 (N_17914,N_15467,N_14329);
or U17915 (N_17915,N_15584,N_14971);
nor U17916 (N_17916,N_14943,N_14324);
xor U17917 (N_17917,N_15488,N_15537);
and U17918 (N_17918,N_15957,N_14520);
or U17919 (N_17919,N_14689,N_15152);
nor U17920 (N_17920,N_15147,N_15214);
xor U17921 (N_17921,N_15455,N_14266);
nand U17922 (N_17922,N_15669,N_15450);
nand U17923 (N_17923,N_14973,N_14736);
nor U17924 (N_17924,N_14410,N_15159);
xor U17925 (N_17925,N_14688,N_14063);
nor U17926 (N_17926,N_15366,N_15035);
xor U17927 (N_17927,N_14641,N_15398);
and U17928 (N_17928,N_14059,N_14615);
or U17929 (N_17929,N_15255,N_14880);
or U17930 (N_17930,N_14431,N_14314);
xnor U17931 (N_17931,N_14513,N_15252);
xnor U17932 (N_17932,N_15796,N_15914);
and U17933 (N_17933,N_15607,N_14472);
nor U17934 (N_17934,N_14310,N_14589);
xor U17935 (N_17935,N_15213,N_14511);
and U17936 (N_17936,N_15687,N_14252);
and U17937 (N_17937,N_15342,N_14549);
and U17938 (N_17938,N_15171,N_15205);
and U17939 (N_17939,N_15604,N_15217);
nand U17940 (N_17940,N_14191,N_15586);
xor U17941 (N_17941,N_15904,N_14100);
xnor U17942 (N_17942,N_14831,N_14405);
nor U17943 (N_17943,N_15513,N_15866);
nand U17944 (N_17944,N_15401,N_14763);
and U17945 (N_17945,N_15626,N_15515);
nor U17946 (N_17946,N_14278,N_15564);
and U17947 (N_17947,N_14897,N_14110);
or U17948 (N_17948,N_15770,N_14568);
nand U17949 (N_17949,N_14182,N_14699);
nand U17950 (N_17950,N_14117,N_14144);
nor U17951 (N_17951,N_14587,N_14470);
or U17952 (N_17952,N_15100,N_15253);
and U17953 (N_17953,N_14409,N_14763);
and U17954 (N_17954,N_15816,N_14725);
xnor U17955 (N_17955,N_15419,N_15408);
or U17956 (N_17956,N_15476,N_14690);
or U17957 (N_17957,N_15681,N_15435);
xor U17958 (N_17958,N_14653,N_14852);
nand U17959 (N_17959,N_15015,N_14909);
and U17960 (N_17960,N_14202,N_15415);
xor U17961 (N_17961,N_15661,N_14433);
nor U17962 (N_17962,N_15112,N_14877);
xor U17963 (N_17963,N_15161,N_14482);
nor U17964 (N_17964,N_14819,N_15494);
nor U17965 (N_17965,N_15353,N_14984);
nor U17966 (N_17966,N_15540,N_15467);
nor U17967 (N_17967,N_14175,N_14718);
or U17968 (N_17968,N_14571,N_15176);
xnor U17969 (N_17969,N_14109,N_15960);
xnor U17970 (N_17970,N_15494,N_14926);
or U17971 (N_17971,N_15835,N_14169);
nand U17972 (N_17972,N_15860,N_15231);
nor U17973 (N_17973,N_15359,N_15450);
nand U17974 (N_17974,N_14362,N_14294);
nor U17975 (N_17975,N_15499,N_15530);
and U17976 (N_17976,N_14816,N_15529);
or U17977 (N_17977,N_14826,N_15759);
nand U17978 (N_17978,N_14696,N_15872);
nand U17979 (N_17979,N_15027,N_14927);
nor U17980 (N_17980,N_14760,N_15962);
or U17981 (N_17981,N_14086,N_14337);
nor U17982 (N_17982,N_15349,N_15080);
nor U17983 (N_17983,N_15130,N_15815);
nor U17984 (N_17984,N_15250,N_14430);
and U17985 (N_17985,N_15622,N_14364);
and U17986 (N_17986,N_14583,N_14325);
and U17987 (N_17987,N_15922,N_15085);
xor U17988 (N_17988,N_15525,N_14667);
xor U17989 (N_17989,N_15789,N_15346);
and U17990 (N_17990,N_15055,N_15881);
and U17991 (N_17991,N_14785,N_14941);
or U17992 (N_17992,N_14174,N_14575);
nand U17993 (N_17993,N_14901,N_14004);
nand U17994 (N_17994,N_14767,N_14891);
nand U17995 (N_17995,N_15102,N_15674);
or U17996 (N_17996,N_14264,N_14917);
or U17997 (N_17997,N_14766,N_15367);
nor U17998 (N_17998,N_15595,N_14621);
nor U17999 (N_17999,N_14419,N_15348);
nand U18000 (N_18000,N_17634,N_17311);
xor U18001 (N_18001,N_16008,N_17074);
and U18002 (N_18002,N_16402,N_16853);
or U18003 (N_18003,N_17374,N_17265);
nand U18004 (N_18004,N_16208,N_17336);
xor U18005 (N_18005,N_16078,N_17671);
xor U18006 (N_18006,N_16443,N_17240);
or U18007 (N_18007,N_16495,N_17703);
nand U18008 (N_18008,N_17011,N_16704);
or U18009 (N_18009,N_17591,N_16745);
xnor U18010 (N_18010,N_17224,N_17155);
or U18011 (N_18011,N_17093,N_17307);
or U18012 (N_18012,N_16445,N_16293);
or U18013 (N_18013,N_17954,N_17613);
and U18014 (N_18014,N_17053,N_16786);
or U18015 (N_18015,N_16081,N_17501);
nor U18016 (N_18016,N_16496,N_17745);
xnor U18017 (N_18017,N_17179,N_16720);
or U18018 (N_18018,N_16998,N_17459);
and U18019 (N_18019,N_17712,N_16325);
or U18020 (N_18020,N_17489,N_16071);
nor U18021 (N_18021,N_17231,N_17604);
and U18022 (N_18022,N_16881,N_17857);
and U18023 (N_18023,N_16089,N_16501);
or U18024 (N_18024,N_17095,N_16905);
xor U18025 (N_18025,N_17827,N_17452);
nand U18026 (N_18026,N_16876,N_16957);
nor U18027 (N_18027,N_17366,N_16614);
or U18028 (N_18028,N_17960,N_17235);
xnor U18029 (N_18029,N_16085,N_17792);
or U18030 (N_18030,N_16392,N_16479);
nand U18031 (N_18031,N_16234,N_17414);
or U18032 (N_18032,N_16269,N_17565);
and U18033 (N_18033,N_17953,N_16301);
nand U18034 (N_18034,N_17503,N_17525);
or U18035 (N_18035,N_17124,N_17207);
xor U18036 (N_18036,N_16139,N_16152);
xnor U18037 (N_18037,N_17025,N_16473);
nor U18038 (N_18038,N_16682,N_16251);
or U18039 (N_18039,N_17123,N_17623);
nand U18040 (N_18040,N_16581,N_17728);
nand U18041 (N_18041,N_17079,N_17014);
or U18042 (N_18042,N_16137,N_17068);
or U18043 (N_18043,N_17361,N_16757);
or U18044 (N_18044,N_16449,N_16116);
nor U18045 (N_18045,N_16361,N_16332);
and U18046 (N_18046,N_17154,N_16554);
nand U18047 (N_18047,N_16342,N_16742);
nand U18048 (N_18048,N_17873,N_16994);
nor U18049 (N_18049,N_17210,N_17164);
and U18050 (N_18050,N_17814,N_17756);
or U18051 (N_18051,N_17127,N_16611);
nand U18052 (N_18052,N_17335,N_17901);
or U18053 (N_18053,N_17135,N_17602);
nor U18054 (N_18054,N_17196,N_17746);
xor U18055 (N_18055,N_17077,N_17139);
and U18056 (N_18056,N_16435,N_16290);
nand U18057 (N_18057,N_16926,N_16803);
nand U18058 (N_18058,N_16668,N_16934);
and U18059 (N_18059,N_16558,N_17449);
xnor U18060 (N_18060,N_16337,N_17642);
nor U18061 (N_18061,N_16698,N_17805);
nand U18062 (N_18062,N_16799,N_16056);
xor U18063 (N_18063,N_17845,N_16255);
and U18064 (N_18064,N_17568,N_16945);
and U18065 (N_18065,N_17800,N_17580);
nand U18066 (N_18066,N_17151,N_16442);
xnor U18067 (N_18067,N_16930,N_17447);
xnor U18068 (N_18068,N_16741,N_16666);
nand U18069 (N_18069,N_16002,N_16621);
nand U18070 (N_18070,N_16419,N_16055);
nand U18071 (N_18071,N_16266,N_17573);
and U18072 (N_18072,N_16047,N_16919);
xor U18073 (N_18073,N_17474,N_16220);
xnor U18074 (N_18074,N_16430,N_17888);
and U18075 (N_18075,N_16936,N_17847);
nor U18076 (N_18076,N_17719,N_16235);
nor U18077 (N_18077,N_17698,N_16223);
nand U18078 (N_18078,N_16578,N_16816);
or U18079 (N_18079,N_17665,N_17567);
xnor U18080 (N_18080,N_16535,N_17523);
and U18081 (N_18081,N_17092,N_16005);
or U18082 (N_18082,N_16670,N_16846);
or U18083 (N_18083,N_17789,N_17770);
or U18084 (N_18084,N_17026,N_17056);
nor U18085 (N_18085,N_16871,N_16677);
and U18086 (N_18086,N_16317,N_17247);
or U18087 (N_18087,N_17578,N_16333);
nor U18088 (N_18088,N_17003,N_17650);
and U18089 (N_18089,N_16952,N_16190);
or U18090 (N_18090,N_17484,N_17941);
nand U18091 (N_18091,N_17669,N_16972);
nand U18092 (N_18092,N_16692,N_17097);
nand U18093 (N_18093,N_17028,N_17391);
or U18094 (N_18094,N_17212,N_16583);
xor U18095 (N_18095,N_17007,N_17933);
nor U18096 (N_18096,N_17148,N_17664);
or U18097 (N_18097,N_16792,N_16789);
nand U18098 (N_18098,N_17463,N_16397);
or U18099 (N_18099,N_16010,N_16405);
nand U18100 (N_18100,N_16570,N_17673);
nor U18101 (N_18101,N_17475,N_17152);
nor U18102 (N_18102,N_16159,N_16236);
nor U18103 (N_18103,N_16519,N_17736);
or U18104 (N_18104,N_17334,N_16077);
nand U18105 (N_18105,N_17248,N_17275);
xnor U18106 (N_18106,N_17040,N_17004);
nor U18107 (N_18107,N_16557,N_17396);
or U18108 (N_18108,N_17258,N_16748);
xnor U18109 (N_18109,N_16591,N_16689);
nand U18110 (N_18110,N_16347,N_16633);
and U18111 (N_18111,N_16831,N_16962);
nand U18112 (N_18112,N_17246,N_17588);
or U18113 (N_18113,N_16469,N_16609);
and U18114 (N_18114,N_16695,N_16316);
and U18115 (N_18115,N_17538,N_17510);
or U18116 (N_18116,N_17957,N_16801);
nand U18117 (N_18117,N_17683,N_16123);
xor U18118 (N_18118,N_16487,N_17296);
or U18119 (N_18119,N_17773,N_17967);
or U18120 (N_18120,N_16475,N_17601);
nand U18121 (N_18121,N_16192,N_17462);
and U18122 (N_18122,N_16737,N_17812);
and U18123 (N_18123,N_16630,N_16599);
or U18124 (N_18124,N_16140,N_16894);
nand U18125 (N_18125,N_17997,N_16640);
nor U18126 (N_18126,N_16088,N_16303);
or U18127 (N_18127,N_17401,N_17036);
xor U18128 (N_18128,N_17104,N_16768);
xnor U18129 (N_18129,N_16855,N_16766);
and U18130 (N_18130,N_16702,N_16477);
nand U18131 (N_18131,N_16713,N_17754);
or U18132 (N_18132,N_16587,N_17570);
nor U18133 (N_18133,N_16451,N_17122);
and U18134 (N_18134,N_17279,N_17998);
nor U18135 (N_18135,N_16204,N_16369);
xor U18136 (N_18136,N_16462,N_16354);
nor U18137 (N_18137,N_16341,N_17631);
or U18138 (N_18138,N_17558,N_17149);
nand U18139 (N_18139,N_17498,N_17750);
nor U18140 (N_18140,N_16328,N_16087);
nand U18141 (N_18141,N_16358,N_17765);
and U18142 (N_18142,N_17267,N_16901);
or U18143 (N_18143,N_17211,N_17821);
and U18144 (N_18144,N_17958,N_17522);
nand U18145 (N_18145,N_17255,N_16020);
xor U18146 (N_18146,N_17426,N_16539);
nor U18147 (N_18147,N_16153,N_17595);
xor U18148 (N_18148,N_16463,N_17915);
or U18149 (N_18149,N_17017,N_17706);
nor U18150 (N_18150,N_16113,N_16749);
nand U18151 (N_18151,N_17860,N_16458);
xnor U18152 (N_18152,N_17238,N_16434);
nor U18153 (N_18153,N_17696,N_16067);
and U18154 (N_18154,N_17778,N_16909);
or U18155 (N_18155,N_16016,N_17944);
xnor U18156 (N_18156,N_17536,N_17024);
nand U18157 (N_18157,N_16158,N_17174);
nand U18158 (N_18158,N_16559,N_17397);
or U18159 (N_18159,N_17759,N_16657);
nor U18160 (N_18160,N_16108,N_16194);
or U18161 (N_18161,N_16176,N_16650);
and U18162 (N_18162,N_16149,N_17194);
nor U18163 (N_18163,N_17083,N_16572);
xor U18164 (N_18164,N_17514,N_16438);
nand U18165 (N_18165,N_17672,N_17136);
or U18166 (N_18166,N_16517,N_17315);
or U18167 (N_18167,N_16605,N_16944);
nand U18168 (N_18168,N_16980,N_16798);
and U18169 (N_18169,N_17477,N_17994);
or U18170 (N_18170,N_17911,N_16017);
nor U18171 (N_18171,N_16925,N_16610);
nand U18172 (N_18172,N_16765,N_17084);
or U18173 (N_18173,N_16384,N_16672);
nor U18174 (N_18174,N_17422,N_16750);
nand U18175 (N_18175,N_16117,N_16838);
nand U18176 (N_18176,N_17547,N_17768);
and U18177 (N_18177,N_17724,N_16093);
nor U18178 (N_18178,N_16995,N_16270);
nor U18179 (N_18179,N_17629,N_17362);
nor U18180 (N_18180,N_17098,N_16996);
nor U18181 (N_18181,N_17897,N_17395);
and U18182 (N_18182,N_17882,N_16125);
or U18183 (N_18183,N_17368,N_17242);
and U18184 (N_18184,N_16439,N_17909);
nand U18185 (N_18185,N_16004,N_16773);
xnor U18186 (N_18186,N_17892,N_16310);
nand U18187 (N_18187,N_17013,N_17912);
nor U18188 (N_18188,N_16225,N_17418);
and U18189 (N_18189,N_16910,N_17150);
or U18190 (N_18190,N_16965,N_17569);
xor U18191 (N_18191,N_17991,N_16858);
nor U18192 (N_18192,N_17332,N_16180);
and U18193 (N_18193,N_16634,N_16009);
xnor U18194 (N_18194,N_16506,N_17886);
and U18195 (N_18195,N_17561,N_16186);
or U18196 (N_18196,N_16191,N_17229);
xor U18197 (N_18197,N_16025,N_17303);
xnor U18198 (N_18198,N_17572,N_16026);
and U18199 (N_18199,N_17584,N_16437);
xor U18200 (N_18200,N_17293,N_16282);
xor U18201 (N_18201,N_16883,N_17468);
and U18202 (N_18202,N_16331,N_17114);
and U18203 (N_18203,N_17078,N_17627);
nand U18204 (N_18204,N_16367,N_17813);
nor U18205 (N_18205,N_17282,N_17505);
nor U18206 (N_18206,N_16814,N_17281);
or U18207 (N_18207,N_17290,N_16507);
or U18208 (N_18208,N_17730,N_17801);
and U18209 (N_18209,N_16121,N_16997);
and U18210 (N_18210,N_17497,N_17437);
nand U18211 (N_18211,N_16807,N_17980);
nand U18212 (N_18212,N_17617,N_17316);
xnor U18213 (N_18213,N_16033,N_17541);
nor U18214 (N_18214,N_16759,N_17337);
nand U18215 (N_18215,N_16850,N_16619);
and U18216 (N_18216,N_17284,N_17702);
nand U18217 (N_18217,N_16400,N_16642);
or U18218 (N_18218,N_16529,N_17715);
nand U18219 (N_18219,N_16351,N_17320);
xor U18220 (N_18220,N_17389,N_17520);
and U18221 (N_18221,N_17478,N_17137);
nand U18222 (N_18222,N_17379,N_16497);
xnor U18223 (N_18223,N_16508,N_16527);
xnor U18224 (N_18224,N_16064,N_16521);
and U18225 (N_18225,N_17461,N_17701);
or U18226 (N_18226,N_16963,N_16305);
or U18227 (N_18227,N_16373,N_16848);
nand U18228 (N_18228,N_17039,N_17767);
nand U18229 (N_18229,N_17637,N_17470);
and U18230 (N_18230,N_16021,N_16385);
or U18231 (N_18231,N_17542,N_16143);
nand U18232 (N_18232,N_16329,N_17632);
xor U18233 (N_18233,N_17609,N_16012);
or U18234 (N_18234,N_17167,N_16170);
xnor U18235 (N_18235,N_16688,N_16623);
xor U18236 (N_18236,N_17908,N_16567);
nand U18237 (N_18237,N_17775,N_16511);
nand U18238 (N_18238,N_16870,N_16075);
or U18239 (N_18239,N_16074,N_16415);
nor U18240 (N_18240,N_16062,N_16272);
and U18241 (N_18241,N_17041,N_16107);
and U18242 (N_18242,N_16218,N_16694);
nor U18243 (N_18243,N_16168,N_16514);
and U18244 (N_18244,N_17030,N_17914);
xnor U18245 (N_18245,N_17180,N_17118);
or U18246 (N_18246,N_17657,N_17199);
nor U18247 (N_18247,N_16857,N_17670);
nor U18248 (N_18248,N_16904,N_16806);
nor U18249 (N_18249,N_16835,N_16700);
or U18250 (N_18250,N_16345,N_16526);
or U18251 (N_18251,N_17818,N_17057);
nor U18252 (N_18252,N_16724,N_17987);
xnor U18253 (N_18253,N_17791,N_17681);
nor U18254 (N_18254,N_16933,N_16491);
nor U18255 (N_18255,N_16092,N_16863);
and U18256 (N_18256,N_16110,N_16822);
or U18257 (N_18257,N_17215,N_17896);
nand U18258 (N_18258,N_16481,N_16073);
nand U18259 (N_18259,N_16263,N_17063);
nand U18260 (N_18260,N_17716,N_17688);
nand U18261 (N_18261,N_17250,N_17469);
xnor U18262 (N_18262,N_16907,N_16461);
and U18263 (N_18263,N_17015,N_16032);
nand U18264 (N_18264,N_16524,N_16566);
nor U18265 (N_18265,N_16388,N_16631);
and U18266 (N_18266,N_16243,N_17298);
nand U18267 (N_18267,N_16346,N_16947);
xnor U18268 (N_18268,N_16311,N_17407);
nor U18269 (N_18269,N_16141,N_17974);
nand U18270 (N_18270,N_17722,N_16543);
or U18271 (N_18271,N_16752,N_17817);
and U18272 (N_18272,N_17667,N_16146);
or U18273 (N_18273,N_17370,N_17710);
or U18274 (N_18274,N_16761,N_16277);
xor U18275 (N_18275,N_17863,N_16289);
nor U18276 (N_18276,N_16841,N_17300);
xnor U18277 (N_18277,N_17556,N_17738);
or U18278 (N_18278,N_17012,N_16364);
nand U18279 (N_18279,N_17988,N_17492);
nand U18280 (N_18280,N_17921,N_17594);
xnor U18281 (N_18281,N_16776,N_17090);
nor U18282 (N_18282,N_16523,N_16828);
nor U18283 (N_18283,N_17338,N_16880);
or U18284 (N_18284,N_17844,N_16760);
xor U18285 (N_18285,N_17810,N_16536);
and U18286 (N_18286,N_17831,N_17192);
and U18287 (N_18287,N_16097,N_16826);
nand U18288 (N_18288,N_17985,N_16129);
nor U18289 (N_18289,N_17061,N_17635);
xnor U18290 (N_18290,N_16315,N_16183);
and U18291 (N_18291,N_16472,N_16426);
xor U18292 (N_18292,N_17984,N_16375);
xnor U18293 (N_18293,N_17540,N_17209);
xor U18294 (N_18294,N_17564,N_17159);
nand U18295 (N_18295,N_16410,N_16249);
or U18296 (N_18296,N_16770,N_17947);
nor U18297 (N_18297,N_16549,N_17979);
nor U18298 (N_18298,N_17128,N_17718);
nand U18299 (N_18299,N_17927,N_16932);
nor U18300 (N_18300,N_17530,N_16716);
and U18301 (N_18301,N_17254,N_16057);
nor U18302 (N_18302,N_16649,N_16890);
nor U18303 (N_18303,N_16307,N_17867);
xnor U18304 (N_18304,N_16979,N_17589);
nor U18305 (N_18305,N_17108,N_17431);
nor U18306 (N_18306,N_16321,N_16987);
nand U18307 (N_18307,N_16959,N_16112);
nor U18308 (N_18308,N_16457,N_16573);
nor U18309 (N_18309,N_17112,N_16124);
nor U18310 (N_18310,N_17067,N_16164);
nand U18311 (N_18311,N_17741,N_16476);
and U18312 (N_18312,N_17910,N_16120);
nand U18313 (N_18313,N_16780,N_17643);
nor U18314 (N_18314,N_16271,N_17232);
xor U18315 (N_18315,N_17619,N_17100);
nand U18316 (N_18316,N_16733,N_16387);
nand U18317 (N_18317,N_17377,N_17292);
and U18318 (N_18318,N_17203,N_17417);
and U18319 (N_18319,N_17913,N_16040);
and U18320 (N_18320,N_16478,N_16774);
or U18321 (N_18321,N_16132,N_17404);
xor U18322 (N_18322,N_16136,N_16096);
or U18323 (N_18323,N_16804,N_16372);
and U18324 (N_18324,N_17782,N_17271);
or U18325 (N_18325,N_16825,N_17195);
xor U18326 (N_18326,N_16399,N_17113);
and U18327 (N_18327,N_16753,N_16635);
nor U18328 (N_18328,N_16992,N_17824);
and U18329 (N_18329,N_16050,N_16882);
nand U18330 (N_18330,N_17156,N_17239);
nor U18331 (N_18331,N_16955,N_16340);
xor U18332 (N_18332,N_16663,N_17900);
xor U18333 (N_18333,N_16178,N_16797);
nand U18334 (N_18334,N_16576,N_17644);
nor U18335 (N_18335,N_16195,N_17763);
and U18336 (N_18336,N_16823,N_17218);
nor U18337 (N_18337,N_17605,N_16349);
and U18338 (N_18338,N_16296,N_17309);
nand U18339 (N_18339,N_16624,N_17950);
nand U18340 (N_18340,N_17021,N_17828);
and U18341 (N_18341,N_17811,N_17555);
and U18342 (N_18342,N_17682,N_16179);
and U18343 (N_18343,N_17432,N_17064);
xnor U18344 (N_18344,N_17717,N_16242);
or U18345 (N_18345,N_17943,N_17858);
nor U18346 (N_18346,N_16382,N_16974);
nor U18347 (N_18347,N_17226,N_17852);
nor U18348 (N_18348,N_16468,N_16589);
or U18349 (N_18349,N_17052,N_16532);
xnor U18350 (N_18350,N_17472,N_16466);
or U18351 (N_18351,N_16363,N_17663);
xnor U18352 (N_18352,N_17270,N_17380);
nand U18353 (N_18353,N_16412,N_16515);
xnor U18354 (N_18354,N_16128,N_17324);
and U18355 (N_18355,N_17109,N_16245);
xor U18356 (N_18356,N_16313,N_17798);
and U18357 (N_18357,N_17721,N_16082);
or U18358 (N_18358,N_16708,N_16887);
nor U18359 (N_18359,N_17725,N_17096);
and U18360 (N_18360,N_17088,N_16083);
or U18361 (N_18361,N_17173,N_17935);
and U18362 (N_18362,N_16893,N_17513);
nand U18363 (N_18363,N_17333,N_16066);
xor U18364 (N_18364,N_16498,N_17575);
or U18365 (N_18365,N_17557,N_17005);
nand U18366 (N_18366,N_16456,N_17420);
nor U18367 (N_18367,N_17170,N_16394);
xnor U18368 (N_18368,N_17582,N_16884);
nand U18369 (N_18369,N_16027,N_17883);
or U18370 (N_18370,N_17952,N_17214);
or U18371 (N_18371,N_17051,N_17859);
and U18372 (N_18372,N_16983,N_16134);
nor U18373 (N_18373,N_17115,N_17286);
nand U18374 (N_18374,N_17185,N_16416);
nor U18375 (N_18375,N_16685,N_16203);
and U18376 (N_18376,N_17949,N_17652);
xnor U18377 (N_18377,N_16182,N_17964);
xnor U18378 (N_18378,N_17168,N_16480);
or U18379 (N_18379,N_16028,N_17802);
xnor U18380 (N_18380,N_17393,N_17237);
nand U18381 (N_18381,N_17382,N_16683);
nor U18382 (N_18382,N_16673,N_17408);
nand U18383 (N_18383,N_16785,N_16811);
nor U18384 (N_18384,N_17799,N_16209);
and U18385 (N_18385,N_17851,N_17651);
or U18386 (N_18386,N_17329,N_16034);
nor U18387 (N_18387,N_17260,N_17976);
nand U18388 (N_18388,N_17948,N_17043);
nand U18389 (N_18389,N_17826,N_16546);
nor U18390 (N_18390,N_16701,N_17607);
and U18391 (N_18391,N_16157,N_16058);
and U18392 (N_18392,N_17073,N_16793);
and U18393 (N_18393,N_17638,N_17055);
xnor U18394 (N_18394,N_17321,N_17516);
or U18395 (N_18395,N_16199,N_17328);
nand U18396 (N_18396,N_16122,N_16678);
nor U18397 (N_18397,N_16181,N_17111);
nand U18398 (N_18398,N_17630,N_17546);
nor U18399 (N_18399,N_16184,N_16420);
and U18400 (N_18400,N_16898,N_16035);
and U18401 (N_18401,N_17989,N_17848);
nand U18402 (N_18402,N_16403,N_16258);
nand U18403 (N_18403,N_16632,N_16739);
nand U18404 (N_18404,N_16031,N_17448);
nor U18405 (N_18405,N_16731,N_16404);
or U18406 (N_18406,N_17121,N_17781);
and U18407 (N_18407,N_16395,N_17843);
and U18408 (N_18408,N_16928,N_17415);
nor U18409 (N_18409,N_17839,N_17225);
or U18410 (N_18410,N_17116,N_16975);
xor U18411 (N_18411,N_17714,N_16764);
nand U18412 (N_18412,N_16503,N_16743);
nand U18413 (N_18413,N_17543,N_16101);
nand U18414 (N_18414,N_16794,N_17624);
xnor U18415 (N_18415,N_17243,N_16784);
nand U18416 (N_18416,N_17126,N_17739);
xnor U18417 (N_18417,N_17842,N_17598);
nand U18418 (N_18418,N_17069,N_16844);
and U18419 (N_18419,N_17940,N_16460);
or U18420 (N_18420,N_16655,N_17434);
nor U18421 (N_18421,N_16571,N_17198);
xor U18422 (N_18422,N_17257,N_17268);
nor U18423 (N_18423,N_17027,N_16726);
nor U18424 (N_18424,N_16467,N_17744);
nor U18425 (N_18425,N_17752,N_16641);
or U18426 (N_18426,N_17502,N_17455);
or U18427 (N_18427,N_16989,N_17038);
xor U18428 (N_18428,N_17628,N_17878);
nor U18429 (N_18429,N_16569,N_17369);
xor U18430 (N_18430,N_17454,N_17228);
or U18431 (N_18431,N_16492,N_16448);
or U18432 (N_18432,N_16528,N_16275);
xor U18433 (N_18433,N_16795,N_17453);
nor U18434 (N_18434,N_17599,N_16039);
nand U18435 (N_18435,N_17691,N_16232);
or U18436 (N_18436,N_16604,N_17481);
or U18437 (N_18437,N_17022,N_16915);
and U18438 (N_18438,N_17733,N_16485);
or U18439 (N_18439,N_17587,N_16086);
and U18440 (N_18440,N_17936,N_17992);
nor U18441 (N_18441,N_16348,N_17533);
nor U18442 (N_18442,N_17134,N_16665);
or U18443 (N_18443,N_16019,N_16982);
xor U18444 (N_18444,N_16046,N_16555);
nand U18445 (N_18445,N_16411,N_16206);
xnor U18446 (N_18446,N_17836,N_16585);
and U18447 (N_18447,N_17085,N_17266);
or U18448 (N_18448,N_17512,N_16431);
or U18449 (N_18449,N_17485,N_16261);
and U18450 (N_18450,N_17029,N_16590);
xor U18451 (N_18451,N_17807,N_17458);
nand U18452 (N_18452,N_16114,N_16284);
and U18453 (N_18453,N_16849,N_16579);
xor U18454 (N_18454,N_17346,N_17054);
and U18455 (N_18455,N_16586,N_17165);
nor U18456 (N_18456,N_17310,N_16993);
or U18457 (N_18457,N_17131,N_16868);
xnor U18458 (N_18458,N_17425,N_17956);
xor U18459 (N_18459,N_16072,N_16043);
or U18460 (N_18460,N_16544,N_17072);
nor U18461 (N_18461,N_17130,N_16376);
and U18462 (N_18462,N_17592,N_16727);
and U18463 (N_18463,N_16254,N_17059);
xor U18464 (N_18464,N_16600,N_17586);
xor U18465 (N_18465,N_17668,N_16864);
nand U18466 (N_18466,N_17327,N_17189);
nor U18467 (N_18467,N_16187,N_16628);
or U18468 (N_18468,N_17600,N_16253);
nor U18469 (N_18469,N_16295,N_17330);
xor U18470 (N_18470,N_16484,N_16493);
xor U18471 (N_18471,N_17045,N_17313);
nand U18472 (N_18472,N_17143,N_17413);
or U18473 (N_18473,N_17995,N_16903);
nor U18474 (N_18474,N_17687,N_16705);
or U18475 (N_18475,N_17815,N_16440);
and U18476 (N_18476,N_16059,N_17274);
nand U18477 (N_18477,N_16777,N_17879);
and U18478 (N_18478,N_17089,N_17436);
nor U18479 (N_18479,N_16219,N_17119);
nand U18480 (N_18480,N_16175,N_16732);
xor U18481 (N_18481,N_17732,N_17511);
nor U18482 (N_18482,N_16030,N_16118);
nor U18483 (N_18483,N_17375,N_17507);
and U18484 (N_18484,N_16297,N_17087);
nor U18485 (N_18485,N_17438,N_16730);
and U18486 (N_18486,N_16091,N_16895);
and U18487 (N_18487,N_16450,N_17190);
and U18488 (N_18488,N_16336,N_17476);
and U18489 (N_18489,N_17806,N_17480);
and U18490 (N_18490,N_17264,N_16740);
or U18491 (N_18491,N_16725,N_16424);
nand U18492 (N_18492,N_17008,N_16264);
nor U18493 (N_18493,N_17145,N_16827);
and U18494 (N_18494,N_16309,N_17363);
nor U18495 (N_18495,N_17709,N_17539);
or U18496 (N_18496,N_16189,N_17625);
nand U18497 (N_18497,N_16279,N_17982);
nor U18498 (N_18498,N_16565,N_17986);
and U18499 (N_18499,N_17521,N_17220);
nor U18500 (N_18500,N_16499,N_16425);
xor U18501 (N_18501,N_17550,N_16818);
nand U18502 (N_18502,N_16418,N_16001);
or U18503 (N_18503,N_16287,N_16343);
nor U18504 (N_18504,N_17753,N_17419);
nand U18505 (N_18505,N_16645,N_17349);
or U18506 (N_18506,N_17659,N_16106);
nor U18507 (N_18507,N_17343,N_16875);
and U18508 (N_18508,N_16984,N_17340);
and U18509 (N_18509,N_17387,N_17094);
and U18510 (N_18510,N_17693,N_16080);
xnor U18511 (N_18511,N_16935,N_16892);
and U18512 (N_18512,N_16659,N_17433);
nor U18513 (N_18513,N_17776,N_17531);
and U18514 (N_18514,N_16252,N_16697);
nor U18515 (N_18515,N_16652,N_17383);
nor U18516 (N_18516,N_17518,N_16154);
nor U18517 (N_18517,N_16562,N_16281);
or U18518 (N_18518,N_17790,N_17705);
nand U18519 (N_18519,N_17450,N_16699);
and U18520 (N_18520,N_16422,N_16474);
and U18521 (N_18521,N_16246,N_17708);
xnor U18522 (N_18522,N_17653,N_16548);
nand U18523 (N_18523,N_16888,N_16432);
nor U18524 (N_18524,N_17972,N_17169);
or U18525 (N_18525,N_17692,N_17922);
and U18526 (N_18526,N_16537,N_16629);
and U18527 (N_18527,N_17576,N_16015);
and U18528 (N_18528,N_17748,N_16862);
nor U18529 (N_18529,N_17889,N_17062);
and U18530 (N_18530,N_16833,N_16217);
nand U18531 (N_18531,N_17158,N_17585);
nor U18532 (N_18532,N_16891,N_17144);
nor U18533 (N_18533,N_17352,N_17685);
or U18534 (N_18534,N_16755,N_17376);
or U18535 (N_18535,N_17784,N_17399);
or U18536 (N_18536,N_17545,N_17772);
xor U18537 (N_18537,N_17552,N_16126);
nand U18538 (N_18538,N_17978,N_17506);
nand U18539 (N_18539,N_16094,N_16148);
nor U18540 (N_18540,N_16355,N_16593);
xor U18541 (N_18541,N_17285,N_17755);
and U18542 (N_18542,N_17217,N_17785);
nor U18543 (N_18543,N_17101,N_17891);
nor U18544 (N_18544,N_16049,N_17559);
nand U18545 (N_18545,N_16886,N_16772);
and U18546 (N_18546,N_17299,N_17367);
nand U18547 (N_18547,N_17661,N_16455);
or U18548 (N_18548,N_16371,N_17381);
nor U18549 (N_18549,N_16398,N_16428);
nor U18550 (N_18550,N_16969,N_17907);
nand U18551 (N_18551,N_17795,N_16262);
xor U18552 (N_18552,N_16656,N_16185);
nand U18553 (N_18553,N_17862,N_17904);
or U18554 (N_18554,N_17304,N_17658);
or U18555 (N_18555,N_16454,N_17884);
nand U18556 (N_18556,N_17677,N_16912);
xnor U18557 (N_18557,N_16646,N_17726);
nor U18558 (N_18558,N_17430,N_17429);
xnor U18559 (N_18559,N_17193,N_17633);
xnor U18560 (N_18560,N_17856,N_17044);
or U18561 (N_18561,N_16174,N_16409);
nand U18562 (N_18562,N_17230,N_17918);
or U18563 (N_18563,N_16029,N_16651);
and U18564 (N_18564,N_17655,N_16247);
or U18565 (N_18565,N_17794,N_17339);
and U18566 (N_18566,N_17162,N_17622);
and U18567 (N_18567,N_17009,N_17872);
nor U18568 (N_18568,N_16946,N_16130);
nand U18569 (N_18569,N_16553,N_17487);
or U18570 (N_18570,N_17854,N_16250);
or U18571 (N_18571,N_17326,N_17641);
nor U18572 (N_18572,N_16224,N_17973);
xnor U18573 (N_18573,N_16389,N_17147);
xnor U18574 (N_18574,N_17747,N_16714);
or U18575 (N_18575,N_16335,N_17962);
or U18576 (N_18576,N_16937,N_17219);
or U18577 (N_18577,N_16324,N_17186);
or U18578 (N_18578,N_17849,N_16592);
xor U18579 (N_18579,N_16464,N_17649);
xor U18580 (N_18580,N_17205,N_16201);
nor U18581 (N_18581,N_17846,N_17660);
nor U18582 (N_18582,N_16778,N_16210);
xor U18583 (N_18583,N_16837,N_17675);
nand U18584 (N_18584,N_16661,N_16960);
nand U18585 (N_18585,N_17384,N_17466);
or U18586 (N_18586,N_16791,N_16552);
and U18587 (N_18587,N_17553,N_17354);
nor U18588 (N_18588,N_16374,N_17331);
nor U18589 (N_18589,N_16541,N_16815);
and U18590 (N_18590,N_16636,N_16941);
or U18591 (N_18591,N_17797,N_17966);
or U18592 (N_18592,N_17086,N_16676);
xnor U18593 (N_18593,N_17855,N_17351);
nand U18594 (N_18594,N_16861,N_16444);
and U18595 (N_18595,N_17163,N_16684);
and U18596 (N_18596,N_16390,N_17451);
nand U18597 (N_18597,N_17704,N_16362);
xor U18598 (N_18598,N_16736,N_17925);
or U18599 (N_18599,N_17680,N_16800);
nand U18600 (N_18600,N_16734,N_17227);
xnor U18601 (N_18601,N_17251,N_17876);
and U18602 (N_18602,N_16259,N_16356);
nand U18603 (N_18603,N_17942,N_17175);
nand U18604 (N_18604,N_16988,N_17581);
and U18605 (N_18605,N_17837,N_17171);
nand U18606 (N_18606,N_16830,N_17050);
and U18607 (N_18607,N_17486,N_16423);
or U18608 (N_18608,N_16977,N_17779);
and U18609 (N_18609,N_17639,N_17493);
nand U18610 (N_18610,N_16504,N_16824);
nand U18611 (N_18611,N_17646,N_17133);
nand U18612 (N_18612,N_17647,N_16486);
and U18613 (N_18613,N_16929,N_16417);
nor U18614 (N_18614,N_16260,N_16365);
xnor U18615 (N_18615,N_16360,N_16896);
nand U18616 (N_18616,N_16924,N_17833);
or U18617 (N_18617,N_16545,N_16522);
or U18618 (N_18618,N_17280,N_16353);
nand U18619 (N_18619,N_16885,N_16421);
xor U18620 (N_18620,N_17830,N_17551);
and U18621 (N_18621,N_16268,N_16131);
or U18622 (N_18622,N_16986,N_17146);
and U18623 (N_18623,N_16339,N_16860);
nand U18624 (N_18624,N_17494,N_17920);
xor U18625 (N_18625,N_17483,N_17504);
nand U18626 (N_18626,N_17924,N_16805);
nor U18627 (N_18627,N_17287,N_17042);
nand U18628 (N_18628,N_16240,N_17959);
or U18629 (N_18629,N_17233,N_17482);
or U18630 (N_18630,N_16256,N_16267);
or U18631 (N_18631,N_17838,N_16691);
and U18632 (N_18632,N_16169,N_17990);
nand U18633 (N_18633,N_17928,N_17560);
or U18634 (N_18634,N_16441,N_17829);
and U18635 (N_18635,N_16735,N_16568);
nand U18636 (N_18636,N_17517,N_16618);
nor U18637 (N_18637,N_16715,N_16913);
and U18638 (N_18638,N_16003,N_16285);
or U18639 (N_18639,N_16214,N_16228);
nand U18640 (N_18640,N_16867,N_17405);
xor U18641 (N_18641,N_16564,N_16639);
nand U18642 (N_18642,N_17188,N_17465);
and U18643 (N_18643,N_17269,N_17932);
nor U18644 (N_18644,N_17977,N_17697);
xor U18645 (N_18645,N_16729,N_16298);
xnor U18646 (N_18646,N_17887,N_16832);
or U18647 (N_18647,N_17727,N_16921);
nor U18648 (N_18648,N_16105,N_16173);
xor U18649 (N_18649,N_17780,N_17378);
nand U18650 (N_18650,N_17993,N_17252);
xor U18651 (N_18651,N_17766,N_16014);
and U18652 (N_18652,N_16065,N_17082);
and U18653 (N_18653,N_16207,N_16099);
nor U18654 (N_18654,N_16872,N_17816);
nor U18655 (N_18655,N_17048,N_17945);
nor U18656 (N_18656,N_16300,N_16582);
xnor U18657 (N_18657,N_16205,N_17342);
nand U18658 (N_18658,N_17373,N_16244);
and U18659 (N_18659,N_17969,N_16447);
nand U18660 (N_18660,N_16510,N_16707);
nand U18661 (N_18661,N_16407,N_17519);
xor U18662 (N_18662,N_17107,N_17662);
xor U18663 (N_18663,N_16230,N_16233);
and U18664 (N_18664,N_17182,N_17877);
xnor U18665 (N_18665,N_16045,N_17406);
nor U18666 (N_18666,N_16166,N_16563);
xnor U18667 (N_18667,N_17305,N_16095);
xor U18668 (N_18668,N_16312,N_16278);
and U18669 (N_18669,N_16626,N_16709);
or U18670 (N_18670,N_16308,N_16429);
xor U18671 (N_18671,N_16048,N_17656);
nand U18672 (N_18672,N_17412,N_17526);
and U18673 (N_18673,N_17308,N_16370);
nor U18674 (N_18674,N_16783,N_16821);
or U18675 (N_18675,N_17700,N_17184);
and U18676 (N_18676,N_17614,N_17442);
nor U18677 (N_18677,N_16637,N_16314);
and U18678 (N_18678,N_17996,N_17364);
or U18679 (N_18679,N_16177,N_16165);
or U18680 (N_18680,N_17047,N_17645);
nor U18681 (N_18681,N_17968,N_17318);
nor U18682 (N_18682,N_16908,N_16248);
nor U18683 (N_18683,N_17018,N_17016);
nand U18684 (N_18684,N_17861,N_16967);
nor U18685 (N_18685,N_16396,N_16840);
nor U18686 (N_18686,N_17793,N_16839);
or U18687 (N_18687,N_17975,N_16693);
or U18688 (N_18688,N_16712,N_17394);
nor U18689 (N_18689,N_17689,N_17105);
xor U18690 (N_18690,N_17983,N_16007);
xnor U18691 (N_18691,N_16820,N_16810);
nor U18692 (N_18692,N_16155,N_16273);
nor U18693 (N_18693,N_16115,N_16221);
and U18694 (N_18694,N_17758,N_17259);
nor U18695 (N_18695,N_16648,N_17306);
and U18696 (N_18696,N_16763,N_16151);
xnor U18697 (N_18697,N_17490,N_17201);
and U18698 (N_18698,N_16943,N_16939);
nor U18699 (N_18699,N_17388,N_16851);
nand U18700 (N_18700,N_16238,N_17216);
nand U18701 (N_18701,N_17749,N_17153);
or U18702 (N_18702,N_16856,N_17937);
nor U18703 (N_18703,N_16041,N_16069);
or U18704 (N_18704,N_17441,N_17762);
or U18705 (N_18705,N_17832,N_17919);
xnor U18706 (N_18706,N_17106,N_17010);
xor U18707 (N_18707,N_17890,N_17488);
xnor U18708 (N_18708,N_16809,N_16516);
nand U18709 (N_18709,N_17603,N_16111);
or U18710 (N_18710,N_17365,N_16446);
xor U18711 (N_18711,N_17694,N_17223);
nand U18712 (N_18712,N_17020,N_16494);
nand U18713 (N_18713,N_16500,N_16291);
or U18714 (N_18714,N_16436,N_16874);
xor U18715 (N_18715,N_16227,N_16023);
or U18716 (N_18716,N_16938,N_17544);
nand U18717 (N_18717,N_16150,N_17729);
or U18718 (N_18718,N_16326,N_16013);
nor U18719 (N_18719,N_17620,N_17035);
xnor U18720 (N_18720,N_17938,N_16954);
nand U18721 (N_18721,N_17110,N_17853);
or U18722 (N_18722,N_17288,N_17325);
and U18723 (N_18723,N_17930,N_17496);
xor U18724 (N_18724,N_16459,N_16603);
xnor U18725 (N_18725,N_17464,N_17272);
xor U18726 (N_18726,N_17000,N_17593);
and U18727 (N_18727,N_16401,N_17058);
nor U18728 (N_18728,N_17019,N_17562);
nand U18729 (N_18729,N_17777,N_16718);
nand U18730 (N_18730,N_17262,N_16196);
and U18731 (N_18731,N_17963,N_17263);
and U18732 (N_18732,N_17864,N_16200);
nand U18733 (N_18733,N_16231,N_16520);
or U18734 (N_18734,N_16981,N_17640);
xor U18735 (N_18735,N_17253,N_17283);
nand U18736 (N_18736,N_16728,N_17611);
or U18737 (N_18737,N_17033,N_17616);
nand U18738 (N_18738,N_17788,N_16834);
and U18739 (N_18739,N_16951,N_16971);
xor U18740 (N_18740,N_16771,N_17353);
and U18741 (N_18741,N_17241,N_16453);
xnor U18742 (N_18742,N_16547,N_17868);
nor U18743 (N_18743,N_16350,N_17961);
or U18744 (N_18744,N_17786,N_16703);
nor U18745 (N_18745,N_17294,N_16973);
and U18746 (N_18746,N_17446,N_17202);
nand U18747 (N_18747,N_16999,N_17181);
xnor U18748 (N_18748,N_16744,N_17400);
nand U18749 (N_18749,N_16530,N_17618);
nand U18750 (N_18750,N_16662,N_17428);
nor U18751 (N_18751,N_17245,N_17899);
and U18752 (N_18752,N_16280,N_17360);
and U18753 (N_18753,N_17161,N_17583);
or U18754 (N_18754,N_17579,N_17636);
or U18755 (N_18755,N_17323,N_17467);
or U18756 (N_18756,N_16163,N_16580);
xnor U18757 (N_18757,N_16953,N_17841);
and U18758 (N_18758,N_16352,N_17783);
nor U18759 (N_18759,N_16669,N_17206);
xor U18760 (N_18760,N_16968,N_16393);
nor U18761 (N_18761,N_16292,N_16036);
or U18762 (N_18762,N_17166,N_17301);
xnor U18763 (N_18763,N_16540,N_17256);
xor U18764 (N_18764,N_17500,N_17905);
or U18765 (N_18765,N_16294,N_17129);
or U18766 (N_18766,N_16241,N_16819);
nand U18767 (N_18767,N_16024,N_16775);
nor U18768 (N_18768,N_16127,N_16601);
or U18769 (N_18769,N_17917,N_17445);
and U18770 (N_18770,N_16911,N_17495);
nor U18771 (N_18771,N_17322,N_17537);
nor U18772 (N_18772,N_16427,N_16471);
or U18773 (N_18773,N_17473,N_17764);
xnor U18774 (N_18774,N_16627,N_16061);
nor U18775 (N_18775,N_17200,N_16900);
or U18776 (N_18776,N_17534,N_17183);
and U18777 (N_18777,N_17902,N_17970);
nor U18778 (N_18778,N_16171,N_17874);
or U18779 (N_18779,N_16808,N_17597);
or U18780 (N_18780,N_17676,N_17674);
nor U18781 (N_18781,N_16643,N_17787);
or U18782 (N_18782,N_16406,N_16193);
or U18783 (N_18783,N_16845,N_16160);
and U18784 (N_18784,N_16950,N_16550);
and U18785 (N_18785,N_16257,N_17699);
nand U18786 (N_18786,N_16836,N_16076);
xor U18787 (N_18787,N_16681,N_16751);
or U18788 (N_18788,N_16873,N_17177);
and U18789 (N_18789,N_16758,N_17178);
and U18790 (N_18790,N_17080,N_16162);
and U18791 (N_18791,N_16319,N_16202);
nor U18792 (N_18792,N_16288,N_17939);
and U18793 (N_18793,N_17527,N_17099);
or U18794 (N_18794,N_17999,N_17577);
nand U18795 (N_18795,N_17678,N_16687);
or U18796 (N_18796,N_16653,N_17757);
xnor U18797 (N_18797,N_16829,N_16859);
nand U18798 (N_18798,N_17031,N_16961);
xnor U18799 (N_18799,N_16079,N_16381);
nor U18800 (N_18800,N_16063,N_17160);
or U18801 (N_18801,N_16738,N_16878);
and U18802 (N_18802,N_16664,N_16710);
or U18803 (N_18803,N_16302,N_17034);
nor U18804 (N_18804,N_16414,N_16144);
or U18805 (N_18805,N_17125,N_16518);
nand U18806 (N_18806,N_16000,N_16696);
xor U18807 (N_18807,N_17713,N_17679);
nand U18808 (N_18808,N_17385,N_17348);
or U18809 (N_18809,N_16386,N_17344);
or U18810 (N_18810,N_16433,N_17172);
nand U18811 (N_18811,N_16145,N_16606);
xnor U18812 (N_18812,N_17946,N_16889);
and U18813 (N_18813,N_16133,N_17532);
and U18814 (N_18814,N_16239,N_16368);
or U18815 (N_18815,N_16940,N_17424);
and U18816 (N_18816,N_17898,N_17140);
and U18817 (N_18817,N_16161,N_16679);
xnor U18818 (N_18818,N_17317,N_16920);
and U18819 (N_18819,N_17648,N_17204);
nor U18820 (N_18820,N_17931,N_17695);
nor U18821 (N_18821,N_17596,N_16817);
or U18822 (N_18822,N_17440,N_16502);
xnor U18823 (N_18823,N_16746,N_16286);
or U18824 (N_18824,N_17141,N_16304);
nand U18825 (N_18825,N_16613,N_16525);
and U18826 (N_18826,N_16706,N_17347);
xnor U18827 (N_18827,N_16899,N_17070);
or U18828 (N_18828,N_16671,N_17965);
and U18829 (N_18829,N_17191,N_16542);
nor U18830 (N_18830,N_16879,N_16534);
and U18831 (N_18831,N_16070,N_17213);
and U18832 (N_18832,N_17423,N_16877);
nand U18833 (N_18833,N_17261,N_17612);
nand U18834 (N_18834,N_17359,N_16237);
nand U18835 (N_18835,N_16320,N_16942);
or U18836 (N_18836,N_17421,N_17471);
and U18837 (N_18837,N_16103,N_17769);
xor U18838 (N_18838,N_16533,N_17529);
nand U18839 (N_18839,N_16596,N_16383);
or U18840 (N_18840,N_17731,N_16813);
nand U18841 (N_18841,N_16667,N_16711);
and U18842 (N_18842,N_16966,N_17479);
or U18843 (N_18843,N_17402,N_17302);
nand U18844 (N_18844,N_16577,N_17001);
or U18845 (N_18845,N_16054,N_17723);
nand U18846 (N_18846,N_16338,N_17132);
or U18847 (N_18847,N_16377,N_16616);
and U18848 (N_18848,N_17923,N_17737);
nor U18849 (N_18849,N_17803,N_16531);
and U18850 (N_18850,N_17081,N_16051);
nand U18851 (N_18851,N_17865,N_17075);
nand U18852 (N_18852,N_16897,N_16391);
nand U18853 (N_18853,N_17457,N_17906);
nor U18854 (N_18854,N_17187,N_16654);
nor U18855 (N_18855,N_16607,N_16917);
or U18856 (N_18856,N_16923,N_17684);
xor U18857 (N_18857,N_16602,N_16318);
and U18858 (N_18858,N_17870,N_16212);
or U18859 (N_18859,N_16721,N_16090);
or U18860 (N_18860,N_16147,N_16767);
nor U18861 (N_18861,N_17971,N_17666);
nand U18862 (N_18862,N_16538,N_17751);
nor U18863 (N_18863,N_17439,N_16647);
nor U18864 (N_18864,N_17574,N_17435);
xnor U18865 (N_18865,N_17499,N_16098);
and U18866 (N_18866,N_16991,N_17197);
xnor U18867 (N_18867,N_16594,N_16638);
and U18868 (N_18868,N_17735,N_16595);
xor U18869 (N_18869,N_17819,N_17023);
or U18870 (N_18870,N_16068,N_16781);
nand U18871 (N_18871,N_17743,N_17289);
nor U18872 (N_18872,N_16226,N_17916);
or U18873 (N_18873,N_16584,N_17372);
nand U18874 (N_18874,N_16588,N_17796);
nand U18875 (N_18875,N_17740,N_17345);
or U18876 (N_18876,N_16802,N_16680);
nand U18877 (N_18877,N_16842,N_17548);
nand U18878 (N_18878,N_17835,N_17895);
xnor U18879 (N_18879,N_16018,N_16380);
xnor U18880 (N_18880,N_16812,N_16918);
nor U18881 (N_18881,N_17295,N_16675);
xor U18882 (N_18882,N_17760,N_16022);
nor U18883 (N_18883,N_17297,N_17690);
and U18884 (N_18884,N_16970,N_17822);
nor U18885 (N_18885,N_16927,N_16330);
and U18886 (N_18886,N_16483,N_16102);
xor U18887 (N_18887,N_17820,N_16958);
and U18888 (N_18888,N_16779,N_17276);
nand U18889 (N_18889,N_17208,N_17102);
xor U18890 (N_18890,N_16044,N_16188);
or U18891 (N_18891,N_16104,N_16560);
and U18892 (N_18892,N_17711,N_16265);
nand U18893 (N_18893,N_16413,N_17761);
or U18894 (N_18894,N_17142,N_16843);
nand U18895 (N_18895,N_17460,N_16598);
nor U18896 (N_18896,N_17885,N_16620);
nor U18897 (N_18897,N_17808,N_17875);
and U18898 (N_18898,N_16723,N_16658);
nand U18899 (N_18899,N_16167,N_16978);
nor U18900 (N_18900,N_16379,N_17608);
nor U18901 (N_18901,N_17392,N_17456);
and U18902 (N_18902,N_16100,N_17626);
or U18903 (N_18903,N_16322,N_16053);
xnor U18904 (N_18904,N_17871,N_16756);
and U18905 (N_18905,N_16084,N_16902);
and U18906 (N_18906,N_16914,N_16615);
nand U18907 (N_18907,N_16722,N_17403);
or U18908 (N_18908,N_16790,N_17071);
or U18909 (N_18909,N_17356,N_16489);
xor U18910 (N_18910,N_16866,N_17371);
and U18911 (N_18911,N_17427,N_16574);
or U18912 (N_18912,N_16575,N_16597);
nand U18913 (N_18913,N_16197,N_16283);
xor U18914 (N_18914,N_16949,N_16006);
nand U18915 (N_18915,N_16215,N_17076);
nand U18916 (N_18916,N_16674,N_17866);
or U18917 (N_18917,N_17742,N_17686);
nor U18918 (N_18918,N_17117,N_17893);
and U18919 (N_18919,N_17654,N_17444);
xnor U18920 (N_18920,N_16138,N_16985);
and U18921 (N_18921,N_16306,N_17929);
nor U18922 (N_18922,N_16490,N_16276);
or U18923 (N_18923,N_17312,N_17357);
xor U18924 (N_18924,N_17002,N_17410);
xnor U18925 (N_18925,N_16644,N_17509);
and U18926 (N_18926,N_16211,N_16787);
nor U18927 (N_18927,N_17610,N_17006);
nand U18928 (N_18928,N_17409,N_17804);
nor U18929 (N_18929,N_17951,N_17222);
nor U18930 (N_18930,N_16847,N_16408);
nand U18931 (N_18931,N_16109,N_17176);
and U18932 (N_18932,N_17411,N_17341);
nand U18933 (N_18933,N_17390,N_17120);
and U18934 (N_18934,N_17955,N_17236);
nor U18935 (N_18935,N_16509,N_16660);
or U18936 (N_18936,N_16344,N_17065);
or U18937 (N_18937,N_16327,N_16052);
xor U18938 (N_18938,N_16916,N_17278);
nor U18939 (N_18939,N_16482,N_17491);
and U18940 (N_18940,N_17244,N_16686);
nor U18941 (N_18941,N_16556,N_16060);
or U18942 (N_18942,N_17707,N_17515);
nor U18943 (N_18943,N_16135,N_16229);
or U18944 (N_18944,N_17066,N_16038);
xnor U18945 (N_18945,N_17443,N_17881);
nand U18946 (N_18946,N_17566,N_17355);
xor U18947 (N_18947,N_16625,N_17981);
xor U18948 (N_18948,N_16869,N_17049);
nor U18949 (N_18949,N_17571,N_16119);
nor U18950 (N_18950,N_16299,N_16172);
nor U18951 (N_18951,N_16617,N_17771);
nor U18952 (N_18952,N_16782,N_16852);
nand U18953 (N_18953,N_16274,N_16690);
nor U18954 (N_18954,N_17903,N_17249);
or U18955 (N_18955,N_16222,N_17720);
and U18956 (N_18956,N_17157,N_17358);
or U18957 (N_18957,N_16505,N_16865);
and U18958 (N_18958,N_17869,N_17528);
nand U18959 (N_18959,N_17615,N_17934);
nor U18960 (N_18960,N_17037,N_16323);
nor U18961 (N_18961,N_16359,N_17809);
nor U18962 (N_18962,N_16213,N_17535);
or U18963 (N_18963,N_17823,N_16608);
xnor U18964 (N_18964,N_17416,N_17234);
xor U18965 (N_18965,N_16976,N_17291);
xnor U18966 (N_18966,N_17091,N_17046);
or U18967 (N_18967,N_16357,N_17032);
and U18968 (N_18968,N_16788,N_17590);
nor U18969 (N_18969,N_17221,N_16042);
or U18970 (N_18970,N_16378,N_16964);
nand U18971 (N_18971,N_17606,N_17840);
or U18972 (N_18972,N_17273,N_16366);
nor U18973 (N_18973,N_17734,N_16931);
nand U18974 (N_18974,N_17563,N_16796);
nand U18975 (N_18975,N_17825,N_17774);
nand U18976 (N_18976,N_16334,N_17138);
and U18977 (N_18977,N_17621,N_16769);
and U18978 (N_18978,N_17554,N_17386);
or U18979 (N_18979,N_17524,N_16488);
xnor U18980 (N_18980,N_17350,N_16948);
xnor U18981 (N_18981,N_17277,N_16906);
nor U18982 (N_18982,N_17103,N_16561);
xor U18983 (N_18983,N_16198,N_16717);
xnor U18984 (N_18984,N_16465,N_16216);
nor U18985 (N_18985,N_17926,N_17894);
nor U18986 (N_18986,N_17880,N_16612);
and U18987 (N_18987,N_17319,N_16551);
and U18988 (N_18988,N_17314,N_16922);
xor U18989 (N_18989,N_17850,N_16747);
nor U18990 (N_18990,N_17508,N_17398);
and U18991 (N_18991,N_16156,N_16011);
nand U18992 (N_18992,N_16452,N_16470);
and U18993 (N_18993,N_16142,N_16854);
and U18994 (N_18994,N_17549,N_16513);
nor U18995 (N_18995,N_16037,N_16956);
or U18996 (N_18996,N_16719,N_16622);
nand U18997 (N_18997,N_17060,N_16990);
xnor U18998 (N_18998,N_16762,N_17834);
nor U18999 (N_18999,N_16754,N_16512);
nand U19000 (N_19000,N_16245,N_17946);
or U19001 (N_19001,N_16101,N_17153);
nor U19002 (N_19002,N_17654,N_17222);
nand U19003 (N_19003,N_16792,N_16575);
nor U19004 (N_19004,N_17878,N_17883);
and U19005 (N_19005,N_17300,N_17071);
nor U19006 (N_19006,N_17665,N_17240);
and U19007 (N_19007,N_16588,N_17062);
or U19008 (N_19008,N_16799,N_17510);
xnor U19009 (N_19009,N_16195,N_16118);
or U19010 (N_19010,N_17766,N_16389);
xnor U19011 (N_19011,N_17805,N_17732);
nand U19012 (N_19012,N_16978,N_16640);
and U19013 (N_19013,N_17367,N_17977);
and U19014 (N_19014,N_17594,N_16033);
and U19015 (N_19015,N_16421,N_17581);
and U19016 (N_19016,N_17647,N_17282);
or U19017 (N_19017,N_16784,N_17248);
nand U19018 (N_19018,N_16948,N_17850);
nand U19019 (N_19019,N_17940,N_17826);
nor U19020 (N_19020,N_16004,N_17957);
and U19021 (N_19021,N_17105,N_16277);
nor U19022 (N_19022,N_16197,N_17328);
nand U19023 (N_19023,N_16717,N_17142);
and U19024 (N_19024,N_17784,N_17788);
and U19025 (N_19025,N_17280,N_16788);
nor U19026 (N_19026,N_16710,N_17915);
or U19027 (N_19027,N_17887,N_16926);
and U19028 (N_19028,N_16747,N_17990);
or U19029 (N_19029,N_17997,N_17522);
and U19030 (N_19030,N_17748,N_17276);
and U19031 (N_19031,N_16439,N_16915);
or U19032 (N_19032,N_16747,N_17439);
nor U19033 (N_19033,N_16849,N_17197);
and U19034 (N_19034,N_17434,N_16561);
nand U19035 (N_19035,N_16549,N_16618);
or U19036 (N_19036,N_17809,N_17946);
and U19037 (N_19037,N_17246,N_16959);
or U19038 (N_19038,N_17270,N_17410);
or U19039 (N_19039,N_17146,N_16291);
or U19040 (N_19040,N_17158,N_17680);
or U19041 (N_19041,N_17781,N_17355);
and U19042 (N_19042,N_16322,N_17808);
nand U19043 (N_19043,N_17424,N_17037);
nor U19044 (N_19044,N_17414,N_16813);
nand U19045 (N_19045,N_17110,N_16420);
nor U19046 (N_19046,N_17637,N_16077);
nor U19047 (N_19047,N_17768,N_17959);
nand U19048 (N_19048,N_17381,N_17814);
nand U19049 (N_19049,N_17198,N_16583);
or U19050 (N_19050,N_16818,N_17662);
nand U19051 (N_19051,N_16914,N_16836);
or U19052 (N_19052,N_16631,N_17191);
or U19053 (N_19053,N_17292,N_17106);
xor U19054 (N_19054,N_16804,N_17288);
nor U19055 (N_19055,N_16598,N_17806);
nor U19056 (N_19056,N_16718,N_16790);
nor U19057 (N_19057,N_16670,N_17672);
or U19058 (N_19058,N_16024,N_17447);
xor U19059 (N_19059,N_17288,N_16047);
and U19060 (N_19060,N_16246,N_16490);
and U19061 (N_19061,N_17225,N_16988);
and U19062 (N_19062,N_17325,N_17022);
xnor U19063 (N_19063,N_16047,N_16048);
and U19064 (N_19064,N_16651,N_16413);
or U19065 (N_19065,N_17957,N_17711);
or U19066 (N_19066,N_17055,N_17216);
and U19067 (N_19067,N_17260,N_16618);
or U19068 (N_19068,N_17800,N_16579);
and U19069 (N_19069,N_16816,N_16294);
nor U19070 (N_19070,N_16537,N_17874);
or U19071 (N_19071,N_17718,N_17836);
nand U19072 (N_19072,N_17439,N_17142);
or U19073 (N_19073,N_17123,N_17609);
and U19074 (N_19074,N_17433,N_16919);
or U19075 (N_19075,N_16710,N_16133);
and U19076 (N_19076,N_17521,N_17948);
nand U19077 (N_19077,N_17806,N_17484);
nand U19078 (N_19078,N_16515,N_17455);
xor U19079 (N_19079,N_17675,N_16159);
and U19080 (N_19080,N_17705,N_16973);
nor U19081 (N_19081,N_16412,N_17425);
nand U19082 (N_19082,N_16163,N_16126);
nand U19083 (N_19083,N_17636,N_17496);
nand U19084 (N_19084,N_17043,N_16703);
or U19085 (N_19085,N_17734,N_17319);
nand U19086 (N_19086,N_16439,N_17147);
xor U19087 (N_19087,N_16217,N_16913);
and U19088 (N_19088,N_16137,N_16329);
nor U19089 (N_19089,N_17582,N_16750);
nor U19090 (N_19090,N_16381,N_17525);
or U19091 (N_19091,N_16651,N_16367);
and U19092 (N_19092,N_17690,N_16570);
nor U19093 (N_19093,N_17490,N_16174);
or U19094 (N_19094,N_17704,N_16115);
and U19095 (N_19095,N_17641,N_17658);
or U19096 (N_19096,N_17012,N_16257);
and U19097 (N_19097,N_17685,N_17149);
nor U19098 (N_19098,N_16596,N_17586);
and U19099 (N_19099,N_16095,N_16759);
or U19100 (N_19100,N_17468,N_16063);
or U19101 (N_19101,N_17135,N_16650);
nor U19102 (N_19102,N_17826,N_17365);
nor U19103 (N_19103,N_17355,N_17659);
or U19104 (N_19104,N_17822,N_16646);
nor U19105 (N_19105,N_16602,N_16460);
or U19106 (N_19106,N_16981,N_17095);
xnor U19107 (N_19107,N_16046,N_16079);
or U19108 (N_19108,N_17584,N_16247);
or U19109 (N_19109,N_17801,N_16762);
and U19110 (N_19110,N_16155,N_16446);
and U19111 (N_19111,N_16912,N_16734);
or U19112 (N_19112,N_16504,N_16458);
xnor U19113 (N_19113,N_16208,N_17534);
and U19114 (N_19114,N_16684,N_17473);
or U19115 (N_19115,N_17104,N_17639);
xnor U19116 (N_19116,N_17813,N_16598);
nor U19117 (N_19117,N_16589,N_16427);
nor U19118 (N_19118,N_17865,N_17258);
nand U19119 (N_19119,N_17835,N_17769);
nor U19120 (N_19120,N_16087,N_16572);
xnor U19121 (N_19121,N_16033,N_16614);
and U19122 (N_19122,N_16742,N_17758);
nand U19123 (N_19123,N_16247,N_17606);
nor U19124 (N_19124,N_17427,N_16884);
nor U19125 (N_19125,N_17117,N_16819);
xnor U19126 (N_19126,N_16429,N_16673);
nand U19127 (N_19127,N_17724,N_17602);
xor U19128 (N_19128,N_17527,N_16240);
nand U19129 (N_19129,N_16003,N_16259);
nor U19130 (N_19130,N_17109,N_17382);
nand U19131 (N_19131,N_16439,N_17781);
nand U19132 (N_19132,N_17562,N_16958);
nand U19133 (N_19133,N_16569,N_17263);
and U19134 (N_19134,N_17082,N_16871);
nand U19135 (N_19135,N_17736,N_17217);
nand U19136 (N_19136,N_17773,N_16774);
or U19137 (N_19137,N_17850,N_16290);
and U19138 (N_19138,N_17138,N_17340);
and U19139 (N_19139,N_16296,N_17528);
nor U19140 (N_19140,N_17977,N_17117);
or U19141 (N_19141,N_16542,N_17744);
or U19142 (N_19142,N_17993,N_17648);
nand U19143 (N_19143,N_17848,N_16211);
nand U19144 (N_19144,N_17531,N_16033);
nand U19145 (N_19145,N_17154,N_17636);
nand U19146 (N_19146,N_16854,N_17081);
or U19147 (N_19147,N_16969,N_16669);
and U19148 (N_19148,N_17609,N_16958);
xor U19149 (N_19149,N_16275,N_16249);
and U19150 (N_19150,N_17969,N_16146);
xor U19151 (N_19151,N_16054,N_17182);
nand U19152 (N_19152,N_17788,N_16048);
and U19153 (N_19153,N_16361,N_16883);
xnor U19154 (N_19154,N_16049,N_16061);
nor U19155 (N_19155,N_16080,N_16940);
nor U19156 (N_19156,N_16016,N_17604);
nor U19157 (N_19157,N_17221,N_17061);
nor U19158 (N_19158,N_16049,N_16606);
or U19159 (N_19159,N_16016,N_17395);
and U19160 (N_19160,N_16557,N_16597);
or U19161 (N_19161,N_17256,N_17191);
xor U19162 (N_19162,N_17636,N_17087);
nor U19163 (N_19163,N_16644,N_16247);
xor U19164 (N_19164,N_17333,N_16544);
xnor U19165 (N_19165,N_16079,N_16795);
or U19166 (N_19166,N_17137,N_16343);
xor U19167 (N_19167,N_17154,N_16738);
nand U19168 (N_19168,N_16770,N_17412);
or U19169 (N_19169,N_16778,N_16943);
or U19170 (N_19170,N_16444,N_17205);
nand U19171 (N_19171,N_17936,N_16253);
xnor U19172 (N_19172,N_17267,N_17980);
or U19173 (N_19173,N_17612,N_17765);
and U19174 (N_19174,N_17248,N_16123);
nor U19175 (N_19175,N_17652,N_16503);
nand U19176 (N_19176,N_16332,N_17322);
nor U19177 (N_19177,N_16781,N_17729);
or U19178 (N_19178,N_17835,N_17142);
and U19179 (N_19179,N_17085,N_17425);
and U19180 (N_19180,N_16608,N_16355);
nor U19181 (N_19181,N_16526,N_16365);
or U19182 (N_19182,N_16115,N_16570);
nor U19183 (N_19183,N_16522,N_16299);
and U19184 (N_19184,N_16369,N_17604);
xor U19185 (N_19185,N_17556,N_16971);
and U19186 (N_19186,N_16369,N_17475);
nand U19187 (N_19187,N_17171,N_17703);
and U19188 (N_19188,N_17747,N_16241);
or U19189 (N_19189,N_16773,N_16901);
xnor U19190 (N_19190,N_17961,N_17651);
nor U19191 (N_19191,N_16371,N_16675);
nand U19192 (N_19192,N_17839,N_16312);
nor U19193 (N_19193,N_16784,N_16598);
xnor U19194 (N_19194,N_16480,N_16168);
or U19195 (N_19195,N_16652,N_16833);
nor U19196 (N_19196,N_16759,N_17726);
and U19197 (N_19197,N_16455,N_16666);
nor U19198 (N_19198,N_17731,N_16215);
nor U19199 (N_19199,N_17635,N_16780);
nand U19200 (N_19200,N_17559,N_17676);
nor U19201 (N_19201,N_17183,N_16483);
xnor U19202 (N_19202,N_16455,N_17535);
xnor U19203 (N_19203,N_17544,N_16732);
nand U19204 (N_19204,N_16390,N_16188);
or U19205 (N_19205,N_16779,N_16665);
and U19206 (N_19206,N_17193,N_16036);
xnor U19207 (N_19207,N_17269,N_17539);
nand U19208 (N_19208,N_16130,N_16969);
nor U19209 (N_19209,N_16196,N_16235);
xnor U19210 (N_19210,N_16959,N_16381);
and U19211 (N_19211,N_17950,N_16621);
xor U19212 (N_19212,N_17202,N_16914);
or U19213 (N_19213,N_17469,N_17656);
nand U19214 (N_19214,N_16706,N_16182);
and U19215 (N_19215,N_17891,N_16799);
nand U19216 (N_19216,N_16437,N_16442);
and U19217 (N_19217,N_16634,N_16935);
or U19218 (N_19218,N_16783,N_17904);
and U19219 (N_19219,N_17745,N_17115);
or U19220 (N_19220,N_17627,N_17733);
nor U19221 (N_19221,N_17432,N_17186);
or U19222 (N_19222,N_16133,N_17547);
and U19223 (N_19223,N_17657,N_17907);
or U19224 (N_19224,N_17030,N_16036);
xor U19225 (N_19225,N_16144,N_17117);
or U19226 (N_19226,N_17155,N_17957);
nand U19227 (N_19227,N_16628,N_16613);
or U19228 (N_19228,N_16062,N_17902);
nor U19229 (N_19229,N_17732,N_17487);
and U19230 (N_19230,N_17688,N_17975);
nor U19231 (N_19231,N_17501,N_16204);
or U19232 (N_19232,N_17012,N_16221);
nor U19233 (N_19233,N_17403,N_17510);
and U19234 (N_19234,N_17589,N_17137);
nand U19235 (N_19235,N_17907,N_17546);
nand U19236 (N_19236,N_17456,N_17120);
xnor U19237 (N_19237,N_17704,N_16658);
nor U19238 (N_19238,N_17848,N_16178);
nor U19239 (N_19239,N_17241,N_16294);
or U19240 (N_19240,N_17764,N_16735);
nor U19241 (N_19241,N_16293,N_17941);
nor U19242 (N_19242,N_16540,N_16407);
nand U19243 (N_19243,N_17647,N_16752);
nor U19244 (N_19244,N_17602,N_17594);
xor U19245 (N_19245,N_16656,N_16913);
nor U19246 (N_19246,N_17592,N_16501);
and U19247 (N_19247,N_17502,N_17935);
nand U19248 (N_19248,N_16565,N_17684);
nand U19249 (N_19249,N_17084,N_16484);
and U19250 (N_19250,N_16007,N_17007);
and U19251 (N_19251,N_17476,N_16996);
or U19252 (N_19252,N_17512,N_17041);
nor U19253 (N_19253,N_16302,N_17890);
nor U19254 (N_19254,N_16274,N_17202);
xnor U19255 (N_19255,N_16666,N_16529);
nor U19256 (N_19256,N_17461,N_17032);
nand U19257 (N_19257,N_17094,N_16388);
nand U19258 (N_19258,N_17263,N_17455);
nand U19259 (N_19259,N_16183,N_16311);
and U19260 (N_19260,N_17505,N_17720);
nor U19261 (N_19261,N_17696,N_16208);
nand U19262 (N_19262,N_16328,N_17828);
xnor U19263 (N_19263,N_17514,N_16039);
nor U19264 (N_19264,N_17344,N_17345);
nor U19265 (N_19265,N_17515,N_17908);
or U19266 (N_19266,N_17638,N_17798);
or U19267 (N_19267,N_17030,N_16726);
nand U19268 (N_19268,N_16687,N_17372);
and U19269 (N_19269,N_16641,N_17884);
and U19270 (N_19270,N_16301,N_16929);
nor U19271 (N_19271,N_17119,N_16242);
nand U19272 (N_19272,N_17408,N_17109);
xnor U19273 (N_19273,N_16307,N_17945);
or U19274 (N_19274,N_16434,N_17862);
or U19275 (N_19275,N_17521,N_17549);
nand U19276 (N_19276,N_16961,N_17876);
and U19277 (N_19277,N_17912,N_16568);
and U19278 (N_19278,N_16099,N_17991);
or U19279 (N_19279,N_17070,N_17656);
or U19280 (N_19280,N_17856,N_17788);
nor U19281 (N_19281,N_16622,N_17472);
xnor U19282 (N_19282,N_17392,N_16553);
nor U19283 (N_19283,N_17558,N_16175);
and U19284 (N_19284,N_17545,N_17366);
nand U19285 (N_19285,N_17840,N_16051);
nor U19286 (N_19286,N_16155,N_17379);
nor U19287 (N_19287,N_17346,N_17707);
or U19288 (N_19288,N_16007,N_17251);
nand U19289 (N_19289,N_17822,N_16401);
nand U19290 (N_19290,N_16749,N_16710);
xnor U19291 (N_19291,N_17047,N_17232);
or U19292 (N_19292,N_17714,N_16781);
nor U19293 (N_19293,N_17534,N_16503);
and U19294 (N_19294,N_17446,N_17909);
and U19295 (N_19295,N_16703,N_17074);
xnor U19296 (N_19296,N_16670,N_16949);
or U19297 (N_19297,N_16462,N_16980);
or U19298 (N_19298,N_17995,N_16197);
or U19299 (N_19299,N_17744,N_17923);
or U19300 (N_19300,N_16000,N_17502);
nor U19301 (N_19301,N_16789,N_16928);
xor U19302 (N_19302,N_17564,N_17487);
nor U19303 (N_19303,N_17000,N_16043);
nor U19304 (N_19304,N_17987,N_17901);
nand U19305 (N_19305,N_17315,N_17554);
or U19306 (N_19306,N_16563,N_17404);
and U19307 (N_19307,N_17065,N_17254);
nand U19308 (N_19308,N_17418,N_16240);
nand U19309 (N_19309,N_17877,N_16316);
nand U19310 (N_19310,N_17670,N_17992);
xnor U19311 (N_19311,N_17777,N_17141);
and U19312 (N_19312,N_17166,N_17967);
and U19313 (N_19313,N_16576,N_17763);
nor U19314 (N_19314,N_16290,N_16276);
and U19315 (N_19315,N_16034,N_16608);
or U19316 (N_19316,N_16407,N_16989);
and U19317 (N_19317,N_17433,N_17147);
xnor U19318 (N_19318,N_16253,N_17151);
nand U19319 (N_19319,N_16414,N_16430);
xnor U19320 (N_19320,N_16697,N_17789);
nand U19321 (N_19321,N_16189,N_17172);
xnor U19322 (N_19322,N_16833,N_17845);
nand U19323 (N_19323,N_16322,N_16418);
or U19324 (N_19324,N_17440,N_17098);
nand U19325 (N_19325,N_16750,N_16945);
or U19326 (N_19326,N_16598,N_17759);
nor U19327 (N_19327,N_16104,N_16357);
nand U19328 (N_19328,N_16083,N_16782);
nand U19329 (N_19329,N_16395,N_17745);
and U19330 (N_19330,N_16900,N_17296);
or U19331 (N_19331,N_16527,N_17180);
and U19332 (N_19332,N_17723,N_17502);
nand U19333 (N_19333,N_17680,N_16870);
nand U19334 (N_19334,N_16828,N_17944);
nor U19335 (N_19335,N_16876,N_16128);
nand U19336 (N_19336,N_16200,N_17212);
xor U19337 (N_19337,N_17745,N_16387);
nand U19338 (N_19338,N_16629,N_16479);
or U19339 (N_19339,N_17631,N_16109);
or U19340 (N_19340,N_16087,N_16178);
or U19341 (N_19341,N_16957,N_16782);
or U19342 (N_19342,N_16755,N_16815);
nor U19343 (N_19343,N_16318,N_17255);
nor U19344 (N_19344,N_16750,N_16582);
nor U19345 (N_19345,N_16847,N_17780);
nor U19346 (N_19346,N_16834,N_16181);
nand U19347 (N_19347,N_17907,N_16707);
xor U19348 (N_19348,N_17019,N_17854);
nand U19349 (N_19349,N_17441,N_17100);
nor U19350 (N_19350,N_17015,N_16959);
nand U19351 (N_19351,N_16519,N_16469);
nand U19352 (N_19352,N_17532,N_16857);
or U19353 (N_19353,N_17804,N_16891);
nor U19354 (N_19354,N_16866,N_16560);
or U19355 (N_19355,N_16701,N_16676);
or U19356 (N_19356,N_17010,N_17035);
xor U19357 (N_19357,N_16088,N_16198);
nor U19358 (N_19358,N_16354,N_16882);
xor U19359 (N_19359,N_16481,N_17607);
and U19360 (N_19360,N_17039,N_16043);
xor U19361 (N_19361,N_16752,N_16231);
xnor U19362 (N_19362,N_16322,N_16756);
or U19363 (N_19363,N_16477,N_16511);
or U19364 (N_19364,N_16179,N_16312);
nor U19365 (N_19365,N_16985,N_17623);
and U19366 (N_19366,N_16316,N_16110);
or U19367 (N_19367,N_17115,N_17531);
nand U19368 (N_19368,N_17866,N_17842);
and U19369 (N_19369,N_17074,N_17759);
nand U19370 (N_19370,N_17916,N_17029);
nor U19371 (N_19371,N_16686,N_16325);
xor U19372 (N_19372,N_17038,N_17848);
or U19373 (N_19373,N_16381,N_16350);
and U19374 (N_19374,N_16356,N_17943);
xor U19375 (N_19375,N_16123,N_17626);
or U19376 (N_19376,N_16272,N_16759);
and U19377 (N_19377,N_17665,N_17824);
xnor U19378 (N_19378,N_17989,N_16548);
or U19379 (N_19379,N_17500,N_16516);
nor U19380 (N_19380,N_17177,N_17677);
or U19381 (N_19381,N_17689,N_16214);
xnor U19382 (N_19382,N_16875,N_17110);
nor U19383 (N_19383,N_17330,N_17456);
or U19384 (N_19384,N_16586,N_17063);
nand U19385 (N_19385,N_17611,N_17751);
nand U19386 (N_19386,N_16791,N_17415);
nand U19387 (N_19387,N_17193,N_16778);
and U19388 (N_19388,N_16787,N_16244);
xnor U19389 (N_19389,N_16706,N_17237);
and U19390 (N_19390,N_16665,N_17171);
nor U19391 (N_19391,N_16182,N_16775);
xor U19392 (N_19392,N_17553,N_16486);
xor U19393 (N_19393,N_17244,N_17986);
nor U19394 (N_19394,N_17032,N_17604);
and U19395 (N_19395,N_16606,N_17851);
nor U19396 (N_19396,N_16206,N_17805);
xor U19397 (N_19397,N_16240,N_17560);
and U19398 (N_19398,N_17983,N_16814);
nand U19399 (N_19399,N_16429,N_16152);
nor U19400 (N_19400,N_17586,N_16346);
and U19401 (N_19401,N_17932,N_16954);
xor U19402 (N_19402,N_17973,N_17711);
or U19403 (N_19403,N_16312,N_17777);
xnor U19404 (N_19404,N_16443,N_16673);
nand U19405 (N_19405,N_17977,N_17201);
nand U19406 (N_19406,N_16611,N_17832);
nor U19407 (N_19407,N_17972,N_17229);
nor U19408 (N_19408,N_16867,N_17543);
nand U19409 (N_19409,N_16188,N_17668);
xnor U19410 (N_19410,N_16110,N_17344);
xnor U19411 (N_19411,N_16039,N_16747);
or U19412 (N_19412,N_17871,N_16986);
or U19413 (N_19413,N_16715,N_16710);
and U19414 (N_19414,N_17195,N_17663);
nor U19415 (N_19415,N_17347,N_16156);
and U19416 (N_19416,N_16060,N_16305);
nor U19417 (N_19417,N_17389,N_17952);
xnor U19418 (N_19418,N_16559,N_17927);
xor U19419 (N_19419,N_16108,N_17816);
xor U19420 (N_19420,N_17110,N_16715);
nor U19421 (N_19421,N_17814,N_16244);
or U19422 (N_19422,N_17156,N_17089);
or U19423 (N_19423,N_16651,N_16073);
xor U19424 (N_19424,N_17832,N_17906);
xor U19425 (N_19425,N_17479,N_16722);
nor U19426 (N_19426,N_17379,N_17577);
nand U19427 (N_19427,N_17216,N_16867);
or U19428 (N_19428,N_16856,N_17570);
xnor U19429 (N_19429,N_16218,N_16061);
nand U19430 (N_19430,N_16900,N_17002);
and U19431 (N_19431,N_16406,N_17340);
nor U19432 (N_19432,N_17123,N_17957);
or U19433 (N_19433,N_17628,N_17499);
or U19434 (N_19434,N_16318,N_17698);
and U19435 (N_19435,N_17073,N_16259);
xor U19436 (N_19436,N_16951,N_16027);
nand U19437 (N_19437,N_17685,N_16025);
or U19438 (N_19438,N_17031,N_17725);
nand U19439 (N_19439,N_17993,N_17099);
xnor U19440 (N_19440,N_17220,N_17637);
nor U19441 (N_19441,N_16228,N_17943);
and U19442 (N_19442,N_16426,N_16901);
nor U19443 (N_19443,N_17422,N_16715);
nand U19444 (N_19444,N_17954,N_16815);
and U19445 (N_19445,N_17999,N_17886);
nor U19446 (N_19446,N_16537,N_16167);
nand U19447 (N_19447,N_17807,N_16638);
or U19448 (N_19448,N_16382,N_17394);
and U19449 (N_19449,N_17888,N_16601);
or U19450 (N_19450,N_16585,N_16508);
and U19451 (N_19451,N_17751,N_17733);
and U19452 (N_19452,N_16481,N_16415);
nand U19453 (N_19453,N_16382,N_17576);
or U19454 (N_19454,N_16910,N_16357);
or U19455 (N_19455,N_16134,N_17591);
or U19456 (N_19456,N_17750,N_16579);
and U19457 (N_19457,N_17173,N_17400);
nor U19458 (N_19458,N_16262,N_17556);
and U19459 (N_19459,N_16989,N_17150);
or U19460 (N_19460,N_16890,N_17829);
xnor U19461 (N_19461,N_16050,N_17578);
or U19462 (N_19462,N_17278,N_16515);
and U19463 (N_19463,N_17666,N_17294);
xnor U19464 (N_19464,N_17166,N_17035);
nor U19465 (N_19465,N_17823,N_16699);
nand U19466 (N_19466,N_16685,N_17211);
xnor U19467 (N_19467,N_17057,N_16898);
or U19468 (N_19468,N_16901,N_16052);
nand U19469 (N_19469,N_17265,N_16858);
or U19470 (N_19470,N_16373,N_17111);
nand U19471 (N_19471,N_16691,N_17443);
or U19472 (N_19472,N_16080,N_17084);
nor U19473 (N_19473,N_16393,N_16079);
nor U19474 (N_19474,N_17016,N_17890);
nor U19475 (N_19475,N_17085,N_16003);
nor U19476 (N_19476,N_17568,N_17691);
nand U19477 (N_19477,N_16186,N_16552);
nand U19478 (N_19478,N_17882,N_17173);
nand U19479 (N_19479,N_17488,N_16354);
xor U19480 (N_19480,N_16672,N_16841);
or U19481 (N_19481,N_16862,N_17659);
nand U19482 (N_19482,N_17517,N_17264);
xor U19483 (N_19483,N_16081,N_17225);
nor U19484 (N_19484,N_17073,N_17434);
xnor U19485 (N_19485,N_17277,N_17492);
or U19486 (N_19486,N_16390,N_17447);
and U19487 (N_19487,N_16931,N_16490);
or U19488 (N_19488,N_16358,N_16209);
and U19489 (N_19489,N_16221,N_16026);
nor U19490 (N_19490,N_16462,N_17523);
and U19491 (N_19491,N_16826,N_17530);
xnor U19492 (N_19492,N_17183,N_17770);
and U19493 (N_19493,N_16137,N_17371);
and U19494 (N_19494,N_16624,N_17527);
xor U19495 (N_19495,N_16589,N_17642);
or U19496 (N_19496,N_16575,N_17664);
and U19497 (N_19497,N_17943,N_17668);
and U19498 (N_19498,N_16978,N_17777);
xor U19499 (N_19499,N_16642,N_16364);
and U19500 (N_19500,N_16649,N_16099);
or U19501 (N_19501,N_16511,N_17894);
xnor U19502 (N_19502,N_17208,N_16997);
or U19503 (N_19503,N_16774,N_16207);
nand U19504 (N_19504,N_16951,N_17061);
nand U19505 (N_19505,N_17172,N_17961);
and U19506 (N_19506,N_17337,N_16995);
nor U19507 (N_19507,N_16869,N_17303);
and U19508 (N_19508,N_16116,N_17494);
xnor U19509 (N_19509,N_17395,N_16614);
nand U19510 (N_19510,N_17148,N_16998);
or U19511 (N_19511,N_16532,N_17928);
xnor U19512 (N_19512,N_16139,N_17893);
nand U19513 (N_19513,N_17841,N_16830);
xor U19514 (N_19514,N_17770,N_17993);
or U19515 (N_19515,N_16325,N_16459);
or U19516 (N_19516,N_17028,N_16636);
nor U19517 (N_19517,N_17863,N_16661);
and U19518 (N_19518,N_16155,N_16536);
xor U19519 (N_19519,N_17697,N_17854);
and U19520 (N_19520,N_17567,N_17445);
and U19521 (N_19521,N_17319,N_16479);
nand U19522 (N_19522,N_17034,N_16717);
nor U19523 (N_19523,N_17765,N_17431);
nand U19524 (N_19524,N_16087,N_16219);
or U19525 (N_19525,N_16485,N_17395);
or U19526 (N_19526,N_17746,N_16651);
or U19527 (N_19527,N_16241,N_17377);
and U19528 (N_19528,N_17060,N_17972);
xor U19529 (N_19529,N_17807,N_17751);
nor U19530 (N_19530,N_17884,N_16480);
and U19531 (N_19531,N_16498,N_16435);
xnor U19532 (N_19532,N_16442,N_16528);
nand U19533 (N_19533,N_16625,N_17860);
nor U19534 (N_19534,N_17820,N_16820);
or U19535 (N_19535,N_16962,N_16182);
or U19536 (N_19536,N_17577,N_17239);
nor U19537 (N_19537,N_17057,N_16681);
nand U19538 (N_19538,N_17554,N_17695);
nor U19539 (N_19539,N_17294,N_16465);
and U19540 (N_19540,N_17959,N_17552);
and U19541 (N_19541,N_17904,N_16499);
nand U19542 (N_19542,N_17086,N_16305);
nand U19543 (N_19543,N_16186,N_16511);
nor U19544 (N_19544,N_16634,N_17178);
and U19545 (N_19545,N_16020,N_16613);
and U19546 (N_19546,N_17835,N_17180);
xor U19547 (N_19547,N_16932,N_17128);
nor U19548 (N_19548,N_16522,N_16382);
nand U19549 (N_19549,N_16611,N_17777);
or U19550 (N_19550,N_17325,N_17834);
or U19551 (N_19551,N_17927,N_17966);
nand U19552 (N_19552,N_16246,N_16356);
or U19553 (N_19553,N_16589,N_16500);
nor U19554 (N_19554,N_17159,N_16285);
nand U19555 (N_19555,N_17672,N_17525);
xor U19556 (N_19556,N_17466,N_16981);
and U19557 (N_19557,N_16798,N_17539);
or U19558 (N_19558,N_17999,N_16561);
or U19559 (N_19559,N_16449,N_16172);
nand U19560 (N_19560,N_16371,N_16729);
or U19561 (N_19561,N_16564,N_17269);
and U19562 (N_19562,N_16923,N_17258);
or U19563 (N_19563,N_16637,N_16880);
nor U19564 (N_19564,N_17288,N_17410);
or U19565 (N_19565,N_17873,N_16120);
xnor U19566 (N_19566,N_16476,N_17575);
nor U19567 (N_19567,N_16455,N_17620);
nor U19568 (N_19568,N_17147,N_17215);
nand U19569 (N_19569,N_16739,N_17179);
xor U19570 (N_19570,N_16250,N_17819);
or U19571 (N_19571,N_16292,N_17162);
nor U19572 (N_19572,N_16133,N_16160);
xnor U19573 (N_19573,N_17909,N_16463);
and U19574 (N_19574,N_16425,N_17676);
nor U19575 (N_19575,N_16087,N_17817);
nand U19576 (N_19576,N_16769,N_16679);
xor U19577 (N_19577,N_16704,N_16729);
or U19578 (N_19578,N_16628,N_17817);
or U19579 (N_19579,N_17718,N_17048);
or U19580 (N_19580,N_17645,N_16617);
nand U19581 (N_19581,N_17389,N_17390);
or U19582 (N_19582,N_16853,N_16364);
nand U19583 (N_19583,N_17126,N_16856);
nand U19584 (N_19584,N_17699,N_16811);
or U19585 (N_19585,N_16596,N_16305);
xor U19586 (N_19586,N_17533,N_17528);
and U19587 (N_19587,N_17691,N_17472);
nand U19588 (N_19588,N_16551,N_16087);
nand U19589 (N_19589,N_17227,N_16682);
or U19590 (N_19590,N_17790,N_17627);
xor U19591 (N_19591,N_16867,N_16341);
xnor U19592 (N_19592,N_16580,N_17383);
nor U19593 (N_19593,N_17180,N_17043);
nand U19594 (N_19594,N_17658,N_17578);
or U19595 (N_19595,N_16660,N_17224);
or U19596 (N_19596,N_16720,N_17167);
and U19597 (N_19597,N_17910,N_17397);
and U19598 (N_19598,N_16433,N_16039);
nor U19599 (N_19599,N_17764,N_16516);
or U19600 (N_19600,N_17843,N_16264);
and U19601 (N_19601,N_17737,N_17189);
nand U19602 (N_19602,N_16649,N_16833);
and U19603 (N_19603,N_16957,N_16572);
nor U19604 (N_19604,N_17591,N_17681);
nor U19605 (N_19605,N_17529,N_16676);
nand U19606 (N_19606,N_17578,N_16191);
nor U19607 (N_19607,N_17478,N_16987);
xnor U19608 (N_19608,N_17141,N_17485);
xor U19609 (N_19609,N_16272,N_16886);
nor U19610 (N_19610,N_16214,N_16294);
or U19611 (N_19611,N_16791,N_17554);
and U19612 (N_19612,N_16275,N_17557);
or U19613 (N_19613,N_16876,N_16955);
and U19614 (N_19614,N_16311,N_16111);
nor U19615 (N_19615,N_17959,N_17782);
nor U19616 (N_19616,N_17680,N_17496);
nand U19617 (N_19617,N_16973,N_17429);
nand U19618 (N_19618,N_16761,N_16532);
or U19619 (N_19619,N_17503,N_17174);
nand U19620 (N_19620,N_16797,N_17278);
xor U19621 (N_19621,N_16317,N_17672);
and U19622 (N_19622,N_16418,N_17683);
or U19623 (N_19623,N_16771,N_17189);
and U19624 (N_19624,N_17805,N_16618);
nor U19625 (N_19625,N_16405,N_17730);
nand U19626 (N_19626,N_16511,N_17218);
and U19627 (N_19627,N_17872,N_16007);
nand U19628 (N_19628,N_16590,N_16334);
and U19629 (N_19629,N_17824,N_17851);
nor U19630 (N_19630,N_17560,N_16517);
or U19631 (N_19631,N_17481,N_16952);
and U19632 (N_19632,N_17549,N_16447);
nand U19633 (N_19633,N_16659,N_17700);
nor U19634 (N_19634,N_16129,N_17460);
nor U19635 (N_19635,N_17225,N_17310);
nor U19636 (N_19636,N_16735,N_16924);
nand U19637 (N_19637,N_16227,N_16167);
or U19638 (N_19638,N_16026,N_17648);
or U19639 (N_19639,N_17030,N_17715);
and U19640 (N_19640,N_16659,N_17632);
or U19641 (N_19641,N_17236,N_16381);
and U19642 (N_19642,N_17652,N_16915);
nand U19643 (N_19643,N_17849,N_16348);
or U19644 (N_19644,N_17474,N_17506);
or U19645 (N_19645,N_17282,N_16802);
xnor U19646 (N_19646,N_16978,N_16455);
nor U19647 (N_19647,N_16621,N_16335);
or U19648 (N_19648,N_16110,N_16260);
or U19649 (N_19649,N_17591,N_16683);
or U19650 (N_19650,N_17599,N_16213);
nand U19651 (N_19651,N_17194,N_16157);
nand U19652 (N_19652,N_16415,N_16034);
or U19653 (N_19653,N_16403,N_16518);
nand U19654 (N_19654,N_16933,N_16778);
nor U19655 (N_19655,N_17682,N_16164);
or U19656 (N_19656,N_16252,N_16288);
or U19657 (N_19657,N_16643,N_16930);
nor U19658 (N_19658,N_17673,N_16463);
nor U19659 (N_19659,N_16836,N_17578);
or U19660 (N_19660,N_16183,N_17097);
nand U19661 (N_19661,N_16068,N_16061);
nor U19662 (N_19662,N_16377,N_17411);
nand U19663 (N_19663,N_16921,N_17498);
nand U19664 (N_19664,N_17283,N_16848);
nor U19665 (N_19665,N_17143,N_16817);
xor U19666 (N_19666,N_16389,N_16224);
or U19667 (N_19667,N_16240,N_17419);
nand U19668 (N_19668,N_16019,N_16636);
and U19669 (N_19669,N_17379,N_17648);
or U19670 (N_19670,N_16213,N_17839);
xor U19671 (N_19671,N_16725,N_17115);
nor U19672 (N_19672,N_17545,N_17094);
xnor U19673 (N_19673,N_16652,N_16093);
nand U19674 (N_19674,N_16868,N_17446);
or U19675 (N_19675,N_16873,N_16262);
nor U19676 (N_19676,N_16111,N_16920);
nand U19677 (N_19677,N_16220,N_16672);
or U19678 (N_19678,N_17451,N_17436);
or U19679 (N_19679,N_16589,N_17454);
nor U19680 (N_19680,N_16819,N_16384);
nand U19681 (N_19681,N_17819,N_17448);
xnor U19682 (N_19682,N_16942,N_16975);
and U19683 (N_19683,N_17397,N_17110);
and U19684 (N_19684,N_16356,N_16112);
nand U19685 (N_19685,N_17093,N_17730);
nor U19686 (N_19686,N_16717,N_16852);
nand U19687 (N_19687,N_16843,N_17216);
and U19688 (N_19688,N_16427,N_17249);
nor U19689 (N_19689,N_16993,N_16204);
nand U19690 (N_19690,N_17805,N_17583);
and U19691 (N_19691,N_16688,N_16354);
nand U19692 (N_19692,N_17823,N_16690);
nand U19693 (N_19693,N_17026,N_16708);
xnor U19694 (N_19694,N_16412,N_16602);
nand U19695 (N_19695,N_17059,N_17278);
or U19696 (N_19696,N_16764,N_17553);
or U19697 (N_19697,N_16353,N_17456);
xor U19698 (N_19698,N_16198,N_17794);
xor U19699 (N_19699,N_17059,N_16723);
or U19700 (N_19700,N_16239,N_17550);
and U19701 (N_19701,N_16111,N_16444);
xor U19702 (N_19702,N_16604,N_16885);
nand U19703 (N_19703,N_16133,N_17161);
xnor U19704 (N_19704,N_16168,N_17763);
nor U19705 (N_19705,N_17928,N_16165);
and U19706 (N_19706,N_17188,N_17931);
nor U19707 (N_19707,N_16829,N_16860);
xnor U19708 (N_19708,N_17209,N_17570);
and U19709 (N_19709,N_16958,N_17952);
or U19710 (N_19710,N_17826,N_17079);
xor U19711 (N_19711,N_16813,N_17316);
nand U19712 (N_19712,N_16781,N_16202);
or U19713 (N_19713,N_16201,N_17430);
nand U19714 (N_19714,N_17011,N_16202);
xnor U19715 (N_19715,N_16006,N_16681);
xor U19716 (N_19716,N_17912,N_16860);
nand U19717 (N_19717,N_17992,N_17274);
and U19718 (N_19718,N_17732,N_16242);
or U19719 (N_19719,N_17583,N_17465);
and U19720 (N_19720,N_16599,N_17864);
nand U19721 (N_19721,N_16552,N_16201);
nand U19722 (N_19722,N_17452,N_17693);
nor U19723 (N_19723,N_17113,N_16104);
or U19724 (N_19724,N_17010,N_17919);
xor U19725 (N_19725,N_16300,N_16918);
or U19726 (N_19726,N_17249,N_16955);
nor U19727 (N_19727,N_17344,N_17166);
nor U19728 (N_19728,N_16051,N_16810);
xnor U19729 (N_19729,N_16584,N_17188);
and U19730 (N_19730,N_17095,N_17809);
or U19731 (N_19731,N_17620,N_17451);
and U19732 (N_19732,N_17206,N_16076);
xnor U19733 (N_19733,N_17035,N_17693);
xor U19734 (N_19734,N_17686,N_17664);
nand U19735 (N_19735,N_17023,N_17073);
nor U19736 (N_19736,N_17461,N_17039);
xor U19737 (N_19737,N_16059,N_16632);
xnor U19738 (N_19738,N_16260,N_16462);
xor U19739 (N_19739,N_16671,N_16436);
xnor U19740 (N_19740,N_16397,N_17833);
and U19741 (N_19741,N_17178,N_17180);
nor U19742 (N_19742,N_17529,N_17396);
or U19743 (N_19743,N_17086,N_16186);
nand U19744 (N_19744,N_16335,N_17273);
nand U19745 (N_19745,N_16797,N_16509);
nand U19746 (N_19746,N_16920,N_16784);
nor U19747 (N_19747,N_16859,N_16297);
or U19748 (N_19748,N_16436,N_17001);
nand U19749 (N_19749,N_17802,N_16426);
xor U19750 (N_19750,N_17138,N_16278);
nand U19751 (N_19751,N_16075,N_17682);
nor U19752 (N_19752,N_17653,N_17361);
and U19753 (N_19753,N_17866,N_17331);
nand U19754 (N_19754,N_17262,N_17030);
and U19755 (N_19755,N_16580,N_17923);
and U19756 (N_19756,N_17268,N_17841);
or U19757 (N_19757,N_16718,N_17597);
xor U19758 (N_19758,N_17479,N_17110);
xor U19759 (N_19759,N_17447,N_17937);
xnor U19760 (N_19760,N_16799,N_16939);
xnor U19761 (N_19761,N_16362,N_17324);
and U19762 (N_19762,N_16892,N_17189);
xor U19763 (N_19763,N_16846,N_16885);
nand U19764 (N_19764,N_16568,N_17184);
and U19765 (N_19765,N_17966,N_17771);
nor U19766 (N_19766,N_17864,N_16442);
nor U19767 (N_19767,N_16521,N_17976);
xor U19768 (N_19768,N_16408,N_17288);
xor U19769 (N_19769,N_16348,N_17813);
xnor U19770 (N_19770,N_16517,N_16002);
and U19771 (N_19771,N_17349,N_16317);
or U19772 (N_19772,N_16883,N_16202);
nor U19773 (N_19773,N_17912,N_17632);
and U19774 (N_19774,N_17761,N_16393);
nor U19775 (N_19775,N_16820,N_16138);
nand U19776 (N_19776,N_16706,N_17325);
or U19777 (N_19777,N_16066,N_16012);
nand U19778 (N_19778,N_16989,N_16283);
or U19779 (N_19779,N_17931,N_16045);
nand U19780 (N_19780,N_16717,N_16008);
nand U19781 (N_19781,N_17974,N_17577);
and U19782 (N_19782,N_17762,N_16041);
nand U19783 (N_19783,N_16882,N_16676);
and U19784 (N_19784,N_17934,N_17566);
nand U19785 (N_19785,N_16247,N_17773);
and U19786 (N_19786,N_17515,N_17677);
xor U19787 (N_19787,N_17142,N_16873);
nand U19788 (N_19788,N_16501,N_17377);
and U19789 (N_19789,N_16442,N_17297);
or U19790 (N_19790,N_16062,N_17337);
or U19791 (N_19791,N_17341,N_17441);
and U19792 (N_19792,N_16717,N_16174);
or U19793 (N_19793,N_16077,N_16624);
nor U19794 (N_19794,N_16642,N_16014);
and U19795 (N_19795,N_17273,N_16775);
xnor U19796 (N_19796,N_16977,N_17567);
and U19797 (N_19797,N_17714,N_16860);
nand U19798 (N_19798,N_17564,N_16967);
and U19799 (N_19799,N_17445,N_17847);
nor U19800 (N_19800,N_16490,N_17660);
or U19801 (N_19801,N_17744,N_16102);
nand U19802 (N_19802,N_16803,N_17840);
and U19803 (N_19803,N_16019,N_16548);
or U19804 (N_19804,N_17648,N_17921);
or U19805 (N_19805,N_16416,N_17599);
nand U19806 (N_19806,N_16533,N_16385);
and U19807 (N_19807,N_17789,N_16239);
or U19808 (N_19808,N_16171,N_16509);
nor U19809 (N_19809,N_16997,N_17061);
or U19810 (N_19810,N_17767,N_17176);
and U19811 (N_19811,N_16816,N_17991);
or U19812 (N_19812,N_16147,N_17502);
and U19813 (N_19813,N_16940,N_17676);
nor U19814 (N_19814,N_17400,N_16365);
or U19815 (N_19815,N_16337,N_17263);
or U19816 (N_19816,N_17256,N_17400);
xor U19817 (N_19817,N_16111,N_17641);
nand U19818 (N_19818,N_16609,N_17551);
and U19819 (N_19819,N_16631,N_17315);
xor U19820 (N_19820,N_17379,N_17046);
and U19821 (N_19821,N_17042,N_16906);
nand U19822 (N_19822,N_17233,N_16720);
nor U19823 (N_19823,N_16305,N_17594);
xnor U19824 (N_19824,N_17647,N_17184);
and U19825 (N_19825,N_17156,N_16552);
nand U19826 (N_19826,N_16268,N_17598);
or U19827 (N_19827,N_16655,N_16153);
or U19828 (N_19828,N_16483,N_16640);
and U19829 (N_19829,N_17543,N_17032);
xnor U19830 (N_19830,N_16311,N_17696);
nor U19831 (N_19831,N_16210,N_17864);
nor U19832 (N_19832,N_17610,N_16885);
or U19833 (N_19833,N_17301,N_16738);
xnor U19834 (N_19834,N_17452,N_17670);
or U19835 (N_19835,N_16861,N_17830);
nand U19836 (N_19836,N_17734,N_17575);
or U19837 (N_19837,N_17852,N_16327);
nand U19838 (N_19838,N_16198,N_17418);
or U19839 (N_19839,N_17997,N_17197);
and U19840 (N_19840,N_17344,N_16162);
or U19841 (N_19841,N_16086,N_16797);
or U19842 (N_19842,N_16832,N_16330);
and U19843 (N_19843,N_17947,N_16766);
nor U19844 (N_19844,N_16848,N_16413);
nor U19845 (N_19845,N_16950,N_17664);
or U19846 (N_19846,N_17797,N_16536);
or U19847 (N_19847,N_17474,N_17243);
nor U19848 (N_19848,N_17840,N_16989);
nand U19849 (N_19849,N_17019,N_17252);
nand U19850 (N_19850,N_16606,N_17009);
nor U19851 (N_19851,N_17996,N_16939);
nor U19852 (N_19852,N_17109,N_16627);
and U19853 (N_19853,N_16096,N_17276);
or U19854 (N_19854,N_17113,N_17690);
or U19855 (N_19855,N_17964,N_17691);
nor U19856 (N_19856,N_16785,N_16200);
and U19857 (N_19857,N_17781,N_17947);
xor U19858 (N_19858,N_16512,N_17191);
and U19859 (N_19859,N_16196,N_17123);
nor U19860 (N_19860,N_16689,N_16780);
nand U19861 (N_19861,N_17985,N_17651);
or U19862 (N_19862,N_17639,N_16604);
and U19863 (N_19863,N_16796,N_17734);
and U19864 (N_19864,N_16845,N_17867);
or U19865 (N_19865,N_16843,N_17300);
nor U19866 (N_19866,N_17049,N_16406);
and U19867 (N_19867,N_17093,N_17246);
xor U19868 (N_19868,N_16950,N_16825);
nor U19869 (N_19869,N_16286,N_17190);
nor U19870 (N_19870,N_16881,N_17142);
nand U19871 (N_19871,N_16887,N_17023);
nand U19872 (N_19872,N_16501,N_17394);
xnor U19873 (N_19873,N_16238,N_17001);
nor U19874 (N_19874,N_16536,N_17964);
nor U19875 (N_19875,N_17867,N_16559);
nand U19876 (N_19876,N_17330,N_17575);
nand U19877 (N_19877,N_16085,N_17244);
xor U19878 (N_19878,N_16818,N_16393);
nor U19879 (N_19879,N_16372,N_16924);
xor U19880 (N_19880,N_16722,N_16430);
and U19881 (N_19881,N_16406,N_16423);
nand U19882 (N_19882,N_16780,N_17655);
or U19883 (N_19883,N_16910,N_17307);
and U19884 (N_19884,N_17107,N_17775);
nor U19885 (N_19885,N_16312,N_16036);
nor U19886 (N_19886,N_17046,N_17713);
or U19887 (N_19887,N_16451,N_17281);
nor U19888 (N_19888,N_17207,N_17958);
and U19889 (N_19889,N_17150,N_16591);
nand U19890 (N_19890,N_17168,N_17249);
nor U19891 (N_19891,N_16783,N_17884);
nor U19892 (N_19892,N_16017,N_17438);
nor U19893 (N_19893,N_17150,N_16474);
or U19894 (N_19894,N_17948,N_17296);
nor U19895 (N_19895,N_16193,N_16083);
nand U19896 (N_19896,N_16466,N_17525);
or U19897 (N_19897,N_16695,N_16623);
or U19898 (N_19898,N_16668,N_16512);
nor U19899 (N_19899,N_16328,N_17786);
xnor U19900 (N_19900,N_16655,N_16549);
or U19901 (N_19901,N_16400,N_17824);
nand U19902 (N_19902,N_17802,N_17094);
nor U19903 (N_19903,N_16269,N_16066);
nor U19904 (N_19904,N_17138,N_16989);
xor U19905 (N_19905,N_16969,N_17980);
xor U19906 (N_19906,N_16350,N_16550);
or U19907 (N_19907,N_16344,N_17371);
or U19908 (N_19908,N_17648,N_17003);
nand U19909 (N_19909,N_16557,N_16544);
or U19910 (N_19910,N_17805,N_17309);
and U19911 (N_19911,N_17501,N_17293);
nand U19912 (N_19912,N_16964,N_17671);
and U19913 (N_19913,N_16905,N_16641);
xor U19914 (N_19914,N_17098,N_16262);
nand U19915 (N_19915,N_16062,N_16090);
xnor U19916 (N_19916,N_17188,N_17717);
xor U19917 (N_19917,N_17969,N_17647);
or U19918 (N_19918,N_17948,N_17992);
nand U19919 (N_19919,N_17037,N_17481);
or U19920 (N_19920,N_17236,N_17079);
nand U19921 (N_19921,N_17098,N_17924);
and U19922 (N_19922,N_16693,N_16857);
nand U19923 (N_19923,N_16758,N_17328);
and U19924 (N_19924,N_17798,N_16461);
nor U19925 (N_19925,N_16271,N_16699);
nand U19926 (N_19926,N_16500,N_17615);
nor U19927 (N_19927,N_16281,N_16103);
nor U19928 (N_19928,N_17330,N_17124);
or U19929 (N_19929,N_16587,N_17089);
nand U19930 (N_19930,N_16605,N_17263);
or U19931 (N_19931,N_17678,N_16455);
nand U19932 (N_19932,N_16520,N_17059);
and U19933 (N_19933,N_17611,N_16816);
nor U19934 (N_19934,N_17744,N_16626);
and U19935 (N_19935,N_16229,N_16055);
or U19936 (N_19936,N_16209,N_16205);
and U19937 (N_19937,N_16065,N_16155);
and U19938 (N_19938,N_17932,N_17563);
and U19939 (N_19939,N_17922,N_16654);
and U19940 (N_19940,N_16100,N_16054);
and U19941 (N_19941,N_16751,N_17007);
and U19942 (N_19942,N_17030,N_17101);
nor U19943 (N_19943,N_17176,N_17890);
nor U19944 (N_19944,N_17474,N_16001);
nand U19945 (N_19945,N_16171,N_17644);
nor U19946 (N_19946,N_17236,N_17776);
nand U19947 (N_19947,N_16276,N_17993);
or U19948 (N_19948,N_16569,N_17454);
xor U19949 (N_19949,N_16566,N_17266);
nand U19950 (N_19950,N_16791,N_17328);
nand U19951 (N_19951,N_16256,N_16236);
xnor U19952 (N_19952,N_17067,N_16835);
xor U19953 (N_19953,N_17170,N_17275);
nor U19954 (N_19954,N_16994,N_17904);
nor U19955 (N_19955,N_17287,N_17103);
or U19956 (N_19956,N_17078,N_17330);
nor U19957 (N_19957,N_16153,N_17827);
nand U19958 (N_19958,N_17922,N_17758);
xnor U19959 (N_19959,N_16682,N_16745);
or U19960 (N_19960,N_17688,N_16128);
nor U19961 (N_19961,N_17409,N_16754);
xnor U19962 (N_19962,N_16355,N_16989);
xnor U19963 (N_19963,N_16476,N_16223);
nand U19964 (N_19964,N_17678,N_16603);
xor U19965 (N_19965,N_17045,N_16172);
xnor U19966 (N_19966,N_17163,N_16234);
and U19967 (N_19967,N_17571,N_17417);
or U19968 (N_19968,N_17946,N_17070);
and U19969 (N_19969,N_16087,N_17138);
nor U19970 (N_19970,N_17780,N_16529);
and U19971 (N_19971,N_17484,N_17531);
or U19972 (N_19972,N_17068,N_16013);
or U19973 (N_19973,N_16209,N_16645);
and U19974 (N_19974,N_17160,N_17218);
xor U19975 (N_19975,N_16171,N_16098);
nand U19976 (N_19976,N_17428,N_17536);
nand U19977 (N_19977,N_17286,N_16349);
nor U19978 (N_19978,N_17443,N_17930);
or U19979 (N_19979,N_17852,N_16148);
nor U19980 (N_19980,N_17955,N_17934);
or U19981 (N_19981,N_16630,N_17139);
nand U19982 (N_19982,N_17337,N_17389);
and U19983 (N_19983,N_17004,N_17371);
nor U19984 (N_19984,N_16573,N_16479);
nor U19985 (N_19985,N_16233,N_16418);
nor U19986 (N_19986,N_16100,N_16312);
or U19987 (N_19987,N_17613,N_16655);
nor U19988 (N_19988,N_16366,N_16724);
nor U19989 (N_19989,N_17666,N_17504);
and U19990 (N_19990,N_17270,N_17918);
nand U19991 (N_19991,N_16726,N_17947);
nand U19992 (N_19992,N_17031,N_17302);
or U19993 (N_19993,N_16021,N_16983);
and U19994 (N_19994,N_16129,N_17330);
nor U19995 (N_19995,N_17998,N_16726);
or U19996 (N_19996,N_17121,N_16514);
or U19997 (N_19997,N_17697,N_16170);
xnor U19998 (N_19998,N_16210,N_17254);
xor U19999 (N_19999,N_17398,N_17397);
nand U20000 (N_20000,N_19379,N_19864);
and U20001 (N_20001,N_19048,N_19870);
nand U20002 (N_20002,N_18473,N_18225);
and U20003 (N_20003,N_19543,N_18222);
xor U20004 (N_20004,N_19767,N_18462);
xor U20005 (N_20005,N_19112,N_18638);
nand U20006 (N_20006,N_19797,N_18962);
and U20007 (N_20007,N_19440,N_18488);
and U20008 (N_20008,N_19574,N_19737);
or U20009 (N_20009,N_19537,N_18074);
nand U20010 (N_20010,N_18677,N_18387);
nor U20011 (N_20011,N_18291,N_18773);
or U20012 (N_20012,N_18315,N_18292);
nor U20013 (N_20013,N_18851,N_19142);
nor U20014 (N_20014,N_19776,N_19289);
and U20015 (N_20015,N_18525,N_19041);
or U20016 (N_20016,N_18517,N_18068);
or U20017 (N_20017,N_19255,N_18153);
and U20018 (N_20018,N_18922,N_19400);
nor U20019 (N_20019,N_19403,N_18701);
xor U20020 (N_20020,N_19113,N_18665);
or U20021 (N_20021,N_19661,N_18166);
nand U20022 (N_20022,N_18944,N_18937);
and U20023 (N_20023,N_18800,N_18644);
xnor U20024 (N_20024,N_18618,N_18147);
and U20025 (N_20025,N_18847,N_18231);
nand U20026 (N_20026,N_19907,N_19587);
nand U20027 (N_20027,N_18359,N_19016);
nand U20028 (N_20028,N_19830,N_19828);
nand U20029 (N_20029,N_18641,N_19798);
nor U20030 (N_20030,N_18753,N_18588);
xor U20031 (N_20031,N_19866,N_19770);
and U20032 (N_20032,N_18293,N_19415);
nor U20033 (N_20033,N_18016,N_19003);
or U20034 (N_20034,N_18109,N_18894);
nor U20035 (N_20035,N_18828,N_18207);
nor U20036 (N_20036,N_19859,N_19634);
xor U20037 (N_20037,N_18341,N_18816);
nor U20038 (N_20038,N_18725,N_18782);
and U20039 (N_20039,N_19629,N_18549);
nand U20040 (N_20040,N_19957,N_19512);
nor U20041 (N_20041,N_19410,N_18660);
or U20042 (N_20042,N_18758,N_19580);
nand U20043 (N_20043,N_19244,N_19817);
and U20044 (N_20044,N_19692,N_18880);
and U20045 (N_20045,N_18324,N_18986);
xor U20046 (N_20046,N_19758,N_18072);
nand U20047 (N_20047,N_19240,N_19678);
nor U20048 (N_20048,N_19900,N_19356);
nor U20049 (N_20049,N_19560,N_19811);
nor U20050 (N_20050,N_19052,N_18904);
xor U20051 (N_20051,N_18430,N_19098);
and U20052 (N_20052,N_19691,N_19838);
and U20053 (N_20053,N_19931,N_18846);
or U20054 (N_20054,N_18999,N_19852);
nor U20055 (N_20055,N_18289,N_19552);
nor U20056 (N_20056,N_18557,N_18502);
or U20057 (N_20057,N_18251,N_19844);
nor U20058 (N_20058,N_19597,N_18426);
and U20059 (N_20059,N_18405,N_19999);
and U20060 (N_20060,N_18746,N_19087);
nor U20061 (N_20061,N_18843,N_19382);
or U20062 (N_20062,N_18622,N_19605);
and U20063 (N_20063,N_19502,N_18181);
nor U20064 (N_20064,N_19687,N_19210);
nor U20065 (N_20065,N_18331,N_19668);
nor U20066 (N_20066,N_18516,N_18531);
and U20067 (N_20067,N_19059,N_18271);
and U20068 (N_20068,N_19395,N_18204);
or U20069 (N_20069,N_19173,N_19461);
xnor U20070 (N_20070,N_19856,N_18952);
xor U20071 (N_20071,N_18757,N_19677);
or U20072 (N_20072,N_19444,N_19071);
nor U20073 (N_20073,N_18939,N_19082);
xnor U20074 (N_20074,N_18185,N_19810);
xnor U20075 (N_20075,N_18711,N_18739);
and U20076 (N_20076,N_18724,N_18945);
and U20077 (N_20077,N_19008,N_19463);
or U20078 (N_20078,N_18110,N_19279);
or U20079 (N_20079,N_18871,N_19219);
or U20080 (N_20080,N_19061,N_19997);
xor U20081 (N_20081,N_18955,N_18336);
nor U20082 (N_20082,N_19841,N_18447);
nand U20083 (N_20083,N_18888,N_18223);
or U20084 (N_20084,N_18610,N_18813);
or U20085 (N_20085,N_19062,N_18522);
nand U20086 (N_20086,N_18442,N_19096);
xnor U20087 (N_20087,N_19660,N_18551);
nand U20088 (N_20088,N_18797,N_18138);
nand U20089 (N_20089,N_19871,N_19419);
nand U20090 (N_20090,N_19386,N_19753);
nand U20091 (N_20091,N_18221,N_19538);
nor U20092 (N_20092,N_18314,N_19044);
nand U20093 (N_20093,N_18349,N_19187);
xnor U20094 (N_20094,N_19066,N_19357);
xnor U20095 (N_20095,N_18056,N_18587);
or U20096 (N_20096,N_18268,N_19249);
nand U20097 (N_20097,N_19088,N_19441);
and U20098 (N_20098,N_18506,N_18270);
or U20099 (N_20099,N_18450,N_18694);
or U20100 (N_20100,N_19092,N_18403);
nor U20101 (N_20101,N_18055,N_19134);
xor U20102 (N_20102,N_19254,N_18855);
and U20103 (N_20103,N_19701,N_18135);
and U20104 (N_20104,N_18494,N_18862);
or U20105 (N_20105,N_18479,N_18564);
and U20106 (N_20106,N_18500,N_19328);
or U20107 (N_20107,N_18371,N_19268);
or U20108 (N_20108,N_19780,N_19839);
xor U20109 (N_20109,N_18111,N_19887);
or U20110 (N_20110,N_18358,N_18712);
nor U20111 (N_20111,N_18678,N_18234);
nand U20112 (N_20112,N_19028,N_18614);
nand U20113 (N_20113,N_19936,N_19848);
xnor U20114 (N_20114,N_19332,N_18714);
nor U20115 (N_20115,N_18383,N_18240);
and U20116 (N_20116,N_18467,N_19821);
xor U20117 (N_20117,N_19026,N_19968);
and U20118 (N_20118,N_18495,N_18245);
or U20119 (N_20119,N_19470,N_19034);
xnor U20120 (N_20120,N_18584,N_19509);
or U20121 (N_20121,N_19773,N_19290);
nor U20122 (N_20122,N_19549,N_19032);
nand U20123 (N_20123,N_19104,N_18187);
nand U20124 (N_20124,N_19796,N_18217);
xor U20125 (N_20125,N_19202,N_18049);
xnor U20126 (N_20126,N_19081,N_19937);
nand U20127 (N_20127,N_19731,N_18446);
or U20128 (N_20128,N_19133,N_19638);
xnor U20129 (N_20129,N_18202,N_19438);
xor U20130 (N_20130,N_19238,N_19570);
xnor U20131 (N_20131,N_18316,N_18449);
nand U20132 (N_20132,N_18091,N_19909);
or U20133 (N_20133,N_18784,N_18670);
nor U20134 (N_20134,N_19364,N_19732);
nand U20135 (N_20135,N_18415,N_18378);
nor U20136 (N_20136,N_19013,N_19805);
nand U20137 (N_20137,N_18968,N_19948);
nand U20138 (N_20138,N_19884,N_18076);
xor U20139 (N_20139,N_19945,N_19788);
and U20140 (N_20140,N_19488,N_18444);
and U20141 (N_20141,N_19644,N_19453);
nand U20142 (N_20142,N_19327,N_19212);
nand U20143 (N_20143,N_18421,N_19380);
and U20144 (N_20144,N_19342,N_19895);
nand U20145 (N_20145,N_18157,N_18377);
nor U20146 (N_20146,N_18553,N_19695);
and U20147 (N_20147,N_19194,N_18794);
nor U20148 (N_20148,N_19850,N_19611);
xor U20149 (N_20149,N_19954,N_19733);
nor U20150 (N_20150,N_19860,N_19103);
and U20151 (N_20151,N_19037,N_19992);
nand U20152 (N_20152,N_18640,N_18165);
nand U20153 (N_20153,N_18134,N_18485);
nand U20154 (N_20154,N_19829,N_18063);
and U20155 (N_20155,N_18875,N_19426);
nor U20156 (N_20156,N_19744,N_18649);
xnor U20157 (N_20157,N_18560,N_18713);
nand U20158 (N_20158,N_18869,N_19741);
xor U20159 (N_20159,N_18342,N_19506);
and U20160 (N_20160,N_19961,N_19130);
and U20161 (N_20161,N_19431,N_18154);
and U20162 (N_20162,N_19083,N_19736);
nand U20163 (N_20163,N_18936,N_19181);
xor U20164 (N_20164,N_19647,N_19162);
xnor U20165 (N_20165,N_18353,N_19681);
or U20166 (N_20166,N_19861,N_18152);
and U20167 (N_20167,N_18589,N_19942);
and U20168 (N_20168,N_18868,N_18681);
nand U20169 (N_20169,N_18770,N_19529);
nor U20170 (N_20170,N_18971,N_19418);
and U20171 (N_20171,N_19216,N_18745);
or U20172 (N_20172,N_18991,N_18642);
or U20173 (N_20173,N_18018,N_19685);
and U20174 (N_20174,N_18008,N_18386);
xor U20175 (N_20175,N_18989,N_18831);
nor U20176 (N_20176,N_19778,N_18747);
xnor U20177 (N_20177,N_18893,N_18651);
and U20178 (N_20178,N_19427,N_18431);
nor U20179 (N_20179,N_18535,N_18071);
or U20180 (N_20180,N_18585,N_18212);
nand U20181 (N_20181,N_18059,N_18634);
nor U20182 (N_20182,N_18252,N_18572);
xnor U20183 (N_20183,N_19117,N_18174);
nand U20184 (N_20184,N_19513,N_18787);
and U20185 (N_20185,N_19399,N_19054);
xnor U20186 (N_20186,N_18227,N_19190);
nor U20187 (N_20187,N_19609,N_18464);
or U20188 (N_20188,N_18329,N_18710);
or U20189 (N_20189,N_18605,N_18092);
and U20190 (N_20190,N_19304,N_18633);
xnor U20191 (N_20191,N_18379,N_18674);
nand U20192 (N_20192,N_19696,N_19703);
nand U20193 (N_20193,N_19458,N_19094);
or U20194 (N_20194,N_18086,N_18796);
and U20195 (N_20195,N_19141,N_18445);
nor U20196 (N_20196,N_19152,N_18775);
and U20197 (N_20197,N_19772,N_18598);
or U20198 (N_20198,N_18900,N_19667);
and U20199 (N_20199,N_18139,N_19230);
nand U20200 (N_20200,N_18244,N_18041);
nor U20201 (N_20201,N_19205,N_19110);
nor U20202 (N_20202,N_19613,N_18285);
and U20203 (N_20203,N_19006,N_18256);
nand U20204 (N_20204,N_18934,N_19734);
xnor U20205 (N_20205,N_18106,N_19567);
and U20206 (N_20206,N_18366,N_18057);
or U20207 (N_20207,N_19336,N_18304);
or U20208 (N_20208,N_19615,N_19793);
and U20209 (N_20209,N_18803,N_18399);
nand U20210 (N_20210,N_19000,N_18509);
or U20211 (N_20211,N_18006,N_19873);
nand U20212 (N_20212,N_19697,N_18484);
nand U20213 (N_20213,N_18514,N_19686);
and U20214 (N_20214,N_18909,N_19376);
and U20215 (N_20215,N_18410,N_18695);
nor U20216 (N_20216,N_18566,N_18707);
nor U20217 (N_20217,N_19921,N_18015);
nand U20218 (N_20218,N_19656,N_18312);
xor U20219 (N_20219,N_19755,N_19989);
or U20220 (N_20220,N_18873,N_18249);
xnor U20221 (N_20221,N_19524,N_19282);
nand U20222 (N_20222,N_18308,N_19060);
nand U20223 (N_20223,N_19265,N_19339);
xor U20224 (N_20224,N_19294,N_19497);
xnor U20225 (N_20225,N_19739,N_19479);
xor U20226 (N_20226,N_18084,N_18302);
nand U20227 (N_20227,N_18103,N_19349);
or U20228 (N_20228,N_18740,N_19366);
xor U20229 (N_20229,N_19639,N_18480);
or U20230 (N_20230,N_19757,N_18077);
nand U20231 (N_20231,N_18288,N_18951);
xnor U20232 (N_20232,N_18810,N_18919);
and U20233 (N_20233,N_19771,N_18114);
nand U20234 (N_20234,N_19180,N_19531);
and U20235 (N_20235,N_18806,N_18173);
nor U20236 (N_20236,N_18096,N_18849);
nor U20237 (N_20237,N_18481,N_18956);
or U20238 (N_20238,N_18150,N_19407);
and U20239 (N_20239,N_18958,N_18735);
xnor U20240 (N_20240,N_18688,N_18239);
xor U20241 (N_20241,N_19106,N_19835);
and U20242 (N_20242,N_18503,N_18263);
xor U20243 (N_20243,N_18456,N_18137);
and U20244 (N_20244,N_19214,N_19457);
and U20245 (N_20245,N_18942,N_19974);
nor U20246 (N_20246,N_19649,N_18088);
and U20247 (N_20247,N_19978,N_18631);
nand U20248 (N_20248,N_19775,N_19532);
or U20249 (N_20249,N_18172,N_19122);
and U20250 (N_20250,N_19953,N_18408);
nor U20251 (N_20251,N_18295,N_18839);
or U20252 (N_20252,N_19789,N_18053);
nor U20253 (N_20253,N_18422,N_18929);
nand U20254 (N_20254,N_18930,N_18065);
and U20255 (N_20255,N_19179,N_19562);
or U20256 (N_20256,N_18539,N_19160);
nor U20257 (N_20257,N_18976,N_18544);
xnor U20258 (N_20258,N_19726,N_18125);
or U20259 (N_20259,N_19099,N_19551);
nand U20260 (N_20260,N_18460,N_18363);
nand U20261 (N_20261,N_19143,N_19442);
or U20262 (N_20262,N_19408,N_19120);
or U20263 (N_20263,N_18734,N_18339);
xnor U20264 (N_20264,N_19046,N_19960);
or U20265 (N_20265,N_19161,N_18453);
xor U20266 (N_20266,N_19618,N_19598);
xor U20267 (N_20267,N_19228,N_18933);
nor U20268 (N_20268,N_18443,N_19700);
nand U20269 (N_20269,N_19322,N_19675);
xor U20270 (N_20270,N_18624,N_19807);
and U20271 (N_20271,N_18507,N_19541);
nand U20272 (N_20272,N_19827,N_19890);
xnor U20273 (N_20273,N_18505,N_19146);
nor U20274 (N_20274,N_19257,N_19991);
nor U20275 (N_20275,N_19448,N_19706);
nor U20276 (N_20276,N_18297,N_19865);
nand U20277 (N_20277,N_19522,N_18558);
or U20278 (N_20278,N_19582,N_18033);
xor U20279 (N_20279,N_18769,N_18026);
nor U20280 (N_20280,N_18298,N_18556);
nand U20281 (N_20281,N_19548,N_19335);
xnor U20282 (N_20282,N_19417,N_19910);
and U20283 (N_20283,N_18402,N_19801);
nor U20284 (N_20284,N_18483,N_18184);
or U20285 (N_20285,N_18042,N_19138);
nand U20286 (N_20286,N_18143,N_19836);
xnor U20287 (N_20287,N_19510,N_18941);
or U20288 (N_20288,N_19164,N_19471);
xor U20289 (N_20289,N_19220,N_19221);
xnor U20290 (N_20290,N_19102,N_18540);
or U20291 (N_20291,N_18542,N_18801);
or U20292 (N_20292,N_18393,N_18477);
nand U20293 (N_20293,N_18917,N_19704);
nor U20294 (N_20294,N_18927,N_19191);
nand U20295 (N_20295,N_18680,N_19934);
nor U20296 (N_20296,N_19804,N_18023);
nand U20297 (N_20297,N_18579,N_18984);
or U20298 (N_20298,N_19280,N_18140);
nand U20299 (N_20299,N_18616,N_18783);
nand U20300 (N_20300,N_19875,N_18455);
nand U20301 (N_20301,N_19435,N_19188);
or U20302 (N_20302,N_19456,N_18602);
nor U20303 (N_20303,N_18776,N_19420);
nor U20304 (N_20304,N_18198,N_18357);
nand U20305 (N_20305,N_18538,N_18699);
or U20306 (N_20306,N_18716,N_18645);
xnor U20307 (N_20307,N_19939,N_19481);
or U20308 (N_20308,N_19746,N_18168);
and U20309 (N_20309,N_18755,N_18596);
xnor U20310 (N_20310,N_18113,N_19545);
and U20311 (N_20311,N_19837,N_19330);
or U20312 (N_20312,N_19447,N_18940);
nand U20313 (N_20313,N_18612,N_19595);
and U20314 (N_20314,N_18620,N_19702);
and U20315 (N_20315,N_19915,N_18265);
nand U20316 (N_20316,N_19990,N_19646);
xnor U20317 (N_20317,N_19925,N_18030);
and U20318 (N_20318,N_18692,N_19779);
xor U20319 (N_20319,N_18466,N_18176);
xnor U20320 (N_20320,N_19284,N_19462);
and U20321 (N_20321,N_19825,N_18160);
or U20322 (N_20322,N_19367,N_18727);
and U20323 (N_20323,N_19657,N_18279);
xnor U20324 (N_20324,N_19955,N_18521);
or U20325 (N_20325,N_18788,N_18728);
or U20326 (N_20326,N_18290,N_19519);
xor U20327 (N_20327,N_19967,N_18913);
nor U20328 (N_20328,N_19454,N_18419);
nand U20329 (N_20329,N_19303,N_19912);
nand U20330 (N_20330,N_19154,N_18253);
or U20331 (N_20331,N_18044,N_19014);
or U20332 (N_20332,N_18732,N_19411);
or U20333 (N_20333,N_19520,N_18567);
and U20334 (N_20334,N_18350,N_19636);
or U20335 (N_20335,N_19058,N_18412);
nor U20336 (N_20336,N_19119,N_19833);
and U20337 (N_20337,N_18630,N_19321);
xnor U20338 (N_20338,N_18209,N_19387);
nor U20339 (N_20339,N_18733,N_18179);
and U20340 (N_20340,N_18148,N_18237);
or U20341 (N_20341,N_18205,N_18195);
nor U20342 (N_20342,N_18510,N_19949);
or U20343 (N_20343,N_18577,N_18513);
xor U20344 (N_20344,N_18391,N_19816);
nor U20345 (N_20345,N_19662,N_19168);
nand U20346 (N_20346,N_18872,N_18347);
nor U20347 (N_20347,N_19150,N_18987);
nor U20348 (N_20348,N_19437,N_18731);
and U20349 (N_20349,N_19293,N_19129);
or U20350 (N_20350,N_18272,N_18802);
or U20351 (N_20351,N_19874,N_19576);
or U20352 (N_20352,N_18617,N_19012);
xnor U20353 (N_20353,N_18025,N_19005);
or U20354 (N_20354,N_19347,N_19226);
nor U20355 (N_20355,N_19786,N_19302);
and U20356 (N_20356,N_19985,N_18523);
nor U20357 (N_20357,N_18452,N_18574);
nor U20358 (N_20358,N_18365,N_19822);
and U20359 (N_20359,N_19108,N_19325);
and U20360 (N_20360,N_18867,N_18409);
or U20361 (N_20361,N_19577,N_19449);
xor U20362 (N_20362,N_19252,N_19105);
or U20363 (N_20363,N_19213,N_18395);
nand U20364 (N_20364,N_18451,N_19988);
and U20365 (N_20365,N_19247,N_19475);
and U20366 (N_20366,N_18394,N_18623);
and U20367 (N_20367,N_19785,N_19927);
xor U20368 (N_20368,N_18441,N_18648);
and U20369 (N_20369,N_18967,N_19503);
xnor U20370 (N_20370,N_19902,N_19039);
nor U20371 (N_20371,N_19218,N_19869);
nor U20372 (N_20372,N_18764,N_19787);
nand U20373 (N_20373,N_18582,N_19429);
or U20374 (N_20374,N_19260,N_18211);
nand U20375 (N_20375,N_19705,N_19195);
and U20376 (N_20376,N_19561,N_19197);
or U20377 (N_20377,N_19752,N_19472);
or U20378 (N_20378,N_18685,N_18317);
nand U20379 (N_20379,N_19315,N_18899);
nor U20380 (N_20380,N_18673,N_19631);
nor U20381 (N_20381,N_19288,N_18957);
xnor U20382 (N_20382,N_19625,N_19619);
nand U20383 (N_20383,N_19664,N_18382);
or U20384 (N_20384,N_19359,N_19116);
nor U20385 (N_20385,N_18262,N_18693);
nor U20386 (N_20386,N_19224,N_18062);
xnor U20387 (N_20387,N_18335,N_18156);
or U20388 (N_20388,N_19211,N_18001);
and U20389 (N_20389,N_19259,N_18895);
xor U20390 (N_20390,N_19819,N_19067);
nor U20391 (N_20391,N_18974,N_18375);
nor U20392 (N_20392,N_19682,N_19521);
nand U20393 (N_20393,N_19467,N_19883);
nand U20394 (N_20394,N_19064,N_18715);
nor U20395 (N_20395,N_18778,N_18250);
and U20396 (N_20396,N_18051,N_18532);
nor U20397 (N_20397,N_19579,N_18492);
nor U20398 (N_20398,N_18879,N_18811);
nand U20399 (N_20399,N_19422,N_19964);
nor U20400 (N_20400,N_19882,N_19078);
nor U20401 (N_20401,N_19745,N_19151);
or U20402 (N_20402,N_18625,N_19423);
nor U20403 (N_20403,N_18283,N_19149);
and U20404 (N_20404,N_18427,N_18276);
or U20405 (N_20405,N_19140,N_18098);
nor U20406 (N_20406,N_19035,N_19396);
xnor U20407 (N_20407,N_18918,N_19941);
xor U20408 (N_20408,N_19095,N_19728);
xnor U20409 (N_20409,N_18180,N_18552);
and U20410 (N_20410,N_18122,N_18085);
nor U20411 (N_20411,N_19893,N_19049);
and U20412 (N_20412,N_18213,N_18812);
and U20413 (N_20413,N_19478,N_18932);
nor U20414 (N_20414,N_19490,N_18530);
nor U20415 (N_20415,N_19076,N_18562);
xor U20416 (N_20416,N_18206,N_19671);
nor U20417 (N_20417,N_19017,N_19845);
xor U20418 (N_20418,N_19225,N_19975);
and U20419 (N_20419,N_18116,N_19425);
nor U20420 (N_20420,N_19077,N_18814);
and U20421 (N_20421,N_19145,N_19352);
nand U20422 (N_20422,N_18144,N_19633);
xor U20423 (N_20423,N_18301,N_19267);
nand U20424 (N_20424,N_19201,N_18876);
or U20425 (N_20425,N_19792,N_19868);
nor U20426 (N_20426,N_18241,N_18889);
xnor U20427 (N_20427,N_19069,N_18960);
xnor U20428 (N_20428,N_19283,N_18609);
nand U20429 (N_20429,N_19832,N_18722);
nand U20430 (N_20430,N_18857,N_19621);
and U20431 (N_20431,N_18397,N_19606);
and U20432 (N_20432,N_19234,N_19446);
nor U20433 (N_20433,N_18534,N_19716);
xor U20434 (N_20434,N_18723,N_19672);
xnor U20435 (N_20435,N_19433,N_18474);
nor U20436 (N_20436,N_18533,N_19192);
nor U20437 (N_20437,N_19484,N_18229);
nor U20438 (N_20438,N_19765,N_19275);
nor U20439 (N_20439,N_19341,N_19546);
xor U20440 (N_20440,N_18461,N_18177);
and U20441 (N_20441,N_19670,N_18193);
or U20442 (N_20442,N_19178,N_19555);
and U20443 (N_20443,N_18832,N_18498);
nand U20444 (N_20444,N_19620,N_18914);
nor U20445 (N_20445,N_18860,N_18002);
and U20446 (N_20446,N_19476,N_18892);
nand U20447 (N_20447,N_18928,N_18823);
nand U20448 (N_20448,N_18654,N_19445);
xor U20449 (N_20449,N_19977,N_18182);
nand U20450 (N_20450,N_18896,N_18081);
nand U20451 (N_20451,N_19274,N_18170);
nor U20452 (N_20452,N_19209,N_18751);
xnor U20453 (N_20453,N_19652,N_18031);
nand U20454 (N_20454,N_18490,N_19867);
nor U20455 (N_20455,N_18489,N_19851);
nor U20456 (N_20456,N_19107,N_19051);
nand U20457 (N_20457,N_18721,N_19065);
nor U20458 (N_20458,N_19648,N_18550);
xor U20459 (N_20459,N_18012,N_18017);
or U20460 (N_20460,N_19100,N_18963);
and U20461 (N_20461,N_19324,N_19971);
and U20462 (N_20462,N_18493,N_19876);
xor U20463 (N_20463,N_19679,N_19928);
nand U20464 (N_20464,N_19914,N_18664);
nor U20465 (N_20465,N_18682,N_19232);
nand U20466 (N_20466,N_19235,N_19944);
nor U20467 (N_20467,N_18501,N_18511);
xor U20468 (N_20468,N_19299,N_18362);
nand U20469 (N_20469,N_18908,N_19430);
or U20470 (N_20470,N_18569,N_19713);
xnor U20471 (N_20471,N_18856,N_18320);
nand U20472 (N_20472,N_19808,N_19655);
and U20473 (N_20473,N_18155,N_18975);
nor U20474 (N_20474,N_18021,N_19952);
and U20475 (N_20475,N_19849,N_19127);
and U20476 (N_20476,N_19243,N_19200);
and U20477 (N_20477,N_19536,N_19610);
and U20478 (N_20478,N_19908,N_18303);
nor U20479 (N_20479,N_18756,N_18646);
nor U20480 (N_20480,N_18982,N_18635);
nand U20481 (N_20481,N_18171,N_18436);
nand U20482 (N_20482,N_18512,N_18555);
xor U20483 (N_20483,N_19820,N_19761);
nand U20484 (N_20484,N_19604,N_19306);
nand U20485 (N_20485,N_18066,N_19163);
nand U20486 (N_20486,N_18804,N_18175);
xnor U20487 (N_20487,N_18330,N_19270);
nand U20488 (N_20488,N_19698,N_18998);
nor U20489 (N_20489,N_18718,N_19913);
nor U20490 (N_20490,N_18476,N_19183);
xnor U20491 (N_20491,N_18189,N_19578);
and U20492 (N_20492,N_18668,N_19297);
nor U20493 (N_20493,N_19564,N_19452);
and U20494 (N_20494,N_18658,N_19405);
nor U20495 (N_20495,N_18844,N_18547);
nor U20496 (N_20496,N_18161,N_18995);
nand U20497 (N_20497,N_18127,N_19055);
and U20498 (N_20498,N_18861,N_19434);
nand U20499 (N_20499,N_18311,N_19938);
nand U20500 (N_20500,N_18126,N_19590);
xnor U20501 (N_20501,N_18417,N_19040);
nor U20502 (N_20502,N_19215,N_19858);
and U20503 (N_20503,N_18647,N_18361);
or U20504 (N_20504,N_19015,N_18827);
or U20505 (N_20505,N_19233,N_19569);
or U20506 (N_20506,N_18924,N_19591);
nand U20507 (N_20507,N_18425,N_18822);
and U20508 (N_20508,N_18864,N_18970);
xnor U20509 (N_20509,N_19599,N_19586);
or U20510 (N_20510,N_19372,N_19653);
and U20511 (N_20511,N_19782,N_19473);
xor U20512 (N_20512,N_19459,N_18931);
nor U20513 (N_20513,N_19222,N_18705);
xnor U20514 (N_20514,N_19922,N_19432);
and U20515 (N_20515,N_18226,N_19353);
nand U20516 (N_20516,N_19568,N_18254);
xnor U20517 (N_20517,N_18576,N_18519);
or U20518 (N_20518,N_19635,N_19998);
nand U20519 (N_20519,N_18003,N_18121);
or U20520 (N_20520,N_18826,N_19394);
and U20521 (N_20521,N_19389,N_18067);
or U20522 (N_20522,N_19428,N_19715);
or U20523 (N_20523,N_18216,N_18080);
xor U20524 (N_20524,N_19170,N_18159);
or U20525 (N_20525,N_19754,N_19528);
or U20526 (N_20526,N_18906,N_19919);
nand U20527 (N_20527,N_18659,N_18465);
xnor U20528 (N_20528,N_19223,N_18518);
nor U20529 (N_20529,N_18454,N_18458);
nand U20530 (N_20530,N_19684,N_18497);
or U20531 (N_20531,N_18420,N_18369);
or U20532 (N_20532,N_19717,N_19346);
or U20533 (N_20533,N_19862,N_18591);
xnor U20534 (N_20534,N_18197,N_18400);
nor U20535 (N_20535,N_18130,N_19565);
or U20536 (N_20536,N_18273,N_18628);
or U20537 (N_20537,N_18563,N_19409);
nor U20538 (N_20538,N_18457,N_19371);
xnor U20539 (N_20539,N_18352,N_18194);
or U20540 (N_20540,N_19320,N_19489);
nand U20541 (N_20541,N_19157,N_18837);
xor U20542 (N_20542,N_19995,N_19169);
or U20543 (N_20543,N_19641,N_18966);
nor U20544 (N_20544,N_18321,N_18281);
xnor U20545 (N_20545,N_19258,N_19466);
or U20546 (N_20546,N_18087,N_18679);
nand U20547 (N_20547,N_19318,N_18313);
or U20548 (N_20548,N_18977,N_19916);
nor U20549 (N_20549,N_19947,N_19718);
xnor U20550 (N_20550,N_18959,N_19720);
and U20551 (N_20551,N_19759,N_19943);
nor U20552 (N_20552,N_19074,N_18435);
xnor U20553 (N_20553,N_19508,N_18786);
xor U20554 (N_20554,N_18355,N_19021);
nor U20555 (N_20555,N_18310,N_18275);
and U20556 (N_20556,N_18613,N_18798);
nand U20557 (N_20557,N_19128,N_19374);
or U20558 (N_20558,N_19443,N_18719);
nand U20559 (N_20559,N_19033,N_18655);
nand U20560 (N_20560,N_18842,N_18190);
nor U20561 (N_20561,N_19043,N_19622);
and U20562 (N_20562,N_18912,N_19378);
nor U20563 (N_20563,N_19027,N_18287);
and U20564 (N_20564,N_18592,N_18604);
or U20565 (N_20565,N_18606,N_18459);
xnor U20566 (N_20566,N_19643,N_18107);
nor U20567 (N_20567,N_18792,N_18702);
and U20568 (N_20568,N_18005,N_18554);
or U20569 (N_20569,N_19311,N_19460);
nor U20570 (N_20570,N_18866,N_18762);
and U20571 (N_20571,N_19314,N_19010);
nor U20572 (N_20572,N_19091,N_18404);
nor U20573 (N_20573,N_19707,N_18601);
xor U20574 (N_20574,N_19217,N_19803);
nor U20575 (N_20575,N_19547,N_18978);
nor U20576 (N_20576,N_18368,N_18019);
and U20577 (N_20577,N_19198,N_18095);
and U20578 (N_20578,N_19384,N_19756);
xnor U20579 (N_20579,N_19126,N_18299);
nor U20580 (N_20580,N_18423,N_19121);
and U20581 (N_20581,N_19401,N_19879);
and U20582 (N_20582,N_19455,N_19897);
and U20583 (N_20583,N_18657,N_19558);
or U20584 (N_20584,N_19139,N_18323);
xor U20585 (N_20585,N_19514,N_19155);
and U20586 (N_20586,N_18414,N_18499);
nand U20587 (N_20587,N_19504,N_18145);
and U20588 (N_20588,N_19727,N_18819);
and U20589 (N_20589,N_18090,N_19421);
nor U20590 (N_20590,N_19024,N_18992);
nand U20591 (N_20591,N_18850,N_18034);
xnor U20592 (N_20592,N_18075,N_19227);
and U20593 (N_20593,N_19053,N_18413);
xnor U20594 (N_20594,N_19397,N_18230);
nand U20595 (N_20595,N_18997,N_18151);
xor U20596 (N_20596,N_19581,N_19189);
xnor U20597 (N_20597,N_18996,N_18590);
nor U20598 (N_20598,N_18749,N_18133);
nand U20599 (N_20599,N_18024,N_18169);
and U20600 (N_20600,N_19329,N_19263);
xor U20601 (N_20601,N_18973,N_18282);
xnor U20602 (N_20602,N_18717,N_18780);
and U20603 (N_20603,N_19296,N_19554);
nor U20604 (N_20604,N_19632,N_19333);
or U20605 (N_20605,N_18656,N_18840);
nor U20606 (N_20606,N_19465,N_19385);
or U20607 (N_20607,N_18853,N_18407);
xor U20608 (N_20608,N_19507,N_18039);
xor U20609 (N_20609,N_18385,N_19167);
xor U20610 (N_20610,N_19553,N_19093);
nor U20611 (N_20611,N_18201,N_18639);
nand U20612 (N_20612,N_19388,N_18529);
and U20613 (N_20613,N_19261,N_19674);
nor U20614 (N_20614,N_18208,N_18911);
nand U20615 (N_20615,N_19735,N_18687);
and U20616 (N_20616,N_19603,N_19823);
nand U20617 (N_20617,N_18491,N_19063);
or U20618 (N_20618,N_18504,N_19530);
or U20619 (N_20619,N_19959,N_19888);
nand U20620 (N_20620,N_19777,N_19594);
nand U20621 (N_20621,N_19111,N_18662);
xnor U20622 (N_20622,N_18938,N_18332);
and U20623 (N_20623,N_19499,N_18653);
or U20624 (N_20624,N_18730,N_19023);
nor U20625 (N_20625,N_19525,N_19918);
nor U20626 (N_20626,N_18073,N_18428);
or U20627 (N_20627,N_18188,N_19962);
nor U20628 (N_20628,N_19031,N_18101);
xor U20629 (N_20629,N_19144,N_19413);
nor U20630 (N_20630,N_19326,N_18752);
and U20631 (N_20631,N_18570,N_18046);
nor U20632 (N_20632,N_19799,N_19588);
nor U20633 (N_20633,N_19710,N_18200);
nand U20634 (N_20634,N_18667,N_18218);
and U20635 (N_20635,N_18891,N_18210);
xor U20636 (N_20636,N_19906,N_19904);
and U20637 (N_20637,N_18136,N_18354);
nor U20638 (N_20638,N_19148,N_19535);
xnor U20639 (N_20639,N_19979,N_18520);
nor U20640 (N_20640,N_19711,N_19794);
xor U20641 (N_20641,N_19348,N_19250);
or U20642 (N_20642,N_18672,N_19301);
or U20643 (N_20643,N_18683,N_18337);
and U20644 (N_20644,N_19640,N_19047);
and U20645 (N_20645,N_18830,N_19287);
and U20646 (N_20646,N_19886,N_18475);
xor U20647 (N_20647,N_18528,N_18286);
nand U20648 (N_20648,N_18817,N_18104);
and U20649 (N_20649,N_18704,N_19946);
nor U20650 (N_20650,N_18920,N_18744);
nand U20651 (N_20651,N_19950,N_18548);
xor U20652 (N_20652,N_18946,N_18146);
nor U20653 (N_20653,N_19956,N_18326);
or U20654 (N_20654,N_18586,N_19714);
and U20655 (N_20655,N_19312,N_18907);
xor U20656 (N_20656,N_18578,N_19343);
nor U20657 (N_20657,N_19207,N_19885);
and U20658 (N_20658,N_19182,N_18219);
nor U20659 (N_20659,N_19036,N_18708);
and U20660 (N_20660,N_19784,N_18750);
nand U20661 (N_20661,N_18004,N_19450);
nor U20662 (N_20662,N_18037,N_19612);
and U20663 (N_20663,N_19791,N_18196);
xor U20664 (N_20664,N_19370,N_19766);
nor U20665 (N_20665,N_19176,N_18777);
nand U20666 (N_20666,N_19184,N_18985);
or U20667 (N_20667,N_19439,N_18345);
or U20668 (N_20668,N_19073,N_19768);
and U20669 (N_20669,N_18611,N_19911);
and U20670 (N_20670,N_18424,N_19935);
and U20671 (N_20671,N_19136,N_19295);
xor U20672 (N_20672,N_19650,N_18779);
or U20673 (N_20673,N_19086,N_18902);
xnor U20674 (N_20674,N_19589,N_18568);
xnor U20675 (N_20675,N_19983,N_18666);
and U20676 (N_20676,N_19831,N_19940);
xnor U20677 (N_20677,N_19350,N_18926);
and U20678 (N_20678,N_19045,N_19511);
and U20679 (N_20679,N_18325,N_18619);
and U20680 (N_20680,N_19239,N_18167);
xnor U20681 (N_20681,N_18838,N_19894);
or U20682 (N_20682,N_19050,N_19617);
or U20683 (N_20683,N_19468,N_18709);
or U20684 (N_20684,N_18079,N_19355);
and U20685 (N_20685,N_18470,N_18115);
nand U20686 (N_20686,N_19571,N_19491);
nor U20687 (N_20687,N_18482,N_18972);
or U20688 (N_20688,N_19085,N_18040);
nand U20689 (N_20689,N_18527,N_18990);
and U20690 (N_20690,N_18013,N_18434);
xor U20691 (N_20691,N_18858,N_19665);
and U20692 (N_20692,N_18881,N_18344);
nand U20693 (N_20693,N_19251,N_19079);
xor U20694 (N_20694,N_18684,N_18690);
or U20695 (N_20695,N_19001,N_19742);
nor U20696 (N_20696,N_18950,N_19666);
and U20697 (N_20697,N_19690,N_18761);
or U20698 (N_20698,N_19156,N_19932);
and U20699 (N_20699,N_18949,N_19291);
nand U20700 (N_20700,N_18691,N_19236);
or U20701 (N_20701,N_18748,N_19593);
nor U20702 (N_20702,N_18022,N_19402);
and U20703 (N_20703,N_19689,N_18636);
and U20704 (N_20704,N_18980,N_18050);
nor U20705 (N_20705,N_19800,N_18496);
xnor U20706 (N_20706,N_19624,N_18669);
nand U20707 (N_20707,N_19627,N_19237);
or U20708 (N_20708,N_19132,N_19334);
nand U20709 (N_20709,N_19847,N_19248);
nand U20710 (N_20710,N_19492,N_19924);
and U20711 (N_20711,N_19826,N_19602);
xnor U20712 (N_20712,N_18112,N_19109);
xnor U20713 (N_20713,N_19501,N_18319);
xnor U20714 (N_20714,N_18398,N_19317);
nor U20715 (N_20715,N_19242,N_19933);
nor U20716 (N_20716,N_18440,N_18781);
or U20717 (N_20717,N_18874,N_18338);
or U20718 (N_20718,N_18545,N_18854);
nand U20719 (N_20719,N_18300,N_19137);
nand U20720 (N_20720,N_18736,N_18608);
nand U20721 (N_20721,N_18266,N_19680);
and U20722 (N_20722,N_19986,N_18228);
or U20723 (N_20723,N_19814,N_19889);
and U20724 (N_20724,N_19601,N_18124);
nor U20725 (N_20725,N_18627,N_18260);
nor U20726 (N_20726,N_19813,N_18356);
nand U20727 (N_20727,N_18010,N_18248);
and U20728 (N_20728,N_19469,N_19769);
or U20729 (N_20729,N_18094,N_19628);
xor U20730 (N_20730,N_18389,N_18267);
or U20731 (N_20731,N_19375,N_18789);
or U20732 (N_20732,N_18448,N_19286);
xnor U20733 (N_20733,N_18626,N_18790);
nor U20734 (N_20734,N_18469,N_18865);
nand U20735 (N_20735,N_19307,N_18859);
nand U20736 (N_20736,N_19651,N_18988);
xor U20737 (N_20737,N_18772,N_19748);
or U20738 (N_20738,N_18726,N_19313);
or U20739 (N_20739,N_18054,N_18360);
xor U20740 (N_20740,N_19038,N_18132);
nor U20741 (N_20741,N_18675,N_19527);
or U20742 (N_20742,N_19795,N_19654);
nor U20743 (N_20743,N_19483,N_19451);
xor U20744 (N_20744,N_18047,N_19544);
nor U20745 (N_20745,N_18011,N_19171);
nand U20746 (N_20746,N_18343,N_18573);
and U20747 (N_20747,N_18191,N_19072);
and U20748 (N_20748,N_19203,N_18953);
or U20749 (N_20749,N_19751,N_19515);
nor U20750 (N_20750,N_18333,N_19901);
nor U20751 (N_20751,N_19892,N_19373);
nor U20752 (N_20752,N_18035,N_18841);
xnor U20753 (N_20753,N_18760,N_19241);
nor U20754 (N_20754,N_19377,N_18877);
xnor U20755 (N_20755,N_19658,N_19009);
nor U20756 (N_20756,N_18700,N_18439);
or U20757 (N_20757,N_18437,N_19723);
or U20758 (N_20758,N_18032,N_18069);
xnor U20759 (N_20759,N_18910,N_18809);
xnor U20760 (N_20760,N_19084,N_18524);
or U20761 (N_20761,N_18089,N_19958);
xnor U20762 (N_20762,N_19269,N_19029);
or U20763 (N_20763,N_19592,N_19896);
nor U20764 (N_20764,N_19763,N_19101);
or U20765 (N_20765,N_19694,N_18921);
nor U20766 (N_20766,N_18852,N_18661);
xor U20767 (N_20767,N_19369,N_19300);
nand U20768 (N_20768,N_19493,N_18767);
or U20769 (N_20769,N_18280,N_18119);
nand U20770 (N_20770,N_19774,N_19708);
nand U20771 (N_20771,N_18246,N_18559);
nor U20772 (N_20772,N_19404,N_19750);
nand U20773 (N_20773,N_19966,N_18027);
or U20774 (N_20774,N_19266,N_18581);
and U20775 (N_20775,N_18575,N_18508);
nor U20776 (N_20776,N_19563,N_18141);
nor U20777 (N_20777,N_19185,N_18029);
or U20778 (N_20778,N_19278,N_18526);
nor U20779 (N_20779,N_19174,N_19669);
xnor U20780 (N_20780,N_18793,N_19846);
nand U20781 (N_20781,N_18243,N_18763);
xor U20782 (N_20782,N_18334,N_18433);
nand U20783 (N_20783,N_19920,N_18468);
and U20784 (N_20784,N_18294,N_18142);
or U20785 (N_20785,N_18961,N_18833);
nor U20786 (N_20786,N_18805,N_19663);
xnor U20787 (N_20787,N_19982,N_18935);
or U20788 (N_20788,N_19608,N_18370);
and U20789 (N_20789,N_18236,N_19976);
xnor U20790 (N_20790,N_18807,N_18045);
and U20791 (N_20791,N_18048,N_19645);
or U20792 (N_20792,N_19319,N_19994);
and U20793 (N_20793,N_18824,N_19354);
nand U20794 (N_20794,N_19204,N_19323);
nor U20795 (N_20795,N_18367,N_18247);
xor U20796 (N_20796,N_19824,N_18597);
nand U20797 (N_20797,N_18981,N_19480);
nor U20798 (N_20798,N_18128,N_19505);
or U20799 (N_20799,N_18632,N_19004);
and U20800 (N_20800,N_18993,N_19996);
and U20801 (N_20801,N_18808,N_18183);
xor U20802 (N_20802,N_18948,N_19020);
xor U20803 (N_20803,N_18815,N_18203);
or U20804 (N_20804,N_19246,N_18697);
nor U20805 (N_20805,N_19516,N_18737);
nand U20806 (N_20806,N_19358,N_18220);
xnor U20807 (N_20807,N_19486,N_19626);
nand U20808 (N_20808,N_19980,N_18309);
xor U20809 (N_20809,N_19973,N_18214);
nor U20810 (N_20810,N_18759,N_18372);
and U20811 (N_20811,N_19496,N_19676);
xnor U20812 (N_20812,N_18698,N_19338);
nor U20813 (N_20813,N_19709,N_19984);
nand U20814 (N_20814,N_19464,N_18836);
and U20815 (N_20815,N_18818,N_18364);
and U20816 (N_20816,N_19526,N_18870);
xnor U20817 (N_20817,N_18060,N_19724);
nor U20818 (N_20818,N_18322,N_19068);
nor U20819 (N_20819,N_19972,N_19474);
and U20820 (N_20820,N_18593,N_19970);
xor U20821 (N_20821,N_19880,N_18390);
xor U20822 (N_20822,N_19781,N_18599);
nor U20823 (N_20823,N_18117,N_18607);
and U20824 (N_20824,N_19930,N_18061);
nand U20825 (N_20825,N_18384,N_19523);
nand U20826 (N_20826,N_19412,N_19123);
and U20827 (N_20827,N_19166,N_19722);
xor U20828 (N_20828,N_19007,N_19256);
or U20829 (N_20829,N_19498,N_18515);
nor U20830 (N_20830,N_19719,N_19843);
and U20831 (N_20831,N_18123,N_18255);
nor U20832 (N_20832,N_18901,N_18546);
or U20833 (N_20833,N_18883,N_18903);
xnor U20834 (N_20834,N_18274,N_19316);
xor U20835 (N_20835,N_18192,N_18820);
nor U20836 (N_20836,N_18429,N_19637);
or U20837 (N_20837,N_18829,N_19271);
and U20838 (N_20838,N_19186,N_18432);
and U20839 (N_20839,N_19929,N_18346);
nor U20840 (N_20840,N_19818,N_18374);
nor U20841 (N_20841,N_19575,N_19556);
nor U20842 (N_20842,N_19760,N_19135);
and U20843 (N_20843,N_18318,N_19196);
or U20844 (N_20844,N_19056,N_19533);
or U20845 (N_20845,N_19131,N_19878);
nand U20846 (N_20846,N_19693,N_19534);
nor U20847 (N_20847,N_19208,N_18038);
nand U20848 (N_20848,N_19175,N_18093);
nand U20849 (N_20849,N_19500,N_19917);
nor U20850 (N_20850,N_19057,N_19877);
xor U20851 (N_20851,N_19743,N_19368);
and U20852 (N_20852,N_18768,N_18009);
and U20853 (N_20853,N_18848,N_18178);
or U20854 (N_20854,N_18845,N_18232);
nor U20855 (N_20855,N_18954,N_19253);
xnor U20856 (N_20856,N_19229,N_19729);
nor U20857 (N_20857,N_18215,N_19018);
xor U20858 (N_20858,N_18296,N_18105);
and U20859 (N_20859,N_18663,N_18676);
nand U20860 (N_20860,N_19262,N_18887);
and U20861 (N_20861,N_18791,N_19361);
or U20862 (N_20862,N_18706,N_19659);
xor U20863 (N_20863,N_18381,N_19557);
or U20864 (N_20864,N_18392,N_18863);
or U20865 (N_20865,N_19264,N_19688);
or U20866 (N_20866,N_19495,N_18158);
or U20867 (N_20867,N_18541,N_19344);
or U20868 (N_20868,N_19573,N_19310);
and U20869 (N_20869,N_19097,N_19642);
xnor U20870 (N_20870,N_19273,N_19390);
or U20871 (N_20871,N_19360,N_19392);
nor U20872 (N_20872,N_18083,N_18487);
or U20873 (N_20873,N_18411,N_19485);
and U20874 (N_20874,N_19725,N_19969);
nor U20875 (N_20875,N_18595,N_19298);
or U20876 (N_20876,N_19414,N_19699);
and U20877 (N_20877,N_18058,N_18478);
or U20878 (N_20878,N_18129,N_18327);
nor U20879 (N_20879,N_18923,N_19623);
or U20880 (N_20880,N_19406,N_19783);
and U20881 (N_20881,N_18915,N_18795);
or U20882 (N_20882,N_18406,N_18603);
nand U20883 (N_20883,N_18186,N_19308);
nor U20884 (N_20884,N_18082,N_18652);
nand U20885 (N_20885,N_18766,N_19030);
and U20886 (N_20886,N_18258,N_19738);
nor U20887 (N_20887,N_19153,N_19542);
nor U20888 (N_20888,N_19863,N_19762);
or U20889 (N_20889,N_18885,N_19383);
nand U20890 (N_20890,N_18561,N_18979);
and U20891 (N_20891,N_18774,N_18905);
xor U20892 (N_20892,N_19309,N_18162);
or U20893 (N_20893,N_19276,N_19903);
xnor U20894 (N_20894,N_19905,N_18994);
nand U20895 (N_20895,N_19550,N_18418);
xnor U20896 (N_20896,N_18689,N_19436);
nand U20897 (N_20897,N_19199,N_18486);
xor U20898 (N_20898,N_19080,N_19673);
nor U20899 (N_20899,N_19834,N_19231);
or U20900 (N_20900,N_18565,N_18882);
nand U20901 (N_20901,N_19019,N_18064);
xor U20902 (N_20902,N_18771,N_19124);
nand U20903 (N_20903,N_19393,N_19721);
or U20904 (N_20904,N_19987,N_19070);
nand U20905 (N_20905,N_19115,N_18278);
xor U20906 (N_20906,N_19812,N_18388);
nor U20907 (N_20907,N_18964,N_19011);
and U20908 (N_20908,N_19749,N_19740);
or U20909 (N_20909,N_18000,N_19881);
xor U20910 (N_20910,N_18834,N_18729);
nor U20911 (N_20911,N_19730,N_18264);
nand U20912 (N_20912,N_18277,N_19272);
nor U20913 (N_20913,N_19075,N_19285);
or U20914 (N_20914,N_18238,N_19381);
nor U20915 (N_20915,N_19362,N_19365);
xnor U20916 (N_20916,N_18537,N_18118);
nor U20917 (N_20917,N_19854,N_19002);
xnor U20918 (N_20918,N_19853,N_18373);
nor U20919 (N_20919,N_19790,N_19281);
nand U20920 (N_20920,N_18305,N_18328);
nor U20921 (N_20921,N_18100,N_19345);
and U20922 (N_20922,N_18738,N_18380);
nand U20923 (N_20923,N_18348,N_19809);
or U20924 (N_20924,N_18259,N_18261);
nand U20925 (N_20925,N_19855,N_18108);
nand U20926 (N_20926,N_18307,N_19583);
nor U20927 (N_20927,N_18965,N_19572);
or U20928 (N_20928,N_19616,N_19963);
nor U20929 (N_20929,N_19584,N_18401);
xor U20930 (N_20930,N_19022,N_19614);
xnor U20931 (N_20931,N_18671,N_18615);
and U20932 (N_20932,N_18235,N_18878);
xor U20933 (N_20933,N_18799,N_18257);
nand U20934 (N_20934,N_18742,N_19872);
nand U20935 (N_20935,N_18163,N_18916);
nand U20936 (N_20936,N_18898,N_19891);
and U20937 (N_20937,N_18925,N_19683);
nor U20938 (N_20938,N_18007,N_19477);
nand U20939 (N_20939,N_18743,N_19926);
or U20940 (N_20940,N_19042,N_18703);
nand U20941 (N_20941,N_19337,N_18720);
nand U20942 (N_20942,N_18643,N_18340);
or U20943 (N_20943,N_18629,N_18014);
or U20944 (N_20944,N_19482,N_18164);
or U20945 (N_20945,N_19965,N_19600);
nor U20946 (N_20946,N_18078,N_19159);
nor U20947 (N_20947,N_18472,N_19114);
xor U20948 (N_20948,N_19566,N_19398);
nor U20949 (N_20949,N_18637,N_18120);
nor U20950 (N_20950,N_19540,N_18438);
or U20951 (N_20951,N_19089,N_19559);
nor U20952 (N_20952,N_18650,N_19292);
and U20953 (N_20953,N_18580,N_18884);
nand U20954 (N_20954,N_19090,N_18131);
or U20955 (N_20955,N_18070,N_19118);
nor U20956 (N_20956,N_18102,N_19840);
xor U20957 (N_20957,N_18835,N_19340);
xor U20958 (N_20958,N_18621,N_19923);
nand U20959 (N_20959,N_18571,N_19416);
xnor U20960 (N_20960,N_19747,N_19424);
nor U20961 (N_20961,N_18983,N_19806);
or U20962 (N_20962,N_19815,N_19518);
nor U20963 (N_20963,N_19025,N_19596);
nor U20964 (N_20964,N_19206,N_18020);
nand U20965 (N_20965,N_19993,N_18825);
nor U20966 (N_20966,N_19165,N_19147);
and U20967 (N_20967,N_18052,N_19125);
or U20968 (N_20968,N_18686,N_18269);
xor U20969 (N_20969,N_19391,N_18351);
nand U20970 (N_20970,N_18416,N_19802);
nand U20971 (N_20971,N_18886,N_19193);
and U20972 (N_20972,N_18594,N_18043);
nand U20973 (N_20973,N_19630,N_18099);
xnor U20974 (N_20974,N_18821,N_18897);
xor U20975 (N_20975,N_18765,N_19158);
nand U20976 (N_20976,N_18696,N_19487);
xor U20977 (N_20977,N_18028,N_18199);
or U20978 (N_20978,N_18396,N_19951);
nand U20979 (N_20979,N_19764,N_19177);
nor U20980 (N_20980,N_19899,N_19981);
xor U20981 (N_20981,N_19539,N_18376);
nor U20982 (N_20982,N_19245,N_18543);
xor U20983 (N_20983,N_19517,N_19172);
or U20984 (N_20984,N_19842,N_18754);
xnor U20985 (N_20985,N_18306,N_18224);
nor U20986 (N_20986,N_19277,N_19494);
and U20987 (N_20987,N_18233,N_18583);
nand U20988 (N_20988,N_18036,N_18600);
or U20989 (N_20989,N_18947,N_19898);
nand U20990 (N_20990,N_18149,N_18785);
nor U20991 (N_20991,N_18536,N_18943);
or U20992 (N_20992,N_19305,N_18969);
and U20993 (N_20993,N_18284,N_18471);
or U20994 (N_20994,N_19331,N_19351);
nand U20995 (N_20995,N_19712,N_19857);
or U20996 (N_20996,N_19585,N_18463);
and U20997 (N_20997,N_18097,N_19607);
or U20998 (N_20998,N_19363,N_18741);
nand U20999 (N_20999,N_18242,N_18890);
nor U21000 (N_21000,N_18328,N_18439);
nor U21001 (N_21001,N_19481,N_18602);
and U21002 (N_21002,N_19620,N_18556);
nor U21003 (N_21003,N_19733,N_19368);
nor U21004 (N_21004,N_18778,N_18349);
and U21005 (N_21005,N_19948,N_18836);
xor U21006 (N_21006,N_18731,N_18969);
or U21007 (N_21007,N_19398,N_18064);
nand U21008 (N_21008,N_19275,N_18969);
nand U21009 (N_21009,N_19170,N_19871);
and U21010 (N_21010,N_18528,N_18081);
and U21011 (N_21011,N_18755,N_18420);
and U21012 (N_21012,N_18662,N_18054);
nor U21013 (N_21013,N_18635,N_18026);
nor U21014 (N_21014,N_18701,N_18504);
nand U21015 (N_21015,N_18990,N_19038);
and U21016 (N_21016,N_19229,N_18846);
xor U21017 (N_21017,N_19551,N_18513);
nor U21018 (N_21018,N_18500,N_19819);
xnor U21019 (N_21019,N_18003,N_19162);
xnor U21020 (N_21020,N_19829,N_19863);
xor U21021 (N_21021,N_18972,N_18839);
nand U21022 (N_21022,N_18308,N_18020);
and U21023 (N_21023,N_18265,N_18109);
nand U21024 (N_21024,N_18534,N_18595);
xor U21025 (N_21025,N_19130,N_18347);
xor U21026 (N_21026,N_18872,N_19897);
nand U21027 (N_21027,N_19690,N_19629);
or U21028 (N_21028,N_18760,N_19298);
nor U21029 (N_21029,N_19166,N_19557);
xnor U21030 (N_21030,N_18329,N_18806);
and U21031 (N_21031,N_18911,N_19257);
and U21032 (N_21032,N_19923,N_19364);
nor U21033 (N_21033,N_18475,N_19929);
or U21034 (N_21034,N_19986,N_19316);
and U21035 (N_21035,N_19072,N_18502);
nand U21036 (N_21036,N_18318,N_19238);
or U21037 (N_21037,N_19649,N_19597);
and U21038 (N_21038,N_18173,N_18056);
nand U21039 (N_21039,N_18118,N_19495);
nor U21040 (N_21040,N_19545,N_18244);
nor U21041 (N_21041,N_19013,N_18969);
nand U21042 (N_21042,N_18495,N_18285);
and U21043 (N_21043,N_18916,N_18366);
nor U21044 (N_21044,N_18423,N_18364);
nand U21045 (N_21045,N_19761,N_19117);
nor U21046 (N_21046,N_18822,N_19634);
nor U21047 (N_21047,N_18059,N_18355);
or U21048 (N_21048,N_18741,N_19255);
nand U21049 (N_21049,N_19504,N_18655);
or U21050 (N_21050,N_19014,N_18307);
or U21051 (N_21051,N_19518,N_18705);
and U21052 (N_21052,N_19039,N_19445);
xnor U21053 (N_21053,N_18467,N_18330);
nor U21054 (N_21054,N_19675,N_19781);
nor U21055 (N_21055,N_19234,N_19123);
and U21056 (N_21056,N_19471,N_19223);
and U21057 (N_21057,N_18865,N_18489);
nor U21058 (N_21058,N_18949,N_19119);
and U21059 (N_21059,N_19845,N_18925);
nand U21060 (N_21060,N_18298,N_18109);
and U21061 (N_21061,N_18341,N_18825);
nor U21062 (N_21062,N_18889,N_18015);
or U21063 (N_21063,N_18019,N_18259);
xor U21064 (N_21064,N_18492,N_19711);
nor U21065 (N_21065,N_18974,N_18540);
xor U21066 (N_21066,N_19077,N_19434);
and U21067 (N_21067,N_19522,N_18062);
or U21068 (N_21068,N_18937,N_19510);
nor U21069 (N_21069,N_18087,N_18401);
or U21070 (N_21070,N_18850,N_19180);
nor U21071 (N_21071,N_18677,N_18669);
nand U21072 (N_21072,N_18141,N_19899);
nor U21073 (N_21073,N_18739,N_18301);
xnor U21074 (N_21074,N_18189,N_18160);
and U21075 (N_21075,N_19103,N_18905);
xor U21076 (N_21076,N_18675,N_19465);
nor U21077 (N_21077,N_18871,N_19820);
xnor U21078 (N_21078,N_18023,N_18374);
and U21079 (N_21079,N_19295,N_18599);
xor U21080 (N_21080,N_19625,N_19290);
or U21081 (N_21081,N_19857,N_19846);
or U21082 (N_21082,N_19811,N_19454);
nor U21083 (N_21083,N_18806,N_18667);
nor U21084 (N_21084,N_18332,N_18701);
and U21085 (N_21085,N_19515,N_19803);
nand U21086 (N_21086,N_19836,N_19708);
nand U21087 (N_21087,N_18369,N_18912);
and U21088 (N_21088,N_18923,N_19993);
nand U21089 (N_21089,N_19955,N_19389);
or U21090 (N_21090,N_18690,N_18802);
or U21091 (N_21091,N_18662,N_19234);
xnor U21092 (N_21092,N_18975,N_19495);
or U21093 (N_21093,N_18278,N_18090);
or U21094 (N_21094,N_19766,N_19954);
nor U21095 (N_21095,N_19478,N_19842);
nand U21096 (N_21096,N_18496,N_19791);
xnor U21097 (N_21097,N_18813,N_18191);
nor U21098 (N_21098,N_19930,N_19320);
and U21099 (N_21099,N_19092,N_18803);
nand U21100 (N_21100,N_19758,N_18731);
xnor U21101 (N_21101,N_18984,N_19062);
and U21102 (N_21102,N_19464,N_18215);
or U21103 (N_21103,N_18230,N_18703);
nand U21104 (N_21104,N_19280,N_19238);
nand U21105 (N_21105,N_18008,N_18241);
xnor U21106 (N_21106,N_18726,N_19572);
nand U21107 (N_21107,N_19991,N_19560);
and U21108 (N_21108,N_19242,N_18865);
xor U21109 (N_21109,N_18993,N_18975);
nor U21110 (N_21110,N_19228,N_18089);
nand U21111 (N_21111,N_18050,N_19253);
xor U21112 (N_21112,N_18528,N_18228);
and U21113 (N_21113,N_19169,N_19249);
nor U21114 (N_21114,N_18699,N_18379);
xor U21115 (N_21115,N_19714,N_19730);
or U21116 (N_21116,N_19174,N_19821);
nor U21117 (N_21117,N_18507,N_19916);
or U21118 (N_21118,N_18501,N_18241);
and U21119 (N_21119,N_19039,N_19283);
xnor U21120 (N_21120,N_18962,N_18156);
xor U21121 (N_21121,N_18323,N_19113);
and U21122 (N_21122,N_18649,N_18856);
and U21123 (N_21123,N_18749,N_18829);
nor U21124 (N_21124,N_18302,N_18959);
xor U21125 (N_21125,N_19379,N_19512);
xor U21126 (N_21126,N_18351,N_18960);
nor U21127 (N_21127,N_18755,N_18176);
or U21128 (N_21128,N_19080,N_19927);
xnor U21129 (N_21129,N_18887,N_19573);
nor U21130 (N_21130,N_19075,N_19784);
nor U21131 (N_21131,N_18382,N_19758);
xor U21132 (N_21132,N_19275,N_19063);
or U21133 (N_21133,N_18214,N_18876);
and U21134 (N_21134,N_18410,N_19448);
and U21135 (N_21135,N_19049,N_19071);
or U21136 (N_21136,N_18888,N_19109);
nand U21137 (N_21137,N_19073,N_18969);
and U21138 (N_21138,N_19926,N_18665);
and U21139 (N_21139,N_18444,N_19999);
or U21140 (N_21140,N_18693,N_18106);
nor U21141 (N_21141,N_19352,N_18096);
nor U21142 (N_21142,N_19768,N_19145);
and U21143 (N_21143,N_19690,N_18695);
nor U21144 (N_21144,N_19855,N_19975);
nand U21145 (N_21145,N_19234,N_18196);
nand U21146 (N_21146,N_19922,N_19757);
and U21147 (N_21147,N_19789,N_19759);
or U21148 (N_21148,N_19488,N_19963);
nor U21149 (N_21149,N_19770,N_19735);
nand U21150 (N_21150,N_19132,N_19809);
xor U21151 (N_21151,N_19166,N_18937);
nand U21152 (N_21152,N_18220,N_18944);
nand U21153 (N_21153,N_18005,N_19369);
xnor U21154 (N_21154,N_18895,N_19302);
xor U21155 (N_21155,N_19836,N_19612);
and U21156 (N_21156,N_19364,N_18772);
nor U21157 (N_21157,N_19663,N_19728);
nor U21158 (N_21158,N_19930,N_19052);
xor U21159 (N_21159,N_18635,N_18049);
nor U21160 (N_21160,N_19083,N_19615);
nor U21161 (N_21161,N_19578,N_19914);
xor U21162 (N_21162,N_19177,N_19251);
nor U21163 (N_21163,N_18721,N_18265);
xor U21164 (N_21164,N_19766,N_18118);
nor U21165 (N_21165,N_18886,N_19594);
nand U21166 (N_21166,N_18152,N_18467);
xnor U21167 (N_21167,N_19314,N_18386);
or U21168 (N_21168,N_19532,N_19527);
nand U21169 (N_21169,N_18217,N_19424);
or U21170 (N_21170,N_18292,N_19357);
xnor U21171 (N_21171,N_19877,N_18265);
and U21172 (N_21172,N_19708,N_19375);
nor U21173 (N_21173,N_18458,N_19488);
and U21174 (N_21174,N_19437,N_19518);
xor U21175 (N_21175,N_19031,N_18091);
nand U21176 (N_21176,N_18731,N_18070);
or U21177 (N_21177,N_18702,N_19996);
or U21178 (N_21178,N_19013,N_19933);
nor U21179 (N_21179,N_18306,N_19782);
nand U21180 (N_21180,N_19530,N_19575);
xnor U21181 (N_21181,N_19408,N_18422);
or U21182 (N_21182,N_19526,N_18815);
xnor U21183 (N_21183,N_19194,N_18527);
nor U21184 (N_21184,N_18746,N_19787);
nor U21185 (N_21185,N_18880,N_19593);
or U21186 (N_21186,N_19236,N_18329);
or U21187 (N_21187,N_19983,N_19786);
nand U21188 (N_21188,N_19330,N_18006);
xnor U21189 (N_21189,N_18487,N_19680);
xnor U21190 (N_21190,N_18516,N_18971);
nand U21191 (N_21191,N_19969,N_19923);
nor U21192 (N_21192,N_19724,N_18632);
and U21193 (N_21193,N_18967,N_19663);
nor U21194 (N_21194,N_19756,N_19533);
xor U21195 (N_21195,N_18529,N_18950);
nand U21196 (N_21196,N_19545,N_19728);
or U21197 (N_21197,N_19608,N_19738);
xor U21198 (N_21198,N_18204,N_18933);
nor U21199 (N_21199,N_19982,N_19527);
nor U21200 (N_21200,N_18183,N_18638);
or U21201 (N_21201,N_18352,N_18929);
nor U21202 (N_21202,N_18656,N_19175);
nand U21203 (N_21203,N_19164,N_18472);
nand U21204 (N_21204,N_18384,N_19130);
nand U21205 (N_21205,N_19742,N_19459);
nor U21206 (N_21206,N_18007,N_19655);
xor U21207 (N_21207,N_18732,N_19583);
nor U21208 (N_21208,N_18522,N_19015);
nor U21209 (N_21209,N_18211,N_18773);
nand U21210 (N_21210,N_19462,N_19346);
nand U21211 (N_21211,N_18775,N_18105);
and U21212 (N_21212,N_19531,N_18039);
or U21213 (N_21213,N_19858,N_18361);
and U21214 (N_21214,N_18727,N_19704);
and U21215 (N_21215,N_19448,N_19820);
nand U21216 (N_21216,N_18053,N_19395);
and U21217 (N_21217,N_18697,N_18407);
and U21218 (N_21218,N_18072,N_18088);
nand U21219 (N_21219,N_19017,N_19711);
or U21220 (N_21220,N_18248,N_19469);
nand U21221 (N_21221,N_19350,N_18409);
xnor U21222 (N_21222,N_18351,N_18721);
or U21223 (N_21223,N_18080,N_19494);
nor U21224 (N_21224,N_19641,N_18460);
xor U21225 (N_21225,N_19499,N_19064);
nand U21226 (N_21226,N_18689,N_18408);
xnor U21227 (N_21227,N_18723,N_18457);
nor U21228 (N_21228,N_19314,N_18409);
xnor U21229 (N_21229,N_18347,N_18224);
nor U21230 (N_21230,N_18625,N_19526);
and U21231 (N_21231,N_19815,N_18131);
and U21232 (N_21232,N_19738,N_18038);
or U21233 (N_21233,N_18001,N_19328);
nand U21234 (N_21234,N_19690,N_19178);
nand U21235 (N_21235,N_19496,N_19252);
or U21236 (N_21236,N_19261,N_18834);
nor U21237 (N_21237,N_19693,N_19504);
and U21238 (N_21238,N_19702,N_19154);
or U21239 (N_21239,N_18483,N_18158);
nor U21240 (N_21240,N_18810,N_19875);
or U21241 (N_21241,N_19851,N_19955);
and U21242 (N_21242,N_19211,N_18355);
nand U21243 (N_21243,N_19222,N_18570);
and U21244 (N_21244,N_19299,N_19203);
nor U21245 (N_21245,N_18494,N_18603);
and U21246 (N_21246,N_18968,N_19379);
xnor U21247 (N_21247,N_18295,N_19543);
and U21248 (N_21248,N_19518,N_19775);
xor U21249 (N_21249,N_18673,N_18250);
nand U21250 (N_21250,N_19959,N_19926);
or U21251 (N_21251,N_19790,N_18509);
and U21252 (N_21252,N_18019,N_18660);
nor U21253 (N_21253,N_18718,N_18506);
nand U21254 (N_21254,N_18981,N_18157);
nor U21255 (N_21255,N_19272,N_18661);
xor U21256 (N_21256,N_19920,N_18593);
xor U21257 (N_21257,N_18023,N_19042);
nand U21258 (N_21258,N_18653,N_19780);
xor U21259 (N_21259,N_18936,N_19493);
nand U21260 (N_21260,N_18737,N_18381);
xor U21261 (N_21261,N_19438,N_19353);
and U21262 (N_21262,N_18265,N_18395);
xnor U21263 (N_21263,N_18006,N_18280);
and U21264 (N_21264,N_18187,N_18060);
nor U21265 (N_21265,N_19574,N_19163);
nor U21266 (N_21266,N_18197,N_19716);
and U21267 (N_21267,N_18308,N_19808);
and U21268 (N_21268,N_19202,N_18270);
nor U21269 (N_21269,N_18627,N_19220);
nand U21270 (N_21270,N_18628,N_18868);
nor U21271 (N_21271,N_18710,N_19009);
or U21272 (N_21272,N_19583,N_18083);
or U21273 (N_21273,N_19057,N_18261);
nor U21274 (N_21274,N_18710,N_18968);
xnor U21275 (N_21275,N_18428,N_18314);
xor U21276 (N_21276,N_18392,N_19304);
or U21277 (N_21277,N_19323,N_18637);
nand U21278 (N_21278,N_19633,N_19958);
xor U21279 (N_21279,N_19156,N_19987);
nand U21280 (N_21280,N_18273,N_18793);
and U21281 (N_21281,N_19076,N_19586);
xor U21282 (N_21282,N_19685,N_19150);
or U21283 (N_21283,N_19176,N_18117);
nor U21284 (N_21284,N_18611,N_19196);
xor U21285 (N_21285,N_19449,N_18840);
nor U21286 (N_21286,N_18886,N_19382);
nor U21287 (N_21287,N_19385,N_19268);
nor U21288 (N_21288,N_18556,N_19938);
and U21289 (N_21289,N_18633,N_18681);
nand U21290 (N_21290,N_19116,N_18198);
xor U21291 (N_21291,N_19509,N_19457);
nand U21292 (N_21292,N_18158,N_19117);
nor U21293 (N_21293,N_19774,N_18413);
and U21294 (N_21294,N_19873,N_19004);
xor U21295 (N_21295,N_18305,N_18843);
nor U21296 (N_21296,N_18990,N_18699);
nand U21297 (N_21297,N_19249,N_19129);
nor U21298 (N_21298,N_18354,N_18241);
nand U21299 (N_21299,N_19718,N_18253);
or U21300 (N_21300,N_18374,N_19063);
nand U21301 (N_21301,N_19293,N_18798);
xnor U21302 (N_21302,N_18042,N_18515);
or U21303 (N_21303,N_19815,N_18310);
and U21304 (N_21304,N_18608,N_18002);
nand U21305 (N_21305,N_19367,N_18238);
nand U21306 (N_21306,N_19498,N_19337);
and U21307 (N_21307,N_19308,N_18512);
nor U21308 (N_21308,N_18801,N_19674);
or U21309 (N_21309,N_19287,N_19176);
xor U21310 (N_21310,N_18007,N_19858);
nand U21311 (N_21311,N_18571,N_18846);
xnor U21312 (N_21312,N_19893,N_18889);
nand U21313 (N_21313,N_18555,N_18604);
nor U21314 (N_21314,N_18596,N_18572);
nand U21315 (N_21315,N_19162,N_19406);
and U21316 (N_21316,N_18202,N_18933);
nand U21317 (N_21317,N_19132,N_18000);
xor U21318 (N_21318,N_18334,N_18630);
nand U21319 (N_21319,N_18829,N_18093);
and U21320 (N_21320,N_19596,N_19894);
and U21321 (N_21321,N_19347,N_18677);
nand U21322 (N_21322,N_19358,N_19167);
and U21323 (N_21323,N_18780,N_19067);
nor U21324 (N_21324,N_18410,N_19914);
and U21325 (N_21325,N_19042,N_19620);
nand U21326 (N_21326,N_19566,N_19412);
xor U21327 (N_21327,N_18256,N_19917);
nor U21328 (N_21328,N_18092,N_19880);
nor U21329 (N_21329,N_18323,N_18503);
nand U21330 (N_21330,N_19805,N_19251);
or U21331 (N_21331,N_18617,N_19959);
or U21332 (N_21332,N_19507,N_18383);
nand U21333 (N_21333,N_19023,N_19927);
nor U21334 (N_21334,N_19411,N_18773);
nor U21335 (N_21335,N_18748,N_19075);
and U21336 (N_21336,N_18012,N_18334);
or U21337 (N_21337,N_18456,N_19615);
nor U21338 (N_21338,N_19064,N_18685);
xor U21339 (N_21339,N_19795,N_19116);
xnor U21340 (N_21340,N_19506,N_19275);
xnor U21341 (N_21341,N_19315,N_18901);
xnor U21342 (N_21342,N_19991,N_18796);
or U21343 (N_21343,N_18310,N_18501);
or U21344 (N_21344,N_19940,N_19133);
xor U21345 (N_21345,N_18255,N_19646);
or U21346 (N_21346,N_18149,N_19925);
or U21347 (N_21347,N_19796,N_18366);
nor U21348 (N_21348,N_19643,N_19060);
nand U21349 (N_21349,N_18118,N_19442);
xor U21350 (N_21350,N_18528,N_19614);
xnor U21351 (N_21351,N_18978,N_19179);
xnor U21352 (N_21352,N_19403,N_18506);
nand U21353 (N_21353,N_19967,N_19401);
or U21354 (N_21354,N_19810,N_19646);
or U21355 (N_21355,N_19687,N_18763);
xnor U21356 (N_21356,N_18308,N_19291);
xnor U21357 (N_21357,N_18034,N_18024);
nand U21358 (N_21358,N_19889,N_18794);
nand U21359 (N_21359,N_18503,N_18521);
xnor U21360 (N_21360,N_18326,N_19102);
xor U21361 (N_21361,N_19838,N_19604);
and U21362 (N_21362,N_19761,N_18163);
nor U21363 (N_21363,N_19947,N_18891);
nor U21364 (N_21364,N_19469,N_18102);
nand U21365 (N_21365,N_19087,N_18018);
and U21366 (N_21366,N_18847,N_18977);
and U21367 (N_21367,N_18566,N_18312);
nor U21368 (N_21368,N_19722,N_19304);
xor U21369 (N_21369,N_18775,N_19894);
nor U21370 (N_21370,N_19463,N_19816);
and U21371 (N_21371,N_18464,N_19913);
nand U21372 (N_21372,N_19827,N_18403);
and U21373 (N_21373,N_18234,N_18843);
and U21374 (N_21374,N_19525,N_19553);
or U21375 (N_21375,N_19372,N_19883);
xnor U21376 (N_21376,N_18258,N_18077);
and U21377 (N_21377,N_19283,N_19138);
or U21378 (N_21378,N_18602,N_19497);
or U21379 (N_21379,N_19242,N_18116);
nor U21380 (N_21380,N_19879,N_18051);
xor U21381 (N_21381,N_18854,N_19154);
xor U21382 (N_21382,N_18680,N_18850);
xor U21383 (N_21383,N_18137,N_18854);
and U21384 (N_21384,N_19714,N_18702);
nand U21385 (N_21385,N_18949,N_19624);
or U21386 (N_21386,N_19697,N_19840);
and U21387 (N_21387,N_18082,N_19961);
nand U21388 (N_21388,N_19533,N_18995);
or U21389 (N_21389,N_18339,N_19294);
or U21390 (N_21390,N_18695,N_18210);
nand U21391 (N_21391,N_18509,N_18190);
xnor U21392 (N_21392,N_18213,N_18699);
or U21393 (N_21393,N_18260,N_18517);
xor U21394 (N_21394,N_19762,N_19401);
nand U21395 (N_21395,N_18918,N_18161);
xnor U21396 (N_21396,N_19183,N_19884);
and U21397 (N_21397,N_19055,N_19442);
nand U21398 (N_21398,N_18599,N_18908);
nand U21399 (N_21399,N_18452,N_19464);
xnor U21400 (N_21400,N_18613,N_19000);
xor U21401 (N_21401,N_18169,N_18981);
and U21402 (N_21402,N_18344,N_18758);
and U21403 (N_21403,N_19776,N_19925);
xor U21404 (N_21404,N_18603,N_18832);
nand U21405 (N_21405,N_19256,N_18185);
xor U21406 (N_21406,N_19922,N_19148);
and U21407 (N_21407,N_19795,N_18213);
and U21408 (N_21408,N_18050,N_19161);
nor U21409 (N_21409,N_18639,N_18980);
or U21410 (N_21410,N_19741,N_19173);
or U21411 (N_21411,N_19079,N_18260);
xnor U21412 (N_21412,N_18625,N_19174);
xor U21413 (N_21413,N_18520,N_18187);
xor U21414 (N_21414,N_19544,N_19250);
nor U21415 (N_21415,N_18839,N_18668);
and U21416 (N_21416,N_19480,N_19269);
or U21417 (N_21417,N_18761,N_19867);
and U21418 (N_21418,N_18165,N_19092);
nand U21419 (N_21419,N_19065,N_18726);
or U21420 (N_21420,N_18737,N_18137);
nor U21421 (N_21421,N_18509,N_18204);
xnor U21422 (N_21422,N_19985,N_19440);
nor U21423 (N_21423,N_19031,N_19850);
nor U21424 (N_21424,N_19091,N_19987);
xnor U21425 (N_21425,N_19052,N_18013);
and U21426 (N_21426,N_18153,N_19609);
nor U21427 (N_21427,N_18209,N_18234);
xor U21428 (N_21428,N_19496,N_19450);
or U21429 (N_21429,N_18564,N_19862);
nand U21430 (N_21430,N_19086,N_18576);
nor U21431 (N_21431,N_19751,N_19227);
or U21432 (N_21432,N_19832,N_19461);
or U21433 (N_21433,N_18698,N_19001);
or U21434 (N_21434,N_19566,N_19287);
or U21435 (N_21435,N_19872,N_18756);
or U21436 (N_21436,N_18311,N_18546);
and U21437 (N_21437,N_19100,N_18124);
or U21438 (N_21438,N_19532,N_18347);
or U21439 (N_21439,N_19968,N_18080);
or U21440 (N_21440,N_18489,N_18639);
nand U21441 (N_21441,N_18883,N_19097);
nor U21442 (N_21442,N_18926,N_18648);
or U21443 (N_21443,N_18160,N_18784);
or U21444 (N_21444,N_19355,N_18934);
xnor U21445 (N_21445,N_18942,N_18586);
xnor U21446 (N_21446,N_19726,N_19739);
or U21447 (N_21447,N_18890,N_18267);
nand U21448 (N_21448,N_19753,N_19683);
nor U21449 (N_21449,N_18031,N_18819);
xor U21450 (N_21450,N_19077,N_19868);
and U21451 (N_21451,N_19559,N_19129);
nor U21452 (N_21452,N_19243,N_18402);
xor U21453 (N_21453,N_19954,N_19252);
nor U21454 (N_21454,N_19700,N_19194);
xnor U21455 (N_21455,N_19951,N_18287);
nand U21456 (N_21456,N_19381,N_18000);
or U21457 (N_21457,N_18566,N_19282);
or U21458 (N_21458,N_19444,N_19615);
nor U21459 (N_21459,N_18551,N_18983);
nand U21460 (N_21460,N_19369,N_19381);
nor U21461 (N_21461,N_18504,N_18279);
or U21462 (N_21462,N_19444,N_19352);
nor U21463 (N_21463,N_19417,N_18197);
nor U21464 (N_21464,N_19404,N_19864);
xnor U21465 (N_21465,N_18926,N_18303);
and U21466 (N_21466,N_19351,N_19722);
nor U21467 (N_21467,N_18601,N_18841);
nand U21468 (N_21468,N_19873,N_19923);
nor U21469 (N_21469,N_18850,N_18990);
xor U21470 (N_21470,N_18688,N_19461);
or U21471 (N_21471,N_19096,N_18464);
or U21472 (N_21472,N_18534,N_19776);
and U21473 (N_21473,N_18764,N_19890);
xor U21474 (N_21474,N_19450,N_19822);
or U21475 (N_21475,N_19465,N_19251);
xor U21476 (N_21476,N_18508,N_19667);
xor U21477 (N_21477,N_19792,N_18253);
and U21478 (N_21478,N_19604,N_19898);
and U21479 (N_21479,N_18318,N_18986);
nor U21480 (N_21480,N_18388,N_19293);
nand U21481 (N_21481,N_19033,N_18705);
nand U21482 (N_21482,N_19255,N_19229);
nor U21483 (N_21483,N_19213,N_18841);
nand U21484 (N_21484,N_19161,N_19628);
nand U21485 (N_21485,N_19543,N_18938);
nand U21486 (N_21486,N_19425,N_19173);
and U21487 (N_21487,N_19481,N_19979);
or U21488 (N_21488,N_18743,N_18284);
xor U21489 (N_21489,N_19683,N_19419);
xnor U21490 (N_21490,N_19384,N_19800);
xor U21491 (N_21491,N_19536,N_19918);
nor U21492 (N_21492,N_18730,N_19693);
nor U21493 (N_21493,N_19768,N_19662);
nand U21494 (N_21494,N_19662,N_19682);
and U21495 (N_21495,N_19300,N_18827);
or U21496 (N_21496,N_19939,N_18124);
or U21497 (N_21497,N_18511,N_19760);
and U21498 (N_21498,N_18147,N_19866);
and U21499 (N_21499,N_18017,N_19923);
nor U21500 (N_21500,N_18263,N_18578);
xnor U21501 (N_21501,N_19478,N_19347);
nand U21502 (N_21502,N_18220,N_18241);
nor U21503 (N_21503,N_19844,N_18379);
nand U21504 (N_21504,N_18346,N_19457);
or U21505 (N_21505,N_19876,N_19569);
and U21506 (N_21506,N_18036,N_18211);
xnor U21507 (N_21507,N_18960,N_18622);
and U21508 (N_21508,N_18742,N_18210);
nand U21509 (N_21509,N_19504,N_18874);
and U21510 (N_21510,N_18491,N_19197);
nor U21511 (N_21511,N_19036,N_19593);
or U21512 (N_21512,N_19201,N_18267);
xnor U21513 (N_21513,N_19755,N_18867);
xor U21514 (N_21514,N_19156,N_18077);
and U21515 (N_21515,N_19600,N_19968);
and U21516 (N_21516,N_19525,N_19591);
or U21517 (N_21517,N_18399,N_19610);
nor U21518 (N_21518,N_18186,N_18076);
nor U21519 (N_21519,N_19153,N_18430);
nand U21520 (N_21520,N_18054,N_19968);
or U21521 (N_21521,N_19559,N_18014);
nand U21522 (N_21522,N_18401,N_18855);
nand U21523 (N_21523,N_19901,N_18783);
nor U21524 (N_21524,N_19036,N_18532);
xnor U21525 (N_21525,N_19096,N_19163);
or U21526 (N_21526,N_19122,N_18326);
nand U21527 (N_21527,N_18184,N_19667);
nor U21528 (N_21528,N_18784,N_19672);
nor U21529 (N_21529,N_18892,N_19465);
nand U21530 (N_21530,N_19155,N_19593);
and U21531 (N_21531,N_18663,N_19805);
nand U21532 (N_21532,N_19267,N_19746);
or U21533 (N_21533,N_19142,N_19419);
or U21534 (N_21534,N_18068,N_19182);
xor U21535 (N_21535,N_19249,N_19243);
or U21536 (N_21536,N_19764,N_19276);
or U21537 (N_21537,N_18377,N_18184);
or U21538 (N_21538,N_19632,N_18370);
or U21539 (N_21539,N_18420,N_18828);
or U21540 (N_21540,N_18242,N_18423);
or U21541 (N_21541,N_19121,N_19792);
nand U21542 (N_21542,N_19774,N_18230);
xnor U21543 (N_21543,N_19258,N_19257);
or U21544 (N_21544,N_18277,N_18997);
and U21545 (N_21545,N_19295,N_19042);
and U21546 (N_21546,N_18620,N_18640);
and U21547 (N_21547,N_19908,N_19653);
nand U21548 (N_21548,N_18455,N_19583);
nand U21549 (N_21549,N_18395,N_18867);
or U21550 (N_21550,N_18126,N_18128);
nor U21551 (N_21551,N_18164,N_18179);
nor U21552 (N_21552,N_19849,N_19843);
and U21553 (N_21553,N_18919,N_19716);
nor U21554 (N_21554,N_19182,N_18971);
nand U21555 (N_21555,N_18847,N_19518);
xor U21556 (N_21556,N_19622,N_19139);
xnor U21557 (N_21557,N_19727,N_19968);
nand U21558 (N_21558,N_19100,N_18367);
and U21559 (N_21559,N_18740,N_19353);
or U21560 (N_21560,N_19551,N_19797);
or U21561 (N_21561,N_19920,N_19472);
xnor U21562 (N_21562,N_18860,N_19606);
nand U21563 (N_21563,N_19579,N_18428);
or U21564 (N_21564,N_19442,N_19652);
and U21565 (N_21565,N_19791,N_19255);
and U21566 (N_21566,N_18593,N_19035);
or U21567 (N_21567,N_19958,N_19206);
xnor U21568 (N_21568,N_19889,N_19340);
nor U21569 (N_21569,N_19645,N_18959);
xnor U21570 (N_21570,N_19826,N_19450);
nand U21571 (N_21571,N_19842,N_19731);
nand U21572 (N_21572,N_19956,N_19065);
or U21573 (N_21573,N_18450,N_19745);
or U21574 (N_21574,N_19722,N_18194);
and U21575 (N_21575,N_18656,N_18904);
xor U21576 (N_21576,N_18486,N_19329);
nand U21577 (N_21577,N_18279,N_19331);
xnor U21578 (N_21578,N_18880,N_19918);
or U21579 (N_21579,N_19529,N_18126);
nor U21580 (N_21580,N_19158,N_19040);
xnor U21581 (N_21581,N_18067,N_18238);
nand U21582 (N_21582,N_18277,N_19717);
xor U21583 (N_21583,N_19528,N_18951);
nand U21584 (N_21584,N_19684,N_19525);
and U21585 (N_21585,N_19379,N_19672);
nor U21586 (N_21586,N_19836,N_18566);
or U21587 (N_21587,N_18845,N_19477);
nor U21588 (N_21588,N_19189,N_19092);
or U21589 (N_21589,N_18073,N_19186);
and U21590 (N_21590,N_18661,N_19540);
nand U21591 (N_21591,N_18575,N_18391);
and U21592 (N_21592,N_19512,N_18129);
nand U21593 (N_21593,N_19144,N_18435);
and U21594 (N_21594,N_19338,N_19961);
nand U21595 (N_21595,N_18133,N_19869);
nand U21596 (N_21596,N_18562,N_18861);
xor U21597 (N_21597,N_19516,N_19341);
or U21598 (N_21598,N_18682,N_19969);
nand U21599 (N_21599,N_19902,N_18522);
or U21600 (N_21600,N_18059,N_19016);
and U21601 (N_21601,N_19391,N_18239);
xor U21602 (N_21602,N_18527,N_18182);
or U21603 (N_21603,N_18100,N_18487);
and U21604 (N_21604,N_19428,N_18374);
or U21605 (N_21605,N_18494,N_19510);
nor U21606 (N_21606,N_19350,N_19292);
nand U21607 (N_21607,N_18511,N_18418);
and U21608 (N_21608,N_19525,N_19185);
xnor U21609 (N_21609,N_18968,N_19623);
nor U21610 (N_21610,N_19936,N_18561);
xor U21611 (N_21611,N_19627,N_18926);
nand U21612 (N_21612,N_19177,N_19621);
nor U21613 (N_21613,N_19119,N_19009);
or U21614 (N_21614,N_18507,N_19859);
nand U21615 (N_21615,N_18085,N_18914);
xnor U21616 (N_21616,N_18250,N_19380);
xor U21617 (N_21617,N_18596,N_19704);
and U21618 (N_21618,N_19533,N_18788);
and U21619 (N_21619,N_19939,N_19225);
nand U21620 (N_21620,N_18232,N_18717);
nand U21621 (N_21621,N_19008,N_18482);
xor U21622 (N_21622,N_18729,N_18089);
xor U21623 (N_21623,N_18017,N_19196);
and U21624 (N_21624,N_19627,N_19309);
or U21625 (N_21625,N_18365,N_18205);
nor U21626 (N_21626,N_19722,N_18721);
and U21627 (N_21627,N_18569,N_19659);
nor U21628 (N_21628,N_19364,N_19798);
xor U21629 (N_21629,N_18391,N_18858);
xnor U21630 (N_21630,N_18814,N_19861);
or U21631 (N_21631,N_19418,N_19353);
nor U21632 (N_21632,N_19068,N_18240);
nand U21633 (N_21633,N_19832,N_19680);
nand U21634 (N_21634,N_19747,N_19151);
or U21635 (N_21635,N_18914,N_18862);
xor U21636 (N_21636,N_19097,N_18798);
and U21637 (N_21637,N_19209,N_19838);
xnor U21638 (N_21638,N_19899,N_18143);
nand U21639 (N_21639,N_19894,N_18058);
xor U21640 (N_21640,N_19819,N_19193);
xnor U21641 (N_21641,N_18065,N_19475);
nand U21642 (N_21642,N_18457,N_18875);
or U21643 (N_21643,N_18187,N_19866);
xnor U21644 (N_21644,N_18754,N_19446);
and U21645 (N_21645,N_18649,N_19293);
nor U21646 (N_21646,N_19153,N_18680);
nor U21647 (N_21647,N_18064,N_18697);
or U21648 (N_21648,N_18644,N_19180);
nand U21649 (N_21649,N_19684,N_19775);
or U21650 (N_21650,N_18909,N_18764);
nor U21651 (N_21651,N_19898,N_18580);
nor U21652 (N_21652,N_19445,N_19683);
or U21653 (N_21653,N_18352,N_19617);
xor U21654 (N_21654,N_19561,N_19199);
or U21655 (N_21655,N_19686,N_18767);
and U21656 (N_21656,N_18145,N_18861);
or U21657 (N_21657,N_19111,N_18899);
or U21658 (N_21658,N_19945,N_18279);
nand U21659 (N_21659,N_18039,N_18063);
nor U21660 (N_21660,N_19977,N_18542);
and U21661 (N_21661,N_18171,N_19002);
or U21662 (N_21662,N_18939,N_19701);
and U21663 (N_21663,N_18601,N_18739);
nand U21664 (N_21664,N_18315,N_18212);
or U21665 (N_21665,N_18249,N_18031);
nor U21666 (N_21666,N_18223,N_19430);
xnor U21667 (N_21667,N_18275,N_18744);
or U21668 (N_21668,N_18319,N_18270);
or U21669 (N_21669,N_18899,N_18968);
xor U21670 (N_21670,N_18595,N_18548);
xor U21671 (N_21671,N_18190,N_18320);
nand U21672 (N_21672,N_19790,N_18530);
or U21673 (N_21673,N_19642,N_19356);
xor U21674 (N_21674,N_18004,N_18795);
and U21675 (N_21675,N_18294,N_18907);
xnor U21676 (N_21676,N_18662,N_18576);
or U21677 (N_21677,N_18978,N_18735);
nand U21678 (N_21678,N_18011,N_19738);
nor U21679 (N_21679,N_18015,N_18808);
nor U21680 (N_21680,N_19743,N_18757);
nor U21681 (N_21681,N_18899,N_19643);
or U21682 (N_21682,N_19918,N_18293);
xnor U21683 (N_21683,N_18386,N_18958);
or U21684 (N_21684,N_19830,N_18264);
nor U21685 (N_21685,N_18166,N_18236);
nand U21686 (N_21686,N_18421,N_18955);
nand U21687 (N_21687,N_18241,N_19668);
nand U21688 (N_21688,N_18522,N_18221);
and U21689 (N_21689,N_18394,N_18832);
nor U21690 (N_21690,N_19062,N_18649);
nor U21691 (N_21691,N_19489,N_19042);
nor U21692 (N_21692,N_18308,N_18579);
nor U21693 (N_21693,N_18640,N_18548);
or U21694 (N_21694,N_18391,N_18226);
and U21695 (N_21695,N_18054,N_18293);
nand U21696 (N_21696,N_19243,N_19725);
xnor U21697 (N_21697,N_18676,N_18959);
and U21698 (N_21698,N_18121,N_18462);
xor U21699 (N_21699,N_18098,N_19587);
nand U21700 (N_21700,N_18212,N_18907);
and U21701 (N_21701,N_19046,N_19744);
xor U21702 (N_21702,N_19562,N_18506);
xor U21703 (N_21703,N_18780,N_18594);
nor U21704 (N_21704,N_18467,N_19891);
nand U21705 (N_21705,N_18538,N_18591);
nor U21706 (N_21706,N_19932,N_19620);
nor U21707 (N_21707,N_19041,N_18613);
xnor U21708 (N_21708,N_19238,N_19431);
nand U21709 (N_21709,N_18690,N_18326);
xor U21710 (N_21710,N_18631,N_19497);
xnor U21711 (N_21711,N_19789,N_19805);
xnor U21712 (N_21712,N_18485,N_19278);
xnor U21713 (N_21713,N_18874,N_19050);
and U21714 (N_21714,N_18686,N_19429);
or U21715 (N_21715,N_19713,N_18920);
nor U21716 (N_21716,N_19211,N_18583);
and U21717 (N_21717,N_18051,N_18460);
or U21718 (N_21718,N_19981,N_19069);
xor U21719 (N_21719,N_18989,N_18382);
nand U21720 (N_21720,N_18547,N_19032);
and U21721 (N_21721,N_19501,N_19564);
xor U21722 (N_21722,N_19811,N_18588);
and U21723 (N_21723,N_18464,N_18509);
nand U21724 (N_21724,N_18896,N_18300);
or U21725 (N_21725,N_18843,N_18129);
and U21726 (N_21726,N_19913,N_18559);
and U21727 (N_21727,N_19321,N_19747);
xor U21728 (N_21728,N_19424,N_18778);
and U21729 (N_21729,N_19077,N_19198);
nand U21730 (N_21730,N_19171,N_19386);
and U21731 (N_21731,N_18168,N_18609);
nor U21732 (N_21732,N_18288,N_18385);
nor U21733 (N_21733,N_19142,N_19679);
xnor U21734 (N_21734,N_19113,N_19354);
or U21735 (N_21735,N_19752,N_18381);
or U21736 (N_21736,N_18773,N_18741);
nor U21737 (N_21737,N_19332,N_19046);
xor U21738 (N_21738,N_18139,N_18207);
or U21739 (N_21739,N_19301,N_18641);
nand U21740 (N_21740,N_19023,N_18878);
and U21741 (N_21741,N_18441,N_18013);
or U21742 (N_21742,N_19148,N_18601);
or U21743 (N_21743,N_18927,N_18543);
xor U21744 (N_21744,N_18961,N_18600);
xor U21745 (N_21745,N_19003,N_18734);
or U21746 (N_21746,N_19079,N_18699);
nand U21747 (N_21747,N_18050,N_18317);
and U21748 (N_21748,N_19644,N_19232);
or U21749 (N_21749,N_19075,N_19402);
nor U21750 (N_21750,N_19773,N_19753);
and U21751 (N_21751,N_18325,N_18713);
and U21752 (N_21752,N_19958,N_18726);
nor U21753 (N_21753,N_18850,N_19781);
or U21754 (N_21754,N_19597,N_19888);
xnor U21755 (N_21755,N_19675,N_19056);
and U21756 (N_21756,N_18073,N_19904);
or U21757 (N_21757,N_18061,N_18072);
xnor U21758 (N_21758,N_18433,N_18726);
xor U21759 (N_21759,N_18389,N_19100);
xor U21760 (N_21760,N_19508,N_19362);
and U21761 (N_21761,N_18205,N_18169);
and U21762 (N_21762,N_19937,N_19457);
and U21763 (N_21763,N_18952,N_18633);
xnor U21764 (N_21764,N_18377,N_19519);
and U21765 (N_21765,N_19929,N_18616);
xnor U21766 (N_21766,N_19116,N_18561);
xnor U21767 (N_21767,N_19850,N_19308);
and U21768 (N_21768,N_18567,N_18896);
nand U21769 (N_21769,N_19240,N_18131);
nor U21770 (N_21770,N_19043,N_19797);
nand U21771 (N_21771,N_19618,N_18001);
nor U21772 (N_21772,N_18501,N_19152);
xnor U21773 (N_21773,N_18787,N_19469);
and U21774 (N_21774,N_19141,N_18237);
nand U21775 (N_21775,N_18707,N_19734);
or U21776 (N_21776,N_19785,N_19757);
and U21777 (N_21777,N_18895,N_19409);
and U21778 (N_21778,N_18496,N_19131);
or U21779 (N_21779,N_18342,N_19239);
nand U21780 (N_21780,N_18976,N_19105);
nand U21781 (N_21781,N_19301,N_19880);
or U21782 (N_21782,N_19488,N_18251);
and U21783 (N_21783,N_19883,N_19899);
nand U21784 (N_21784,N_18412,N_19689);
xnor U21785 (N_21785,N_18491,N_18953);
nor U21786 (N_21786,N_19515,N_19621);
xnor U21787 (N_21787,N_19233,N_19332);
xor U21788 (N_21788,N_19958,N_19585);
nor U21789 (N_21789,N_18306,N_18741);
or U21790 (N_21790,N_18292,N_18466);
xor U21791 (N_21791,N_18314,N_18424);
nand U21792 (N_21792,N_19969,N_19639);
nor U21793 (N_21793,N_18864,N_19710);
nand U21794 (N_21794,N_18116,N_18831);
nor U21795 (N_21795,N_19307,N_18599);
or U21796 (N_21796,N_19732,N_19893);
and U21797 (N_21797,N_19415,N_18087);
or U21798 (N_21798,N_19534,N_18060);
and U21799 (N_21799,N_19441,N_19422);
xnor U21800 (N_21800,N_18809,N_19360);
xor U21801 (N_21801,N_18140,N_19550);
nor U21802 (N_21802,N_18205,N_18624);
and U21803 (N_21803,N_18928,N_19436);
nand U21804 (N_21804,N_19937,N_19540);
xor U21805 (N_21805,N_19891,N_18461);
xor U21806 (N_21806,N_18295,N_19259);
nor U21807 (N_21807,N_18351,N_19793);
and U21808 (N_21808,N_18594,N_18901);
and U21809 (N_21809,N_18802,N_18209);
nor U21810 (N_21810,N_19158,N_18948);
nand U21811 (N_21811,N_19557,N_18811);
or U21812 (N_21812,N_19388,N_19365);
nand U21813 (N_21813,N_19982,N_19615);
or U21814 (N_21814,N_19169,N_19209);
xor U21815 (N_21815,N_18218,N_19363);
xnor U21816 (N_21816,N_18436,N_18347);
nor U21817 (N_21817,N_18787,N_19994);
xnor U21818 (N_21818,N_18806,N_18709);
and U21819 (N_21819,N_19468,N_18428);
nor U21820 (N_21820,N_19355,N_19580);
and U21821 (N_21821,N_19939,N_18961);
xor U21822 (N_21822,N_18288,N_19426);
or U21823 (N_21823,N_18621,N_19638);
or U21824 (N_21824,N_19217,N_18598);
nor U21825 (N_21825,N_19395,N_18826);
xnor U21826 (N_21826,N_19534,N_19025);
and U21827 (N_21827,N_19636,N_18307);
nand U21828 (N_21828,N_19058,N_18023);
or U21829 (N_21829,N_19840,N_19229);
and U21830 (N_21830,N_18589,N_19763);
xor U21831 (N_21831,N_19427,N_19367);
xnor U21832 (N_21832,N_18192,N_19248);
and U21833 (N_21833,N_18841,N_19212);
or U21834 (N_21834,N_18248,N_19283);
xnor U21835 (N_21835,N_19965,N_19619);
nand U21836 (N_21836,N_18787,N_19500);
xnor U21837 (N_21837,N_19336,N_18810);
nand U21838 (N_21838,N_18066,N_19206);
nand U21839 (N_21839,N_18817,N_19146);
or U21840 (N_21840,N_19029,N_19378);
nand U21841 (N_21841,N_18674,N_18940);
and U21842 (N_21842,N_19196,N_19426);
nor U21843 (N_21843,N_19357,N_18808);
or U21844 (N_21844,N_19860,N_19295);
or U21845 (N_21845,N_18123,N_19867);
nand U21846 (N_21846,N_19961,N_19249);
nor U21847 (N_21847,N_19410,N_18391);
nor U21848 (N_21848,N_18860,N_19050);
and U21849 (N_21849,N_19581,N_19275);
nand U21850 (N_21850,N_18240,N_19916);
or U21851 (N_21851,N_19399,N_18323);
nand U21852 (N_21852,N_18349,N_18996);
or U21853 (N_21853,N_18964,N_18458);
xnor U21854 (N_21854,N_18223,N_18522);
or U21855 (N_21855,N_18933,N_18660);
and U21856 (N_21856,N_18498,N_18117);
nand U21857 (N_21857,N_19175,N_19656);
or U21858 (N_21858,N_18275,N_18781);
and U21859 (N_21859,N_18346,N_18893);
and U21860 (N_21860,N_19260,N_19482);
xor U21861 (N_21861,N_18138,N_19831);
xor U21862 (N_21862,N_18278,N_19526);
nand U21863 (N_21863,N_18960,N_19516);
xnor U21864 (N_21864,N_18618,N_19570);
nand U21865 (N_21865,N_19042,N_19019);
xor U21866 (N_21866,N_19758,N_18990);
xnor U21867 (N_21867,N_19564,N_18403);
nand U21868 (N_21868,N_18842,N_18150);
or U21869 (N_21869,N_19259,N_19396);
or U21870 (N_21870,N_18119,N_18187);
or U21871 (N_21871,N_19170,N_19947);
nor U21872 (N_21872,N_19185,N_19493);
xnor U21873 (N_21873,N_18005,N_18140);
nand U21874 (N_21874,N_18321,N_19163);
nor U21875 (N_21875,N_18759,N_18440);
or U21876 (N_21876,N_18777,N_18825);
xnor U21877 (N_21877,N_18635,N_18085);
nor U21878 (N_21878,N_19064,N_18446);
and U21879 (N_21879,N_18080,N_18430);
nor U21880 (N_21880,N_19556,N_18940);
xor U21881 (N_21881,N_19373,N_19399);
or U21882 (N_21882,N_19451,N_18468);
and U21883 (N_21883,N_18562,N_18324);
nor U21884 (N_21884,N_18916,N_19713);
xor U21885 (N_21885,N_19113,N_19503);
nor U21886 (N_21886,N_18938,N_18961);
nor U21887 (N_21887,N_18560,N_18866);
and U21888 (N_21888,N_18634,N_19662);
nor U21889 (N_21889,N_18685,N_18687);
or U21890 (N_21890,N_19494,N_19896);
nor U21891 (N_21891,N_19400,N_19372);
or U21892 (N_21892,N_18285,N_19179);
or U21893 (N_21893,N_19328,N_19084);
nor U21894 (N_21894,N_19437,N_19422);
and U21895 (N_21895,N_19919,N_18008);
xor U21896 (N_21896,N_18068,N_19435);
or U21897 (N_21897,N_19270,N_18866);
xor U21898 (N_21898,N_19175,N_18933);
nor U21899 (N_21899,N_18596,N_18413);
nor U21900 (N_21900,N_19920,N_19402);
nand U21901 (N_21901,N_18345,N_19376);
and U21902 (N_21902,N_18262,N_19500);
and U21903 (N_21903,N_19549,N_19477);
or U21904 (N_21904,N_18589,N_18579);
nand U21905 (N_21905,N_18434,N_18160);
and U21906 (N_21906,N_19961,N_18505);
nand U21907 (N_21907,N_19786,N_19705);
nor U21908 (N_21908,N_18835,N_18913);
and U21909 (N_21909,N_18675,N_18346);
xnor U21910 (N_21910,N_19203,N_19611);
and U21911 (N_21911,N_19571,N_18466);
xnor U21912 (N_21912,N_18806,N_19203);
nand U21913 (N_21913,N_19938,N_18380);
and U21914 (N_21914,N_18074,N_18963);
or U21915 (N_21915,N_18244,N_19100);
and U21916 (N_21916,N_19018,N_18937);
xnor U21917 (N_21917,N_19034,N_19373);
xor U21918 (N_21918,N_18174,N_18856);
nand U21919 (N_21919,N_19186,N_19334);
nand U21920 (N_21920,N_18096,N_18268);
or U21921 (N_21921,N_19621,N_18616);
and U21922 (N_21922,N_19474,N_18067);
nor U21923 (N_21923,N_18747,N_18638);
xor U21924 (N_21924,N_19828,N_18681);
xor U21925 (N_21925,N_19708,N_19243);
nor U21926 (N_21926,N_18948,N_18690);
nor U21927 (N_21927,N_19417,N_19590);
nor U21928 (N_21928,N_19260,N_19616);
nand U21929 (N_21929,N_18193,N_18797);
or U21930 (N_21930,N_19868,N_19758);
and U21931 (N_21931,N_19330,N_18923);
and U21932 (N_21932,N_19651,N_19428);
nand U21933 (N_21933,N_18035,N_18117);
nand U21934 (N_21934,N_19113,N_19248);
nor U21935 (N_21935,N_18804,N_18783);
and U21936 (N_21936,N_19572,N_18912);
nor U21937 (N_21937,N_19876,N_18823);
or U21938 (N_21938,N_18957,N_18832);
nor U21939 (N_21939,N_19468,N_19821);
xor U21940 (N_21940,N_18537,N_18151);
or U21941 (N_21941,N_18465,N_19221);
xor U21942 (N_21942,N_18741,N_19687);
and U21943 (N_21943,N_18106,N_18636);
or U21944 (N_21944,N_19658,N_19707);
nor U21945 (N_21945,N_18129,N_19397);
and U21946 (N_21946,N_19531,N_18542);
nor U21947 (N_21947,N_19311,N_19832);
nor U21948 (N_21948,N_18341,N_19584);
xor U21949 (N_21949,N_18506,N_19544);
nand U21950 (N_21950,N_19939,N_18429);
or U21951 (N_21951,N_19019,N_18400);
nor U21952 (N_21952,N_18325,N_18940);
xnor U21953 (N_21953,N_18819,N_19554);
and U21954 (N_21954,N_19077,N_19632);
and U21955 (N_21955,N_19092,N_19340);
and U21956 (N_21956,N_18100,N_19342);
and U21957 (N_21957,N_18340,N_19084);
xor U21958 (N_21958,N_18668,N_19722);
xor U21959 (N_21959,N_19946,N_18854);
or U21960 (N_21960,N_18429,N_18512);
nand U21961 (N_21961,N_18098,N_18922);
nor U21962 (N_21962,N_18815,N_19693);
nand U21963 (N_21963,N_18617,N_19198);
nor U21964 (N_21964,N_18370,N_18219);
and U21965 (N_21965,N_19568,N_19609);
nor U21966 (N_21966,N_19498,N_18680);
or U21967 (N_21967,N_19274,N_18958);
and U21968 (N_21968,N_19826,N_18586);
or U21969 (N_21969,N_18480,N_18652);
and U21970 (N_21970,N_18969,N_18787);
xor U21971 (N_21971,N_18665,N_19482);
xnor U21972 (N_21972,N_19440,N_18428);
xor U21973 (N_21973,N_18822,N_18229);
xnor U21974 (N_21974,N_18774,N_19624);
and U21975 (N_21975,N_18172,N_18454);
and U21976 (N_21976,N_19233,N_19564);
nand U21977 (N_21977,N_19956,N_19153);
and U21978 (N_21978,N_18317,N_18037);
nand U21979 (N_21979,N_19638,N_18596);
nand U21980 (N_21980,N_19257,N_18405);
nand U21981 (N_21981,N_18221,N_18450);
nand U21982 (N_21982,N_19367,N_18424);
xnor U21983 (N_21983,N_18161,N_18959);
and U21984 (N_21984,N_18450,N_18045);
xor U21985 (N_21985,N_18242,N_18624);
xor U21986 (N_21986,N_19340,N_18701);
and U21987 (N_21987,N_18703,N_19835);
xnor U21988 (N_21988,N_19095,N_19065);
nand U21989 (N_21989,N_18320,N_19272);
or U21990 (N_21990,N_18009,N_19419);
nor U21991 (N_21991,N_19288,N_18424);
nand U21992 (N_21992,N_18458,N_18091);
nor U21993 (N_21993,N_19074,N_19825);
xnor U21994 (N_21994,N_19531,N_18189);
xor U21995 (N_21995,N_18941,N_18147);
xnor U21996 (N_21996,N_19540,N_18370);
or U21997 (N_21997,N_19540,N_19404);
nand U21998 (N_21998,N_18741,N_18738);
nor U21999 (N_21999,N_19977,N_19326);
xnor U22000 (N_22000,N_20159,N_20839);
and U22001 (N_22001,N_21534,N_21618);
and U22002 (N_22002,N_20547,N_20079);
or U22003 (N_22003,N_21375,N_20946);
nand U22004 (N_22004,N_20738,N_21461);
nor U22005 (N_22005,N_20324,N_21174);
or U22006 (N_22006,N_21969,N_20377);
nor U22007 (N_22007,N_20838,N_21412);
xnor U22008 (N_22008,N_20729,N_21398);
nor U22009 (N_22009,N_21465,N_21466);
xnor U22010 (N_22010,N_21245,N_20970);
xor U22011 (N_22011,N_20577,N_21148);
or U22012 (N_22012,N_21057,N_21274);
nand U22013 (N_22013,N_20129,N_20570);
nand U22014 (N_22014,N_20501,N_20048);
nor U22015 (N_22015,N_20020,N_21912);
or U22016 (N_22016,N_21389,N_20600);
or U22017 (N_22017,N_20447,N_21202);
xor U22018 (N_22018,N_21304,N_20574);
nor U22019 (N_22019,N_21681,N_20031);
or U22020 (N_22020,N_21471,N_20780);
or U22021 (N_22021,N_20393,N_20268);
xor U22022 (N_22022,N_20597,N_20016);
xnor U22023 (N_22023,N_21998,N_21509);
xor U22024 (N_22024,N_21716,N_20476);
or U22025 (N_22025,N_21635,N_20845);
or U22026 (N_22026,N_21826,N_20110);
and U22027 (N_22027,N_20088,N_20170);
xor U22028 (N_22028,N_20892,N_21033);
and U22029 (N_22029,N_20888,N_20550);
or U22030 (N_22030,N_20921,N_20056);
and U22031 (N_22031,N_20227,N_21450);
nand U22032 (N_22032,N_21090,N_21076);
and U22033 (N_22033,N_21356,N_20701);
and U22034 (N_22034,N_21967,N_21833);
nor U22035 (N_22035,N_21871,N_20144);
xnor U22036 (N_22036,N_21229,N_21013);
nor U22037 (N_22037,N_21919,N_21032);
nand U22038 (N_22038,N_21784,N_20622);
and U22039 (N_22039,N_21844,N_21539);
or U22040 (N_22040,N_20416,N_21141);
and U22041 (N_22041,N_20638,N_21879);
nand U22042 (N_22042,N_20741,N_20230);
xor U22043 (N_22043,N_20601,N_20507);
xnor U22044 (N_22044,N_21880,N_20090);
xnor U22045 (N_22045,N_20074,N_21649);
or U22046 (N_22046,N_21042,N_21055);
and U22047 (N_22047,N_20042,N_21593);
and U22048 (N_22048,N_21532,N_20906);
xor U22049 (N_22049,N_21894,N_21080);
nand U22050 (N_22050,N_21835,N_20357);
xnor U22051 (N_22051,N_20339,N_21469);
and U22052 (N_22052,N_21902,N_20855);
nand U22053 (N_22053,N_20382,N_20512);
and U22054 (N_22054,N_20288,N_20976);
or U22055 (N_22055,N_20718,N_21194);
and U22056 (N_22056,N_20967,N_20938);
or U22057 (N_22057,N_21993,N_20896);
nor U22058 (N_22058,N_20665,N_21648);
or U22059 (N_22059,N_21801,N_20030);
and U22060 (N_22060,N_21711,N_20289);
nand U22061 (N_22061,N_21438,N_20717);
nor U22062 (N_22062,N_21143,N_21665);
or U22063 (N_22063,N_21760,N_21212);
nand U22064 (N_22064,N_21232,N_20740);
nor U22065 (N_22065,N_20290,N_21970);
nor U22066 (N_22066,N_20522,N_20829);
nor U22067 (N_22067,N_20452,N_20531);
and U22068 (N_22068,N_21875,N_21252);
xnor U22069 (N_22069,N_21577,N_21052);
and U22070 (N_22070,N_20878,N_20397);
nor U22071 (N_22071,N_20980,N_20140);
or U22072 (N_22072,N_21776,N_20508);
or U22073 (N_22073,N_20702,N_20524);
nand U22074 (N_22074,N_20361,N_20007);
or U22075 (N_22075,N_20637,N_20295);
and U22076 (N_22076,N_21581,N_21300);
and U22077 (N_22077,N_21311,N_20802);
nand U22078 (N_22078,N_20883,N_20891);
xnor U22079 (N_22079,N_20242,N_21876);
nand U22080 (N_22080,N_20816,N_21280);
nor U22081 (N_22081,N_20109,N_20605);
and U22082 (N_22082,N_21161,N_20572);
nand U22083 (N_22083,N_20441,N_20486);
nor U22084 (N_22084,N_21035,N_21462);
and U22085 (N_22085,N_20199,N_21775);
xnor U22086 (N_22086,N_21866,N_20279);
xnor U22087 (N_22087,N_21359,N_21120);
and U22088 (N_22088,N_20443,N_21060);
nor U22089 (N_22089,N_20058,N_21352);
or U22090 (N_22090,N_20472,N_20205);
or U22091 (N_22091,N_21854,N_20478);
and U22092 (N_22092,N_20984,N_20898);
and U22093 (N_22093,N_21504,N_21544);
nor U22094 (N_22094,N_21510,N_21059);
or U22095 (N_22095,N_20352,N_21246);
nor U22096 (N_22096,N_20540,N_21432);
and U22097 (N_22097,N_20419,N_20315);
nand U22098 (N_22098,N_21550,N_20425);
or U22099 (N_22099,N_21898,N_20530);
or U22100 (N_22100,N_20787,N_21038);
and U22101 (N_22101,N_21627,N_21315);
or U22102 (N_22102,N_20463,N_20911);
and U22103 (N_22103,N_21123,N_20889);
xor U22104 (N_22104,N_20256,N_20971);
and U22105 (N_22105,N_21044,N_21028);
or U22106 (N_22106,N_20364,N_21870);
nand U22107 (N_22107,N_21022,N_20111);
nand U22108 (N_22108,N_21670,N_21363);
nor U22109 (N_22109,N_21354,N_20498);
xor U22110 (N_22110,N_20595,N_20826);
or U22111 (N_22111,N_21702,N_20102);
or U22112 (N_22112,N_20859,N_21977);
or U22113 (N_22113,N_20591,N_20190);
or U22114 (N_22114,N_21507,N_21522);
xor U22115 (N_22115,N_20615,N_20618);
nor U22116 (N_22116,N_20006,N_21523);
and U22117 (N_22117,N_20026,N_21454);
nand U22118 (N_22118,N_20342,N_21756);
or U22119 (N_22119,N_20143,N_21125);
or U22120 (N_22120,N_21139,N_20621);
or U22121 (N_22121,N_21477,N_21690);
and U22122 (N_22122,N_21424,N_21473);
nor U22123 (N_22123,N_21547,N_20926);
nor U22124 (N_22124,N_20582,N_21804);
and U22125 (N_22125,N_20499,N_21700);
and U22126 (N_22126,N_20163,N_21335);
xnor U22127 (N_22127,N_21272,N_21641);
nor U22128 (N_22128,N_21346,N_21049);
nor U22129 (N_22129,N_20487,N_21892);
or U22130 (N_22130,N_21831,N_21347);
and U22131 (N_22131,N_20010,N_20843);
nand U22132 (N_22132,N_21843,N_20861);
nand U22133 (N_22133,N_21572,N_21338);
nor U22134 (N_22134,N_21034,N_21147);
and U22135 (N_22135,N_20220,N_20022);
and U22136 (N_22136,N_20602,N_20917);
xnor U22137 (N_22137,N_21729,N_20726);
xnor U22138 (N_22138,N_21185,N_20100);
xnor U22139 (N_22139,N_21806,N_20756);
and U22140 (N_22140,N_21789,N_20142);
and U22141 (N_22141,N_20505,N_21312);
or U22142 (N_22142,N_21910,N_20520);
nand U22143 (N_22143,N_21231,N_21759);
and U22144 (N_22144,N_20837,N_20690);
and U22145 (N_22145,N_21289,N_21554);
or U22146 (N_22146,N_21786,N_20616);
nor U22147 (N_22147,N_21286,N_21269);
xor U22148 (N_22148,N_21561,N_21193);
nor U22149 (N_22149,N_20387,N_20404);
nor U22150 (N_22150,N_21737,N_20977);
xor U22151 (N_22151,N_20529,N_21241);
xor U22152 (N_22152,N_20200,N_20626);
xnor U22153 (N_22153,N_21939,N_21991);
and U22154 (N_22154,N_21244,N_21658);
or U22155 (N_22155,N_20224,N_20293);
or U22156 (N_22156,N_20745,N_20444);
or U22157 (N_22157,N_20092,N_21719);
nand U22158 (N_22158,N_21883,N_20354);
or U22159 (N_22159,N_20960,N_20502);
and U22160 (N_22160,N_21137,N_21221);
xnor U22161 (N_22161,N_21739,N_20484);
or U22162 (N_22162,N_21294,N_21376);
xor U22163 (N_22163,N_21230,N_20536);
nand U22164 (N_22164,N_21934,N_21004);
xor U22165 (N_22165,N_20932,N_20687);
or U22166 (N_22166,N_20933,N_21330);
xor U22167 (N_22167,N_20796,N_20306);
and U22168 (N_22168,N_20269,N_21911);
and U22169 (N_22169,N_21131,N_20617);
xor U22170 (N_22170,N_21515,N_21606);
and U22171 (N_22171,N_20019,N_21390);
nand U22172 (N_22172,N_20045,N_21021);
nor U22173 (N_22173,N_20321,N_21345);
and U22174 (N_22174,N_21811,N_20211);
nand U22175 (N_22175,N_20203,N_20824);
and U22176 (N_22176,N_21709,N_21565);
and U22177 (N_22177,N_20251,N_21855);
nand U22178 (N_22178,N_20981,N_21130);
xor U22179 (N_22179,N_20335,N_20396);
or U22180 (N_22180,N_21698,N_21985);
nand U22181 (N_22181,N_20809,N_20271);
nand U22182 (N_22182,N_21132,N_20852);
nor U22183 (N_22183,N_20332,N_21490);
and U22184 (N_22184,N_20465,N_20997);
or U22185 (N_22185,N_20681,N_20526);
and U22186 (N_22186,N_21845,N_21113);
nor U22187 (N_22187,N_21749,N_20510);
and U22188 (N_22188,N_20316,N_20871);
and U22189 (N_22189,N_21521,N_20669);
or U22190 (N_22190,N_21664,N_21195);
xnor U22191 (N_22191,N_20453,N_20732);
or U22192 (N_22192,N_20018,N_21418);
or U22193 (N_22193,N_20151,N_20746);
and U22194 (N_22194,N_21543,N_20770);
nor U22195 (N_22195,N_21429,N_21236);
nor U22196 (N_22196,N_21582,N_21434);
or U22197 (N_22197,N_20059,N_20327);
xnor U22198 (N_22198,N_21552,N_20811);
nand U22199 (N_22199,N_20978,N_21571);
and U22200 (N_22200,N_20947,N_21407);
nor U22201 (N_22201,N_21520,N_20781);
nand U22202 (N_22202,N_21744,N_21814);
or U22203 (N_22203,N_21129,N_21180);
nor U22204 (N_22204,N_20473,N_21400);
nor U22205 (N_22205,N_21247,N_20683);
xnor U22206 (N_22206,N_21107,N_21783);
nand U22207 (N_22207,N_20937,N_21896);
nor U22208 (N_22208,N_21667,N_21134);
or U22209 (N_22209,N_20614,N_21943);
nand U22210 (N_22210,N_21440,N_20189);
nand U22211 (N_22211,N_20180,N_21070);
or U22212 (N_22212,N_21301,N_20710);
and U22213 (N_22213,N_21358,N_21607);
xor U22214 (N_22214,N_20334,N_21474);
nor U22215 (N_22215,N_21036,N_20231);
nor U22216 (N_22216,N_21858,N_20401);
nand U22217 (N_22217,N_20875,N_21106);
nor U22218 (N_22218,N_21039,N_21248);
nand U22219 (N_22219,N_20500,N_20901);
nor U22220 (N_22220,N_20558,N_21094);
and U22221 (N_22221,N_21742,N_20655);
nor U22222 (N_22222,N_20094,N_21923);
xor U22223 (N_22223,N_21045,N_21672);
nand U22224 (N_22224,N_20281,N_20175);
nand U22225 (N_22225,N_21388,N_21478);
nand U22226 (N_22226,N_20751,N_21209);
nor U22227 (N_22227,N_21256,N_21483);
or U22228 (N_22228,N_20286,N_21242);
or U22229 (N_22229,N_20709,N_20069);
or U22230 (N_22230,N_20713,N_20928);
nor U22231 (N_22231,N_21747,N_20674);
nor U22232 (N_22232,N_20158,N_21529);
xnor U22233 (N_22233,N_20696,N_21973);
nor U22234 (N_22234,N_20183,N_20569);
xor U22235 (N_22235,N_21463,N_21839);
and U22236 (N_22236,N_20988,N_20262);
xnor U22237 (N_22237,N_20439,N_20095);
or U22238 (N_22238,N_20238,N_21965);
xnor U22239 (N_22239,N_21992,N_21030);
or U22240 (N_22240,N_20044,N_20769);
nand U22241 (N_22241,N_20370,N_21237);
and U22242 (N_22242,N_20273,N_21159);
nor U22243 (N_22243,N_20025,N_20842);
nand U22244 (N_22244,N_20579,N_21476);
xnor U22245 (N_22245,N_20821,N_21733);
xor U22246 (N_22246,N_20834,N_20098);
or U22247 (N_22247,N_21083,N_20897);
xnor U22248 (N_22248,N_20803,N_20840);
nand U22249 (N_22249,N_21266,N_20194);
xnor U22250 (N_22250,N_20649,N_20849);
nand U22251 (N_22251,N_20137,N_20765);
or U22252 (N_22252,N_21095,N_20503);
and U22253 (N_22253,N_21740,N_20879);
xnor U22254 (N_22254,N_21608,N_21546);
nand U22255 (N_22255,N_21753,N_20394);
and U22256 (N_22256,N_20552,N_20373);
nor U22257 (N_22257,N_20658,N_21995);
and U22258 (N_22258,N_20749,N_20676);
or U22259 (N_22259,N_20688,N_20504);
nand U22260 (N_22260,N_21428,N_21941);
nor U22261 (N_22261,N_21367,N_20122);
nand U22262 (N_22262,N_21555,N_21084);
and U22263 (N_22263,N_21479,N_21575);
nor U22264 (N_22264,N_20551,N_20403);
nor U22265 (N_22265,N_21284,N_21817);
nor U22266 (N_22266,N_21932,N_20703);
nor U22267 (N_22267,N_20454,N_20790);
nand U22268 (N_22268,N_21423,N_20073);
nand U22269 (N_22269,N_20483,N_21558);
nor U22270 (N_22270,N_21344,N_20351);
and U22271 (N_22271,N_21173,N_20877);
xnor U22272 (N_22272,N_21903,N_20544);
nand U22273 (N_22273,N_20784,N_21708);
and U22274 (N_22274,N_21926,N_21278);
nor U22275 (N_22275,N_20645,N_21500);
nand U22276 (N_22276,N_21172,N_20167);
nand U22277 (N_22277,N_21947,N_20436);
nand U22278 (N_22278,N_21974,N_21836);
nand U22279 (N_22279,N_21798,N_21767);
xor U22280 (N_22280,N_20782,N_21273);
xnor U22281 (N_22281,N_20931,N_21018);
nor U22282 (N_22282,N_20263,N_21309);
nor U22283 (N_22283,N_21891,N_21647);
nor U22284 (N_22284,N_21368,N_21701);
nand U22285 (N_22285,N_20722,N_21907);
xnor U22286 (N_22286,N_20598,N_20154);
nand U22287 (N_22287,N_20868,N_21815);
nand U22288 (N_22288,N_21818,N_21730);
xor U22289 (N_22289,N_20402,N_21766);
or U22290 (N_22290,N_20319,N_20525);
and U22291 (N_22291,N_20573,N_21852);
or U22292 (N_22292,N_20982,N_20628);
nand U22293 (N_22293,N_20236,N_20232);
and U22294 (N_22294,N_20280,N_20580);
nand U22295 (N_22295,N_21240,N_21557);
or U22296 (N_22296,N_20185,N_21986);
and U22297 (N_22297,N_21849,N_21255);
and U22298 (N_22298,N_21206,N_21218);
xnor U22299 (N_22299,N_20858,N_21570);
nor U22300 (N_22300,N_20479,N_20715);
and U22301 (N_22301,N_21366,N_21638);
or U22302 (N_22302,N_20862,N_21408);
nor U22303 (N_22303,N_21937,N_20378);
xor U22304 (N_22304,N_20623,N_21614);
nand U22305 (N_22305,N_20777,N_20139);
nor U22306 (N_22306,N_21645,N_21679);
xor U22307 (N_22307,N_21281,N_20533);
nand U22308 (N_22308,N_21293,N_21303);
nand U22309 (N_22309,N_20046,N_21207);
and U22310 (N_22310,N_21054,N_20063);
and U22311 (N_22311,N_20460,N_21204);
or U22312 (N_22312,N_21097,N_20193);
and U22313 (N_22313,N_21167,N_21292);
nand U22314 (N_22314,N_21014,N_21600);
or U22315 (N_22315,N_20349,N_20346);
and U22316 (N_22316,N_21596,N_21601);
xnor U22317 (N_22317,N_21000,N_20944);
and U22318 (N_22318,N_21168,N_20797);
and U22319 (N_22319,N_21545,N_20663);
or U22320 (N_22320,N_21769,N_20241);
and U22321 (N_22321,N_20664,N_21928);
or U22322 (N_22322,N_20055,N_20548);
and U22323 (N_22323,N_21685,N_21604);
nor U22324 (N_22324,N_20390,N_21074);
nor U22325 (N_22325,N_21401,N_21020);
nor U22326 (N_22326,N_21897,N_20651);
or U22327 (N_22327,N_21830,N_20107);
nand U22328 (N_22328,N_20958,N_21961);
xor U22329 (N_22329,N_21707,N_20927);
nand U22330 (N_22330,N_20358,N_20596);
nand U22331 (N_22331,N_21517,N_21265);
nand U22332 (N_22332,N_20792,N_20174);
nand U22333 (N_22333,N_20913,N_21427);
or U22334 (N_22334,N_21287,N_20712);
or U22335 (N_22335,N_20819,N_21157);
or U22336 (N_22336,N_21290,N_21153);
or U22337 (N_22337,N_20311,N_21958);
xnor U22338 (N_22338,N_21693,N_21512);
xor U22339 (N_22339,N_21873,N_21436);
or U22340 (N_22340,N_21187,N_20461);
and U22341 (N_22341,N_21689,N_21069);
nand U22342 (N_22342,N_20607,N_21164);
or U22343 (N_22343,N_20034,N_21151);
nor U22344 (N_22344,N_20497,N_21444);
nor U22345 (N_22345,N_20283,N_20996);
and U22346 (N_22346,N_21372,N_20294);
and U22347 (N_22347,N_20310,N_20767);
xnor U22348 (N_22348,N_21043,N_20458);
and U22349 (N_22349,N_21816,N_20642);
nor U22350 (N_22350,N_20320,N_21752);
and U22351 (N_22351,N_21082,N_20631);
nor U22352 (N_22352,N_21703,N_20060);
and U22353 (N_22353,N_20491,N_20630);
and U22354 (N_22354,N_21111,N_21340);
xor U22355 (N_22355,N_21807,N_20089);
and U22356 (N_22356,N_20993,N_20455);
nand U22357 (N_22357,N_20347,N_20736);
or U22358 (N_22358,N_21940,N_20920);
nand U22359 (N_22359,N_21735,N_20537);
nor U22360 (N_22360,N_20994,N_21223);
and U22361 (N_22361,N_20559,N_20150);
nor U22362 (N_22362,N_21396,N_20429);
xor U22363 (N_22363,N_21334,N_21813);
xnor U22364 (N_22364,N_20495,N_21254);
or U22365 (N_22365,N_21562,N_20894);
nand U22366 (N_22366,N_21109,N_20935);
xor U22367 (N_22367,N_20388,N_21373);
nor U22368 (N_22368,N_21015,N_20748);
or U22369 (N_22369,N_20005,N_21659);
or U22370 (N_22370,N_20851,N_21380);
or U22371 (N_22371,N_21331,N_20481);
nand U22372 (N_22372,N_20274,N_20808);
nor U22373 (N_22373,N_21738,N_21307);
nor U22374 (N_22374,N_21761,N_20583);
or U22375 (N_22375,N_21683,N_21694);
or U22376 (N_22376,N_21640,N_20235);
nor U22377 (N_22377,N_21633,N_20934);
and U22378 (N_22378,N_21857,N_21598);
nand U22379 (N_22379,N_21644,N_21416);
or U22380 (N_22380,N_21224,N_20385);
xor U22381 (N_22381,N_20684,N_21771);
nor U22382 (N_22382,N_21096,N_21364);
nor U22383 (N_22383,N_21916,N_20517);
and U22384 (N_22384,N_20433,N_20575);
or U22385 (N_22385,N_20365,N_21175);
nand U22386 (N_22386,N_20023,N_21170);
and U22387 (N_22387,N_21104,N_20774);
xnor U22388 (N_22388,N_21895,N_20966);
xor U22389 (N_22389,N_20881,N_21397);
nor U22390 (N_22390,N_21486,N_20204);
nand U22391 (N_22391,N_21990,N_20490);
xor U22392 (N_22392,N_20693,N_21182);
nand U22393 (N_22393,N_20082,N_20084);
nand U22394 (N_22394,N_20253,N_21877);
nand U22395 (N_22395,N_20719,N_20817);
or U22396 (N_22396,N_20188,N_21727);
or U22397 (N_22397,N_20141,N_20181);
nor U22398 (N_22398,N_20820,N_21442);
and U22399 (N_22399,N_20314,N_20954);
and U22400 (N_22400,N_21800,N_20964);
xnor U22401 (N_22401,N_21395,N_20219);
nor U22402 (N_22402,N_20431,N_20720);
and U22403 (N_22403,N_20379,N_20240);
nor U22404 (N_22404,N_21447,N_20768);
and U22405 (N_22405,N_21865,N_21646);
or U22406 (N_22406,N_20187,N_20343);
xnor U22407 (N_22407,N_20223,N_21446);
and U22408 (N_22408,N_20835,N_20773);
and U22409 (N_22409,N_21503,N_21092);
nor U22410 (N_22410,N_20576,N_21488);
nand U22411 (N_22411,N_20196,N_21636);
nand U22412 (N_22412,N_20940,N_20610);
and U22413 (N_22413,N_20474,N_20534);
and U22414 (N_22414,N_21580,N_21122);
xnor U22415 (N_22415,N_20519,N_21119);
xor U22416 (N_22416,N_20899,N_20359);
nor U22417 (N_22417,N_20671,N_21467);
or U22418 (N_22418,N_20822,N_21656);
and U22419 (N_22419,N_20606,N_20698);
nand U22420 (N_22420,N_20105,N_20113);
and U22421 (N_22421,N_20305,N_20376);
or U22422 (N_22422,N_20832,N_20677);
or U22423 (N_22423,N_21812,N_20162);
nor U22424 (N_22424,N_20567,N_20884);
and U22425 (N_22425,N_21056,N_21513);
xnor U22426 (N_22426,N_20653,N_21868);
xor U22427 (N_22427,N_20764,N_21590);
nand U22428 (N_22428,N_20226,N_20087);
nand U22429 (N_22429,N_20426,N_21688);
nand U22430 (N_22430,N_21920,N_21313);
xor U22431 (N_22431,N_21603,N_21979);
xnor U22432 (N_22432,N_21699,N_21305);
nor U22433 (N_22433,N_20662,N_21774);
xor U22434 (N_22434,N_20369,N_21653);
and U22435 (N_22435,N_20915,N_21142);
nand U22436 (N_22436,N_20644,N_21861);
and U22437 (N_22437,N_20147,N_21795);
xor U22438 (N_22438,N_20846,N_20464);
nor U22439 (N_22439,N_21799,N_20728);
nor U22440 (N_22440,N_21960,N_20000);
or U22441 (N_22441,N_20656,N_21628);
nand U22442 (N_22442,N_20560,N_21382);
xnor U22443 (N_22443,N_20149,N_20914);
or U22444 (N_22444,N_20130,N_20546);
nand U22445 (N_22445,N_20998,N_20075);
and U22446 (N_22446,N_20116,N_21867);
xor U22447 (N_22447,N_21549,N_21900);
nor U22448 (N_22448,N_21150,N_21158);
and U22449 (N_22449,N_21211,N_21631);
or U22450 (N_22450,N_21415,N_20912);
nor U22451 (N_22451,N_20260,N_21654);
and U22452 (N_22452,N_21073,N_20833);
nor U22453 (N_22453,N_20890,N_21351);
and U22454 (N_22454,N_20318,N_20568);
or U22455 (N_22455,N_21062,N_21944);
and U22456 (N_22456,N_21957,N_20864);
nor U22457 (N_22457,N_21921,N_21984);
xnor U22458 (N_22458,N_21959,N_20024);
or U22459 (N_22459,N_21085,N_21797);
nor U22460 (N_22460,N_21061,N_21077);
nor U22461 (N_22461,N_21361,N_20789);
and U22462 (N_22462,N_20104,N_21189);
nand U22463 (N_22463,N_21922,N_20788);
or U22464 (N_22464,N_20356,N_20424);
xnor U22465 (N_22465,N_21827,N_21115);
or U22466 (N_22466,N_21384,N_20353);
nor U22467 (N_22467,N_20523,N_21181);
xnor U22468 (N_22468,N_20636,N_20077);
or U22469 (N_22469,N_20731,N_20697);
and U22470 (N_22470,N_21594,N_21793);
nand U22471 (N_22471,N_20872,N_21611);
xnor U22472 (N_22472,N_20571,N_20776);
nor U22473 (N_22473,N_20620,N_21671);
and U22474 (N_22474,N_21160,N_20345);
nand U22475 (N_22475,N_20527,N_20654);
nand U22476 (N_22476,N_21715,N_21299);
or U22477 (N_22477,N_20017,N_21502);
nand U22478 (N_22478,N_20292,N_21001);
nor U22479 (N_22479,N_21726,N_20735);
xnor U22480 (N_22480,N_20064,N_20905);
or U22481 (N_22481,N_20250,N_20750);
xnor U22482 (N_22482,N_21791,N_21832);
nor U22483 (N_22483,N_20166,N_21149);
xor U22484 (N_22484,N_21751,N_20032);
or U22485 (N_22485,N_20818,N_21893);
xor U22486 (N_22486,N_20033,N_20801);
nor U22487 (N_22487,N_20435,N_21528);
xnor U22488 (N_22488,N_21525,N_21283);
xnor U22489 (N_22489,N_21560,N_20036);
xor U22490 (N_22490,N_20153,N_21632);
and U22491 (N_22491,N_21821,N_20778);
and U22492 (N_22492,N_20682,N_20067);
nand U22493 (N_22493,N_20867,N_20057);
nor U22494 (N_22494,N_21864,N_20282);
or U22495 (N_22495,N_20066,N_20350);
nand U22496 (N_22496,N_21101,N_20309);
nand U22497 (N_22497,N_20374,N_20930);
nand U22498 (N_22498,N_21841,N_20593);
xor U22499 (N_22499,N_20065,N_20229);
and U22500 (N_22500,N_21110,N_20672);
nor U22501 (N_22501,N_20969,N_21714);
nor U22502 (N_22502,N_20420,N_20027);
and U22503 (N_22503,N_21621,N_20856);
nand U22504 (N_22504,N_20277,N_21612);
and U22505 (N_22505,N_21064,N_20155);
or U22506 (N_22506,N_20909,N_20737);
xor U22507 (N_22507,N_20611,N_20668);
xor U22508 (N_22508,N_21963,N_21288);
and U22509 (N_22509,N_20168,N_21277);
or U22510 (N_22510,N_20513,N_20307);
and U22511 (N_22511,N_20613,N_20308);
nand U22512 (N_22512,N_20953,N_21297);
nand U22513 (N_22513,N_20705,N_21578);
and U22514 (N_22514,N_20480,N_20156);
nand U22515 (N_22515,N_21810,N_21012);
and U22516 (N_22516,N_21099,N_20120);
and U22517 (N_22517,N_21378,N_20265);
or U22518 (N_22518,N_21010,N_20708);
nand U22519 (N_22519,N_21950,N_21720);
or U22520 (N_22520,N_21494,N_20667);
nor U22521 (N_22521,N_21426,N_20366);
and U22522 (N_22522,N_21834,N_20923);
nor U22523 (N_22523,N_21322,N_20699);
or U22524 (N_22524,N_20152,N_20791);
nand U22525 (N_22525,N_20249,N_20206);
or U22526 (N_22526,N_20371,N_21197);
and U22527 (N_22527,N_21417,N_21696);
nand U22528 (N_22528,N_20794,N_20902);
nand U22529 (N_22529,N_21904,N_21091);
or U22530 (N_22530,N_21135,N_20689);
or U22531 (N_22531,N_21296,N_20015);
and U22532 (N_22532,N_21677,N_20603);
xor U22533 (N_22533,N_21484,N_21165);
and U22534 (N_22534,N_21765,N_20564);
nor U22535 (N_22535,N_21457,N_21946);
and U22536 (N_22536,N_20108,N_20297);
xor U22537 (N_22537,N_20979,N_21349);
nand U22538 (N_22538,N_20355,N_20210);
or U22539 (N_22539,N_21456,N_21933);
or U22540 (N_22540,N_20001,N_21409);
and U22541 (N_22541,N_21952,N_20103);
nor U22542 (N_22542,N_20521,N_21262);
or U22543 (N_22543,N_20325,N_20068);
nand U22544 (N_22544,N_20565,N_21126);
or U22545 (N_22545,N_20952,N_21433);
or U22546 (N_22546,N_21216,N_21050);
or U22547 (N_22547,N_21208,N_21178);
or U22548 (N_22548,N_20442,N_21410);
or U22549 (N_22549,N_21850,N_20301);
and U22550 (N_22550,N_21673,N_20395);
nand U22551 (N_22551,N_21661,N_21615);
nand U22552 (N_22552,N_21200,N_21697);
and U22553 (N_22553,N_20853,N_20164);
and U22554 (N_22554,N_20400,N_20258);
and U22555 (N_22555,N_20272,N_21710);
or U22556 (N_22556,N_21177,N_20259);
xor U22557 (N_22557,N_21078,N_20002);
and U22558 (N_22558,N_21355,N_20112);
or U22559 (N_22559,N_20038,N_20640);
xnor U22560 (N_22560,N_21823,N_20910);
or U22561 (N_22561,N_20267,N_20929);
nand U22562 (N_22562,N_20762,N_20956);
xnor U22563 (N_22563,N_21972,N_21140);
nand U22564 (N_22564,N_20885,N_21680);
xor U22565 (N_22565,N_21981,N_21279);
nor U22566 (N_22566,N_20178,N_20752);
nand U22567 (N_22567,N_21746,N_20456);
and U22568 (N_22568,N_21994,N_21383);
and U22569 (N_22569,N_21337,N_21163);
xnor U22570 (N_22570,N_21267,N_21437);
and U22571 (N_22571,N_20641,N_20173);
nor U22572 (N_22572,N_21291,N_21837);
nor U22573 (N_22573,N_20866,N_20806);
xnor U22574 (N_22574,N_21176,N_21329);
xor U22575 (N_22575,N_20961,N_20115);
nor U22576 (N_22576,N_21553,N_21687);
nand U22577 (N_22577,N_20438,N_20753);
and U22578 (N_22578,N_20398,N_21421);
and U22579 (N_22579,N_20860,N_20485);
nand U22580 (N_22580,N_20423,N_20805);
and U22581 (N_22581,N_21102,N_21002);
nor U22582 (N_22582,N_20643,N_20870);
or U22583 (N_22583,N_21381,N_20865);
nor U22584 (N_22584,N_20963,N_20261);
nand U22585 (N_22585,N_20989,N_20903);
and U22586 (N_22586,N_21238,N_21838);
xor U22587 (N_22587,N_20882,N_20135);
xnor U22588 (N_22588,N_21138,N_21588);
nand U22589 (N_22589,N_21316,N_21650);
nand U22590 (N_22590,N_20647,N_21772);
xor U22591 (N_22591,N_21538,N_20471);
nand U22592 (N_22592,N_21495,N_21519);
or U22593 (N_22593,N_21188,N_21531);
or U22594 (N_22594,N_20907,N_21443);
nand U22595 (N_22595,N_21736,N_21319);
xor U22596 (N_22596,N_21805,N_21526);
and U22597 (N_22597,N_21127,N_20828);
nand U22598 (N_22598,N_20904,N_21435);
nor U22599 (N_22599,N_21705,N_20375);
and U22600 (N_22600,N_20123,N_20589);
nor U22601 (N_22601,N_20131,N_20202);
or U22602 (N_22602,N_20218,N_20650);
or U22603 (N_22603,N_21885,N_21712);
or U22604 (N_22604,N_20133,N_20772);
or U22605 (N_22605,N_21302,N_21828);
or U22606 (N_22606,N_21201,N_20421);
and U22607 (N_22607,N_21259,N_21324);
xnor U22608 (N_22608,N_21533,N_21341);
nand U22609 (N_22609,N_20086,N_20604);
nor U22610 (N_22610,N_20758,N_21924);
nand U22611 (N_22611,N_21501,N_20711);
and U22612 (N_22612,N_20417,N_21362);
xnor U22613 (N_22613,N_21980,N_21124);
nand U22614 (N_22614,N_20012,N_20854);
nor U22615 (N_22615,N_20434,N_20581);
xnor U22616 (N_22616,N_21662,N_20047);
nand U22617 (N_22617,N_20459,N_21226);
nor U22618 (N_22618,N_20657,N_20275);
or U22619 (N_22619,N_21482,N_20543);
xor U22620 (N_22620,N_21802,N_20841);
xnor U22621 (N_22621,N_20449,N_21956);
or U22622 (N_22622,N_21118,N_21385);
nor U22623 (N_22623,N_21121,N_21152);
nand U22624 (N_22624,N_20679,N_21327);
and U22625 (N_22625,N_20962,N_21874);
or U22626 (N_22626,N_21487,N_20266);
or U22627 (N_22627,N_20625,N_20814);
nor U22628 (N_22628,N_21913,N_20363);
nor U22629 (N_22629,N_20234,N_21451);
nor U22630 (N_22630,N_21067,N_20209);
and U22631 (N_22631,N_21190,N_20594);
nand U22632 (N_22632,N_20469,N_20161);
xnor U22633 (N_22633,N_21430,N_21087);
nor U22634 (N_22634,N_21942,N_21643);
nand U22635 (N_22635,N_20243,N_20078);
xor U22636 (N_22636,N_20172,N_20739);
xor U22637 (N_22637,N_20704,N_20959);
xnor U22638 (N_22638,N_20813,N_20329);
xnor U22639 (N_22639,N_21564,N_21745);
and U22640 (N_22640,N_20128,N_21007);
nor U22641 (N_22641,N_21318,N_20197);
or U22642 (N_22642,N_21624,N_21684);
nand U22643 (N_22643,N_21198,N_21086);
or U22644 (N_22644,N_21955,N_20239);
xnor U22645 (N_22645,N_21732,N_21785);
and U22646 (N_22646,N_21472,N_20496);
xnor U22647 (N_22647,N_21445,N_21754);
xor U22648 (N_22648,N_21308,N_20848);
and U22649 (N_22649,N_20121,N_21093);
or U22650 (N_22650,N_20221,N_21718);
xor U22651 (N_22651,N_21982,N_21787);
or U22652 (N_22652,N_21750,N_20857);
xor U22653 (N_22653,N_20132,N_20244);
nand U22654 (N_22654,N_21887,N_21788);
and U22655 (N_22655,N_20072,N_21411);
xnor U22656 (N_22656,N_20405,N_21089);
or U22657 (N_22657,N_21037,N_21071);
nand U22658 (N_22658,N_20285,N_20222);
xnor U22659 (N_22659,N_20409,N_20184);
or U22660 (N_22660,N_20312,N_21333);
nor U22661 (N_22661,N_20844,N_21249);
or U22662 (N_22662,N_20987,N_20730);
and U22663 (N_22663,N_20539,N_20700);
or U22664 (N_22664,N_21537,N_21915);
and U22665 (N_22665,N_21987,N_21100);
or U22666 (N_22666,N_20389,N_21088);
xnor U22667 (N_22667,N_21489,N_20076);
nand U22668 (N_22668,N_20945,N_20632);
xnor U22669 (N_22669,N_21599,N_20542);
or U22670 (N_22670,N_21660,N_21348);
nor U22671 (N_22671,N_20380,N_21630);
and U22672 (N_22672,N_20052,N_20985);
nand U22673 (N_22673,N_21610,N_21899);
or U22674 (N_22674,N_20475,N_21260);
and U22675 (N_22675,N_21773,N_21203);
nor U22676 (N_22676,N_20381,N_20660);
or U22677 (N_22677,N_21270,N_20414);
nand U22678 (N_22678,N_21377,N_20299);
nand U22679 (N_22679,N_21623,N_20744);
nand U22680 (N_22680,N_21326,N_20716);
nand U22681 (N_22681,N_21758,N_21452);
nand U22682 (N_22682,N_21524,N_21448);
nor U22683 (N_22683,N_20886,N_20916);
or U22684 (N_22684,N_20541,N_20418);
and U22685 (N_22685,N_21387,N_21586);
or U22686 (N_22686,N_20627,N_20608);
nor U22687 (N_22687,N_20302,N_21996);
nor U22688 (N_22688,N_21505,N_21449);
and U22689 (N_22689,N_20252,N_20326);
nand U22690 (N_22690,N_20586,N_21205);
or U22691 (N_22691,N_20673,N_21652);
and U22692 (N_22692,N_21566,N_21927);
nand U22693 (N_22693,N_20028,N_20812);
or U22694 (N_22694,N_21276,N_20093);
and U22695 (N_22695,N_21493,N_21511);
and U22696 (N_22696,N_21869,N_20492);
nand U22697 (N_22697,N_21770,N_20943);
or U22698 (N_22698,N_21320,N_21214);
nor U22699 (N_22699,N_20695,N_20743);
and U22700 (N_22700,N_21780,N_20724);
nor U22701 (N_22701,N_21851,N_20422);
or U22702 (N_22702,N_21336,N_20733);
nor U22703 (N_22703,N_20528,N_21595);
and U22704 (N_22704,N_21183,N_21353);
nand U22705 (N_22705,N_20494,N_21029);
xor U22706 (N_22706,N_21399,N_21548);
and U22707 (N_22707,N_21325,N_20119);
nand U22708 (N_22708,N_20215,N_21485);
or U22709 (N_22709,N_20298,N_20538);
nand U22710 (N_22710,N_21413,N_21882);
nand U22711 (N_22711,N_21068,N_21460);
or U22712 (N_22712,N_21453,N_21764);
nor U22713 (N_22713,N_21343,N_20054);
or U22714 (N_22714,N_21629,N_21339);
nor U22715 (N_22715,N_21605,N_21053);
nor U22716 (N_22716,N_20384,N_20563);
or U22717 (N_22717,N_21041,N_21006);
nand U22718 (N_22718,N_20341,N_20639);
or U22719 (N_22719,N_21762,N_21574);
and U22720 (N_22720,N_21782,N_21455);
nor U22721 (N_22721,N_21579,N_21306);
or U22722 (N_22722,N_21234,N_20317);
and U22723 (N_22723,N_20430,N_21859);
or U22724 (N_22724,N_20493,N_20330);
xnor U22725 (N_22725,N_20488,N_21964);
nor U22726 (N_22726,N_20313,N_21365);
or U22727 (N_22727,N_21757,N_20195);
nand U22728 (N_22728,N_20553,N_21597);
nor U22729 (N_22729,N_20284,N_20827);
or U22730 (N_22730,N_21728,N_20440);
or U22731 (N_22731,N_20633,N_20096);
nor U22732 (N_22732,N_21976,N_20050);
nor U22733 (N_22733,N_21862,N_21978);
xor U22734 (N_22734,N_21763,N_20214);
nand U22735 (N_22735,N_21951,N_20014);
nor U22736 (N_22736,N_20127,N_20470);
nand U22737 (N_22737,N_20372,N_20659);
nor U22738 (N_22738,N_21930,N_21253);
nor U22739 (N_22739,N_21542,N_21983);
and U22740 (N_22740,N_20083,N_20331);
nand U22741 (N_22741,N_20759,N_20707);
nor U22742 (N_22742,N_20775,N_21458);
nand U22743 (N_22743,N_20925,N_20136);
nor U22744 (N_22744,N_21268,N_21988);
xnor U22745 (N_22745,N_21321,N_21065);
or U22746 (N_22746,N_21962,N_21569);
nand U22747 (N_22747,N_21475,N_20893);
and U22748 (N_22748,N_21027,N_20815);
and U22749 (N_22749,N_21108,N_20763);
nand U22750 (N_22750,N_20091,N_21116);
nor U22751 (N_22751,N_20179,N_20450);
nand U22752 (N_22752,N_20287,N_21948);
or U22753 (N_22753,N_20201,N_20957);
nand U22754 (N_22754,N_21017,N_20506);
and U22755 (N_22755,N_21379,N_20383);
and U22756 (N_22756,N_20599,N_20468);
xor U22757 (N_22757,N_20830,N_20831);
and U22758 (N_22758,N_20410,N_21225);
nor U22759 (N_22759,N_21243,N_20208);
or U22760 (N_22760,N_21394,N_20691);
nand U22761 (N_22761,N_20922,N_21820);
nand U22762 (N_22762,N_21144,N_21796);
xnor U22763 (N_22763,N_20680,N_20694);
nor U22764 (N_22764,N_21704,N_21019);
or U22765 (N_22765,N_21779,N_20924);
nand U22766 (N_22766,N_20304,N_21184);
or U22767 (N_22767,N_21228,N_21508);
and U22768 (N_22768,N_20392,N_20585);
xnor U22769 (N_22769,N_20509,N_21162);
nand U22770 (N_22770,N_21692,N_21999);
nor U22771 (N_22771,N_20836,N_21989);
nand U22772 (N_22772,N_21881,N_20990);
nand U22773 (N_22773,N_20873,N_20367);
and U22774 (N_22774,N_20457,N_21717);
and U22775 (N_22775,N_21748,N_21210);
or U22776 (N_22776,N_21724,N_21233);
and U22777 (N_22777,N_21264,N_20013);
nand U22778 (N_22778,N_20941,N_21808);
or U22779 (N_22779,N_20800,N_21731);
nor U22780 (N_22780,N_21098,N_20991);
and U22781 (N_22781,N_21369,N_21938);
and U22782 (N_22782,N_20432,N_20192);
xor U22783 (N_22783,N_20255,N_21496);
nand U22784 (N_22784,N_20992,N_21676);
nor U22785 (N_22785,N_21192,N_20761);
xor U22786 (N_22786,N_20021,N_20646);
nor U22787 (N_22787,N_21809,N_20338);
nor U22788 (N_22788,N_20176,N_20408);
xor U22789 (N_22789,N_21722,N_21568);
nand U22790 (N_22790,N_21741,N_21713);
and U22791 (N_22791,N_21657,N_21402);
nor U22792 (N_22792,N_20535,N_21251);
nor U22793 (N_22793,N_20437,N_21171);
xor U22794 (N_22794,N_20246,N_21439);
nor U22795 (N_22795,N_20634,N_21263);
and U22796 (N_22796,N_20071,N_20549);
nor U22797 (N_22797,N_20029,N_21674);
nor U22798 (N_22798,N_21853,N_20566);
nor U22799 (N_22799,N_21622,N_21755);
nand U22800 (N_22800,N_20685,N_21506);
and U22801 (N_22801,N_21317,N_21016);
and U22802 (N_22802,N_20675,N_20182);
and U22803 (N_22803,N_21166,N_21949);
or U22804 (N_22804,N_20466,N_21156);
nand U22805 (N_22805,N_20648,N_21066);
nor U22806 (N_22806,N_21403,N_21642);
and U22807 (N_22807,N_21105,N_21953);
nand U22808 (N_22808,N_20725,N_21768);
and U22809 (N_22809,N_21825,N_20661);
and U22810 (N_22810,N_21619,N_20785);
and U22811 (N_22811,N_20555,N_21393);
xor U22812 (N_22812,N_21023,N_20973);
nor U22813 (N_22813,N_20968,N_20847);
and U22814 (N_22814,N_21235,N_21971);
nand U22815 (N_22815,N_21258,N_21310);
or U22816 (N_22816,N_20245,N_20237);
nand U22817 (N_22817,N_21058,N_20995);
and U22818 (N_22818,N_20134,N_20254);
nor U22819 (N_22819,N_20248,N_20177);
and U22820 (N_22820,N_20278,N_21563);
or U22821 (N_22821,N_20983,N_21406);
or U22822 (N_22822,N_20165,N_20948);
or U22823 (N_22823,N_21499,N_21350);
or U22824 (N_22824,N_21541,N_21392);
and U22825 (N_22825,N_20257,N_21169);
nand U22826 (N_22826,N_21824,N_21261);
nand U22827 (N_22827,N_20887,N_21592);
nor U22828 (N_22828,N_21540,N_20562);
and U22829 (N_22829,N_20757,N_20918);
and U22830 (N_22830,N_21051,N_20099);
nor U22831 (N_22831,N_21282,N_20692);
or U22832 (N_22832,N_21048,N_21551);
nor U22833 (N_22833,N_20554,N_20415);
nor U22834 (N_22834,N_20062,N_20391);
nand U22835 (N_22835,N_21040,N_20514);
nor U22836 (N_22836,N_20869,N_21846);
or U22837 (N_22837,N_21556,N_21602);
or U22838 (N_22838,N_20368,N_20747);
nor U22839 (N_22839,N_21968,N_21514);
and U22840 (N_22840,N_20412,N_21220);
xnor U22841 (N_22841,N_21675,N_20670);
and U22842 (N_22842,N_20999,N_21199);
or U22843 (N_22843,N_21257,N_20041);
xor U22844 (N_22844,N_20264,N_21295);
nor U22845 (N_22845,N_21275,N_20053);
nand U22846 (N_22846,N_20186,N_20706);
xnor U22847 (N_22847,N_21966,N_21906);
nand U22848 (N_22848,N_21332,N_21154);
or U22849 (N_22849,N_20798,N_21425);
nor U22850 (N_22850,N_20516,N_21239);
nor U22851 (N_22851,N_21298,N_20515);
nand U22852 (N_22852,N_20734,N_20721);
xor U22853 (N_22853,N_21031,N_20635);
and U22854 (N_22854,N_21009,N_20588);
nand U22855 (N_22855,N_21370,N_20198);
xnor U22856 (N_22856,N_21975,N_21271);
xnor U22857 (N_22857,N_20106,N_21559);
nand U22858 (N_22858,N_20270,N_20951);
or U22859 (N_22859,N_20445,N_21872);
xnor U22860 (N_22860,N_20880,N_20247);
or U22861 (N_22861,N_21822,N_20169);
or U22862 (N_22862,N_20584,N_21481);
nor U22863 (N_22863,N_20942,N_20011);
and U22864 (N_22864,N_20360,N_20043);
xnor U22865 (N_22865,N_20138,N_20587);
xnor U22866 (N_22866,N_21133,N_20532);
or U22867 (N_22867,N_20986,N_20779);
or U22868 (N_22868,N_21587,N_20727);
nand U22869 (N_22869,N_21079,N_20386);
xnor U22870 (N_22870,N_21840,N_20296);
or U22871 (N_22871,N_20080,N_20793);
xnor U22872 (N_22872,N_20876,N_21527);
and U22873 (N_22873,N_20101,N_20037);
or U22874 (N_22874,N_20771,N_21567);
nor U22875 (N_22875,N_20863,N_21723);
or U22876 (N_22876,N_20974,N_21498);
and U22877 (N_22877,N_21918,N_21617);
xnor U22878 (N_22878,N_21468,N_20766);
nand U22879 (N_22879,N_20328,N_20850);
or U22880 (N_22880,N_21145,N_20955);
nand U22881 (N_22881,N_20097,N_21075);
xnor U22882 (N_22882,N_20825,N_21925);
nand U22883 (N_22883,N_21794,N_21637);
and U22884 (N_22884,N_20362,N_20482);
nand U22885 (N_22885,N_20467,N_21047);
nor U22886 (N_22886,N_21008,N_21848);
and U22887 (N_22887,N_20874,N_20070);
nor U22888 (N_22888,N_21691,N_20652);
and U22889 (N_22889,N_20760,N_21491);
xor U22890 (N_22890,N_20323,N_21777);
nand U22891 (N_22891,N_21917,N_21081);
and U22892 (N_22892,N_20804,N_21583);
or U22893 (N_22893,N_21706,N_21191);
nand U22894 (N_22894,N_20666,N_20157);
nand U22895 (N_22895,N_20609,N_20035);
nor U22896 (N_22896,N_21929,N_21781);
or U22897 (N_22897,N_20126,N_20061);
nor U22898 (N_22898,N_20754,N_20117);
or U22899 (N_22899,N_21878,N_21155);
or U22900 (N_22900,N_20900,N_20612);
or U22901 (N_22901,N_20276,N_21046);
xnor U22902 (N_22902,N_21530,N_20578);
nor U22903 (N_22903,N_20009,N_21404);
nand U22904 (N_22904,N_20561,N_20742);
nor U22905 (N_22905,N_20413,N_20303);
nand U22906 (N_22906,N_21725,N_21186);
nor U22907 (N_22907,N_20411,N_21585);
nor U22908 (N_22908,N_21516,N_20300);
and U22909 (N_22909,N_21935,N_20786);
nand U22910 (N_22910,N_21860,N_20114);
and U22911 (N_22911,N_21217,N_20755);
nor U22912 (N_22912,N_21792,N_21227);
nor U22913 (N_22913,N_20511,N_21616);
and U22914 (N_22914,N_20216,N_20146);
or U22915 (N_22915,N_21734,N_21589);
nor U22916 (N_22916,N_21374,N_20406);
xor U22917 (N_22917,N_21063,N_21908);
nand U22918 (N_22918,N_21323,N_21414);
nor U22919 (N_22919,N_21222,N_21856);
nor U22920 (N_22920,N_21655,N_20004);
nand U22921 (N_22921,N_21884,N_21117);
nand U22922 (N_22922,N_21497,N_20590);
or U22923 (N_22923,N_21342,N_21431);
and U22924 (N_22924,N_21829,N_21613);
nor U22925 (N_22925,N_21179,N_20556);
xor U22926 (N_22926,N_20919,N_21103);
nor U22927 (N_22927,N_21905,N_20619);
nor U22928 (N_22928,N_21591,N_21011);
and U22929 (N_22929,N_20518,N_21863);
nor U22930 (N_22930,N_20592,N_20049);
nor U22931 (N_22931,N_20348,N_20191);
or U22932 (N_22932,N_20160,N_20950);
xnor U22933 (N_22933,N_21819,N_20333);
or U22934 (N_22934,N_20462,N_21576);
and U22935 (N_22935,N_20936,N_21931);
xnor U22936 (N_22936,N_20939,N_21743);
xnor U22937 (N_22937,N_21954,N_21609);
or U22938 (N_22938,N_20118,N_20629);
and U22939 (N_22939,N_21112,N_20148);
or U22940 (N_22940,N_21888,N_20545);
nor U22941 (N_22941,N_20233,N_21620);
nand U22942 (N_22942,N_21215,N_20399);
and U22943 (N_22943,N_21573,N_21386);
xnor U22944 (N_22944,N_20810,N_20008);
and U22945 (N_22945,N_21464,N_21420);
and U22946 (N_22946,N_20428,N_20489);
xnor U22947 (N_22947,N_21669,N_20344);
xor U22948 (N_22948,N_21666,N_21128);
nand U22949 (N_22949,N_21026,N_21847);
or U22950 (N_22950,N_21405,N_20124);
nand U22951 (N_22951,N_20686,N_20783);
xnor U22952 (N_22952,N_20407,N_21072);
and U22953 (N_22953,N_21584,N_20427);
or U22954 (N_22954,N_21936,N_21886);
or U22955 (N_22955,N_21997,N_21778);
nor U22956 (N_22956,N_20145,N_21470);
nor U22957 (N_22957,N_20217,N_20795);
nand U22958 (N_22958,N_20624,N_21146);
nand U22959 (N_22959,N_21678,N_20477);
and U22960 (N_22960,N_20451,N_21842);
or U22961 (N_22961,N_21536,N_21250);
or U22962 (N_22962,N_21024,N_21285);
nor U22963 (N_22963,N_21945,N_21213);
and U22964 (N_22964,N_20895,N_21668);
nor U22965 (N_22965,N_20322,N_21518);
and U22966 (N_22966,N_20949,N_21025);
or U22967 (N_22967,N_21914,N_21328);
or U22968 (N_22968,N_20171,N_20039);
and U22969 (N_22969,N_20051,N_21890);
and U22970 (N_22970,N_21314,N_20714);
or U22971 (N_22971,N_21909,N_20212);
or U22972 (N_22972,N_20337,N_20799);
nand U22973 (N_22973,N_21695,N_20723);
and U22974 (N_22974,N_21005,N_21419);
nand U22975 (N_22975,N_20965,N_21371);
nand U22976 (N_22976,N_21360,N_20972);
xor U22977 (N_22977,N_21391,N_21651);
nand U22978 (N_22978,N_20213,N_20975);
nand U22979 (N_22979,N_21196,N_20081);
and U22980 (N_22980,N_21803,N_21480);
and U22981 (N_22981,N_21626,N_21790);
and U22982 (N_22982,N_21219,N_20340);
nand U22983 (N_22983,N_20291,N_20085);
xnor U22984 (N_22984,N_20336,N_21114);
nor U22985 (N_22985,N_21422,N_20207);
nand U22986 (N_22986,N_21663,N_20678);
or U22987 (N_22987,N_20125,N_21357);
or U22988 (N_22988,N_21459,N_21492);
xnor U22989 (N_22989,N_21441,N_20040);
nand U22990 (N_22990,N_21136,N_21682);
nor U22991 (N_22991,N_21721,N_20446);
nand U22992 (N_22992,N_20448,N_20228);
xor U22993 (N_22993,N_20003,N_20908);
nor U22994 (N_22994,N_21634,N_21901);
or U22995 (N_22995,N_21686,N_20557);
nor U22996 (N_22996,N_21889,N_20807);
nand U22997 (N_22997,N_21639,N_20823);
and U22998 (N_22998,N_21003,N_20225);
nand U22999 (N_22999,N_21535,N_21625);
or U23000 (N_23000,N_21917,N_20885);
nor U23001 (N_23001,N_21436,N_20277);
xor U23002 (N_23002,N_20958,N_20213);
nor U23003 (N_23003,N_20431,N_21066);
xor U23004 (N_23004,N_21377,N_21965);
or U23005 (N_23005,N_20354,N_21533);
or U23006 (N_23006,N_20455,N_21537);
nor U23007 (N_23007,N_20470,N_21931);
nor U23008 (N_23008,N_21153,N_20156);
and U23009 (N_23009,N_21622,N_20290);
nand U23010 (N_23010,N_21320,N_20921);
nor U23011 (N_23011,N_21141,N_20529);
or U23012 (N_23012,N_20717,N_20643);
xor U23013 (N_23013,N_20416,N_21985);
nand U23014 (N_23014,N_20593,N_20555);
and U23015 (N_23015,N_20621,N_20491);
or U23016 (N_23016,N_21948,N_20992);
xor U23017 (N_23017,N_20935,N_20488);
nor U23018 (N_23018,N_21807,N_20501);
xnor U23019 (N_23019,N_20159,N_21841);
or U23020 (N_23020,N_20372,N_21150);
or U23021 (N_23021,N_20164,N_21699);
or U23022 (N_23022,N_21540,N_20367);
xor U23023 (N_23023,N_21879,N_21562);
nand U23024 (N_23024,N_20918,N_21964);
or U23025 (N_23025,N_20693,N_21255);
nor U23026 (N_23026,N_21911,N_21332);
and U23027 (N_23027,N_20973,N_21442);
xor U23028 (N_23028,N_21371,N_20171);
nand U23029 (N_23029,N_21239,N_20197);
nand U23030 (N_23030,N_21067,N_21856);
and U23031 (N_23031,N_20813,N_20373);
xnor U23032 (N_23032,N_20608,N_21595);
xor U23033 (N_23033,N_20327,N_21273);
and U23034 (N_23034,N_21510,N_20849);
and U23035 (N_23035,N_21813,N_20876);
xnor U23036 (N_23036,N_20552,N_21097);
xor U23037 (N_23037,N_21583,N_20770);
or U23038 (N_23038,N_20621,N_21217);
or U23039 (N_23039,N_20543,N_20395);
xnor U23040 (N_23040,N_21973,N_20668);
and U23041 (N_23041,N_21164,N_21888);
xnor U23042 (N_23042,N_20330,N_20537);
and U23043 (N_23043,N_20019,N_20284);
nor U23044 (N_23044,N_21323,N_20125);
or U23045 (N_23045,N_20572,N_20404);
nor U23046 (N_23046,N_21914,N_21101);
or U23047 (N_23047,N_21171,N_21595);
nor U23048 (N_23048,N_21109,N_21621);
and U23049 (N_23049,N_20485,N_21038);
xnor U23050 (N_23050,N_21488,N_20753);
or U23051 (N_23051,N_20725,N_21736);
nor U23052 (N_23052,N_21272,N_20463);
nor U23053 (N_23053,N_20529,N_21522);
xor U23054 (N_23054,N_21621,N_21805);
xor U23055 (N_23055,N_20174,N_21115);
and U23056 (N_23056,N_21068,N_20883);
nand U23057 (N_23057,N_20629,N_21455);
xnor U23058 (N_23058,N_20787,N_21043);
or U23059 (N_23059,N_21373,N_21700);
nand U23060 (N_23060,N_21272,N_20986);
xor U23061 (N_23061,N_20874,N_21513);
or U23062 (N_23062,N_21950,N_21589);
or U23063 (N_23063,N_21836,N_20942);
nor U23064 (N_23064,N_20037,N_21791);
and U23065 (N_23065,N_20869,N_21954);
nand U23066 (N_23066,N_21854,N_20113);
and U23067 (N_23067,N_21453,N_21693);
or U23068 (N_23068,N_20386,N_20350);
or U23069 (N_23069,N_21545,N_21441);
xor U23070 (N_23070,N_21252,N_20749);
or U23071 (N_23071,N_20282,N_20668);
nor U23072 (N_23072,N_20741,N_21444);
or U23073 (N_23073,N_21965,N_21727);
nand U23074 (N_23074,N_21393,N_20039);
xor U23075 (N_23075,N_21840,N_21675);
and U23076 (N_23076,N_20935,N_20609);
nand U23077 (N_23077,N_21646,N_21540);
nand U23078 (N_23078,N_21863,N_20852);
and U23079 (N_23079,N_21462,N_20827);
nor U23080 (N_23080,N_21808,N_20469);
and U23081 (N_23081,N_20604,N_21397);
xor U23082 (N_23082,N_20299,N_20079);
nor U23083 (N_23083,N_20601,N_21318);
nor U23084 (N_23084,N_20661,N_21915);
and U23085 (N_23085,N_21748,N_21291);
xnor U23086 (N_23086,N_21109,N_21461);
nor U23087 (N_23087,N_20347,N_20801);
nor U23088 (N_23088,N_21673,N_21330);
or U23089 (N_23089,N_21721,N_20098);
and U23090 (N_23090,N_20858,N_21134);
xor U23091 (N_23091,N_20253,N_21856);
nand U23092 (N_23092,N_21654,N_20629);
xnor U23093 (N_23093,N_20682,N_20714);
nor U23094 (N_23094,N_21648,N_20853);
xor U23095 (N_23095,N_20297,N_20258);
xor U23096 (N_23096,N_20469,N_21991);
nand U23097 (N_23097,N_21565,N_20252);
xnor U23098 (N_23098,N_21820,N_21378);
xnor U23099 (N_23099,N_20789,N_20640);
nand U23100 (N_23100,N_20551,N_20619);
and U23101 (N_23101,N_21401,N_21787);
xnor U23102 (N_23102,N_21891,N_20584);
and U23103 (N_23103,N_20086,N_20659);
or U23104 (N_23104,N_21085,N_20832);
nor U23105 (N_23105,N_20703,N_20752);
or U23106 (N_23106,N_20533,N_21155);
or U23107 (N_23107,N_20838,N_20037);
xnor U23108 (N_23108,N_20517,N_20506);
nor U23109 (N_23109,N_21619,N_21016);
nor U23110 (N_23110,N_21032,N_20330);
nand U23111 (N_23111,N_20558,N_20496);
nand U23112 (N_23112,N_20389,N_21754);
xnor U23113 (N_23113,N_21151,N_21220);
nand U23114 (N_23114,N_21758,N_20615);
xor U23115 (N_23115,N_20413,N_20468);
and U23116 (N_23116,N_20708,N_20720);
nand U23117 (N_23117,N_21380,N_21053);
xor U23118 (N_23118,N_21616,N_21589);
nor U23119 (N_23119,N_20419,N_21686);
and U23120 (N_23120,N_21839,N_21665);
nand U23121 (N_23121,N_21484,N_21865);
nor U23122 (N_23122,N_20900,N_21106);
nand U23123 (N_23123,N_20824,N_21055);
and U23124 (N_23124,N_21526,N_20722);
and U23125 (N_23125,N_20457,N_20945);
xor U23126 (N_23126,N_20001,N_21383);
nor U23127 (N_23127,N_21921,N_20132);
nor U23128 (N_23128,N_21112,N_20800);
or U23129 (N_23129,N_20911,N_20959);
and U23130 (N_23130,N_21572,N_21337);
and U23131 (N_23131,N_21147,N_20082);
and U23132 (N_23132,N_21373,N_20190);
or U23133 (N_23133,N_21130,N_21482);
nor U23134 (N_23134,N_20373,N_21440);
nor U23135 (N_23135,N_21229,N_20779);
nand U23136 (N_23136,N_21121,N_20532);
nand U23137 (N_23137,N_20745,N_20071);
or U23138 (N_23138,N_20039,N_21454);
xor U23139 (N_23139,N_20186,N_20307);
nand U23140 (N_23140,N_21372,N_21714);
or U23141 (N_23141,N_20621,N_21546);
nand U23142 (N_23142,N_20498,N_21812);
and U23143 (N_23143,N_20414,N_20880);
nor U23144 (N_23144,N_20085,N_20904);
xnor U23145 (N_23145,N_21517,N_21505);
and U23146 (N_23146,N_20164,N_21147);
or U23147 (N_23147,N_21836,N_20497);
nand U23148 (N_23148,N_21045,N_21561);
nor U23149 (N_23149,N_21305,N_20322);
or U23150 (N_23150,N_20590,N_20631);
xor U23151 (N_23151,N_20044,N_20887);
or U23152 (N_23152,N_21859,N_21975);
and U23153 (N_23153,N_21095,N_21313);
nand U23154 (N_23154,N_20489,N_20881);
or U23155 (N_23155,N_20275,N_21224);
and U23156 (N_23156,N_21120,N_20069);
and U23157 (N_23157,N_21265,N_21913);
nand U23158 (N_23158,N_20422,N_21889);
nor U23159 (N_23159,N_20567,N_20998);
nor U23160 (N_23160,N_21034,N_21597);
or U23161 (N_23161,N_20559,N_20938);
nor U23162 (N_23162,N_21938,N_20613);
nor U23163 (N_23163,N_21319,N_20008);
or U23164 (N_23164,N_20552,N_20574);
nor U23165 (N_23165,N_21921,N_21756);
nor U23166 (N_23166,N_20315,N_21744);
and U23167 (N_23167,N_21781,N_21163);
or U23168 (N_23168,N_21758,N_20100);
xor U23169 (N_23169,N_20434,N_20284);
nand U23170 (N_23170,N_20178,N_21985);
nor U23171 (N_23171,N_20006,N_20471);
and U23172 (N_23172,N_21982,N_21805);
xnor U23173 (N_23173,N_21433,N_20520);
or U23174 (N_23174,N_20269,N_21985);
or U23175 (N_23175,N_21250,N_21676);
nor U23176 (N_23176,N_20572,N_20110);
xor U23177 (N_23177,N_20431,N_20628);
xor U23178 (N_23178,N_20217,N_20299);
nand U23179 (N_23179,N_20437,N_21767);
and U23180 (N_23180,N_21696,N_21631);
nand U23181 (N_23181,N_21327,N_20920);
or U23182 (N_23182,N_20877,N_21771);
or U23183 (N_23183,N_21699,N_21774);
nand U23184 (N_23184,N_20886,N_20861);
nor U23185 (N_23185,N_20837,N_20013);
nor U23186 (N_23186,N_21174,N_21131);
nor U23187 (N_23187,N_21139,N_21769);
or U23188 (N_23188,N_20524,N_20150);
nor U23189 (N_23189,N_20207,N_21164);
nand U23190 (N_23190,N_21821,N_20301);
or U23191 (N_23191,N_21477,N_21845);
nand U23192 (N_23192,N_21822,N_20484);
nand U23193 (N_23193,N_20545,N_20239);
nor U23194 (N_23194,N_21915,N_21362);
or U23195 (N_23195,N_21512,N_21536);
xor U23196 (N_23196,N_21417,N_21250);
and U23197 (N_23197,N_21476,N_21266);
nand U23198 (N_23198,N_20763,N_20641);
nand U23199 (N_23199,N_20979,N_21709);
nand U23200 (N_23200,N_21842,N_20015);
xnor U23201 (N_23201,N_20537,N_21813);
nor U23202 (N_23202,N_21898,N_21309);
nor U23203 (N_23203,N_21235,N_21026);
nand U23204 (N_23204,N_20393,N_20523);
nor U23205 (N_23205,N_20797,N_21595);
and U23206 (N_23206,N_20539,N_21179);
nand U23207 (N_23207,N_20859,N_21802);
and U23208 (N_23208,N_21549,N_21107);
xor U23209 (N_23209,N_20037,N_20088);
nand U23210 (N_23210,N_20612,N_21537);
nand U23211 (N_23211,N_21600,N_20727);
nand U23212 (N_23212,N_20198,N_21974);
nand U23213 (N_23213,N_20233,N_20935);
or U23214 (N_23214,N_20754,N_20751);
and U23215 (N_23215,N_21275,N_20704);
and U23216 (N_23216,N_21719,N_21263);
xnor U23217 (N_23217,N_20992,N_20127);
nand U23218 (N_23218,N_21481,N_20517);
xor U23219 (N_23219,N_20471,N_21242);
nand U23220 (N_23220,N_21941,N_21569);
nor U23221 (N_23221,N_21185,N_21925);
or U23222 (N_23222,N_21907,N_21692);
and U23223 (N_23223,N_20522,N_20891);
or U23224 (N_23224,N_21689,N_21072);
or U23225 (N_23225,N_21225,N_21226);
or U23226 (N_23226,N_20764,N_21133);
or U23227 (N_23227,N_20773,N_20845);
xnor U23228 (N_23228,N_20474,N_21672);
nor U23229 (N_23229,N_20246,N_21981);
nand U23230 (N_23230,N_21693,N_21021);
and U23231 (N_23231,N_21323,N_20701);
xor U23232 (N_23232,N_21843,N_20402);
xor U23233 (N_23233,N_20311,N_21256);
nand U23234 (N_23234,N_20852,N_20126);
nor U23235 (N_23235,N_21026,N_21577);
xor U23236 (N_23236,N_21253,N_20878);
nor U23237 (N_23237,N_20211,N_20161);
nor U23238 (N_23238,N_20100,N_21440);
and U23239 (N_23239,N_21236,N_20182);
and U23240 (N_23240,N_21443,N_20414);
or U23241 (N_23241,N_20847,N_21787);
and U23242 (N_23242,N_20742,N_21655);
xor U23243 (N_23243,N_21270,N_20773);
and U23244 (N_23244,N_20855,N_21896);
and U23245 (N_23245,N_21721,N_20633);
and U23246 (N_23246,N_20760,N_20032);
and U23247 (N_23247,N_21998,N_20553);
nand U23248 (N_23248,N_20519,N_20077);
and U23249 (N_23249,N_20487,N_20129);
nor U23250 (N_23250,N_21655,N_20317);
or U23251 (N_23251,N_21502,N_21010);
and U23252 (N_23252,N_20102,N_21589);
nor U23253 (N_23253,N_20726,N_21978);
and U23254 (N_23254,N_21818,N_20337);
and U23255 (N_23255,N_20776,N_20628);
nand U23256 (N_23256,N_21895,N_20454);
xnor U23257 (N_23257,N_20414,N_21774);
nand U23258 (N_23258,N_21011,N_20838);
and U23259 (N_23259,N_20490,N_20483);
nand U23260 (N_23260,N_20894,N_21811);
or U23261 (N_23261,N_20239,N_20868);
and U23262 (N_23262,N_20257,N_20024);
and U23263 (N_23263,N_21153,N_20026);
nand U23264 (N_23264,N_20702,N_20395);
and U23265 (N_23265,N_21659,N_21316);
nand U23266 (N_23266,N_20195,N_21342);
or U23267 (N_23267,N_21678,N_21022);
or U23268 (N_23268,N_21269,N_21719);
and U23269 (N_23269,N_20603,N_21631);
xnor U23270 (N_23270,N_20738,N_21829);
xor U23271 (N_23271,N_20146,N_21016);
or U23272 (N_23272,N_21013,N_21829);
nand U23273 (N_23273,N_20494,N_21540);
xnor U23274 (N_23274,N_20575,N_21029);
nand U23275 (N_23275,N_21090,N_20843);
and U23276 (N_23276,N_21481,N_21659);
or U23277 (N_23277,N_21457,N_20168);
xor U23278 (N_23278,N_21780,N_20550);
nor U23279 (N_23279,N_21071,N_20456);
and U23280 (N_23280,N_20348,N_21106);
nand U23281 (N_23281,N_21325,N_21475);
and U23282 (N_23282,N_21459,N_20936);
or U23283 (N_23283,N_20706,N_21209);
and U23284 (N_23284,N_21355,N_21514);
xor U23285 (N_23285,N_20327,N_20308);
xnor U23286 (N_23286,N_20104,N_20441);
nand U23287 (N_23287,N_21306,N_20155);
nor U23288 (N_23288,N_21517,N_20337);
or U23289 (N_23289,N_20528,N_20427);
xor U23290 (N_23290,N_21882,N_21989);
nor U23291 (N_23291,N_20901,N_20567);
or U23292 (N_23292,N_21191,N_21176);
nor U23293 (N_23293,N_21716,N_20876);
nor U23294 (N_23294,N_20787,N_21072);
xnor U23295 (N_23295,N_20709,N_21881);
and U23296 (N_23296,N_20775,N_21443);
or U23297 (N_23297,N_21752,N_21588);
nand U23298 (N_23298,N_20320,N_21574);
and U23299 (N_23299,N_20103,N_21280);
nor U23300 (N_23300,N_21867,N_21241);
nand U23301 (N_23301,N_21651,N_20228);
nand U23302 (N_23302,N_20734,N_21872);
nor U23303 (N_23303,N_20875,N_20517);
nand U23304 (N_23304,N_20618,N_21732);
xor U23305 (N_23305,N_21055,N_20406);
xnor U23306 (N_23306,N_20460,N_21467);
nor U23307 (N_23307,N_21967,N_20555);
xor U23308 (N_23308,N_20767,N_20315);
or U23309 (N_23309,N_20242,N_20724);
xnor U23310 (N_23310,N_21471,N_21902);
and U23311 (N_23311,N_20647,N_20383);
nand U23312 (N_23312,N_20191,N_21148);
xor U23313 (N_23313,N_20194,N_21640);
nor U23314 (N_23314,N_21356,N_21810);
nor U23315 (N_23315,N_20725,N_20095);
nand U23316 (N_23316,N_20681,N_20612);
or U23317 (N_23317,N_20551,N_20025);
nor U23318 (N_23318,N_20735,N_20044);
nand U23319 (N_23319,N_20938,N_20824);
nor U23320 (N_23320,N_21824,N_20678);
or U23321 (N_23321,N_21873,N_21839);
and U23322 (N_23322,N_20756,N_20702);
xnor U23323 (N_23323,N_20928,N_20576);
and U23324 (N_23324,N_20827,N_21808);
or U23325 (N_23325,N_21165,N_20725);
nor U23326 (N_23326,N_21636,N_21766);
xnor U23327 (N_23327,N_21393,N_21987);
nand U23328 (N_23328,N_21528,N_21847);
or U23329 (N_23329,N_20486,N_21813);
and U23330 (N_23330,N_21249,N_21461);
or U23331 (N_23331,N_21168,N_20895);
xor U23332 (N_23332,N_20317,N_21631);
xnor U23333 (N_23333,N_21913,N_21854);
and U23334 (N_23334,N_21387,N_21832);
xor U23335 (N_23335,N_20479,N_21187);
nand U23336 (N_23336,N_20415,N_21827);
nor U23337 (N_23337,N_21102,N_20623);
or U23338 (N_23338,N_21388,N_21121);
nor U23339 (N_23339,N_20760,N_20544);
or U23340 (N_23340,N_21844,N_21369);
or U23341 (N_23341,N_21340,N_20889);
xor U23342 (N_23342,N_20652,N_21348);
xor U23343 (N_23343,N_21717,N_20641);
and U23344 (N_23344,N_21037,N_20434);
xnor U23345 (N_23345,N_21017,N_21689);
xor U23346 (N_23346,N_21590,N_21674);
nand U23347 (N_23347,N_21000,N_20834);
xnor U23348 (N_23348,N_21718,N_20320);
xnor U23349 (N_23349,N_21382,N_20395);
xnor U23350 (N_23350,N_21887,N_20167);
nor U23351 (N_23351,N_20560,N_20835);
nand U23352 (N_23352,N_21338,N_20561);
or U23353 (N_23353,N_20697,N_20711);
nand U23354 (N_23354,N_21717,N_21427);
nand U23355 (N_23355,N_21945,N_20900);
nor U23356 (N_23356,N_20735,N_21067);
xnor U23357 (N_23357,N_20812,N_21000);
and U23358 (N_23358,N_21637,N_20745);
nor U23359 (N_23359,N_21544,N_21992);
nor U23360 (N_23360,N_20778,N_21961);
nand U23361 (N_23361,N_21924,N_20658);
or U23362 (N_23362,N_21403,N_20966);
xnor U23363 (N_23363,N_20690,N_20495);
nor U23364 (N_23364,N_21861,N_21328);
xnor U23365 (N_23365,N_21752,N_20377);
and U23366 (N_23366,N_20205,N_21156);
xnor U23367 (N_23367,N_20413,N_20436);
nor U23368 (N_23368,N_21394,N_20074);
nand U23369 (N_23369,N_21308,N_21691);
nor U23370 (N_23370,N_20290,N_20847);
or U23371 (N_23371,N_21429,N_21090);
nor U23372 (N_23372,N_21922,N_21875);
nor U23373 (N_23373,N_20292,N_21961);
and U23374 (N_23374,N_20781,N_20240);
and U23375 (N_23375,N_21093,N_21179);
or U23376 (N_23376,N_20419,N_21287);
nand U23377 (N_23377,N_20302,N_21012);
and U23378 (N_23378,N_20861,N_20343);
and U23379 (N_23379,N_20977,N_21437);
and U23380 (N_23380,N_21189,N_20109);
and U23381 (N_23381,N_20798,N_20870);
or U23382 (N_23382,N_21851,N_21954);
and U23383 (N_23383,N_21531,N_21323);
nor U23384 (N_23384,N_21708,N_20821);
nand U23385 (N_23385,N_21623,N_20298);
xnor U23386 (N_23386,N_21696,N_20955);
nand U23387 (N_23387,N_21932,N_20044);
nand U23388 (N_23388,N_21208,N_20414);
nor U23389 (N_23389,N_20615,N_21646);
or U23390 (N_23390,N_20519,N_21763);
xnor U23391 (N_23391,N_20434,N_21760);
and U23392 (N_23392,N_21172,N_21868);
nor U23393 (N_23393,N_21809,N_21655);
xnor U23394 (N_23394,N_21050,N_21313);
xor U23395 (N_23395,N_20061,N_21482);
nand U23396 (N_23396,N_21365,N_20840);
xor U23397 (N_23397,N_20186,N_20874);
nand U23398 (N_23398,N_20854,N_21460);
nor U23399 (N_23399,N_21551,N_20555);
nand U23400 (N_23400,N_20773,N_20432);
nand U23401 (N_23401,N_20844,N_21484);
or U23402 (N_23402,N_20746,N_20908);
or U23403 (N_23403,N_21941,N_21293);
nand U23404 (N_23404,N_21676,N_20870);
xnor U23405 (N_23405,N_20858,N_20656);
nand U23406 (N_23406,N_21219,N_20119);
or U23407 (N_23407,N_21175,N_21986);
nor U23408 (N_23408,N_20083,N_21779);
xnor U23409 (N_23409,N_21161,N_20078);
or U23410 (N_23410,N_20403,N_20459);
and U23411 (N_23411,N_20783,N_21471);
and U23412 (N_23412,N_20542,N_21506);
xor U23413 (N_23413,N_20433,N_21254);
nand U23414 (N_23414,N_21684,N_21426);
and U23415 (N_23415,N_21634,N_21305);
nand U23416 (N_23416,N_20206,N_20974);
and U23417 (N_23417,N_20164,N_20498);
and U23418 (N_23418,N_20675,N_21950);
or U23419 (N_23419,N_20814,N_21427);
and U23420 (N_23420,N_20443,N_20877);
xnor U23421 (N_23421,N_20494,N_21905);
or U23422 (N_23422,N_21115,N_21918);
nand U23423 (N_23423,N_21861,N_20030);
and U23424 (N_23424,N_21538,N_20588);
or U23425 (N_23425,N_20184,N_21088);
nand U23426 (N_23426,N_20412,N_20205);
nor U23427 (N_23427,N_20957,N_21749);
nor U23428 (N_23428,N_21751,N_21091);
and U23429 (N_23429,N_21216,N_20603);
or U23430 (N_23430,N_21625,N_21132);
nand U23431 (N_23431,N_21047,N_21740);
xor U23432 (N_23432,N_20174,N_21515);
nor U23433 (N_23433,N_20616,N_21024);
xor U23434 (N_23434,N_20826,N_20658);
nor U23435 (N_23435,N_20245,N_20239);
nand U23436 (N_23436,N_20751,N_20308);
xnor U23437 (N_23437,N_20047,N_21572);
or U23438 (N_23438,N_20114,N_21099);
or U23439 (N_23439,N_21668,N_21726);
xnor U23440 (N_23440,N_21331,N_21426);
nand U23441 (N_23441,N_21590,N_20155);
nand U23442 (N_23442,N_21950,N_20602);
xnor U23443 (N_23443,N_21453,N_20607);
nand U23444 (N_23444,N_20031,N_20071);
nor U23445 (N_23445,N_20087,N_20622);
or U23446 (N_23446,N_21357,N_21625);
and U23447 (N_23447,N_20678,N_21662);
nand U23448 (N_23448,N_20644,N_20788);
or U23449 (N_23449,N_21020,N_20745);
nor U23450 (N_23450,N_21723,N_21115);
and U23451 (N_23451,N_20056,N_20404);
nand U23452 (N_23452,N_21275,N_21886);
nand U23453 (N_23453,N_20047,N_21224);
or U23454 (N_23454,N_21746,N_20196);
xor U23455 (N_23455,N_21643,N_21181);
nor U23456 (N_23456,N_20521,N_21869);
xor U23457 (N_23457,N_20670,N_20410);
xnor U23458 (N_23458,N_20008,N_21085);
nor U23459 (N_23459,N_20728,N_21999);
xor U23460 (N_23460,N_21424,N_21905);
nor U23461 (N_23461,N_20902,N_21245);
xnor U23462 (N_23462,N_21687,N_20666);
and U23463 (N_23463,N_21314,N_20046);
or U23464 (N_23464,N_20644,N_21513);
nand U23465 (N_23465,N_21756,N_20300);
nor U23466 (N_23466,N_20835,N_21968);
xor U23467 (N_23467,N_20184,N_21247);
nand U23468 (N_23468,N_20978,N_21878);
and U23469 (N_23469,N_21075,N_20041);
and U23470 (N_23470,N_21951,N_20957);
nand U23471 (N_23471,N_21500,N_21961);
nor U23472 (N_23472,N_21318,N_21798);
or U23473 (N_23473,N_21677,N_20934);
xnor U23474 (N_23474,N_21049,N_20398);
nor U23475 (N_23475,N_20226,N_21031);
and U23476 (N_23476,N_20381,N_21419);
and U23477 (N_23477,N_20812,N_20342);
or U23478 (N_23478,N_21982,N_21598);
and U23479 (N_23479,N_20060,N_21740);
nor U23480 (N_23480,N_21647,N_21810);
xnor U23481 (N_23481,N_20671,N_21367);
or U23482 (N_23482,N_20685,N_21263);
nor U23483 (N_23483,N_21708,N_20833);
nor U23484 (N_23484,N_20537,N_21176);
or U23485 (N_23485,N_21916,N_20299);
nand U23486 (N_23486,N_20711,N_21171);
nand U23487 (N_23487,N_21642,N_20221);
nor U23488 (N_23488,N_21055,N_21144);
or U23489 (N_23489,N_20237,N_20693);
and U23490 (N_23490,N_21468,N_21189);
xor U23491 (N_23491,N_20901,N_20918);
or U23492 (N_23492,N_20965,N_20145);
nor U23493 (N_23493,N_20560,N_20643);
or U23494 (N_23494,N_21362,N_21314);
and U23495 (N_23495,N_20077,N_20274);
nand U23496 (N_23496,N_20084,N_20883);
nor U23497 (N_23497,N_20661,N_20779);
or U23498 (N_23498,N_21067,N_21594);
nand U23499 (N_23499,N_21755,N_21770);
nor U23500 (N_23500,N_21976,N_21984);
nand U23501 (N_23501,N_20442,N_21782);
nor U23502 (N_23502,N_20338,N_20604);
nor U23503 (N_23503,N_20244,N_21323);
nor U23504 (N_23504,N_20897,N_20525);
nand U23505 (N_23505,N_20787,N_21859);
and U23506 (N_23506,N_21514,N_20949);
nand U23507 (N_23507,N_21045,N_20616);
nand U23508 (N_23508,N_21379,N_21186);
xnor U23509 (N_23509,N_21461,N_21377);
nand U23510 (N_23510,N_20419,N_20440);
and U23511 (N_23511,N_21033,N_20750);
xor U23512 (N_23512,N_21821,N_20259);
or U23513 (N_23513,N_20054,N_20601);
or U23514 (N_23514,N_21039,N_21571);
and U23515 (N_23515,N_21529,N_20189);
xor U23516 (N_23516,N_20046,N_21748);
nand U23517 (N_23517,N_20130,N_21569);
nor U23518 (N_23518,N_21665,N_21715);
and U23519 (N_23519,N_20395,N_20557);
nor U23520 (N_23520,N_21624,N_21763);
and U23521 (N_23521,N_21438,N_20472);
nor U23522 (N_23522,N_20378,N_21659);
and U23523 (N_23523,N_21143,N_21520);
and U23524 (N_23524,N_20098,N_21855);
nand U23525 (N_23525,N_21439,N_20973);
or U23526 (N_23526,N_21112,N_20255);
xor U23527 (N_23527,N_21668,N_20377);
and U23528 (N_23528,N_20420,N_21031);
and U23529 (N_23529,N_21114,N_20271);
nor U23530 (N_23530,N_20657,N_20093);
nand U23531 (N_23531,N_20378,N_21485);
xor U23532 (N_23532,N_21173,N_20093);
nor U23533 (N_23533,N_21901,N_20146);
and U23534 (N_23534,N_21030,N_20996);
xor U23535 (N_23535,N_20935,N_21244);
and U23536 (N_23536,N_21029,N_21832);
nand U23537 (N_23537,N_21337,N_21829);
and U23538 (N_23538,N_20343,N_20139);
nor U23539 (N_23539,N_21492,N_20862);
or U23540 (N_23540,N_20954,N_21204);
and U23541 (N_23541,N_20501,N_20735);
nand U23542 (N_23542,N_20073,N_20922);
and U23543 (N_23543,N_21198,N_21657);
nor U23544 (N_23544,N_21159,N_20163);
xnor U23545 (N_23545,N_20258,N_20275);
nor U23546 (N_23546,N_20213,N_20614);
or U23547 (N_23547,N_21471,N_20474);
xnor U23548 (N_23548,N_20844,N_21059);
xor U23549 (N_23549,N_21242,N_20678);
or U23550 (N_23550,N_20395,N_21578);
nor U23551 (N_23551,N_21730,N_21914);
xnor U23552 (N_23552,N_21691,N_20250);
xor U23553 (N_23553,N_20278,N_21808);
nor U23554 (N_23554,N_20545,N_20448);
nor U23555 (N_23555,N_21077,N_20726);
and U23556 (N_23556,N_21026,N_20794);
nor U23557 (N_23557,N_21357,N_21103);
nand U23558 (N_23558,N_21516,N_20863);
nand U23559 (N_23559,N_21779,N_20531);
xor U23560 (N_23560,N_21454,N_21101);
xnor U23561 (N_23561,N_20204,N_20932);
xor U23562 (N_23562,N_21136,N_20098);
xnor U23563 (N_23563,N_21607,N_20514);
nand U23564 (N_23564,N_20392,N_21138);
or U23565 (N_23565,N_21165,N_20461);
and U23566 (N_23566,N_20589,N_21553);
and U23567 (N_23567,N_21237,N_20582);
nand U23568 (N_23568,N_21463,N_20797);
and U23569 (N_23569,N_20144,N_21723);
nor U23570 (N_23570,N_20750,N_20549);
xnor U23571 (N_23571,N_20645,N_21635);
or U23572 (N_23572,N_21195,N_21608);
nand U23573 (N_23573,N_20342,N_20709);
and U23574 (N_23574,N_20988,N_21447);
xor U23575 (N_23575,N_20620,N_21613);
and U23576 (N_23576,N_21452,N_20697);
and U23577 (N_23577,N_21975,N_21210);
xnor U23578 (N_23578,N_21221,N_21346);
and U23579 (N_23579,N_21006,N_20596);
nand U23580 (N_23580,N_20438,N_21393);
xnor U23581 (N_23581,N_21750,N_21261);
nand U23582 (N_23582,N_21986,N_21594);
nand U23583 (N_23583,N_20964,N_20160);
nor U23584 (N_23584,N_20877,N_21179);
nor U23585 (N_23585,N_20875,N_20559);
nor U23586 (N_23586,N_21492,N_20543);
nand U23587 (N_23587,N_20578,N_20615);
xnor U23588 (N_23588,N_20772,N_21110);
or U23589 (N_23589,N_20448,N_21440);
xnor U23590 (N_23590,N_20364,N_20303);
nand U23591 (N_23591,N_21562,N_21443);
or U23592 (N_23592,N_21453,N_21835);
or U23593 (N_23593,N_20486,N_20096);
nand U23594 (N_23594,N_20792,N_21009);
xnor U23595 (N_23595,N_21825,N_21338);
and U23596 (N_23596,N_20952,N_21836);
nand U23597 (N_23597,N_21324,N_21954);
and U23598 (N_23598,N_20189,N_20379);
or U23599 (N_23599,N_20975,N_20419);
and U23600 (N_23600,N_21051,N_20337);
xnor U23601 (N_23601,N_20031,N_21936);
and U23602 (N_23602,N_20559,N_20743);
xnor U23603 (N_23603,N_20697,N_21311);
or U23604 (N_23604,N_20431,N_21054);
and U23605 (N_23605,N_21354,N_21801);
xor U23606 (N_23606,N_20134,N_20694);
or U23607 (N_23607,N_20059,N_21868);
nand U23608 (N_23608,N_20495,N_21526);
nor U23609 (N_23609,N_21125,N_20192);
or U23610 (N_23610,N_21660,N_20821);
or U23611 (N_23611,N_21226,N_21912);
xnor U23612 (N_23612,N_20262,N_21950);
and U23613 (N_23613,N_20482,N_21393);
or U23614 (N_23614,N_20700,N_21757);
nand U23615 (N_23615,N_20824,N_21811);
nand U23616 (N_23616,N_20479,N_20657);
or U23617 (N_23617,N_21239,N_20951);
xor U23618 (N_23618,N_20489,N_21765);
nor U23619 (N_23619,N_20353,N_20831);
and U23620 (N_23620,N_20056,N_20519);
xor U23621 (N_23621,N_20445,N_20056);
nor U23622 (N_23622,N_21940,N_20730);
nand U23623 (N_23623,N_20432,N_20060);
or U23624 (N_23624,N_21562,N_20708);
or U23625 (N_23625,N_21555,N_21077);
nor U23626 (N_23626,N_21813,N_20907);
nor U23627 (N_23627,N_21063,N_21412);
nor U23628 (N_23628,N_20453,N_20508);
nor U23629 (N_23629,N_20351,N_20667);
xnor U23630 (N_23630,N_20892,N_21723);
and U23631 (N_23631,N_21761,N_21127);
nand U23632 (N_23632,N_21438,N_21399);
and U23633 (N_23633,N_20774,N_20638);
nor U23634 (N_23634,N_21974,N_20411);
nand U23635 (N_23635,N_20982,N_21844);
and U23636 (N_23636,N_21398,N_21285);
and U23637 (N_23637,N_20226,N_20868);
nor U23638 (N_23638,N_21405,N_20512);
xor U23639 (N_23639,N_21701,N_21214);
xnor U23640 (N_23640,N_21243,N_21876);
nor U23641 (N_23641,N_21695,N_20835);
xnor U23642 (N_23642,N_21612,N_21824);
nand U23643 (N_23643,N_21480,N_20908);
or U23644 (N_23644,N_21803,N_21605);
or U23645 (N_23645,N_21894,N_21236);
nor U23646 (N_23646,N_20562,N_20778);
nor U23647 (N_23647,N_21001,N_21060);
nor U23648 (N_23648,N_20555,N_21708);
nand U23649 (N_23649,N_20397,N_21828);
or U23650 (N_23650,N_20504,N_20203);
xnor U23651 (N_23651,N_21786,N_21501);
or U23652 (N_23652,N_20821,N_21229);
nand U23653 (N_23653,N_21811,N_20929);
xnor U23654 (N_23654,N_20329,N_21231);
xnor U23655 (N_23655,N_20544,N_20131);
xnor U23656 (N_23656,N_21031,N_20016);
xor U23657 (N_23657,N_21152,N_20836);
and U23658 (N_23658,N_20696,N_21312);
nand U23659 (N_23659,N_21813,N_20062);
and U23660 (N_23660,N_20818,N_20017);
and U23661 (N_23661,N_21068,N_20842);
or U23662 (N_23662,N_21437,N_20823);
nand U23663 (N_23663,N_21527,N_21372);
nand U23664 (N_23664,N_20679,N_20774);
and U23665 (N_23665,N_21275,N_21131);
and U23666 (N_23666,N_20724,N_21908);
xnor U23667 (N_23667,N_20694,N_20544);
nor U23668 (N_23668,N_21906,N_21696);
and U23669 (N_23669,N_20264,N_20592);
xor U23670 (N_23670,N_21831,N_21326);
and U23671 (N_23671,N_21667,N_21665);
nor U23672 (N_23672,N_20552,N_20785);
nor U23673 (N_23673,N_20596,N_21915);
and U23674 (N_23674,N_21179,N_20231);
or U23675 (N_23675,N_21801,N_20634);
xor U23676 (N_23676,N_21245,N_20792);
and U23677 (N_23677,N_20722,N_20891);
and U23678 (N_23678,N_21460,N_20911);
nor U23679 (N_23679,N_21780,N_21817);
and U23680 (N_23680,N_20189,N_20670);
nor U23681 (N_23681,N_20644,N_21807);
or U23682 (N_23682,N_20712,N_20177);
nand U23683 (N_23683,N_21983,N_21893);
or U23684 (N_23684,N_20598,N_20822);
or U23685 (N_23685,N_20837,N_20763);
nand U23686 (N_23686,N_21708,N_21275);
xnor U23687 (N_23687,N_20255,N_21303);
nand U23688 (N_23688,N_20774,N_20512);
xor U23689 (N_23689,N_20945,N_21854);
nand U23690 (N_23690,N_21479,N_20456);
nand U23691 (N_23691,N_20758,N_21228);
nand U23692 (N_23692,N_20202,N_20995);
xor U23693 (N_23693,N_20013,N_21130);
nor U23694 (N_23694,N_21378,N_20203);
nor U23695 (N_23695,N_21935,N_20802);
xor U23696 (N_23696,N_21653,N_21037);
xor U23697 (N_23697,N_21185,N_21186);
xor U23698 (N_23698,N_21649,N_21329);
nand U23699 (N_23699,N_20304,N_20599);
nor U23700 (N_23700,N_20323,N_20800);
or U23701 (N_23701,N_20590,N_20051);
nand U23702 (N_23702,N_21265,N_20640);
xnor U23703 (N_23703,N_21772,N_20615);
nand U23704 (N_23704,N_21321,N_20257);
and U23705 (N_23705,N_21790,N_20702);
or U23706 (N_23706,N_20289,N_20247);
nor U23707 (N_23707,N_20519,N_21357);
nand U23708 (N_23708,N_20925,N_20684);
nand U23709 (N_23709,N_20637,N_21235);
nand U23710 (N_23710,N_21977,N_21589);
and U23711 (N_23711,N_21545,N_21095);
xnor U23712 (N_23712,N_21057,N_21865);
and U23713 (N_23713,N_21206,N_20573);
xnor U23714 (N_23714,N_20084,N_21014);
or U23715 (N_23715,N_21971,N_21119);
nand U23716 (N_23716,N_20969,N_21497);
or U23717 (N_23717,N_20855,N_20397);
xor U23718 (N_23718,N_20127,N_20839);
and U23719 (N_23719,N_20612,N_20684);
nand U23720 (N_23720,N_20363,N_21762);
and U23721 (N_23721,N_20109,N_20159);
or U23722 (N_23722,N_20277,N_21113);
or U23723 (N_23723,N_20334,N_21390);
xor U23724 (N_23724,N_21782,N_21797);
or U23725 (N_23725,N_20476,N_21092);
xor U23726 (N_23726,N_20376,N_20452);
nand U23727 (N_23727,N_21565,N_20740);
nor U23728 (N_23728,N_21934,N_20755);
and U23729 (N_23729,N_21114,N_20488);
and U23730 (N_23730,N_20005,N_21334);
or U23731 (N_23731,N_21889,N_20474);
xnor U23732 (N_23732,N_20945,N_21724);
xor U23733 (N_23733,N_21706,N_20807);
and U23734 (N_23734,N_21443,N_21190);
nor U23735 (N_23735,N_21012,N_21016);
and U23736 (N_23736,N_20051,N_20006);
or U23737 (N_23737,N_20164,N_20769);
nand U23738 (N_23738,N_21187,N_20175);
nand U23739 (N_23739,N_21294,N_20749);
nor U23740 (N_23740,N_21770,N_20298);
nand U23741 (N_23741,N_20900,N_20806);
nand U23742 (N_23742,N_20222,N_21397);
nor U23743 (N_23743,N_20409,N_21174);
xnor U23744 (N_23744,N_21168,N_21603);
or U23745 (N_23745,N_20265,N_20362);
and U23746 (N_23746,N_21296,N_21278);
or U23747 (N_23747,N_20768,N_21474);
or U23748 (N_23748,N_21834,N_21548);
nor U23749 (N_23749,N_20763,N_21334);
or U23750 (N_23750,N_21126,N_20848);
and U23751 (N_23751,N_21011,N_21576);
and U23752 (N_23752,N_21165,N_21491);
xnor U23753 (N_23753,N_20262,N_20761);
nand U23754 (N_23754,N_20238,N_20828);
nand U23755 (N_23755,N_21498,N_21074);
nand U23756 (N_23756,N_20354,N_20204);
xnor U23757 (N_23757,N_21952,N_21203);
nand U23758 (N_23758,N_20317,N_20390);
and U23759 (N_23759,N_20362,N_21231);
nor U23760 (N_23760,N_21673,N_21943);
and U23761 (N_23761,N_20261,N_21161);
nor U23762 (N_23762,N_21391,N_21823);
and U23763 (N_23763,N_20229,N_20714);
nand U23764 (N_23764,N_21138,N_21096);
or U23765 (N_23765,N_20226,N_20686);
nand U23766 (N_23766,N_20446,N_21553);
nor U23767 (N_23767,N_21489,N_20036);
xnor U23768 (N_23768,N_20612,N_21819);
or U23769 (N_23769,N_21181,N_21912);
nor U23770 (N_23770,N_21496,N_21794);
nor U23771 (N_23771,N_21853,N_21002);
and U23772 (N_23772,N_20922,N_20148);
nand U23773 (N_23773,N_20104,N_20043);
xnor U23774 (N_23774,N_20852,N_20689);
nor U23775 (N_23775,N_20496,N_20453);
nor U23776 (N_23776,N_21461,N_20118);
and U23777 (N_23777,N_20934,N_21629);
nor U23778 (N_23778,N_21882,N_21307);
xor U23779 (N_23779,N_21412,N_20036);
and U23780 (N_23780,N_20968,N_21364);
and U23781 (N_23781,N_20980,N_21351);
or U23782 (N_23782,N_20792,N_20571);
xnor U23783 (N_23783,N_21015,N_20704);
and U23784 (N_23784,N_21029,N_20210);
nor U23785 (N_23785,N_20863,N_21127);
and U23786 (N_23786,N_21909,N_20341);
or U23787 (N_23787,N_21931,N_20265);
nor U23788 (N_23788,N_20170,N_21853);
or U23789 (N_23789,N_20712,N_20096);
xor U23790 (N_23790,N_21492,N_20957);
or U23791 (N_23791,N_21073,N_20398);
nand U23792 (N_23792,N_20271,N_20982);
and U23793 (N_23793,N_21855,N_20054);
nand U23794 (N_23794,N_21738,N_20665);
nor U23795 (N_23795,N_20890,N_21532);
xor U23796 (N_23796,N_21935,N_20798);
xor U23797 (N_23797,N_21397,N_20474);
or U23798 (N_23798,N_20045,N_21638);
nor U23799 (N_23799,N_20952,N_21323);
and U23800 (N_23800,N_21607,N_21369);
nor U23801 (N_23801,N_21811,N_21212);
nand U23802 (N_23802,N_20579,N_20654);
and U23803 (N_23803,N_20576,N_20282);
nor U23804 (N_23804,N_21182,N_21745);
xor U23805 (N_23805,N_21985,N_20855);
nor U23806 (N_23806,N_21477,N_20170);
nand U23807 (N_23807,N_20184,N_20871);
nor U23808 (N_23808,N_20583,N_20445);
or U23809 (N_23809,N_20333,N_21853);
or U23810 (N_23810,N_20510,N_21812);
or U23811 (N_23811,N_20261,N_21861);
and U23812 (N_23812,N_20391,N_21889);
nand U23813 (N_23813,N_20112,N_20024);
xnor U23814 (N_23814,N_21333,N_21371);
nand U23815 (N_23815,N_21355,N_21212);
nand U23816 (N_23816,N_21560,N_20413);
xor U23817 (N_23817,N_20641,N_21018);
or U23818 (N_23818,N_20526,N_21402);
xor U23819 (N_23819,N_20637,N_20174);
nor U23820 (N_23820,N_20224,N_21864);
and U23821 (N_23821,N_20426,N_21423);
xor U23822 (N_23822,N_21653,N_20288);
or U23823 (N_23823,N_21205,N_20303);
xor U23824 (N_23824,N_20959,N_20142);
nand U23825 (N_23825,N_21205,N_20734);
or U23826 (N_23826,N_20030,N_20098);
nand U23827 (N_23827,N_21969,N_21066);
xor U23828 (N_23828,N_21401,N_21489);
and U23829 (N_23829,N_20919,N_20942);
or U23830 (N_23830,N_21358,N_20727);
nor U23831 (N_23831,N_20085,N_21640);
and U23832 (N_23832,N_21233,N_21733);
nand U23833 (N_23833,N_20291,N_20730);
or U23834 (N_23834,N_21347,N_21003);
xnor U23835 (N_23835,N_21597,N_20071);
nor U23836 (N_23836,N_21470,N_21953);
or U23837 (N_23837,N_21493,N_20145);
xnor U23838 (N_23838,N_20975,N_20833);
and U23839 (N_23839,N_20782,N_20944);
nor U23840 (N_23840,N_21804,N_21534);
or U23841 (N_23841,N_21847,N_21537);
and U23842 (N_23842,N_20476,N_21078);
nor U23843 (N_23843,N_20721,N_20009);
and U23844 (N_23844,N_20558,N_20834);
or U23845 (N_23845,N_20598,N_20635);
nand U23846 (N_23846,N_20986,N_20989);
nand U23847 (N_23847,N_21457,N_20802);
nor U23848 (N_23848,N_21878,N_21776);
nand U23849 (N_23849,N_21184,N_20922);
or U23850 (N_23850,N_20647,N_21418);
and U23851 (N_23851,N_21494,N_20331);
or U23852 (N_23852,N_21878,N_21994);
xnor U23853 (N_23853,N_20733,N_20687);
xnor U23854 (N_23854,N_20577,N_20886);
or U23855 (N_23855,N_21411,N_20852);
nor U23856 (N_23856,N_21391,N_21724);
or U23857 (N_23857,N_20693,N_20099);
xor U23858 (N_23858,N_20664,N_20180);
or U23859 (N_23859,N_21437,N_20169);
nor U23860 (N_23860,N_20240,N_20569);
nor U23861 (N_23861,N_21243,N_21294);
nand U23862 (N_23862,N_20697,N_21301);
xor U23863 (N_23863,N_21224,N_20740);
or U23864 (N_23864,N_20349,N_20408);
and U23865 (N_23865,N_20837,N_21925);
xnor U23866 (N_23866,N_21880,N_21271);
or U23867 (N_23867,N_21083,N_21829);
and U23868 (N_23868,N_20243,N_20818);
nor U23869 (N_23869,N_21443,N_20954);
xnor U23870 (N_23870,N_21888,N_20025);
nor U23871 (N_23871,N_20410,N_20336);
nand U23872 (N_23872,N_21701,N_20582);
nand U23873 (N_23873,N_20304,N_20571);
or U23874 (N_23874,N_21805,N_21773);
nand U23875 (N_23875,N_20387,N_21844);
and U23876 (N_23876,N_21486,N_20251);
nand U23877 (N_23877,N_21231,N_20208);
xnor U23878 (N_23878,N_21169,N_20346);
and U23879 (N_23879,N_21038,N_20828);
and U23880 (N_23880,N_20289,N_21191);
xor U23881 (N_23881,N_21594,N_21357);
xnor U23882 (N_23882,N_21743,N_20471);
and U23883 (N_23883,N_20841,N_20201);
or U23884 (N_23884,N_20748,N_21961);
xnor U23885 (N_23885,N_21243,N_20581);
nand U23886 (N_23886,N_20744,N_21436);
nor U23887 (N_23887,N_20879,N_21378);
and U23888 (N_23888,N_20103,N_20438);
nor U23889 (N_23889,N_21719,N_20322);
and U23890 (N_23890,N_21585,N_20516);
nand U23891 (N_23891,N_21146,N_21198);
nor U23892 (N_23892,N_20143,N_20200);
and U23893 (N_23893,N_20365,N_20095);
and U23894 (N_23894,N_21152,N_21620);
or U23895 (N_23895,N_21151,N_20931);
xor U23896 (N_23896,N_21906,N_20325);
or U23897 (N_23897,N_21957,N_21873);
and U23898 (N_23898,N_20960,N_21648);
xor U23899 (N_23899,N_21497,N_21236);
or U23900 (N_23900,N_21735,N_21178);
and U23901 (N_23901,N_20787,N_21592);
nand U23902 (N_23902,N_21057,N_21619);
xor U23903 (N_23903,N_21877,N_20521);
nand U23904 (N_23904,N_21337,N_21862);
xnor U23905 (N_23905,N_21260,N_20390);
xor U23906 (N_23906,N_20151,N_20650);
nand U23907 (N_23907,N_20352,N_20535);
or U23908 (N_23908,N_20329,N_20574);
nor U23909 (N_23909,N_21419,N_20992);
xnor U23910 (N_23910,N_20563,N_20891);
and U23911 (N_23911,N_21076,N_21329);
and U23912 (N_23912,N_21755,N_21370);
nor U23913 (N_23913,N_21719,N_21564);
or U23914 (N_23914,N_21908,N_20815);
nand U23915 (N_23915,N_20822,N_20964);
nor U23916 (N_23916,N_20160,N_21066);
and U23917 (N_23917,N_20261,N_21846);
nor U23918 (N_23918,N_20593,N_20868);
nand U23919 (N_23919,N_21750,N_21764);
and U23920 (N_23920,N_20832,N_21109);
and U23921 (N_23921,N_21542,N_20802);
or U23922 (N_23922,N_21370,N_20190);
nand U23923 (N_23923,N_21429,N_20625);
nor U23924 (N_23924,N_20651,N_20361);
xnor U23925 (N_23925,N_20968,N_20314);
and U23926 (N_23926,N_21555,N_20439);
or U23927 (N_23927,N_20161,N_21024);
xnor U23928 (N_23928,N_21203,N_21110);
xnor U23929 (N_23929,N_21653,N_20086);
nand U23930 (N_23930,N_20547,N_20817);
or U23931 (N_23931,N_21309,N_20282);
or U23932 (N_23932,N_21060,N_20655);
nand U23933 (N_23933,N_20140,N_21408);
or U23934 (N_23934,N_21973,N_20412);
nor U23935 (N_23935,N_21307,N_21752);
or U23936 (N_23936,N_20466,N_21220);
nor U23937 (N_23937,N_21505,N_21676);
xor U23938 (N_23938,N_20562,N_20757);
or U23939 (N_23939,N_21190,N_21196);
or U23940 (N_23940,N_21167,N_20810);
nor U23941 (N_23941,N_20726,N_21660);
nor U23942 (N_23942,N_20069,N_21911);
nor U23943 (N_23943,N_21876,N_20995);
nand U23944 (N_23944,N_21920,N_20873);
xor U23945 (N_23945,N_21952,N_20727);
nor U23946 (N_23946,N_20946,N_21995);
or U23947 (N_23947,N_21837,N_21370);
xnor U23948 (N_23948,N_20123,N_21629);
and U23949 (N_23949,N_20828,N_21297);
or U23950 (N_23950,N_20002,N_20586);
nand U23951 (N_23951,N_21465,N_21952);
nand U23952 (N_23952,N_21767,N_21289);
nand U23953 (N_23953,N_20496,N_21507);
nor U23954 (N_23954,N_21355,N_20102);
nor U23955 (N_23955,N_20639,N_21004);
and U23956 (N_23956,N_21214,N_20143);
nor U23957 (N_23957,N_21704,N_21469);
nand U23958 (N_23958,N_21478,N_20167);
nor U23959 (N_23959,N_20904,N_21283);
nand U23960 (N_23960,N_20228,N_20849);
nor U23961 (N_23961,N_20036,N_20335);
or U23962 (N_23962,N_20432,N_21436);
nand U23963 (N_23963,N_20601,N_20669);
and U23964 (N_23964,N_21631,N_20447);
xnor U23965 (N_23965,N_20822,N_20052);
and U23966 (N_23966,N_20861,N_21838);
or U23967 (N_23967,N_21507,N_20121);
and U23968 (N_23968,N_21677,N_21213);
and U23969 (N_23969,N_20442,N_20534);
or U23970 (N_23970,N_21193,N_20604);
xnor U23971 (N_23971,N_20791,N_21423);
nor U23972 (N_23972,N_20118,N_21860);
or U23973 (N_23973,N_21424,N_20576);
nand U23974 (N_23974,N_20535,N_20948);
or U23975 (N_23975,N_20570,N_21379);
or U23976 (N_23976,N_20174,N_21222);
nor U23977 (N_23977,N_21702,N_20954);
nor U23978 (N_23978,N_21070,N_21536);
nor U23979 (N_23979,N_21293,N_20007);
and U23980 (N_23980,N_20795,N_21384);
nand U23981 (N_23981,N_20667,N_20452);
or U23982 (N_23982,N_20205,N_21678);
nor U23983 (N_23983,N_21849,N_21667);
or U23984 (N_23984,N_21342,N_21280);
or U23985 (N_23985,N_21245,N_20145);
nor U23986 (N_23986,N_20525,N_21888);
nor U23987 (N_23987,N_21507,N_21986);
or U23988 (N_23988,N_21196,N_21667);
xnor U23989 (N_23989,N_21144,N_21275);
nor U23990 (N_23990,N_21411,N_21136);
or U23991 (N_23991,N_21728,N_20330);
and U23992 (N_23992,N_20633,N_21925);
or U23993 (N_23993,N_21097,N_20512);
xnor U23994 (N_23994,N_20552,N_20898);
nand U23995 (N_23995,N_20077,N_21435);
and U23996 (N_23996,N_21972,N_21334);
nand U23997 (N_23997,N_20379,N_20838);
nand U23998 (N_23998,N_20607,N_20269);
or U23999 (N_23999,N_20827,N_20707);
or U24000 (N_24000,N_23508,N_23947);
xor U24001 (N_24001,N_23825,N_23635);
xnor U24002 (N_24002,N_22451,N_22523);
nand U24003 (N_24003,N_22093,N_22872);
nor U24004 (N_24004,N_22146,N_23402);
nand U24005 (N_24005,N_23221,N_23095);
xor U24006 (N_24006,N_22740,N_23180);
and U24007 (N_24007,N_23854,N_23621);
and U24008 (N_24008,N_23866,N_23557);
xor U24009 (N_24009,N_23566,N_23423);
nor U24010 (N_24010,N_23116,N_22348);
nor U24011 (N_24011,N_23534,N_22486);
and U24012 (N_24012,N_22737,N_22324);
xor U24013 (N_24013,N_23269,N_22404);
and U24014 (N_24014,N_23043,N_23084);
and U24015 (N_24015,N_23175,N_23259);
or U24016 (N_24016,N_22558,N_22668);
nand U24017 (N_24017,N_22898,N_22521);
nor U24018 (N_24018,N_22956,N_23222);
xnor U24019 (N_24019,N_22206,N_22647);
xor U24020 (N_24020,N_22722,N_22595);
nor U24021 (N_24021,N_22813,N_23634);
or U24022 (N_24022,N_23442,N_23161);
xnor U24023 (N_24023,N_23928,N_23348);
or U24024 (N_24024,N_22625,N_23837);
nor U24025 (N_24025,N_23802,N_22336);
nor U24026 (N_24026,N_23716,N_23686);
nand U24027 (N_24027,N_23698,N_22251);
nand U24028 (N_24028,N_23968,N_22752);
xnor U24029 (N_24029,N_22084,N_23005);
nor U24030 (N_24030,N_23248,N_23464);
xor U24031 (N_24031,N_23579,N_22860);
or U24032 (N_24032,N_23395,N_23963);
or U24033 (N_24033,N_22703,N_23048);
nand U24034 (N_24034,N_23450,N_22353);
nor U24035 (N_24035,N_23561,N_23559);
nor U24036 (N_24036,N_22712,N_22401);
nor U24037 (N_24037,N_23551,N_23233);
and U24038 (N_24038,N_23598,N_23030);
or U24039 (N_24039,N_23040,N_22108);
and U24040 (N_24040,N_22914,N_22731);
and U24041 (N_24041,N_22407,N_23230);
nor U24042 (N_24042,N_22545,N_23618);
xor U24043 (N_24043,N_23893,N_22017);
xnor U24044 (N_24044,N_22091,N_22476);
or U24045 (N_24045,N_23009,N_22276);
nand U24046 (N_24046,N_23115,N_22958);
nor U24047 (N_24047,N_23125,N_23096);
or U24048 (N_24048,N_22425,N_22998);
xor U24049 (N_24049,N_23637,N_22380);
and U24050 (N_24050,N_23504,N_23465);
nand U24051 (N_24051,N_23266,N_23571);
xnor U24052 (N_24052,N_22779,N_23822);
nand U24053 (N_24053,N_22411,N_22540);
nand U24054 (N_24054,N_23904,N_22579);
and U24055 (N_24055,N_22855,N_22924);
nor U24056 (N_24056,N_23517,N_22697);
nand U24057 (N_24057,N_22052,N_23282);
xnor U24058 (N_24058,N_22531,N_23304);
or U24059 (N_24059,N_22641,N_23328);
nor U24060 (N_24060,N_22562,N_23372);
or U24061 (N_24061,N_23117,N_22143);
nand U24062 (N_24062,N_23946,N_23432);
nand U24063 (N_24063,N_22297,N_23017);
and U24064 (N_24064,N_23341,N_23952);
nor U24065 (N_24065,N_22717,N_22213);
or U24066 (N_24066,N_22462,N_22196);
or U24067 (N_24067,N_22505,N_23872);
nand U24068 (N_24068,N_23717,N_23001);
nand U24069 (N_24069,N_22663,N_22071);
and U24070 (N_24070,N_22002,N_23056);
nor U24071 (N_24071,N_23940,N_22575);
nor U24072 (N_24072,N_22508,N_23624);
and U24073 (N_24073,N_22314,N_22217);
xor U24074 (N_24074,N_23424,N_22601);
nor U24075 (N_24075,N_22271,N_23629);
or U24076 (N_24076,N_23858,N_23882);
or U24077 (N_24077,N_22605,N_23871);
nand U24078 (N_24078,N_22238,N_22820);
xnor U24079 (N_24079,N_22205,N_23315);
and U24080 (N_24080,N_22804,N_22742);
and U24081 (N_24081,N_22946,N_23536);
xor U24082 (N_24082,N_22332,N_23948);
nand U24083 (N_24083,N_22285,N_22194);
nor U24084 (N_24084,N_23285,N_23604);
or U24085 (N_24085,N_22098,N_22927);
or U24086 (N_24086,N_22392,N_22319);
and U24087 (N_24087,N_22948,N_22607);
xor U24088 (N_24088,N_23167,N_23581);
or U24089 (N_24089,N_23857,N_23232);
nand U24090 (N_24090,N_23473,N_23436);
nor U24091 (N_24091,N_23687,N_23061);
xor U24092 (N_24092,N_22773,N_23648);
nand U24093 (N_24093,N_22784,N_23414);
xnor U24094 (N_24094,N_22096,N_23879);
nor U24095 (N_24095,N_23234,N_22802);
and U24096 (N_24096,N_23038,N_22879);
nand U24097 (N_24097,N_23933,N_22999);
or U24098 (N_24098,N_23205,N_23470);
nor U24099 (N_24099,N_23358,N_23950);
and U24100 (N_24100,N_22799,N_23141);
nand U24101 (N_24101,N_22550,N_22408);
nand U24102 (N_24102,N_23626,N_22049);
or U24103 (N_24103,N_23092,N_23885);
nand U24104 (N_24104,N_22051,N_22788);
or U24105 (N_24105,N_23615,N_22274);
or U24106 (N_24106,N_23365,N_23861);
nor U24107 (N_24107,N_22874,N_23573);
nand U24108 (N_24108,N_22995,N_22387);
or U24109 (N_24109,N_22710,N_22258);
and U24110 (N_24110,N_23251,N_23331);
nor U24111 (N_24111,N_23601,N_23123);
and U24112 (N_24112,N_23216,N_22756);
nor U24113 (N_24113,N_22242,N_22282);
xnor U24114 (N_24114,N_23699,N_22959);
xor U24115 (N_24115,N_23146,N_23409);
or U24116 (N_24116,N_22437,N_22526);
nor U24117 (N_24117,N_22553,N_23823);
and U24118 (N_24118,N_22092,N_22787);
nor U24119 (N_24119,N_22878,N_23462);
nand U24120 (N_24120,N_22480,N_23741);
and U24121 (N_24121,N_22546,N_23463);
xor U24122 (N_24122,N_22800,N_23862);
or U24123 (N_24123,N_23889,N_22608);
nor U24124 (N_24124,N_22653,N_22357);
nand U24125 (N_24125,N_22805,N_22844);
nor U24126 (N_24126,N_23630,N_22597);
nand U24127 (N_24127,N_22381,N_23769);
or U24128 (N_24128,N_22181,N_22384);
xor U24129 (N_24129,N_23090,N_22635);
nor U24130 (N_24130,N_22750,N_22603);
or U24131 (N_24131,N_22340,N_22485);
and U24132 (N_24132,N_23712,N_22645);
or U24133 (N_24133,N_22247,N_23770);
or U24134 (N_24134,N_22309,N_22280);
xor U24135 (N_24135,N_22024,N_23976);
and U24136 (N_24136,N_23931,N_22130);
nand U24137 (N_24137,N_22629,N_23327);
or U24138 (N_24138,N_23909,N_23758);
nor U24139 (N_24139,N_22970,N_22846);
xor U24140 (N_24140,N_23786,N_23826);
nand U24141 (N_24141,N_23787,N_23429);
xnor U24142 (N_24142,N_22424,N_23632);
nor U24143 (N_24143,N_23468,N_23294);
xnor U24144 (N_24144,N_22266,N_23800);
nor U24145 (N_24145,N_22236,N_23939);
nor U24146 (N_24146,N_23135,N_22237);
or U24147 (N_24147,N_23736,N_23188);
nor U24148 (N_24148,N_23670,N_22836);
or U24149 (N_24149,N_22957,N_22871);
nor U24150 (N_24150,N_22079,N_22207);
or U24151 (N_24151,N_23509,N_22382);
or U24152 (N_24152,N_22661,N_23359);
nand U24153 (N_24153,N_23367,N_23132);
and U24154 (N_24154,N_23268,N_22839);
and U24155 (N_24155,N_22479,N_23446);
nand U24156 (N_24156,N_23776,N_22287);
or U24157 (N_24157,N_22515,N_23431);
nand U24158 (N_24158,N_23695,N_23452);
and U24159 (N_24159,N_22222,N_22517);
nor U24160 (N_24160,N_22857,N_23318);
xnor U24161 (N_24161,N_22250,N_22907);
xnor U24162 (N_24162,N_22027,N_22151);
nor U24163 (N_24163,N_22159,N_23671);
xnor U24164 (N_24164,N_22911,N_23720);
nor U24165 (N_24165,N_23015,N_23320);
nor U24166 (N_24166,N_23605,N_22869);
nand U24167 (N_24167,N_23788,N_23426);
or U24168 (N_24168,N_22818,N_23196);
xor U24169 (N_24169,N_23214,N_23789);
xnor U24170 (N_24170,N_22997,N_23192);
nand U24171 (N_24171,N_22056,N_23869);
nand U24172 (N_24172,N_22125,N_22041);
xnor U24173 (N_24173,N_23599,N_23591);
nand U24174 (N_24174,N_22322,N_23984);
nand U24175 (N_24175,N_22106,N_23708);
nor U24176 (N_24176,N_22708,N_22815);
nor U24177 (N_24177,N_22606,N_22650);
xor U24178 (N_24178,N_23026,N_22524);
and U24179 (N_24179,N_22239,N_23875);
xor U24180 (N_24180,N_23403,N_22436);
or U24181 (N_24181,N_23245,N_23199);
or U24182 (N_24182,N_22721,N_23541);
and U24183 (N_24183,N_23730,N_23021);
and U24184 (N_24184,N_22054,N_22442);
and U24185 (N_24185,N_22269,N_23845);
and U24186 (N_24186,N_23992,N_23790);
nand U24187 (N_24187,N_23820,N_22256);
nor U24188 (N_24188,N_22067,N_22578);
and U24189 (N_24189,N_22665,N_23377);
and U24190 (N_24190,N_23673,N_23903);
xnor U24191 (N_24191,N_23891,N_23779);
nor U24192 (N_24192,N_23439,N_23526);
nand U24193 (N_24193,N_22918,N_23032);
nor U24194 (N_24194,N_23956,N_22583);
xnor U24195 (N_24195,N_22267,N_23018);
nor U24196 (N_24196,N_22749,N_23515);
nor U24197 (N_24197,N_22050,N_23053);
and U24198 (N_24198,N_22011,N_23636);
and U24199 (N_24199,N_22539,N_23128);
or U24200 (N_24200,N_23916,N_23025);
and U24201 (N_24201,N_23838,N_22028);
nand U24202 (N_24202,N_22964,N_23937);
or U24203 (N_24203,N_22377,N_22230);
and U24204 (N_24204,N_22718,N_22134);
and U24205 (N_24205,N_23198,N_22853);
nand U24206 (N_24206,N_23548,N_23554);
nor U24207 (N_24207,N_23189,N_22952);
nor U24208 (N_24208,N_23070,N_23485);
nand U24209 (N_24209,N_23839,N_22528);
and U24210 (N_24210,N_23537,N_22154);
or U24211 (N_24211,N_22156,N_23610);
or U24212 (N_24212,N_23574,N_23643);
or U24213 (N_24213,N_23801,N_23731);
or U24214 (N_24214,N_23994,N_22249);
nor U24215 (N_24215,N_23997,N_22840);
and U24216 (N_24216,N_23420,N_22277);
xnor U24217 (N_24217,N_22358,N_22789);
or U24218 (N_24218,N_23512,N_23475);
or U24219 (N_24219,N_22337,N_23979);
nand U24220 (N_24220,N_22488,N_23973);
xnor U24221 (N_24221,N_23142,N_23533);
and U24222 (N_24222,N_22817,N_22592);
and U24223 (N_24223,N_23772,N_23104);
and U24224 (N_24224,N_23980,N_22669);
nand U24225 (N_24225,N_23576,N_23796);
and U24226 (N_24226,N_23710,N_22199);
or U24227 (N_24227,N_22430,N_22930);
or U24228 (N_24228,N_23706,N_22568);
nand U24229 (N_24229,N_22925,N_23531);
xor U24230 (N_24230,N_23612,N_22178);
xor U24231 (N_24231,N_22630,N_22754);
nor U24232 (N_24232,N_23258,N_23703);
nor U24233 (N_24233,N_22715,N_23210);
or U24234 (N_24234,N_23276,N_23363);
nand U24235 (N_24235,N_23682,N_23572);
xor U24236 (N_24236,N_23927,N_22417);
or U24237 (N_24237,N_23926,N_22573);
xor U24238 (N_24238,N_22803,N_22983);
and U24239 (N_24239,N_23521,N_22620);
xor U24240 (N_24240,N_22262,N_23352);
or U24241 (N_24241,N_23166,N_23316);
nand U24242 (N_24242,N_22720,N_22498);
or U24243 (N_24243,N_22499,N_23919);
nor U24244 (N_24244,N_23003,N_23784);
nor U24245 (N_24245,N_22455,N_22363);
nor U24246 (N_24246,N_22910,N_23203);
and U24247 (N_24247,N_22219,N_23074);
nand U24248 (N_24248,N_22509,N_23549);
and U24249 (N_24249,N_22748,N_22954);
or U24250 (N_24250,N_22281,N_23811);
and U24251 (N_24251,N_22210,N_23191);
and U24252 (N_24252,N_22456,N_23150);
nor U24253 (N_24253,N_22117,N_22667);
xnor U24254 (N_24254,N_23317,N_22723);
nor U24255 (N_24255,N_23588,N_23303);
or U24256 (N_24256,N_23727,N_22006);
and U24257 (N_24257,N_22938,N_23944);
xnor U24258 (N_24258,N_23649,N_23081);
xnor U24259 (N_24259,N_23865,N_23479);
or U24260 (N_24260,N_23564,N_22637);
xnor U24261 (N_24261,N_22313,N_23676);
and U24262 (N_24262,N_23754,N_23490);
or U24263 (N_24263,N_22713,N_22689);
xor U24264 (N_24264,N_22652,N_23842);
xor U24265 (N_24265,N_22776,N_23181);
nor U24266 (N_24266,N_22899,N_22126);
nand U24267 (N_24267,N_23783,N_22687);
nor U24268 (N_24268,N_23019,N_22851);
and U24269 (N_24269,N_22989,N_23121);
or U24270 (N_24270,N_22015,N_23740);
nand U24271 (N_24271,N_23087,N_23575);
or U24272 (N_24272,N_22868,N_22293);
nand U24273 (N_24273,N_23982,N_22588);
nand U24274 (N_24274,N_22478,N_22691);
or U24275 (N_24275,N_23350,N_22842);
nor U24276 (N_24276,N_23611,N_22881);
or U24277 (N_24277,N_23340,N_23281);
and U24278 (N_24278,N_23287,N_22681);
xor U24279 (N_24279,N_22591,N_23308);
nand U24280 (N_24280,N_22057,N_22174);
nand U24281 (N_24281,N_23035,N_22039);
or U24282 (N_24282,N_22438,N_22140);
xnor U24283 (N_24283,N_23714,N_22321);
xnor U24284 (N_24284,N_23284,N_22435);
and U24285 (N_24285,N_23413,N_23388);
or U24286 (N_24286,N_22235,N_22987);
nand U24287 (N_24287,N_23407,N_22876);
nor U24288 (N_24288,N_22116,N_22968);
nor U24289 (N_24289,N_23065,N_22504);
or U24290 (N_24290,N_23457,N_22596);
nor U24291 (N_24291,N_23739,N_23428);
nand U24292 (N_24292,N_22428,N_22613);
and U24293 (N_24293,N_22413,N_22530);
nand U24294 (N_24294,N_22229,N_23664);
xnor U24295 (N_24295,N_22942,N_23400);
xnor U24296 (N_24296,N_22201,N_23466);
or U24297 (N_24297,N_22825,N_22894);
and U24298 (N_24298,N_22111,N_22137);
or U24299 (N_24299,N_23832,N_22204);
or U24300 (N_24300,N_23532,N_22360);
or U24301 (N_24301,N_22311,N_23160);
xor U24302 (N_24302,N_23288,N_22295);
and U24303 (N_24303,N_22094,N_23323);
nand U24304 (N_24304,N_23384,N_23438);
and U24305 (N_24305,N_22974,N_22753);
nand U24306 (N_24306,N_23808,N_22099);
nor U24307 (N_24307,N_23502,N_22105);
and U24308 (N_24308,N_23067,N_22906);
nor U24309 (N_24309,N_23041,N_22757);
or U24310 (N_24310,N_22810,N_22030);
xnor U24311 (N_24311,N_22383,N_23332);
nand U24312 (N_24312,N_23989,N_22169);
nor U24313 (N_24313,N_22537,N_22474);
or U24314 (N_24314,N_23828,N_22215);
nand U24315 (N_24315,N_23349,N_22985);
and U24316 (N_24316,N_23397,N_22160);
nand U24317 (N_24317,N_22439,N_23505);
nand U24318 (N_24318,N_22762,N_22496);
or U24319 (N_24319,N_23277,N_23672);
or U24320 (N_24320,N_22795,N_23737);
nor U24321 (N_24321,N_23237,N_23492);
or U24322 (N_24322,N_23645,N_22122);
xnor U24323 (N_24323,N_23763,N_23362);
and U24324 (N_24324,N_22316,N_22263);
and U24325 (N_24325,N_22355,N_22070);
nor U24326 (N_24326,N_23228,N_22443);
xor U24327 (N_24327,N_22714,N_23692);
and U24328 (N_24328,N_22088,N_22136);
or U24329 (N_24329,N_23254,N_23729);
or U24330 (N_24330,N_23638,N_22761);
xnor U24331 (N_24331,N_22612,N_22555);
xor U24332 (N_24332,N_23155,N_22211);
and U24333 (N_24333,N_23625,N_23456);
and U24334 (N_24334,N_23392,N_22100);
and U24335 (N_24335,N_23212,N_23333);
xnor U24336 (N_24336,N_23380,N_23435);
nor U24337 (N_24337,N_22388,N_22253);
xor U24338 (N_24338,N_22915,N_23088);
nor U24339 (N_24339,N_23631,N_23242);
or U24340 (N_24340,N_23220,N_22935);
or U24341 (N_24341,N_22241,N_23079);
or U24342 (N_24342,N_23778,N_23208);
nand U24343 (N_24343,N_22228,N_22566);
or U24344 (N_24344,N_22415,N_22586);
xnor U24345 (N_24345,N_23910,N_22170);
nor U24346 (N_24346,N_23724,N_22829);
xnor U24347 (N_24347,N_23745,N_23360);
nand U24348 (N_24348,N_22976,N_22529);
nand U24349 (N_24349,N_23013,N_23239);
and U24350 (N_24350,N_22705,N_23295);
or U24351 (N_24351,N_23831,N_23934);
nand U24352 (N_24352,N_22240,N_22768);
xor U24353 (N_24353,N_23097,N_22138);
and U24354 (N_24354,N_23883,N_22335);
nor U24355 (N_24355,N_22943,N_23908);
nand U24356 (N_24356,N_22621,N_22278);
nand U24357 (N_24357,N_22986,N_23217);
nor U24358 (N_24358,N_23182,N_23346);
nor U24359 (N_24359,N_22859,N_22038);
nand U24360 (N_24360,N_22863,N_22640);
or U24361 (N_24361,N_23105,N_22197);
nand U24362 (N_24362,N_23306,N_23183);
xor U24363 (N_24363,N_23039,N_22157);
nor U24364 (N_24364,N_22864,N_23033);
or U24365 (N_24365,N_22089,N_23998);
and U24366 (N_24366,N_23766,N_22007);
and U24367 (N_24367,N_23179,N_23905);
and U24368 (N_24368,N_22127,N_22895);
or U24369 (N_24369,N_23393,N_22385);
and U24370 (N_24370,N_23119,N_22484);
xnor U24371 (N_24371,N_23412,N_22245);
nand U24372 (N_24372,N_22808,N_23586);
and U24373 (N_24373,N_23036,N_22203);
or U24374 (N_24374,N_22464,N_22090);
nand U24375 (N_24375,N_22048,N_23775);
xnor U24376 (N_24376,N_23522,N_22678);
xnor U24377 (N_24377,N_23723,N_22374);
nand U24378 (N_24378,N_23733,N_23165);
xnor U24379 (N_24379,N_22359,N_22511);
xor U24380 (N_24380,N_23153,N_22043);
nand U24381 (N_24381,N_23404,N_22153);
or U24382 (N_24382,N_23029,N_23725);
and U24383 (N_24383,N_22312,N_23034);
and U24384 (N_24384,N_22945,N_22164);
xor U24385 (N_24385,N_23793,N_22135);
nand U24386 (N_24386,N_22701,N_22725);
and U24387 (N_24387,N_23964,N_23007);
nor U24388 (N_24388,N_22457,N_22128);
nor U24389 (N_24389,N_22738,N_23164);
or U24390 (N_24390,N_22195,N_23978);
xnor U24391 (N_24391,N_23197,N_22448);
and U24392 (N_24392,N_22124,N_22900);
xnor U24393 (N_24393,N_22171,N_23028);
or U24394 (N_24394,N_22260,N_22264);
and U24395 (N_24395,N_23818,N_23925);
or U24396 (N_24396,N_22921,N_23113);
xnor U24397 (N_24397,N_22719,N_23840);
or U24398 (N_24398,N_22421,N_23836);
xnor U24399 (N_24399,N_22631,N_23523);
xor U24400 (N_24400,N_23897,N_23051);
nor U24401 (N_24401,N_23678,N_23109);
nand U24402 (N_24402,N_22660,N_23681);
nor U24403 (N_24403,N_22520,N_22040);
or U24404 (N_24404,N_23675,N_23370);
nand U24405 (N_24405,N_22065,N_23609);
and U24406 (N_24406,N_23941,N_22232);
nand U24407 (N_24407,N_22074,N_22554);
xnor U24408 (N_24408,N_23083,N_22165);
nand U24409 (N_24409,N_23815,N_22931);
and U24410 (N_24410,N_22590,N_23550);
nand U24411 (N_24411,N_22783,N_22150);
nor U24412 (N_24412,N_23791,N_22345);
and U24413 (N_24413,N_23623,N_22390);
nor U24414 (N_24414,N_22533,N_22822);
nor U24415 (N_24415,N_22699,N_22809);
xnor U24416 (N_24416,N_22996,N_22941);
and U24417 (N_24417,N_22163,N_23487);
nand U24418 (N_24418,N_23353,N_22473);
nand U24419 (N_24419,N_22780,N_23050);
nor U24420 (N_24420,N_22564,N_22744);
xnor U24421 (N_24421,N_22110,N_23231);
xnor U24422 (N_24422,N_23726,N_23507);
xnor U24423 (N_24423,N_23218,N_22962);
nand U24424 (N_24424,N_23915,N_23158);
xor U24425 (N_24425,N_23660,N_23722);
nor U24426 (N_24426,N_23345,N_22702);
and U24427 (N_24427,N_22330,N_22979);
and U24428 (N_24428,N_22598,N_22600);
nor U24429 (N_24429,N_22624,N_22080);
or U24430 (N_24430,N_22131,N_23339);
and U24431 (N_24431,N_22212,N_22676);
or U24432 (N_24432,N_22402,N_22323);
or U24433 (N_24433,N_22535,N_23954);
xnor U24434 (N_24434,N_23480,N_22189);
nor U24435 (N_24435,N_23577,N_23369);
and U24436 (N_24436,N_23765,N_22097);
xor U24437 (N_24437,N_23555,N_23062);
and U24438 (N_24438,N_23274,N_23387);
nand U24439 (N_24439,N_23149,N_23416);
and U24440 (N_24440,N_22187,N_23540);
nand U24441 (N_24441,N_23782,N_22183);
nor U24442 (N_24442,N_23140,N_22409);
xor U24443 (N_24443,N_22977,N_22549);
xor U24444 (N_24444,N_23356,N_22463);
xor U24445 (N_24445,N_22349,N_23064);
or U24446 (N_24446,N_22231,N_23873);
and U24447 (N_24447,N_22303,N_22690);
xnor U24448 (N_24448,N_22410,N_22685);
and U24449 (N_24449,N_23024,N_22939);
and U24450 (N_24450,N_22279,N_22045);
nand U24451 (N_24451,N_23443,N_22830);
and U24452 (N_24452,N_23411,N_23949);
or U24453 (N_24453,N_23816,N_22350);
or U24454 (N_24454,N_23371,N_23874);
and U24455 (N_24455,N_22082,N_23073);
and U24456 (N_24456,N_22730,N_23995);
or U24457 (N_24457,N_22465,N_22733);
and U24458 (N_24458,N_23653,N_23817);
xor U24459 (N_24459,N_22534,N_23658);
xnor U24460 (N_24460,N_22774,N_22066);
nand U24461 (N_24461,N_22862,N_23488);
or U24462 (N_24462,N_23361,N_22837);
and U24463 (N_24463,N_22882,N_22142);
xor U24464 (N_24464,N_22577,N_22400);
and U24465 (N_24465,N_22364,N_22492);
nor U24466 (N_24466,N_23215,N_23595);
nand U24467 (N_24467,N_22014,N_23415);
or U24468 (N_24468,N_23528,N_23746);
or U24469 (N_24469,N_22420,N_23898);
xor U24470 (N_24470,N_23107,N_23434);
and U24471 (N_24471,N_22695,N_23513);
xor U24472 (N_24472,N_23589,N_23603);
nor U24473 (N_24473,N_22192,N_22732);
and U24474 (N_24474,N_23810,N_23880);
and U24475 (N_24475,N_23923,N_22929);
nand U24476 (N_24476,N_23441,N_23760);
xnor U24477 (N_24477,N_23538,N_23476);
xor U24478 (N_24478,N_23619,N_22467);
xor U24479 (N_24479,N_23535,N_22866);
and U24480 (N_24480,N_23843,N_23847);
xnor U24481 (N_24481,N_23265,N_23511);
nor U24482 (N_24482,N_23799,N_23560);
nor U24483 (N_24483,N_22755,N_23342);
nor U24484 (N_24484,N_23558,N_22729);
or U24485 (N_24485,N_23986,N_22471);
and U24486 (N_24486,N_23386,N_22901);
nor U24487 (N_24487,N_23319,N_23211);
nor U24488 (N_24488,N_23827,N_23145);
xnor U24489 (N_24489,N_23855,N_22763);
or U24490 (N_24490,N_23958,N_22046);
xor U24491 (N_24491,N_23546,N_22460);
or U24492 (N_24492,N_22843,N_22643);
nor U24493 (N_24493,N_22767,N_22461);
xor U24494 (N_24494,N_22396,N_23493);
xor U24495 (N_24495,N_22967,N_22759);
and U24496 (N_24496,N_23974,N_22419);
nand U24497 (N_24497,N_22162,N_22516);
nand U24498 (N_24498,N_23674,N_23641);
nand U24499 (N_24499,N_22481,N_23633);
nand U24500 (N_24500,N_23685,N_23756);
xnor U24501 (N_24501,N_22746,N_23884);
xor U24502 (N_24502,N_23309,N_23835);
nand U24503 (N_24503,N_23750,N_22398);
nor U24504 (N_24504,N_22922,N_23644);
and U24505 (N_24505,N_22917,N_23850);
nor U24506 (N_24506,N_23103,N_23795);
and U24507 (N_24507,N_22031,N_22771);
and U24508 (N_24508,N_23713,N_23144);
xnor U24509 (N_24509,N_22184,N_23814);
nor U24510 (N_24510,N_22944,N_22684);
nand U24511 (N_24511,N_22431,N_22812);
or U24512 (N_24512,N_22543,N_22819);
and U24513 (N_24513,N_23467,N_23565);
xnor U24514 (N_24514,N_23496,N_23008);
nor U24515 (N_24515,N_23556,N_23170);
nor U24516 (N_24516,N_22781,N_23172);
or U24517 (N_24517,N_23497,N_22429);
nor U24518 (N_24518,N_23094,N_23616);
xor U24519 (N_24519,N_23448,N_23562);
nand U24520 (N_24520,N_23798,N_22622);
or U24521 (N_24521,N_22955,N_22261);
xnor U24522 (N_24522,N_23298,N_22365);
xnor U24523 (N_24523,N_22167,N_22386);
or U24524 (N_24524,N_22626,N_23803);
and U24525 (N_24525,N_22102,N_23344);
or U24526 (N_24526,N_23100,N_22892);
xnor U24527 (N_24527,N_23410,N_23852);
nand U24528 (N_24528,N_23955,N_23190);
nor U24529 (N_24529,N_23668,N_23914);
and U24530 (N_24530,N_23136,N_23206);
xnor U24531 (N_24531,N_22833,N_23876);
or U24532 (N_24532,N_22908,N_22452);
or U24533 (N_24533,N_23390,N_22877);
and U24534 (N_24534,N_23291,N_22772);
xor U24535 (N_24535,N_23525,N_23499);
nor U24536 (N_24536,N_23768,N_23099);
nor U24537 (N_24537,N_22887,N_22841);
or U24538 (N_24538,N_23449,N_22994);
xor U24539 (N_24539,N_22422,N_23398);
xnor U24540 (N_24540,N_23299,N_23972);
nor U24541 (N_24541,N_23283,N_22512);
xnor U24542 (N_24542,N_22447,N_22797);
nor U24543 (N_24543,N_22475,N_22491);
or U24544 (N_24544,N_23510,N_23280);
or U24545 (N_24545,N_22727,N_22379);
nand U24546 (N_24546,N_22778,N_23759);
nand U24547 (N_24547,N_23489,N_23743);
and U24548 (N_24548,N_22328,N_23622);
and U24549 (N_24549,N_22785,N_22490);
and U24550 (N_24550,N_22814,N_23454);
and U24551 (N_24551,N_23702,N_23357);
nor U24552 (N_24552,N_22766,N_23697);
or U24553 (N_24553,N_23744,N_23004);
and U24554 (N_24554,N_23124,N_23707);
xor U24555 (N_24555,N_23651,N_23620);
nand U24556 (N_24556,N_22406,N_23921);
xor U24557 (N_24557,N_22777,N_22694);
xor U24558 (N_24558,N_22570,N_23614);
nand U24559 (N_24559,N_23981,N_22806);
and U24560 (N_24560,N_23133,N_23023);
or U24561 (N_24561,N_23901,N_22270);
and U24562 (N_24562,N_23406,N_23469);
nand U24563 (N_24563,N_23262,N_22551);
and U24564 (N_24564,N_23628,N_23011);
or U24565 (N_24565,N_22304,N_23241);
and U24566 (N_24566,N_23223,N_23461);
nand U24567 (N_24567,N_22120,N_23657);
and U24568 (N_24568,N_23684,N_22648);
nor U24569 (N_24569,N_23042,N_22299);
xor U24570 (N_24570,N_22704,N_23325);
xnor U24571 (N_24571,N_23310,N_23755);
and U24572 (N_24572,N_23286,N_23993);
or U24573 (N_24573,N_22642,N_23545);
and U24574 (N_24574,N_23547,N_22152);
nor U24575 (N_24575,N_23924,N_23157);
or U24576 (N_24576,N_22794,N_22688);
nor U24577 (N_24577,N_22831,N_22707);
xor U24578 (N_24578,N_23516,N_22619);
nand U24579 (N_24579,N_23263,N_22114);
and U24580 (N_24580,N_23728,N_23243);
and U24581 (N_24581,N_23389,N_23296);
and U24582 (N_24582,N_22107,N_23260);
nand U24583 (N_24583,N_23225,N_22611);
nand U24584 (N_24584,N_23596,N_23031);
and U24585 (N_24585,N_22832,N_23202);
and U24586 (N_24586,N_22651,N_23126);
xor U24587 (N_24587,N_23227,N_22556);
nor U24588 (N_24588,N_23137,N_23383);
or U24589 (N_24589,N_22234,N_22101);
and U24590 (N_24590,N_23364,N_23878);
or U24591 (N_24591,N_23679,N_23396);
nand U24592 (N_24592,N_23690,N_23195);
xor U24593 (N_24593,N_23762,N_22272);
or U24594 (N_24594,N_23892,N_23552);
nand U24595 (N_24595,N_23143,N_22670);
nand U24596 (N_24596,N_23700,N_22993);
nor U24597 (N_24597,N_22224,N_23127);
and U24598 (N_24598,N_23580,N_23747);
nor U24599 (N_24599,N_22376,N_23060);
or U24600 (N_24600,N_22765,N_22459);
or U24601 (N_24601,N_22072,N_22283);
nand U24602 (N_24602,N_23683,N_22141);
and U24603 (N_24603,N_23322,N_23147);
and U24604 (N_24604,N_22905,N_23646);
or U24605 (N_24605,N_22064,N_23689);
nor U24606 (N_24606,N_22019,N_23527);
and U24607 (N_24607,N_23985,N_22284);
or U24608 (N_24608,N_23235,N_23886);
nand U24609 (N_24609,N_22320,N_23066);
or U24610 (N_24610,N_23076,N_23951);
nor U24611 (N_24611,N_22155,N_22850);
and U24612 (N_24612,N_23696,N_22086);
nor U24613 (N_24613,N_22728,N_22338);
nor U24614 (N_24614,N_22115,N_23661);
or U24615 (N_24615,N_23055,N_22483);
xor U24616 (N_24616,N_22268,N_22903);
nor U24617 (N_24617,N_23022,N_22623);
or U24618 (N_24618,N_23273,N_22497);
and U24619 (N_24619,N_23337,N_23351);
and U24620 (N_24620,N_23821,N_22811);
and U24621 (N_24621,N_23486,N_22683);
or U24622 (N_24622,N_22741,N_23264);
xor U24623 (N_24623,N_22933,N_23355);
xor U24624 (N_24624,N_23935,N_23809);
or U24625 (N_24625,N_22414,N_23394);
and U24626 (N_24626,N_22300,N_22920);
nor U24627 (N_24627,N_22209,N_23639);
and U24628 (N_24628,N_22173,N_23932);
nor U24629 (N_24629,N_22724,N_22037);
nor U24630 (N_24630,N_22033,N_23627);
nand U24631 (N_24631,N_22133,N_22518);
and U24632 (N_24632,N_23279,N_22012);
and U24633 (N_24633,N_22658,N_23544);
nand U24634 (N_24634,N_22453,N_22633);
nor U24635 (N_24635,N_23715,N_22301);
xor U24636 (N_24636,N_23058,N_22609);
or U24637 (N_24637,N_23000,N_22602);
nor U24638 (N_24638,N_23292,N_22023);
nor U24639 (N_24639,N_23860,N_22190);
nor U24640 (N_24640,N_22904,N_22427);
xnor U24641 (N_24641,N_22791,N_23806);
and U24642 (N_24642,N_22121,N_22351);
nand U24643 (N_24643,N_22580,N_22032);
and U24644 (N_24644,N_23797,N_23379);
nand U24645 (N_24645,N_23688,N_23666);
xor U24646 (N_24646,N_22928,N_23961);
or U24647 (N_24647,N_23072,N_23311);
nor U24648 (N_24648,N_23709,N_22674);
xnor U24649 (N_24649,N_22886,N_22405);
xnor U24650 (N_24650,N_22888,N_22760);
nor U24651 (N_24651,N_22827,N_22403);
nor U24652 (N_24652,N_22493,N_23159);
nor U24653 (N_24653,N_23694,N_22541);
and U24654 (N_24654,N_23122,N_23642);
nand U24655 (N_24655,N_23863,N_23045);
or U24656 (N_24656,N_22992,N_23999);
or U24657 (N_24657,N_23193,N_22883);
and U24658 (N_24658,N_23849,N_22616);
nor U24659 (N_24659,N_22078,N_22307);
nand U24660 (N_24660,N_22610,N_22807);
nor U24661 (N_24661,N_22161,N_22000);
or U24662 (N_24662,N_22333,N_23255);
nor U24663 (N_24663,N_22971,N_22978);
and U24664 (N_24664,N_22593,N_22144);
nand U24665 (N_24665,N_23261,N_22560);
nor U24666 (N_24666,N_22062,N_23922);
nor U24667 (N_24667,N_22824,N_22369);
nand U24668 (N_24668,N_22584,N_23059);
xnor U24669 (N_24669,N_23991,N_23888);
nand U24670 (N_24670,N_23911,N_22826);
xnor U24671 (N_24671,N_23173,N_22325);
nand U24672 (N_24672,N_23867,N_22389);
nand U24673 (N_24673,N_22440,N_22506);
nor U24674 (N_24674,N_22004,N_22835);
nor U24675 (N_24675,N_23204,N_22188);
nand U24676 (N_24676,N_23419,N_23110);
nand U24677 (N_24677,N_23738,N_23474);
nor U24678 (N_24678,N_22472,N_22739);
nand U24679 (N_24679,N_23659,N_23481);
nor U24680 (N_24680,N_22225,N_22639);
xor U24681 (N_24681,N_23098,N_23101);
nand U24682 (N_24682,N_23721,N_23347);
and U24683 (N_24683,N_23752,N_22123);
and U24684 (N_24684,N_22649,N_23408);
nor U24685 (N_24685,N_22692,N_22775);
or U24686 (N_24686,N_22845,N_22769);
nand U24687 (N_24687,N_23417,N_23494);
or U24688 (N_24688,N_22973,N_22654);
nor U24689 (N_24689,N_23049,N_23338);
nand U24690 (N_24690,N_22361,N_22449);
xor U24691 (N_24691,N_23600,N_23329);
nand U24692 (N_24692,N_22960,N_23037);
or U24693 (N_24693,N_22937,N_22706);
nand U24694 (N_24694,N_23174,N_23895);
nand U24695 (N_24695,N_23987,N_22891);
nand U24696 (N_24696,N_23229,N_23794);
xnor U24697 (N_24697,N_22902,N_23771);
nand U24698 (N_24698,N_22148,N_23929);
nand U24699 (N_24699,N_23376,N_22145);
or U24700 (N_24700,N_23014,N_22426);
nor U24701 (N_24701,N_23270,N_22003);
or U24702 (N_24702,N_23830,N_23613);
nor U24703 (N_24703,N_22318,N_22947);
nand U24704 (N_24704,N_23002,N_22139);
nand U24705 (N_24705,N_22068,N_23774);
xnor U24706 (N_24706,N_22265,N_22934);
nor U24707 (N_24707,N_23764,N_22507);
nor U24708 (N_24708,N_22790,N_22202);
xnor U24709 (N_24709,N_22112,N_23201);
xnor U24710 (N_24710,N_23082,N_23594);
nor U24711 (N_24711,N_23890,N_22200);
nor U24712 (N_24712,N_22950,N_22013);
nor U24713 (N_24713,N_23902,N_22470);
nor U24714 (N_24714,N_22468,N_23324);
xnor U24715 (N_24715,N_22604,N_22305);
nand U24716 (N_24716,N_23401,N_23334);
nor U24717 (N_24717,N_23792,N_22227);
or U24718 (N_24718,N_22378,N_22501);
or U24719 (N_24719,N_22916,N_23819);
xnor U24720 (N_24720,N_22288,N_22961);
and U24721 (N_24721,N_23271,N_22659);
and U24722 (N_24722,N_23289,N_23156);
or U24723 (N_24723,N_23881,N_23272);
nand U24724 (N_24724,N_22984,N_23607);
or U24725 (N_24725,N_23020,N_23300);
nand U24726 (N_24726,N_22662,N_22394);
and U24727 (N_24727,N_22675,N_22341);
and U24728 (N_24728,N_22975,N_23213);
nor U24729 (N_24729,N_22758,N_23877);
nand U24730 (N_24730,N_23427,N_22965);
nor U24731 (N_24731,N_23455,N_22576);
xnor U24732 (N_24732,N_23735,N_23335);
or U24733 (N_24733,N_22821,N_22949);
or U24734 (N_24734,N_23518,N_22214);
nand U24735 (N_24735,N_22828,N_22770);
and U24736 (N_24736,N_22334,N_22873);
xnor U24737 (N_24737,N_23399,N_22849);
and U24738 (N_24738,N_22890,N_23118);
or U24739 (N_24739,N_22366,N_22252);
nor U24740 (N_24740,N_23187,N_23458);
nand U24741 (N_24741,N_23938,N_22061);
or U24742 (N_24742,N_22193,N_22709);
or U24743 (N_24743,N_22798,N_22693);
and U24744 (N_24744,N_22393,N_22001);
nand U24745 (N_24745,N_22180,N_22617);
xor U24746 (N_24746,N_23965,N_22801);
xor U24747 (N_24747,N_22542,N_22119);
or U24748 (N_24748,N_22680,N_23054);
and U24749 (N_24749,N_23374,N_22344);
nor U24750 (N_24750,N_22191,N_23907);
and U24751 (N_24751,N_22454,N_22244);
and U24752 (N_24752,N_23134,N_23495);
nor U24753 (N_24753,N_22571,N_22208);
xor U24754 (N_24754,N_22147,N_23430);
or U24755 (N_24755,N_23224,N_22848);
nand U24756 (N_24756,N_23177,N_22412);
xor U24757 (N_24757,N_22035,N_23336);
or U24758 (N_24758,N_23382,N_23662);
or U24759 (N_24759,N_23027,N_22433);
nand U24760 (N_24760,N_22343,N_22919);
nand U24761 (N_24761,N_22073,N_22988);
and U24762 (N_24762,N_22372,N_22548);
or U24763 (N_24763,N_22168,N_23590);
or U24764 (N_24764,N_23373,N_22434);
or U24765 (N_24765,N_22646,N_23829);
or U24766 (N_24766,N_22221,N_22527);
nor U24767 (N_24767,N_22021,N_23046);
and U24768 (N_24768,N_22482,N_23962);
or U24769 (N_24769,N_22103,N_23864);
and U24770 (N_24770,N_22896,N_23701);
nand U24771 (N_24771,N_22615,N_22450);
xnor U24772 (N_24772,N_22025,N_23314);
and U24773 (N_24773,N_23868,N_23529);
nor U24774 (N_24774,N_23500,N_23693);
xor U24775 (N_24775,N_23563,N_23186);
and U24776 (N_24776,N_23920,N_23063);
xor U24777 (N_24777,N_23044,N_23491);
and U24778 (N_24778,N_22743,N_23734);
and U24779 (N_24779,N_23781,N_22286);
xnor U24780 (N_24780,N_22854,N_22022);
and U24781 (N_24781,N_22638,N_22682);
and U24782 (N_24782,N_23757,N_23085);
and U24783 (N_24783,N_22634,N_22216);
xor U24784 (N_24784,N_22317,N_22255);
nand U24785 (N_24785,N_22834,N_23148);
nor U24786 (N_24786,N_22246,N_22792);
and U24787 (N_24787,N_23592,N_23969);
and U24788 (N_24788,N_22514,N_22346);
nand U24789 (N_24789,N_23343,N_22736);
xnor U24790 (N_24790,N_23080,N_23749);
xnor U24791 (N_24791,N_22503,N_22290);
nand U24792 (N_24792,N_23751,N_22696);
xor U24793 (N_24793,N_22302,N_23841);
or U24794 (N_24794,N_22567,N_23078);
or U24795 (N_24795,N_23071,N_22132);
or U24796 (N_24796,N_22081,N_22599);
xnor U24797 (N_24797,N_23075,N_23278);
xor U24798 (N_24798,N_23016,N_22734);
and U24799 (N_24799,N_23899,N_23767);
xor U24800 (N_24800,N_22926,N_23246);
nand U24801 (N_24801,N_22963,N_22458);
and U24802 (N_24802,N_23483,N_23163);
or U24803 (N_24803,N_23257,N_23584);
nand U24804 (N_24804,N_23977,N_22175);
nand U24805 (N_24805,N_22327,N_23602);
xnor U24806 (N_24806,N_22852,N_23501);
nor U24807 (N_24807,N_23139,N_23129);
or U24808 (N_24808,N_23677,N_22513);
and U24809 (N_24809,N_23851,N_22352);
nor U24810 (N_24810,N_23418,N_23375);
nand U24811 (N_24811,N_22129,N_22018);
or U24812 (N_24812,N_22373,N_22525);
nor U24813 (N_24813,N_23975,N_23942);
nor U24814 (N_24814,N_22275,N_23543);
nand U24815 (N_24815,N_22880,N_22306);
or U24816 (N_24816,N_22700,N_22273);
and U24817 (N_24817,N_23477,N_22569);
xnor U24818 (N_24818,N_23996,N_23777);
or U24819 (N_24819,N_23256,N_22786);
xnor U24820 (N_24820,N_22053,N_22489);
nand U24821 (N_24821,N_23321,N_22069);
xnor U24822 (N_24822,N_23514,N_23154);
or U24823 (N_24823,N_22793,N_23447);
xnor U24824 (N_24824,N_22932,N_22044);
nor U24825 (N_24825,N_23267,N_22289);
nand U24826 (N_24826,N_23240,N_22370);
and U24827 (N_24827,N_22923,N_22870);
nor U24828 (N_24828,N_22047,N_23667);
or U24829 (N_24829,N_22655,N_22559);
or U24830 (N_24830,N_23983,N_22469);
xnor U24831 (N_24831,N_22889,N_22445);
nand U24832 (N_24832,N_23597,N_23953);
and U24833 (N_24833,N_23542,N_23293);
xnor U24834 (N_24834,N_23244,N_22747);
nor U24835 (N_24835,N_23219,N_22565);
nand U24836 (N_24836,N_22572,N_23569);
xnor U24837 (N_24837,N_22875,N_23753);
and U24838 (N_24838,N_23894,N_23275);
nand U24839 (N_24839,N_23290,N_23052);
or U24840 (N_24840,N_23805,N_23669);
nor U24841 (N_24841,N_23650,N_22254);
or U24842 (N_24842,N_23691,N_22856);
nand U24843 (N_24843,N_22673,N_23959);
nand U24844 (N_24844,N_23471,N_22444);
or U24845 (N_24845,N_22494,N_23047);
or U24846 (N_24846,N_23966,N_22294);
and U24847 (N_24847,N_23366,N_22118);
nor U24848 (N_24848,N_22315,N_22331);
or U24849 (N_24849,N_22618,N_23433);
or U24850 (N_24850,N_23853,N_23169);
or U24851 (N_24851,N_22823,N_22182);
nand U24852 (N_24852,N_22672,N_22395);
xor U24853 (N_24853,N_22418,N_22679);
nand U24854 (N_24854,N_22686,N_22502);
or U24855 (N_24855,N_23568,N_22671);
nor U24856 (N_24856,N_23010,N_23459);
xnor U24857 (N_24857,N_23106,N_23326);
and U24858 (N_24858,N_22951,N_22166);
or U24859 (N_24859,N_23704,N_23918);
or U24860 (N_24860,N_22367,N_22764);
xnor U24861 (N_24861,N_23761,N_22574);
xnor U24862 (N_24862,N_22636,N_23151);
xnor U24863 (N_24863,N_23617,N_22104);
or U24864 (N_24864,N_22716,N_22594);
or U24865 (N_24865,N_22368,N_22711);
nor U24866 (N_24866,N_23570,N_22909);
and U24867 (N_24867,N_22177,N_22186);
and U24868 (N_24868,N_23870,N_23250);
xor U24869 (N_24869,N_22627,N_23093);
and U24870 (N_24870,N_22375,N_22557);
nor U24871 (N_24871,N_23138,N_22009);
or U24872 (N_24872,N_23524,N_22522);
and U24873 (N_24873,N_22538,N_22310);
xnor U24874 (N_24874,N_22897,N_23520);
or U24875 (N_24875,N_23578,N_22446);
and U24876 (N_24876,N_23069,N_22745);
xnor U24877 (N_24877,N_22113,N_22008);
or U24878 (N_24878,N_22614,N_22953);
nor U24879 (N_24879,N_23732,N_22342);
nand U24880 (N_24880,N_22582,N_22063);
nand U24881 (N_24881,N_22176,N_22059);
nand U24882 (N_24882,N_23742,N_23453);
or U24883 (N_24883,N_22060,N_23844);
nand U24884 (N_24884,N_23444,N_23833);
xor U24885 (N_24885,N_23391,N_23553);
nor U24886 (N_24886,N_23381,N_23705);
nor U24887 (N_24887,N_23068,N_23773);
and U24888 (N_24888,N_23185,N_23503);
nor U24889 (N_24889,N_22042,N_22536);
or U24890 (N_24890,N_23785,N_23567);
nor U24891 (N_24891,N_23091,N_23654);
xor U24892 (N_24892,N_22083,N_22561);
or U24893 (N_24893,N_22257,N_23824);
nor U24894 (N_24894,N_22029,N_22326);
nand U24895 (N_24895,N_22020,N_22329);
or U24896 (N_24896,N_23655,N_23200);
xor U24897 (N_24897,N_22632,N_22371);
nand U24898 (N_24898,N_22861,N_22095);
and U24899 (N_24899,N_22149,N_22677);
nand U24900 (N_24900,N_23582,N_23719);
nor U24901 (N_24901,N_23077,N_23089);
or U24902 (N_24902,N_23451,N_22466);
and U24903 (N_24903,N_23807,N_23111);
xor U24904 (N_24904,N_22005,N_22519);
xor U24905 (N_24905,N_22397,N_22587);
or U24906 (N_24906,N_22198,N_23108);
or U24907 (N_24907,N_23957,N_22010);
or U24908 (N_24908,N_23647,N_22735);
nand U24909 (N_24909,N_23368,N_23307);
nor U24910 (N_24910,N_22223,N_23057);
nor U24911 (N_24911,N_23130,N_22885);
or U24912 (N_24912,N_23478,N_22751);
or U24913 (N_24913,N_22259,N_23120);
and U24914 (N_24914,N_22058,N_22087);
and U24915 (N_24915,N_22865,N_22980);
or U24916 (N_24916,N_23887,N_23184);
and U24917 (N_24917,N_23930,N_22179);
or U24918 (N_24918,N_23472,N_22666);
nor U24919 (N_24919,N_22016,N_22838);
nand U24920 (N_24920,N_22589,N_23171);
xor U24921 (N_24921,N_22796,N_22354);
nor U24922 (N_24922,N_23330,N_22399);
or U24923 (N_24923,N_23405,N_23945);
or U24924 (N_24924,N_22893,N_23813);
nand U24925 (N_24925,N_23606,N_22782);
and U24926 (N_24926,N_22510,N_22657);
or U24927 (N_24927,N_22969,N_22544);
xor U24928 (N_24928,N_22391,N_22991);
and U24929 (N_24929,N_23988,N_23297);
nor U24930 (N_24930,N_22726,N_22581);
and U24931 (N_24931,N_23168,N_23587);
xor U24932 (N_24932,N_23354,N_23593);
xor U24933 (N_24933,N_23253,N_23896);
nor U24934 (N_24934,N_23112,N_23301);
nor U24935 (N_24935,N_23422,N_22940);
xnor U24936 (N_24936,N_22296,N_23608);
nor U24937 (N_24937,N_23238,N_23226);
and U24938 (N_24938,N_22243,N_23834);
and U24939 (N_24939,N_23804,N_23460);
xnor U24940 (N_24940,N_22936,N_22085);
or U24941 (N_24941,N_23917,N_23665);
xor U24942 (N_24942,N_23385,N_22291);
or U24943 (N_24943,N_22477,N_22172);
or U24944 (N_24944,N_22308,N_22298);
nor U24945 (N_24945,N_22218,N_23312);
nand U24946 (N_24946,N_22628,N_23680);
or U24947 (N_24947,N_23640,N_22972);
and U24948 (N_24948,N_23152,N_23484);
and U24949 (N_24949,N_23006,N_23656);
xnor U24950 (N_24950,N_22185,N_23990);
or U24951 (N_24951,N_22220,N_22867);
or U24952 (N_24952,N_22858,N_22816);
nor U24953 (N_24953,N_22158,N_23131);
xor U24954 (N_24954,N_23176,N_23519);
nand U24955 (N_24955,N_22966,N_23102);
nand U24956 (N_24956,N_22077,N_22055);
xor U24957 (N_24957,N_22912,N_23313);
and U24958 (N_24958,N_22441,N_23967);
and U24959 (N_24959,N_22233,N_22036);
nand U24960 (N_24960,N_23530,N_23912);
nand U24961 (N_24961,N_22248,N_22109);
nand U24962 (N_24962,N_22500,N_23207);
or U24963 (N_24963,N_22362,N_22698);
nand U24964 (N_24964,N_23425,N_22075);
xor U24965 (N_24965,N_22664,N_23718);
and U24966 (N_24966,N_23913,N_23971);
xnor U24967 (N_24967,N_23378,N_23445);
or U24968 (N_24968,N_23086,N_23943);
nand U24969 (N_24969,N_23585,N_23848);
and U24970 (N_24970,N_22982,N_23900);
nor U24971 (N_24971,N_23012,N_23506);
xnor U24972 (N_24972,N_23482,N_22990);
and U24973 (N_24973,N_23970,N_22076);
and U24974 (N_24974,N_23711,N_22487);
xor U24975 (N_24975,N_23252,N_23780);
and U24976 (N_24976,N_22347,N_22432);
and U24977 (N_24977,N_23162,N_23305);
xor U24978 (N_24978,N_22563,N_23302);
and U24979 (N_24979,N_23583,N_22026);
and U24980 (N_24980,N_23856,N_22416);
or U24981 (N_24981,N_22339,N_23209);
xor U24982 (N_24982,N_22552,N_23236);
and U24983 (N_24983,N_22884,N_22423);
and U24984 (N_24984,N_22034,N_23440);
nand U24985 (N_24985,N_22356,N_23249);
and U24986 (N_24986,N_23247,N_22226);
xor U24987 (N_24987,N_22644,N_22913);
nor U24988 (N_24988,N_23437,N_23846);
nand U24989 (N_24989,N_22981,N_23652);
xor U24990 (N_24990,N_22847,N_23194);
or U24991 (N_24991,N_23498,N_23906);
nor U24992 (N_24992,N_23960,N_23812);
and U24993 (N_24993,N_23859,N_23539);
and U24994 (N_24994,N_22495,N_23936);
or U24995 (N_24995,N_23114,N_22532);
or U24996 (N_24996,N_23178,N_22585);
nand U24997 (N_24997,N_22292,N_23663);
xnor U24998 (N_24998,N_23748,N_23421);
xnor U24999 (N_24999,N_22656,N_22547);
nand U25000 (N_25000,N_22948,N_23504);
or U25001 (N_25001,N_23088,N_22522);
nand U25002 (N_25002,N_22136,N_22001);
and U25003 (N_25003,N_23410,N_23787);
nor U25004 (N_25004,N_22607,N_22551);
or U25005 (N_25005,N_22789,N_22138);
nor U25006 (N_25006,N_22464,N_22430);
xor U25007 (N_25007,N_22667,N_23339);
xnor U25008 (N_25008,N_23909,N_22055);
nor U25009 (N_25009,N_22801,N_22930);
and U25010 (N_25010,N_23141,N_23155);
nand U25011 (N_25011,N_23953,N_22369);
xor U25012 (N_25012,N_22396,N_23544);
or U25013 (N_25013,N_22011,N_22607);
xnor U25014 (N_25014,N_23577,N_22303);
and U25015 (N_25015,N_23083,N_22388);
nor U25016 (N_25016,N_22493,N_22091);
and U25017 (N_25017,N_23585,N_22696);
nand U25018 (N_25018,N_22458,N_22101);
or U25019 (N_25019,N_22029,N_23668);
xor U25020 (N_25020,N_23959,N_23411);
and U25021 (N_25021,N_23200,N_23836);
nor U25022 (N_25022,N_22118,N_22374);
and U25023 (N_25023,N_22208,N_22890);
or U25024 (N_25024,N_22078,N_22378);
xor U25025 (N_25025,N_22104,N_22648);
xor U25026 (N_25026,N_23649,N_23620);
xnor U25027 (N_25027,N_22760,N_23519);
or U25028 (N_25028,N_22914,N_22561);
nand U25029 (N_25029,N_22573,N_23386);
nand U25030 (N_25030,N_22073,N_23363);
xor U25031 (N_25031,N_23250,N_23288);
and U25032 (N_25032,N_22052,N_23919);
nand U25033 (N_25033,N_22001,N_23533);
or U25034 (N_25034,N_22325,N_23085);
xnor U25035 (N_25035,N_23808,N_22149);
nor U25036 (N_25036,N_23611,N_23032);
or U25037 (N_25037,N_23562,N_22701);
or U25038 (N_25038,N_22129,N_23358);
nand U25039 (N_25039,N_22952,N_23601);
and U25040 (N_25040,N_22493,N_22076);
and U25041 (N_25041,N_23916,N_22235);
xnor U25042 (N_25042,N_23529,N_22676);
xnor U25043 (N_25043,N_23354,N_22885);
and U25044 (N_25044,N_23909,N_22613);
nor U25045 (N_25045,N_22564,N_22349);
or U25046 (N_25046,N_22166,N_23894);
or U25047 (N_25047,N_22590,N_23259);
nor U25048 (N_25048,N_22306,N_23368);
and U25049 (N_25049,N_22684,N_22868);
xor U25050 (N_25050,N_22169,N_22320);
nand U25051 (N_25051,N_23116,N_23361);
nand U25052 (N_25052,N_23012,N_23510);
nor U25053 (N_25053,N_23837,N_23654);
and U25054 (N_25054,N_23148,N_23943);
or U25055 (N_25055,N_23843,N_23296);
or U25056 (N_25056,N_23316,N_23506);
and U25057 (N_25057,N_23085,N_23963);
or U25058 (N_25058,N_22431,N_23820);
nor U25059 (N_25059,N_23873,N_22675);
or U25060 (N_25060,N_23825,N_22810);
nand U25061 (N_25061,N_23203,N_23281);
nand U25062 (N_25062,N_23395,N_22237);
nand U25063 (N_25063,N_22423,N_23101);
xnor U25064 (N_25064,N_23712,N_22871);
nor U25065 (N_25065,N_22774,N_22043);
or U25066 (N_25066,N_23219,N_22063);
nand U25067 (N_25067,N_23390,N_22587);
nor U25068 (N_25068,N_23579,N_23922);
nand U25069 (N_25069,N_23673,N_22941);
xor U25070 (N_25070,N_22495,N_22352);
xnor U25071 (N_25071,N_22616,N_23320);
or U25072 (N_25072,N_23551,N_22775);
xnor U25073 (N_25073,N_23519,N_22981);
nor U25074 (N_25074,N_23497,N_22550);
or U25075 (N_25075,N_22685,N_23016);
or U25076 (N_25076,N_22711,N_22303);
and U25077 (N_25077,N_22729,N_23670);
nor U25078 (N_25078,N_22704,N_22806);
nand U25079 (N_25079,N_23283,N_23210);
xor U25080 (N_25080,N_22967,N_22156);
or U25081 (N_25081,N_22223,N_22185);
nor U25082 (N_25082,N_23887,N_23144);
nand U25083 (N_25083,N_23946,N_23367);
and U25084 (N_25084,N_23373,N_23866);
or U25085 (N_25085,N_23454,N_22092);
nand U25086 (N_25086,N_23800,N_22942);
or U25087 (N_25087,N_22693,N_23060);
or U25088 (N_25088,N_23222,N_22959);
nor U25089 (N_25089,N_22079,N_22178);
and U25090 (N_25090,N_23356,N_23632);
nor U25091 (N_25091,N_23872,N_23143);
or U25092 (N_25092,N_22660,N_23512);
nand U25093 (N_25093,N_23216,N_22796);
nor U25094 (N_25094,N_22233,N_22145);
xnor U25095 (N_25095,N_22111,N_23046);
nor U25096 (N_25096,N_22747,N_22174);
and U25097 (N_25097,N_23336,N_22252);
xnor U25098 (N_25098,N_22500,N_23654);
and U25099 (N_25099,N_23845,N_22417);
nand U25100 (N_25100,N_23475,N_23226);
nand U25101 (N_25101,N_23522,N_23550);
nand U25102 (N_25102,N_22336,N_23058);
and U25103 (N_25103,N_23835,N_22848);
nor U25104 (N_25104,N_23551,N_23337);
nand U25105 (N_25105,N_22264,N_22759);
nand U25106 (N_25106,N_23555,N_23117);
xor U25107 (N_25107,N_23213,N_23898);
nor U25108 (N_25108,N_23526,N_22508);
and U25109 (N_25109,N_23201,N_22393);
nor U25110 (N_25110,N_22746,N_23016);
nand U25111 (N_25111,N_22930,N_23169);
or U25112 (N_25112,N_23516,N_22158);
or U25113 (N_25113,N_23459,N_23574);
nand U25114 (N_25114,N_22614,N_23352);
nand U25115 (N_25115,N_23734,N_23727);
nand U25116 (N_25116,N_22063,N_22537);
and U25117 (N_25117,N_22271,N_22509);
or U25118 (N_25118,N_23508,N_23415);
or U25119 (N_25119,N_23506,N_23197);
and U25120 (N_25120,N_22856,N_23118);
nand U25121 (N_25121,N_22885,N_23930);
nand U25122 (N_25122,N_23231,N_22900);
nand U25123 (N_25123,N_23587,N_22706);
and U25124 (N_25124,N_22093,N_22459);
xnor U25125 (N_25125,N_22839,N_22274);
nand U25126 (N_25126,N_23752,N_23811);
xor U25127 (N_25127,N_22655,N_23345);
and U25128 (N_25128,N_23373,N_22717);
nand U25129 (N_25129,N_23446,N_22722);
xor U25130 (N_25130,N_22946,N_22553);
and U25131 (N_25131,N_22773,N_23950);
nand U25132 (N_25132,N_23808,N_22523);
or U25133 (N_25133,N_23970,N_23252);
xor U25134 (N_25134,N_22175,N_22204);
and U25135 (N_25135,N_23544,N_22769);
xnor U25136 (N_25136,N_23988,N_22498);
xnor U25137 (N_25137,N_23374,N_22528);
nand U25138 (N_25138,N_23634,N_23782);
or U25139 (N_25139,N_23551,N_22576);
nor U25140 (N_25140,N_23143,N_22352);
and U25141 (N_25141,N_23224,N_23655);
or U25142 (N_25142,N_23296,N_22862);
and U25143 (N_25143,N_23698,N_22270);
nand U25144 (N_25144,N_23988,N_22683);
nor U25145 (N_25145,N_23195,N_23897);
xor U25146 (N_25146,N_22680,N_23358);
or U25147 (N_25147,N_22340,N_23039);
nor U25148 (N_25148,N_22963,N_22626);
and U25149 (N_25149,N_22129,N_23023);
xnor U25150 (N_25150,N_22734,N_23058);
or U25151 (N_25151,N_22392,N_22691);
nor U25152 (N_25152,N_23301,N_22115);
nand U25153 (N_25153,N_23493,N_22309);
nor U25154 (N_25154,N_23068,N_22492);
nand U25155 (N_25155,N_23916,N_22372);
nand U25156 (N_25156,N_22983,N_23137);
and U25157 (N_25157,N_22820,N_23424);
and U25158 (N_25158,N_23634,N_22080);
nand U25159 (N_25159,N_23094,N_23170);
nor U25160 (N_25160,N_22132,N_23286);
and U25161 (N_25161,N_23308,N_22985);
nor U25162 (N_25162,N_23319,N_23414);
or U25163 (N_25163,N_22326,N_23061);
nand U25164 (N_25164,N_23506,N_22956);
xnor U25165 (N_25165,N_23734,N_23632);
and U25166 (N_25166,N_22182,N_22483);
and U25167 (N_25167,N_22457,N_22482);
nand U25168 (N_25168,N_23012,N_23230);
nand U25169 (N_25169,N_23782,N_22327);
nor U25170 (N_25170,N_22679,N_23367);
nand U25171 (N_25171,N_23661,N_23756);
or U25172 (N_25172,N_23844,N_23503);
or U25173 (N_25173,N_23340,N_22446);
or U25174 (N_25174,N_23571,N_23944);
nor U25175 (N_25175,N_23360,N_22904);
and U25176 (N_25176,N_23937,N_23505);
nand U25177 (N_25177,N_23725,N_22372);
nor U25178 (N_25178,N_22006,N_23324);
or U25179 (N_25179,N_23815,N_22786);
nand U25180 (N_25180,N_23207,N_22439);
and U25181 (N_25181,N_22612,N_23605);
and U25182 (N_25182,N_22796,N_22088);
nand U25183 (N_25183,N_22344,N_22747);
nor U25184 (N_25184,N_23546,N_22054);
or U25185 (N_25185,N_22302,N_23906);
or U25186 (N_25186,N_22801,N_22538);
nand U25187 (N_25187,N_23944,N_22243);
or U25188 (N_25188,N_22335,N_23479);
nor U25189 (N_25189,N_22825,N_22981);
and U25190 (N_25190,N_23136,N_23780);
and U25191 (N_25191,N_23549,N_23215);
nand U25192 (N_25192,N_22853,N_22374);
and U25193 (N_25193,N_23436,N_23211);
nor U25194 (N_25194,N_23602,N_23489);
and U25195 (N_25195,N_23095,N_23342);
or U25196 (N_25196,N_22868,N_22636);
nor U25197 (N_25197,N_22910,N_23695);
or U25198 (N_25198,N_22640,N_22112);
and U25199 (N_25199,N_22583,N_22475);
nor U25200 (N_25200,N_23374,N_22430);
xor U25201 (N_25201,N_23194,N_22297);
nand U25202 (N_25202,N_23975,N_22635);
nor U25203 (N_25203,N_23704,N_22056);
nor U25204 (N_25204,N_23524,N_22904);
xnor U25205 (N_25205,N_22197,N_23893);
xor U25206 (N_25206,N_23186,N_23301);
or U25207 (N_25207,N_22561,N_23843);
or U25208 (N_25208,N_22372,N_23075);
nor U25209 (N_25209,N_22609,N_23650);
and U25210 (N_25210,N_23199,N_22238);
or U25211 (N_25211,N_22063,N_22958);
or U25212 (N_25212,N_22900,N_23822);
nor U25213 (N_25213,N_22451,N_22110);
and U25214 (N_25214,N_22399,N_22532);
or U25215 (N_25215,N_22665,N_22530);
and U25216 (N_25216,N_23705,N_22542);
or U25217 (N_25217,N_23948,N_23408);
or U25218 (N_25218,N_23942,N_22933);
and U25219 (N_25219,N_22521,N_22489);
and U25220 (N_25220,N_22272,N_22431);
xnor U25221 (N_25221,N_22195,N_22458);
or U25222 (N_25222,N_22701,N_22843);
nor U25223 (N_25223,N_23985,N_23017);
nand U25224 (N_25224,N_22765,N_23294);
nor U25225 (N_25225,N_23032,N_23715);
nand U25226 (N_25226,N_22136,N_22226);
nor U25227 (N_25227,N_22176,N_23269);
xnor U25228 (N_25228,N_22283,N_22292);
nor U25229 (N_25229,N_22586,N_23343);
and U25230 (N_25230,N_23316,N_23240);
xor U25231 (N_25231,N_23300,N_23319);
and U25232 (N_25232,N_23573,N_23657);
xor U25233 (N_25233,N_22461,N_22238);
nand U25234 (N_25234,N_22436,N_22060);
xnor U25235 (N_25235,N_22288,N_23408);
and U25236 (N_25236,N_23142,N_23683);
or U25237 (N_25237,N_22619,N_22531);
nand U25238 (N_25238,N_22457,N_23082);
nand U25239 (N_25239,N_22969,N_22884);
nand U25240 (N_25240,N_22085,N_22786);
and U25241 (N_25241,N_22411,N_22986);
or U25242 (N_25242,N_22254,N_23435);
or U25243 (N_25243,N_22328,N_23233);
nor U25244 (N_25244,N_22900,N_23545);
nor U25245 (N_25245,N_22368,N_22250);
nor U25246 (N_25246,N_22624,N_23099);
xor U25247 (N_25247,N_22609,N_22058);
or U25248 (N_25248,N_22924,N_23784);
and U25249 (N_25249,N_23086,N_23582);
xnor U25250 (N_25250,N_22402,N_23721);
xnor U25251 (N_25251,N_23162,N_23040);
xnor U25252 (N_25252,N_23536,N_22444);
nand U25253 (N_25253,N_22288,N_22260);
nor U25254 (N_25254,N_22170,N_23131);
or U25255 (N_25255,N_22153,N_22856);
or U25256 (N_25256,N_22604,N_22752);
or U25257 (N_25257,N_23899,N_22781);
or U25258 (N_25258,N_22129,N_23335);
nand U25259 (N_25259,N_23436,N_22336);
and U25260 (N_25260,N_23117,N_22159);
and U25261 (N_25261,N_23225,N_22912);
xor U25262 (N_25262,N_22144,N_23454);
and U25263 (N_25263,N_22042,N_23317);
nor U25264 (N_25264,N_23159,N_22304);
nor U25265 (N_25265,N_23295,N_23565);
or U25266 (N_25266,N_23952,N_23866);
nand U25267 (N_25267,N_23820,N_22449);
nand U25268 (N_25268,N_22433,N_22004);
nor U25269 (N_25269,N_22018,N_23162);
nor U25270 (N_25270,N_23093,N_23118);
nand U25271 (N_25271,N_23528,N_22944);
nand U25272 (N_25272,N_23363,N_23931);
nand U25273 (N_25273,N_23144,N_23607);
nand U25274 (N_25274,N_22345,N_23145);
nand U25275 (N_25275,N_22751,N_23472);
and U25276 (N_25276,N_23127,N_22313);
nor U25277 (N_25277,N_23386,N_23443);
and U25278 (N_25278,N_22261,N_22811);
nand U25279 (N_25279,N_23421,N_22398);
nor U25280 (N_25280,N_22374,N_22168);
nor U25281 (N_25281,N_22129,N_22959);
xnor U25282 (N_25282,N_23172,N_22245);
or U25283 (N_25283,N_22507,N_22228);
or U25284 (N_25284,N_22775,N_23603);
or U25285 (N_25285,N_23229,N_23522);
and U25286 (N_25286,N_22204,N_23285);
nand U25287 (N_25287,N_22464,N_22841);
nor U25288 (N_25288,N_23441,N_22127);
or U25289 (N_25289,N_22750,N_22039);
nor U25290 (N_25290,N_23158,N_23794);
nand U25291 (N_25291,N_23268,N_23042);
xnor U25292 (N_25292,N_22125,N_23666);
or U25293 (N_25293,N_22652,N_22422);
nand U25294 (N_25294,N_22591,N_23244);
and U25295 (N_25295,N_23673,N_23615);
nor U25296 (N_25296,N_22326,N_23722);
nor U25297 (N_25297,N_22800,N_22407);
and U25298 (N_25298,N_22455,N_22669);
xnor U25299 (N_25299,N_23944,N_22183);
xor U25300 (N_25300,N_22838,N_23039);
or U25301 (N_25301,N_23220,N_22198);
xor U25302 (N_25302,N_22570,N_23915);
nand U25303 (N_25303,N_22792,N_23561);
and U25304 (N_25304,N_22565,N_23587);
and U25305 (N_25305,N_23253,N_22032);
xnor U25306 (N_25306,N_23864,N_22694);
or U25307 (N_25307,N_22991,N_22594);
and U25308 (N_25308,N_22386,N_23769);
nor U25309 (N_25309,N_23222,N_22725);
and U25310 (N_25310,N_22873,N_23740);
or U25311 (N_25311,N_23804,N_22496);
xnor U25312 (N_25312,N_23030,N_23333);
and U25313 (N_25313,N_23818,N_23579);
and U25314 (N_25314,N_23864,N_23190);
nand U25315 (N_25315,N_23797,N_23058);
nor U25316 (N_25316,N_23712,N_23456);
and U25317 (N_25317,N_22631,N_22353);
or U25318 (N_25318,N_22549,N_22758);
xor U25319 (N_25319,N_22867,N_23242);
xor U25320 (N_25320,N_23966,N_23021);
or U25321 (N_25321,N_23106,N_22234);
xor U25322 (N_25322,N_22414,N_22946);
nand U25323 (N_25323,N_22741,N_23641);
or U25324 (N_25324,N_23619,N_23607);
and U25325 (N_25325,N_23408,N_23756);
or U25326 (N_25326,N_22323,N_22528);
nor U25327 (N_25327,N_23799,N_22227);
xnor U25328 (N_25328,N_23102,N_23427);
and U25329 (N_25329,N_23122,N_23572);
or U25330 (N_25330,N_23904,N_22904);
nand U25331 (N_25331,N_23834,N_23559);
or U25332 (N_25332,N_23690,N_23767);
and U25333 (N_25333,N_23003,N_23498);
nor U25334 (N_25334,N_22455,N_23630);
nor U25335 (N_25335,N_23459,N_23401);
nor U25336 (N_25336,N_23184,N_22261);
xnor U25337 (N_25337,N_23986,N_23621);
xor U25338 (N_25338,N_22712,N_23413);
nand U25339 (N_25339,N_23484,N_23593);
nand U25340 (N_25340,N_23746,N_22430);
and U25341 (N_25341,N_23710,N_23469);
and U25342 (N_25342,N_22319,N_23983);
and U25343 (N_25343,N_22958,N_23963);
nand U25344 (N_25344,N_22584,N_22171);
or U25345 (N_25345,N_23980,N_22615);
nand U25346 (N_25346,N_22067,N_23842);
and U25347 (N_25347,N_23619,N_22229);
and U25348 (N_25348,N_23961,N_23778);
nor U25349 (N_25349,N_22647,N_22616);
xnor U25350 (N_25350,N_22586,N_23497);
and U25351 (N_25351,N_23570,N_22405);
nor U25352 (N_25352,N_23197,N_22680);
or U25353 (N_25353,N_23862,N_23176);
nand U25354 (N_25354,N_23282,N_22109);
or U25355 (N_25355,N_23361,N_23263);
or U25356 (N_25356,N_22422,N_22980);
or U25357 (N_25357,N_23865,N_23746);
or U25358 (N_25358,N_23532,N_22839);
nand U25359 (N_25359,N_22598,N_22864);
nor U25360 (N_25360,N_23057,N_23827);
nor U25361 (N_25361,N_22861,N_23138);
nand U25362 (N_25362,N_23041,N_23706);
xnor U25363 (N_25363,N_22271,N_23361);
xor U25364 (N_25364,N_23495,N_23865);
or U25365 (N_25365,N_22041,N_23868);
nand U25366 (N_25366,N_22077,N_23714);
nor U25367 (N_25367,N_23256,N_23875);
xnor U25368 (N_25368,N_23801,N_23853);
nor U25369 (N_25369,N_22638,N_22130);
xor U25370 (N_25370,N_23276,N_23619);
and U25371 (N_25371,N_22512,N_23517);
xnor U25372 (N_25372,N_23637,N_22276);
nand U25373 (N_25373,N_22830,N_22485);
nor U25374 (N_25374,N_22901,N_22795);
and U25375 (N_25375,N_23354,N_22847);
xor U25376 (N_25376,N_22173,N_23456);
xnor U25377 (N_25377,N_22754,N_23650);
or U25378 (N_25378,N_23292,N_22457);
xor U25379 (N_25379,N_22745,N_23795);
nand U25380 (N_25380,N_22228,N_22138);
nor U25381 (N_25381,N_22326,N_23304);
xnor U25382 (N_25382,N_22546,N_22601);
xnor U25383 (N_25383,N_22398,N_23114);
nor U25384 (N_25384,N_23807,N_23832);
nand U25385 (N_25385,N_22232,N_23377);
and U25386 (N_25386,N_23742,N_22105);
nand U25387 (N_25387,N_22214,N_22079);
nand U25388 (N_25388,N_22179,N_22962);
xnor U25389 (N_25389,N_22762,N_23318);
nor U25390 (N_25390,N_22006,N_22927);
nand U25391 (N_25391,N_22332,N_22064);
xor U25392 (N_25392,N_22903,N_22800);
nor U25393 (N_25393,N_23351,N_22852);
and U25394 (N_25394,N_23534,N_23511);
xnor U25395 (N_25395,N_22150,N_22830);
xor U25396 (N_25396,N_22402,N_23180);
nor U25397 (N_25397,N_23149,N_22742);
and U25398 (N_25398,N_23328,N_22246);
or U25399 (N_25399,N_23327,N_22915);
xnor U25400 (N_25400,N_23278,N_22905);
nor U25401 (N_25401,N_22506,N_22839);
nor U25402 (N_25402,N_23431,N_23802);
nor U25403 (N_25403,N_23254,N_22791);
nand U25404 (N_25404,N_23408,N_22404);
and U25405 (N_25405,N_23846,N_23175);
or U25406 (N_25406,N_23342,N_23158);
and U25407 (N_25407,N_23111,N_23796);
or U25408 (N_25408,N_22086,N_23727);
nor U25409 (N_25409,N_22173,N_23398);
and U25410 (N_25410,N_23981,N_23748);
nand U25411 (N_25411,N_22981,N_23725);
xnor U25412 (N_25412,N_22385,N_22784);
and U25413 (N_25413,N_22081,N_23127);
and U25414 (N_25414,N_23941,N_23412);
and U25415 (N_25415,N_22035,N_22063);
xor U25416 (N_25416,N_22372,N_23793);
xnor U25417 (N_25417,N_22428,N_23304);
nor U25418 (N_25418,N_23153,N_22016);
and U25419 (N_25419,N_22379,N_23080);
or U25420 (N_25420,N_23247,N_23182);
nand U25421 (N_25421,N_23893,N_22124);
or U25422 (N_25422,N_23419,N_22475);
nor U25423 (N_25423,N_23535,N_22564);
or U25424 (N_25424,N_23230,N_22069);
or U25425 (N_25425,N_22268,N_23703);
nor U25426 (N_25426,N_22890,N_23453);
and U25427 (N_25427,N_22048,N_22689);
or U25428 (N_25428,N_23345,N_22369);
or U25429 (N_25429,N_23347,N_22151);
or U25430 (N_25430,N_22356,N_22771);
or U25431 (N_25431,N_22547,N_22408);
nor U25432 (N_25432,N_23208,N_22645);
xor U25433 (N_25433,N_23882,N_23225);
or U25434 (N_25434,N_23078,N_23543);
and U25435 (N_25435,N_22780,N_23900);
nor U25436 (N_25436,N_22884,N_23491);
or U25437 (N_25437,N_22026,N_23428);
and U25438 (N_25438,N_23663,N_23112);
or U25439 (N_25439,N_22867,N_22756);
xor U25440 (N_25440,N_23503,N_23495);
xor U25441 (N_25441,N_23491,N_22875);
and U25442 (N_25442,N_23543,N_22714);
xor U25443 (N_25443,N_23501,N_22040);
or U25444 (N_25444,N_22807,N_22526);
nor U25445 (N_25445,N_22618,N_22747);
xnor U25446 (N_25446,N_22454,N_23252);
or U25447 (N_25447,N_22518,N_23842);
or U25448 (N_25448,N_22577,N_23960);
or U25449 (N_25449,N_23257,N_23042);
nand U25450 (N_25450,N_23242,N_23269);
nand U25451 (N_25451,N_23736,N_22955);
and U25452 (N_25452,N_23120,N_22545);
nand U25453 (N_25453,N_22103,N_22192);
or U25454 (N_25454,N_23538,N_22312);
nand U25455 (N_25455,N_23846,N_22073);
or U25456 (N_25456,N_22903,N_23037);
or U25457 (N_25457,N_23256,N_22882);
nor U25458 (N_25458,N_23313,N_23656);
and U25459 (N_25459,N_23556,N_23622);
or U25460 (N_25460,N_22783,N_23225);
nor U25461 (N_25461,N_23620,N_22441);
nor U25462 (N_25462,N_22094,N_23599);
nor U25463 (N_25463,N_22138,N_22524);
nor U25464 (N_25464,N_23509,N_23917);
nand U25465 (N_25465,N_23404,N_22148);
or U25466 (N_25466,N_23621,N_23871);
nand U25467 (N_25467,N_23329,N_23259);
and U25468 (N_25468,N_22965,N_23219);
or U25469 (N_25469,N_22005,N_22884);
xor U25470 (N_25470,N_22504,N_22734);
nor U25471 (N_25471,N_23552,N_23817);
or U25472 (N_25472,N_23926,N_22536);
xor U25473 (N_25473,N_23283,N_23161);
nor U25474 (N_25474,N_22477,N_22699);
or U25475 (N_25475,N_22834,N_23618);
or U25476 (N_25476,N_22407,N_22567);
and U25477 (N_25477,N_22660,N_23768);
or U25478 (N_25478,N_22332,N_23060);
nand U25479 (N_25479,N_22816,N_23054);
nand U25480 (N_25480,N_23293,N_23246);
nor U25481 (N_25481,N_22245,N_22552);
nand U25482 (N_25482,N_23690,N_23274);
and U25483 (N_25483,N_22592,N_22788);
and U25484 (N_25484,N_23770,N_22404);
and U25485 (N_25485,N_23215,N_22475);
or U25486 (N_25486,N_23236,N_22511);
or U25487 (N_25487,N_22494,N_22574);
and U25488 (N_25488,N_22831,N_23716);
xnor U25489 (N_25489,N_22962,N_23970);
nor U25490 (N_25490,N_23911,N_22936);
nor U25491 (N_25491,N_23185,N_22585);
nand U25492 (N_25492,N_23868,N_22400);
nor U25493 (N_25493,N_23247,N_23909);
xnor U25494 (N_25494,N_22606,N_22557);
nand U25495 (N_25495,N_23657,N_22414);
xnor U25496 (N_25496,N_22250,N_22686);
and U25497 (N_25497,N_22240,N_23761);
and U25498 (N_25498,N_22041,N_23969);
xor U25499 (N_25499,N_23370,N_23243);
and U25500 (N_25500,N_22567,N_22203);
and U25501 (N_25501,N_22727,N_23221);
and U25502 (N_25502,N_22881,N_22350);
nor U25503 (N_25503,N_23730,N_23241);
xor U25504 (N_25504,N_22051,N_23038);
and U25505 (N_25505,N_23263,N_23078);
or U25506 (N_25506,N_23988,N_22078);
xor U25507 (N_25507,N_22875,N_23824);
and U25508 (N_25508,N_23228,N_23498);
and U25509 (N_25509,N_22416,N_22508);
xnor U25510 (N_25510,N_23145,N_22721);
and U25511 (N_25511,N_22025,N_22437);
nand U25512 (N_25512,N_23885,N_22503);
or U25513 (N_25513,N_23277,N_22597);
and U25514 (N_25514,N_22804,N_22440);
nor U25515 (N_25515,N_23157,N_22099);
or U25516 (N_25516,N_23764,N_22294);
and U25517 (N_25517,N_22232,N_22119);
and U25518 (N_25518,N_22505,N_23186);
xnor U25519 (N_25519,N_23839,N_23849);
or U25520 (N_25520,N_22265,N_23922);
xor U25521 (N_25521,N_22572,N_23148);
nand U25522 (N_25522,N_23465,N_23570);
xnor U25523 (N_25523,N_23069,N_23672);
nand U25524 (N_25524,N_23672,N_22087);
xor U25525 (N_25525,N_22984,N_23137);
nand U25526 (N_25526,N_23990,N_23704);
nor U25527 (N_25527,N_23948,N_23660);
nor U25528 (N_25528,N_22889,N_23066);
and U25529 (N_25529,N_22290,N_22912);
and U25530 (N_25530,N_23966,N_22774);
or U25531 (N_25531,N_22236,N_22578);
nor U25532 (N_25532,N_23857,N_22057);
nor U25533 (N_25533,N_22357,N_23086);
nor U25534 (N_25534,N_23657,N_23077);
xnor U25535 (N_25535,N_22193,N_22149);
or U25536 (N_25536,N_23091,N_23120);
and U25537 (N_25537,N_23091,N_23845);
or U25538 (N_25538,N_23094,N_23023);
or U25539 (N_25539,N_22557,N_23970);
nor U25540 (N_25540,N_22685,N_22937);
or U25541 (N_25541,N_23981,N_22637);
nor U25542 (N_25542,N_23878,N_22990);
or U25543 (N_25543,N_22098,N_23107);
or U25544 (N_25544,N_23371,N_22586);
or U25545 (N_25545,N_22854,N_23276);
xor U25546 (N_25546,N_23334,N_22774);
nand U25547 (N_25547,N_22710,N_22017);
and U25548 (N_25548,N_23341,N_22875);
xor U25549 (N_25549,N_23823,N_22565);
xor U25550 (N_25550,N_23507,N_22078);
nor U25551 (N_25551,N_22424,N_23763);
xnor U25552 (N_25552,N_22134,N_22827);
nor U25553 (N_25553,N_22549,N_22419);
or U25554 (N_25554,N_22924,N_22228);
nand U25555 (N_25555,N_23902,N_22973);
nand U25556 (N_25556,N_23077,N_23360);
xnor U25557 (N_25557,N_23452,N_22611);
or U25558 (N_25558,N_22023,N_22266);
xor U25559 (N_25559,N_22155,N_23789);
or U25560 (N_25560,N_22133,N_23336);
nor U25561 (N_25561,N_22395,N_23418);
nand U25562 (N_25562,N_22724,N_23716);
nand U25563 (N_25563,N_23200,N_22539);
or U25564 (N_25564,N_23098,N_23686);
nand U25565 (N_25565,N_23438,N_22297);
and U25566 (N_25566,N_23903,N_22331);
nand U25567 (N_25567,N_23072,N_22273);
nor U25568 (N_25568,N_22911,N_22980);
xor U25569 (N_25569,N_22298,N_23741);
or U25570 (N_25570,N_22823,N_22839);
nor U25571 (N_25571,N_23408,N_23335);
xor U25572 (N_25572,N_22398,N_22389);
nor U25573 (N_25573,N_22659,N_22453);
xor U25574 (N_25574,N_23755,N_22192);
nand U25575 (N_25575,N_23005,N_23510);
and U25576 (N_25576,N_22452,N_22921);
nand U25577 (N_25577,N_22137,N_22808);
and U25578 (N_25578,N_22768,N_22341);
and U25579 (N_25579,N_22573,N_23798);
nor U25580 (N_25580,N_22019,N_23197);
nor U25581 (N_25581,N_23735,N_23087);
or U25582 (N_25582,N_23921,N_23745);
xor U25583 (N_25583,N_22362,N_23736);
xor U25584 (N_25584,N_23644,N_23688);
xor U25585 (N_25585,N_22006,N_23423);
nor U25586 (N_25586,N_22593,N_22818);
or U25587 (N_25587,N_22740,N_23502);
nor U25588 (N_25588,N_22918,N_23004);
xnor U25589 (N_25589,N_22632,N_23909);
nand U25590 (N_25590,N_22310,N_22259);
and U25591 (N_25591,N_22194,N_22928);
and U25592 (N_25592,N_23662,N_23035);
or U25593 (N_25593,N_22883,N_22730);
nand U25594 (N_25594,N_23186,N_23608);
xnor U25595 (N_25595,N_23655,N_22297);
and U25596 (N_25596,N_22260,N_22603);
nor U25597 (N_25597,N_22513,N_23552);
nor U25598 (N_25598,N_23239,N_23348);
and U25599 (N_25599,N_22395,N_22408);
nand U25600 (N_25600,N_23218,N_22264);
xnor U25601 (N_25601,N_23372,N_22131);
nand U25602 (N_25602,N_23125,N_22573);
nor U25603 (N_25603,N_22233,N_22062);
nand U25604 (N_25604,N_23033,N_22916);
or U25605 (N_25605,N_23538,N_23723);
xnor U25606 (N_25606,N_22404,N_22874);
nor U25607 (N_25607,N_23671,N_22812);
nand U25608 (N_25608,N_22852,N_22641);
nor U25609 (N_25609,N_23123,N_23928);
and U25610 (N_25610,N_22793,N_22401);
nor U25611 (N_25611,N_22918,N_22874);
nor U25612 (N_25612,N_22625,N_23143);
xor U25613 (N_25613,N_22665,N_22463);
nor U25614 (N_25614,N_23664,N_22252);
xor U25615 (N_25615,N_23473,N_23672);
and U25616 (N_25616,N_22996,N_22822);
xor U25617 (N_25617,N_23621,N_22789);
nor U25618 (N_25618,N_23084,N_22926);
or U25619 (N_25619,N_23823,N_22107);
nand U25620 (N_25620,N_22733,N_22441);
nor U25621 (N_25621,N_23040,N_22587);
and U25622 (N_25622,N_23337,N_23766);
xor U25623 (N_25623,N_22715,N_22009);
or U25624 (N_25624,N_22896,N_23863);
nand U25625 (N_25625,N_22418,N_23697);
nand U25626 (N_25626,N_23142,N_22059);
nand U25627 (N_25627,N_22436,N_23225);
xor U25628 (N_25628,N_22410,N_23243);
nor U25629 (N_25629,N_22432,N_22973);
nor U25630 (N_25630,N_22676,N_22817);
nor U25631 (N_25631,N_23306,N_23453);
or U25632 (N_25632,N_22424,N_23593);
or U25633 (N_25633,N_23212,N_22138);
xnor U25634 (N_25634,N_22090,N_23889);
and U25635 (N_25635,N_23672,N_23512);
and U25636 (N_25636,N_22122,N_22022);
nor U25637 (N_25637,N_23905,N_23835);
xor U25638 (N_25638,N_22956,N_22421);
and U25639 (N_25639,N_22134,N_22729);
nand U25640 (N_25640,N_23276,N_23998);
nand U25641 (N_25641,N_22447,N_22080);
and U25642 (N_25642,N_23193,N_22326);
xnor U25643 (N_25643,N_23884,N_23786);
nand U25644 (N_25644,N_22968,N_22211);
or U25645 (N_25645,N_23123,N_23023);
and U25646 (N_25646,N_23321,N_22910);
or U25647 (N_25647,N_23644,N_23410);
and U25648 (N_25648,N_23486,N_23586);
or U25649 (N_25649,N_23192,N_23535);
nor U25650 (N_25650,N_22323,N_22873);
nor U25651 (N_25651,N_23795,N_23696);
and U25652 (N_25652,N_22013,N_23422);
and U25653 (N_25653,N_22268,N_22060);
and U25654 (N_25654,N_23863,N_23802);
nor U25655 (N_25655,N_22421,N_22480);
and U25656 (N_25656,N_22138,N_23625);
and U25657 (N_25657,N_23054,N_22315);
and U25658 (N_25658,N_23376,N_22727);
and U25659 (N_25659,N_23966,N_22997);
nand U25660 (N_25660,N_23936,N_23488);
nand U25661 (N_25661,N_23088,N_23868);
or U25662 (N_25662,N_23919,N_23814);
nand U25663 (N_25663,N_23459,N_22475);
xnor U25664 (N_25664,N_22841,N_23745);
nand U25665 (N_25665,N_23806,N_22084);
nor U25666 (N_25666,N_22113,N_22255);
nand U25667 (N_25667,N_23612,N_22306);
nor U25668 (N_25668,N_22910,N_23706);
and U25669 (N_25669,N_23651,N_23746);
nor U25670 (N_25670,N_23219,N_22327);
or U25671 (N_25671,N_22287,N_22051);
xnor U25672 (N_25672,N_22933,N_22977);
xor U25673 (N_25673,N_23774,N_22846);
nand U25674 (N_25674,N_23236,N_23332);
or U25675 (N_25675,N_22781,N_22280);
nor U25676 (N_25676,N_23241,N_22132);
or U25677 (N_25677,N_22866,N_23437);
and U25678 (N_25678,N_23984,N_22029);
and U25679 (N_25679,N_22399,N_23111);
and U25680 (N_25680,N_22207,N_22465);
or U25681 (N_25681,N_22989,N_23901);
xor U25682 (N_25682,N_22714,N_23636);
or U25683 (N_25683,N_22993,N_22500);
xor U25684 (N_25684,N_23154,N_22922);
nor U25685 (N_25685,N_22923,N_23995);
nand U25686 (N_25686,N_22908,N_22573);
or U25687 (N_25687,N_22460,N_23300);
or U25688 (N_25688,N_23351,N_23010);
xor U25689 (N_25689,N_23547,N_23100);
xnor U25690 (N_25690,N_22920,N_23273);
or U25691 (N_25691,N_22099,N_23508);
nor U25692 (N_25692,N_22066,N_22820);
and U25693 (N_25693,N_23192,N_23269);
and U25694 (N_25694,N_23371,N_23596);
and U25695 (N_25695,N_22905,N_22247);
or U25696 (N_25696,N_23965,N_22760);
nand U25697 (N_25697,N_23413,N_22670);
and U25698 (N_25698,N_23374,N_22453);
xor U25699 (N_25699,N_22427,N_23058);
nand U25700 (N_25700,N_23482,N_23808);
nand U25701 (N_25701,N_23873,N_23823);
nand U25702 (N_25702,N_23902,N_22939);
xor U25703 (N_25703,N_23917,N_23219);
or U25704 (N_25704,N_23274,N_22568);
or U25705 (N_25705,N_23999,N_23391);
or U25706 (N_25706,N_22304,N_23534);
or U25707 (N_25707,N_23201,N_23435);
or U25708 (N_25708,N_22856,N_22778);
or U25709 (N_25709,N_22937,N_23664);
or U25710 (N_25710,N_22882,N_22538);
and U25711 (N_25711,N_23883,N_22394);
or U25712 (N_25712,N_22559,N_23400);
nand U25713 (N_25713,N_23043,N_23840);
and U25714 (N_25714,N_23823,N_22663);
or U25715 (N_25715,N_22979,N_23372);
and U25716 (N_25716,N_22241,N_22123);
xnor U25717 (N_25717,N_23810,N_23950);
and U25718 (N_25718,N_22267,N_22394);
xnor U25719 (N_25719,N_23182,N_23044);
nand U25720 (N_25720,N_22439,N_22907);
nor U25721 (N_25721,N_22539,N_23224);
or U25722 (N_25722,N_23786,N_23297);
nor U25723 (N_25723,N_23201,N_22736);
or U25724 (N_25724,N_22645,N_23424);
or U25725 (N_25725,N_22643,N_22067);
nor U25726 (N_25726,N_23737,N_22733);
or U25727 (N_25727,N_22281,N_23721);
nor U25728 (N_25728,N_23115,N_22106);
and U25729 (N_25729,N_22166,N_22887);
xnor U25730 (N_25730,N_22618,N_22191);
or U25731 (N_25731,N_22024,N_22945);
nor U25732 (N_25732,N_22075,N_22122);
nand U25733 (N_25733,N_23709,N_22455);
and U25734 (N_25734,N_22573,N_22440);
or U25735 (N_25735,N_22360,N_22641);
xor U25736 (N_25736,N_22106,N_23933);
nand U25737 (N_25737,N_23103,N_22076);
nand U25738 (N_25738,N_23233,N_23349);
xnor U25739 (N_25739,N_23975,N_22801);
nor U25740 (N_25740,N_22561,N_22421);
nand U25741 (N_25741,N_22911,N_22375);
and U25742 (N_25742,N_23198,N_22263);
nand U25743 (N_25743,N_23590,N_22454);
nor U25744 (N_25744,N_22282,N_22248);
xnor U25745 (N_25745,N_23612,N_22805);
xor U25746 (N_25746,N_22345,N_23461);
or U25747 (N_25747,N_23128,N_23745);
or U25748 (N_25748,N_22280,N_22354);
and U25749 (N_25749,N_22731,N_22048);
xor U25750 (N_25750,N_23087,N_22029);
nor U25751 (N_25751,N_23533,N_23310);
xor U25752 (N_25752,N_23249,N_22073);
or U25753 (N_25753,N_22703,N_22656);
xor U25754 (N_25754,N_23115,N_22641);
nand U25755 (N_25755,N_22672,N_22304);
nand U25756 (N_25756,N_22893,N_23828);
nor U25757 (N_25757,N_22114,N_23826);
nand U25758 (N_25758,N_23508,N_23334);
xor U25759 (N_25759,N_23370,N_23184);
xor U25760 (N_25760,N_22273,N_22391);
and U25761 (N_25761,N_23843,N_23001);
or U25762 (N_25762,N_22447,N_22610);
nand U25763 (N_25763,N_22151,N_23889);
or U25764 (N_25764,N_22663,N_22743);
and U25765 (N_25765,N_22676,N_23728);
xor U25766 (N_25766,N_23527,N_23295);
and U25767 (N_25767,N_23761,N_23815);
and U25768 (N_25768,N_22948,N_22312);
xor U25769 (N_25769,N_22343,N_23887);
nand U25770 (N_25770,N_23243,N_23918);
nor U25771 (N_25771,N_23582,N_23778);
xnor U25772 (N_25772,N_23895,N_22839);
xor U25773 (N_25773,N_23720,N_23770);
xnor U25774 (N_25774,N_22054,N_23443);
xor U25775 (N_25775,N_22250,N_22466);
or U25776 (N_25776,N_23539,N_23781);
nand U25777 (N_25777,N_22196,N_23022);
nor U25778 (N_25778,N_23940,N_22720);
or U25779 (N_25779,N_22643,N_23440);
nor U25780 (N_25780,N_23401,N_22768);
and U25781 (N_25781,N_22497,N_22656);
nand U25782 (N_25782,N_22805,N_23625);
and U25783 (N_25783,N_22105,N_22277);
xor U25784 (N_25784,N_23503,N_23680);
nand U25785 (N_25785,N_22231,N_23031);
xor U25786 (N_25786,N_22254,N_23940);
xnor U25787 (N_25787,N_23872,N_23324);
and U25788 (N_25788,N_22730,N_23491);
xnor U25789 (N_25789,N_23209,N_22502);
or U25790 (N_25790,N_22268,N_22869);
xor U25791 (N_25791,N_22666,N_23770);
and U25792 (N_25792,N_22265,N_23147);
xnor U25793 (N_25793,N_22084,N_22108);
and U25794 (N_25794,N_22872,N_22904);
or U25795 (N_25795,N_22654,N_23479);
nand U25796 (N_25796,N_22836,N_23638);
or U25797 (N_25797,N_22301,N_22458);
xnor U25798 (N_25798,N_22280,N_23932);
and U25799 (N_25799,N_22663,N_22474);
xnor U25800 (N_25800,N_23760,N_22370);
and U25801 (N_25801,N_23139,N_22441);
and U25802 (N_25802,N_23071,N_22666);
xnor U25803 (N_25803,N_23141,N_22814);
nor U25804 (N_25804,N_22315,N_22533);
nor U25805 (N_25805,N_23999,N_22253);
xor U25806 (N_25806,N_22323,N_22682);
and U25807 (N_25807,N_23615,N_22205);
or U25808 (N_25808,N_22111,N_22662);
xnor U25809 (N_25809,N_23285,N_23380);
nand U25810 (N_25810,N_23795,N_22038);
nand U25811 (N_25811,N_22297,N_23979);
nor U25812 (N_25812,N_23641,N_23365);
nand U25813 (N_25813,N_22140,N_23488);
xnor U25814 (N_25814,N_23223,N_23969);
and U25815 (N_25815,N_22346,N_23945);
or U25816 (N_25816,N_23168,N_23442);
or U25817 (N_25817,N_23454,N_22511);
and U25818 (N_25818,N_22381,N_22103);
and U25819 (N_25819,N_22345,N_22432);
xor U25820 (N_25820,N_22187,N_22446);
nor U25821 (N_25821,N_23744,N_22393);
xor U25822 (N_25822,N_23458,N_22614);
xor U25823 (N_25823,N_23344,N_23185);
nor U25824 (N_25824,N_23355,N_22712);
nand U25825 (N_25825,N_23293,N_22506);
and U25826 (N_25826,N_23400,N_23248);
and U25827 (N_25827,N_23936,N_22483);
xor U25828 (N_25828,N_23951,N_22134);
xnor U25829 (N_25829,N_22285,N_23797);
or U25830 (N_25830,N_23682,N_22723);
nand U25831 (N_25831,N_23877,N_22507);
and U25832 (N_25832,N_23812,N_23980);
nand U25833 (N_25833,N_22779,N_23752);
and U25834 (N_25834,N_22362,N_22890);
or U25835 (N_25835,N_22400,N_23118);
and U25836 (N_25836,N_22766,N_23260);
or U25837 (N_25837,N_23511,N_22733);
and U25838 (N_25838,N_22160,N_22086);
or U25839 (N_25839,N_23600,N_23681);
nand U25840 (N_25840,N_22351,N_23306);
nand U25841 (N_25841,N_23621,N_22455);
or U25842 (N_25842,N_22445,N_23415);
nand U25843 (N_25843,N_22731,N_23016);
nand U25844 (N_25844,N_23496,N_23210);
and U25845 (N_25845,N_22311,N_22365);
xnor U25846 (N_25846,N_22735,N_22170);
nand U25847 (N_25847,N_22774,N_22590);
xor U25848 (N_25848,N_22625,N_23751);
nor U25849 (N_25849,N_22354,N_22166);
xnor U25850 (N_25850,N_23776,N_23725);
nand U25851 (N_25851,N_22306,N_22152);
or U25852 (N_25852,N_23126,N_22867);
and U25853 (N_25853,N_23083,N_23167);
nor U25854 (N_25854,N_23774,N_23931);
and U25855 (N_25855,N_22597,N_22549);
and U25856 (N_25856,N_22675,N_22798);
and U25857 (N_25857,N_23203,N_22657);
xnor U25858 (N_25858,N_22387,N_23499);
xnor U25859 (N_25859,N_22511,N_23121);
xor U25860 (N_25860,N_22334,N_22271);
nand U25861 (N_25861,N_22027,N_22255);
nand U25862 (N_25862,N_22059,N_23945);
xor U25863 (N_25863,N_23436,N_22027);
or U25864 (N_25864,N_22790,N_23040);
and U25865 (N_25865,N_23347,N_23523);
and U25866 (N_25866,N_23467,N_23955);
nand U25867 (N_25867,N_22527,N_23205);
nor U25868 (N_25868,N_22851,N_22559);
nand U25869 (N_25869,N_23755,N_23919);
nor U25870 (N_25870,N_22228,N_22012);
xor U25871 (N_25871,N_23264,N_23821);
and U25872 (N_25872,N_23005,N_22135);
nor U25873 (N_25873,N_22132,N_22726);
nor U25874 (N_25874,N_22830,N_22938);
nor U25875 (N_25875,N_23477,N_22461);
nand U25876 (N_25876,N_23052,N_23143);
and U25877 (N_25877,N_23314,N_22573);
xnor U25878 (N_25878,N_22522,N_22352);
or U25879 (N_25879,N_23488,N_23887);
or U25880 (N_25880,N_22874,N_23266);
and U25881 (N_25881,N_23745,N_22131);
nand U25882 (N_25882,N_22405,N_22724);
and U25883 (N_25883,N_22458,N_23133);
and U25884 (N_25884,N_23975,N_22970);
nor U25885 (N_25885,N_23276,N_23910);
and U25886 (N_25886,N_22689,N_23117);
nor U25887 (N_25887,N_23187,N_23799);
xnor U25888 (N_25888,N_23068,N_22823);
xnor U25889 (N_25889,N_22024,N_23518);
xor U25890 (N_25890,N_23567,N_23047);
and U25891 (N_25891,N_22403,N_23199);
nor U25892 (N_25892,N_22573,N_22138);
or U25893 (N_25893,N_23663,N_22437);
or U25894 (N_25894,N_22560,N_23675);
and U25895 (N_25895,N_23629,N_22299);
or U25896 (N_25896,N_22551,N_22008);
xor U25897 (N_25897,N_22360,N_22807);
nand U25898 (N_25898,N_22356,N_22232);
nand U25899 (N_25899,N_22155,N_22693);
and U25900 (N_25900,N_23712,N_23292);
nand U25901 (N_25901,N_23477,N_22702);
xnor U25902 (N_25902,N_23699,N_22344);
and U25903 (N_25903,N_22078,N_22869);
nand U25904 (N_25904,N_22718,N_22687);
or U25905 (N_25905,N_23976,N_23494);
or U25906 (N_25906,N_23785,N_22922);
nor U25907 (N_25907,N_23071,N_22155);
or U25908 (N_25908,N_23199,N_23919);
xor U25909 (N_25909,N_22602,N_22279);
nor U25910 (N_25910,N_23957,N_22188);
nor U25911 (N_25911,N_22838,N_22262);
xor U25912 (N_25912,N_23011,N_22590);
or U25913 (N_25913,N_23524,N_23495);
and U25914 (N_25914,N_23199,N_23812);
nor U25915 (N_25915,N_23403,N_23354);
xor U25916 (N_25916,N_22917,N_22516);
nor U25917 (N_25917,N_22874,N_23365);
or U25918 (N_25918,N_22865,N_22768);
nand U25919 (N_25919,N_22484,N_23299);
nand U25920 (N_25920,N_23714,N_22180);
nor U25921 (N_25921,N_22100,N_23952);
xor U25922 (N_25922,N_23517,N_23875);
or U25923 (N_25923,N_23570,N_22101);
xnor U25924 (N_25924,N_22782,N_23610);
or U25925 (N_25925,N_23450,N_23090);
xnor U25926 (N_25926,N_23328,N_23818);
xnor U25927 (N_25927,N_23509,N_23538);
or U25928 (N_25928,N_23467,N_23066);
nand U25929 (N_25929,N_23298,N_22860);
nor U25930 (N_25930,N_22860,N_22855);
nor U25931 (N_25931,N_23667,N_22376);
or U25932 (N_25932,N_23450,N_23123);
xnor U25933 (N_25933,N_22253,N_22069);
xnor U25934 (N_25934,N_23622,N_22896);
xnor U25935 (N_25935,N_22452,N_23681);
or U25936 (N_25936,N_22214,N_23874);
nor U25937 (N_25937,N_22978,N_23977);
and U25938 (N_25938,N_23408,N_22930);
nor U25939 (N_25939,N_22450,N_22205);
xnor U25940 (N_25940,N_22225,N_23973);
xor U25941 (N_25941,N_23543,N_23630);
or U25942 (N_25942,N_23058,N_22862);
xor U25943 (N_25943,N_23143,N_22578);
nor U25944 (N_25944,N_22748,N_22588);
nand U25945 (N_25945,N_22067,N_22564);
or U25946 (N_25946,N_22455,N_23930);
xor U25947 (N_25947,N_23643,N_22474);
and U25948 (N_25948,N_23674,N_23146);
and U25949 (N_25949,N_22141,N_22465);
nand U25950 (N_25950,N_22669,N_23255);
nor U25951 (N_25951,N_23286,N_23504);
or U25952 (N_25952,N_23115,N_23740);
nand U25953 (N_25953,N_23120,N_23611);
xnor U25954 (N_25954,N_22139,N_22231);
xor U25955 (N_25955,N_23453,N_22716);
xnor U25956 (N_25956,N_22462,N_23689);
nand U25957 (N_25957,N_22883,N_23258);
or U25958 (N_25958,N_23423,N_22274);
or U25959 (N_25959,N_22327,N_22208);
or U25960 (N_25960,N_22349,N_23476);
xor U25961 (N_25961,N_22924,N_23646);
nand U25962 (N_25962,N_23058,N_23921);
and U25963 (N_25963,N_22020,N_23630);
xnor U25964 (N_25964,N_22269,N_23553);
nand U25965 (N_25965,N_22995,N_23660);
or U25966 (N_25966,N_23108,N_23232);
nor U25967 (N_25967,N_22673,N_23309);
and U25968 (N_25968,N_23178,N_22355);
nor U25969 (N_25969,N_23111,N_22768);
or U25970 (N_25970,N_23045,N_23687);
or U25971 (N_25971,N_23518,N_22029);
xor U25972 (N_25972,N_22618,N_23156);
nor U25973 (N_25973,N_22361,N_23403);
or U25974 (N_25974,N_22078,N_22251);
and U25975 (N_25975,N_23409,N_22598);
nand U25976 (N_25976,N_22437,N_23761);
xnor U25977 (N_25977,N_22625,N_22953);
nor U25978 (N_25978,N_23225,N_23277);
nor U25979 (N_25979,N_22926,N_23161);
nand U25980 (N_25980,N_23564,N_23796);
and U25981 (N_25981,N_23590,N_23930);
and U25982 (N_25982,N_22694,N_22796);
or U25983 (N_25983,N_22942,N_23063);
xnor U25984 (N_25984,N_22727,N_23436);
nand U25985 (N_25985,N_22308,N_22364);
nand U25986 (N_25986,N_22767,N_23274);
or U25987 (N_25987,N_23584,N_22974);
and U25988 (N_25988,N_22781,N_23090);
xnor U25989 (N_25989,N_23395,N_22756);
nor U25990 (N_25990,N_23742,N_23223);
nand U25991 (N_25991,N_22645,N_22602);
nand U25992 (N_25992,N_23468,N_22488);
xnor U25993 (N_25993,N_23091,N_23507);
or U25994 (N_25994,N_22428,N_23871);
nor U25995 (N_25995,N_22149,N_22904);
or U25996 (N_25996,N_22252,N_23989);
nand U25997 (N_25997,N_23007,N_23489);
or U25998 (N_25998,N_22102,N_23630);
or U25999 (N_25999,N_23204,N_22796);
nor U26000 (N_26000,N_25841,N_24667);
and U26001 (N_26001,N_25474,N_25060);
nand U26002 (N_26002,N_24162,N_25146);
nand U26003 (N_26003,N_25909,N_24619);
nand U26004 (N_26004,N_25508,N_24399);
xnor U26005 (N_26005,N_25512,N_25201);
or U26006 (N_26006,N_25237,N_24472);
nor U26007 (N_26007,N_24509,N_24705);
nand U26008 (N_26008,N_25916,N_25231);
and U26009 (N_26009,N_25156,N_24878);
and U26010 (N_26010,N_25453,N_24304);
and U26011 (N_26011,N_25264,N_25406);
nand U26012 (N_26012,N_25690,N_25248);
nand U26013 (N_26013,N_25731,N_24531);
or U26014 (N_26014,N_25280,N_25509);
nor U26015 (N_26015,N_25135,N_24672);
and U26016 (N_26016,N_25739,N_24676);
xor U26017 (N_26017,N_24929,N_25853);
nor U26018 (N_26018,N_25399,N_24490);
xor U26019 (N_26019,N_25669,N_24152);
or U26020 (N_26020,N_24328,N_24961);
and U26021 (N_26021,N_24376,N_24319);
xor U26022 (N_26022,N_24639,N_24147);
nand U26023 (N_26023,N_25210,N_24566);
and U26024 (N_26024,N_25151,N_25796);
nand U26025 (N_26025,N_24471,N_24335);
nand U26026 (N_26026,N_24284,N_24589);
nand U26027 (N_26027,N_25548,N_24675);
nand U26028 (N_26028,N_24151,N_25945);
xor U26029 (N_26029,N_25689,N_25500);
nand U26030 (N_26030,N_24287,N_25554);
or U26031 (N_26031,N_25794,N_25908);
nor U26032 (N_26032,N_24167,N_25461);
or U26033 (N_26033,N_24852,N_25137);
or U26034 (N_26034,N_24489,N_25769);
nor U26035 (N_26035,N_25953,N_25995);
and U26036 (N_26036,N_25486,N_25812);
and U26037 (N_26037,N_25779,N_25589);
and U26038 (N_26038,N_25318,N_24880);
nand U26039 (N_26039,N_24032,N_24617);
xnor U26040 (N_26040,N_24782,N_25714);
or U26041 (N_26041,N_24160,N_24945);
and U26042 (N_26042,N_24495,N_25143);
and U26043 (N_26043,N_24336,N_25692);
nor U26044 (N_26044,N_24425,N_24468);
or U26045 (N_26045,N_25417,N_25282);
xor U26046 (N_26046,N_25829,N_24516);
and U26047 (N_26047,N_25907,N_25065);
xor U26048 (N_26048,N_25362,N_24819);
nor U26049 (N_26049,N_25022,N_25054);
xor U26050 (N_26050,N_25418,N_24135);
or U26051 (N_26051,N_24383,N_25895);
nand U26052 (N_26052,N_24792,N_25090);
or U26053 (N_26053,N_25860,N_25477);
xor U26054 (N_26054,N_24749,N_25758);
xor U26055 (N_26055,N_25064,N_24657);
or U26056 (N_26056,N_25420,N_25899);
xnor U26057 (N_26057,N_24753,N_24706);
and U26058 (N_26058,N_24751,N_24034);
xor U26059 (N_26059,N_25943,N_24913);
nor U26060 (N_26060,N_25319,N_25212);
nor U26061 (N_26061,N_25638,N_24708);
and U26062 (N_26062,N_25034,N_24485);
nand U26063 (N_26063,N_24189,N_24626);
or U26064 (N_26064,N_24402,N_25506);
nand U26065 (N_26065,N_25541,N_24208);
and U26066 (N_26066,N_25504,N_24111);
xor U26067 (N_26067,N_25973,N_24642);
nor U26068 (N_26068,N_24637,N_25910);
nand U26069 (N_26069,N_24380,N_24165);
or U26070 (N_26070,N_25425,N_25919);
xor U26071 (N_26071,N_24567,N_24652);
nor U26072 (N_26072,N_24312,N_24501);
or U26073 (N_26073,N_24584,N_25685);
and U26074 (N_26074,N_25701,N_24768);
nor U26075 (N_26075,N_25781,N_25936);
or U26076 (N_26076,N_24858,N_25178);
nor U26077 (N_26077,N_25869,N_24901);
and U26078 (N_26078,N_25791,N_25481);
nand U26079 (N_26079,N_24272,N_25790);
or U26080 (N_26080,N_24222,N_24552);
xor U26081 (N_26081,N_24663,N_25242);
xnor U26082 (N_26082,N_24710,N_25507);
and U26083 (N_26083,N_25476,N_24839);
or U26084 (N_26084,N_24213,N_24220);
nand U26085 (N_26085,N_25235,N_25009);
nor U26086 (N_26086,N_24510,N_24930);
or U26087 (N_26087,N_25094,N_24403);
and U26088 (N_26088,N_25160,N_24551);
xor U26089 (N_26089,N_24983,N_25302);
nor U26090 (N_26090,N_24294,N_24178);
nor U26091 (N_26091,N_24291,N_24175);
and U26092 (N_26092,N_25691,N_24799);
nor U26093 (N_26093,N_25587,N_24355);
xor U26094 (N_26094,N_24440,N_25913);
xor U26095 (N_26095,N_24326,N_25566);
and U26096 (N_26096,N_24217,N_24354);
xnor U26097 (N_26097,N_24124,N_25260);
nand U26098 (N_26098,N_25838,N_24201);
nand U26099 (N_26099,N_25753,N_25165);
and U26100 (N_26100,N_24691,N_25721);
or U26101 (N_26101,N_25658,N_24150);
nand U26102 (N_26102,N_24816,N_25882);
and U26103 (N_26103,N_25357,N_25815);
or U26104 (N_26104,N_24451,N_24070);
nand U26105 (N_26105,N_24965,N_24919);
nor U26106 (N_26106,N_25710,N_24997);
xor U26107 (N_26107,N_24194,N_25773);
and U26108 (N_26108,N_24862,N_25540);
and U26109 (N_26109,N_25098,N_25141);
and U26110 (N_26110,N_25778,N_25674);
or U26111 (N_26111,N_25881,N_24163);
and U26112 (N_26112,N_24948,N_24814);
nor U26113 (N_26113,N_24624,N_24779);
nand U26114 (N_26114,N_25407,N_24288);
xor U26115 (N_26115,N_24352,N_24685);
xnor U26116 (N_26116,N_25513,N_24851);
or U26117 (N_26117,N_24716,N_24736);
xor U26118 (N_26118,N_24558,N_25561);
xor U26119 (N_26119,N_24737,N_24271);
and U26120 (N_26120,N_24121,N_25615);
nor U26121 (N_26121,N_25804,N_24726);
nand U26122 (N_26122,N_24683,N_25765);
xnor U26123 (N_26123,N_25965,N_24992);
xor U26124 (N_26124,N_25074,N_25050);
or U26125 (N_26125,N_25107,N_24955);
nand U26126 (N_26126,N_25670,N_25221);
or U26127 (N_26127,N_25680,N_25783);
xnor U26128 (N_26128,N_25777,N_25263);
nand U26129 (N_26129,N_24023,N_25770);
xor U26130 (N_26130,N_24803,N_25432);
nand U26131 (N_26131,N_25331,N_24231);
nand U26132 (N_26132,N_24800,N_24872);
nor U26133 (N_26133,N_24718,N_25787);
and U26134 (N_26134,N_25904,N_24105);
nand U26135 (N_26135,N_24944,N_24068);
xor U26136 (N_26136,N_24266,N_25459);
nor U26137 (N_26137,N_24798,N_25121);
and U26138 (N_26138,N_24921,N_25660);
and U26139 (N_26139,N_25713,N_25194);
nand U26140 (N_26140,N_25093,N_25903);
and U26141 (N_26141,N_24707,N_25768);
or U26142 (N_26142,N_25693,N_25188);
nor U26143 (N_26143,N_24602,N_24957);
xor U26144 (N_26144,N_25682,N_25257);
nor U26145 (N_26145,N_25799,N_25709);
nor U26146 (N_26146,N_24596,N_25169);
xor U26147 (N_26147,N_25468,N_24137);
and U26148 (N_26148,N_24869,N_24534);
nor U26149 (N_26149,N_24661,N_24318);
nand U26150 (N_26150,N_24140,N_24629);
nand U26151 (N_26151,N_24313,N_24416);
xnor U26152 (N_26152,N_25401,N_24607);
and U26153 (N_26153,N_25600,N_25035);
or U26154 (N_26154,N_24190,N_24917);
xnor U26155 (N_26155,N_25300,N_24553);
nor U26156 (N_26156,N_24073,N_24112);
xor U26157 (N_26157,N_24606,N_24592);
or U26158 (N_26158,N_24755,N_25197);
xnor U26159 (N_26159,N_25549,N_24679);
nor U26160 (N_26160,N_24181,N_25364);
nor U26161 (N_26161,N_24006,N_24384);
nand U26162 (N_26162,N_25752,N_25346);
nor U26163 (N_26163,N_25352,N_24184);
xnor U26164 (N_26164,N_25464,N_24806);
nor U26165 (N_26165,N_24229,N_25819);
xnor U26166 (N_26166,N_25048,N_25493);
xor U26167 (N_26167,N_25012,N_24963);
or U26168 (N_26168,N_24420,N_25593);
or U26169 (N_26169,N_24035,N_24258);
and U26170 (N_26170,N_25326,N_24082);
nand U26171 (N_26171,N_25440,N_24940);
xor U26172 (N_26172,N_25342,N_25077);
or U26173 (N_26173,N_24842,N_24568);
or U26174 (N_26174,N_25075,N_24655);
and U26175 (N_26175,N_24476,N_25411);
and U26176 (N_26176,N_24537,N_24456);
nand U26177 (N_26177,N_25457,N_24808);
nand U26178 (N_26178,N_25792,N_24115);
nor U26179 (N_26179,N_24954,N_24107);
nor U26180 (N_26180,N_25848,N_25643);
nand U26181 (N_26181,N_25351,N_24359);
and U26182 (N_26182,N_25213,N_25890);
nor U26183 (N_26183,N_25944,N_24462);
nor U26184 (N_26184,N_24833,N_25705);
nor U26185 (N_26185,N_25536,N_24583);
nand U26186 (N_26186,N_24500,N_24226);
and U26187 (N_26187,N_24702,N_25488);
nor U26188 (N_26188,N_25884,N_24109);
nor U26189 (N_26189,N_25332,N_25422);
nand U26190 (N_26190,N_25855,N_24891);
and U26191 (N_26191,N_25544,N_25533);
xor U26192 (N_26192,N_24039,N_25738);
nand U26193 (N_26193,N_25298,N_24021);
nor U26194 (N_26194,N_24804,N_25746);
nand U26195 (N_26195,N_25708,N_24245);
or U26196 (N_26196,N_24993,N_24450);
nand U26197 (N_26197,N_25595,N_25619);
or U26198 (N_26198,N_25455,N_25754);
xnor U26199 (N_26199,N_24243,N_25272);
or U26200 (N_26200,N_24656,N_24988);
and U26201 (N_26201,N_25238,N_25633);
xor U26202 (N_26202,N_24106,N_24925);
xor U26203 (N_26203,N_25313,N_24457);
nand U26204 (N_26204,N_25874,N_24766);
nand U26205 (N_26205,N_25664,N_25623);
or U26206 (N_26206,N_25545,N_24677);
xor U26207 (N_26207,N_25396,N_24196);
and U26208 (N_26208,N_24216,N_25419);
nor U26209 (N_26209,N_24465,N_25940);
nor U26210 (N_26210,N_25501,N_25303);
and U26211 (N_26211,N_24888,N_24850);
and U26212 (N_26212,N_25412,N_24191);
nor U26213 (N_26213,N_25228,N_24091);
nor U26214 (N_26214,N_25484,N_25467);
nor U26215 (N_26215,N_25546,N_24368);
and U26216 (N_26216,N_24904,N_25384);
nor U26217 (N_26217,N_24484,N_24733);
nor U26218 (N_26218,N_24396,N_24999);
nor U26219 (N_26219,N_24414,N_24406);
and U26220 (N_26220,N_24769,N_25808);
xnor U26221 (N_26221,N_25555,N_24002);
and U26222 (N_26222,N_25030,N_24704);
nor U26223 (N_26223,N_24660,N_25003);
xnor U26224 (N_26224,N_25538,N_24311);
nor U26225 (N_26225,N_24700,N_24273);
or U26226 (N_26226,N_24978,N_24459);
and U26227 (N_26227,N_24877,N_24517);
nand U26228 (N_26228,N_24846,N_24518);
and U26229 (N_26229,N_25911,N_24267);
or U26230 (N_26230,N_25284,N_24787);
xnor U26231 (N_26231,N_25800,N_24236);
nand U26232 (N_26232,N_25743,N_24487);
and U26233 (N_26233,N_25523,N_25058);
nand U26234 (N_26234,N_24762,N_24204);
xnor U26235 (N_26235,N_25154,N_24906);
and U26236 (N_26236,N_25214,N_24156);
or U26237 (N_26237,N_24934,N_24281);
or U26238 (N_26238,N_24829,N_25328);
nand U26239 (N_26239,N_25458,N_24036);
nor U26240 (N_26240,N_24514,N_24237);
and U26241 (N_26241,N_24131,N_24280);
nand U26242 (N_26242,N_24316,N_24364);
and U26243 (N_26243,N_24911,N_25158);
nor U26244 (N_26244,N_25993,N_25671);
xor U26245 (N_26245,N_24269,N_24812);
xor U26246 (N_26246,N_25439,N_24047);
or U26247 (N_26247,N_24681,N_24289);
nor U26248 (N_26248,N_25620,N_25469);
nand U26249 (N_26249,N_25253,N_24722);
xor U26250 (N_26250,N_24224,N_25901);
nor U26251 (N_26251,N_24274,N_24964);
or U26252 (N_26252,N_24446,N_25551);
nor U26253 (N_26253,N_25703,N_25842);
nor U26254 (N_26254,N_25915,N_24473);
xnor U26255 (N_26255,N_24659,N_25363);
and U26256 (N_26256,N_25409,N_25797);
xnor U26257 (N_26257,N_25834,N_25644);
and U26258 (N_26258,N_25949,N_25597);
nor U26259 (N_26259,N_25049,N_24775);
or U26260 (N_26260,N_24429,N_25722);
and U26261 (N_26261,N_25485,N_25846);
and U26262 (N_26262,N_24735,N_24576);
and U26263 (N_26263,N_25081,N_24654);
and U26264 (N_26264,N_25001,N_24099);
and U26265 (N_26265,N_24306,N_25498);
nor U26266 (N_26266,N_25938,N_24620);
nor U26267 (N_26267,N_24444,N_25125);
nand U26268 (N_26268,N_25816,N_24969);
or U26269 (N_26269,N_24242,N_24025);
nor U26270 (N_26270,N_25301,N_25027);
nand U26271 (N_26271,N_24522,N_24729);
xor U26272 (N_26272,N_24599,N_24563);
xor U26273 (N_26273,N_25159,N_25937);
nand U26274 (N_26274,N_24747,N_25594);
nor U26275 (N_26275,N_25479,N_24562);
nor U26276 (N_26276,N_25870,N_24096);
xor U26277 (N_26277,N_25341,N_25558);
xnor U26278 (N_26278,N_24122,N_24161);
and U26279 (N_26279,N_25496,N_24665);
and U26280 (N_26280,N_25252,N_25347);
and U26281 (N_26281,N_24283,N_25278);
xor U26282 (N_26282,N_24461,N_24918);
nor U26283 (N_26283,N_25312,N_25651);
nor U26284 (N_26284,N_25330,N_24603);
xor U26285 (N_26285,N_25310,N_24350);
nor U26286 (N_26286,N_25337,N_24981);
nor U26287 (N_26287,N_24356,N_25951);
nand U26288 (N_26288,N_25138,N_25495);
and U26289 (N_26289,N_25957,N_25462);
nand U26290 (N_26290,N_25217,N_24690);
nand U26291 (N_26291,N_24253,N_25851);
xnor U26292 (N_26292,N_24118,N_25866);
or U26293 (N_26293,N_24057,N_24223);
nor U26294 (N_26294,N_25774,N_24613);
and U26295 (N_26295,N_25696,N_24010);
nor U26296 (N_26296,N_25698,N_24859);
or U26297 (N_26297,N_25450,N_24048);
xnor U26298 (N_26298,N_25837,N_24805);
nor U26299 (N_26299,N_25921,N_25408);
or U26300 (N_26300,N_24895,N_25822);
and U26301 (N_26301,N_25489,N_24044);
nor U26302 (N_26302,N_25243,N_24561);
nand U26303 (N_26303,N_25127,N_25031);
nand U26304 (N_26304,N_24541,N_25071);
or U26305 (N_26305,N_25567,N_24028);
xor U26306 (N_26306,N_24867,N_24774);
nand U26307 (N_26307,N_24086,N_25315);
xnor U26308 (N_26308,N_24741,N_24971);
xnor U26309 (N_26309,N_24832,N_24689);
or U26310 (N_26310,N_24116,N_25656);
or U26311 (N_26311,N_24315,N_25707);
or U26312 (N_26312,N_24387,N_25499);
xnor U26313 (N_26313,N_24767,N_24815);
and U26314 (N_26314,N_25416,N_24012);
and U26315 (N_26315,N_24834,N_25490);
nand U26316 (N_26316,N_25066,N_25684);
or U26317 (N_26317,N_25627,N_25483);
and U26318 (N_26318,N_25126,N_25423);
nand U26319 (N_26319,N_24030,N_24638);
and U26320 (N_26320,N_24907,N_24669);
and U26321 (N_26321,N_24866,N_25618);
and U26322 (N_26322,N_24317,N_24171);
nand U26323 (N_26323,N_25274,N_25149);
nor U26324 (N_26324,N_24952,N_25992);
xor U26325 (N_26325,N_25675,N_24830);
and U26326 (N_26326,N_24225,N_24197);
or U26327 (N_26327,N_24174,N_24323);
and U26328 (N_26328,N_24348,N_25581);
xor U26329 (N_26329,N_24045,N_24776);
nor U26330 (N_26330,N_24664,N_25532);
or U26331 (N_26331,N_25964,N_25321);
nand U26332 (N_26332,N_25080,N_24653);
and U26333 (N_26333,N_25520,N_24452);
nand U26334 (N_26334,N_24721,N_25963);
nor U26335 (N_26335,N_24670,N_24912);
or U26336 (N_26336,N_24154,N_24662);
nand U26337 (N_26337,N_24513,N_24329);
nor U26338 (N_26338,N_25270,N_25478);
and U26339 (N_26339,N_24539,N_24909);
or U26340 (N_26340,N_25572,N_25088);
nand U26341 (N_26341,N_24532,N_25570);
xnor U26342 (N_26342,N_25218,N_24786);
nor U26343 (N_26343,N_24784,N_24410);
and U26344 (N_26344,N_25123,N_24615);
nor U26345 (N_26345,N_25706,N_24277);
or U26346 (N_26346,N_24052,N_25099);
nand U26347 (N_26347,N_25198,N_25780);
nor U26348 (N_26348,N_24321,N_25959);
and U26349 (N_26349,N_25124,N_25932);
or U26350 (N_26350,N_25255,N_24865);
xnor U26351 (N_26351,N_24475,N_25515);
xnor U26352 (N_26352,N_24533,N_24011);
xnor U26353 (N_26353,N_24324,N_25592);
and U26354 (N_26354,N_24234,N_25983);
or U26355 (N_26355,N_25108,N_25767);
nor U26356 (N_26356,N_25616,N_25268);
and U26357 (N_26357,N_24478,N_25905);
xor U26358 (N_26358,N_24479,N_25441);
nand U26359 (N_26359,N_25877,N_25266);
xnor U26360 (N_26360,N_24835,N_25199);
nor U26361 (N_26361,N_25475,N_24578);
or U26362 (N_26362,N_24182,N_24439);
nand U26363 (N_26363,N_25550,N_24104);
and U26364 (N_26364,N_24334,N_24419);
and U26365 (N_26365,N_24292,N_24976);
nand U26366 (N_26366,N_25044,N_24764);
and U26367 (N_26367,N_24990,N_25211);
nor U26368 (N_26368,N_25206,N_24038);
and U26369 (N_26369,N_25152,N_25832);
xor U26370 (N_26370,N_25262,N_24300);
nor U26371 (N_26371,N_25234,N_25116);
and U26372 (N_26372,N_24211,N_25795);
and U26373 (N_26373,N_25926,N_24571);
and U26374 (N_26374,N_24825,N_25233);
or U26375 (N_26375,N_25451,N_24719);
xnor U26376 (N_26376,N_24405,N_25535);
xnor U26377 (N_26377,N_25091,N_24732);
or U26378 (N_26378,N_24697,N_24823);
xor U26379 (N_26379,N_24628,N_25854);
nor U26380 (N_26380,N_24612,N_24185);
and U26381 (N_26381,N_25209,N_24477);
or U26382 (N_26382,N_24295,N_25029);
and U26383 (N_26383,N_25148,N_25497);
xnor U26384 (N_26384,N_24203,N_25695);
nand U26385 (N_26385,N_25374,N_25437);
and U26386 (N_26386,N_24481,N_24986);
xor U26387 (N_26387,N_24873,N_25747);
and U26388 (N_26388,N_24515,N_24235);
nor U26389 (N_26389,N_24040,N_24605);
nand U26390 (N_26390,N_25923,N_25429);
xnor U26391 (N_26391,N_25365,N_25751);
or U26392 (N_26392,N_25744,N_24523);
nor U26393 (N_26393,N_24232,N_24297);
nor U26394 (N_26394,N_25192,N_25977);
and U26395 (N_26395,N_25287,N_24159);
and U26396 (N_26396,N_25358,N_24788);
xnor U26397 (N_26397,N_25875,N_25818);
xnor U26398 (N_26398,N_24678,N_24279);
nand U26399 (N_26399,N_25805,N_24133);
xnor U26400 (N_26400,N_24029,N_24007);
xor U26401 (N_26401,N_24157,N_24856);
nor U26402 (N_26402,N_25249,N_24727);
nand U26403 (N_26403,N_25334,N_24868);
and U26404 (N_26404,N_24188,N_24301);
xor U26405 (N_26405,N_25859,N_25840);
nor U26406 (N_26406,N_25607,N_25517);
nand U26407 (N_26407,N_25117,N_25906);
or U26408 (N_26408,N_25171,N_24899);
nor U26409 (N_26409,N_24199,N_24759);
or U26410 (N_26410,N_25529,N_25036);
nor U26411 (N_26411,N_24467,N_25985);
xor U26412 (N_26412,N_24801,N_24395);
nand U26413 (N_26413,N_24424,N_24960);
nand U26414 (N_26414,N_25974,N_24586);
and U26415 (N_26415,N_25543,N_25991);
or U26416 (N_26416,N_24366,N_24585);
nor U26417 (N_26417,N_25087,N_24388);
xor U26418 (N_26418,N_24724,N_25299);
nand U26419 (N_26419,N_25062,N_25433);
or U26420 (N_26420,N_24095,N_25927);
and U26421 (N_26421,N_25547,N_25952);
or U26422 (N_26422,N_24202,N_24975);
xor U26423 (N_26423,N_24031,N_24346);
nand U26424 (N_26424,N_25205,N_24666);
or U26425 (N_26425,N_24627,N_24360);
xnor U26426 (N_26426,N_24996,N_24296);
nand U26427 (N_26427,N_24443,N_24557);
xor U26428 (N_26428,N_24363,N_25111);
nand U26429 (N_26429,N_24144,N_24339);
nand U26430 (N_26430,N_25614,N_24897);
xnor U26431 (N_26431,N_24530,N_24148);
and U26432 (N_26432,N_25021,N_25082);
nand U26433 (N_26433,N_25762,N_24286);
nand U26434 (N_26434,N_24341,N_25646);
nor U26435 (N_26435,N_25858,N_25687);
xor U26436 (N_26436,N_24264,N_25017);
or U26437 (N_26437,N_25518,N_25635);
xor U26438 (N_26438,N_24389,N_24227);
nand U26439 (N_26439,N_24098,N_25608);
xor U26440 (N_26440,N_24371,N_25307);
or U26441 (N_26441,N_24694,N_24087);
and U26442 (N_26442,N_25069,N_24093);
and U26443 (N_26443,N_24838,N_25380);
or U26444 (N_26444,N_24062,N_25702);
nand U26445 (N_26445,N_24195,N_24646);
nor U26446 (N_26446,N_24949,N_25224);
and U26447 (N_26447,N_24590,N_24588);
nand U26448 (N_26448,N_25293,N_25011);
nand U26449 (N_26449,N_24881,N_25460);
nor U26450 (N_26450,N_24889,N_25824);
nand U26451 (N_26451,N_25527,N_24695);
nor U26452 (N_26452,N_25622,N_25059);
nand U26453 (N_26453,N_24059,N_24249);
nor U26454 (N_26454,N_24361,N_24857);
nand U26455 (N_26455,N_24746,N_25184);
nor U26456 (N_26456,N_25606,N_25244);
xnor U26457 (N_26457,N_24139,N_24244);
xnor U26458 (N_26458,N_24018,N_25394);
and U26459 (N_26459,N_24141,N_25132);
nand U26460 (N_26460,N_25917,N_25704);
nor U26461 (N_26461,N_24894,N_24372);
and U26462 (N_26462,N_25871,N_25880);
and U26463 (N_26463,N_25240,N_24454);
or U26464 (N_26464,N_25922,N_24458);
and U26465 (N_26465,N_25865,N_25577);
xnor U26466 (N_26466,N_24421,N_25491);
xnor U26467 (N_26467,N_25878,N_24555);
or U26468 (N_26468,N_25897,N_25955);
nand U26469 (N_26469,N_25986,N_24902);
nor U26470 (N_26470,N_25285,N_24520);
nor U26471 (N_26471,N_25361,N_24432);
and U26472 (N_26472,N_24003,N_25097);
or U26473 (N_26473,N_25482,N_24827);
xnor U26474 (N_26474,N_24703,N_25018);
and U26475 (N_26475,N_24001,N_24063);
or U26476 (N_26476,N_25072,N_24298);
nor U26477 (N_26477,N_24543,N_25560);
nor U26478 (N_26478,N_25603,N_24861);
and U26479 (N_26479,N_24915,N_25809);
nor U26480 (N_26480,N_24821,N_25979);
and U26481 (N_26481,N_24756,N_25246);
and U26482 (N_26482,N_25170,N_24179);
nor U26483 (N_26483,N_24408,N_24575);
nor U26484 (N_26484,N_25220,N_24643);
xor U26485 (N_26485,N_25311,N_24645);
xnor U26486 (N_26486,N_24598,N_24594);
or U26487 (N_26487,N_25789,N_24246);
and U26488 (N_26488,N_24079,N_25305);
or U26489 (N_26489,N_25360,N_25324);
nor U26490 (N_26490,N_24673,N_24065);
nor U26491 (N_26491,N_24092,N_25665);
nand U26492 (N_26492,N_24340,N_25898);
and U26493 (N_26493,N_24170,N_25987);
xor U26494 (N_26494,N_24075,N_24709);
xnor U26495 (N_26495,N_25424,N_25613);
xnor U26496 (N_26496,N_25186,N_25645);
nand U26497 (N_26497,N_25005,N_25250);
xor U26498 (N_26498,N_24053,N_24228);
nand U26499 (N_26499,N_25999,N_25850);
nor U26500 (N_26500,N_24305,N_24742);
or U26501 (N_26501,N_25344,N_25686);
nor U26502 (N_26502,N_24207,N_25338);
nor U26503 (N_26503,N_25325,N_24840);
nor U26504 (N_26504,N_24847,N_24337);
nor U26505 (N_26505,N_25449,N_24460);
nand U26506 (N_26506,N_24056,N_24544);
nor U26507 (N_26507,N_24401,N_25956);
nand U26508 (N_26508,N_24119,N_24824);
nor U26509 (N_26509,N_24939,N_24442);
nand U26510 (N_26510,N_24290,N_24134);
nor U26511 (N_26511,N_25174,N_24331);
nand U26512 (N_26512,N_24885,N_24166);
or U26513 (N_26513,N_24418,N_25813);
nand U26514 (N_26514,N_24998,N_24597);
xor U26515 (N_26515,N_25759,N_24307);
and U26516 (N_26516,N_24577,N_25694);
or U26517 (N_26517,N_25978,N_25008);
and U26518 (N_26518,N_24146,N_25026);
and U26519 (N_26519,N_24125,N_25207);
nor U26520 (N_26520,N_25172,N_25076);
xnor U26521 (N_26521,N_25892,N_25265);
xnor U26522 (N_26522,N_25112,N_24545);
nor U26523 (N_26523,N_25864,N_24777);
xnor U26524 (N_26524,N_25887,N_25755);
nand U26525 (N_26525,N_24916,N_25678);
nor U26526 (N_26526,N_24609,N_25176);
nor U26527 (N_26527,N_25920,N_25914);
or U26528 (N_26528,N_25389,N_24221);
xor U26529 (N_26529,N_25227,N_25379);
or U26530 (N_26530,N_24750,N_24649);
nor U26531 (N_26531,N_24535,N_25862);
nand U26532 (N_26532,N_24240,N_25007);
xnor U26533 (N_26533,N_24037,N_25195);
xor U26534 (N_26534,N_24081,N_24282);
nor U26535 (N_26535,N_25975,N_24275);
xnor U26536 (N_26536,N_25356,N_25750);
or U26537 (N_26537,N_24569,N_25223);
nor U26538 (N_26538,N_24914,N_24950);
or U26539 (N_26539,N_24113,N_24754);
or U26540 (N_26540,N_24186,N_24547);
and U26541 (N_26541,N_24077,N_25579);
and U26542 (N_26542,N_24958,N_25637);
nor U26543 (N_26543,N_25388,N_24344);
nand U26544 (N_26544,N_24494,N_25624);
or U26545 (N_26545,N_24320,N_25273);
nand U26546 (N_26546,N_25084,N_24138);
nor U26547 (N_26547,N_24076,N_24309);
and U26548 (N_26548,N_24072,N_25131);
nand U26549 (N_26549,N_25225,N_24169);
xor U26550 (N_26550,N_25390,N_24977);
or U26551 (N_26551,N_24415,N_25133);
nand U26552 (N_26552,N_24778,N_25110);
xor U26553 (N_26553,N_25510,N_24693);
or U26554 (N_26554,N_25586,N_24658);
nand U26555 (N_26555,N_25398,N_25041);
xor U26556 (N_26556,N_25241,N_25621);
nand U26557 (N_26557,N_24844,N_25784);
xor U26558 (N_26558,N_24466,N_24241);
xnor U26559 (N_26559,N_24353,N_25766);
nor U26560 (N_26560,N_24200,N_24430);
xor U26561 (N_26561,N_25802,N_24610);
xor U26562 (N_26562,N_25203,N_24760);
nand U26563 (N_26563,N_25004,N_25827);
xnor U26564 (N_26564,N_24123,N_25292);
nand U26565 (N_26565,N_24641,N_25202);
or U26566 (N_26566,N_25630,N_25668);
xor U26567 (N_26567,N_24651,N_25229);
xor U26568 (N_26568,N_24254,N_25718);
nor U26569 (N_26569,N_25793,N_24020);
and U26570 (N_26570,N_25584,N_25814);
xor U26571 (N_26571,N_25836,N_24927);
nor U26572 (N_26572,N_24579,N_25430);
xnor U26573 (N_26573,N_24682,N_24008);
xnor U26574 (N_26574,N_25256,N_25573);
nand U26575 (N_26575,N_24126,N_24362);
xor U26576 (N_26576,N_25688,N_24966);
nor U26577 (N_26577,N_25935,N_24470);
and U26578 (N_26578,N_24392,N_25304);
nand U26579 (N_26579,N_25655,N_24512);
and U26580 (N_26580,N_25336,N_25283);
xnor U26581 (N_26581,N_24941,N_24097);
or U26582 (N_26582,N_25542,N_25051);
or U26583 (N_26583,N_25902,N_25745);
nand U26584 (N_26584,N_24164,N_25894);
and U26585 (N_26585,N_24818,N_25037);
or U26586 (N_26586,N_25296,N_24771);
or U26587 (N_26587,N_25130,N_24896);
nand U26588 (N_26588,N_25820,N_24900);
xnor U26589 (N_26589,N_25119,N_25322);
and U26590 (N_26590,N_25314,N_25839);
and U26591 (N_26591,N_25355,N_25990);
nor U26592 (N_26592,N_24390,N_24453);
xor U26593 (N_26593,N_24303,N_25431);
xnor U26594 (N_26594,N_25562,N_24480);
and U26595 (N_26595,N_24205,N_25677);
or U26596 (N_26596,N_24632,N_25428);
or U26597 (N_26597,N_24822,N_25640);
and U26598 (N_26598,N_25254,N_24449);
nor U26599 (N_26599,N_24644,N_24299);
nand U26600 (N_26600,N_24631,N_24230);
nor U26601 (N_26601,N_25930,N_25359);
or U26602 (N_26602,N_24042,N_24400);
or U26603 (N_26603,N_24728,N_24209);
and U26604 (N_26604,N_24193,N_25447);
xor U26605 (N_26605,N_24074,N_25631);
and U26606 (N_26606,N_24187,N_25960);
or U26607 (N_26607,N_25239,N_24625);
nor U26608 (N_26608,N_25306,N_24635);
nor U26609 (N_26609,N_25697,N_25068);
and U26610 (N_26610,N_25873,N_25817);
or U26611 (N_26611,N_24369,N_24935);
and U26612 (N_26612,N_25845,N_25281);
or U26613 (N_26613,N_24504,N_25934);
xnor U26614 (N_26614,N_25492,N_25969);
nand U26615 (N_26615,N_25025,N_25599);
nor U26616 (N_26616,N_25267,N_25729);
xnor U26617 (N_26617,N_25654,N_25525);
nand U26618 (N_26618,N_25556,N_25590);
nand U26619 (N_26619,N_25967,N_25672);
nand U26620 (N_26620,N_24278,N_24293);
nor U26621 (N_26621,N_24474,N_25370);
nand U26622 (N_26622,N_25775,N_25868);
and U26623 (N_26623,N_24854,N_24026);
nor U26624 (N_26624,N_25610,N_25602);
xnor U26625 (N_26625,N_24936,N_24218);
and U26626 (N_26626,N_25382,N_25055);
or U26627 (N_26627,N_25442,N_24373);
xnor U26628 (N_26628,N_24668,N_24618);
nand U26629 (N_26629,N_24745,N_25748);
nand U26630 (N_26630,N_24849,N_24370);
and U26631 (N_26631,N_24860,N_24375);
and U26632 (N_26632,N_25166,N_24050);
nand U26633 (N_26633,N_25271,N_25933);
nand U26634 (N_26634,N_25730,N_24593);
xnor U26635 (N_26635,N_25317,N_25724);
or U26636 (N_26636,N_25950,N_24469);
nor U26637 (N_26637,N_24114,N_24382);
or U26638 (N_26638,N_24422,N_25772);
nor U26639 (N_26639,N_25155,N_24951);
or U26640 (N_26640,N_25378,N_24855);
xnor U26641 (N_26641,N_25245,N_24738);
and U26642 (N_26642,N_25652,N_24974);
or U26643 (N_26643,N_25961,N_25182);
nor U26644 (N_26644,N_25371,N_25288);
nand U26645 (N_26645,N_25931,N_24411);
or U26646 (N_26646,N_24061,N_24505);
or U26647 (N_26647,N_24455,N_24714);
nand U26648 (N_26648,N_25727,N_24101);
and U26649 (N_26649,N_24995,N_24720);
nor U26650 (N_26650,N_24765,N_24503);
or U26651 (N_26651,N_25580,N_25663);
and U26652 (N_26652,N_25410,N_25596);
nand U26653 (N_26653,N_24884,N_24143);
or U26654 (N_26654,N_24616,N_25200);
and U26655 (N_26655,N_25539,N_24351);
or U26656 (N_26656,N_25385,N_25988);
and U26657 (N_26657,N_25989,N_25187);
and U26658 (N_26658,N_24781,N_25177);
nand U26659 (N_26659,N_24447,N_24251);
nand U26660 (N_26660,N_24365,N_24013);
and U26661 (N_26661,N_25786,N_25377);
and U26662 (N_26662,N_25830,N_25070);
xor U26663 (N_26663,N_25526,N_24117);
xnor U26664 (N_26664,N_24711,N_25835);
nand U26665 (N_26665,N_25582,N_24102);
nand U26666 (N_26666,N_25067,N_24060);
and U26667 (N_26667,N_24397,N_24206);
xor U26668 (N_26668,N_25144,N_25373);
nand U26669 (N_26669,N_25737,N_24066);
nor U26670 (N_26670,N_24623,N_24496);
nand U26671 (N_26671,N_24084,N_25002);
and U26672 (N_26672,N_24582,N_24094);
or U26673 (N_26673,N_24548,N_25741);
nand U26674 (N_26674,N_24717,N_24772);
nor U26675 (N_26675,N_24875,N_25316);
nor U26676 (N_26676,N_25946,N_24549);
nor U26677 (N_26677,N_24250,N_25653);
xor U26678 (N_26678,N_25598,N_24426);
nor U26679 (N_26679,N_24252,N_25405);
and U26680 (N_26680,N_24431,N_25095);
or U26681 (N_26681,N_24611,N_25046);
nor U26682 (N_26682,N_25208,N_25466);
or U26683 (N_26683,N_25487,N_25648);
nand U26684 (N_26684,N_25289,N_25764);
xnor U26685 (N_26685,N_25962,N_24796);
xor U26686 (N_26686,N_25448,N_25641);
and U26687 (N_26687,N_24740,N_24790);
nand U26688 (N_26688,N_25601,N_24845);
and U26689 (N_26689,N_25335,N_24428);
xnor U26690 (N_26690,N_24308,N_25153);
and U26691 (N_26691,N_24559,N_25251);
xor U26692 (N_26692,N_24879,N_25716);
xor U26693 (N_26693,N_24239,N_25052);
or U26694 (N_26694,N_25503,N_24342);
nand U26695 (N_26695,N_24595,N_25391);
or U26696 (N_26696,N_24078,N_24831);
nor U26697 (N_26697,N_25115,N_25395);
nor U26698 (N_26698,N_25998,N_25247);
nor U26699 (N_26699,N_24962,N_25168);
nand U26700 (N_26700,N_25861,N_24024);
nor U26701 (N_26701,N_25333,N_25454);
nor U26702 (N_26702,N_24634,N_25522);
xnor U26703 (N_26703,N_25806,N_25844);
or U26704 (N_26704,N_24744,N_24811);
nor U26705 (N_26705,N_25444,N_25972);
and U26706 (N_26706,N_25279,N_25386);
and U26707 (N_26707,N_25717,N_24176);
nand U26708 (N_26708,N_24928,N_25700);
or U26709 (N_26709,N_24255,N_24922);
and U26710 (N_26710,N_25040,N_25565);
or U26711 (N_26711,N_24270,N_25516);
nand U26712 (N_26712,N_24893,N_24019);
nand U26713 (N_26713,N_25900,N_25142);
xor U26714 (N_26714,N_24908,N_25628);
xor U26715 (N_26715,N_24570,N_24265);
nor U26716 (N_26716,N_24874,N_24581);
and U26717 (N_26717,N_24041,N_24268);
and U26718 (N_26718,N_25826,N_25219);
xnor U26719 (N_26719,N_25569,N_25000);
nand U26720 (N_26720,N_25470,N_25323);
and U26721 (N_26721,N_25735,N_24937);
xor U26722 (N_26722,N_24546,N_24183);
nand U26723 (N_26723,N_24173,N_24502);
nand U26724 (N_26724,N_24979,N_24043);
and U26725 (N_26725,N_24493,N_24734);
xnor U26726 (N_26726,N_25147,N_25657);
nor U26727 (N_26727,N_24793,N_25981);
and U26728 (N_26728,N_25984,N_24445);
nand U26729 (N_26729,N_25381,N_24448);
or U26730 (N_26730,N_25397,N_25291);
nand U26731 (N_26731,N_24572,N_24302);
xnor U26732 (N_26732,N_25102,N_25366);
nand U26733 (N_26733,N_24991,N_25375);
and U26734 (N_26734,N_24180,N_25277);
nand U26735 (N_26735,N_25340,N_24177);
xnor U26736 (N_26736,N_25929,N_24723);
xnor U26737 (N_26737,N_24743,N_25699);
xnor U26738 (N_26738,N_24887,N_24560);
or U26739 (N_26739,N_24276,N_25505);
nor U26740 (N_26740,N_24000,N_24322);
and U26741 (N_26741,N_25494,N_25885);
nand U26742 (N_26742,N_25015,N_25114);
or U26743 (N_26743,N_25020,N_24674);
or U26744 (N_26744,N_25023,N_25715);
nand U26745 (N_26745,N_24347,N_25642);
and U26746 (N_26746,N_24155,N_25553);
nand U26747 (N_26747,N_24049,N_24386);
and U26748 (N_26748,N_24985,N_25327);
nand U26749 (N_26749,N_25636,N_25427);
or U26750 (N_26750,N_24325,N_25673);
or U26751 (N_26751,N_25079,N_24055);
and U26752 (N_26752,N_25258,N_24587);
nand U26753 (N_26753,N_24809,N_24972);
or U26754 (N_26754,N_25402,N_24980);
nor U26755 (N_26755,N_24486,N_25353);
and U26756 (N_26756,N_25736,N_24149);
and U26757 (N_26757,N_25828,N_24058);
nor U26758 (N_26758,N_24920,N_24464);
and U26759 (N_26759,N_24015,N_25354);
or U26760 (N_26760,N_24876,N_24033);
nor U26761 (N_26761,N_24946,N_25434);
or U26762 (N_26762,N_25139,N_25966);
or U26763 (N_26763,N_24404,N_24614);
and U26764 (N_26764,N_24198,N_24017);
xnor U26765 (N_26765,N_24982,N_25073);
or U26766 (N_26766,N_24943,N_25039);
or U26767 (N_26767,N_25083,N_24526);
nand U26768 (N_26768,N_24650,N_25383);
nor U26769 (N_26769,N_24938,N_24870);
xnor U26770 (N_26770,N_24820,N_25626);
and U26771 (N_26771,N_25276,N_24892);
xnor U26772 (N_26772,N_25463,N_25413);
and U26773 (N_26773,N_24698,N_24550);
nand U26774 (N_26774,N_25104,N_25275);
and U26775 (N_26775,N_24519,N_24409);
xor U26776 (N_26776,N_25290,N_25103);
nand U26777 (N_26777,N_25297,N_25106);
or U26778 (N_26778,N_25308,N_24129);
and U26779 (N_26779,N_24120,N_25609);
nor U26780 (N_26780,N_25857,N_25376);
xor U26781 (N_26781,N_24761,N_24524);
or U26782 (N_26782,N_24492,N_25528);
nand U26783 (N_26783,N_25810,N_24374);
nand U26784 (N_26784,N_24438,N_25847);
or U26785 (N_26785,N_25958,N_25345);
and U26786 (N_26786,N_24752,N_25183);
nor U26787 (N_26787,N_25650,N_25605);
and U26788 (N_26788,N_25888,N_24871);
and U26789 (N_26789,N_24314,N_25575);
or U26790 (N_26790,N_24497,N_25712);
nand U26791 (N_26791,N_25530,N_24338);
or U26792 (N_26792,N_25028,N_24926);
or U26793 (N_26793,N_25876,N_25471);
nor U26794 (N_26794,N_25456,N_25807);
nand U26795 (N_26795,N_25173,N_25191);
and U26796 (N_26796,N_24247,N_24511);
xor U26797 (N_26797,N_24932,N_24540);
xor U26798 (N_26798,N_25118,N_24412);
nand U26799 (N_26799,N_24730,N_24521);
xnor U26800 (N_26800,N_25179,N_25421);
nand U26801 (N_26801,N_24256,N_25997);
nand U26802 (N_26802,N_24441,N_24947);
or U26803 (N_26803,N_25588,N_24083);
and U26804 (N_26804,N_24886,N_25404);
xor U26805 (N_26805,N_24508,N_25563);
nand U26806 (N_26806,N_25728,N_24686);
xnor U26807 (N_26807,N_25968,N_25928);
nand U26808 (N_26808,N_24843,N_25889);
nor U26809 (N_26809,N_25032,N_25134);
and U26810 (N_26810,N_25180,N_24014);
and U26811 (N_26811,N_25339,N_25831);
xor U26812 (N_26812,N_25216,N_24813);
nand U26813 (N_26813,N_25612,N_25013);
xor U26814 (N_26814,N_25939,N_25521);
or U26815 (N_26815,N_25446,N_25891);
xor U26816 (N_26816,N_24715,N_24574);
nor U26817 (N_26817,N_25033,N_24005);
or U26818 (N_26818,N_24600,N_25970);
nor U26819 (N_26819,N_24071,N_24491);
or U26820 (N_26820,N_25604,N_25122);
nor U26821 (N_26821,N_24433,N_25982);
and U26822 (N_26822,N_24498,N_24836);
nand U26823 (N_26823,N_25415,N_24699);
nand U26824 (N_26824,N_24795,N_25092);
and U26825 (N_26825,N_24345,N_25480);
nand U26826 (N_26826,N_25667,N_25006);
nand U26827 (N_26827,N_24262,N_25591);
nor U26828 (N_26828,N_24580,N_25879);
or U26829 (N_26829,N_25426,N_25849);
nor U26830 (N_26830,N_25825,N_25942);
and U26831 (N_26831,N_25740,N_25617);
and U26832 (N_26832,N_24529,N_24817);
or U26833 (N_26833,N_24748,N_25661);
nand U26834 (N_26834,N_24989,N_25368);
or U26835 (N_26835,N_24046,N_24378);
and U26836 (N_26836,N_25534,N_25105);
xnor U26837 (N_26837,N_24630,N_24863);
and U26838 (N_26838,N_25061,N_24482);
xor U26839 (N_26839,N_25204,N_25723);
nand U26840 (N_26840,N_24393,N_25259);
or U26841 (N_26841,N_25843,N_24330);
or U26842 (N_26842,N_25823,N_24103);
xnor U26843 (N_26843,N_25679,N_25742);
nor U26844 (N_26844,N_24882,N_25443);
nor U26845 (N_26845,N_25683,N_24785);
xnor U26846 (N_26846,N_25733,N_25167);
xnor U26847 (N_26847,N_25732,N_25996);
nor U26848 (N_26848,N_24413,N_25100);
nor U26849 (N_26849,N_24692,N_24128);
or U26850 (N_26850,N_25863,N_25954);
or U26851 (N_26851,N_25531,N_24757);
or U26852 (N_26852,N_24219,N_25348);
or U26853 (N_26853,N_24883,N_24488);
xnor U26854 (N_26854,N_25856,N_25350);
nand U26855 (N_26855,N_25803,N_25578);
or U26856 (N_26856,N_25472,N_25557);
xor U26857 (N_26857,N_25145,N_25294);
nand U26858 (N_26858,N_24090,N_24192);
nor U26859 (N_26859,N_24332,N_24385);
xnor U26860 (N_26860,N_24349,N_25625);
or U26861 (N_26861,N_25175,N_25896);
nor U26862 (N_26862,N_24381,N_24647);
nor U26863 (N_26863,N_25393,N_25681);
xor U26864 (N_26864,N_24687,N_24507);
xnor U26865 (N_26865,N_25833,N_24528);
or U26866 (N_26866,N_25585,N_24601);
nand U26867 (N_26867,N_25502,N_24636);
nand U26868 (N_26868,N_25010,N_24343);
nor U26869 (N_26869,N_25445,N_25634);
xor U26870 (N_26870,N_25096,N_24648);
nand U26871 (N_26871,N_24100,N_24970);
and U26872 (N_26872,N_25976,N_25947);
xor U26873 (N_26873,N_24994,N_25024);
xnor U26874 (N_26874,N_25511,N_24248);
nor U26875 (N_26875,N_24701,N_24051);
nand U26876 (N_26876,N_25016,N_24773);
nand U26877 (N_26877,N_24696,N_24127);
nor U26878 (N_26878,N_25392,N_25196);
and U26879 (N_26879,N_24259,N_24136);
nand U26880 (N_26880,N_25886,N_25089);
and U26881 (N_26881,N_24621,N_25632);
nor U26882 (N_26882,N_25236,N_24260);
xnor U26883 (N_26883,N_24130,N_24142);
and U26884 (N_26884,N_25047,N_25971);
and U26885 (N_26885,N_24398,N_24987);
and U26886 (N_26886,N_25452,N_24069);
nand U26887 (N_26887,N_24848,N_24333);
or U26888 (N_26888,N_24713,N_24903);
or U26889 (N_26889,N_25559,N_24089);
nor U26890 (N_26890,N_25161,N_25760);
and U26891 (N_26891,N_25136,N_24427);
nand U26892 (N_26892,N_24263,N_24864);
nand U26893 (N_26893,N_25666,N_24933);
nor U26894 (N_26894,N_24358,N_24783);
and U26895 (N_26895,N_25163,N_24794);
nor U26896 (N_26896,N_24841,N_24022);
nor U26897 (N_26897,N_24680,N_25811);
xor U26898 (N_26898,N_24789,N_25821);
xor U26899 (N_26899,N_24168,N_24212);
and U26900 (N_26900,N_25042,N_25726);
nand U26901 (N_26901,N_25519,N_24633);
nor U26902 (N_26902,N_24731,N_24210);
xor U26903 (N_26903,N_25190,N_25109);
nand U26904 (N_26904,N_25053,N_24285);
nand U26905 (N_26905,N_25776,N_24391);
or U26906 (N_26906,N_24640,N_25771);
and U26907 (N_26907,N_24604,N_24556);
and U26908 (N_26908,N_25436,N_24310);
or U26909 (N_26909,N_25941,N_25564);
or U26910 (N_26910,N_24725,N_24780);
or U26911 (N_26911,N_25568,N_25893);
xnor U26912 (N_26912,N_25761,N_25162);
xor U26913 (N_26913,N_24542,N_24853);
nand U26914 (N_26914,N_25320,N_25140);
and U26915 (N_26915,N_24671,N_25085);
nand U26916 (N_26916,N_24080,N_25181);
or U26917 (N_26917,N_25086,N_25286);
and U26918 (N_26918,N_24009,N_24967);
xor U26919 (N_26919,N_25215,N_24684);
or U26920 (N_26920,N_25924,N_24483);
nor U26921 (N_26921,N_24973,N_24407);
nor U26922 (N_26922,N_24377,N_25537);
and U26923 (N_26923,N_24797,N_24923);
nand U26924 (N_26924,N_25261,N_25948);
and U26925 (N_26925,N_24565,N_25343);
nor U26926 (N_26926,N_24527,N_25367);
or U26927 (N_26927,N_24807,N_25725);
or U26928 (N_26928,N_24145,N_25514);
xnor U26929 (N_26929,N_25649,N_24436);
nand U26930 (N_26930,N_24257,N_24890);
xnor U26931 (N_26931,N_25269,N_25157);
and U26932 (N_26932,N_24536,N_24108);
xnor U26933 (N_26933,N_24379,N_24802);
nor U26934 (N_26934,N_24088,N_25435);
and U26935 (N_26935,N_25719,N_25647);
nand U26936 (N_26936,N_25101,N_25756);
or U26937 (N_26937,N_25369,N_24931);
nor U26938 (N_26938,N_24898,N_25749);
xnor U26939 (N_26939,N_24153,N_25785);
and U26940 (N_26940,N_24591,N_24506);
xnor U26941 (N_26941,N_25659,N_25925);
xor U26942 (N_26942,N_25403,N_24158);
or U26943 (N_26943,N_25014,N_25583);
nand U26944 (N_26944,N_25045,N_24215);
and U26945 (N_26945,N_24791,N_25867);
and U26946 (N_26946,N_25129,N_25414);
and U26947 (N_26947,N_24238,N_24110);
xnor U26948 (N_26948,N_25128,N_25734);
nor U26949 (N_26949,N_24214,N_25222);
nor U26950 (N_26950,N_25295,N_24233);
nand U26951 (N_26951,N_25782,N_24435);
xnor U26952 (N_26952,N_25711,N_24924);
and U26953 (N_26953,N_24739,N_25676);
or U26954 (N_26954,N_24027,N_25639);
xnor U26955 (N_26955,N_25552,N_24837);
nor U26956 (N_26956,N_24327,N_25372);
xnor U26957 (N_26957,N_24261,N_24064);
xor U26958 (N_26958,N_25883,N_24622);
xor U26959 (N_26959,N_24942,N_25629);
nand U26960 (N_26960,N_24688,N_25019);
or U26961 (N_26961,N_25329,N_24712);
nand U26962 (N_26962,N_24905,N_25150);
nor U26963 (N_26963,N_25524,N_24828);
and U26964 (N_26964,N_24953,N_24417);
xor U26965 (N_26965,N_25078,N_24770);
nor U26966 (N_26966,N_24054,N_24423);
or U26967 (N_26967,N_24810,N_25400);
and U26968 (N_26968,N_25465,N_25120);
and U26969 (N_26969,N_25980,N_24910);
and U26970 (N_26970,N_25309,N_24538);
and U26971 (N_26971,N_25571,N_25387);
nand U26972 (N_26972,N_25193,N_25763);
or U26973 (N_26973,N_24067,N_25063);
or U26974 (N_26974,N_24763,N_25189);
nand U26975 (N_26975,N_24437,N_24826);
or U26976 (N_26976,N_24357,N_25757);
xnor U26977 (N_26977,N_25438,N_25798);
nor U26978 (N_26978,N_25043,N_24525);
xnor U26979 (N_26979,N_24573,N_24394);
or U26980 (N_26980,N_25576,N_25038);
and U26981 (N_26981,N_24758,N_25912);
or U26982 (N_26982,N_25473,N_25164);
nor U26983 (N_26983,N_25056,N_25801);
and U26984 (N_26984,N_25226,N_24367);
nand U26985 (N_26985,N_25611,N_24132);
xnor U26986 (N_26986,N_24004,N_25113);
xor U26987 (N_26987,N_25994,N_25720);
or U26988 (N_26988,N_24564,N_25574);
and U26989 (N_26989,N_24085,N_25057);
and U26990 (N_26990,N_25918,N_24959);
and U26991 (N_26991,N_24984,N_25230);
nand U26992 (N_26992,N_25662,N_24554);
xnor U26993 (N_26993,N_24016,N_25872);
nor U26994 (N_26994,N_24956,N_24172);
xor U26995 (N_26995,N_24968,N_25349);
or U26996 (N_26996,N_24463,N_24434);
nand U26997 (N_26997,N_24608,N_25185);
xnor U26998 (N_26998,N_24499,N_25232);
nor U26999 (N_26999,N_25852,N_25788);
nand U27000 (N_27000,N_25973,N_24300);
xnor U27001 (N_27001,N_24213,N_24995);
nor U27002 (N_27002,N_24301,N_25462);
nor U27003 (N_27003,N_24714,N_24960);
nor U27004 (N_27004,N_25627,N_25906);
and U27005 (N_27005,N_24436,N_24117);
nor U27006 (N_27006,N_24977,N_24069);
or U27007 (N_27007,N_25822,N_25566);
or U27008 (N_27008,N_24228,N_24563);
xnor U27009 (N_27009,N_25184,N_24697);
or U27010 (N_27010,N_25042,N_25205);
and U27011 (N_27011,N_24888,N_24444);
nor U27012 (N_27012,N_24674,N_25609);
xor U27013 (N_27013,N_24286,N_25321);
nor U27014 (N_27014,N_24675,N_24505);
or U27015 (N_27015,N_25818,N_24570);
or U27016 (N_27016,N_25035,N_25571);
xnor U27017 (N_27017,N_25770,N_24810);
nand U27018 (N_27018,N_25165,N_25013);
xor U27019 (N_27019,N_25263,N_24489);
and U27020 (N_27020,N_25670,N_25925);
nor U27021 (N_27021,N_25114,N_24195);
and U27022 (N_27022,N_25865,N_25294);
xor U27023 (N_27023,N_25875,N_24476);
or U27024 (N_27024,N_24559,N_25946);
or U27025 (N_27025,N_25700,N_24624);
and U27026 (N_27026,N_24076,N_25674);
nand U27027 (N_27027,N_25723,N_25208);
nor U27028 (N_27028,N_24473,N_25026);
nor U27029 (N_27029,N_25552,N_24733);
nand U27030 (N_27030,N_25730,N_24648);
and U27031 (N_27031,N_24464,N_25744);
or U27032 (N_27032,N_24508,N_25228);
and U27033 (N_27033,N_24553,N_24047);
or U27034 (N_27034,N_24358,N_24672);
nor U27035 (N_27035,N_25637,N_24770);
nor U27036 (N_27036,N_24119,N_25297);
nor U27037 (N_27037,N_25608,N_25429);
xnor U27038 (N_27038,N_25412,N_25268);
xnor U27039 (N_27039,N_24370,N_24571);
nor U27040 (N_27040,N_25926,N_24394);
xnor U27041 (N_27041,N_25428,N_24477);
or U27042 (N_27042,N_24983,N_25534);
nor U27043 (N_27043,N_24856,N_25441);
xnor U27044 (N_27044,N_25871,N_24129);
nand U27045 (N_27045,N_24889,N_24146);
and U27046 (N_27046,N_24138,N_25403);
nand U27047 (N_27047,N_24806,N_24550);
and U27048 (N_27048,N_25948,N_24072);
nand U27049 (N_27049,N_25940,N_25158);
nand U27050 (N_27050,N_24728,N_25868);
or U27051 (N_27051,N_24923,N_24122);
nor U27052 (N_27052,N_25981,N_25700);
nand U27053 (N_27053,N_25141,N_25549);
and U27054 (N_27054,N_25168,N_24899);
xor U27055 (N_27055,N_25157,N_24419);
xor U27056 (N_27056,N_24612,N_25790);
or U27057 (N_27057,N_25392,N_25825);
nor U27058 (N_27058,N_25598,N_25941);
nor U27059 (N_27059,N_24075,N_25734);
xnor U27060 (N_27060,N_25407,N_25111);
and U27061 (N_27061,N_24821,N_24397);
nor U27062 (N_27062,N_24669,N_24347);
nand U27063 (N_27063,N_24383,N_24356);
nand U27064 (N_27064,N_24545,N_24788);
nand U27065 (N_27065,N_24923,N_25978);
or U27066 (N_27066,N_25997,N_25251);
or U27067 (N_27067,N_24152,N_24702);
and U27068 (N_27068,N_25799,N_24760);
nor U27069 (N_27069,N_24813,N_24805);
nor U27070 (N_27070,N_25757,N_25841);
and U27071 (N_27071,N_24562,N_25392);
xor U27072 (N_27072,N_24459,N_25851);
nor U27073 (N_27073,N_24270,N_25948);
and U27074 (N_27074,N_24702,N_24912);
and U27075 (N_27075,N_24341,N_24854);
and U27076 (N_27076,N_24610,N_25277);
or U27077 (N_27077,N_24775,N_24153);
or U27078 (N_27078,N_24405,N_25415);
and U27079 (N_27079,N_25366,N_24959);
xor U27080 (N_27080,N_25863,N_25667);
nand U27081 (N_27081,N_24364,N_24163);
xnor U27082 (N_27082,N_25314,N_25290);
nand U27083 (N_27083,N_24558,N_25718);
nand U27084 (N_27084,N_25843,N_24263);
nor U27085 (N_27085,N_25815,N_25283);
nand U27086 (N_27086,N_25976,N_25410);
nand U27087 (N_27087,N_25911,N_25438);
or U27088 (N_27088,N_24169,N_24666);
nor U27089 (N_27089,N_25689,N_24193);
and U27090 (N_27090,N_25917,N_24441);
xnor U27091 (N_27091,N_25648,N_25952);
nor U27092 (N_27092,N_25006,N_24517);
xor U27093 (N_27093,N_25263,N_24148);
xnor U27094 (N_27094,N_24856,N_24096);
or U27095 (N_27095,N_24204,N_24572);
nor U27096 (N_27096,N_24090,N_25723);
xor U27097 (N_27097,N_25262,N_25791);
and U27098 (N_27098,N_24732,N_25581);
and U27099 (N_27099,N_24130,N_24104);
nor U27100 (N_27100,N_25174,N_25041);
nand U27101 (N_27101,N_25382,N_25986);
and U27102 (N_27102,N_25791,N_24355);
nor U27103 (N_27103,N_24260,N_24869);
xor U27104 (N_27104,N_25031,N_25012);
nor U27105 (N_27105,N_24996,N_25399);
xor U27106 (N_27106,N_25676,N_24530);
or U27107 (N_27107,N_24720,N_24051);
and U27108 (N_27108,N_24327,N_24330);
xnor U27109 (N_27109,N_25324,N_25044);
xor U27110 (N_27110,N_25446,N_24625);
and U27111 (N_27111,N_25834,N_24465);
xnor U27112 (N_27112,N_25569,N_24891);
and U27113 (N_27113,N_25544,N_24025);
and U27114 (N_27114,N_24999,N_25752);
and U27115 (N_27115,N_25691,N_24757);
nor U27116 (N_27116,N_24497,N_24625);
xnor U27117 (N_27117,N_25682,N_24645);
xnor U27118 (N_27118,N_25224,N_25767);
or U27119 (N_27119,N_24073,N_24661);
or U27120 (N_27120,N_25103,N_25073);
and U27121 (N_27121,N_24585,N_25794);
nand U27122 (N_27122,N_24576,N_25242);
and U27123 (N_27123,N_24960,N_24297);
nand U27124 (N_27124,N_25248,N_25894);
and U27125 (N_27125,N_24887,N_24073);
and U27126 (N_27126,N_24048,N_24879);
xnor U27127 (N_27127,N_25159,N_25636);
nor U27128 (N_27128,N_24858,N_24361);
or U27129 (N_27129,N_25680,N_24069);
and U27130 (N_27130,N_25073,N_25586);
nor U27131 (N_27131,N_24887,N_24251);
xnor U27132 (N_27132,N_25022,N_25957);
or U27133 (N_27133,N_25836,N_25958);
nand U27134 (N_27134,N_25467,N_25794);
or U27135 (N_27135,N_24726,N_25464);
xor U27136 (N_27136,N_24305,N_24609);
xnor U27137 (N_27137,N_25094,N_24958);
and U27138 (N_27138,N_24054,N_25699);
and U27139 (N_27139,N_24001,N_24689);
xnor U27140 (N_27140,N_24743,N_24101);
nand U27141 (N_27141,N_24640,N_25456);
or U27142 (N_27142,N_24522,N_24909);
xor U27143 (N_27143,N_24723,N_24175);
and U27144 (N_27144,N_25404,N_25304);
xnor U27145 (N_27145,N_24035,N_24037);
and U27146 (N_27146,N_24618,N_25974);
nor U27147 (N_27147,N_24673,N_25673);
and U27148 (N_27148,N_24888,N_25115);
and U27149 (N_27149,N_24577,N_24304);
nand U27150 (N_27150,N_25359,N_25025);
or U27151 (N_27151,N_25035,N_25299);
and U27152 (N_27152,N_25462,N_24732);
or U27153 (N_27153,N_25711,N_24331);
nor U27154 (N_27154,N_25786,N_24666);
xnor U27155 (N_27155,N_24271,N_24580);
nand U27156 (N_27156,N_25731,N_24613);
nand U27157 (N_27157,N_25349,N_24030);
xor U27158 (N_27158,N_25712,N_25759);
nand U27159 (N_27159,N_25498,N_24398);
and U27160 (N_27160,N_25444,N_25975);
or U27161 (N_27161,N_25351,N_25585);
nand U27162 (N_27162,N_24748,N_25043);
and U27163 (N_27163,N_25100,N_25572);
and U27164 (N_27164,N_25061,N_25972);
and U27165 (N_27165,N_24068,N_25956);
nor U27166 (N_27166,N_24984,N_24232);
or U27167 (N_27167,N_25164,N_25104);
xnor U27168 (N_27168,N_24652,N_24117);
nor U27169 (N_27169,N_25061,N_25532);
xnor U27170 (N_27170,N_25584,N_24563);
and U27171 (N_27171,N_25712,N_25426);
nor U27172 (N_27172,N_24895,N_25877);
or U27173 (N_27173,N_25917,N_24587);
xor U27174 (N_27174,N_24751,N_25812);
xor U27175 (N_27175,N_24888,N_24356);
nor U27176 (N_27176,N_24770,N_25195);
xnor U27177 (N_27177,N_24639,N_24716);
nand U27178 (N_27178,N_25652,N_25045);
nor U27179 (N_27179,N_25501,N_24225);
nand U27180 (N_27180,N_24157,N_25648);
nand U27181 (N_27181,N_25180,N_25174);
or U27182 (N_27182,N_25620,N_24913);
nor U27183 (N_27183,N_24725,N_25033);
and U27184 (N_27184,N_25093,N_25793);
nor U27185 (N_27185,N_24204,N_24570);
nand U27186 (N_27186,N_24612,N_24553);
or U27187 (N_27187,N_25070,N_25028);
and U27188 (N_27188,N_24298,N_24365);
or U27189 (N_27189,N_25679,N_24001);
nand U27190 (N_27190,N_25222,N_25083);
nor U27191 (N_27191,N_24291,N_24767);
and U27192 (N_27192,N_25557,N_24274);
or U27193 (N_27193,N_25052,N_25270);
and U27194 (N_27194,N_24858,N_25725);
nand U27195 (N_27195,N_25701,N_24922);
nand U27196 (N_27196,N_24238,N_24569);
nand U27197 (N_27197,N_25192,N_24601);
nor U27198 (N_27198,N_25382,N_25910);
nand U27199 (N_27199,N_25313,N_25677);
nand U27200 (N_27200,N_24786,N_24075);
nor U27201 (N_27201,N_24810,N_25952);
and U27202 (N_27202,N_24654,N_24220);
xnor U27203 (N_27203,N_24286,N_24024);
nor U27204 (N_27204,N_25042,N_24218);
or U27205 (N_27205,N_24722,N_24850);
and U27206 (N_27206,N_24515,N_24043);
and U27207 (N_27207,N_24508,N_25631);
or U27208 (N_27208,N_25865,N_24831);
nor U27209 (N_27209,N_25974,N_25807);
or U27210 (N_27210,N_24086,N_24717);
and U27211 (N_27211,N_25564,N_24814);
xor U27212 (N_27212,N_25882,N_25867);
nand U27213 (N_27213,N_25780,N_24892);
and U27214 (N_27214,N_24687,N_24212);
and U27215 (N_27215,N_25926,N_25292);
xor U27216 (N_27216,N_24066,N_25511);
and U27217 (N_27217,N_25511,N_25691);
and U27218 (N_27218,N_25103,N_25048);
nor U27219 (N_27219,N_25070,N_25312);
and U27220 (N_27220,N_24543,N_24631);
xor U27221 (N_27221,N_24860,N_24680);
nand U27222 (N_27222,N_24906,N_24820);
xor U27223 (N_27223,N_24885,N_25526);
nand U27224 (N_27224,N_25316,N_24309);
nand U27225 (N_27225,N_25479,N_25597);
nand U27226 (N_27226,N_24978,N_24683);
nand U27227 (N_27227,N_24269,N_25023);
and U27228 (N_27228,N_24839,N_24488);
or U27229 (N_27229,N_24917,N_24624);
or U27230 (N_27230,N_24738,N_24703);
and U27231 (N_27231,N_25776,N_25239);
or U27232 (N_27232,N_25615,N_24500);
nand U27233 (N_27233,N_25489,N_25977);
nand U27234 (N_27234,N_24000,N_24914);
nand U27235 (N_27235,N_25027,N_25552);
nand U27236 (N_27236,N_24048,N_24500);
nor U27237 (N_27237,N_25138,N_25080);
and U27238 (N_27238,N_24382,N_24289);
xor U27239 (N_27239,N_24448,N_25643);
xnor U27240 (N_27240,N_25312,N_25841);
xor U27241 (N_27241,N_25305,N_25263);
or U27242 (N_27242,N_24086,N_25493);
nand U27243 (N_27243,N_25858,N_25562);
or U27244 (N_27244,N_25427,N_25454);
or U27245 (N_27245,N_25517,N_25127);
nor U27246 (N_27246,N_25229,N_24129);
nand U27247 (N_27247,N_24743,N_25295);
and U27248 (N_27248,N_24008,N_25217);
and U27249 (N_27249,N_24681,N_24450);
xor U27250 (N_27250,N_25385,N_24513);
xor U27251 (N_27251,N_24909,N_25207);
nand U27252 (N_27252,N_24340,N_25895);
xnor U27253 (N_27253,N_25492,N_25617);
nor U27254 (N_27254,N_25644,N_24151);
xnor U27255 (N_27255,N_25720,N_24129);
and U27256 (N_27256,N_25332,N_24858);
and U27257 (N_27257,N_25184,N_24028);
and U27258 (N_27258,N_25514,N_25933);
or U27259 (N_27259,N_24712,N_25696);
xnor U27260 (N_27260,N_25597,N_25760);
nand U27261 (N_27261,N_25573,N_24018);
and U27262 (N_27262,N_24437,N_25904);
nor U27263 (N_27263,N_24629,N_24771);
xor U27264 (N_27264,N_25846,N_24879);
nor U27265 (N_27265,N_24353,N_25539);
xor U27266 (N_27266,N_24024,N_24944);
xnor U27267 (N_27267,N_25267,N_24211);
or U27268 (N_27268,N_24434,N_24577);
and U27269 (N_27269,N_25379,N_24996);
and U27270 (N_27270,N_25227,N_25072);
xnor U27271 (N_27271,N_25748,N_24329);
nor U27272 (N_27272,N_24479,N_24276);
nor U27273 (N_27273,N_25195,N_25525);
nand U27274 (N_27274,N_24883,N_25403);
xor U27275 (N_27275,N_24379,N_25384);
and U27276 (N_27276,N_24467,N_25255);
nand U27277 (N_27277,N_24364,N_25170);
nand U27278 (N_27278,N_25566,N_25108);
nand U27279 (N_27279,N_25533,N_24387);
xnor U27280 (N_27280,N_24876,N_25089);
nand U27281 (N_27281,N_25344,N_24295);
nand U27282 (N_27282,N_25566,N_24401);
or U27283 (N_27283,N_25112,N_24219);
nand U27284 (N_27284,N_25482,N_24751);
and U27285 (N_27285,N_25286,N_24874);
and U27286 (N_27286,N_24424,N_24833);
and U27287 (N_27287,N_24511,N_25306);
nor U27288 (N_27288,N_25395,N_25013);
nor U27289 (N_27289,N_25067,N_24242);
nand U27290 (N_27290,N_24744,N_24095);
xor U27291 (N_27291,N_25428,N_24502);
and U27292 (N_27292,N_24907,N_25089);
xnor U27293 (N_27293,N_24665,N_24401);
nand U27294 (N_27294,N_25783,N_25303);
nor U27295 (N_27295,N_25864,N_24875);
and U27296 (N_27296,N_24039,N_24811);
or U27297 (N_27297,N_25696,N_24291);
and U27298 (N_27298,N_25516,N_25904);
xnor U27299 (N_27299,N_25876,N_24624);
xnor U27300 (N_27300,N_24033,N_24055);
or U27301 (N_27301,N_25479,N_25948);
nand U27302 (N_27302,N_24399,N_25441);
nor U27303 (N_27303,N_24005,N_25612);
nand U27304 (N_27304,N_24003,N_24461);
xnor U27305 (N_27305,N_24636,N_25747);
or U27306 (N_27306,N_24493,N_24935);
or U27307 (N_27307,N_25386,N_25927);
xnor U27308 (N_27308,N_25378,N_24121);
and U27309 (N_27309,N_24790,N_24695);
and U27310 (N_27310,N_25695,N_25898);
xor U27311 (N_27311,N_25614,N_25490);
nor U27312 (N_27312,N_24754,N_24237);
xnor U27313 (N_27313,N_24011,N_25882);
nand U27314 (N_27314,N_24012,N_25970);
or U27315 (N_27315,N_25424,N_24816);
xor U27316 (N_27316,N_24015,N_25452);
and U27317 (N_27317,N_25862,N_25994);
xnor U27318 (N_27318,N_25369,N_25094);
xnor U27319 (N_27319,N_24451,N_24207);
or U27320 (N_27320,N_24621,N_24922);
or U27321 (N_27321,N_24326,N_24254);
and U27322 (N_27322,N_25040,N_24602);
and U27323 (N_27323,N_24985,N_25359);
and U27324 (N_27324,N_24978,N_24038);
or U27325 (N_27325,N_25394,N_24684);
or U27326 (N_27326,N_25235,N_24477);
or U27327 (N_27327,N_24104,N_24881);
nor U27328 (N_27328,N_25833,N_24640);
nand U27329 (N_27329,N_24049,N_24905);
and U27330 (N_27330,N_25088,N_25204);
or U27331 (N_27331,N_24591,N_25145);
and U27332 (N_27332,N_25273,N_25566);
and U27333 (N_27333,N_24567,N_24160);
or U27334 (N_27334,N_25710,N_24714);
and U27335 (N_27335,N_24260,N_25032);
or U27336 (N_27336,N_24787,N_24039);
nand U27337 (N_27337,N_24227,N_24352);
nand U27338 (N_27338,N_24174,N_25999);
nand U27339 (N_27339,N_24000,N_24993);
or U27340 (N_27340,N_24454,N_24441);
nor U27341 (N_27341,N_24199,N_25599);
nand U27342 (N_27342,N_25079,N_24750);
nor U27343 (N_27343,N_24884,N_24158);
xor U27344 (N_27344,N_25108,N_25685);
or U27345 (N_27345,N_24305,N_25940);
xor U27346 (N_27346,N_25184,N_24060);
nand U27347 (N_27347,N_25883,N_24390);
nand U27348 (N_27348,N_24644,N_25906);
xnor U27349 (N_27349,N_24336,N_24682);
or U27350 (N_27350,N_25317,N_24671);
or U27351 (N_27351,N_24451,N_24819);
and U27352 (N_27352,N_25224,N_24169);
or U27353 (N_27353,N_25408,N_24905);
xnor U27354 (N_27354,N_24927,N_25317);
and U27355 (N_27355,N_25236,N_24677);
or U27356 (N_27356,N_25388,N_24309);
or U27357 (N_27357,N_25926,N_25811);
nor U27358 (N_27358,N_24287,N_25833);
xor U27359 (N_27359,N_24406,N_24045);
or U27360 (N_27360,N_25152,N_24791);
nand U27361 (N_27361,N_25090,N_25155);
or U27362 (N_27362,N_25900,N_24703);
or U27363 (N_27363,N_24348,N_24599);
nor U27364 (N_27364,N_24932,N_25970);
and U27365 (N_27365,N_25001,N_24344);
nand U27366 (N_27366,N_24270,N_25736);
and U27367 (N_27367,N_24040,N_24400);
xnor U27368 (N_27368,N_24764,N_25285);
xnor U27369 (N_27369,N_25666,N_25227);
nor U27370 (N_27370,N_25775,N_25191);
xnor U27371 (N_27371,N_25259,N_24597);
and U27372 (N_27372,N_24540,N_25278);
xor U27373 (N_27373,N_24301,N_25919);
nor U27374 (N_27374,N_25527,N_25034);
nor U27375 (N_27375,N_24230,N_25114);
xnor U27376 (N_27376,N_24898,N_25865);
or U27377 (N_27377,N_25941,N_25687);
xnor U27378 (N_27378,N_25902,N_25996);
or U27379 (N_27379,N_24949,N_24379);
and U27380 (N_27380,N_24452,N_24290);
nor U27381 (N_27381,N_24012,N_24957);
and U27382 (N_27382,N_25920,N_25282);
or U27383 (N_27383,N_25686,N_24772);
or U27384 (N_27384,N_24821,N_25528);
nor U27385 (N_27385,N_24438,N_25061);
nor U27386 (N_27386,N_25585,N_24696);
or U27387 (N_27387,N_24026,N_25413);
or U27388 (N_27388,N_24987,N_24842);
nand U27389 (N_27389,N_24818,N_25690);
nand U27390 (N_27390,N_25204,N_25511);
nand U27391 (N_27391,N_25049,N_25400);
xor U27392 (N_27392,N_25332,N_24917);
and U27393 (N_27393,N_24051,N_25242);
xor U27394 (N_27394,N_25437,N_25331);
or U27395 (N_27395,N_24925,N_24360);
nor U27396 (N_27396,N_25828,N_24697);
xor U27397 (N_27397,N_25244,N_25898);
or U27398 (N_27398,N_24171,N_24504);
or U27399 (N_27399,N_24035,N_25527);
nand U27400 (N_27400,N_24501,N_24411);
nand U27401 (N_27401,N_25691,N_24713);
xor U27402 (N_27402,N_24273,N_25089);
xor U27403 (N_27403,N_24337,N_24407);
xnor U27404 (N_27404,N_24400,N_25110);
or U27405 (N_27405,N_24612,N_24484);
or U27406 (N_27406,N_24130,N_24254);
nor U27407 (N_27407,N_25152,N_24013);
xor U27408 (N_27408,N_24262,N_25050);
nand U27409 (N_27409,N_24009,N_25918);
and U27410 (N_27410,N_25954,N_24874);
nor U27411 (N_27411,N_25533,N_25279);
nor U27412 (N_27412,N_25625,N_25098);
and U27413 (N_27413,N_25680,N_25052);
and U27414 (N_27414,N_25474,N_24723);
or U27415 (N_27415,N_25856,N_25245);
nor U27416 (N_27416,N_24399,N_25251);
and U27417 (N_27417,N_25099,N_25246);
nand U27418 (N_27418,N_25542,N_25441);
nand U27419 (N_27419,N_25937,N_25957);
and U27420 (N_27420,N_25293,N_24227);
xor U27421 (N_27421,N_24871,N_24806);
nand U27422 (N_27422,N_25854,N_24350);
nor U27423 (N_27423,N_24022,N_25854);
and U27424 (N_27424,N_25583,N_24014);
and U27425 (N_27425,N_25421,N_24874);
and U27426 (N_27426,N_24943,N_25170);
or U27427 (N_27427,N_25898,N_25096);
nor U27428 (N_27428,N_25794,N_25081);
or U27429 (N_27429,N_24679,N_25188);
nand U27430 (N_27430,N_24194,N_24465);
nand U27431 (N_27431,N_24569,N_24976);
nand U27432 (N_27432,N_25944,N_25326);
nor U27433 (N_27433,N_24279,N_25115);
xor U27434 (N_27434,N_24207,N_24684);
and U27435 (N_27435,N_25042,N_24479);
and U27436 (N_27436,N_24703,N_24754);
or U27437 (N_27437,N_25749,N_25974);
nor U27438 (N_27438,N_24358,N_25493);
nor U27439 (N_27439,N_25269,N_25373);
nor U27440 (N_27440,N_24565,N_25969);
nor U27441 (N_27441,N_25633,N_25942);
nor U27442 (N_27442,N_25378,N_25402);
nand U27443 (N_27443,N_24788,N_25255);
xnor U27444 (N_27444,N_25528,N_25818);
or U27445 (N_27445,N_25020,N_25973);
nand U27446 (N_27446,N_24383,N_25058);
nand U27447 (N_27447,N_24721,N_25630);
nor U27448 (N_27448,N_25562,N_24025);
xnor U27449 (N_27449,N_25188,N_24163);
nand U27450 (N_27450,N_25351,N_24617);
nand U27451 (N_27451,N_25441,N_25955);
nand U27452 (N_27452,N_25937,N_25201);
and U27453 (N_27453,N_25193,N_24972);
or U27454 (N_27454,N_25508,N_25099);
xnor U27455 (N_27455,N_24308,N_25995);
nor U27456 (N_27456,N_25387,N_25567);
nor U27457 (N_27457,N_24120,N_24466);
nor U27458 (N_27458,N_24027,N_25503);
or U27459 (N_27459,N_24708,N_24967);
nand U27460 (N_27460,N_24964,N_24733);
and U27461 (N_27461,N_24644,N_24762);
xnor U27462 (N_27462,N_24810,N_25566);
xnor U27463 (N_27463,N_25582,N_25445);
nor U27464 (N_27464,N_25775,N_25391);
xor U27465 (N_27465,N_25681,N_25114);
nor U27466 (N_27466,N_24746,N_24539);
nor U27467 (N_27467,N_25783,N_25336);
or U27468 (N_27468,N_24779,N_24304);
nor U27469 (N_27469,N_25425,N_25785);
and U27470 (N_27470,N_24034,N_25883);
nor U27471 (N_27471,N_24438,N_25633);
or U27472 (N_27472,N_24586,N_24280);
nand U27473 (N_27473,N_25161,N_24157);
or U27474 (N_27474,N_25526,N_25360);
xnor U27475 (N_27475,N_25791,N_24583);
nand U27476 (N_27476,N_25296,N_24101);
and U27477 (N_27477,N_25304,N_25312);
or U27478 (N_27478,N_25586,N_24378);
nor U27479 (N_27479,N_25420,N_25610);
or U27480 (N_27480,N_25684,N_25848);
xnor U27481 (N_27481,N_24212,N_24067);
nor U27482 (N_27482,N_24552,N_25726);
nor U27483 (N_27483,N_25515,N_25539);
and U27484 (N_27484,N_24292,N_24963);
or U27485 (N_27485,N_25094,N_24946);
nand U27486 (N_27486,N_25224,N_25646);
and U27487 (N_27487,N_25843,N_24226);
and U27488 (N_27488,N_25901,N_24324);
nor U27489 (N_27489,N_25099,N_25926);
nor U27490 (N_27490,N_25952,N_24512);
or U27491 (N_27491,N_25819,N_24779);
nor U27492 (N_27492,N_24083,N_24842);
nand U27493 (N_27493,N_24039,N_24006);
nand U27494 (N_27494,N_24630,N_24741);
or U27495 (N_27495,N_24411,N_24705);
nand U27496 (N_27496,N_24860,N_24949);
nand U27497 (N_27497,N_24936,N_24815);
nor U27498 (N_27498,N_24595,N_25515);
and U27499 (N_27499,N_25273,N_25236);
or U27500 (N_27500,N_24835,N_25319);
nor U27501 (N_27501,N_24732,N_24620);
xor U27502 (N_27502,N_24622,N_25038);
or U27503 (N_27503,N_25645,N_24629);
and U27504 (N_27504,N_24310,N_25118);
and U27505 (N_27505,N_24146,N_25257);
or U27506 (N_27506,N_25820,N_25858);
or U27507 (N_27507,N_24710,N_24006);
nand U27508 (N_27508,N_24665,N_24055);
or U27509 (N_27509,N_25043,N_24294);
or U27510 (N_27510,N_25765,N_25154);
nor U27511 (N_27511,N_24316,N_25221);
and U27512 (N_27512,N_24888,N_25696);
nand U27513 (N_27513,N_25733,N_24736);
or U27514 (N_27514,N_24295,N_24376);
nand U27515 (N_27515,N_25588,N_24304);
or U27516 (N_27516,N_25476,N_25339);
nor U27517 (N_27517,N_24082,N_25019);
nor U27518 (N_27518,N_24568,N_25801);
or U27519 (N_27519,N_24392,N_24258);
and U27520 (N_27520,N_25613,N_24953);
and U27521 (N_27521,N_25974,N_25810);
and U27522 (N_27522,N_25522,N_25634);
xnor U27523 (N_27523,N_25999,N_25887);
xor U27524 (N_27524,N_24846,N_24264);
nand U27525 (N_27525,N_25135,N_25124);
and U27526 (N_27526,N_24657,N_24953);
and U27527 (N_27527,N_24773,N_25153);
and U27528 (N_27528,N_25200,N_25025);
and U27529 (N_27529,N_24072,N_25902);
nor U27530 (N_27530,N_25694,N_25735);
and U27531 (N_27531,N_25226,N_25132);
or U27532 (N_27532,N_25402,N_25801);
or U27533 (N_27533,N_25950,N_25240);
or U27534 (N_27534,N_25737,N_25243);
xor U27535 (N_27535,N_25007,N_24344);
xor U27536 (N_27536,N_24393,N_25982);
and U27537 (N_27537,N_25763,N_25527);
nand U27538 (N_27538,N_25060,N_25196);
nand U27539 (N_27539,N_25675,N_24954);
nand U27540 (N_27540,N_25150,N_24736);
xor U27541 (N_27541,N_24599,N_25335);
or U27542 (N_27542,N_25102,N_25862);
xor U27543 (N_27543,N_24995,N_24797);
nor U27544 (N_27544,N_24538,N_24626);
xnor U27545 (N_27545,N_24111,N_25369);
xnor U27546 (N_27546,N_25227,N_24549);
xor U27547 (N_27547,N_24212,N_25671);
or U27548 (N_27548,N_24305,N_24773);
or U27549 (N_27549,N_25189,N_25266);
nor U27550 (N_27550,N_25304,N_24360);
xor U27551 (N_27551,N_25050,N_25501);
nand U27552 (N_27552,N_25577,N_25064);
nand U27553 (N_27553,N_25531,N_25438);
and U27554 (N_27554,N_25145,N_25459);
or U27555 (N_27555,N_24210,N_25837);
or U27556 (N_27556,N_24690,N_24026);
nor U27557 (N_27557,N_24635,N_24164);
xnor U27558 (N_27558,N_25106,N_25387);
nor U27559 (N_27559,N_25783,N_24500);
and U27560 (N_27560,N_25614,N_25073);
nor U27561 (N_27561,N_24858,N_24320);
or U27562 (N_27562,N_25183,N_24075);
nand U27563 (N_27563,N_25324,N_24374);
nor U27564 (N_27564,N_24651,N_25471);
nor U27565 (N_27565,N_24652,N_25136);
nor U27566 (N_27566,N_25406,N_25502);
nand U27567 (N_27567,N_25683,N_25667);
nand U27568 (N_27568,N_24188,N_25934);
nand U27569 (N_27569,N_25226,N_24398);
and U27570 (N_27570,N_24078,N_24833);
nand U27571 (N_27571,N_24068,N_24676);
nand U27572 (N_27572,N_24531,N_24076);
nand U27573 (N_27573,N_25255,N_25987);
nand U27574 (N_27574,N_25190,N_25250);
nor U27575 (N_27575,N_25674,N_25235);
and U27576 (N_27576,N_25140,N_25018);
nor U27577 (N_27577,N_24336,N_24720);
nand U27578 (N_27578,N_24911,N_24170);
or U27579 (N_27579,N_24575,N_24578);
xnor U27580 (N_27580,N_24155,N_24543);
and U27581 (N_27581,N_24203,N_25885);
and U27582 (N_27582,N_25069,N_24094);
nand U27583 (N_27583,N_25476,N_25526);
nor U27584 (N_27584,N_24513,N_24240);
nor U27585 (N_27585,N_25092,N_24832);
nor U27586 (N_27586,N_25428,N_24309);
and U27587 (N_27587,N_24284,N_25301);
nor U27588 (N_27588,N_24893,N_25990);
nand U27589 (N_27589,N_25094,N_24912);
and U27590 (N_27590,N_25341,N_24660);
xor U27591 (N_27591,N_25465,N_24391);
or U27592 (N_27592,N_25842,N_24302);
xor U27593 (N_27593,N_24237,N_24482);
or U27594 (N_27594,N_25816,N_25451);
nor U27595 (N_27595,N_25930,N_24712);
nor U27596 (N_27596,N_24017,N_25468);
xor U27597 (N_27597,N_25391,N_25462);
nand U27598 (N_27598,N_25398,N_25380);
nand U27599 (N_27599,N_24107,N_24270);
xor U27600 (N_27600,N_25082,N_25390);
nor U27601 (N_27601,N_25475,N_24899);
and U27602 (N_27602,N_24933,N_25889);
or U27603 (N_27603,N_24578,N_24205);
and U27604 (N_27604,N_24933,N_24593);
nand U27605 (N_27605,N_25541,N_24619);
or U27606 (N_27606,N_25100,N_24232);
and U27607 (N_27607,N_24589,N_25546);
nand U27608 (N_27608,N_25418,N_24032);
xnor U27609 (N_27609,N_24496,N_25616);
or U27610 (N_27610,N_24728,N_24350);
and U27611 (N_27611,N_24438,N_24956);
nand U27612 (N_27612,N_24613,N_25288);
nand U27613 (N_27613,N_24126,N_24363);
nand U27614 (N_27614,N_25265,N_25411);
xor U27615 (N_27615,N_25084,N_24912);
xnor U27616 (N_27616,N_24131,N_24041);
xor U27617 (N_27617,N_24105,N_25585);
nor U27618 (N_27618,N_24372,N_24010);
nor U27619 (N_27619,N_25686,N_25854);
and U27620 (N_27620,N_25618,N_24071);
and U27621 (N_27621,N_24058,N_25176);
and U27622 (N_27622,N_25529,N_25911);
and U27623 (N_27623,N_25764,N_25281);
xnor U27624 (N_27624,N_24865,N_24414);
nand U27625 (N_27625,N_24711,N_25878);
and U27626 (N_27626,N_25524,N_24705);
nand U27627 (N_27627,N_25459,N_25896);
nor U27628 (N_27628,N_25197,N_25600);
nor U27629 (N_27629,N_25527,N_24193);
xor U27630 (N_27630,N_25071,N_24658);
xor U27631 (N_27631,N_25849,N_25893);
and U27632 (N_27632,N_25487,N_24736);
nor U27633 (N_27633,N_24409,N_24156);
and U27634 (N_27634,N_24022,N_25533);
xor U27635 (N_27635,N_24494,N_25068);
xor U27636 (N_27636,N_24621,N_25888);
xnor U27637 (N_27637,N_24215,N_25824);
xor U27638 (N_27638,N_24982,N_25000);
nand U27639 (N_27639,N_25011,N_24893);
or U27640 (N_27640,N_24029,N_25660);
or U27641 (N_27641,N_25650,N_25240);
nor U27642 (N_27642,N_24069,N_24533);
nand U27643 (N_27643,N_25118,N_25667);
xor U27644 (N_27644,N_24702,N_25987);
nand U27645 (N_27645,N_24027,N_25554);
or U27646 (N_27646,N_25219,N_24194);
and U27647 (N_27647,N_24450,N_24279);
nor U27648 (N_27648,N_25083,N_25488);
xor U27649 (N_27649,N_25574,N_24876);
nor U27650 (N_27650,N_25020,N_24728);
and U27651 (N_27651,N_24900,N_24410);
nor U27652 (N_27652,N_24163,N_24134);
nand U27653 (N_27653,N_24767,N_24779);
and U27654 (N_27654,N_25101,N_24846);
nand U27655 (N_27655,N_24983,N_24587);
xor U27656 (N_27656,N_25844,N_25712);
or U27657 (N_27657,N_25533,N_24856);
nand U27658 (N_27658,N_25561,N_25337);
xor U27659 (N_27659,N_25489,N_25112);
or U27660 (N_27660,N_25567,N_24745);
or U27661 (N_27661,N_24984,N_24829);
nand U27662 (N_27662,N_25284,N_24709);
xor U27663 (N_27663,N_24008,N_24826);
and U27664 (N_27664,N_24965,N_24950);
and U27665 (N_27665,N_25581,N_24654);
nand U27666 (N_27666,N_25482,N_25863);
or U27667 (N_27667,N_25517,N_24802);
and U27668 (N_27668,N_25067,N_25425);
xor U27669 (N_27669,N_24498,N_24958);
or U27670 (N_27670,N_24908,N_25082);
and U27671 (N_27671,N_25912,N_24027);
and U27672 (N_27672,N_25473,N_25827);
nand U27673 (N_27673,N_24538,N_25671);
nor U27674 (N_27674,N_24879,N_25448);
or U27675 (N_27675,N_25526,N_25509);
nand U27676 (N_27676,N_25999,N_24132);
nand U27677 (N_27677,N_24093,N_24849);
nor U27678 (N_27678,N_24758,N_24748);
xor U27679 (N_27679,N_25671,N_25716);
xor U27680 (N_27680,N_25732,N_24412);
nand U27681 (N_27681,N_25302,N_24305);
nor U27682 (N_27682,N_24055,N_24430);
nand U27683 (N_27683,N_24740,N_25957);
and U27684 (N_27684,N_24986,N_25562);
xor U27685 (N_27685,N_25534,N_24087);
or U27686 (N_27686,N_24039,N_24864);
xor U27687 (N_27687,N_24305,N_24537);
nand U27688 (N_27688,N_25225,N_25165);
nand U27689 (N_27689,N_25952,N_25620);
and U27690 (N_27690,N_25554,N_25610);
xor U27691 (N_27691,N_24987,N_25789);
and U27692 (N_27692,N_24365,N_25995);
or U27693 (N_27693,N_24224,N_24308);
xor U27694 (N_27694,N_25931,N_24054);
nand U27695 (N_27695,N_25781,N_25107);
and U27696 (N_27696,N_24806,N_25880);
nand U27697 (N_27697,N_25808,N_25312);
xnor U27698 (N_27698,N_24593,N_24677);
xnor U27699 (N_27699,N_25832,N_24348);
nand U27700 (N_27700,N_25587,N_24816);
and U27701 (N_27701,N_24358,N_24675);
nand U27702 (N_27702,N_25444,N_24630);
nand U27703 (N_27703,N_24080,N_25949);
nor U27704 (N_27704,N_25285,N_24530);
and U27705 (N_27705,N_24536,N_24012);
and U27706 (N_27706,N_24176,N_24940);
xnor U27707 (N_27707,N_24694,N_25292);
xnor U27708 (N_27708,N_24857,N_24688);
nor U27709 (N_27709,N_24113,N_24841);
nor U27710 (N_27710,N_24074,N_24386);
or U27711 (N_27711,N_24219,N_25041);
and U27712 (N_27712,N_25163,N_25949);
nand U27713 (N_27713,N_25984,N_25794);
nor U27714 (N_27714,N_25136,N_24000);
and U27715 (N_27715,N_24255,N_25958);
xor U27716 (N_27716,N_24468,N_24083);
and U27717 (N_27717,N_24552,N_24555);
xor U27718 (N_27718,N_25929,N_25207);
and U27719 (N_27719,N_25421,N_25080);
and U27720 (N_27720,N_25474,N_24887);
nand U27721 (N_27721,N_24145,N_24302);
xnor U27722 (N_27722,N_25723,N_25292);
nand U27723 (N_27723,N_24643,N_24995);
xnor U27724 (N_27724,N_25615,N_25934);
nor U27725 (N_27725,N_25114,N_24210);
or U27726 (N_27726,N_24754,N_25404);
nor U27727 (N_27727,N_24044,N_24253);
and U27728 (N_27728,N_25771,N_24378);
nand U27729 (N_27729,N_24263,N_24312);
and U27730 (N_27730,N_24227,N_24202);
nor U27731 (N_27731,N_25161,N_24087);
nor U27732 (N_27732,N_24571,N_25860);
nand U27733 (N_27733,N_25651,N_25747);
nor U27734 (N_27734,N_24879,N_25755);
and U27735 (N_27735,N_25926,N_24939);
nor U27736 (N_27736,N_25114,N_25582);
xor U27737 (N_27737,N_24411,N_25945);
xnor U27738 (N_27738,N_24388,N_25325);
nand U27739 (N_27739,N_25197,N_24314);
or U27740 (N_27740,N_25285,N_24798);
and U27741 (N_27741,N_25885,N_24471);
or U27742 (N_27742,N_24509,N_25684);
nor U27743 (N_27743,N_24677,N_25135);
and U27744 (N_27744,N_24909,N_24055);
xnor U27745 (N_27745,N_25462,N_24815);
nand U27746 (N_27746,N_24965,N_24419);
or U27747 (N_27747,N_25512,N_25086);
xnor U27748 (N_27748,N_25881,N_25209);
and U27749 (N_27749,N_24929,N_24387);
nor U27750 (N_27750,N_24966,N_24343);
nor U27751 (N_27751,N_25707,N_24922);
nor U27752 (N_27752,N_25634,N_25268);
xor U27753 (N_27753,N_24907,N_25778);
and U27754 (N_27754,N_25863,N_24678);
xnor U27755 (N_27755,N_24782,N_25982);
nand U27756 (N_27756,N_25650,N_24761);
and U27757 (N_27757,N_24084,N_24161);
or U27758 (N_27758,N_24171,N_25100);
nor U27759 (N_27759,N_24837,N_25822);
nand U27760 (N_27760,N_24548,N_25138);
or U27761 (N_27761,N_25110,N_25713);
or U27762 (N_27762,N_24275,N_25523);
nand U27763 (N_27763,N_25555,N_25846);
nor U27764 (N_27764,N_25574,N_24937);
and U27765 (N_27765,N_25399,N_24737);
nor U27766 (N_27766,N_25777,N_25323);
or U27767 (N_27767,N_25662,N_25309);
nor U27768 (N_27768,N_24937,N_25249);
or U27769 (N_27769,N_24653,N_25820);
xor U27770 (N_27770,N_25325,N_24564);
xor U27771 (N_27771,N_24457,N_25031);
and U27772 (N_27772,N_24185,N_25446);
xor U27773 (N_27773,N_24829,N_24368);
and U27774 (N_27774,N_25798,N_25600);
or U27775 (N_27775,N_24020,N_24111);
nor U27776 (N_27776,N_24546,N_25002);
nand U27777 (N_27777,N_24500,N_24972);
and U27778 (N_27778,N_25493,N_25990);
and U27779 (N_27779,N_25812,N_25736);
and U27780 (N_27780,N_25805,N_24472);
nor U27781 (N_27781,N_24085,N_25808);
xor U27782 (N_27782,N_24504,N_25821);
nor U27783 (N_27783,N_24562,N_24963);
nand U27784 (N_27784,N_24816,N_25430);
and U27785 (N_27785,N_24268,N_24088);
or U27786 (N_27786,N_25012,N_24881);
xor U27787 (N_27787,N_25914,N_25481);
or U27788 (N_27788,N_25459,N_25836);
and U27789 (N_27789,N_25525,N_25413);
xnor U27790 (N_27790,N_25900,N_25201);
xor U27791 (N_27791,N_25833,N_25603);
or U27792 (N_27792,N_24232,N_25377);
and U27793 (N_27793,N_25158,N_25622);
nor U27794 (N_27794,N_25731,N_25755);
nor U27795 (N_27795,N_24725,N_25676);
and U27796 (N_27796,N_24568,N_25003);
and U27797 (N_27797,N_25564,N_25451);
xnor U27798 (N_27798,N_24864,N_24976);
nor U27799 (N_27799,N_25463,N_24841);
and U27800 (N_27800,N_25637,N_25554);
or U27801 (N_27801,N_24965,N_25229);
nor U27802 (N_27802,N_24954,N_25018);
and U27803 (N_27803,N_24938,N_25370);
nand U27804 (N_27804,N_25725,N_24911);
nand U27805 (N_27805,N_24038,N_25545);
or U27806 (N_27806,N_25876,N_24866);
or U27807 (N_27807,N_25820,N_25350);
xor U27808 (N_27808,N_25738,N_25482);
or U27809 (N_27809,N_25488,N_25122);
or U27810 (N_27810,N_25787,N_24496);
nor U27811 (N_27811,N_25782,N_25033);
nand U27812 (N_27812,N_24375,N_25319);
xor U27813 (N_27813,N_25272,N_24457);
nor U27814 (N_27814,N_25298,N_24486);
and U27815 (N_27815,N_24987,N_25620);
nor U27816 (N_27816,N_24270,N_24502);
nand U27817 (N_27817,N_24834,N_24559);
nor U27818 (N_27818,N_24157,N_24233);
nor U27819 (N_27819,N_25934,N_24945);
xor U27820 (N_27820,N_25053,N_24299);
or U27821 (N_27821,N_24273,N_25675);
xor U27822 (N_27822,N_25260,N_24132);
and U27823 (N_27823,N_25191,N_24059);
or U27824 (N_27824,N_25285,N_24369);
nor U27825 (N_27825,N_25621,N_25374);
nor U27826 (N_27826,N_25381,N_25085);
nor U27827 (N_27827,N_25063,N_24412);
or U27828 (N_27828,N_24017,N_24960);
nor U27829 (N_27829,N_24235,N_25093);
nand U27830 (N_27830,N_24766,N_24482);
nand U27831 (N_27831,N_25808,N_24378);
nor U27832 (N_27832,N_25696,N_25358);
and U27833 (N_27833,N_24554,N_24472);
xor U27834 (N_27834,N_24622,N_24395);
and U27835 (N_27835,N_24577,N_25101);
and U27836 (N_27836,N_24893,N_24580);
nand U27837 (N_27837,N_24888,N_24917);
xor U27838 (N_27838,N_24769,N_24935);
and U27839 (N_27839,N_24190,N_24713);
or U27840 (N_27840,N_25011,N_25274);
or U27841 (N_27841,N_24467,N_24820);
or U27842 (N_27842,N_25343,N_24389);
or U27843 (N_27843,N_25167,N_24287);
and U27844 (N_27844,N_25832,N_25157);
nor U27845 (N_27845,N_25355,N_25220);
xnor U27846 (N_27846,N_24652,N_24615);
nand U27847 (N_27847,N_24681,N_24510);
and U27848 (N_27848,N_25896,N_25265);
xor U27849 (N_27849,N_24137,N_24856);
nor U27850 (N_27850,N_24565,N_25803);
or U27851 (N_27851,N_25047,N_25583);
nor U27852 (N_27852,N_25872,N_25069);
xor U27853 (N_27853,N_24837,N_25347);
or U27854 (N_27854,N_24876,N_25108);
nand U27855 (N_27855,N_24252,N_24183);
and U27856 (N_27856,N_24280,N_25189);
and U27857 (N_27857,N_25841,N_25584);
xnor U27858 (N_27858,N_25137,N_25839);
nand U27859 (N_27859,N_25786,N_25862);
xnor U27860 (N_27860,N_24596,N_24559);
and U27861 (N_27861,N_25605,N_25165);
and U27862 (N_27862,N_24659,N_24420);
nor U27863 (N_27863,N_25217,N_24570);
and U27864 (N_27864,N_24874,N_24496);
nor U27865 (N_27865,N_24370,N_24193);
and U27866 (N_27866,N_25458,N_25948);
nand U27867 (N_27867,N_24990,N_24534);
nand U27868 (N_27868,N_25765,N_25943);
nand U27869 (N_27869,N_25893,N_24159);
xnor U27870 (N_27870,N_25651,N_24528);
xor U27871 (N_27871,N_25968,N_24447);
nor U27872 (N_27872,N_24588,N_24387);
xnor U27873 (N_27873,N_25650,N_25559);
nor U27874 (N_27874,N_25161,N_25222);
nand U27875 (N_27875,N_25006,N_24818);
nand U27876 (N_27876,N_24671,N_25778);
and U27877 (N_27877,N_25004,N_24834);
nand U27878 (N_27878,N_25083,N_25273);
nand U27879 (N_27879,N_24082,N_24246);
nor U27880 (N_27880,N_25749,N_24529);
and U27881 (N_27881,N_24887,N_24417);
xor U27882 (N_27882,N_24031,N_24528);
or U27883 (N_27883,N_25873,N_24094);
and U27884 (N_27884,N_25902,N_24672);
nor U27885 (N_27885,N_25415,N_25300);
and U27886 (N_27886,N_24127,N_25431);
and U27887 (N_27887,N_25287,N_25741);
and U27888 (N_27888,N_24550,N_25556);
and U27889 (N_27889,N_25433,N_25037);
xor U27890 (N_27890,N_25235,N_24705);
nand U27891 (N_27891,N_24809,N_24817);
xor U27892 (N_27892,N_25239,N_24867);
nand U27893 (N_27893,N_25503,N_24410);
and U27894 (N_27894,N_25848,N_24209);
xnor U27895 (N_27895,N_24233,N_24119);
or U27896 (N_27896,N_24387,N_24108);
nor U27897 (N_27897,N_24494,N_24631);
nand U27898 (N_27898,N_25961,N_24961);
and U27899 (N_27899,N_24265,N_25788);
nand U27900 (N_27900,N_25028,N_24057);
xnor U27901 (N_27901,N_25596,N_24976);
xnor U27902 (N_27902,N_24180,N_24133);
or U27903 (N_27903,N_24598,N_24825);
nand U27904 (N_27904,N_24708,N_25710);
and U27905 (N_27905,N_25513,N_25329);
and U27906 (N_27906,N_25602,N_24167);
nor U27907 (N_27907,N_25836,N_25859);
or U27908 (N_27908,N_24972,N_24033);
nor U27909 (N_27909,N_24281,N_24732);
nor U27910 (N_27910,N_25893,N_24293);
nor U27911 (N_27911,N_25751,N_24750);
xor U27912 (N_27912,N_25388,N_24520);
or U27913 (N_27913,N_25430,N_24459);
or U27914 (N_27914,N_24224,N_24916);
nor U27915 (N_27915,N_25962,N_25303);
and U27916 (N_27916,N_25495,N_25442);
xnor U27917 (N_27917,N_24893,N_24669);
nor U27918 (N_27918,N_25867,N_24896);
nor U27919 (N_27919,N_24274,N_25790);
nand U27920 (N_27920,N_25806,N_25601);
xnor U27921 (N_27921,N_24073,N_25139);
nor U27922 (N_27922,N_25669,N_25455);
nor U27923 (N_27923,N_25276,N_24420);
nand U27924 (N_27924,N_24025,N_25437);
nor U27925 (N_27925,N_25847,N_24780);
nand U27926 (N_27926,N_24961,N_24296);
nor U27927 (N_27927,N_24258,N_24612);
nand U27928 (N_27928,N_24184,N_25446);
nor U27929 (N_27929,N_25152,N_24549);
nor U27930 (N_27930,N_25389,N_24484);
nor U27931 (N_27931,N_24419,N_25215);
and U27932 (N_27932,N_25018,N_24203);
nor U27933 (N_27933,N_24940,N_24774);
and U27934 (N_27934,N_25088,N_25031);
xor U27935 (N_27935,N_25930,N_25360);
nor U27936 (N_27936,N_24478,N_24645);
nor U27937 (N_27937,N_24427,N_25539);
nor U27938 (N_27938,N_24811,N_25289);
or U27939 (N_27939,N_25364,N_25463);
or U27940 (N_27940,N_24108,N_24624);
and U27941 (N_27941,N_24614,N_25546);
xor U27942 (N_27942,N_24407,N_24574);
nand U27943 (N_27943,N_24243,N_25248);
nand U27944 (N_27944,N_25534,N_25103);
or U27945 (N_27945,N_25770,N_25868);
or U27946 (N_27946,N_25155,N_25550);
nor U27947 (N_27947,N_25571,N_24694);
and U27948 (N_27948,N_25956,N_25872);
and U27949 (N_27949,N_25768,N_25534);
and U27950 (N_27950,N_25101,N_25303);
and U27951 (N_27951,N_25849,N_24243);
and U27952 (N_27952,N_24693,N_24511);
nand U27953 (N_27953,N_24170,N_24553);
or U27954 (N_27954,N_24508,N_24110);
nand U27955 (N_27955,N_24606,N_25859);
nor U27956 (N_27956,N_25098,N_24337);
or U27957 (N_27957,N_25558,N_25130);
nor U27958 (N_27958,N_25304,N_24070);
nand U27959 (N_27959,N_25233,N_25903);
or U27960 (N_27960,N_24772,N_24808);
nand U27961 (N_27961,N_25512,N_25847);
nand U27962 (N_27962,N_24136,N_24024);
nand U27963 (N_27963,N_24340,N_25015);
or U27964 (N_27964,N_24949,N_24712);
and U27965 (N_27965,N_24122,N_24665);
or U27966 (N_27966,N_24505,N_24758);
xor U27967 (N_27967,N_25108,N_25860);
nor U27968 (N_27968,N_24559,N_24988);
nor U27969 (N_27969,N_25636,N_24988);
nor U27970 (N_27970,N_24497,N_24577);
xnor U27971 (N_27971,N_25321,N_24715);
xnor U27972 (N_27972,N_24098,N_24206);
nor U27973 (N_27973,N_24651,N_25217);
and U27974 (N_27974,N_25637,N_25809);
or U27975 (N_27975,N_24989,N_24340);
nand U27976 (N_27976,N_25877,N_25105);
or U27977 (N_27977,N_24355,N_25652);
nand U27978 (N_27978,N_24726,N_24661);
and U27979 (N_27979,N_25803,N_25868);
xor U27980 (N_27980,N_25044,N_25988);
or U27981 (N_27981,N_24285,N_25336);
nor U27982 (N_27982,N_25737,N_25421);
xnor U27983 (N_27983,N_24213,N_25451);
nor U27984 (N_27984,N_25948,N_25129);
xor U27985 (N_27985,N_25884,N_25131);
or U27986 (N_27986,N_24193,N_24649);
xnor U27987 (N_27987,N_25685,N_24928);
nor U27988 (N_27988,N_24762,N_24399);
or U27989 (N_27989,N_25133,N_25371);
nor U27990 (N_27990,N_25436,N_25172);
and U27991 (N_27991,N_25276,N_24388);
xnor U27992 (N_27992,N_24839,N_24030);
or U27993 (N_27993,N_24740,N_25722);
and U27994 (N_27994,N_25511,N_25954);
nand U27995 (N_27995,N_25832,N_24372);
or U27996 (N_27996,N_24086,N_24060);
nand U27997 (N_27997,N_25189,N_24605);
nor U27998 (N_27998,N_25807,N_24843);
nand U27999 (N_27999,N_25307,N_24132);
nand U28000 (N_28000,N_26760,N_26083);
or U28001 (N_28001,N_26017,N_27337);
and U28002 (N_28002,N_26196,N_26957);
or U28003 (N_28003,N_26146,N_26874);
or U28004 (N_28004,N_27178,N_26549);
xnor U28005 (N_28005,N_27701,N_26664);
nand U28006 (N_28006,N_26561,N_26851);
nand U28007 (N_28007,N_27738,N_26013);
and U28008 (N_28008,N_26216,N_26953);
xnor U28009 (N_28009,N_27101,N_26456);
nor U28010 (N_28010,N_26705,N_27276);
and U28011 (N_28011,N_27064,N_27507);
and U28012 (N_28012,N_26039,N_27732);
or U28013 (N_28013,N_26995,N_27857);
xnor U28014 (N_28014,N_27791,N_27497);
or U28015 (N_28015,N_27348,N_27063);
nand U28016 (N_28016,N_26623,N_27242);
nand U28017 (N_28017,N_26562,N_27524);
and U28018 (N_28018,N_27047,N_26936);
nor U28019 (N_28019,N_26527,N_26532);
or U28020 (N_28020,N_26053,N_27014);
or U28021 (N_28021,N_26949,N_26708);
or U28022 (N_28022,N_27926,N_27071);
nor U28023 (N_28023,N_27540,N_26704);
xnor U28024 (N_28024,N_26648,N_27457);
xor U28025 (N_28025,N_26480,N_26076);
nor U28026 (N_28026,N_26597,N_26344);
nand U28027 (N_28027,N_27140,N_27604);
nor U28028 (N_28028,N_26822,N_27325);
nand U28029 (N_28029,N_26087,N_27621);
nor U28030 (N_28030,N_26449,N_27870);
nor U28031 (N_28031,N_26534,N_26033);
xor U28032 (N_28032,N_27441,N_26180);
xnor U28033 (N_28033,N_27269,N_26389);
xnor U28034 (N_28034,N_26155,N_27534);
nor U28035 (N_28035,N_26903,N_27544);
nor U28036 (N_28036,N_27765,N_27702);
nor U28037 (N_28037,N_27288,N_26284);
and U28038 (N_28038,N_26699,N_27158);
or U28039 (N_28039,N_27301,N_27145);
xor U28040 (N_28040,N_26899,N_27387);
and U28041 (N_28041,N_26621,N_27032);
and U28042 (N_28042,N_27149,N_27107);
nand U28043 (N_28043,N_26917,N_26012);
nor U28044 (N_28044,N_26599,N_26864);
or U28045 (N_28045,N_26598,N_26572);
and U28046 (N_28046,N_27247,N_27517);
nor U28047 (N_28047,N_26732,N_26673);
xor U28048 (N_28048,N_27129,N_26045);
xor U28049 (N_28049,N_27662,N_27108);
and U28050 (N_28050,N_27386,N_26502);
xnor U28051 (N_28051,N_27827,N_26394);
nor U28052 (N_28052,N_26789,N_27307);
nor U28053 (N_28053,N_26674,N_27938);
nor U28054 (N_28054,N_26210,N_26361);
nor U28055 (N_28055,N_26579,N_26762);
xor U28056 (N_28056,N_27249,N_27279);
nand U28057 (N_28057,N_26072,N_26154);
or U28058 (N_28058,N_27162,N_27959);
and U28059 (N_28059,N_26927,N_26835);
or U28060 (N_28060,N_26435,N_26228);
nand U28061 (N_28061,N_27277,N_26962);
nand U28062 (N_28062,N_26318,N_27389);
xnor U28063 (N_28063,N_27576,N_27244);
nand U28064 (N_28064,N_27635,N_26776);
xor U28065 (N_28065,N_26457,N_27123);
xor U28066 (N_28066,N_26029,N_27437);
or U28067 (N_28067,N_26023,N_26236);
nor U28068 (N_28068,N_26731,N_27263);
or U28069 (N_28069,N_27718,N_26867);
and U28070 (N_28070,N_27464,N_27282);
xnor U28071 (N_28071,N_27271,N_27142);
nand U28072 (N_28072,N_27931,N_27548);
xor U28073 (N_28073,N_26245,N_27556);
and U28074 (N_28074,N_27763,N_27589);
nor U28075 (N_28075,N_26671,N_26589);
or U28076 (N_28076,N_27838,N_27020);
nand U28077 (N_28077,N_27099,N_27969);
or U28078 (N_28078,N_26861,N_26870);
and U28079 (N_28079,N_27639,N_26299);
nor U28080 (N_28080,N_27204,N_27267);
xor U28081 (N_28081,N_26031,N_26459);
nor U28082 (N_28082,N_26624,N_27550);
or U28083 (N_28083,N_26727,N_26741);
or U28084 (N_28084,N_26307,N_27953);
nor U28085 (N_28085,N_26665,N_27824);
or U28086 (N_28086,N_26571,N_27503);
or U28087 (N_28087,N_27111,N_27281);
nand U28088 (N_28088,N_26877,N_26445);
xnor U28089 (N_28089,N_27042,N_27153);
nand U28090 (N_28090,N_27316,N_26928);
and U28091 (N_28091,N_26909,N_26353);
nand U28092 (N_28092,N_26998,N_26296);
or U28093 (N_28093,N_27318,N_27382);
nor U28094 (N_28094,N_27947,N_27114);
xor U28095 (N_28095,N_26551,N_27500);
nand U28096 (N_28096,N_27211,N_27365);
and U28097 (N_28097,N_27780,N_26792);
nand U28098 (N_28098,N_26733,N_27707);
xnor U28099 (N_28099,N_26659,N_27935);
and U28100 (N_28100,N_27414,N_26988);
nand U28101 (N_28101,N_27169,N_27802);
or U28102 (N_28102,N_26439,N_27481);
and U28103 (N_28103,N_26497,N_27641);
or U28104 (N_28104,N_26696,N_26747);
nand U28105 (N_28105,N_26478,N_26518);
nor U28106 (N_28106,N_26935,N_27061);
and U28107 (N_28107,N_27504,N_26912);
or U28108 (N_28108,N_26157,N_27364);
nand U28109 (N_28109,N_26918,N_26440);
nor U28110 (N_28110,N_26043,N_27894);
and U28111 (N_28111,N_26088,N_26213);
or U28112 (N_28112,N_26565,N_27498);
or U28113 (N_28113,N_27104,N_27424);
nand U28114 (N_28114,N_26417,N_27823);
nand U28115 (N_28115,N_27186,N_26639);
xor U28116 (N_28116,N_27102,N_26186);
nor U28117 (N_28117,N_26050,N_26379);
nand U28118 (N_28118,N_26887,N_27110);
xnor U28119 (N_28119,N_27214,N_27367);
nor U28120 (N_28120,N_27274,N_26225);
nand U28121 (N_28121,N_26368,N_26377);
and U28122 (N_28122,N_26192,N_26413);
nand U28123 (N_28123,N_26484,N_26635);
and U28124 (N_28124,N_26931,N_26686);
nor U28125 (N_28125,N_26205,N_26770);
and U28126 (N_28126,N_26801,N_27744);
xnor U28127 (N_28127,N_27160,N_27484);
or U28128 (N_28128,N_27619,N_26925);
xnor U28129 (N_28129,N_27459,N_27361);
nand U28130 (N_28130,N_27817,N_26896);
and U28131 (N_28131,N_26947,N_27650);
or U28132 (N_28132,N_27860,N_26657);
xor U28133 (N_28133,N_26716,N_26193);
xor U28134 (N_28134,N_27176,N_27597);
and U28135 (N_28135,N_26488,N_27858);
and U28136 (N_28136,N_26622,N_26983);
and U28137 (N_28137,N_27516,N_26794);
nand U28138 (N_28138,N_26848,N_27036);
nor U28139 (N_28139,N_27625,N_27917);
and U28140 (N_28140,N_27353,N_27239);
and U28141 (N_28141,N_26923,N_26577);
or U28142 (N_28142,N_27351,N_26090);
or U28143 (N_28143,N_26107,N_27560);
nor U28144 (N_28144,N_27837,N_27002);
nor U28145 (N_28145,N_27687,N_26566);
xor U28146 (N_28146,N_27741,N_26952);
and U28147 (N_28147,N_26127,N_26514);
nor U28148 (N_28148,N_27322,N_27444);
xor U28149 (N_28149,N_27175,N_27596);
or U28150 (N_28150,N_26730,N_27854);
xnor U28151 (N_28151,N_27469,N_26841);
nor U28152 (N_28152,N_27254,N_26365);
and U28153 (N_28153,N_27808,N_26218);
xor U28154 (N_28154,N_27182,N_26140);
and U28155 (N_28155,N_27394,N_27486);
xnor U28156 (N_28156,N_26481,N_27167);
nand U28157 (N_28157,N_27717,N_27343);
nor U28158 (N_28158,N_26317,N_26676);
xnor U28159 (N_28159,N_26366,N_26712);
nor U28160 (N_28160,N_27742,N_26955);
xnor U28161 (N_28161,N_26474,N_26181);
nor U28162 (N_28162,N_27120,N_26486);
nor U28163 (N_28163,N_26123,N_27474);
nand U28164 (N_28164,N_26914,N_26024);
nor U28165 (N_28165,N_26150,N_27033);
xnor U28166 (N_28166,N_26086,N_26859);
nand U28167 (N_28167,N_26825,N_27373);
nor U28168 (N_28168,N_26134,N_26625);
nand U28169 (N_28169,N_27506,N_27647);
nand U28170 (N_28170,N_26616,N_26702);
nand U28171 (N_28171,N_26177,N_27831);
and U28172 (N_28172,N_26306,N_27697);
nand U28173 (N_28173,N_26901,N_27058);
nor U28174 (N_28174,N_26267,N_26424);
or U28175 (N_28175,N_26409,N_27927);
and U28176 (N_28176,N_26226,N_27374);
and U28177 (N_28177,N_27069,N_26243);
nand U28178 (N_28178,N_26349,N_27202);
or U28179 (N_28179,N_27849,N_27115);
and U28180 (N_28180,N_26994,N_27190);
and U28181 (N_28181,N_27892,N_27725);
xor U28182 (N_28182,N_26185,N_27118);
nand U28183 (N_28183,N_26465,N_26883);
nor U28184 (N_28184,N_27172,N_26726);
nand U28185 (N_28185,N_26187,N_27755);
and U28186 (N_28186,N_27347,N_27131);
nand U28187 (N_28187,N_26386,N_27406);
nor U28188 (N_28188,N_26334,N_26051);
nand U28189 (N_28189,N_27331,N_26037);
or U28190 (N_28190,N_27843,N_26278);
nand U28191 (N_28191,N_26507,N_27303);
and U28192 (N_28192,N_26373,N_27566);
xor U28193 (N_28193,N_27593,N_27180);
nor U28194 (N_28194,N_27028,N_27944);
nor U28195 (N_28195,N_26611,N_26437);
nand U28196 (N_28196,N_26725,N_26108);
xor U28197 (N_28197,N_26643,N_27358);
xor U28198 (N_28198,N_26371,N_26158);
nor U28199 (N_28199,N_27159,N_27633);
xor U28200 (N_28200,N_27308,N_27630);
xor U28201 (N_28201,N_27574,N_27585);
nand U28202 (N_28202,N_27022,N_27710);
nor U28203 (N_28203,N_26057,N_26159);
nor U28204 (N_28204,N_26764,N_26084);
or U28205 (N_28205,N_26009,N_27393);
xor U28206 (N_28206,N_26052,N_26775);
nand U28207 (N_28207,N_27914,N_26438);
or U28208 (N_28208,N_27094,N_26946);
or U28209 (N_28209,N_26554,N_26189);
or U28210 (N_28210,N_27958,N_26911);
nor U28211 (N_28211,N_27624,N_27166);
or U28212 (N_28212,N_26436,N_26504);
nor U28213 (N_28213,N_27411,N_26374);
nor U28214 (N_28214,N_26869,N_26961);
xnor U28215 (N_28215,N_26402,N_26168);
nor U28216 (N_28216,N_26836,N_27525);
and U28217 (N_28217,N_27217,N_26683);
xor U28218 (N_28218,N_26182,N_26924);
or U28219 (N_28219,N_27258,N_27005);
or U28220 (N_28220,N_26063,N_26241);
xnor U28221 (N_28221,N_26629,N_26281);
and U28222 (N_28222,N_27880,N_26717);
xor U28223 (N_28223,N_27752,N_26008);
or U28224 (N_28224,N_26746,N_27476);
nand U28225 (N_28225,N_27615,N_27181);
xnor U28226 (N_28226,N_26512,N_26685);
nor U28227 (N_28227,N_27652,N_26370);
xor U28228 (N_28228,N_27825,N_27598);
nand U28229 (N_28229,N_26410,N_27930);
xor U28230 (N_28230,N_27897,N_26425);
and U28231 (N_28231,N_27998,N_27868);
xnor U28232 (N_28232,N_27966,N_26604);
or U28233 (N_28233,N_26346,N_26384);
xor U28234 (N_28234,N_27979,N_27971);
and U28235 (N_28235,N_27019,N_26414);
nor U28236 (N_28236,N_27177,N_27888);
and U28237 (N_28237,N_27344,N_27773);
or U28238 (N_28238,N_26645,N_27026);
nand U28239 (N_28239,N_27098,N_26980);
xnor U28240 (N_28240,N_26843,N_27179);
and U28241 (N_28241,N_26420,N_26030);
xor U28242 (N_28242,N_26120,N_27762);
xor U28243 (N_28243,N_27737,N_27809);
and U28244 (N_28244,N_26845,N_26580);
and U28245 (N_28245,N_27000,N_26056);
and U28246 (N_28246,N_27851,N_26319);
nor U28247 (N_28247,N_27960,N_26412);
xnor U28248 (N_28248,N_27287,N_26133);
and U28249 (N_28249,N_27139,N_26833);
or U28250 (N_28250,N_26894,N_26007);
xnor U28251 (N_28251,N_26244,N_26526);
or U28252 (N_28252,N_26541,N_27079);
nand U28253 (N_28253,N_26498,N_27312);
nand U28254 (N_28254,N_27007,N_26838);
xor U28255 (N_28255,N_27694,N_26944);
nor U28256 (N_28256,N_26206,N_26634);
xnor U28257 (N_28257,N_26419,N_26913);
or U28258 (N_28258,N_27487,N_26965);
nand U28259 (N_28259,N_26546,N_27168);
and U28260 (N_28260,N_27943,N_27342);
xor U28261 (N_28261,N_26074,N_26173);
nor U28262 (N_28262,N_27200,N_27677);
nand U28263 (N_28263,N_26668,N_27561);
nor U28264 (N_28264,N_26954,N_26662);
nand U28265 (N_28265,N_26711,N_26508);
xor U28266 (N_28266,N_27820,N_27221);
nor U28267 (N_28267,N_27753,N_26807);
xnor U28268 (N_28268,N_26289,N_27103);
xor U28269 (N_28269,N_26477,N_26511);
xnor U28270 (N_28270,N_26336,N_26989);
nand U28271 (N_28271,N_27764,N_26695);
and U28272 (N_28272,N_27970,N_27654);
xnor U28273 (N_28273,N_26431,N_26496);
nand U28274 (N_28274,N_27488,N_26253);
and U28275 (N_28275,N_27077,N_27038);
and U28276 (N_28276,N_26866,N_27613);
and U28277 (N_28277,N_27747,N_26382);
or U28278 (N_28278,N_26203,N_27439);
nor U28279 (N_28279,N_26248,N_26416);
nand U28280 (N_28280,N_26096,N_26547);
nor U28281 (N_28281,N_26517,N_26678);
nor U28282 (N_28282,N_26658,N_27940);
nand U28283 (N_28283,N_27612,N_27573);
xor U28284 (N_28284,N_26889,N_27402);
and U28285 (N_28285,N_26058,N_26128);
xor U28286 (N_28286,N_27018,N_27017);
and U28287 (N_28287,N_27156,N_26904);
and U28288 (N_28288,N_27097,N_27196);
nor U28289 (N_28289,N_27392,N_27473);
or U28290 (N_28290,N_27495,N_27731);
nand U28291 (N_28291,N_26315,N_26006);
nor U28292 (N_28292,N_27852,N_27853);
and U28293 (N_28293,N_26609,N_27904);
xor U28294 (N_28294,N_27091,N_27578);
nor U28295 (N_28295,N_27203,N_27724);
and U28296 (N_28296,N_27674,N_26479);
nor U28297 (N_28297,N_26018,N_27531);
and U28298 (N_28298,N_26321,N_27452);
nand U28299 (N_28299,N_27642,N_27933);
nand U28300 (N_28300,N_27705,N_27499);
xor U28301 (N_28301,N_26688,N_26797);
xor U28302 (N_28302,N_26538,N_27084);
or U28303 (N_28303,N_27378,N_27683);
or U28304 (N_28304,N_26573,N_27083);
or U28305 (N_28305,N_27968,N_26646);
nor U28306 (N_28306,N_27679,N_26467);
nor U28307 (N_28307,N_27928,N_27993);
xor U28308 (N_28308,N_27266,N_26774);
and U28309 (N_28309,N_27783,N_27407);
and U28310 (N_28310,N_27834,N_27165);
or U28311 (N_28311,N_26428,N_27788);
nand U28312 (N_28312,N_27552,N_26537);
nor U28313 (N_28313,N_26804,N_26694);
and U28314 (N_28314,N_27515,N_27999);
nand U28315 (N_28315,N_27936,N_27579);
or U28316 (N_28316,N_26788,N_27434);
xnor U28317 (N_28317,N_27816,N_27082);
nand U28318 (N_28318,N_26719,N_26991);
xnor U28319 (N_28319,N_26882,N_27054);
xor U28320 (N_28320,N_26038,N_27988);
xor U28321 (N_28321,N_26047,N_27680);
xnor U28322 (N_28322,N_27896,N_27541);
nor U28323 (N_28323,N_26454,N_27768);
nand U28324 (N_28324,N_26682,N_27492);
and U28325 (N_28325,N_26908,N_26742);
or U28326 (N_28326,N_26976,N_27025);
nor U28327 (N_28327,N_26145,N_26250);
nor U28328 (N_28328,N_27046,N_27428);
nor U28329 (N_28329,N_27733,N_26888);
or U28330 (N_28330,N_27793,N_27719);
or U28331 (N_28331,N_27865,N_26089);
nor U28332 (N_28332,N_26268,N_27215);
nor U28333 (N_28333,N_26669,N_26079);
or U28334 (N_28334,N_26583,N_26391);
or U28335 (N_28335,N_27219,N_27590);
nor U28336 (N_28336,N_26523,N_27003);
and U28337 (N_28337,N_27087,N_27617);
and U28338 (N_28338,N_26892,N_26415);
nand U28339 (N_28339,N_26300,N_26290);
nor U28340 (N_28340,N_26254,N_26337);
or U28341 (N_28341,N_26879,N_26592);
nor U28342 (N_28342,N_26359,N_26171);
xnor U28343 (N_28343,N_26687,N_27250);
or U28344 (N_28344,N_26555,N_27416);
nor U28345 (N_28345,N_26430,N_27423);
or U28346 (N_28346,N_26821,N_26510);
nand U28347 (N_28347,N_27293,N_27070);
or U28348 (N_28348,N_27676,N_26650);
nand U28349 (N_28349,N_26276,N_27113);
nor U28350 (N_28350,N_27380,N_27096);
nand U28351 (N_28351,N_26900,N_27368);
or U28352 (N_28352,N_26968,N_26396);
nand U28353 (N_28353,N_26001,N_26524);
nand U28354 (N_28354,N_27774,N_26997);
nand U28355 (N_28355,N_26964,N_26846);
nor U28356 (N_28356,N_26333,N_26026);
and U28357 (N_28357,N_27682,N_27869);
nand U28358 (N_28358,N_27664,N_27568);
xnor U28359 (N_28359,N_26544,N_27833);
nand U28360 (N_28360,N_26766,N_26427);
or U28361 (N_28361,N_27886,N_26633);
and U28362 (N_28362,N_27268,N_26692);
xnor U28363 (N_28363,N_26802,N_27466);
nor U28364 (N_28364,N_26945,N_27876);
and U28365 (N_28365,N_26470,N_26138);
xor U28366 (N_28366,N_27882,N_26455);
or U28367 (N_28367,N_27745,N_27209);
nor U28368 (N_28368,N_27171,N_27235);
nor U28369 (N_28369,N_26941,N_27264);
and U28370 (N_28370,N_26104,N_27794);
xor U28371 (N_28371,N_26596,N_27629);
nor U28372 (N_28372,N_26743,N_27784);
nand U28373 (N_28373,N_27907,N_26816);
xor U28374 (N_28374,N_27004,N_26264);
and U28375 (N_28375,N_26765,N_26356);
or U28376 (N_28376,N_27781,N_27405);
nor U28377 (N_28377,N_26197,N_26125);
nand U28378 (N_28378,N_27133,N_26049);
or U28379 (N_28379,N_26109,N_27813);
or U28380 (N_28380,N_26034,N_27921);
or U28381 (N_28381,N_26463,N_27822);
or U28382 (N_28382,N_26175,N_26291);
nand U28383 (N_28383,N_27125,N_26839);
or U28384 (N_28384,N_26447,N_27422);
and U28385 (N_28385,N_27841,N_26570);
nor U28386 (N_28386,N_27826,N_27564);
and U28387 (N_28387,N_26608,N_27449);
xor U28388 (N_28388,N_27357,N_27366);
nand U28389 (N_28389,N_27323,N_26048);
and U28390 (N_28390,N_27539,N_26885);
xor U28391 (N_28391,N_27317,N_26921);
and U28392 (N_28392,N_26491,N_26160);
and U28393 (N_28393,N_26019,N_27805);
xnor U28394 (N_28394,N_27119,N_27299);
nor U28395 (N_28395,N_27549,N_27345);
or U28396 (N_28396,N_26352,N_26853);
and U28397 (N_28397,N_26475,N_27212);
or U28398 (N_28398,N_26626,N_26602);
or U28399 (N_28399,N_27623,N_26933);
xor U28400 (N_28400,N_26505,N_27126);
or U28401 (N_28401,N_26993,N_27643);
nor U28402 (N_28402,N_26973,N_27475);
xnor U28403 (N_28403,N_27977,N_26636);
and U28404 (N_28404,N_27404,N_27163);
nand U28405 (N_28405,N_27313,N_26693);
nor U28406 (N_28406,N_26871,N_26316);
xor U28407 (N_28407,N_27611,N_26385);
xor U28408 (N_28408,N_26640,N_26661);
nand U28409 (N_28409,N_27463,N_27844);
nand U28410 (N_28410,N_26323,N_27272);
xnor U28411 (N_28411,N_26808,N_27489);
xor U28412 (N_28412,N_26355,N_26651);
nand U28413 (N_28413,N_26690,N_26081);
and U28414 (N_28414,N_26458,N_27432);
nor U28415 (N_28415,N_27779,N_26509);
and U28416 (N_28416,N_26002,N_27906);
xor U28417 (N_28417,N_27532,N_26530);
nand U28418 (N_28418,N_27726,N_27972);
nor U28419 (N_28419,N_27758,N_27207);
nor U28420 (N_28420,N_27305,N_26521);
xor U28421 (N_28421,N_26920,N_26347);
or U28422 (N_28422,N_26884,N_27134);
and U28423 (N_28423,N_26073,N_27385);
xor U28424 (N_28424,N_27902,N_27632);
xnor U28425 (N_28425,N_27285,N_26204);
xnor U28426 (N_28426,N_27379,N_27908);
or U28427 (N_28427,N_26363,N_27349);
nand U28428 (N_28428,N_27418,N_26251);
nand U28429 (N_28429,N_27722,N_26441);
xnor U28430 (N_28430,N_27052,N_26466);
xor U28431 (N_28431,N_27580,N_27408);
nand U28432 (N_28432,N_27132,N_26448);
xnor U28433 (N_28433,N_27803,N_26847);
or U28434 (N_28434,N_26684,N_26429);
nand U28435 (N_28435,N_27112,N_26151);
or U28436 (N_28436,N_27651,N_26567);
and U28437 (N_28437,N_26338,N_26040);
nor U28438 (N_28438,N_27105,N_26576);
or U28439 (N_28439,N_27770,N_26501);
or U28440 (N_28440,N_26591,N_27521);
and U28441 (N_28441,N_26397,N_26274);
nor U28442 (N_28442,N_27522,N_26164);
xor U28443 (N_28443,N_27748,N_26938);
nand U28444 (N_28444,N_26027,N_26984);
nor U28445 (N_28445,N_27673,N_27173);
nor U28446 (N_28446,N_26721,N_27716);
nor U28447 (N_28447,N_27360,N_27270);
or U28448 (N_28448,N_26542,N_27554);
xor U28449 (N_28449,N_27045,N_27976);
xnor U28450 (N_28450,N_27567,N_27356);
nand U28451 (N_28451,N_26557,N_27117);
or U28452 (N_28452,N_27205,N_27964);
and U28453 (N_28453,N_26978,N_26375);
nand U28454 (N_28454,N_27789,N_26071);
nand U28455 (N_28455,N_27609,N_27340);
nand U28456 (N_28456,N_27700,N_26085);
xnor U28457 (N_28457,N_27146,N_26139);
nor U28458 (N_28458,N_26630,N_26288);
and U28459 (N_28459,N_27605,N_27206);
or U28460 (N_28460,N_27640,N_27995);
or U28461 (N_28461,N_26793,N_27135);
or U28462 (N_28462,N_26890,N_26055);
nand U28463 (N_28463,N_27950,N_27918);
xnor U28464 (N_28464,N_27245,N_27261);
or U28465 (N_28465,N_26610,N_26806);
xor U28466 (N_28466,N_27542,N_27646);
or U28467 (N_28467,N_27248,N_26649);
and U28468 (N_28468,N_26990,N_26387);
nand U28469 (N_28469,N_26405,N_26032);
and U28470 (N_28470,N_27193,N_26569);
nand U28471 (N_28471,N_27955,N_27213);
or U28472 (N_28472,N_27796,N_27297);
nand U28473 (N_28473,N_26313,N_27199);
and U28474 (N_28474,N_26966,N_26117);
or U28475 (N_28475,N_26540,N_27284);
or U28476 (N_28476,N_26985,N_26285);
and U28477 (N_28477,N_27031,N_26752);
nand U28478 (N_28478,N_26293,N_27924);
or U28479 (N_28479,N_27067,N_26700);
xor U28480 (N_28480,N_27538,N_27100);
xnor U28481 (N_28481,N_27769,N_27335);
nand U28482 (N_28482,N_27138,N_27006);
or U28483 (N_28483,N_27910,N_27581);
nor U28484 (N_28484,N_27300,N_27814);
xnor U28485 (N_28485,N_26873,N_26823);
or U28486 (N_28486,N_26758,N_26860);
or U28487 (N_28487,N_26209,N_27874);
nand U28488 (N_28488,N_27577,N_27470);
or U28489 (N_28489,N_27986,N_26817);
and U28490 (N_28490,N_26574,N_26691);
and U28491 (N_28491,N_27900,N_26739);
xnor U28492 (N_28492,N_26443,N_26273);
or U28493 (N_28493,N_26485,N_27872);
or U28494 (N_28494,N_27638,N_27934);
nor U28495 (N_28495,N_26309,N_26826);
nor U28496 (N_28496,N_26784,N_26595);
xnor U28497 (N_28497,N_26679,N_27866);
xnor U28498 (N_28498,N_26112,N_27491);
and U28499 (N_28499,N_26715,N_26898);
and U28500 (N_28500,N_26229,N_27759);
and U28501 (N_28501,N_27819,N_27903);
and U28502 (N_28502,N_26720,N_27607);
or U28503 (N_28503,N_26269,N_27148);
and U28504 (N_28504,N_26718,N_27218);
or U28505 (N_28505,N_27050,N_27743);
nand U28506 (N_28506,N_27410,N_27399);
and U28507 (N_28507,N_26750,N_26618);
nand U28508 (N_28508,N_26855,N_27571);
nand U28509 (N_28509,N_26584,N_26631);
xnor U28510 (N_28510,N_26824,N_27147);
nand U28511 (N_28511,N_27806,N_26099);
or U28512 (N_28512,N_26487,N_27512);
or U28513 (N_28513,N_27505,N_26943);
nand U28514 (N_28514,N_26462,N_27477);
nor U28515 (N_28515,N_26872,N_26255);
and U28516 (N_28516,N_26937,N_26876);
nor U28517 (N_28517,N_26606,N_27426);
nor U28518 (N_28518,N_26422,N_27291);
and U28519 (N_28519,N_27734,N_26211);
xor U28520 (N_28520,N_26963,N_26638);
and U28521 (N_28521,N_27137,N_27945);
and U28522 (N_28522,N_26744,N_27957);
nor U28523 (N_28523,N_26813,N_27714);
xnor U28524 (N_28524,N_27925,N_27314);
or U28525 (N_28525,N_26383,N_27260);
nand U28526 (N_28526,N_26940,N_27812);
or U28527 (N_28527,N_27842,N_26230);
or U28528 (N_28528,N_27397,N_26653);
or U28529 (N_28529,N_26531,N_27231);
nand U28530 (N_28530,N_26376,N_27983);
nor U28531 (N_28531,N_27893,N_26393);
nand U28532 (N_28532,N_27328,N_27065);
xor U28533 (N_28533,N_26301,N_26221);
nand U28534 (N_28534,N_27161,N_27257);
and U28535 (N_28535,N_27878,N_27233);
xnor U28536 (N_28536,N_26810,N_27591);
nand U28537 (N_28537,N_27425,N_27839);
or U28538 (N_28538,N_26620,N_27222);
nand U28539 (N_28539,N_27320,N_27879);
nand U28540 (N_28540,N_27551,N_26582);
nor U28541 (N_28541,N_26280,N_27447);
and U28542 (N_28542,N_27543,N_26298);
nor U28543 (N_28543,N_26070,N_27772);
nand U28544 (N_28544,N_26489,N_27223);
or U28545 (N_28545,N_26992,N_26875);
nor U28546 (N_28546,N_26796,N_27599);
nor U28547 (N_28547,N_26246,N_27396);
or U28548 (N_28548,N_26198,N_27730);
and U28549 (N_28549,N_26348,N_26709);
nand U28550 (N_28550,N_26680,N_27309);
xnor U28551 (N_28551,N_26539,N_27136);
and U28552 (N_28552,N_27756,N_27355);
and U28553 (N_28553,N_26840,N_26644);
and U28554 (N_28554,N_26232,N_27363);
and U28555 (N_28555,N_26654,N_27056);
nand U28556 (N_28556,N_26600,N_27354);
or U28557 (N_28557,N_26520,N_27592);
or U28558 (N_28558,N_26220,N_27723);
xnor U28559 (N_28559,N_27709,N_27255);
or U28560 (N_28560,N_26106,N_26147);
nand U28561 (N_28561,N_27513,N_27602);
nand U28562 (N_28562,N_26078,N_27419);
or U28563 (N_28563,N_27889,N_26830);
and U28564 (N_28564,N_26627,N_26303);
and U28565 (N_28565,N_26753,N_27594);
nor U28566 (N_28566,N_26722,N_26929);
xnor U28567 (N_28567,N_26261,N_26044);
or U28568 (N_28568,N_27669,N_26310);
or U28569 (N_28569,N_26101,N_27433);
xnor U28570 (N_28570,N_26000,N_26543);
and U28571 (N_28571,N_27736,N_27403);
nor U28572 (N_28572,N_26358,N_27703);
nand U28573 (N_28573,N_26194,N_26380);
nand U28574 (N_28574,N_27949,N_26442);
and U28575 (N_28575,N_27174,N_26503);
or U28576 (N_28576,N_27618,N_26141);
xnor U28577 (N_28577,N_26324,N_27545);
and U28578 (N_28578,N_27610,N_26868);
nor U28579 (N_28579,N_26844,N_27339);
nor U28580 (N_28580,N_27514,N_27040);
nor U28581 (N_28581,N_26647,N_26996);
nand U28582 (N_28582,N_27699,N_27659);
nand U28583 (N_28583,N_27997,N_26115);
and U28584 (N_28584,N_27315,N_27197);
or U28585 (N_28585,N_27124,N_27081);
nor U28586 (N_28586,N_27013,N_27915);
nand U28587 (N_28587,N_27572,N_26490);
and U28588 (N_28588,N_27068,N_26670);
and U28589 (N_28589,N_26433,N_27066);
or U28590 (N_28590,N_27273,N_27471);
nor U28591 (N_28591,N_27089,N_26362);
and U28592 (N_28592,N_26003,N_26237);
nand U28593 (N_28593,N_26460,N_27846);
nor U28594 (N_28594,N_26723,N_27757);
xor U28595 (N_28595,N_27413,N_26062);
and U28596 (N_28596,N_27383,N_27729);
xor U28597 (N_28597,N_26060,N_27338);
nand U28598 (N_28598,N_27708,N_27051);
or U28599 (N_28599,N_26381,N_26240);
and U28600 (N_28600,N_27688,N_26666);
xnor U28601 (N_28601,N_27989,N_27559);
nor U28602 (N_28602,N_26224,N_26262);
nor U28603 (N_28603,N_26897,N_26811);
nand U28604 (N_28604,N_27790,N_26710);
and U28605 (N_28605,N_27251,N_27076);
nor U28606 (N_28606,N_27109,N_27400);
and U28607 (N_28607,N_26880,N_26585);
nor U28608 (N_28608,N_26129,N_27622);
or U28609 (N_28609,N_26343,N_27649);
nand U28610 (N_28610,N_27587,N_26357);
nor U28611 (N_28611,N_27533,N_26239);
or U28612 (N_28612,N_26805,N_27760);
and U28613 (N_28613,N_27384,N_26578);
xor U28614 (N_28614,N_27985,N_27994);
xnor U28615 (N_28615,N_27653,N_26075);
and U28616 (N_28616,N_26818,N_26471);
nor U28617 (N_28617,N_27750,N_26322);
or U28618 (N_28618,N_27230,N_27391);
and U28619 (N_28619,N_26714,N_27294);
or U28620 (N_28620,N_26588,N_27436);
and U28621 (N_28621,N_26215,N_26305);
nand U28622 (N_28622,N_27238,N_26163);
xor U28623 (N_28623,N_27240,N_26736);
xnor U28624 (N_28624,N_26388,N_26506);
nand U28625 (N_28625,N_26190,N_26827);
nand U28626 (N_28626,N_27863,N_26910);
and U28627 (N_28627,N_27446,N_26905);
xor U28628 (N_28628,N_27801,N_26701);
and U28629 (N_28629,N_26513,N_26025);
nor U28630 (N_28630,N_27073,N_27728);
xor U28631 (N_28631,N_27085,N_26516);
xor U28632 (N_28632,N_27275,N_26956);
or U28633 (N_28633,N_26856,N_26932);
nor U28634 (N_28634,N_26091,N_26314);
nand U28635 (N_28635,N_27782,N_26103);
or U28636 (N_28636,N_26950,N_27799);
nor U28637 (N_28637,N_27965,N_27627);
nor U28638 (N_28638,N_26986,N_27128);
nand U28639 (N_28639,N_27427,N_26862);
nand U28640 (N_28640,N_26259,N_26097);
and U28641 (N_28641,N_27398,N_26282);
nand U28642 (N_28642,N_26783,N_26642);
xor U28643 (N_28643,N_27092,N_26041);
or U28644 (N_28644,N_26556,N_27555);
or U28645 (N_28645,N_27749,N_27319);
nor U28646 (N_28646,N_26907,N_26834);
or U28647 (N_28647,N_27535,N_27448);
nor U28648 (N_28648,N_26790,N_26082);
xnor U28649 (N_28649,N_27234,N_27246);
and U28650 (N_28650,N_26335,N_26757);
xor U28651 (N_28651,N_26167,N_27987);
or U28652 (N_28652,N_27375,N_27144);
or U28653 (N_28653,N_27528,N_27048);
or U28654 (N_28654,N_26401,N_26494);
xor U28655 (N_28655,N_26934,N_27053);
xnor U28656 (N_28656,N_27152,N_26751);
nor U28657 (N_28657,N_26587,N_26522);
or U28658 (N_28658,N_27563,N_26558);
or U28659 (N_28659,N_27848,N_27982);
and U28660 (N_28660,N_27057,N_26552);
nand U28661 (N_28661,N_26028,N_27027);
or U28662 (N_28662,N_27043,N_26828);
nor U28663 (N_28663,N_26706,N_27867);
and U28664 (N_28664,N_27429,N_27116);
and U28665 (N_28665,N_27951,N_27981);
nor U28666 (N_28666,N_26672,N_27520);
or U28667 (N_28667,N_26891,N_27438);
xor U28668 (N_28668,N_26729,N_26858);
xnor U28669 (N_28669,N_27302,N_27035);
nand U28670 (N_28670,N_26948,N_26265);
and U28671 (N_28671,N_26779,N_27151);
xor U28672 (N_28672,N_26283,N_27243);
and U28673 (N_28673,N_27766,N_27569);
xnor U28674 (N_28674,N_26119,N_26919);
or U28675 (N_28675,N_27606,N_27795);
xnor U28676 (N_28676,N_27792,N_27530);
and U28677 (N_28677,N_26327,N_27895);
nand U28678 (N_28678,N_27037,N_27586);
nand U28679 (N_28679,N_27671,N_26734);
xor U28680 (N_28680,N_26195,N_26100);
or U28681 (N_28681,N_27324,N_26713);
and U28682 (N_28682,N_27290,N_27929);
xnor U28683 (N_28683,N_26930,N_26242);
xnor U28684 (N_28684,N_26094,N_27616);
xnor U28685 (N_28685,N_27696,N_26656);
nand U28686 (N_28686,N_27485,N_27637);
and U28687 (N_28687,N_26325,N_27106);
or U28688 (N_28688,N_26095,N_27381);
nand U28689 (N_28689,N_26594,N_27376);
and U28690 (N_28690,N_27804,N_27746);
or U28691 (N_28691,N_27456,N_27442);
xor U28692 (N_28692,N_27821,N_26768);
or U28693 (N_28693,N_27835,N_26863);
xnor U28694 (N_28694,N_27948,N_27735);
xor U28695 (N_28695,N_26340,N_27078);
and U28696 (N_28696,N_27656,N_27445);
nor U28697 (N_28697,N_26131,N_27686);
and U28698 (N_28698,N_27310,N_26975);
nor U28699 (N_28699,N_26227,N_26607);
nor U28700 (N_28700,N_27283,N_27015);
xor U28701 (N_28701,N_27600,N_27901);
xor U28702 (N_28702,N_26418,N_26372);
nand U28703 (N_28703,N_26011,N_26550);
nor U28704 (N_28704,N_27891,N_26234);
or U28705 (N_28705,N_27881,N_26113);
and U28706 (N_28706,N_27334,N_27226);
or U28707 (N_28707,N_26791,N_27786);
and U28708 (N_28708,N_26005,N_27628);
and U28709 (N_28709,N_26785,N_27460);
nand U28710 (N_28710,N_26148,N_27519);
nand U28711 (N_28711,N_27864,N_27939);
or U28712 (N_28712,N_26559,N_26972);
nand U28713 (N_28713,N_27295,N_26341);
nor U28714 (N_28714,N_26184,N_27963);
xnor U28715 (N_28715,N_27201,N_26046);
or U28716 (N_28716,N_26495,N_26453);
and U28717 (N_28717,N_26367,N_27899);
nor U28718 (N_28718,N_27996,N_27232);
nand U28719 (N_28719,N_26423,N_27252);
xor U28720 (N_28720,N_27761,N_27684);
xor U28721 (N_28721,N_26500,N_27916);
or U28722 (N_28722,N_26067,N_27009);
nand U28723 (N_28723,N_26328,N_26886);
xor U28724 (N_28724,N_26111,N_27690);
nand U28725 (N_28725,N_27450,N_26426);
and U28726 (N_28726,N_26987,N_27044);
and U28727 (N_28727,N_26021,N_27298);
nand U28728 (N_28728,N_27810,N_26400);
xor U28729 (N_28729,N_27911,N_26902);
and U28730 (N_28730,N_26850,N_26350);
nor U28731 (N_28731,N_27721,N_27648);
or U28732 (N_28732,N_26320,N_27154);
or U28733 (N_28733,N_26548,N_27060);
nand U28734 (N_28734,N_27187,N_27798);
xnor U28735 (N_28735,N_26403,N_26812);
nor U28736 (N_28736,N_27636,N_26165);
or U28737 (N_28737,N_27509,N_26832);
nand U28738 (N_28738,N_26004,N_27562);
xor U28739 (N_28739,N_27890,N_26260);
or U28740 (N_28740,N_27847,N_27713);
xnor U28741 (N_28741,N_26408,N_26110);
nor U28742 (N_28742,N_27468,N_27483);
nand U28743 (N_28743,N_26444,N_27195);
and U28744 (N_28744,N_27237,N_27458);
nand U28745 (N_28745,N_27229,N_27304);
nand U28746 (N_28746,N_26042,N_26476);
nor U28747 (N_28747,N_26249,N_27194);
and U28748 (N_28748,N_27584,N_27455);
and U28749 (N_28749,N_27941,N_27130);
nand U28750 (N_28750,N_27435,N_27286);
nor U28751 (N_28751,N_26728,N_27754);
or U28752 (N_28752,N_26201,N_26767);
xor U28753 (N_28753,N_27157,N_26951);
and U28754 (N_28754,N_27191,N_26178);
or U28755 (N_28755,N_27508,N_27336);
and U28756 (N_28756,N_27691,N_27828);
and U28757 (N_28757,N_27787,N_26342);
or U28758 (N_28758,N_27327,N_26533);
xor U28759 (N_28759,N_26772,N_27660);
and U28760 (N_28760,N_27832,N_27875);
and U28761 (N_28761,N_26312,N_26208);
xor U28762 (N_28762,N_27440,N_26122);
nand U28763 (N_28763,N_27962,N_26593);
nand U28764 (N_28764,N_27075,N_27990);
nor U28765 (N_28765,N_27510,N_26294);
or U28766 (N_28766,N_27785,N_27644);
nor U28767 (N_28767,N_27672,N_27967);
or U28768 (N_28768,N_26446,N_27421);
or U28769 (N_28769,N_26326,N_26660);
xor U28770 (N_28770,N_27420,N_27919);
nor U28771 (N_28771,N_27198,N_27974);
nand U28772 (N_28772,N_27884,N_27634);
or U28773 (N_28773,N_26360,N_27980);
xnor U28774 (N_28774,N_27620,N_26022);
and U28775 (N_28775,N_26737,N_26528);
and U28776 (N_28776,N_26130,N_26613);
nor U28777 (N_28777,N_27973,N_27877);
xnor U28778 (N_28778,N_27954,N_26124);
nand U28779 (N_28779,N_27453,N_27127);
nand U28780 (N_28780,N_27330,N_26499);
or U28781 (N_28781,N_27575,N_26132);
nor U28782 (N_28782,N_26093,N_27216);
and U28783 (N_28783,N_26617,N_26967);
nand U28784 (N_28784,N_27807,N_27024);
xor U28785 (N_28785,N_27923,N_26136);
nand U28786 (N_28786,N_26010,N_26054);
nand U28787 (N_28787,N_26525,N_26999);
xnor U28788 (N_28788,N_27192,N_26615);
and U28789 (N_28789,N_27236,N_27922);
nor U28790 (N_28790,N_26749,N_27346);
nand U28791 (N_28791,N_27074,N_26014);
xnor U28792 (N_28792,N_26974,N_27055);
or U28793 (N_28793,N_26563,N_27306);
xnor U28794 (N_28794,N_27333,N_26581);
or U28795 (N_28795,N_27461,N_26782);
nand U28796 (N_28796,N_26207,N_26162);
or U28797 (N_28797,N_26407,N_27631);
xor U28798 (N_28798,N_26759,N_26667);
or U28799 (N_28799,N_27482,N_26663);
nor U28800 (N_28800,N_27409,N_27332);
nand U28801 (N_28801,N_26590,N_27698);
xor U28802 (N_28802,N_27350,N_27711);
nand U28803 (N_28803,N_26369,N_26971);
or U28804 (N_28804,N_27715,N_26395);
and U28805 (N_28805,N_26781,N_27278);
or U28806 (N_28806,N_27675,N_27210);
xor U28807 (N_28807,N_26069,N_27321);
or U28808 (N_28808,N_26451,N_26803);
nand U28809 (N_28809,N_27008,N_27021);
or U28810 (N_28810,N_27678,N_26212);
and U28811 (N_28811,N_26881,N_27693);
xor U28812 (N_28812,N_27695,N_26698);
or U28813 (N_28813,N_27856,N_26179);
and U28814 (N_28814,N_26786,N_26263);
nor U28815 (N_28815,N_26780,N_27909);
nand U28816 (N_28816,N_27289,N_27546);
nor U28817 (N_28817,N_27706,N_27898);
nand U28818 (N_28818,N_26771,N_26235);
nand U28819 (N_28819,N_26345,N_26748);
or U28820 (N_28820,N_26114,N_26756);
and U28821 (N_28821,N_27241,N_26778);
or U28822 (N_28822,N_26170,N_26247);
nor U28823 (N_28823,N_26619,N_26601);
xnor U28824 (N_28824,N_27090,N_26137);
xor U28825 (N_28825,N_27462,N_26152);
nor U28826 (N_28826,N_27739,N_26258);
nor U28827 (N_28827,N_26161,N_27478);
nand U28828 (N_28828,N_26392,N_26098);
nand U28829 (N_28829,N_27704,N_26286);
and U28830 (N_28830,N_27905,N_26763);
or U28831 (N_28831,N_27871,N_26809);
nand U28832 (N_28832,N_27614,N_27143);
or U28833 (N_28833,N_27666,N_26188);
or U28834 (N_28834,N_26787,N_26219);
and U28835 (N_28835,N_27292,N_27913);
or U28836 (N_28836,N_27184,N_27296);
or U28837 (N_28837,N_26545,N_27685);
or U28838 (N_28838,N_27062,N_27778);
nand U28839 (N_28839,N_26399,N_27415);
nor U28840 (N_28840,N_26575,N_27029);
xor U28841 (N_28841,N_26800,N_27776);
xor U28842 (N_28842,N_27992,N_26755);
and U28843 (N_28843,N_27583,N_26270);
nor U28844 (N_28844,N_26330,N_26969);
nand U28845 (N_28845,N_27311,N_26831);
and U28846 (N_28846,N_26452,N_26461);
nor U28847 (N_28847,N_26837,N_27582);
xor U28848 (N_28848,N_26614,N_26536);
nor U28849 (N_28849,N_27228,N_27829);
or U28850 (N_28850,N_27352,N_27595);
or U28851 (N_28851,N_26172,N_26482);
xnor U28852 (N_28852,N_27946,N_27626);
nand U28853 (N_28853,N_27588,N_26703);
xor U28854 (N_28854,N_27359,N_26331);
xor U28855 (N_28855,N_27262,N_27978);
nor U28856 (N_28856,N_27661,N_27527);
nor U28857 (N_28857,N_26450,N_27185);
xnor U28858 (N_28858,N_27689,N_26979);
xor U28859 (N_28859,N_27093,N_26473);
nand U28860 (N_28860,N_26406,N_26515);
or U28861 (N_28861,N_26176,N_26483);
or U28862 (N_28862,N_26116,N_27164);
nor U28863 (N_28863,N_27553,N_26411);
and U28864 (N_28864,N_26958,N_27861);
nand U28865 (N_28865,N_26799,N_26149);
and U28866 (N_28866,N_27850,N_26257);
nand U28867 (N_28867,N_26773,N_26297);
nand U28868 (N_28868,N_26169,N_26080);
or U28869 (N_28869,N_26819,N_27227);
and U28870 (N_28870,N_27155,N_27665);
nand U28871 (N_28871,N_27692,N_26214);
nand U28872 (N_28872,N_26922,N_26077);
and U28873 (N_28873,N_26960,N_26852);
or U28874 (N_28874,N_26233,N_27412);
nand U28875 (N_28875,N_27727,N_26468);
nor U28876 (N_28876,N_26277,N_26404);
nand U28877 (N_28877,N_27942,N_26641);
and U28878 (N_28878,N_27558,N_27511);
xor U28879 (N_28879,N_27557,N_26529);
nor U28880 (N_28880,N_27465,N_27341);
nand U28881 (N_28881,N_26655,N_26632);
or U28882 (N_28882,N_27547,N_27859);
nor U28883 (N_28883,N_27451,N_26738);
or U28884 (N_28884,N_26560,N_27039);
nand U28885 (N_28885,N_27224,N_26329);
nand U28886 (N_28886,N_27771,N_26398);
xor U28887 (N_28887,N_27961,N_27141);
nand U28888 (N_28888,N_26020,N_26271);
nand U28889 (N_28889,N_27480,N_26144);
xnor U28890 (N_28890,N_26878,N_27188);
nand U28891 (N_28891,N_27845,N_26568);
and U28892 (N_28892,N_27401,N_26865);
nand U28893 (N_28893,N_27170,N_26135);
nor U28894 (N_28894,N_26842,N_27049);
and U28895 (N_28895,N_26798,N_26302);
nand U28896 (N_28896,N_27023,N_26390);
xnor U28897 (N_28897,N_26893,N_26761);
nand U28898 (N_28898,N_27370,N_26652);
or U28899 (N_28899,N_27526,N_26769);
nor U28900 (N_28900,N_27873,N_27658);
nand U28901 (N_28901,N_27208,N_26815);
and U28902 (N_28902,N_26183,N_26553);
and U28903 (N_28903,N_26432,N_26735);
nor U28904 (N_28904,N_26092,N_26814);
nand U28905 (N_28905,N_27645,N_26603);
xor U28906 (N_28906,N_26364,N_27490);
nand U28907 (N_28907,N_27797,N_26354);
nor U28908 (N_28908,N_27059,N_26926);
xor U28909 (N_28909,N_27800,N_26675);
and U28910 (N_28910,N_26942,N_26252);
xnor U28911 (N_28911,N_27280,N_27362);
nor U28912 (N_28912,N_26166,N_26102);
nand U28913 (N_28913,N_26064,N_26724);
and U28914 (N_28914,N_26519,N_26061);
xor U28915 (N_28915,N_27494,N_27885);
nor U28916 (N_28916,N_27265,N_26689);
nor U28917 (N_28917,N_26036,N_27417);
nand U28918 (N_28918,N_27225,N_26681);
nor U28919 (N_28919,N_27608,N_27811);
nand U28920 (N_28920,N_27472,N_26628);
and U28921 (N_28921,N_27189,N_27095);
or U28922 (N_28922,N_26677,N_26915);
and U28923 (N_28923,N_26118,N_26464);
nand U28924 (N_28924,N_26238,N_27991);
or U28925 (N_28925,N_26287,N_27121);
or U28926 (N_28926,N_27259,N_27855);
and U28927 (N_28927,N_26795,N_27001);
xor U28928 (N_28928,N_26586,N_27220);
xor U28929 (N_28929,N_26849,N_26829);
nor U28930 (N_28930,N_26754,N_27493);
nor U28931 (N_28931,N_27467,N_27720);
xnor U28932 (N_28932,N_26854,N_26121);
or U28933 (N_28933,N_27377,N_27010);
nand U28934 (N_28934,N_26707,N_26065);
or U28935 (N_28935,N_27183,N_27016);
and U28936 (N_28936,N_27712,N_27518);
nor U28937 (N_28937,N_27767,N_26016);
and U28938 (N_28938,N_27388,N_26697);
and U28939 (N_28939,N_26143,N_27034);
nor U28940 (N_28940,N_27088,N_26378);
nand U28941 (N_28941,N_26231,N_26191);
nand U28942 (N_28942,N_26059,N_26493);
or U28943 (N_28943,N_27815,N_27030);
nor U28944 (N_28944,N_27080,N_26421);
nor U28945 (N_28945,N_27086,N_27479);
nor U28946 (N_28946,N_27920,N_26126);
xor U28947 (N_28947,N_27501,N_27570);
or U28948 (N_28948,N_26035,N_26339);
nor U28949 (N_28949,N_26916,N_26202);
nand U28950 (N_28950,N_27369,N_27395);
xor U28951 (N_28951,N_27740,N_26612);
or U28952 (N_28952,N_27956,N_27371);
or U28953 (N_28953,N_26222,N_26820);
and U28954 (N_28954,N_27657,N_26981);
nand U28955 (N_28955,N_26351,N_26492);
or U28956 (N_28956,N_27862,N_26066);
nand U28957 (N_28957,N_27751,N_26332);
xor U28958 (N_28958,N_27670,N_27668);
nor U28959 (N_28959,N_27840,N_26266);
or U28960 (N_28960,N_27777,N_26857);
and U28961 (N_28961,N_26142,N_27887);
nand U28962 (N_28962,N_27937,N_27836);
and U28963 (N_28963,N_26906,N_27912);
or U28964 (N_28964,N_27529,N_26740);
xnor U28965 (N_28965,N_27329,N_26068);
and U28966 (N_28966,N_27072,N_26745);
xor U28967 (N_28967,N_26199,N_26308);
nor U28968 (N_28968,N_26977,N_26272);
or U28969 (N_28969,N_26275,N_27883);
nor U28970 (N_28970,N_26434,N_27932);
or U28971 (N_28971,N_27681,N_27603);
nand U28972 (N_28972,N_26637,N_26156);
xnor U28973 (N_28973,N_27537,N_26304);
and U28974 (N_28974,N_27536,N_26279);
nor U28975 (N_28975,N_27150,N_27390);
nand U28976 (N_28976,N_27502,N_27496);
and U28977 (N_28977,N_26564,N_27818);
nor U28978 (N_28978,N_27122,N_27012);
or U28979 (N_28979,N_26895,N_26472);
and U28980 (N_28980,N_26970,N_26295);
nand U28981 (N_28981,N_26469,N_26223);
or U28982 (N_28982,N_27430,N_26200);
nand U28983 (N_28983,N_27372,N_27041);
or U28984 (N_28984,N_26105,N_27523);
nor U28985 (N_28985,N_26959,N_26535);
xor U28986 (N_28986,N_27655,N_27326);
xor U28987 (N_28987,N_27443,N_27975);
xor U28988 (N_28988,N_27253,N_27775);
and U28989 (N_28989,N_27011,N_27601);
nand U28990 (N_28990,N_27565,N_26174);
xor U28991 (N_28991,N_27454,N_27667);
nand U28992 (N_28992,N_27431,N_26777);
nor U28993 (N_28993,N_26217,N_26605);
and U28994 (N_28994,N_27830,N_26939);
nand U28995 (N_28995,N_27984,N_27952);
xor U28996 (N_28996,N_26982,N_26153);
and U28997 (N_28997,N_27663,N_26015);
nor U28998 (N_28998,N_26256,N_26311);
nand U28999 (N_28999,N_27256,N_26292);
or U29000 (N_29000,N_26805,N_27977);
or U29001 (N_29001,N_26676,N_26186);
and U29002 (N_29002,N_26524,N_26846);
nor U29003 (N_29003,N_26687,N_26162);
xnor U29004 (N_29004,N_27003,N_26298);
nand U29005 (N_29005,N_27336,N_27617);
xnor U29006 (N_29006,N_26936,N_27916);
nor U29007 (N_29007,N_27403,N_27511);
xnor U29008 (N_29008,N_26282,N_26572);
nor U29009 (N_29009,N_26444,N_27579);
nor U29010 (N_29010,N_26425,N_27307);
nand U29011 (N_29011,N_26681,N_26104);
and U29012 (N_29012,N_27200,N_27874);
nor U29013 (N_29013,N_27793,N_27128);
xor U29014 (N_29014,N_27676,N_26374);
xor U29015 (N_29015,N_26021,N_27759);
xnor U29016 (N_29016,N_26441,N_27755);
and U29017 (N_29017,N_26609,N_27223);
and U29018 (N_29018,N_27197,N_26302);
or U29019 (N_29019,N_26438,N_27819);
or U29020 (N_29020,N_26948,N_27436);
nor U29021 (N_29021,N_26080,N_26916);
and U29022 (N_29022,N_27102,N_27605);
xnor U29023 (N_29023,N_26123,N_27571);
and U29024 (N_29024,N_27383,N_26739);
xnor U29025 (N_29025,N_26685,N_26438);
and U29026 (N_29026,N_27489,N_26262);
nor U29027 (N_29027,N_26943,N_27890);
nor U29028 (N_29028,N_26525,N_27300);
and U29029 (N_29029,N_26941,N_26672);
nor U29030 (N_29030,N_26369,N_26347);
and U29031 (N_29031,N_27713,N_27163);
and U29032 (N_29032,N_27698,N_27112);
xnor U29033 (N_29033,N_27965,N_26664);
xnor U29034 (N_29034,N_26755,N_26937);
xnor U29035 (N_29035,N_26531,N_27244);
xor U29036 (N_29036,N_26784,N_26467);
nand U29037 (N_29037,N_26991,N_27273);
xor U29038 (N_29038,N_26835,N_26637);
and U29039 (N_29039,N_26885,N_26209);
nand U29040 (N_29040,N_27119,N_26964);
xnor U29041 (N_29041,N_27984,N_26441);
nor U29042 (N_29042,N_26343,N_26652);
and U29043 (N_29043,N_27089,N_26567);
or U29044 (N_29044,N_26389,N_27713);
or U29045 (N_29045,N_27689,N_27991);
or U29046 (N_29046,N_27254,N_26370);
xnor U29047 (N_29047,N_27609,N_27170);
and U29048 (N_29048,N_27634,N_26460);
xnor U29049 (N_29049,N_26088,N_26419);
or U29050 (N_29050,N_26460,N_26314);
or U29051 (N_29051,N_27633,N_26841);
xor U29052 (N_29052,N_27068,N_26330);
xnor U29053 (N_29053,N_26940,N_27536);
or U29054 (N_29054,N_27057,N_27075);
nor U29055 (N_29055,N_26501,N_26055);
or U29056 (N_29056,N_26113,N_27791);
nand U29057 (N_29057,N_26241,N_27724);
xnor U29058 (N_29058,N_26581,N_26269);
nand U29059 (N_29059,N_27916,N_26039);
nand U29060 (N_29060,N_26748,N_26714);
nand U29061 (N_29061,N_26198,N_26011);
or U29062 (N_29062,N_27345,N_27082);
nor U29063 (N_29063,N_26837,N_26707);
nor U29064 (N_29064,N_26678,N_27995);
nor U29065 (N_29065,N_27875,N_26594);
xor U29066 (N_29066,N_27369,N_26363);
nand U29067 (N_29067,N_27020,N_26830);
and U29068 (N_29068,N_26014,N_27180);
or U29069 (N_29069,N_26698,N_27211);
or U29070 (N_29070,N_27445,N_27678);
nand U29071 (N_29071,N_27516,N_26856);
xnor U29072 (N_29072,N_26205,N_26127);
nand U29073 (N_29073,N_27080,N_26500);
nor U29074 (N_29074,N_26139,N_26575);
and U29075 (N_29075,N_26987,N_26563);
nor U29076 (N_29076,N_27346,N_27822);
xnor U29077 (N_29077,N_27155,N_27098);
nor U29078 (N_29078,N_27883,N_27694);
nand U29079 (N_29079,N_26515,N_27616);
or U29080 (N_29080,N_27226,N_26640);
or U29081 (N_29081,N_27617,N_27091);
nand U29082 (N_29082,N_26114,N_27784);
or U29083 (N_29083,N_27553,N_27578);
or U29084 (N_29084,N_26257,N_26612);
xor U29085 (N_29085,N_27031,N_26622);
and U29086 (N_29086,N_27410,N_26785);
nand U29087 (N_29087,N_26175,N_26401);
and U29088 (N_29088,N_26860,N_27957);
and U29089 (N_29089,N_26234,N_27731);
xnor U29090 (N_29090,N_26438,N_26881);
xnor U29091 (N_29091,N_26072,N_27359);
and U29092 (N_29092,N_27885,N_26422);
or U29093 (N_29093,N_27456,N_26127);
and U29094 (N_29094,N_27195,N_26439);
and U29095 (N_29095,N_26103,N_27821);
nor U29096 (N_29096,N_26508,N_26644);
xnor U29097 (N_29097,N_26578,N_26413);
xor U29098 (N_29098,N_27583,N_27205);
and U29099 (N_29099,N_26474,N_27767);
nor U29100 (N_29100,N_27009,N_26257);
nor U29101 (N_29101,N_27661,N_26153);
or U29102 (N_29102,N_26852,N_26381);
nor U29103 (N_29103,N_27500,N_27117);
xnor U29104 (N_29104,N_26309,N_27944);
nor U29105 (N_29105,N_27815,N_27924);
nand U29106 (N_29106,N_27534,N_26004);
nand U29107 (N_29107,N_27178,N_26526);
or U29108 (N_29108,N_26534,N_27426);
nor U29109 (N_29109,N_27567,N_26233);
nand U29110 (N_29110,N_26676,N_27359);
xor U29111 (N_29111,N_27178,N_26887);
and U29112 (N_29112,N_26262,N_27641);
xnor U29113 (N_29113,N_26861,N_27528);
nand U29114 (N_29114,N_26962,N_26611);
or U29115 (N_29115,N_27050,N_27893);
and U29116 (N_29116,N_26070,N_26663);
or U29117 (N_29117,N_27570,N_26877);
nand U29118 (N_29118,N_27195,N_27271);
and U29119 (N_29119,N_27650,N_26887);
xnor U29120 (N_29120,N_26698,N_26855);
nor U29121 (N_29121,N_26609,N_27529);
and U29122 (N_29122,N_27612,N_26267);
nor U29123 (N_29123,N_27938,N_27078);
nand U29124 (N_29124,N_27849,N_26969);
nor U29125 (N_29125,N_27110,N_26772);
xnor U29126 (N_29126,N_26335,N_27949);
or U29127 (N_29127,N_27201,N_26550);
xnor U29128 (N_29128,N_27778,N_26537);
nand U29129 (N_29129,N_27682,N_26587);
and U29130 (N_29130,N_27615,N_27151);
or U29131 (N_29131,N_26046,N_27260);
nand U29132 (N_29132,N_27187,N_27377);
and U29133 (N_29133,N_26143,N_26209);
and U29134 (N_29134,N_26263,N_26417);
xor U29135 (N_29135,N_27737,N_27308);
nand U29136 (N_29136,N_27452,N_27992);
or U29137 (N_29137,N_27869,N_26975);
and U29138 (N_29138,N_27649,N_26563);
xnor U29139 (N_29139,N_26584,N_27856);
xnor U29140 (N_29140,N_26889,N_27902);
or U29141 (N_29141,N_26417,N_27529);
and U29142 (N_29142,N_27399,N_26749);
and U29143 (N_29143,N_26034,N_26378);
nor U29144 (N_29144,N_26534,N_27864);
xnor U29145 (N_29145,N_26500,N_27813);
and U29146 (N_29146,N_27552,N_27408);
xor U29147 (N_29147,N_26175,N_26213);
nand U29148 (N_29148,N_27082,N_26548);
nor U29149 (N_29149,N_26896,N_27179);
and U29150 (N_29150,N_27296,N_26928);
and U29151 (N_29151,N_26821,N_26539);
or U29152 (N_29152,N_27240,N_26372);
nor U29153 (N_29153,N_26543,N_26550);
nand U29154 (N_29154,N_26415,N_27868);
xor U29155 (N_29155,N_26476,N_27248);
xnor U29156 (N_29156,N_26151,N_27890);
nor U29157 (N_29157,N_26588,N_27930);
xor U29158 (N_29158,N_26864,N_26466);
nand U29159 (N_29159,N_26913,N_26288);
xor U29160 (N_29160,N_27426,N_27187);
and U29161 (N_29161,N_26477,N_26389);
xor U29162 (N_29162,N_27558,N_26454);
nand U29163 (N_29163,N_26101,N_26984);
and U29164 (N_29164,N_27421,N_26251);
and U29165 (N_29165,N_27798,N_27339);
xnor U29166 (N_29166,N_26051,N_27222);
xor U29167 (N_29167,N_26091,N_26221);
nand U29168 (N_29168,N_26047,N_26470);
xnor U29169 (N_29169,N_27979,N_27830);
and U29170 (N_29170,N_27091,N_26617);
nand U29171 (N_29171,N_26755,N_26336);
and U29172 (N_29172,N_27822,N_26094);
nor U29173 (N_29173,N_27665,N_26810);
nor U29174 (N_29174,N_26926,N_26636);
or U29175 (N_29175,N_27717,N_26370);
and U29176 (N_29176,N_26539,N_27566);
or U29177 (N_29177,N_27722,N_26884);
nor U29178 (N_29178,N_27004,N_27209);
and U29179 (N_29179,N_27595,N_27041);
nand U29180 (N_29180,N_27224,N_27794);
nand U29181 (N_29181,N_27266,N_26662);
or U29182 (N_29182,N_26484,N_26601);
xor U29183 (N_29183,N_26749,N_27612);
or U29184 (N_29184,N_26047,N_26895);
nand U29185 (N_29185,N_27831,N_27367);
nand U29186 (N_29186,N_26017,N_27867);
nor U29187 (N_29187,N_26464,N_27791);
or U29188 (N_29188,N_27146,N_26604);
or U29189 (N_29189,N_26231,N_26038);
nand U29190 (N_29190,N_26057,N_26442);
xnor U29191 (N_29191,N_26430,N_26040);
nor U29192 (N_29192,N_26074,N_27155);
or U29193 (N_29193,N_27968,N_26608);
xor U29194 (N_29194,N_27024,N_26652);
xor U29195 (N_29195,N_27479,N_26968);
nand U29196 (N_29196,N_27195,N_27057);
or U29197 (N_29197,N_26059,N_26711);
and U29198 (N_29198,N_27514,N_26673);
nor U29199 (N_29199,N_26886,N_26225);
nor U29200 (N_29200,N_26491,N_26518);
nand U29201 (N_29201,N_27449,N_27881);
nand U29202 (N_29202,N_26201,N_27671);
and U29203 (N_29203,N_26462,N_26971);
and U29204 (N_29204,N_26498,N_26703);
xnor U29205 (N_29205,N_27261,N_26479);
and U29206 (N_29206,N_27863,N_27532);
xor U29207 (N_29207,N_27067,N_27504);
xor U29208 (N_29208,N_27571,N_27278);
or U29209 (N_29209,N_27734,N_27165);
and U29210 (N_29210,N_26972,N_26207);
xor U29211 (N_29211,N_26292,N_27886);
nand U29212 (N_29212,N_26440,N_26961);
nor U29213 (N_29213,N_27736,N_27310);
xnor U29214 (N_29214,N_27382,N_26820);
nand U29215 (N_29215,N_27260,N_26232);
xnor U29216 (N_29216,N_27514,N_26357);
nand U29217 (N_29217,N_26732,N_26560);
nor U29218 (N_29218,N_27825,N_26819);
and U29219 (N_29219,N_26776,N_27597);
or U29220 (N_29220,N_26459,N_27416);
and U29221 (N_29221,N_26378,N_27320);
or U29222 (N_29222,N_26932,N_27137);
nand U29223 (N_29223,N_27843,N_27267);
nor U29224 (N_29224,N_27462,N_26428);
xor U29225 (N_29225,N_27001,N_27370);
or U29226 (N_29226,N_27504,N_27858);
or U29227 (N_29227,N_27354,N_27118);
xnor U29228 (N_29228,N_27588,N_27316);
nor U29229 (N_29229,N_26354,N_26271);
or U29230 (N_29230,N_27790,N_26703);
nor U29231 (N_29231,N_26293,N_27600);
nor U29232 (N_29232,N_27518,N_26783);
nor U29233 (N_29233,N_26873,N_26365);
xnor U29234 (N_29234,N_27580,N_27232);
nor U29235 (N_29235,N_27477,N_26995);
nand U29236 (N_29236,N_27807,N_26614);
and U29237 (N_29237,N_26184,N_26896);
or U29238 (N_29238,N_26099,N_27419);
and U29239 (N_29239,N_26399,N_27068);
nor U29240 (N_29240,N_27400,N_26082);
and U29241 (N_29241,N_27339,N_26833);
or U29242 (N_29242,N_27591,N_26643);
and U29243 (N_29243,N_26931,N_26624);
or U29244 (N_29244,N_27068,N_27777);
or U29245 (N_29245,N_27060,N_27578);
or U29246 (N_29246,N_26471,N_26554);
nor U29247 (N_29247,N_27246,N_26894);
nand U29248 (N_29248,N_26262,N_27344);
nor U29249 (N_29249,N_26391,N_26242);
xnor U29250 (N_29250,N_26491,N_27324);
and U29251 (N_29251,N_27232,N_26083);
and U29252 (N_29252,N_27733,N_27217);
or U29253 (N_29253,N_26771,N_26577);
and U29254 (N_29254,N_27107,N_27055);
or U29255 (N_29255,N_27045,N_27565);
nand U29256 (N_29256,N_27091,N_26539);
or U29257 (N_29257,N_26675,N_26464);
xor U29258 (N_29258,N_27413,N_26162);
nand U29259 (N_29259,N_27251,N_27746);
nand U29260 (N_29260,N_26720,N_27234);
nand U29261 (N_29261,N_27823,N_27079);
nand U29262 (N_29262,N_27989,N_27593);
or U29263 (N_29263,N_27957,N_26866);
nor U29264 (N_29264,N_26681,N_27452);
nand U29265 (N_29265,N_26551,N_27427);
or U29266 (N_29266,N_26090,N_26042);
xnor U29267 (N_29267,N_27328,N_27214);
or U29268 (N_29268,N_26046,N_26477);
or U29269 (N_29269,N_26036,N_27818);
nand U29270 (N_29270,N_27957,N_27716);
or U29271 (N_29271,N_27123,N_26904);
and U29272 (N_29272,N_27217,N_27197);
xor U29273 (N_29273,N_26316,N_26407);
nor U29274 (N_29274,N_26262,N_26814);
nand U29275 (N_29275,N_27707,N_27857);
nor U29276 (N_29276,N_27048,N_27456);
nand U29277 (N_29277,N_27880,N_26113);
nand U29278 (N_29278,N_27156,N_26179);
nor U29279 (N_29279,N_27883,N_26566);
xnor U29280 (N_29280,N_27615,N_26641);
xor U29281 (N_29281,N_27225,N_27973);
nand U29282 (N_29282,N_27307,N_27745);
xor U29283 (N_29283,N_26619,N_26384);
xnor U29284 (N_29284,N_27061,N_26998);
xor U29285 (N_29285,N_26203,N_26889);
nor U29286 (N_29286,N_26184,N_27728);
and U29287 (N_29287,N_27393,N_26106);
xor U29288 (N_29288,N_26439,N_27560);
xnor U29289 (N_29289,N_27564,N_27277);
nor U29290 (N_29290,N_27892,N_27582);
and U29291 (N_29291,N_27691,N_27589);
or U29292 (N_29292,N_27226,N_26406);
nand U29293 (N_29293,N_26148,N_27533);
xor U29294 (N_29294,N_27573,N_26043);
or U29295 (N_29295,N_26559,N_26598);
xnor U29296 (N_29296,N_26174,N_26216);
nor U29297 (N_29297,N_27063,N_27639);
and U29298 (N_29298,N_26055,N_27551);
and U29299 (N_29299,N_27512,N_27792);
or U29300 (N_29300,N_26909,N_26820);
nor U29301 (N_29301,N_26535,N_27548);
nand U29302 (N_29302,N_27390,N_27586);
nand U29303 (N_29303,N_26700,N_26937);
nand U29304 (N_29304,N_27100,N_26875);
nand U29305 (N_29305,N_27198,N_27125);
nand U29306 (N_29306,N_26204,N_26307);
nand U29307 (N_29307,N_27512,N_27666);
or U29308 (N_29308,N_26450,N_27109);
nand U29309 (N_29309,N_27230,N_27219);
or U29310 (N_29310,N_27364,N_27414);
nor U29311 (N_29311,N_26228,N_26157);
nor U29312 (N_29312,N_27783,N_27917);
xor U29313 (N_29313,N_26787,N_26619);
or U29314 (N_29314,N_27050,N_26404);
nand U29315 (N_29315,N_26075,N_27889);
or U29316 (N_29316,N_26740,N_26904);
xnor U29317 (N_29317,N_26302,N_26750);
xnor U29318 (N_29318,N_27746,N_26498);
nand U29319 (N_29319,N_26188,N_26968);
or U29320 (N_29320,N_26036,N_26076);
xnor U29321 (N_29321,N_26633,N_26489);
xor U29322 (N_29322,N_27120,N_26337);
nand U29323 (N_29323,N_27408,N_26993);
and U29324 (N_29324,N_27323,N_27788);
nand U29325 (N_29325,N_27062,N_27286);
nor U29326 (N_29326,N_26876,N_26258);
xor U29327 (N_29327,N_27261,N_27573);
or U29328 (N_29328,N_27832,N_26074);
xnor U29329 (N_29329,N_26203,N_27733);
and U29330 (N_29330,N_27437,N_26919);
nor U29331 (N_29331,N_27523,N_26831);
nor U29332 (N_29332,N_27598,N_27014);
xnor U29333 (N_29333,N_27947,N_26713);
nand U29334 (N_29334,N_27558,N_26100);
and U29335 (N_29335,N_27621,N_27000);
or U29336 (N_29336,N_27858,N_26948);
nor U29337 (N_29337,N_26196,N_27984);
nor U29338 (N_29338,N_26295,N_26751);
or U29339 (N_29339,N_27919,N_27912);
xor U29340 (N_29340,N_26280,N_26677);
nor U29341 (N_29341,N_27385,N_26212);
xor U29342 (N_29342,N_26144,N_27626);
and U29343 (N_29343,N_27236,N_27395);
nand U29344 (N_29344,N_27240,N_26040);
nor U29345 (N_29345,N_27333,N_26959);
or U29346 (N_29346,N_27429,N_26739);
nand U29347 (N_29347,N_26860,N_26107);
or U29348 (N_29348,N_26304,N_26110);
nand U29349 (N_29349,N_26766,N_26809);
or U29350 (N_29350,N_26032,N_26869);
nand U29351 (N_29351,N_27347,N_26645);
or U29352 (N_29352,N_26105,N_27986);
and U29353 (N_29353,N_26638,N_26754);
nor U29354 (N_29354,N_26509,N_27270);
or U29355 (N_29355,N_27760,N_26043);
nor U29356 (N_29356,N_27247,N_27209);
and U29357 (N_29357,N_27689,N_27512);
xor U29358 (N_29358,N_27311,N_27496);
xor U29359 (N_29359,N_26756,N_26848);
nor U29360 (N_29360,N_26663,N_27653);
and U29361 (N_29361,N_27532,N_27189);
and U29362 (N_29362,N_27199,N_27429);
nor U29363 (N_29363,N_27697,N_27540);
xor U29364 (N_29364,N_27670,N_27176);
nor U29365 (N_29365,N_27681,N_26140);
or U29366 (N_29366,N_27053,N_27074);
xor U29367 (N_29367,N_26465,N_27380);
nand U29368 (N_29368,N_26771,N_27674);
xnor U29369 (N_29369,N_27308,N_26181);
nand U29370 (N_29370,N_27177,N_26242);
or U29371 (N_29371,N_27682,N_26320);
nand U29372 (N_29372,N_27608,N_27103);
xnor U29373 (N_29373,N_26228,N_26819);
xor U29374 (N_29374,N_26034,N_27881);
xor U29375 (N_29375,N_27992,N_26281);
nand U29376 (N_29376,N_27657,N_26529);
or U29377 (N_29377,N_26883,N_27092);
xor U29378 (N_29378,N_27098,N_27040);
nand U29379 (N_29379,N_26360,N_27884);
nor U29380 (N_29380,N_27221,N_27023);
or U29381 (N_29381,N_26865,N_26694);
nor U29382 (N_29382,N_26878,N_27494);
and U29383 (N_29383,N_27237,N_27888);
nand U29384 (N_29384,N_26523,N_27520);
nor U29385 (N_29385,N_26623,N_26708);
and U29386 (N_29386,N_27818,N_27472);
or U29387 (N_29387,N_26626,N_27788);
nand U29388 (N_29388,N_27218,N_26681);
and U29389 (N_29389,N_26375,N_27445);
xnor U29390 (N_29390,N_27557,N_26009);
xnor U29391 (N_29391,N_27767,N_27883);
xor U29392 (N_29392,N_27157,N_26579);
or U29393 (N_29393,N_27414,N_26921);
xnor U29394 (N_29394,N_27548,N_26270);
nor U29395 (N_29395,N_27552,N_27450);
nor U29396 (N_29396,N_26605,N_26639);
nor U29397 (N_29397,N_26532,N_26434);
and U29398 (N_29398,N_26146,N_27056);
nand U29399 (N_29399,N_27584,N_26635);
or U29400 (N_29400,N_27658,N_26444);
nor U29401 (N_29401,N_27122,N_27287);
or U29402 (N_29402,N_26986,N_26063);
xor U29403 (N_29403,N_26831,N_27878);
nor U29404 (N_29404,N_26491,N_27831);
or U29405 (N_29405,N_27255,N_27503);
or U29406 (N_29406,N_26662,N_26714);
and U29407 (N_29407,N_26709,N_26345);
nand U29408 (N_29408,N_27257,N_27905);
and U29409 (N_29409,N_26723,N_27032);
or U29410 (N_29410,N_26166,N_27838);
and U29411 (N_29411,N_27535,N_27167);
nor U29412 (N_29412,N_26409,N_27015);
nand U29413 (N_29413,N_26135,N_26993);
xor U29414 (N_29414,N_26123,N_26584);
or U29415 (N_29415,N_27838,N_26700);
xor U29416 (N_29416,N_27505,N_27386);
nand U29417 (N_29417,N_26222,N_26350);
nand U29418 (N_29418,N_26591,N_27654);
xnor U29419 (N_29419,N_27825,N_27292);
or U29420 (N_29420,N_26650,N_26598);
nor U29421 (N_29421,N_27828,N_27373);
and U29422 (N_29422,N_27002,N_27938);
xor U29423 (N_29423,N_26513,N_27646);
nor U29424 (N_29424,N_27274,N_26282);
nand U29425 (N_29425,N_27362,N_27028);
and U29426 (N_29426,N_26517,N_27388);
and U29427 (N_29427,N_26746,N_27500);
and U29428 (N_29428,N_27752,N_27146);
or U29429 (N_29429,N_26098,N_27187);
and U29430 (N_29430,N_27491,N_27418);
and U29431 (N_29431,N_27048,N_26673);
or U29432 (N_29432,N_26038,N_26770);
nor U29433 (N_29433,N_27255,N_27180);
and U29434 (N_29434,N_26511,N_26270);
or U29435 (N_29435,N_26131,N_26077);
xor U29436 (N_29436,N_26136,N_26847);
nand U29437 (N_29437,N_27487,N_27389);
and U29438 (N_29438,N_26999,N_26383);
nor U29439 (N_29439,N_27490,N_27128);
nor U29440 (N_29440,N_26476,N_26957);
or U29441 (N_29441,N_26542,N_27664);
and U29442 (N_29442,N_26791,N_26175);
nand U29443 (N_29443,N_27030,N_27319);
nor U29444 (N_29444,N_27382,N_27012);
and U29445 (N_29445,N_26032,N_26684);
and U29446 (N_29446,N_27459,N_26808);
and U29447 (N_29447,N_26052,N_27150);
nor U29448 (N_29448,N_26775,N_27838);
nand U29449 (N_29449,N_26698,N_26738);
nor U29450 (N_29450,N_26054,N_27421);
nand U29451 (N_29451,N_27858,N_27350);
xor U29452 (N_29452,N_27932,N_27154);
or U29453 (N_29453,N_26611,N_26554);
nand U29454 (N_29454,N_27515,N_26409);
nor U29455 (N_29455,N_27759,N_26156);
or U29456 (N_29456,N_27849,N_27556);
nor U29457 (N_29457,N_26990,N_26432);
nor U29458 (N_29458,N_26045,N_26237);
nor U29459 (N_29459,N_27385,N_27515);
nand U29460 (N_29460,N_26285,N_26156);
and U29461 (N_29461,N_27542,N_26546);
xnor U29462 (N_29462,N_27485,N_26740);
and U29463 (N_29463,N_27008,N_26735);
nand U29464 (N_29464,N_27744,N_27136);
and U29465 (N_29465,N_26476,N_27061);
or U29466 (N_29466,N_26709,N_26926);
nor U29467 (N_29467,N_27132,N_26825);
xnor U29468 (N_29468,N_26683,N_26236);
and U29469 (N_29469,N_26850,N_27957);
nand U29470 (N_29470,N_26652,N_26921);
or U29471 (N_29471,N_27470,N_26948);
xnor U29472 (N_29472,N_27461,N_27006);
or U29473 (N_29473,N_27029,N_26592);
or U29474 (N_29474,N_27820,N_26920);
nand U29475 (N_29475,N_27804,N_26746);
xor U29476 (N_29476,N_27749,N_27832);
or U29477 (N_29477,N_26476,N_27620);
and U29478 (N_29478,N_26146,N_27820);
nor U29479 (N_29479,N_26911,N_26262);
and U29480 (N_29480,N_27942,N_27255);
nor U29481 (N_29481,N_26660,N_27433);
nand U29482 (N_29482,N_27962,N_26048);
or U29483 (N_29483,N_27324,N_26441);
or U29484 (N_29484,N_26431,N_26159);
and U29485 (N_29485,N_26918,N_27344);
or U29486 (N_29486,N_26737,N_26681);
nor U29487 (N_29487,N_27938,N_27888);
nand U29488 (N_29488,N_26477,N_26013);
xnor U29489 (N_29489,N_26419,N_27424);
and U29490 (N_29490,N_26887,N_26121);
and U29491 (N_29491,N_26773,N_26000);
nor U29492 (N_29492,N_26297,N_27790);
nor U29493 (N_29493,N_26718,N_26066);
or U29494 (N_29494,N_27765,N_27957);
nor U29495 (N_29495,N_27600,N_27930);
and U29496 (N_29496,N_26048,N_26192);
or U29497 (N_29497,N_27366,N_27922);
xnor U29498 (N_29498,N_26138,N_26075);
xnor U29499 (N_29499,N_27115,N_27269);
nor U29500 (N_29500,N_27427,N_27440);
and U29501 (N_29501,N_26734,N_26321);
nand U29502 (N_29502,N_26668,N_26463);
and U29503 (N_29503,N_27290,N_27909);
nor U29504 (N_29504,N_27698,N_27107);
and U29505 (N_29505,N_26649,N_26083);
and U29506 (N_29506,N_27758,N_27280);
nand U29507 (N_29507,N_27099,N_26627);
or U29508 (N_29508,N_26135,N_27395);
and U29509 (N_29509,N_26770,N_26424);
or U29510 (N_29510,N_27853,N_27879);
or U29511 (N_29511,N_26250,N_27534);
xor U29512 (N_29512,N_26451,N_26163);
and U29513 (N_29513,N_27082,N_26187);
or U29514 (N_29514,N_26808,N_27426);
and U29515 (N_29515,N_27043,N_27256);
nand U29516 (N_29516,N_27550,N_26641);
xnor U29517 (N_29517,N_27688,N_27259);
or U29518 (N_29518,N_27933,N_27515);
nand U29519 (N_29519,N_26941,N_27608);
xnor U29520 (N_29520,N_27881,N_27472);
xor U29521 (N_29521,N_27831,N_27212);
nand U29522 (N_29522,N_27551,N_26369);
nor U29523 (N_29523,N_26104,N_27003);
xor U29524 (N_29524,N_27689,N_27966);
nor U29525 (N_29525,N_26834,N_27006);
nand U29526 (N_29526,N_27629,N_27027);
and U29527 (N_29527,N_27316,N_26643);
nor U29528 (N_29528,N_26175,N_26337);
or U29529 (N_29529,N_26145,N_27934);
and U29530 (N_29530,N_26022,N_26313);
and U29531 (N_29531,N_26749,N_27595);
xnor U29532 (N_29532,N_27493,N_26452);
xor U29533 (N_29533,N_26532,N_27479);
xnor U29534 (N_29534,N_27460,N_27404);
nand U29535 (N_29535,N_26765,N_27446);
nor U29536 (N_29536,N_27501,N_26917);
xor U29537 (N_29537,N_26767,N_27084);
nand U29538 (N_29538,N_27065,N_26291);
xnor U29539 (N_29539,N_26362,N_26499);
nor U29540 (N_29540,N_27126,N_27429);
or U29541 (N_29541,N_26030,N_26583);
nand U29542 (N_29542,N_27840,N_27674);
xnor U29543 (N_29543,N_26977,N_26482);
xor U29544 (N_29544,N_26978,N_27338);
and U29545 (N_29545,N_27459,N_26103);
nand U29546 (N_29546,N_27954,N_26055);
or U29547 (N_29547,N_27830,N_27887);
or U29548 (N_29548,N_27189,N_27009);
nor U29549 (N_29549,N_27925,N_27227);
nor U29550 (N_29550,N_27326,N_27842);
nor U29551 (N_29551,N_27221,N_26524);
nand U29552 (N_29552,N_27386,N_26874);
xor U29553 (N_29553,N_27133,N_27954);
nor U29554 (N_29554,N_27389,N_26794);
nor U29555 (N_29555,N_27200,N_26637);
xnor U29556 (N_29556,N_26403,N_27466);
and U29557 (N_29557,N_27865,N_26417);
nand U29558 (N_29558,N_27119,N_26802);
nand U29559 (N_29559,N_27591,N_27877);
xnor U29560 (N_29560,N_26529,N_26315);
and U29561 (N_29561,N_26339,N_27905);
xor U29562 (N_29562,N_26250,N_26302);
nor U29563 (N_29563,N_27334,N_26112);
or U29564 (N_29564,N_26849,N_27224);
and U29565 (N_29565,N_26077,N_27726);
xnor U29566 (N_29566,N_26432,N_26100);
xnor U29567 (N_29567,N_27503,N_26531);
xnor U29568 (N_29568,N_26097,N_27582);
xnor U29569 (N_29569,N_27226,N_27244);
and U29570 (N_29570,N_27578,N_26456);
and U29571 (N_29571,N_27559,N_27286);
xnor U29572 (N_29572,N_27350,N_26581);
and U29573 (N_29573,N_27780,N_26615);
nor U29574 (N_29574,N_26162,N_26244);
or U29575 (N_29575,N_27932,N_27100);
nand U29576 (N_29576,N_26289,N_27225);
nand U29577 (N_29577,N_26668,N_26499);
or U29578 (N_29578,N_26389,N_26745);
nand U29579 (N_29579,N_27656,N_27951);
and U29580 (N_29580,N_27997,N_26935);
xor U29581 (N_29581,N_27393,N_27889);
xnor U29582 (N_29582,N_26437,N_26051);
xor U29583 (N_29583,N_27333,N_27581);
and U29584 (N_29584,N_26608,N_26857);
or U29585 (N_29585,N_26509,N_27467);
nand U29586 (N_29586,N_26277,N_26737);
and U29587 (N_29587,N_26157,N_27663);
xor U29588 (N_29588,N_26942,N_27928);
nor U29589 (N_29589,N_27340,N_26431);
and U29590 (N_29590,N_26139,N_26024);
nor U29591 (N_29591,N_26414,N_26657);
nor U29592 (N_29592,N_27220,N_27070);
and U29593 (N_29593,N_27084,N_26027);
and U29594 (N_29594,N_26233,N_27982);
nand U29595 (N_29595,N_27714,N_27803);
or U29596 (N_29596,N_26761,N_27448);
nand U29597 (N_29597,N_27829,N_27844);
and U29598 (N_29598,N_27604,N_26076);
nand U29599 (N_29599,N_27315,N_27948);
or U29600 (N_29600,N_27071,N_26825);
nand U29601 (N_29601,N_27974,N_26378);
nand U29602 (N_29602,N_27029,N_26576);
or U29603 (N_29603,N_26811,N_27176);
or U29604 (N_29604,N_27440,N_26242);
nor U29605 (N_29605,N_26199,N_27710);
nor U29606 (N_29606,N_27946,N_27077);
nand U29607 (N_29607,N_27890,N_26295);
and U29608 (N_29608,N_26803,N_27535);
or U29609 (N_29609,N_27308,N_27430);
and U29610 (N_29610,N_27531,N_27944);
xnor U29611 (N_29611,N_26360,N_26420);
or U29612 (N_29612,N_27937,N_27550);
nor U29613 (N_29613,N_27702,N_27207);
and U29614 (N_29614,N_27134,N_26873);
nor U29615 (N_29615,N_27696,N_26835);
or U29616 (N_29616,N_26266,N_26233);
nor U29617 (N_29617,N_27521,N_26166);
nand U29618 (N_29618,N_26783,N_26656);
and U29619 (N_29619,N_27832,N_26947);
nand U29620 (N_29620,N_26968,N_27467);
or U29621 (N_29621,N_27548,N_26308);
xor U29622 (N_29622,N_26841,N_27941);
nor U29623 (N_29623,N_26510,N_27653);
xor U29624 (N_29624,N_26992,N_27218);
nor U29625 (N_29625,N_27309,N_26839);
nand U29626 (N_29626,N_26691,N_26239);
nor U29627 (N_29627,N_27790,N_27358);
and U29628 (N_29628,N_27587,N_27305);
and U29629 (N_29629,N_26113,N_26191);
or U29630 (N_29630,N_27166,N_26691);
or U29631 (N_29631,N_26651,N_27119);
nand U29632 (N_29632,N_27806,N_27523);
nand U29633 (N_29633,N_26801,N_26896);
xnor U29634 (N_29634,N_26663,N_26518);
nor U29635 (N_29635,N_26833,N_26975);
xnor U29636 (N_29636,N_26373,N_26951);
and U29637 (N_29637,N_26542,N_26404);
and U29638 (N_29638,N_26084,N_26218);
nor U29639 (N_29639,N_26301,N_27468);
xnor U29640 (N_29640,N_27709,N_26240);
nor U29641 (N_29641,N_27339,N_26091);
or U29642 (N_29642,N_26080,N_26136);
or U29643 (N_29643,N_26225,N_26349);
nand U29644 (N_29644,N_27842,N_26099);
and U29645 (N_29645,N_27150,N_27001);
nor U29646 (N_29646,N_26133,N_26309);
xor U29647 (N_29647,N_27234,N_27160);
nand U29648 (N_29648,N_27723,N_26526);
nand U29649 (N_29649,N_26260,N_26813);
xnor U29650 (N_29650,N_26419,N_27854);
or U29651 (N_29651,N_26935,N_27725);
and U29652 (N_29652,N_26903,N_27929);
nor U29653 (N_29653,N_26547,N_26858);
xnor U29654 (N_29654,N_26715,N_27436);
nand U29655 (N_29655,N_27046,N_26182);
nand U29656 (N_29656,N_26734,N_26482);
or U29657 (N_29657,N_27034,N_26733);
nor U29658 (N_29658,N_26436,N_26273);
nor U29659 (N_29659,N_26175,N_26811);
and U29660 (N_29660,N_27793,N_26636);
nand U29661 (N_29661,N_27629,N_26569);
or U29662 (N_29662,N_26025,N_26039);
xnor U29663 (N_29663,N_26535,N_27784);
nor U29664 (N_29664,N_26662,N_26065);
or U29665 (N_29665,N_27240,N_27704);
xor U29666 (N_29666,N_27764,N_26832);
nand U29667 (N_29667,N_26255,N_26523);
and U29668 (N_29668,N_26912,N_26874);
and U29669 (N_29669,N_27505,N_27698);
and U29670 (N_29670,N_26380,N_26411);
nor U29671 (N_29671,N_26912,N_26747);
and U29672 (N_29672,N_26673,N_26631);
and U29673 (N_29673,N_26285,N_27475);
nand U29674 (N_29674,N_27722,N_26635);
or U29675 (N_29675,N_26835,N_27474);
nand U29676 (N_29676,N_26772,N_26968);
nor U29677 (N_29677,N_26877,N_27220);
xnor U29678 (N_29678,N_26633,N_27672);
nand U29679 (N_29679,N_26997,N_27845);
and U29680 (N_29680,N_27395,N_26179);
and U29681 (N_29681,N_27485,N_27818);
or U29682 (N_29682,N_27480,N_27976);
nand U29683 (N_29683,N_26203,N_26268);
nor U29684 (N_29684,N_26700,N_26138);
nand U29685 (N_29685,N_26780,N_26935);
xnor U29686 (N_29686,N_27214,N_26933);
or U29687 (N_29687,N_26500,N_27592);
xnor U29688 (N_29688,N_26616,N_26193);
xor U29689 (N_29689,N_27793,N_26959);
nand U29690 (N_29690,N_26288,N_26387);
xnor U29691 (N_29691,N_27421,N_26329);
and U29692 (N_29692,N_26852,N_26384);
xor U29693 (N_29693,N_27560,N_26379);
xor U29694 (N_29694,N_26837,N_27801);
nand U29695 (N_29695,N_26942,N_26227);
or U29696 (N_29696,N_27049,N_26484);
xnor U29697 (N_29697,N_27299,N_27492);
nor U29698 (N_29698,N_27816,N_27698);
and U29699 (N_29699,N_27050,N_27153);
nand U29700 (N_29700,N_27321,N_26187);
and U29701 (N_29701,N_27565,N_27228);
or U29702 (N_29702,N_26733,N_27906);
and U29703 (N_29703,N_27096,N_26467);
xor U29704 (N_29704,N_27047,N_27257);
xor U29705 (N_29705,N_27746,N_27792);
nand U29706 (N_29706,N_26904,N_27404);
nor U29707 (N_29707,N_27159,N_26375);
or U29708 (N_29708,N_27519,N_27645);
xnor U29709 (N_29709,N_26552,N_26159);
and U29710 (N_29710,N_27829,N_26181);
and U29711 (N_29711,N_26613,N_26138);
nand U29712 (N_29712,N_27243,N_27371);
or U29713 (N_29713,N_26915,N_26843);
or U29714 (N_29714,N_27497,N_26219);
nand U29715 (N_29715,N_26005,N_27767);
xor U29716 (N_29716,N_26280,N_27917);
xor U29717 (N_29717,N_26453,N_27991);
or U29718 (N_29718,N_27213,N_26385);
xnor U29719 (N_29719,N_26478,N_26855);
or U29720 (N_29720,N_26948,N_26358);
nand U29721 (N_29721,N_26644,N_26543);
nor U29722 (N_29722,N_27127,N_26311);
nor U29723 (N_29723,N_26152,N_26729);
nand U29724 (N_29724,N_26315,N_26395);
and U29725 (N_29725,N_27204,N_26098);
nand U29726 (N_29726,N_26032,N_27188);
nor U29727 (N_29727,N_26735,N_26822);
or U29728 (N_29728,N_27244,N_26007);
nor U29729 (N_29729,N_27601,N_26318);
xor U29730 (N_29730,N_27685,N_27989);
xor U29731 (N_29731,N_26658,N_26344);
and U29732 (N_29732,N_27698,N_27863);
or U29733 (N_29733,N_27463,N_26698);
and U29734 (N_29734,N_27179,N_26749);
nor U29735 (N_29735,N_26966,N_26376);
nor U29736 (N_29736,N_27965,N_27454);
nand U29737 (N_29737,N_27821,N_27921);
nor U29738 (N_29738,N_26243,N_26443);
nor U29739 (N_29739,N_26800,N_26340);
xor U29740 (N_29740,N_27687,N_26990);
and U29741 (N_29741,N_27157,N_26030);
nor U29742 (N_29742,N_26806,N_26333);
xnor U29743 (N_29743,N_26375,N_26350);
xor U29744 (N_29744,N_26011,N_26445);
xnor U29745 (N_29745,N_27593,N_27796);
xor U29746 (N_29746,N_26229,N_27821);
nand U29747 (N_29747,N_27711,N_27317);
nand U29748 (N_29748,N_26662,N_27937);
xor U29749 (N_29749,N_26278,N_26289);
or U29750 (N_29750,N_27487,N_27419);
nand U29751 (N_29751,N_26826,N_26662);
xor U29752 (N_29752,N_26556,N_27173);
nor U29753 (N_29753,N_27136,N_26000);
nand U29754 (N_29754,N_26060,N_26929);
or U29755 (N_29755,N_27047,N_26866);
nand U29756 (N_29756,N_27890,N_27999);
xor U29757 (N_29757,N_26079,N_27752);
nand U29758 (N_29758,N_27251,N_26907);
and U29759 (N_29759,N_26588,N_27825);
nand U29760 (N_29760,N_27010,N_27310);
nand U29761 (N_29761,N_26694,N_26915);
nor U29762 (N_29762,N_26015,N_27871);
or U29763 (N_29763,N_26816,N_26527);
and U29764 (N_29764,N_27649,N_27593);
nand U29765 (N_29765,N_27794,N_27010);
xor U29766 (N_29766,N_27385,N_27015);
and U29767 (N_29767,N_27434,N_26369);
or U29768 (N_29768,N_26965,N_27828);
xor U29769 (N_29769,N_27963,N_27105);
nor U29770 (N_29770,N_26453,N_26707);
nor U29771 (N_29771,N_26550,N_26727);
nor U29772 (N_29772,N_26023,N_27748);
nand U29773 (N_29773,N_26338,N_27671);
or U29774 (N_29774,N_26183,N_26637);
xor U29775 (N_29775,N_27643,N_27384);
nor U29776 (N_29776,N_27376,N_27952);
nand U29777 (N_29777,N_26969,N_26939);
and U29778 (N_29778,N_26457,N_26660);
nor U29779 (N_29779,N_27238,N_26313);
or U29780 (N_29780,N_26175,N_27522);
and U29781 (N_29781,N_27135,N_26645);
and U29782 (N_29782,N_26743,N_27626);
and U29783 (N_29783,N_27583,N_27459);
nor U29784 (N_29784,N_27083,N_27113);
nor U29785 (N_29785,N_27126,N_26118);
or U29786 (N_29786,N_26455,N_26280);
or U29787 (N_29787,N_27223,N_27896);
or U29788 (N_29788,N_27785,N_27295);
or U29789 (N_29789,N_26583,N_27417);
nor U29790 (N_29790,N_26583,N_27336);
and U29791 (N_29791,N_26004,N_27144);
nor U29792 (N_29792,N_26470,N_26611);
nor U29793 (N_29793,N_26272,N_27311);
nor U29794 (N_29794,N_27603,N_27877);
xnor U29795 (N_29795,N_26195,N_27253);
or U29796 (N_29796,N_27348,N_26951);
or U29797 (N_29797,N_27313,N_27683);
and U29798 (N_29798,N_26736,N_27790);
nor U29799 (N_29799,N_26763,N_26621);
and U29800 (N_29800,N_27646,N_27470);
xor U29801 (N_29801,N_27547,N_26538);
or U29802 (N_29802,N_27344,N_26649);
and U29803 (N_29803,N_27344,N_26902);
or U29804 (N_29804,N_27845,N_26004);
or U29805 (N_29805,N_26223,N_26965);
nand U29806 (N_29806,N_27319,N_26088);
nand U29807 (N_29807,N_27639,N_27860);
nor U29808 (N_29808,N_27046,N_27885);
and U29809 (N_29809,N_26720,N_27436);
xor U29810 (N_29810,N_27907,N_26784);
and U29811 (N_29811,N_26049,N_27628);
xor U29812 (N_29812,N_27055,N_27669);
nor U29813 (N_29813,N_27356,N_26521);
and U29814 (N_29814,N_27191,N_27276);
xor U29815 (N_29815,N_26315,N_27233);
and U29816 (N_29816,N_26975,N_26901);
nor U29817 (N_29817,N_27822,N_27160);
and U29818 (N_29818,N_27913,N_27459);
or U29819 (N_29819,N_27574,N_26908);
and U29820 (N_29820,N_27491,N_27730);
nor U29821 (N_29821,N_27027,N_27258);
or U29822 (N_29822,N_26964,N_27520);
and U29823 (N_29823,N_27907,N_27919);
and U29824 (N_29824,N_26777,N_27841);
nor U29825 (N_29825,N_26120,N_27282);
or U29826 (N_29826,N_27984,N_27317);
or U29827 (N_29827,N_26214,N_27336);
and U29828 (N_29828,N_27623,N_26794);
nor U29829 (N_29829,N_27746,N_27273);
xor U29830 (N_29830,N_26863,N_27589);
xor U29831 (N_29831,N_27166,N_27752);
xnor U29832 (N_29832,N_26728,N_26622);
nor U29833 (N_29833,N_27249,N_26407);
nand U29834 (N_29834,N_27067,N_27794);
nor U29835 (N_29835,N_26837,N_26046);
xnor U29836 (N_29836,N_26884,N_27063);
nand U29837 (N_29837,N_27421,N_26995);
and U29838 (N_29838,N_26645,N_26734);
xnor U29839 (N_29839,N_27578,N_26336);
or U29840 (N_29840,N_26030,N_26039);
or U29841 (N_29841,N_26664,N_27870);
xnor U29842 (N_29842,N_26142,N_27404);
or U29843 (N_29843,N_26765,N_26741);
xnor U29844 (N_29844,N_26028,N_27997);
nor U29845 (N_29845,N_26586,N_26401);
or U29846 (N_29846,N_27989,N_26885);
xnor U29847 (N_29847,N_27458,N_26538);
xor U29848 (N_29848,N_26219,N_26198);
nor U29849 (N_29849,N_27599,N_27479);
nand U29850 (N_29850,N_27904,N_27335);
nor U29851 (N_29851,N_26348,N_27749);
nand U29852 (N_29852,N_27792,N_26753);
or U29853 (N_29853,N_27217,N_26160);
xnor U29854 (N_29854,N_26865,N_27213);
and U29855 (N_29855,N_27914,N_27597);
nand U29856 (N_29856,N_26465,N_27594);
nor U29857 (N_29857,N_27630,N_27021);
and U29858 (N_29858,N_27300,N_26671);
and U29859 (N_29859,N_27517,N_26576);
or U29860 (N_29860,N_26427,N_27141);
and U29861 (N_29861,N_27269,N_27954);
xnor U29862 (N_29862,N_26402,N_26095);
nand U29863 (N_29863,N_26393,N_27058);
and U29864 (N_29864,N_27840,N_27285);
and U29865 (N_29865,N_27822,N_27151);
and U29866 (N_29866,N_27110,N_27112);
xor U29867 (N_29867,N_26652,N_27144);
or U29868 (N_29868,N_27645,N_27295);
and U29869 (N_29869,N_27839,N_27875);
xnor U29870 (N_29870,N_27304,N_27251);
nor U29871 (N_29871,N_26176,N_26525);
or U29872 (N_29872,N_27970,N_26486);
xor U29873 (N_29873,N_26938,N_27402);
nand U29874 (N_29874,N_26390,N_27055);
and U29875 (N_29875,N_27052,N_27518);
nor U29876 (N_29876,N_27497,N_27089);
nor U29877 (N_29877,N_26190,N_27611);
xor U29878 (N_29878,N_26288,N_27799);
and U29879 (N_29879,N_27309,N_27886);
xnor U29880 (N_29880,N_27958,N_27596);
nor U29881 (N_29881,N_27574,N_26768);
xnor U29882 (N_29882,N_27512,N_27811);
nor U29883 (N_29883,N_27640,N_26180);
nor U29884 (N_29884,N_26970,N_27015);
and U29885 (N_29885,N_26191,N_26212);
or U29886 (N_29886,N_27934,N_27855);
and U29887 (N_29887,N_26213,N_27527);
and U29888 (N_29888,N_26564,N_27493);
and U29889 (N_29889,N_27214,N_27069);
nand U29890 (N_29890,N_27767,N_27688);
xnor U29891 (N_29891,N_26073,N_26904);
xnor U29892 (N_29892,N_27701,N_26340);
or U29893 (N_29893,N_27919,N_27392);
nor U29894 (N_29894,N_27592,N_27893);
nor U29895 (N_29895,N_26008,N_26308);
nand U29896 (N_29896,N_26396,N_26223);
xor U29897 (N_29897,N_27313,N_27600);
and U29898 (N_29898,N_26244,N_27015);
or U29899 (N_29899,N_27572,N_26835);
and U29900 (N_29900,N_27292,N_26866);
or U29901 (N_29901,N_27207,N_27542);
nor U29902 (N_29902,N_27589,N_27105);
nor U29903 (N_29903,N_27484,N_27356);
xnor U29904 (N_29904,N_27625,N_26046);
nor U29905 (N_29905,N_27291,N_27456);
or U29906 (N_29906,N_26139,N_27698);
or U29907 (N_29907,N_27024,N_27099);
and U29908 (N_29908,N_27060,N_26921);
or U29909 (N_29909,N_26664,N_26878);
or U29910 (N_29910,N_27129,N_26921);
nor U29911 (N_29911,N_26613,N_26073);
or U29912 (N_29912,N_26061,N_26982);
xor U29913 (N_29913,N_27200,N_26353);
or U29914 (N_29914,N_26703,N_27865);
nor U29915 (N_29915,N_26926,N_27015);
nor U29916 (N_29916,N_26101,N_26611);
nand U29917 (N_29917,N_27108,N_27979);
and U29918 (N_29918,N_27160,N_27597);
or U29919 (N_29919,N_27469,N_27881);
and U29920 (N_29920,N_27564,N_27819);
and U29921 (N_29921,N_27881,N_26378);
nor U29922 (N_29922,N_26429,N_26169);
or U29923 (N_29923,N_27411,N_27492);
nand U29924 (N_29924,N_26364,N_27061);
or U29925 (N_29925,N_26791,N_26415);
and U29926 (N_29926,N_27660,N_27244);
or U29927 (N_29927,N_27051,N_27341);
and U29928 (N_29928,N_26436,N_26885);
nand U29929 (N_29929,N_26604,N_26927);
nand U29930 (N_29930,N_27942,N_26822);
nand U29931 (N_29931,N_27764,N_27402);
or U29932 (N_29932,N_26475,N_27275);
nor U29933 (N_29933,N_26894,N_27571);
or U29934 (N_29934,N_26391,N_27527);
nand U29935 (N_29935,N_27513,N_26008);
nor U29936 (N_29936,N_27844,N_26871);
xnor U29937 (N_29937,N_26280,N_27820);
or U29938 (N_29938,N_26381,N_26474);
nor U29939 (N_29939,N_27443,N_27053);
or U29940 (N_29940,N_26334,N_27592);
or U29941 (N_29941,N_26778,N_26219);
nand U29942 (N_29942,N_26790,N_27953);
xnor U29943 (N_29943,N_27343,N_26715);
nor U29944 (N_29944,N_27683,N_26848);
and U29945 (N_29945,N_26076,N_26302);
xor U29946 (N_29946,N_26839,N_26265);
nand U29947 (N_29947,N_26980,N_26048);
nand U29948 (N_29948,N_27597,N_27924);
xnor U29949 (N_29949,N_26531,N_27124);
nand U29950 (N_29950,N_26566,N_27063);
xnor U29951 (N_29951,N_26751,N_27823);
nand U29952 (N_29952,N_26098,N_26731);
or U29953 (N_29953,N_26329,N_27456);
and U29954 (N_29954,N_26594,N_27506);
or U29955 (N_29955,N_27430,N_26898);
or U29956 (N_29956,N_26008,N_26376);
nand U29957 (N_29957,N_27494,N_27605);
and U29958 (N_29958,N_26214,N_27795);
nand U29959 (N_29959,N_27853,N_26588);
nand U29960 (N_29960,N_27258,N_26904);
nand U29961 (N_29961,N_27801,N_27003);
or U29962 (N_29962,N_27084,N_26096);
nand U29963 (N_29963,N_27730,N_27747);
nor U29964 (N_29964,N_27024,N_27483);
xnor U29965 (N_29965,N_27204,N_26099);
nor U29966 (N_29966,N_27706,N_27130);
xor U29967 (N_29967,N_26277,N_27635);
and U29968 (N_29968,N_26982,N_27451);
and U29969 (N_29969,N_26978,N_27184);
nor U29970 (N_29970,N_27418,N_27605);
nand U29971 (N_29971,N_27186,N_27846);
and U29972 (N_29972,N_26467,N_27625);
nand U29973 (N_29973,N_26643,N_27113);
or U29974 (N_29974,N_26757,N_26291);
or U29975 (N_29975,N_26353,N_27587);
and U29976 (N_29976,N_27028,N_27469);
nor U29977 (N_29977,N_26110,N_26079);
nor U29978 (N_29978,N_26089,N_26325);
or U29979 (N_29979,N_26830,N_27151);
nand U29980 (N_29980,N_27875,N_27591);
nor U29981 (N_29981,N_26142,N_27373);
nand U29982 (N_29982,N_27149,N_27148);
or U29983 (N_29983,N_26958,N_26825);
nand U29984 (N_29984,N_26130,N_27910);
xor U29985 (N_29985,N_26862,N_27213);
or U29986 (N_29986,N_27951,N_27477);
or U29987 (N_29987,N_26741,N_27082);
xor U29988 (N_29988,N_27582,N_26897);
nand U29989 (N_29989,N_27630,N_27508);
xnor U29990 (N_29990,N_27358,N_26689);
and U29991 (N_29991,N_26697,N_27004);
or U29992 (N_29992,N_27900,N_27908);
nand U29993 (N_29993,N_27212,N_27504);
nand U29994 (N_29994,N_27181,N_26485);
and U29995 (N_29995,N_26628,N_27630);
or U29996 (N_29996,N_26227,N_26715);
xor U29997 (N_29997,N_27826,N_27581);
and U29998 (N_29998,N_27590,N_26622);
or U29999 (N_29999,N_26279,N_26184);
xor U30000 (N_30000,N_28566,N_29833);
nor U30001 (N_30001,N_29214,N_29960);
and U30002 (N_30002,N_28750,N_29280);
and U30003 (N_30003,N_28031,N_28667);
nand U30004 (N_30004,N_28076,N_29410);
xnor U30005 (N_30005,N_29897,N_28306);
nand U30006 (N_30006,N_28089,N_29834);
xor U30007 (N_30007,N_28477,N_28513);
or U30008 (N_30008,N_29038,N_29433);
xor U30009 (N_30009,N_29436,N_28167);
nor U30010 (N_30010,N_29297,N_28073);
nand U30011 (N_30011,N_29298,N_29689);
nor U30012 (N_30012,N_28957,N_29509);
or U30013 (N_30013,N_29781,N_28319);
xnor U30014 (N_30014,N_28449,N_29081);
or U30015 (N_30015,N_29123,N_29313);
nand U30016 (N_30016,N_29121,N_28108);
or U30017 (N_30017,N_28168,N_29392);
xnor U30018 (N_30018,N_28583,N_28123);
xnor U30019 (N_30019,N_28913,N_28180);
and U30020 (N_30020,N_29174,N_28880);
nor U30021 (N_30021,N_28453,N_28237);
nand U30022 (N_30022,N_29595,N_29534);
nand U30023 (N_30023,N_29602,N_28998);
xor U30024 (N_30024,N_28402,N_28724);
xor U30025 (N_30025,N_28025,N_28970);
and U30026 (N_30026,N_28469,N_29997);
nor U30027 (N_30027,N_28657,N_28182);
nor U30028 (N_30028,N_28706,N_28087);
and U30029 (N_30029,N_28498,N_28479);
xor U30030 (N_30030,N_28737,N_28769);
nand U30031 (N_30031,N_29265,N_28835);
nor U30032 (N_30032,N_29102,N_28542);
xor U30033 (N_30033,N_28948,N_28568);
nand U30034 (N_30034,N_28183,N_29368);
or U30035 (N_30035,N_28414,N_28050);
nand U30036 (N_30036,N_28891,N_29640);
or U30037 (N_30037,N_29959,N_28576);
and U30038 (N_30038,N_29822,N_28428);
nor U30039 (N_30039,N_29430,N_28783);
or U30040 (N_30040,N_28918,N_29893);
xnor U30041 (N_30041,N_29646,N_29562);
xnor U30042 (N_30042,N_29366,N_28877);
nand U30043 (N_30043,N_28718,N_28756);
nor U30044 (N_30044,N_29796,N_29953);
and U30045 (N_30045,N_28631,N_29309);
or U30046 (N_30046,N_28249,N_28119);
nand U30047 (N_30047,N_28458,N_28127);
and U30048 (N_30048,N_29616,N_28238);
or U30049 (N_30049,N_29262,N_28222);
nand U30050 (N_30050,N_28159,N_29921);
or U30051 (N_30051,N_28003,N_29989);
xor U30052 (N_30052,N_29348,N_29545);
xnor U30053 (N_30053,N_28501,N_29225);
nor U30054 (N_30054,N_28662,N_28446);
or U30055 (N_30055,N_28427,N_28985);
nand U30056 (N_30056,N_28005,N_29066);
and U30057 (N_30057,N_29471,N_28273);
xnor U30058 (N_30058,N_29799,N_28164);
nand U30059 (N_30059,N_28519,N_28190);
or U30060 (N_30060,N_29579,N_29944);
or U30061 (N_30061,N_29342,N_29095);
and U30062 (N_30062,N_28000,N_29065);
nand U30063 (N_30063,N_29766,N_28855);
or U30064 (N_30064,N_28023,N_28690);
nand U30065 (N_30065,N_28202,N_28457);
nor U30066 (N_30066,N_29920,N_28098);
xor U30067 (N_30067,N_28420,N_29895);
xnor U30068 (N_30068,N_28426,N_29282);
nor U30069 (N_30069,N_28949,N_29929);
and U30070 (N_30070,N_29487,N_28214);
and U30071 (N_30071,N_28010,N_29202);
xnor U30072 (N_30072,N_29301,N_28231);
nand U30073 (N_30073,N_28321,N_28215);
nor U30074 (N_30074,N_28083,N_29129);
and U30075 (N_30075,N_28523,N_29937);
and U30076 (N_30076,N_29386,N_28156);
nor U30077 (N_30077,N_29664,N_29777);
nand U30078 (N_30078,N_28613,N_28888);
or U30079 (N_30079,N_29349,N_28391);
nor U30080 (N_30080,N_29031,N_28436);
or U30081 (N_30081,N_28712,N_28324);
and U30082 (N_30082,N_28602,N_28914);
nand U30083 (N_30083,N_28042,N_28032);
nand U30084 (N_30084,N_29707,N_28879);
nor U30085 (N_30085,N_28582,N_29532);
nand U30086 (N_30086,N_29511,N_28471);
or U30087 (N_30087,N_28562,N_29802);
nand U30088 (N_30088,N_29048,N_28130);
nor U30089 (N_30089,N_29050,N_29688);
or U30090 (N_30090,N_29034,N_28377);
and U30091 (N_30091,N_28465,N_29496);
nand U30092 (N_30092,N_29155,N_29134);
or U30093 (N_30093,N_29700,N_28068);
or U30094 (N_30094,N_29200,N_28399);
xor U30095 (N_30095,N_28472,N_28822);
nand U30096 (N_30096,N_29832,N_29945);
or U30097 (N_30097,N_28497,N_28256);
and U30098 (N_30098,N_28551,N_29851);
nand U30099 (N_30099,N_28495,N_28533);
xnor U30100 (N_30100,N_28817,N_28975);
nor U30101 (N_30101,N_29837,N_28894);
nor U30102 (N_30102,N_29105,N_29561);
nand U30103 (N_30103,N_28148,N_29044);
nand U30104 (N_30104,N_28749,N_28837);
xnor U30105 (N_30105,N_29529,N_29680);
nand U30106 (N_30106,N_29100,N_28408);
or U30107 (N_30107,N_28330,N_28702);
nand U30108 (N_30108,N_28524,N_28605);
xor U30109 (N_30109,N_29866,N_28788);
nor U30110 (N_30110,N_28939,N_28419);
xnor U30111 (N_30111,N_29845,N_29933);
nor U30112 (N_30112,N_29150,N_28983);
and U30113 (N_30113,N_29938,N_28612);
xnor U30114 (N_30114,N_29489,N_29890);
xnor U30115 (N_30115,N_29423,N_28862);
and U30116 (N_30116,N_28118,N_28064);
nand U30117 (N_30117,N_28152,N_29513);
and U30118 (N_30118,N_29084,N_28536);
nand U30119 (N_30119,N_28893,N_28990);
and U30120 (N_30120,N_29619,N_28181);
and U30121 (N_30121,N_29473,N_29790);
nor U30122 (N_30122,N_29213,N_28313);
or U30123 (N_30123,N_28364,N_29152);
nor U30124 (N_30124,N_28679,N_29358);
nor U30125 (N_30125,N_28006,N_28113);
or U30126 (N_30126,N_29804,N_29935);
nor U30127 (N_30127,N_29425,N_28697);
nand U30128 (N_30128,N_29934,N_29154);
xor U30129 (N_30129,N_29363,N_29915);
or U30130 (N_30130,N_28716,N_28460);
and U30131 (N_30131,N_29958,N_28302);
nor U30132 (N_30132,N_28410,N_29432);
nand U30133 (N_30133,N_29233,N_28730);
and U30134 (N_30134,N_28384,N_29039);
xnor U30135 (N_30135,N_29465,N_29419);
xnor U30136 (N_30136,N_29306,N_28166);
xnor U30137 (N_30137,N_29228,N_29345);
xor U30138 (N_30138,N_29420,N_29889);
nor U30139 (N_30139,N_28800,N_28303);
nand U30140 (N_30140,N_29042,N_29784);
xor U30141 (N_30141,N_28579,N_28991);
and U30142 (N_30142,N_28223,N_29742);
and U30143 (N_30143,N_29830,N_29903);
xor U30144 (N_30144,N_28394,N_29658);
xor U30145 (N_30145,N_28046,N_28953);
nor U30146 (N_30146,N_28859,N_29312);
nand U30147 (N_30147,N_28857,N_28253);
nand U30148 (N_30148,N_29624,N_29885);
nand U30149 (N_30149,N_28676,N_28935);
and U30150 (N_30150,N_29584,N_29149);
nor U30151 (N_30151,N_29536,N_29782);
nor U30152 (N_30152,N_28581,N_29825);
and U30153 (N_30153,N_28721,N_28351);
nor U30154 (N_30154,N_28356,N_29033);
xnor U30155 (N_30155,N_29001,N_28248);
nor U30156 (N_30156,N_29079,N_28592);
or U30157 (N_30157,N_29126,N_29268);
nand U30158 (N_30158,N_28440,N_29378);
xor U30159 (N_30159,N_29373,N_29441);
nor U30160 (N_30160,N_29682,N_29354);
and U30161 (N_30161,N_29715,N_28423);
nor U30162 (N_30162,N_28165,N_28541);
nor U30163 (N_30163,N_28400,N_29158);
nor U30164 (N_30164,N_28534,N_29090);
xor U30165 (N_30165,N_29672,N_28659);
nor U30166 (N_30166,N_29567,N_29533);
nand U30167 (N_30167,N_29806,N_28139);
and U30168 (N_30168,N_28852,N_29863);
and U30169 (N_30169,N_28208,N_29476);
nor U30170 (N_30170,N_28688,N_28672);
nand U30171 (N_30171,N_29136,N_28374);
nor U30172 (N_30172,N_29021,N_28401);
xor U30173 (N_30173,N_28511,N_29719);
xnor U30174 (N_30174,N_29666,N_28117);
or U30175 (N_30175,N_29006,N_29072);
nor U30176 (N_30176,N_28804,N_29274);
or U30177 (N_30177,N_28318,N_28849);
and U30178 (N_30178,N_29159,N_28481);
nor U30179 (N_30179,N_29405,N_28813);
nand U30180 (N_30180,N_29924,N_29617);
and U30181 (N_30181,N_28392,N_29685);
xnor U30182 (N_30182,N_29146,N_29651);
nand U30183 (N_30183,N_28017,N_29708);
and U30184 (N_30184,N_29950,N_29087);
nor U30185 (N_30185,N_29015,N_28262);
nor U30186 (N_30186,N_28388,N_29492);
nor U30187 (N_30187,N_29745,N_28019);
xor U30188 (N_30188,N_29760,N_29776);
xor U30189 (N_30189,N_28973,N_29647);
and U30190 (N_30190,N_29009,N_28691);
xor U30191 (N_30191,N_29994,N_29482);
and U30192 (N_30192,N_28382,N_29505);
nor U30193 (N_30193,N_28280,N_28096);
or U30194 (N_30194,N_29671,N_29993);
nor U30195 (N_30195,N_28911,N_29325);
nand U30196 (N_30196,N_29726,N_29221);
nand U30197 (N_30197,N_29304,N_29996);
nor U30198 (N_30198,N_29582,N_29367);
xnor U30199 (N_30199,N_29209,N_29218);
nor U30200 (N_30200,N_29638,N_29653);
nor U30201 (N_30201,N_29289,N_28137);
and U30202 (N_30202,N_28065,N_29322);
xnor U30203 (N_30203,N_29181,N_28106);
and U30204 (N_30204,N_28931,N_29428);
or U30205 (N_30205,N_29453,N_28376);
xnor U30206 (N_30206,N_29361,N_29192);
and U30207 (N_30207,N_29674,N_29023);
xnor U30208 (N_30208,N_29278,N_28995);
nand U30209 (N_30209,N_28803,N_28986);
nand U30210 (N_30210,N_28719,N_29445);
nor U30211 (N_30211,N_28580,N_28558);
and U30212 (N_30212,N_29954,N_29503);
nand U30213 (N_30213,N_28878,N_28854);
nand U30214 (N_30214,N_28406,N_29030);
xnor U30215 (N_30215,N_29628,N_28110);
and U30216 (N_30216,N_28230,N_28074);
xnor U30217 (N_30217,N_28194,N_29258);
or U30218 (N_30218,N_28887,N_29794);
and U30219 (N_30219,N_28905,N_28195);
and U30220 (N_30220,N_28978,N_28090);
nand U30221 (N_30221,N_28433,N_29396);
nand U30222 (N_30222,N_29869,N_29722);
xor U30223 (N_30223,N_29376,N_29407);
nand U30224 (N_30224,N_29198,N_28340);
or U30225 (N_30225,N_28075,N_29693);
and U30226 (N_30226,N_29856,N_28638);
nand U30227 (N_30227,N_28114,N_28121);
and U30228 (N_30228,N_28067,N_28596);
nand U30229 (N_30229,N_29694,N_28022);
and U30230 (N_30230,N_28900,N_28082);
nand U30231 (N_30231,N_29712,N_29515);
nor U30232 (N_30232,N_29622,N_29840);
or U30233 (N_30233,N_28304,N_28668);
xor U30234 (N_30234,N_28588,N_29585);
and U30235 (N_30235,N_29069,N_28445);
and U30236 (N_30236,N_29070,N_29077);
nor U30237 (N_30237,N_28785,N_28564);
xnor U30238 (N_30238,N_29369,N_28369);
and U30239 (N_30239,N_28814,N_28902);
nand U30240 (N_30240,N_29743,N_29948);
and U30241 (N_30241,N_28552,N_28526);
and U30242 (N_30242,N_28373,N_28058);
nand U30243 (N_30243,N_29705,N_29696);
and U30244 (N_30244,N_28359,N_29498);
nor U30245 (N_30245,N_29681,N_28004);
nor U30246 (N_30246,N_28595,N_28696);
nor U30247 (N_30247,N_29053,N_29620);
or U30248 (N_30248,N_28241,N_28024);
or U30249 (N_30249,N_29401,N_29642);
and U30250 (N_30250,N_29237,N_28333);
or U30251 (N_30251,N_28996,N_29963);
and U30252 (N_30252,N_29271,N_28654);
xor U30253 (N_30253,N_29475,N_29408);
nand U30254 (N_30254,N_29992,N_29463);
nand U30255 (N_30255,N_29901,N_29556);
or U30256 (N_30256,N_29051,N_29872);
and U30257 (N_30257,N_29379,N_29468);
xor U30258 (N_30258,N_29836,N_28315);
xor U30259 (N_30259,N_29947,N_28487);
nor U30260 (N_30260,N_28790,N_29801);
xnor U30261 (N_30261,N_28958,N_28930);
nor U30262 (N_30262,N_29586,N_28378);
xnor U30263 (N_30263,N_29118,N_29854);
nand U30264 (N_30264,N_28773,N_29484);
nor U30265 (N_30265,N_29524,N_28872);
or U30266 (N_30266,N_28418,N_28634);
or U30267 (N_30267,N_29332,N_28689);
and U30268 (N_30268,N_28499,N_28201);
nor U30269 (N_30269,N_28370,N_28292);
or U30270 (N_30270,N_29673,N_28207);
xor U30271 (N_30271,N_29097,N_29908);
and U30272 (N_30272,N_29769,N_28228);
nor U30273 (N_30273,N_28154,N_29746);
or U30274 (N_30274,N_28928,N_28834);
xor U30275 (N_30275,N_29852,N_28741);
or U30276 (N_30276,N_29493,N_28480);
nor U30277 (N_30277,N_29525,N_29573);
xnor U30278 (N_30278,N_28297,N_29838);
nor U30279 (N_30279,N_28828,N_28559);
xnor U30280 (N_30280,N_29612,N_29093);
xor U30281 (N_30281,N_29199,N_29985);
xnor U30282 (N_30282,N_29623,N_28299);
nand U30283 (N_30283,N_28906,N_29979);
or U30284 (N_30284,N_29085,N_28747);
or U30285 (N_30285,N_29520,N_29189);
or U30286 (N_30286,N_28947,N_28807);
and U30287 (N_30287,N_28677,N_29971);
and U30288 (N_30288,N_28456,N_29451);
and U30289 (N_30289,N_29526,N_29686);
nor U30290 (N_30290,N_28416,N_29815);
nand U30291 (N_30291,N_28992,N_29457);
nor U30292 (N_30292,N_29455,N_28452);
or U30293 (N_30293,N_28786,N_29190);
and U30294 (N_30294,N_28628,N_28831);
or U30295 (N_30295,N_29818,N_29824);
and U30296 (N_30296,N_28671,N_29663);
nor U30297 (N_30297,N_29839,N_29659);
or U30298 (N_30298,N_29397,N_29995);
xor U30299 (N_30299,N_28232,N_28764);
and U30300 (N_30300,N_29942,N_29926);
and U30301 (N_30301,N_28598,N_29111);
xor U30302 (N_30302,N_29522,N_29655);
nand U30303 (N_30303,N_29575,N_29748);
or U30304 (N_30304,N_29870,N_29448);
nand U30305 (N_30305,N_28352,N_28153);
nand U30306 (N_30306,N_28933,N_28779);
or U30307 (N_30307,N_29337,N_28611);
nand U30308 (N_30308,N_29699,N_28964);
nand U30309 (N_30309,N_29283,N_28367);
nand U30310 (N_30310,N_29173,N_28708);
nor U30311 (N_30311,N_28197,N_29601);
nand U30312 (N_30312,N_28021,N_28018);
and U30313 (N_30313,N_28776,N_29454);
xor U30314 (N_30314,N_28826,N_29730);
or U30315 (N_30315,N_29029,N_28188);
and U30316 (N_30316,N_29546,N_28284);
xnor U30317 (N_30317,N_29596,N_28486);
nand U30318 (N_30318,N_28431,N_29194);
nor U30319 (N_30319,N_28221,N_28334);
and U30320 (N_30320,N_29527,N_29259);
and U30321 (N_30321,N_29600,N_29449);
xor U30322 (N_30322,N_29735,N_28839);
and U30323 (N_30323,N_28502,N_29032);
nand U30324 (N_30324,N_28586,N_29918);
xnor U30325 (N_30325,N_29243,N_28972);
nor U30326 (N_30326,N_28185,N_29052);
nor U30327 (N_30327,N_28675,N_28910);
xor U30328 (N_30328,N_28966,N_29565);
or U30329 (N_30329,N_28450,N_29821);
xor U30330 (N_30330,N_28842,N_28390);
or U30331 (N_30331,N_29327,N_29116);
xnor U30332 (N_30332,N_28468,N_29831);
or U30333 (N_30333,N_28685,N_29956);
nor U30334 (N_30334,N_28429,N_28129);
or U30335 (N_30335,N_29654,N_28325);
xor U30336 (N_30336,N_29336,N_28398);
or U30337 (N_30337,N_28723,N_29370);
nand U30338 (N_30338,N_28116,N_29678);
xor U30339 (N_30339,N_28515,N_28821);
nor U30340 (N_30340,N_29521,N_29164);
or U30341 (N_30341,N_29429,N_28577);
nor U30342 (N_30342,N_28864,N_28886);
xor U30343 (N_30343,N_28571,N_29108);
nor U30344 (N_30344,N_29059,N_28805);
xnor U30345 (N_30345,N_28200,N_29975);
nor U30346 (N_30346,N_29417,N_28954);
or U30347 (N_30347,N_29414,N_28909);
nor U30348 (N_30348,N_28293,N_29551);
or U30349 (N_30349,N_28476,N_29151);
or U30350 (N_30350,N_28312,N_28353);
and U30351 (N_30351,N_29559,N_28774);
and U30352 (N_30352,N_28282,N_28439);
or U30353 (N_30353,N_29098,N_29610);
xor U30354 (N_30354,N_28229,N_29549);
and U30355 (N_30355,N_29853,N_29754);
or U30356 (N_30356,N_29881,N_29249);
and U30357 (N_30357,N_29917,N_28069);
or U30358 (N_30358,N_28441,N_28968);
nor U30359 (N_30359,N_29868,N_29676);
nor U30360 (N_30360,N_28368,N_29380);
nand U30361 (N_30361,N_29581,N_28550);
nor U30362 (N_30362,N_28011,N_28257);
or U30363 (N_30363,N_28060,N_28107);
nor U30364 (N_30364,N_28179,N_28138);
and U30365 (N_30365,N_29631,N_28528);
or U30366 (N_30366,N_28002,N_28664);
and U30367 (N_30367,N_29145,N_28043);
xor U30368 (N_30368,N_28122,N_28600);
or U30369 (N_30369,N_29203,N_28625);
xnor U30370 (N_30370,N_28527,N_28833);
and U30371 (N_30371,N_29331,N_28196);
nor U30372 (N_30372,N_29844,N_29107);
or U30373 (N_30373,N_29394,N_28478);
nor U30374 (N_30374,N_28520,N_29269);
or U30375 (N_30375,N_29326,N_28205);
and U30376 (N_30376,N_29731,N_29998);
nand U30377 (N_30377,N_29356,N_28485);
nor U30378 (N_30378,N_28765,N_28296);
nor U30379 (N_30379,N_28357,N_29296);
nand U30380 (N_30380,N_28898,N_29131);
xnor U30381 (N_30381,N_28224,N_29162);
and U30382 (N_30382,N_28213,N_29946);
nor U30383 (N_30383,N_28451,N_29166);
nor U30384 (N_30384,N_28162,N_28361);
and U30385 (N_30385,N_28863,N_28919);
nand U30386 (N_30386,N_28766,N_29091);
and U30387 (N_30387,N_28488,N_29792);
nor U30388 (N_30388,N_29517,N_29716);
and U30389 (N_30389,N_28925,N_28627);
nor U30390 (N_30390,N_28380,N_28874);
xor U30391 (N_30391,N_28337,N_28977);
nand U30392 (N_30392,N_28787,N_28347);
xnor U30393 (N_30393,N_28054,N_28982);
and U30394 (N_30394,N_28781,N_29564);
xor U30395 (N_30395,N_29076,N_29168);
and U30396 (N_30396,N_28404,N_29000);
and U30397 (N_30397,N_29911,N_29952);
or U30398 (N_30398,N_29080,N_29236);
or U30399 (N_30399,N_28120,N_28561);
nand U30400 (N_30400,N_29615,N_29372);
or U30401 (N_30401,N_28088,N_29741);
or U30402 (N_30402,N_28161,N_28802);
and U30403 (N_30403,N_28035,N_29578);
nor U30404 (N_30404,N_28771,N_28870);
nor U30405 (N_30405,N_28673,N_28553);
nand U30406 (N_30406,N_28645,N_29759);
nand U30407 (N_30407,N_29435,N_29867);
or U30408 (N_30408,N_29135,N_28503);
nor U30409 (N_30409,N_28276,N_29577);
nor U30410 (N_30410,N_28882,N_29811);
nand U30411 (N_30411,N_29544,N_28323);
and U30412 (N_30412,N_28198,N_29553);
xor U30413 (N_30413,N_29110,N_28555);
or U30414 (N_30414,N_29240,N_29293);
nand U30415 (N_30415,N_29122,N_29762);
nand U30416 (N_30416,N_29763,N_28994);
nand U30417 (N_30417,N_28866,N_29078);
nand U30418 (N_30418,N_29260,N_28070);
xor U30419 (N_30419,N_29252,N_28403);
and U30420 (N_30420,N_29275,N_28264);
xnor U30421 (N_30421,N_28084,N_29508);
or U30422 (N_30422,N_28823,N_28934);
xor U30423 (N_30423,N_28039,N_29316);
or U30424 (N_30424,N_29375,N_29636);
nand U30425 (N_30425,N_29179,N_29421);
nand U30426 (N_30426,N_29805,N_28525);
xor U30427 (N_30427,N_28331,N_28078);
and U30428 (N_30428,N_28381,N_29205);
xnor U30429 (N_30429,N_29558,N_28832);
and U30430 (N_30430,N_28704,N_28752);
nand U30431 (N_30431,N_29547,N_28365);
or U30432 (N_30432,N_29250,N_28514);
and U30433 (N_30433,N_29882,N_29470);
xnor U30434 (N_30434,N_28999,N_29860);
nor U30435 (N_30435,N_28332,N_28560);
and U30436 (N_30436,N_29864,N_28794);
or U30437 (N_30437,N_28647,N_28434);
and U30438 (N_30438,N_28033,N_29057);
nand U30439 (N_30439,N_28328,N_28097);
nand U30440 (N_30440,N_28554,N_28686);
nand U30441 (N_30441,N_29365,N_29310);
xnor U30442 (N_30442,N_29506,N_29875);
nor U30443 (N_30443,N_28661,N_29244);
or U30444 (N_30444,N_28865,N_29721);
nand U30445 (N_30445,N_29569,N_29466);
nor U30446 (N_30446,N_29808,N_28094);
or U30447 (N_30447,N_28987,N_28722);
or U30448 (N_30448,N_29290,N_29630);
and U30449 (N_30449,N_28455,N_29966);
or U30450 (N_30450,N_29308,N_29127);
xnor U30451 (N_30451,N_28782,N_29813);
nor U30452 (N_30452,N_29014,N_28762);
xnor U30453 (N_30453,N_29294,N_28707);
xnor U30454 (N_30454,N_28665,N_28609);
or U30455 (N_30455,N_28916,N_29017);
nor U30456 (N_30456,N_28643,N_28490);
and U30457 (N_30457,N_29234,N_29467);
and U30458 (N_30458,N_29626,N_28549);
nand U30459 (N_30459,N_28389,N_29385);
xnor U30460 (N_30460,N_28593,N_29055);
and U30461 (N_30461,N_29861,N_28969);
and U30462 (N_30462,N_28989,N_29644);
nor U30463 (N_30463,N_28220,N_28792);
and U30464 (N_30464,N_28760,N_29570);
or U30465 (N_30465,N_28192,N_28030);
xnor U30466 (N_30466,N_29518,N_28698);
or U30467 (N_30467,N_29736,N_28254);
xor U30468 (N_30468,N_28288,N_29896);
nand U30469 (N_30469,N_29073,N_28840);
and U30470 (N_30470,N_29099,N_28473);
nand U30471 (N_30471,N_29962,N_29180);
and U30472 (N_30472,N_28342,N_29292);
nor U30473 (N_30473,N_29266,N_29094);
nor U30474 (N_30474,N_28924,N_29828);
or U30475 (N_30475,N_29062,N_28271);
nor U30476 (N_30476,N_28926,N_28251);
and U30477 (N_30477,N_28875,N_29873);
or U30478 (N_30478,N_29499,N_29286);
nor U30479 (N_30479,N_29176,N_29789);
nand U30480 (N_30480,N_29253,N_29530);
and U30481 (N_30481,N_29027,N_29024);
xor U30482 (N_30482,N_29299,N_28569);
nor U30483 (N_30483,N_28438,N_28177);
and U30484 (N_30484,N_29478,N_28937);
and U30485 (N_30485,N_29669,N_29340);
and U30486 (N_30486,N_29846,N_29063);
or U30487 (N_30487,N_29132,N_29819);
or U30488 (N_30488,N_29188,N_28267);
or U30489 (N_30489,N_29787,N_29751);
or U30490 (N_30490,N_29068,N_28395);
xor U30491 (N_30491,N_28847,N_28830);
xor U30492 (N_30492,N_29714,N_28738);
nand U30493 (N_30493,N_29458,N_29862);
or U30494 (N_30494,N_29501,N_29930);
or U30495 (N_30495,N_29491,N_29263);
nand U30496 (N_30496,N_28134,N_29554);
nor U30497 (N_30497,N_29016,N_28093);
and U30498 (N_30498,N_29495,N_28537);
or U30499 (N_30499,N_28574,N_28505);
nor U30500 (N_30500,N_29961,N_28504);
xnor U30501 (N_30501,N_29598,N_29104);
or U30502 (N_30502,N_29165,N_29691);
and U30503 (N_30503,N_28684,N_28459);
nand U30504 (N_30504,N_29740,N_29061);
xnor U30505 (N_30505,N_29703,N_28063);
xor U30506 (N_30506,N_28085,N_29810);
nor U30507 (N_30507,N_29058,N_28649);
or U30508 (N_30508,N_29210,N_28279);
nand U30509 (N_30509,N_28111,N_29987);
nand U30510 (N_30510,N_29245,N_28815);
nor U30511 (N_30511,N_28186,N_28565);
nor U30512 (N_30512,N_29477,N_29886);
nor U30513 (N_30513,N_28100,N_29255);
or U30514 (N_30514,N_28768,N_29641);
or U30515 (N_30515,N_29986,N_29925);
or U30516 (N_30516,N_28041,N_29888);
and U30517 (N_30517,N_28510,N_29768);
nor U30518 (N_30518,N_29932,N_29607);
nor U30519 (N_30519,N_28917,N_28694);
nand U30520 (N_30520,N_28432,N_28015);
and U30521 (N_30521,N_29758,N_28447);
and U30522 (N_30522,N_29412,N_29172);
xnor U30523 (N_30523,N_28210,N_28016);
nand U30524 (N_30524,N_29711,N_29919);
or U30525 (N_30525,N_28599,N_28020);
nor U30526 (N_30526,N_29148,N_29756);
or U30527 (N_30527,N_28448,N_28710);
xnor U30528 (N_30528,N_29587,N_28980);
nor U30529 (N_30529,N_28620,N_28614);
xor U30530 (N_30530,N_28291,N_28187);
nor U30531 (N_30531,N_29036,N_29803);
nor U30532 (N_30532,N_29724,N_28621);
and U30533 (N_30533,N_28575,N_29542);
xor U30534 (N_30534,N_28104,N_29764);
and U30535 (N_30535,N_28601,N_29519);
nand U30536 (N_30536,N_29723,N_29841);
xor U30537 (N_30537,N_28099,N_28929);
nand U30538 (N_30538,N_28311,N_28780);
or U30539 (N_30539,N_29143,N_29652);
or U30540 (N_30540,N_28799,N_29718);
xnor U30541 (N_30541,N_29898,N_28386);
nor U30542 (N_30542,N_28343,N_29637);
nor U30543 (N_30543,N_28492,N_29725);
or U30544 (N_30544,N_29497,N_28412);
nor U30545 (N_30545,N_29679,N_29778);
xor U30546 (N_30546,N_29605,N_29633);
nand U30547 (N_30547,N_28761,N_28693);
or U30548 (N_30548,N_28409,N_29970);
xnor U30549 (N_30549,N_29067,N_29037);
xor U30550 (N_30550,N_29472,N_29753);
and U30551 (N_30551,N_28430,N_29060);
nand U30552 (N_30552,N_28027,N_29757);
or U30553 (N_30553,N_28538,N_29400);
xnor U30554 (N_30554,N_29439,N_29334);
and U30555 (N_30555,N_28474,N_29238);
or U30556 (N_30556,N_28091,N_28626);
or U30557 (N_30557,N_28467,N_28385);
nor U30558 (N_30558,N_28132,N_28055);
nor U30559 (N_30559,N_28530,N_29418);
nand U30560 (N_30560,N_29964,N_29355);
nand U30561 (N_30561,N_29913,N_28425);
or U30562 (N_30562,N_29749,N_29662);
and U30563 (N_30563,N_28956,N_29291);
nor U30564 (N_30564,N_29229,N_28610);
xor U30565 (N_30565,N_28651,N_29583);
nand U30566 (N_30566,N_28590,N_28618);
or U30567 (N_30567,N_29510,N_28298);
xnor U30568 (N_30568,N_28169,N_29201);
and U30569 (N_30569,N_29775,N_29774);
and U30570 (N_30570,N_29690,N_29071);
nor U30571 (N_30571,N_29469,N_29902);
nand U30572 (N_30572,N_29765,N_28509);
or U30573 (N_30573,N_28335,N_28705);
or U30574 (N_30574,N_29972,N_28507);
or U30575 (N_30575,N_28443,N_29459);
and U30576 (N_30576,N_28464,N_29528);
or U30577 (N_30577,N_28703,N_28726);
or U30578 (N_30578,N_29362,N_29728);
nor U30579 (N_30579,N_29780,N_28124);
xor U30580 (N_30580,N_29347,N_29667);
xor U30581 (N_30581,N_29984,N_28320);
nand U30582 (N_30582,N_29702,N_28713);
nand U30583 (N_30583,N_29732,N_29695);
and U30584 (N_30584,N_29675,N_28529);
nand U30585 (N_30585,N_28797,N_29788);
nand U30586 (N_30586,N_28518,N_29328);
xor U30587 (N_30587,N_28339,N_29704);
and U30588 (N_30588,N_28636,N_28072);
nand U30589 (N_30589,N_29973,N_28682);
and U30590 (N_30590,N_28635,N_28736);
and U30591 (N_30591,N_29580,N_29783);
xnor U30592 (N_30592,N_29706,N_28984);
and U30593 (N_30593,N_29670,N_29339);
nor U30594 (N_30594,N_29446,N_28193);
nand U30595 (N_30595,N_28943,N_29196);
nand U30596 (N_30596,N_28301,N_28172);
or U30597 (N_30597,N_28245,N_29011);
or U30598 (N_30598,N_28744,N_28243);
and U30599 (N_30599,N_29632,N_29197);
nand U30600 (N_30600,N_28081,N_29398);
or U30601 (N_30601,N_29635,N_29481);
and U30602 (N_30602,N_29330,N_29371);
nand U30603 (N_30603,N_28777,N_29843);
xor U30604 (N_30604,N_28731,N_29767);
or U30605 (N_30605,N_28951,N_28290);
and U30606 (N_30606,N_29755,N_28131);
or U30607 (N_30607,N_29563,N_29656);
and U30608 (N_30608,N_29314,N_28250);
or U30609 (N_30609,N_29507,N_28637);
nand U30610 (N_30610,N_29634,N_28355);
and U30611 (N_30611,N_28252,N_28247);
nor U30612 (N_30612,N_29117,N_29256);
and U30613 (N_30613,N_29319,N_28417);
and U30614 (N_30614,N_29474,N_29734);
and U30615 (N_30615,N_29795,N_28798);
or U30616 (N_30616,N_29604,N_28881);
or U30617 (N_30617,N_29949,N_29288);
and U30618 (N_30618,N_29939,N_29812);
and U30619 (N_30619,N_28407,N_29988);
nand U30620 (N_30620,N_28819,N_28300);
nand U30621 (N_30621,N_28850,N_28491);
xor U30622 (N_30622,N_29957,N_28105);
nand U30623 (N_30623,N_29907,N_29981);
and U30624 (N_30624,N_29241,N_29899);
nand U30625 (N_30625,N_28109,N_29054);
nor U30626 (N_30626,N_29103,N_28344);
nor U30627 (N_30627,N_28648,N_29941);
or U30628 (N_30628,N_28988,N_28219);
or U30629 (N_30629,N_29677,N_29648);
and U30630 (N_30630,N_28608,N_28305);
and U30631 (N_30631,N_28244,N_29303);
or U30632 (N_30632,N_29698,N_29089);
or U30633 (N_30633,N_29568,N_28045);
nor U30634 (N_30634,N_28745,N_29003);
and U30635 (N_30635,N_28494,N_28962);
and U30636 (N_30636,N_29022,N_28206);
xnor U30637 (N_30637,N_28714,N_29083);
nand U30638 (N_30638,N_29540,N_28345);
or U30639 (N_30639,N_28674,N_29684);
xnor U30640 (N_30640,N_28287,N_29590);
or U30641 (N_30641,N_28979,N_28475);
and U30642 (N_30642,N_29387,N_29597);
and U30643 (N_30643,N_29974,N_29827);
nand U30644 (N_30644,N_29219,N_29231);
nand U30645 (N_30645,N_28871,N_29649);
xnor U30646 (N_30646,N_28482,N_29223);
xor U30647 (N_30647,N_29609,N_28961);
nor U30648 (N_30648,N_29395,N_28143);
or U30649 (N_30649,N_28885,N_29427);
nor U30650 (N_30650,N_28963,N_28946);
xor U30651 (N_30651,N_29823,N_29490);
and U30652 (N_30652,N_28606,N_29614);
and U30653 (N_30653,N_28836,N_28178);
xor U30654 (N_30654,N_28733,N_29025);
nor U30655 (N_30655,N_29010,N_28522);
xor U30656 (N_30656,N_28348,N_28470);
or U30657 (N_30657,N_29115,N_28263);
nor U30658 (N_30658,N_28701,N_29434);
xor U30659 (N_30659,N_29858,N_28141);
and U30660 (N_30660,N_28655,N_28413);
and U30661 (N_30661,N_29321,N_29940);
or U30662 (N_30662,N_28557,N_28051);
nor U30663 (N_30663,N_29980,N_28140);
nor U30664 (N_30664,N_29285,N_29665);
xor U30665 (N_30665,N_28150,N_28889);
nor U30666 (N_30666,N_28007,N_29295);
nor U30667 (N_30667,N_28317,N_29892);
xnor U30668 (N_30668,N_29217,N_28950);
xnor U30669 (N_30669,N_28489,N_28936);
nand U30670 (N_30670,N_29204,N_29424);
and U30671 (N_30671,N_29660,N_28506);
nor U30672 (N_30672,N_29514,N_28796);
or U30673 (N_30673,N_29208,N_29483);
xor U30674 (N_30674,N_29770,N_29012);
nand U30675 (N_30675,N_28658,N_28720);
or U30676 (N_30676,N_29591,N_29389);
and U30677 (N_30677,N_28895,N_29618);
nand U30678 (N_30678,N_28543,N_28013);
and U30679 (N_30679,N_28508,N_28639);
and U30680 (N_30680,N_29276,N_28816);
nor U30681 (N_30681,N_29594,N_28808);
nor U30682 (N_30682,N_28789,N_29184);
and U30683 (N_30683,N_28128,N_28860);
and U30684 (N_30684,N_28584,N_28077);
xnor U30685 (N_30685,N_29119,N_29112);
xnor U30686 (N_30686,N_29999,N_28818);
and U30687 (N_30687,N_28329,N_28255);
xor U30688 (N_30688,N_28184,N_29415);
xor U30689 (N_30689,N_29814,N_29082);
and U30690 (N_30690,N_29300,N_29462);
and U30691 (N_30691,N_29968,N_29683);
and U30692 (N_30692,N_28540,N_29713);
nand U30693 (N_30693,N_28711,N_28570);
nand U30694 (N_30694,N_29139,N_29138);
nand U30695 (N_30695,N_29157,N_29411);
nand U30696 (N_30696,N_28955,N_28371);
or U30697 (N_30697,N_28544,N_28500);
nor U30698 (N_30698,N_28155,N_28753);
nor U30699 (N_30699,N_28932,N_29900);
xor U30700 (N_30700,N_28056,N_28846);
nor U30701 (N_30701,N_28851,N_29137);
nand U30702 (N_30702,N_28227,N_28012);
xor U30703 (N_30703,N_28709,N_29381);
xnor U30704 (N_30704,N_29261,N_29182);
nand U30705 (N_30705,N_28743,N_29456);
and U30706 (N_30706,N_29539,N_29109);
nor U30707 (N_30707,N_29402,N_28759);
xor U30708 (N_30708,N_28727,N_29923);
or U30709 (N_30709,N_29976,N_29560);
nand U30710 (N_30710,N_28421,N_28217);
and U30711 (N_30711,N_28484,N_29643);
and U30712 (N_30712,N_28354,N_29160);
or U30713 (N_30713,N_28466,N_29357);
nand U30714 (N_30714,N_29625,N_28268);
or U30715 (N_30715,N_28660,N_28189);
xor U30716 (N_30716,N_28294,N_29552);
nor U30717 (N_30717,N_28547,N_29178);
xnor U30718 (N_30718,N_28079,N_28901);
nand U30719 (N_30719,N_28841,N_29388);
xor U30720 (N_30720,N_28563,N_29479);
nand U30721 (N_30721,N_29857,N_29943);
or U30722 (N_30722,N_29916,N_29267);
nor U30723 (N_30723,N_29461,N_28175);
nand U30724 (N_30724,N_29692,N_29113);
and U30725 (N_30725,N_29187,N_28026);
or U30726 (N_30726,N_29785,N_29878);
nand U30727 (N_30727,N_28567,N_28795);
or U30728 (N_30728,N_28278,N_28820);
and U30729 (N_30729,N_28844,N_28008);
nand U30730 (N_30730,N_28038,N_28112);
or U30731 (N_30731,N_28236,N_28307);
and U30732 (N_30732,N_29592,N_29264);
nor U30733 (N_30733,N_29106,N_28483);
xnor U30734 (N_30734,N_29047,N_29817);
nor U30735 (N_30735,N_28556,N_29153);
nor U30736 (N_30736,N_28174,N_29254);
nor U30737 (N_30737,N_29557,N_28442);
nand U30738 (N_30738,N_28546,N_28059);
xnor U30739 (N_30739,N_29018,N_28095);
nor U30740 (N_30740,N_28729,N_29645);
nand U30741 (N_30741,N_29335,N_29464);
nand U30742 (N_30742,N_28861,N_29020);
xnor U30743 (N_30743,N_28829,N_29835);
nand U30744 (N_30744,N_28061,N_28049);
or U30745 (N_30745,N_29125,N_28739);
or U30746 (N_30746,N_28216,N_28585);
xnor U30747 (N_30747,N_28199,N_28806);
or U30748 (N_30748,N_28176,N_28742);
nand U30749 (N_30749,N_28029,N_29701);
and U30750 (N_30750,N_28853,N_29537);
and U30751 (N_30751,N_28454,N_29877);
xor U30752 (N_30752,N_28678,N_29739);
nor U30753 (N_30753,N_29982,N_29351);
xnor U30754 (N_30754,N_28856,N_29793);
nand U30755 (N_30755,N_29571,N_29305);
nand U30756 (N_30756,N_29431,N_28548);
xor U30757 (N_30757,N_29284,N_29611);
nand U30758 (N_30758,N_28572,N_29257);
or U30759 (N_30759,N_28001,N_28062);
nand U30760 (N_30760,N_29485,N_28715);
xor U30761 (N_30761,N_28125,N_28867);
and U30762 (N_30762,N_28212,N_29599);
nor U30763 (N_30763,N_29206,N_29859);
xor U30764 (N_30764,N_28435,N_28009);
xnor U30765 (N_30765,N_29409,N_28053);
or U30766 (N_30766,N_29242,N_29442);
xnor U30767 (N_30767,N_28397,N_28927);
or U30768 (N_30768,N_28687,N_28604);
nand U30769 (N_30769,N_29101,N_29752);
and U30770 (N_30770,N_28892,N_28868);
or U30771 (N_30771,N_28670,N_29738);
xor U30772 (N_30772,N_29922,N_28270);
nand U30773 (N_30773,N_28680,N_28578);
nand U30774 (N_30774,N_29566,N_29232);
xor U30775 (N_30775,N_28366,N_28260);
nor U30776 (N_30776,N_29978,N_28848);
and U30777 (N_30777,N_28629,N_28379);
or U30778 (N_30778,N_29550,N_29891);
nand U30779 (N_30779,N_28173,N_29056);
and U30780 (N_30780,N_28734,N_28521);
or U30781 (N_30781,N_28633,N_29120);
xnor U30782 (N_30782,N_28259,N_28531);
and U30783 (N_30783,N_28493,N_28607);
or U30784 (N_30784,N_28462,N_28619);
and U30785 (N_30785,N_29046,N_28086);
nand U30786 (N_30786,N_28641,N_29186);
and U30787 (N_30787,N_28269,N_28908);
xor U30788 (N_30788,N_29248,N_29175);
nor U30789 (N_30789,N_29004,N_28170);
nand U30790 (N_30790,N_28903,N_29344);
or U30791 (N_30791,N_28763,N_29318);
xnor U30792 (N_30792,N_29391,N_29621);
or U30793 (N_30793,N_28812,N_29969);
and U30794 (N_30794,N_28285,N_28363);
nor U30795 (N_30795,N_28827,N_28163);
nand U30796 (N_30796,N_29816,N_28246);
xor U30797 (N_30797,N_29629,N_29161);
and U30798 (N_30798,N_29171,N_28160);
nor U30799 (N_30799,N_28014,N_29211);
and U30800 (N_30800,N_28239,N_28616);
nand U30801 (N_30801,N_28295,N_28692);
and U30802 (N_30802,N_29613,N_29045);
nand U30803 (N_30803,N_29273,N_28516);
and U30804 (N_30804,N_29317,N_29353);
nor U30805 (N_30805,N_28591,N_28191);
and U30806 (N_30806,N_28904,N_29040);
nand U30807 (N_30807,N_29541,N_28869);
or U30808 (N_30808,N_29761,N_28573);
and U30809 (N_30809,N_28811,N_29849);
and U30810 (N_30810,N_29239,N_28624);
xnor U30811 (N_30811,N_29865,N_28959);
and U30812 (N_30812,N_29727,N_28422);
and U30813 (N_30813,N_29019,N_28411);
or U30814 (N_30814,N_28725,N_29531);
nand U30815 (N_30815,N_28362,N_29965);
and U30816 (N_30816,N_29212,N_28669);
nand U30817 (N_30817,N_28463,N_28346);
xor U30818 (N_30818,N_28883,N_29177);
nor U30819 (N_30819,N_29829,N_29884);
and U30820 (N_30820,N_29215,N_29130);
nor U30821 (N_30821,N_29737,N_29193);
nand U30822 (N_30822,N_29936,N_29404);
nand U30823 (N_30823,N_29697,N_28203);
or U30824 (N_30824,N_29847,N_29488);
or U30825 (N_30825,N_28277,N_29191);
nand U30826 (N_30826,N_28653,N_29931);
nand U30827 (N_30827,N_28920,N_29156);
xor U30828 (N_30828,N_29384,N_28622);
and U30829 (N_30829,N_29043,N_28748);
nand U30830 (N_30830,N_28133,N_29246);
and U30831 (N_30831,N_28272,N_28981);
or U30832 (N_30832,N_29128,N_28415);
and U30833 (N_30833,N_29393,N_28922);
nor U30834 (N_30834,N_28326,N_28405);
nor U30835 (N_30835,N_28594,N_29324);
nand U30836 (N_30836,N_28791,N_29809);
nand U30837 (N_30837,N_29516,N_28071);
nand U30838 (N_30838,N_29876,N_29227);
or U30839 (N_30839,N_29086,N_28623);
or U30840 (N_30840,N_28314,N_28037);
nor U30841 (N_30841,N_29657,N_28286);
nand U30842 (N_30842,N_29927,N_28028);
and U30843 (N_30843,N_29800,N_28890);
nor U30844 (N_30844,N_28681,N_29416);
xor U30845 (N_30845,N_29364,N_29880);
and U30846 (N_30846,N_29438,N_28617);
nor U30847 (N_30847,N_28261,N_29382);
nand U30848 (N_30848,N_28375,N_28144);
and U30849 (N_30849,N_29826,N_28770);
and U30850 (N_30850,N_29413,N_29909);
or U30851 (N_30851,N_29717,N_29235);
and U30852 (N_30852,N_28145,N_29733);
or U30853 (N_30853,N_28057,N_29750);
or U30854 (N_30854,N_28952,N_29399);
or U30855 (N_30855,N_28040,N_28912);
nor U30856 (N_30856,N_29879,N_29374);
nor U30857 (N_30857,N_29311,N_29807);
xnor U30858 (N_30858,N_28751,N_29346);
xnor U30859 (N_30859,N_28283,N_28146);
and U30860 (N_30860,N_29224,N_28915);
nand U30861 (N_30861,N_28640,N_28308);
nand U30862 (N_30862,N_28135,N_29333);
xnor U30863 (N_30863,N_28204,N_29443);
or U30864 (N_30864,N_29850,N_29820);
xor U30865 (N_30865,N_28316,N_28944);
or U30866 (N_30866,N_28387,N_29603);
nor U30867 (N_30867,N_29894,N_29390);
or U30868 (N_30868,N_28532,N_28266);
and U30869 (N_30869,N_28695,N_28136);
nand U30870 (N_30870,N_28993,N_29005);
xnor U30871 (N_30871,N_29088,N_28755);
xnor U30872 (N_30872,N_29302,N_29147);
and U30873 (N_30873,N_29377,N_28225);
or U30874 (N_30874,N_28942,N_28036);
nand U30875 (N_30875,N_28907,N_29773);
and U30876 (N_30876,N_28884,N_29350);
nand U30877 (N_30877,N_29002,N_29270);
or U30878 (N_30878,N_29329,N_28858);
nand U30879 (N_30879,N_29287,N_29744);
nor U30880 (N_30880,N_28338,N_28938);
and U30881 (N_30881,N_28336,N_28218);
or U30882 (N_30882,N_29183,N_28960);
or U30883 (N_30883,N_29230,N_29140);
nor U30884 (N_30884,N_28226,N_29426);
nand U30885 (N_30885,N_29281,N_29064);
and U30886 (N_30886,N_29535,N_28728);
nand U30887 (N_30887,N_28048,N_28615);
xnor U30888 (N_30888,N_29422,N_28240);
nor U30889 (N_30889,N_29352,N_29548);
xnor U30890 (N_30890,N_28845,N_28151);
nand U30891 (N_30891,N_28437,N_28976);
and U30892 (N_30892,N_28103,N_29912);
nor U30893 (N_30893,N_29013,N_28461);
and U30894 (N_30894,N_29910,N_28876);
xor U30895 (N_30895,N_28235,N_29687);
xnor U30896 (N_30896,N_29887,N_29504);
nor U30897 (N_30897,N_28784,N_29452);
nor U30898 (N_30898,N_29871,N_28209);
and U30899 (N_30899,N_28896,N_29883);
xor U30900 (N_30900,N_28242,N_29905);
or U30901 (N_30901,N_28945,N_29207);
nand U30902 (N_30902,N_29220,N_29216);
nor U30903 (N_30903,N_29026,N_29460);
nand U30904 (N_30904,N_29041,N_29842);
nand U30905 (N_30905,N_28372,N_29797);
nor U30906 (N_30906,N_28147,N_28274);
xor U30907 (N_30907,N_28809,N_29169);
or U30908 (N_30908,N_28142,N_28646);
nand U30909 (N_30909,N_28044,N_29906);
xnor U30910 (N_30910,N_28589,N_29028);
xnor U30911 (N_30911,N_28971,N_29772);
or U30912 (N_30912,N_29650,N_28778);
xnor U30913 (N_30913,N_28265,N_28940);
nand U30914 (N_30914,N_28899,N_28735);
nor U30915 (N_30915,N_28102,N_29343);
nor U30916 (N_30916,N_29167,N_29307);
and U30917 (N_30917,N_28700,N_29955);
xnor U30918 (N_30918,N_29272,N_28310);
or U30919 (N_30919,N_28322,N_28233);
xor U30920 (N_30920,N_28897,N_28793);
xor U30921 (N_30921,N_28754,N_28630);
nor U30922 (N_30922,N_28652,N_28997);
nand U30923 (N_30923,N_29447,N_29977);
or U30924 (N_30924,N_28775,N_28539);
nor U30925 (N_30925,N_28309,N_28642);
xnor U30926 (N_30926,N_28157,N_29523);
or U30927 (N_30927,N_29855,N_29543);
or U30928 (N_30928,N_29710,N_28967);
xnor U30929 (N_30929,N_29512,N_28517);
and U30930 (N_30930,N_29074,N_28758);
nand U30931 (N_30931,N_29502,N_28234);
and U30932 (N_30932,N_29720,N_28275);
nor U30933 (N_30933,N_29440,N_29338);
or U30934 (N_30934,N_29075,N_29668);
nand U30935 (N_30935,N_29990,N_28801);
xor U30936 (N_30936,N_29142,N_28327);
nand U30937 (N_30937,N_28587,N_29608);
and U30938 (N_30938,N_28666,N_28115);
or U30939 (N_30939,N_28496,N_29277);
nand U30940 (N_30940,N_29967,N_29008);
or U30941 (N_30941,N_29450,N_28663);
nand U30942 (N_30942,N_29323,N_29588);
nor U30943 (N_30943,N_29341,N_28444);
xor U30944 (N_30944,N_29874,N_28597);
nor U30945 (N_30945,N_28644,N_29144);
xnor U30946 (N_30946,N_29170,N_28732);
nand U30947 (N_30947,N_29589,N_28383);
xor U30948 (N_30948,N_29848,N_29092);
xnor U30949 (N_30949,N_29315,N_29555);
xnor U30950 (N_30950,N_28211,N_28843);
xor U30951 (N_30951,N_29406,N_28535);
nor U30952 (N_30952,N_29486,N_29049);
xor U30953 (N_30953,N_28825,N_29779);
nor U30954 (N_30954,N_28349,N_29798);
nor U30955 (N_30955,N_29035,N_28289);
xnor U30956 (N_30956,N_29709,N_29124);
or U30957 (N_30957,N_28683,N_28092);
or U30958 (N_30958,N_28393,N_29096);
xnor U30959 (N_30959,N_29114,N_29360);
or U30960 (N_30960,N_28149,N_28699);
or U30961 (N_30961,N_29444,N_29320);
or U30962 (N_30962,N_29383,N_28757);
and U30963 (N_30963,N_29163,N_29279);
nor U30964 (N_30964,N_29771,N_29951);
or U30965 (N_30965,N_28080,N_28740);
xor U30966 (N_30966,N_29576,N_28126);
nor U30967 (N_30967,N_29247,N_28923);
nor U30968 (N_30968,N_29928,N_28941);
nor U30969 (N_30969,N_28158,N_28396);
and U30970 (N_30970,N_28545,N_28921);
and U30971 (N_30971,N_28512,N_28656);
nor U30972 (N_30972,N_28772,N_28717);
nor U30973 (N_30973,N_28824,N_29606);
xnor U30974 (N_30974,N_29661,N_29226);
xnor U30975 (N_30975,N_28360,N_29914);
nand U30976 (N_30976,N_28810,N_29141);
xor U30977 (N_30977,N_29538,N_29574);
or U30978 (N_30978,N_28603,N_28171);
xor U30979 (N_30979,N_29747,N_28974);
nor U30980 (N_30980,N_28281,N_28424);
and U30981 (N_30981,N_29639,N_29500);
xnor U30982 (N_30982,N_29593,N_28746);
nor U30983 (N_30983,N_28965,N_28101);
and U30984 (N_30984,N_29480,N_29791);
nor U30985 (N_30985,N_28838,N_28258);
and U30986 (N_30986,N_29195,N_29991);
xnor U30987 (N_30987,N_28873,N_29222);
or U30988 (N_30988,N_28341,N_28358);
nor U30989 (N_30989,N_29007,N_29983);
xnor U30990 (N_30990,N_29572,N_28350);
and U30991 (N_30991,N_29494,N_28047);
xor U30992 (N_30992,N_29133,N_28034);
or U30993 (N_30993,N_28052,N_29786);
nor U30994 (N_30994,N_29359,N_29627);
nor U30995 (N_30995,N_29729,N_29251);
and U30996 (N_30996,N_28767,N_29403);
nand U30997 (N_30997,N_28650,N_28066);
or U30998 (N_30998,N_29904,N_28632);
nor U30999 (N_30999,N_29437,N_29185);
xnor U31000 (N_31000,N_28135,N_29222);
xnor U31001 (N_31001,N_29845,N_28308);
or U31002 (N_31002,N_29383,N_28626);
nand U31003 (N_31003,N_29127,N_29031);
nand U31004 (N_31004,N_28115,N_29502);
xor U31005 (N_31005,N_29544,N_28282);
nor U31006 (N_31006,N_28699,N_29785);
nand U31007 (N_31007,N_28893,N_28152);
or U31008 (N_31008,N_28525,N_29576);
or U31009 (N_31009,N_29521,N_28799);
nor U31010 (N_31010,N_28131,N_28211);
and U31011 (N_31011,N_28181,N_29218);
nand U31012 (N_31012,N_28020,N_29355);
nor U31013 (N_31013,N_28440,N_28570);
xnor U31014 (N_31014,N_29638,N_29505);
xnor U31015 (N_31015,N_29326,N_29251);
and U31016 (N_31016,N_29857,N_28867);
xor U31017 (N_31017,N_28276,N_28577);
nor U31018 (N_31018,N_29035,N_29385);
nor U31019 (N_31019,N_28985,N_28505);
nor U31020 (N_31020,N_28946,N_28034);
nor U31021 (N_31021,N_29955,N_28948);
nand U31022 (N_31022,N_29937,N_29458);
nor U31023 (N_31023,N_29644,N_29344);
or U31024 (N_31024,N_28767,N_28276);
nor U31025 (N_31025,N_29049,N_28012);
or U31026 (N_31026,N_29288,N_29926);
and U31027 (N_31027,N_28509,N_29996);
xor U31028 (N_31028,N_29675,N_28660);
nor U31029 (N_31029,N_29015,N_28950);
xor U31030 (N_31030,N_29154,N_29296);
xor U31031 (N_31031,N_28585,N_28599);
xor U31032 (N_31032,N_29970,N_29478);
nor U31033 (N_31033,N_28981,N_29462);
nor U31034 (N_31034,N_29708,N_28331);
nand U31035 (N_31035,N_28616,N_28425);
xor U31036 (N_31036,N_28097,N_28665);
nand U31037 (N_31037,N_28170,N_28747);
or U31038 (N_31038,N_29139,N_28725);
and U31039 (N_31039,N_28891,N_28915);
nor U31040 (N_31040,N_29640,N_28079);
and U31041 (N_31041,N_28476,N_28984);
and U31042 (N_31042,N_28860,N_28368);
or U31043 (N_31043,N_29176,N_29731);
nor U31044 (N_31044,N_28969,N_28749);
xnor U31045 (N_31045,N_29181,N_29070);
and U31046 (N_31046,N_29460,N_28520);
or U31047 (N_31047,N_28252,N_28368);
or U31048 (N_31048,N_28008,N_29480);
nor U31049 (N_31049,N_29580,N_29961);
nand U31050 (N_31050,N_28284,N_28828);
xor U31051 (N_31051,N_28180,N_29808);
nor U31052 (N_31052,N_29360,N_29134);
and U31053 (N_31053,N_29205,N_28232);
nor U31054 (N_31054,N_29273,N_29259);
xor U31055 (N_31055,N_29356,N_29437);
nand U31056 (N_31056,N_28794,N_29764);
xor U31057 (N_31057,N_29991,N_28089);
xor U31058 (N_31058,N_29147,N_29735);
xnor U31059 (N_31059,N_28049,N_28508);
nor U31060 (N_31060,N_28950,N_29903);
and U31061 (N_31061,N_28205,N_28313);
or U31062 (N_31062,N_28232,N_29907);
or U31063 (N_31063,N_28921,N_28796);
xnor U31064 (N_31064,N_29247,N_29264);
and U31065 (N_31065,N_29585,N_28161);
and U31066 (N_31066,N_29270,N_28902);
nand U31067 (N_31067,N_28159,N_29861);
nand U31068 (N_31068,N_29542,N_29892);
nand U31069 (N_31069,N_28676,N_28175);
and U31070 (N_31070,N_29557,N_28006);
or U31071 (N_31071,N_28197,N_28607);
nand U31072 (N_31072,N_28550,N_28522);
nor U31073 (N_31073,N_29733,N_29979);
or U31074 (N_31074,N_28883,N_29839);
or U31075 (N_31075,N_29588,N_29382);
nor U31076 (N_31076,N_28972,N_29824);
xor U31077 (N_31077,N_29499,N_29804);
xor U31078 (N_31078,N_28444,N_28521);
xnor U31079 (N_31079,N_29314,N_29573);
or U31080 (N_31080,N_28779,N_29102);
xnor U31081 (N_31081,N_29593,N_29224);
xnor U31082 (N_31082,N_28533,N_28739);
nand U31083 (N_31083,N_28522,N_29674);
nor U31084 (N_31084,N_29763,N_28199);
xnor U31085 (N_31085,N_29903,N_29424);
xnor U31086 (N_31086,N_28592,N_29626);
xnor U31087 (N_31087,N_28094,N_29779);
and U31088 (N_31088,N_28125,N_29939);
and U31089 (N_31089,N_28304,N_28010);
and U31090 (N_31090,N_29574,N_28063);
and U31091 (N_31091,N_28754,N_28390);
nor U31092 (N_31092,N_29038,N_28358);
nand U31093 (N_31093,N_29446,N_28221);
nor U31094 (N_31094,N_29827,N_29137);
and U31095 (N_31095,N_28722,N_29952);
xnor U31096 (N_31096,N_29502,N_29839);
nor U31097 (N_31097,N_28017,N_29198);
and U31098 (N_31098,N_28971,N_28224);
or U31099 (N_31099,N_29391,N_28161);
or U31100 (N_31100,N_28778,N_29464);
xor U31101 (N_31101,N_29329,N_28774);
nand U31102 (N_31102,N_28896,N_28130);
xor U31103 (N_31103,N_28806,N_29250);
xor U31104 (N_31104,N_28330,N_29963);
or U31105 (N_31105,N_29566,N_29316);
or U31106 (N_31106,N_28392,N_29393);
and U31107 (N_31107,N_28287,N_28888);
nand U31108 (N_31108,N_28102,N_28012);
or U31109 (N_31109,N_28895,N_28923);
or U31110 (N_31110,N_29490,N_28270);
nand U31111 (N_31111,N_29436,N_28318);
xor U31112 (N_31112,N_29940,N_29479);
xor U31113 (N_31113,N_29610,N_29433);
or U31114 (N_31114,N_28369,N_28872);
nand U31115 (N_31115,N_28906,N_28549);
nor U31116 (N_31116,N_28568,N_28144);
nor U31117 (N_31117,N_29310,N_29489);
or U31118 (N_31118,N_28248,N_28937);
nor U31119 (N_31119,N_28062,N_28600);
or U31120 (N_31120,N_28868,N_28095);
xor U31121 (N_31121,N_29505,N_29318);
nor U31122 (N_31122,N_29824,N_28063);
xor U31123 (N_31123,N_29311,N_29952);
nor U31124 (N_31124,N_29360,N_29290);
or U31125 (N_31125,N_29580,N_29143);
nor U31126 (N_31126,N_29313,N_29007);
xor U31127 (N_31127,N_29518,N_28620);
nand U31128 (N_31128,N_29755,N_29599);
or U31129 (N_31129,N_28451,N_29330);
xnor U31130 (N_31130,N_28221,N_28200);
nor U31131 (N_31131,N_29557,N_29723);
and U31132 (N_31132,N_28685,N_29927);
or U31133 (N_31133,N_28252,N_28549);
and U31134 (N_31134,N_29457,N_29561);
or U31135 (N_31135,N_28462,N_28315);
xnor U31136 (N_31136,N_28291,N_28445);
xnor U31137 (N_31137,N_28159,N_28359);
nand U31138 (N_31138,N_28704,N_28682);
and U31139 (N_31139,N_29953,N_29931);
and U31140 (N_31140,N_29111,N_29462);
xor U31141 (N_31141,N_29645,N_29997);
or U31142 (N_31142,N_28610,N_29015);
or U31143 (N_31143,N_29182,N_28324);
nand U31144 (N_31144,N_28064,N_28409);
and U31145 (N_31145,N_29446,N_28961);
xor U31146 (N_31146,N_28285,N_28978);
nand U31147 (N_31147,N_29167,N_28157);
xor U31148 (N_31148,N_29624,N_29779);
or U31149 (N_31149,N_28275,N_28340);
and U31150 (N_31150,N_28270,N_28067);
nand U31151 (N_31151,N_29401,N_28143);
nor U31152 (N_31152,N_28020,N_29443);
and U31153 (N_31153,N_29304,N_29286);
or U31154 (N_31154,N_28853,N_28247);
or U31155 (N_31155,N_28418,N_29945);
nand U31156 (N_31156,N_29893,N_29332);
nor U31157 (N_31157,N_28349,N_29369);
nor U31158 (N_31158,N_28564,N_29585);
and U31159 (N_31159,N_28449,N_28409);
or U31160 (N_31160,N_29844,N_28398);
or U31161 (N_31161,N_28714,N_28171);
or U31162 (N_31162,N_28289,N_29066);
and U31163 (N_31163,N_29186,N_29362);
nor U31164 (N_31164,N_28873,N_28001);
xnor U31165 (N_31165,N_29078,N_28976);
nor U31166 (N_31166,N_29903,N_28046);
xor U31167 (N_31167,N_28103,N_29900);
xnor U31168 (N_31168,N_29205,N_28962);
nand U31169 (N_31169,N_29552,N_28777);
nor U31170 (N_31170,N_28992,N_28125);
or U31171 (N_31171,N_29520,N_28502);
and U31172 (N_31172,N_28591,N_29158);
and U31173 (N_31173,N_29417,N_29028);
or U31174 (N_31174,N_28940,N_28053);
and U31175 (N_31175,N_28107,N_28339);
nand U31176 (N_31176,N_28510,N_28853);
nand U31177 (N_31177,N_29880,N_29616);
xnor U31178 (N_31178,N_29877,N_29550);
nor U31179 (N_31179,N_29233,N_29468);
and U31180 (N_31180,N_29883,N_29870);
nor U31181 (N_31181,N_28815,N_29567);
xnor U31182 (N_31182,N_29638,N_29696);
nor U31183 (N_31183,N_28446,N_28496);
xor U31184 (N_31184,N_29809,N_28088);
nand U31185 (N_31185,N_29795,N_28198);
nand U31186 (N_31186,N_28885,N_29457);
xor U31187 (N_31187,N_28200,N_29954);
or U31188 (N_31188,N_29105,N_28867);
or U31189 (N_31189,N_29397,N_29725);
or U31190 (N_31190,N_28799,N_28404);
or U31191 (N_31191,N_28417,N_28856);
nand U31192 (N_31192,N_28785,N_28806);
nor U31193 (N_31193,N_29806,N_28494);
or U31194 (N_31194,N_29636,N_28174);
xor U31195 (N_31195,N_29877,N_28605);
nand U31196 (N_31196,N_29930,N_29386);
nand U31197 (N_31197,N_28570,N_28790);
or U31198 (N_31198,N_29404,N_28910);
or U31199 (N_31199,N_29029,N_28121);
nor U31200 (N_31200,N_29452,N_29809);
nand U31201 (N_31201,N_29353,N_29713);
nand U31202 (N_31202,N_29267,N_29315);
nand U31203 (N_31203,N_29189,N_29292);
and U31204 (N_31204,N_29753,N_29151);
nor U31205 (N_31205,N_29489,N_28012);
nor U31206 (N_31206,N_28487,N_28454);
or U31207 (N_31207,N_28635,N_29436);
nor U31208 (N_31208,N_28118,N_28515);
nor U31209 (N_31209,N_28579,N_28219);
nor U31210 (N_31210,N_28646,N_28224);
xor U31211 (N_31211,N_29147,N_29684);
and U31212 (N_31212,N_28886,N_29020);
and U31213 (N_31213,N_28578,N_29869);
xnor U31214 (N_31214,N_28923,N_29255);
or U31215 (N_31215,N_28907,N_29696);
or U31216 (N_31216,N_28456,N_29929);
nand U31217 (N_31217,N_28923,N_29982);
nand U31218 (N_31218,N_29341,N_28849);
nor U31219 (N_31219,N_29680,N_28633);
and U31220 (N_31220,N_29574,N_28447);
xor U31221 (N_31221,N_28263,N_28907);
nor U31222 (N_31222,N_28660,N_28628);
or U31223 (N_31223,N_29275,N_29671);
or U31224 (N_31224,N_28869,N_29472);
nor U31225 (N_31225,N_29629,N_29115);
nor U31226 (N_31226,N_28259,N_29365);
xnor U31227 (N_31227,N_29406,N_28410);
xor U31228 (N_31228,N_29960,N_28565);
and U31229 (N_31229,N_29709,N_28871);
or U31230 (N_31230,N_29237,N_28975);
nor U31231 (N_31231,N_28290,N_29681);
nor U31232 (N_31232,N_28495,N_29588);
and U31233 (N_31233,N_29226,N_28472);
nand U31234 (N_31234,N_28153,N_28005);
or U31235 (N_31235,N_28844,N_29323);
nand U31236 (N_31236,N_28986,N_28656);
nor U31237 (N_31237,N_28667,N_29870);
nor U31238 (N_31238,N_29539,N_28501);
nand U31239 (N_31239,N_29370,N_28401);
nand U31240 (N_31240,N_28318,N_29465);
nor U31241 (N_31241,N_29853,N_28597);
nand U31242 (N_31242,N_29070,N_29872);
nor U31243 (N_31243,N_29850,N_28549);
xor U31244 (N_31244,N_29687,N_29652);
xnor U31245 (N_31245,N_29843,N_28764);
and U31246 (N_31246,N_28863,N_28345);
nor U31247 (N_31247,N_28078,N_29104);
xnor U31248 (N_31248,N_28245,N_29609);
xor U31249 (N_31249,N_29008,N_28646);
nand U31250 (N_31250,N_29084,N_29546);
nor U31251 (N_31251,N_29926,N_28541);
nand U31252 (N_31252,N_28201,N_28978);
xor U31253 (N_31253,N_28711,N_28521);
xnor U31254 (N_31254,N_28698,N_28578);
nor U31255 (N_31255,N_29540,N_28372);
or U31256 (N_31256,N_28938,N_28323);
or U31257 (N_31257,N_29383,N_29009);
nand U31258 (N_31258,N_29965,N_29591);
nand U31259 (N_31259,N_28653,N_28617);
and U31260 (N_31260,N_29653,N_28400);
or U31261 (N_31261,N_28695,N_28332);
and U31262 (N_31262,N_28991,N_28936);
nor U31263 (N_31263,N_29637,N_28030);
nor U31264 (N_31264,N_28663,N_28399);
or U31265 (N_31265,N_28612,N_29459);
nor U31266 (N_31266,N_29229,N_28262);
nand U31267 (N_31267,N_28394,N_28090);
or U31268 (N_31268,N_29178,N_28990);
nand U31269 (N_31269,N_28983,N_29686);
nor U31270 (N_31270,N_28891,N_28736);
nand U31271 (N_31271,N_28249,N_29727);
and U31272 (N_31272,N_28239,N_28424);
nor U31273 (N_31273,N_29090,N_29970);
nor U31274 (N_31274,N_28839,N_29350);
xnor U31275 (N_31275,N_29066,N_28676);
nand U31276 (N_31276,N_28305,N_28715);
nand U31277 (N_31277,N_28238,N_29314);
nand U31278 (N_31278,N_28669,N_29257);
or U31279 (N_31279,N_28782,N_29771);
or U31280 (N_31280,N_28739,N_28471);
nand U31281 (N_31281,N_28045,N_29503);
nor U31282 (N_31282,N_29422,N_28970);
or U31283 (N_31283,N_28254,N_29548);
nor U31284 (N_31284,N_29835,N_29564);
nor U31285 (N_31285,N_29108,N_29825);
or U31286 (N_31286,N_28363,N_29438);
or U31287 (N_31287,N_28233,N_28906);
and U31288 (N_31288,N_28717,N_28739);
xor U31289 (N_31289,N_29411,N_28459);
nand U31290 (N_31290,N_28723,N_29726);
xor U31291 (N_31291,N_28078,N_29924);
and U31292 (N_31292,N_29609,N_28109);
nand U31293 (N_31293,N_28158,N_28114);
nand U31294 (N_31294,N_28696,N_28306);
and U31295 (N_31295,N_29729,N_28674);
xor U31296 (N_31296,N_28363,N_29910);
xnor U31297 (N_31297,N_29111,N_29320);
nand U31298 (N_31298,N_29649,N_29285);
nor U31299 (N_31299,N_28765,N_29390);
and U31300 (N_31300,N_28046,N_28585);
xor U31301 (N_31301,N_29305,N_29096);
or U31302 (N_31302,N_28831,N_29043);
and U31303 (N_31303,N_29303,N_28668);
and U31304 (N_31304,N_28680,N_29368);
nor U31305 (N_31305,N_29227,N_29228);
and U31306 (N_31306,N_28526,N_28371);
nor U31307 (N_31307,N_28221,N_28164);
xnor U31308 (N_31308,N_28794,N_29181);
or U31309 (N_31309,N_29248,N_29971);
xnor U31310 (N_31310,N_29130,N_29118);
and U31311 (N_31311,N_29595,N_29355);
or U31312 (N_31312,N_29023,N_28649);
or U31313 (N_31313,N_28296,N_29606);
or U31314 (N_31314,N_28573,N_28629);
and U31315 (N_31315,N_29989,N_28105);
nand U31316 (N_31316,N_29815,N_28027);
or U31317 (N_31317,N_29274,N_28912);
or U31318 (N_31318,N_29036,N_29101);
or U31319 (N_31319,N_28758,N_29912);
nand U31320 (N_31320,N_28985,N_29630);
xnor U31321 (N_31321,N_29824,N_28510);
nand U31322 (N_31322,N_28678,N_29705);
xor U31323 (N_31323,N_29720,N_29232);
nand U31324 (N_31324,N_28933,N_29994);
nand U31325 (N_31325,N_29412,N_28023);
xnor U31326 (N_31326,N_29667,N_29805);
or U31327 (N_31327,N_29517,N_28799);
nor U31328 (N_31328,N_29109,N_29905);
nor U31329 (N_31329,N_28513,N_29846);
xor U31330 (N_31330,N_28669,N_28742);
or U31331 (N_31331,N_29315,N_28760);
or U31332 (N_31332,N_29865,N_28174);
or U31333 (N_31333,N_28084,N_28274);
nor U31334 (N_31334,N_28996,N_28737);
nor U31335 (N_31335,N_28399,N_28962);
nor U31336 (N_31336,N_28726,N_28456);
nand U31337 (N_31337,N_28704,N_29248);
nand U31338 (N_31338,N_28036,N_29249);
nand U31339 (N_31339,N_29284,N_28468);
xnor U31340 (N_31340,N_28089,N_29016);
nor U31341 (N_31341,N_28365,N_28836);
nand U31342 (N_31342,N_28967,N_28863);
and U31343 (N_31343,N_28959,N_28800);
xnor U31344 (N_31344,N_29019,N_29422);
nor U31345 (N_31345,N_28981,N_28208);
nand U31346 (N_31346,N_29154,N_28603);
and U31347 (N_31347,N_28965,N_28322);
nand U31348 (N_31348,N_28810,N_29730);
nand U31349 (N_31349,N_28967,N_28544);
and U31350 (N_31350,N_28217,N_29728);
xor U31351 (N_31351,N_28281,N_29007);
nand U31352 (N_31352,N_29810,N_29747);
nand U31353 (N_31353,N_28339,N_28210);
nand U31354 (N_31354,N_28831,N_29761);
or U31355 (N_31355,N_28566,N_29566);
nand U31356 (N_31356,N_29652,N_28945);
nor U31357 (N_31357,N_29873,N_28302);
xnor U31358 (N_31358,N_29661,N_29731);
nand U31359 (N_31359,N_29931,N_28428);
or U31360 (N_31360,N_29489,N_28689);
or U31361 (N_31361,N_29101,N_29675);
or U31362 (N_31362,N_28513,N_29339);
and U31363 (N_31363,N_28392,N_28137);
and U31364 (N_31364,N_29768,N_29931);
nor U31365 (N_31365,N_29554,N_29509);
xnor U31366 (N_31366,N_28223,N_29487);
nand U31367 (N_31367,N_28413,N_28577);
or U31368 (N_31368,N_28089,N_28933);
nor U31369 (N_31369,N_29143,N_28195);
and U31370 (N_31370,N_28301,N_28238);
and U31371 (N_31371,N_28175,N_29608);
xnor U31372 (N_31372,N_28406,N_28223);
and U31373 (N_31373,N_29457,N_29255);
nand U31374 (N_31374,N_29168,N_28472);
nand U31375 (N_31375,N_28829,N_29208);
and U31376 (N_31376,N_28207,N_28638);
xnor U31377 (N_31377,N_28329,N_28808);
nor U31378 (N_31378,N_29029,N_29138);
or U31379 (N_31379,N_28619,N_29259);
xnor U31380 (N_31380,N_29586,N_29275);
xnor U31381 (N_31381,N_29728,N_29475);
nor U31382 (N_31382,N_28257,N_28283);
nand U31383 (N_31383,N_29463,N_28243);
nor U31384 (N_31384,N_28916,N_28423);
or U31385 (N_31385,N_28525,N_28543);
and U31386 (N_31386,N_28524,N_28628);
and U31387 (N_31387,N_28049,N_28398);
nand U31388 (N_31388,N_28034,N_29514);
or U31389 (N_31389,N_29354,N_28924);
and U31390 (N_31390,N_28183,N_29322);
nand U31391 (N_31391,N_28761,N_29905);
nand U31392 (N_31392,N_29727,N_28672);
or U31393 (N_31393,N_28223,N_29242);
and U31394 (N_31394,N_28650,N_29189);
and U31395 (N_31395,N_28437,N_28125);
nor U31396 (N_31396,N_29875,N_28873);
or U31397 (N_31397,N_28941,N_29871);
and U31398 (N_31398,N_28121,N_28300);
or U31399 (N_31399,N_28671,N_29734);
or U31400 (N_31400,N_28118,N_29895);
or U31401 (N_31401,N_28530,N_29420);
and U31402 (N_31402,N_29056,N_28365);
nor U31403 (N_31403,N_28781,N_29535);
and U31404 (N_31404,N_29212,N_29149);
or U31405 (N_31405,N_29179,N_29875);
and U31406 (N_31406,N_28092,N_28421);
xor U31407 (N_31407,N_28538,N_28009);
nor U31408 (N_31408,N_29101,N_28589);
and U31409 (N_31409,N_29132,N_29789);
xnor U31410 (N_31410,N_29328,N_28281);
xor U31411 (N_31411,N_28682,N_28270);
or U31412 (N_31412,N_28937,N_28623);
and U31413 (N_31413,N_29177,N_29774);
nand U31414 (N_31414,N_28013,N_28709);
nand U31415 (N_31415,N_29623,N_29507);
xor U31416 (N_31416,N_28321,N_28376);
nor U31417 (N_31417,N_29734,N_29175);
or U31418 (N_31418,N_28417,N_29627);
xor U31419 (N_31419,N_29002,N_29530);
xor U31420 (N_31420,N_28667,N_29318);
and U31421 (N_31421,N_29092,N_29569);
or U31422 (N_31422,N_28459,N_29168);
nand U31423 (N_31423,N_29440,N_28299);
or U31424 (N_31424,N_29617,N_28745);
nor U31425 (N_31425,N_28234,N_28869);
and U31426 (N_31426,N_29844,N_28327);
and U31427 (N_31427,N_29333,N_29120);
or U31428 (N_31428,N_28348,N_28236);
xor U31429 (N_31429,N_29510,N_28436);
and U31430 (N_31430,N_29420,N_29847);
xor U31431 (N_31431,N_28202,N_29648);
nor U31432 (N_31432,N_28983,N_28361);
and U31433 (N_31433,N_28466,N_29275);
nand U31434 (N_31434,N_29753,N_29619);
nor U31435 (N_31435,N_29604,N_28704);
nand U31436 (N_31436,N_28603,N_29998);
and U31437 (N_31437,N_29284,N_28917);
xnor U31438 (N_31438,N_28319,N_28112);
nand U31439 (N_31439,N_29123,N_28632);
or U31440 (N_31440,N_29549,N_28721);
nand U31441 (N_31441,N_29840,N_28041);
nor U31442 (N_31442,N_28434,N_29032);
xnor U31443 (N_31443,N_28002,N_28734);
nand U31444 (N_31444,N_28898,N_29674);
xnor U31445 (N_31445,N_29321,N_29383);
or U31446 (N_31446,N_28191,N_28767);
xor U31447 (N_31447,N_29435,N_28548);
and U31448 (N_31448,N_29244,N_28079);
or U31449 (N_31449,N_29675,N_29122);
xor U31450 (N_31450,N_28244,N_29150);
nand U31451 (N_31451,N_29854,N_29576);
and U31452 (N_31452,N_28344,N_28434);
and U31453 (N_31453,N_29893,N_28781);
nor U31454 (N_31454,N_28142,N_29627);
or U31455 (N_31455,N_28063,N_28402);
nor U31456 (N_31456,N_28972,N_29898);
xnor U31457 (N_31457,N_28100,N_28401);
or U31458 (N_31458,N_28214,N_28121);
nand U31459 (N_31459,N_28979,N_28814);
nand U31460 (N_31460,N_29787,N_29665);
xnor U31461 (N_31461,N_28444,N_28620);
nand U31462 (N_31462,N_28698,N_28651);
nor U31463 (N_31463,N_29543,N_28138);
and U31464 (N_31464,N_29913,N_28010);
and U31465 (N_31465,N_29700,N_28388);
nand U31466 (N_31466,N_28433,N_28096);
and U31467 (N_31467,N_29095,N_28434);
nand U31468 (N_31468,N_28943,N_29138);
or U31469 (N_31469,N_29064,N_28818);
and U31470 (N_31470,N_29062,N_28001);
or U31471 (N_31471,N_28901,N_29556);
nand U31472 (N_31472,N_29016,N_28863);
or U31473 (N_31473,N_28814,N_28707);
and U31474 (N_31474,N_29886,N_28551);
nand U31475 (N_31475,N_29561,N_28315);
or U31476 (N_31476,N_29865,N_29778);
and U31477 (N_31477,N_28124,N_28734);
nor U31478 (N_31478,N_29748,N_29299);
xnor U31479 (N_31479,N_28298,N_29072);
nor U31480 (N_31480,N_29979,N_28929);
xnor U31481 (N_31481,N_28584,N_29543);
xor U31482 (N_31482,N_29890,N_28236);
nand U31483 (N_31483,N_28904,N_29601);
nand U31484 (N_31484,N_28712,N_28743);
and U31485 (N_31485,N_28966,N_28901);
xnor U31486 (N_31486,N_28956,N_28429);
nand U31487 (N_31487,N_28063,N_28632);
or U31488 (N_31488,N_29823,N_28713);
nor U31489 (N_31489,N_28991,N_29980);
xor U31490 (N_31490,N_29368,N_29799);
nor U31491 (N_31491,N_29360,N_28549);
xor U31492 (N_31492,N_28213,N_28339);
and U31493 (N_31493,N_28337,N_28103);
or U31494 (N_31494,N_29723,N_28025);
nand U31495 (N_31495,N_29597,N_28873);
or U31496 (N_31496,N_29949,N_29638);
nor U31497 (N_31497,N_29035,N_28797);
and U31498 (N_31498,N_28712,N_29367);
nand U31499 (N_31499,N_28254,N_29895);
nand U31500 (N_31500,N_29909,N_29735);
or U31501 (N_31501,N_28220,N_29298);
or U31502 (N_31502,N_28517,N_29598);
xor U31503 (N_31503,N_28915,N_29311);
nor U31504 (N_31504,N_29877,N_28099);
nand U31505 (N_31505,N_28512,N_29657);
and U31506 (N_31506,N_29813,N_28088);
xor U31507 (N_31507,N_29248,N_29389);
nand U31508 (N_31508,N_29089,N_28332);
nor U31509 (N_31509,N_28918,N_29725);
nand U31510 (N_31510,N_29851,N_28823);
xnor U31511 (N_31511,N_29571,N_29329);
nand U31512 (N_31512,N_29683,N_29167);
or U31513 (N_31513,N_29394,N_28364);
nor U31514 (N_31514,N_28997,N_28996);
nand U31515 (N_31515,N_29448,N_29980);
nor U31516 (N_31516,N_28949,N_29488);
or U31517 (N_31517,N_29637,N_29972);
nor U31518 (N_31518,N_29704,N_29376);
and U31519 (N_31519,N_29108,N_28896);
nor U31520 (N_31520,N_29100,N_28108);
or U31521 (N_31521,N_28144,N_28479);
nor U31522 (N_31522,N_29994,N_29262);
nand U31523 (N_31523,N_29644,N_28563);
or U31524 (N_31524,N_29574,N_28774);
or U31525 (N_31525,N_29640,N_29225);
xnor U31526 (N_31526,N_28606,N_28153);
nand U31527 (N_31527,N_29391,N_28261);
nor U31528 (N_31528,N_29272,N_29051);
xor U31529 (N_31529,N_29951,N_28960);
xor U31530 (N_31530,N_28743,N_29132);
or U31531 (N_31531,N_28078,N_29365);
nand U31532 (N_31532,N_28053,N_28135);
and U31533 (N_31533,N_28470,N_29623);
xor U31534 (N_31534,N_28156,N_28737);
or U31535 (N_31535,N_29550,N_28681);
nor U31536 (N_31536,N_28278,N_28135);
nor U31537 (N_31537,N_29972,N_28670);
nand U31538 (N_31538,N_29182,N_29130);
and U31539 (N_31539,N_29135,N_29285);
and U31540 (N_31540,N_28478,N_28664);
xnor U31541 (N_31541,N_28264,N_29185);
nor U31542 (N_31542,N_29726,N_28172);
nor U31543 (N_31543,N_28803,N_28987);
or U31544 (N_31544,N_29487,N_29545);
xor U31545 (N_31545,N_28140,N_29347);
xnor U31546 (N_31546,N_29824,N_28372);
or U31547 (N_31547,N_28226,N_29588);
or U31548 (N_31548,N_28976,N_29063);
or U31549 (N_31549,N_29642,N_28578);
nor U31550 (N_31550,N_29855,N_28441);
xnor U31551 (N_31551,N_29938,N_29414);
nand U31552 (N_31552,N_29987,N_28197);
and U31553 (N_31553,N_29107,N_29263);
xor U31554 (N_31554,N_28326,N_28426);
nor U31555 (N_31555,N_28316,N_29451);
and U31556 (N_31556,N_28682,N_28257);
xnor U31557 (N_31557,N_29403,N_29272);
or U31558 (N_31558,N_29565,N_28405);
nor U31559 (N_31559,N_29997,N_28314);
xor U31560 (N_31560,N_29744,N_29614);
nor U31561 (N_31561,N_29323,N_28895);
nor U31562 (N_31562,N_29784,N_28261);
and U31563 (N_31563,N_28483,N_29827);
and U31564 (N_31564,N_29451,N_28256);
nand U31565 (N_31565,N_28086,N_29501);
or U31566 (N_31566,N_28522,N_29174);
nand U31567 (N_31567,N_29797,N_28712);
nor U31568 (N_31568,N_29283,N_28485);
or U31569 (N_31569,N_28972,N_29770);
nand U31570 (N_31570,N_28288,N_29820);
and U31571 (N_31571,N_28731,N_29290);
nor U31572 (N_31572,N_29579,N_29302);
or U31573 (N_31573,N_29616,N_29991);
and U31574 (N_31574,N_29113,N_29227);
or U31575 (N_31575,N_29410,N_28622);
nand U31576 (N_31576,N_29284,N_28123);
nand U31577 (N_31577,N_29164,N_28207);
nor U31578 (N_31578,N_28323,N_28034);
or U31579 (N_31579,N_29215,N_28898);
nand U31580 (N_31580,N_29409,N_29435);
nor U31581 (N_31581,N_29960,N_28120);
nor U31582 (N_31582,N_28618,N_29559);
and U31583 (N_31583,N_28029,N_28639);
xnor U31584 (N_31584,N_28712,N_29139);
nand U31585 (N_31585,N_29140,N_28438);
xnor U31586 (N_31586,N_28923,N_28343);
and U31587 (N_31587,N_29438,N_28249);
xor U31588 (N_31588,N_28866,N_29745);
xor U31589 (N_31589,N_28228,N_29834);
and U31590 (N_31590,N_29926,N_28117);
nor U31591 (N_31591,N_28552,N_29637);
nor U31592 (N_31592,N_28170,N_29409);
or U31593 (N_31593,N_29322,N_28918);
xnor U31594 (N_31594,N_29684,N_29245);
or U31595 (N_31595,N_29220,N_29643);
nor U31596 (N_31596,N_29917,N_29738);
and U31597 (N_31597,N_28687,N_28036);
nor U31598 (N_31598,N_29890,N_29582);
nor U31599 (N_31599,N_29526,N_28003);
nor U31600 (N_31600,N_29155,N_29654);
xor U31601 (N_31601,N_28267,N_29977);
or U31602 (N_31602,N_29097,N_29880);
or U31603 (N_31603,N_29333,N_28173);
nor U31604 (N_31604,N_29014,N_29270);
xnor U31605 (N_31605,N_29763,N_29891);
xor U31606 (N_31606,N_29590,N_28692);
nor U31607 (N_31607,N_29629,N_28381);
xor U31608 (N_31608,N_29688,N_28787);
xor U31609 (N_31609,N_29437,N_29514);
or U31610 (N_31610,N_29032,N_28323);
xnor U31611 (N_31611,N_29059,N_28506);
nand U31612 (N_31612,N_28627,N_29349);
nor U31613 (N_31613,N_29461,N_29011);
nor U31614 (N_31614,N_28420,N_28146);
xor U31615 (N_31615,N_29577,N_28084);
and U31616 (N_31616,N_29529,N_29459);
nor U31617 (N_31617,N_28066,N_28050);
or U31618 (N_31618,N_28767,N_29213);
or U31619 (N_31619,N_29663,N_28379);
xnor U31620 (N_31620,N_28112,N_28975);
or U31621 (N_31621,N_29773,N_29424);
xnor U31622 (N_31622,N_29746,N_29148);
and U31623 (N_31623,N_29100,N_28858);
nand U31624 (N_31624,N_28740,N_29865);
nor U31625 (N_31625,N_28071,N_28107);
xnor U31626 (N_31626,N_29679,N_29714);
nand U31627 (N_31627,N_28003,N_29904);
nand U31628 (N_31628,N_29355,N_29315);
and U31629 (N_31629,N_28393,N_28286);
and U31630 (N_31630,N_29983,N_28154);
nand U31631 (N_31631,N_28598,N_28640);
nor U31632 (N_31632,N_29614,N_29582);
xnor U31633 (N_31633,N_29347,N_28745);
nand U31634 (N_31634,N_28028,N_28802);
and U31635 (N_31635,N_28487,N_28955);
xnor U31636 (N_31636,N_29824,N_29760);
xor U31637 (N_31637,N_28626,N_28274);
or U31638 (N_31638,N_29083,N_28509);
xor U31639 (N_31639,N_28160,N_28370);
or U31640 (N_31640,N_28501,N_28868);
nand U31641 (N_31641,N_28098,N_29716);
xor U31642 (N_31642,N_29788,N_29254);
or U31643 (N_31643,N_29135,N_28309);
nand U31644 (N_31644,N_29158,N_28688);
xnor U31645 (N_31645,N_29923,N_28200);
or U31646 (N_31646,N_28460,N_29986);
nor U31647 (N_31647,N_28240,N_28782);
or U31648 (N_31648,N_29942,N_28765);
and U31649 (N_31649,N_29051,N_29312);
or U31650 (N_31650,N_29622,N_29195);
xnor U31651 (N_31651,N_29143,N_29962);
xnor U31652 (N_31652,N_28009,N_29057);
xnor U31653 (N_31653,N_28456,N_28098);
or U31654 (N_31654,N_28243,N_28848);
nor U31655 (N_31655,N_28613,N_29971);
nand U31656 (N_31656,N_28674,N_29901);
or U31657 (N_31657,N_29933,N_29261);
xnor U31658 (N_31658,N_29315,N_29410);
or U31659 (N_31659,N_29676,N_29590);
xnor U31660 (N_31660,N_29886,N_28505);
nor U31661 (N_31661,N_28177,N_28057);
xnor U31662 (N_31662,N_28237,N_29970);
or U31663 (N_31663,N_29493,N_28725);
nand U31664 (N_31664,N_29490,N_28167);
and U31665 (N_31665,N_29653,N_28999);
or U31666 (N_31666,N_28514,N_28827);
nor U31667 (N_31667,N_29341,N_28630);
xnor U31668 (N_31668,N_28104,N_28145);
and U31669 (N_31669,N_28133,N_29300);
and U31670 (N_31670,N_28355,N_29111);
or U31671 (N_31671,N_28817,N_28693);
and U31672 (N_31672,N_29843,N_29066);
and U31673 (N_31673,N_29843,N_29143);
xnor U31674 (N_31674,N_28723,N_28939);
xor U31675 (N_31675,N_29084,N_29775);
nor U31676 (N_31676,N_28881,N_29275);
or U31677 (N_31677,N_29161,N_29388);
or U31678 (N_31678,N_28636,N_28626);
nand U31679 (N_31679,N_28892,N_28493);
nor U31680 (N_31680,N_28305,N_29051);
nor U31681 (N_31681,N_28941,N_28624);
or U31682 (N_31682,N_28935,N_28667);
nor U31683 (N_31683,N_29736,N_28238);
nor U31684 (N_31684,N_28762,N_28968);
nand U31685 (N_31685,N_29451,N_29727);
or U31686 (N_31686,N_28160,N_29126);
nor U31687 (N_31687,N_29075,N_29800);
or U31688 (N_31688,N_29355,N_29240);
nand U31689 (N_31689,N_28507,N_29675);
or U31690 (N_31690,N_29948,N_28801);
nand U31691 (N_31691,N_28039,N_29605);
or U31692 (N_31692,N_28050,N_28718);
nand U31693 (N_31693,N_28761,N_29352);
nor U31694 (N_31694,N_29038,N_28087);
nand U31695 (N_31695,N_29501,N_29736);
nand U31696 (N_31696,N_28099,N_29793);
nand U31697 (N_31697,N_28974,N_28041);
nor U31698 (N_31698,N_28544,N_29608);
nand U31699 (N_31699,N_28792,N_28736);
xor U31700 (N_31700,N_28736,N_29374);
nand U31701 (N_31701,N_29591,N_29128);
and U31702 (N_31702,N_29186,N_29469);
nor U31703 (N_31703,N_29401,N_28138);
and U31704 (N_31704,N_28910,N_29637);
nor U31705 (N_31705,N_29711,N_28300);
and U31706 (N_31706,N_28965,N_29661);
and U31707 (N_31707,N_28673,N_29859);
nand U31708 (N_31708,N_28150,N_28806);
and U31709 (N_31709,N_28606,N_28394);
nor U31710 (N_31710,N_29556,N_29534);
or U31711 (N_31711,N_28234,N_29620);
nor U31712 (N_31712,N_29716,N_29770);
and U31713 (N_31713,N_29878,N_28846);
or U31714 (N_31714,N_29178,N_29411);
nor U31715 (N_31715,N_28283,N_29702);
and U31716 (N_31716,N_29396,N_28084);
xnor U31717 (N_31717,N_28508,N_28149);
and U31718 (N_31718,N_29780,N_29760);
xor U31719 (N_31719,N_29441,N_29528);
nand U31720 (N_31720,N_29296,N_29504);
nand U31721 (N_31721,N_29674,N_29746);
nor U31722 (N_31722,N_28744,N_28394);
xor U31723 (N_31723,N_29596,N_28043);
or U31724 (N_31724,N_28490,N_29029);
nor U31725 (N_31725,N_28892,N_29105);
xnor U31726 (N_31726,N_28765,N_29334);
nor U31727 (N_31727,N_28594,N_29038);
nor U31728 (N_31728,N_28984,N_28654);
xor U31729 (N_31729,N_29655,N_29934);
or U31730 (N_31730,N_29386,N_29746);
or U31731 (N_31731,N_29644,N_29786);
xor U31732 (N_31732,N_29250,N_29994);
nand U31733 (N_31733,N_29977,N_28601);
xnor U31734 (N_31734,N_29095,N_29962);
nand U31735 (N_31735,N_28836,N_29362);
nand U31736 (N_31736,N_29279,N_29012);
and U31737 (N_31737,N_29422,N_29104);
or U31738 (N_31738,N_29713,N_28679);
or U31739 (N_31739,N_28254,N_28912);
and U31740 (N_31740,N_29732,N_28571);
or U31741 (N_31741,N_29491,N_28721);
and U31742 (N_31742,N_28802,N_28378);
or U31743 (N_31743,N_29786,N_28199);
and U31744 (N_31744,N_29504,N_28576);
nor U31745 (N_31745,N_28527,N_28216);
and U31746 (N_31746,N_28324,N_29216);
nand U31747 (N_31747,N_29883,N_29155);
nand U31748 (N_31748,N_28157,N_28442);
or U31749 (N_31749,N_28698,N_29776);
xor U31750 (N_31750,N_29838,N_28540);
nor U31751 (N_31751,N_28017,N_28303);
and U31752 (N_31752,N_28106,N_29439);
nand U31753 (N_31753,N_28630,N_28281);
and U31754 (N_31754,N_28047,N_28500);
nor U31755 (N_31755,N_28870,N_28189);
or U31756 (N_31756,N_28146,N_29346);
nand U31757 (N_31757,N_29561,N_28482);
nor U31758 (N_31758,N_29232,N_29377);
nand U31759 (N_31759,N_28986,N_29965);
nor U31760 (N_31760,N_28788,N_29289);
or U31761 (N_31761,N_29001,N_28839);
xor U31762 (N_31762,N_29972,N_28295);
xor U31763 (N_31763,N_28958,N_28480);
or U31764 (N_31764,N_28335,N_28570);
or U31765 (N_31765,N_29300,N_29185);
xor U31766 (N_31766,N_29894,N_28189);
xor U31767 (N_31767,N_28504,N_28162);
and U31768 (N_31768,N_28362,N_29762);
or U31769 (N_31769,N_28176,N_28725);
nand U31770 (N_31770,N_29597,N_28486);
xnor U31771 (N_31771,N_28338,N_28897);
and U31772 (N_31772,N_28090,N_28677);
nand U31773 (N_31773,N_29323,N_29441);
nand U31774 (N_31774,N_28351,N_28263);
or U31775 (N_31775,N_28565,N_29336);
and U31776 (N_31776,N_29738,N_29354);
xor U31777 (N_31777,N_28220,N_28931);
or U31778 (N_31778,N_28082,N_28920);
and U31779 (N_31779,N_28494,N_29424);
and U31780 (N_31780,N_29118,N_29978);
nor U31781 (N_31781,N_29703,N_29717);
nor U31782 (N_31782,N_28334,N_29222);
nand U31783 (N_31783,N_29698,N_29839);
or U31784 (N_31784,N_29794,N_28227);
xnor U31785 (N_31785,N_29561,N_29104);
or U31786 (N_31786,N_28245,N_28559);
or U31787 (N_31787,N_28441,N_29770);
xnor U31788 (N_31788,N_28770,N_28254);
xnor U31789 (N_31789,N_29156,N_28228);
nand U31790 (N_31790,N_29147,N_29932);
nor U31791 (N_31791,N_29875,N_29518);
xor U31792 (N_31792,N_28214,N_29006);
or U31793 (N_31793,N_28819,N_28026);
xor U31794 (N_31794,N_29347,N_28119);
or U31795 (N_31795,N_29806,N_29543);
nand U31796 (N_31796,N_28357,N_29349);
and U31797 (N_31797,N_28238,N_28960);
and U31798 (N_31798,N_28984,N_29438);
nor U31799 (N_31799,N_29944,N_29352);
xor U31800 (N_31800,N_28916,N_28263);
nor U31801 (N_31801,N_29316,N_29547);
nor U31802 (N_31802,N_29889,N_29780);
xnor U31803 (N_31803,N_29423,N_29748);
and U31804 (N_31804,N_28646,N_29848);
or U31805 (N_31805,N_29290,N_29200);
nor U31806 (N_31806,N_29545,N_29165);
xor U31807 (N_31807,N_28333,N_29301);
and U31808 (N_31808,N_29613,N_28492);
xor U31809 (N_31809,N_28937,N_28999);
or U31810 (N_31810,N_28892,N_29082);
or U31811 (N_31811,N_29980,N_29684);
or U31812 (N_31812,N_29682,N_28275);
nor U31813 (N_31813,N_28165,N_28028);
nand U31814 (N_31814,N_29695,N_29195);
and U31815 (N_31815,N_29210,N_28477);
nand U31816 (N_31816,N_29446,N_29181);
nor U31817 (N_31817,N_28707,N_28561);
nor U31818 (N_31818,N_29135,N_28371);
and U31819 (N_31819,N_28228,N_28026);
and U31820 (N_31820,N_28284,N_28281);
xor U31821 (N_31821,N_28444,N_28995);
nand U31822 (N_31822,N_28305,N_28179);
xor U31823 (N_31823,N_28485,N_29844);
and U31824 (N_31824,N_28684,N_29692);
xor U31825 (N_31825,N_29675,N_29612);
and U31826 (N_31826,N_28554,N_29088);
nor U31827 (N_31827,N_29170,N_29251);
and U31828 (N_31828,N_28514,N_28414);
nand U31829 (N_31829,N_29833,N_29379);
or U31830 (N_31830,N_28916,N_28981);
or U31831 (N_31831,N_28570,N_28921);
and U31832 (N_31832,N_29583,N_28401);
or U31833 (N_31833,N_28707,N_29786);
and U31834 (N_31834,N_29799,N_29790);
nand U31835 (N_31835,N_28902,N_29059);
xor U31836 (N_31836,N_29435,N_28006);
and U31837 (N_31837,N_29364,N_29990);
nand U31838 (N_31838,N_29620,N_29693);
nor U31839 (N_31839,N_28278,N_28175);
xnor U31840 (N_31840,N_29969,N_29545);
and U31841 (N_31841,N_29423,N_29363);
nor U31842 (N_31842,N_28669,N_28191);
or U31843 (N_31843,N_29969,N_28660);
xor U31844 (N_31844,N_28237,N_28191);
xnor U31845 (N_31845,N_28688,N_28712);
xnor U31846 (N_31846,N_29130,N_29869);
nor U31847 (N_31847,N_29806,N_28596);
and U31848 (N_31848,N_28345,N_28948);
nor U31849 (N_31849,N_28744,N_28575);
nand U31850 (N_31850,N_29004,N_29904);
xor U31851 (N_31851,N_28281,N_28675);
nor U31852 (N_31852,N_28769,N_29286);
nor U31853 (N_31853,N_29016,N_29434);
xnor U31854 (N_31854,N_28433,N_29117);
nor U31855 (N_31855,N_28829,N_28692);
and U31856 (N_31856,N_29629,N_28551);
nor U31857 (N_31857,N_29436,N_28715);
and U31858 (N_31858,N_28378,N_28164);
or U31859 (N_31859,N_28225,N_28910);
and U31860 (N_31860,N_28751,N_29247);
nor U31861 (N_31861,N_28806,N_28059);
nor U31862 (N_31862,N_28384,N_29664);
and U31863 (N_31863,N_28253,N_29026);
or U31864 (N_31864,N_28270,N_29063);
nor U31865 (N_31865,N_28732,N_29114);
nand U31866 (N_31866,N_28049,N_29823);
nand U31867 (N_31867,N_28474,N_28491);
nand U31868 (N_31868,N_29270,N_28994);
or U31869 (N_31869,N_29977,N_28337);
and U31870 (N_31870,N_29949,N_28155);
nor U31871 (N_31871,N_29907,N_28801);
nand U31872 (N_31872,N_29322,N_29413);
or U31873 (N_31873,N_29141,N_28806);
xor U31874 (N_31874,N_28268,N_28062);
xnor U31875 (N_31875,N_28114,N_28319);
nor U31876 (N_31876,N_28048,N_28095);
xor U31877 (N_31877,N_29569,N_28901);
nor U31878 (N_31878,N_29031,N_28239);
and U31879 (N_31879,N_29773,N_28487);
nand U31880 (N_31880,N_28716,N_29930);
or U31881 (N_31881,N_29030,N_28504);
nor U31882 (N_31882,N_28655,N_29587);
nand U31883 (N_31883,N_29553,N_28953);
and U31884 (N_31884,N_29868,N_28471);
xor U31885 (N_31885,N_28440,N_29472);
nor U31886 (N_31886,N_29250,N_29345);
nand U31887 (N_31887,N_28242,N_28880);
and U31888 (N_31888,N_29415,N_29463);
nor U31889 (N_31889,N_28332,N_29018);
nand U31890 (N_31890,N_28072,N_28017);
or U31891 (N_31891,N_29908,N_28083);
nand U31892 (N_31892,N_28367,N_29329);
and U31893 (N_31893,N_28559,N_28830);
nor U31894 (N_31894,N_29710,N_28364);
or U31895 (N_31895,N_28796,N_29024);
or U31896 (N_31896,N_29126,N_28807);
nor U31897 (N_31897,N_28796,N_28368);
or U31898 (N_31898,N_28533,N_29535);
nor U31899 (N_31899,N_28536,N_28937);
and U31900 (N_31900,N_29369,N_29405);
nor U31901 (N_31901,N_29570,N_28376);
or U31902 (N_31902,N_29567,N_28452);
nor U31903 (N_31903,N_29408,N_28044);
or U31904 (N_31904,N_29268,N_28051);
and U31905 (N_31905,N_28010,N_28292);
nand U31906 (N_31906,N_28308,N_29456);
or U31907 (N_31907,N_29009,N_29012);
xnor U31908 (N_31908,N_28785,N_29665);
nand U31909 (N_31909,N_29743,N_28050);
and U31910 (N_31910,N_29812,N_29554);
xnor U31911 (N_31911,N_28825,N_29300);
and U31912 (N_31912,N_29590,N_28894);
or U31913 (N_31913,N_29810,N_29003);
xnor U31914 (N_31914,N_29959,N_29435);
nor U31915 (N_31915,N_28910,N_29965);
nand U31916 (N_31916,N_28686,N_29892);
xor U31917 (N_31917,N_29457,N_28026);
or U31918 (N_31918,N_29624,N_28243);
nor U31919 (N_31919,N_29481,N_28189);
xor U31920 (N_31920,N_28534,N_29932);
and U31921 (N_31921,N_28999,N_28115);
or U31922 (N_31922,N_28481,N_29875);
xor U31923 (N_31923,N_29935,N_29474);
nand U31924 (N_31924,N_29018,N_28229);
and U31925 (N_31925,N_29318,N_29820);
xnor U31926 (N_31926,N_28604,N_28878);
and U31927 (N_31927,N_28267,N_29091);
nand U31928 (N_31928,N_29748,N_28355);
nand U31929 (N_31929,N_29349,N_28568);
nor U31930 (N_31930,N_29103,N_28812);
or U31931 (N_31931,N_28980,N_28949);
nand U31932 (N_31932,N_29946,N_29891);
xor U31933 (N_31933,N_28972,N_29609);
and U31934 (N_31934,N_28383,N_29668);
nand U31935 (N_31935,N_29970,N_28969);
nor U31936 (N_31936,N_29141,N_29778);
or U31937 (N_31937,N_29542,N_29142);
nor U31938 (N_31938,N_29648,N_29817);
nor U31939 (N_31939,N_29165,N_29451);
nand U31940 (N_31940,N_29867,N_29620);
xnor U31941 (N_31941,N_28066,N_28393);
nor U31942 (N_31942,N_28372,N_29798);
nand U31943 (N_31943,N_29352,N_29527);
xnor U31944 (N_31944,N_28485,N_28191);
xor U31945 (N_31945,N_29122,N_28962);
or U31946 (N_31946,N_28961,N_28163);
nand U31947 (N_31947,N_29071,N_28940);
nand U31948 (N_31948,N_28650,N_29947);
or U31949 (N_31949,N_29899,N_28884);
and U31950 (N_31950,N_29247,N_28551);
xnor U31951 (N_31951,N_29184,N_28509);
nor U31952 (N_31952,N_28864,N_28774);
or U31953 (N_31953,N_28762,N_29355);
and U31954 (N_31954,N_29824,N_28113);
or U31955 (N_31955,N_28954,N_29633);
nand U31956 (N_31956,N_28916,N_29174);
xnor U31957 (N_31957,N_28846,N_29149);
xor U31958 (N_31958,N_28033,N_29952);
and U31959 (N_31959,N_29222,N_28213);
or U31960 (N_31960,N_28461,N_28955);
nor U31961 (N_31961,N_29475,N_28505);
or U31962 (N_31962,N_28992,N_28781);
xor U31963 (N_31963,N_29035,N_29384);
nor U31964 (N_31964,N_28936,N_28955);
nor U31965 (N_31965,N_28440,N_28808);
nor U31966 (N_31966,N_29112,N_29837);
and U31967 (N_31967,N_29657,N_29526);
or U31968 (N_31968,N_29386,N_28734);
nor U31969 (N_31969,N_29760,N_28956);
and U31970 (N_31970,N_29661,N_29976);
nand U31971 (N_31971,N_28633,N_28881);
and U31972 (N_31972,N_28966,N_29103);
and U31973 (N_31973,N_29701,N_28741);
xor U31974 (N_31974,N_28872,N_28690);
and U31975 (N_31975,N_29708,N_28594);
or U31976 (N_31976,N_29485,N_29503);
nand U31977 (N_31977,N_29923,N_29795);
nand U31978 (N_31978,N_28100,N_29054);
xnor U31979 (N_31979,N_29256,N_28922);
or U31980 (N_31980,N_29270,N_29840);
or U31981 (N_31981,N_29779,N_29817);
nor U31982 (N_31982,N_28477,N_29616);
and U31983 (N_31983,N_28577,N_29399);
xnor U31984 (N_31984,N_28495,N_29370);
xnor U31985 (N_31985,N_29472,N_29509);
nand U31986 (N_31986,N_28695,N_28035);
or U31987 (N_31987,N_28160,N_29374);
xor U31988 (N_31988,N_28806,N_28042);
or U31989 (N_31989,N_29970,N_28843);
xor U31990 (N_31990,N_29080,N_29360);
or U31991 (N_31991,N_28601,N_28592);
and U31992 (N_31992,N_29625,N_28280);
nand U31993 (N_31993,N_28312,N_29196);
and U31994 (N_31994,N_28294,N_29832);
xnor U31995 (N_31995,N_29937,N_29478);
and U31996 (N_31996,N_28856,N_28427);
and U31997 (N_31997,N_29736,N_28729);
xor U31998 (N_31998,N_29807,N_29307);
or U31999 (N_31999,N_28511,N_28934);
and U32000 (N_32000,N_30837,N_30961);
nor U32001 (N_32001,N_31230,N_31654);
or U32002 (N_32002,N_30149,N_31355);
and U32003 (N_32003,N_30241,N_30739);
and U32004 (N_32004,N_31099,N_30221);
xnor U32005 (N_32005,N_30943,N_31544);
nor U32006 (N_32006,N_31970,N_30403);
xor U32007 (N_32007,N_30572,N_30468);
and U32008 (N_32008,N_30482,N_31601);
and U32009 (N_32009,N_31966,N_31824);
and U32010 (N_32010,N_31320,N_30244);
nor U32011 (N_32011,N_30998,N_30225);
xnor U32012 (N_32012,N_30652,N_30278);
and U32013 (N_32013,N_31663,N_30184);
and U32014 (N_32014,N_31042,N_30439);
nand U32015 (N_32015,N_30028,N_30819);
and U32016 (N_32016,N_30722,N_30190);
nor U32017 (N_32017,N_30196,N_30563);
or U32018 (N_32018,N_30307,N_30164);
nand U32019 (N_32019,N_30878,N_31067);
and U32020 (N_32020,N_31033,N_30104);
xnor U32021 (N_32021,N_31222,N_31009);
nand U32022 (N_32022,N_31831,N_30926);
xor U32023 (N_32023,N_30203,N_30651);
or U32024 (N_32024,N_30134,N_30488);
or U32025 (N_32025,N_31828,N_30779);
and U32026 (N_32026,N_31000,N_31946);
or U32027 (N_32027,N_31579,N_31149);
and U32028 (N_32028,N_31707,N_31240);
nor U32029 (N_32029,N_30747,N_31644);
nand U32030 (N_32030,N_30664,N_30816);
nand U32031 (N_32031,N_31167,N_31259);
nand U32032 (N_32032,N_31311,N_31709);
xor U32033 (N_32033,N_31472,N_30323);
nor U32034 (N_32034,N_30511,N_30084);
nor U32035 (N_32035,N_31781,N_31373);
nand U32036 (N_32036,N_30566,N_31914);
or U32037 (N_32037,N_31368,N_31712);
nor U32038 (N_32038,N_30285,N_30896);
or U32039 (N_32039,N_30767,N_31085);
xnor U32040 (N_32040,N_30718,N_30697);
xor U32041 (N_32041,N_30100,N_31789);
xnor U32042 (N_32042,N_31216,N_31779);
or U32043 (N_32043,N_30841,N_31105);
or U32044 (N_32044,N_31389,N_31207);
xnor U32045 (N_32045,N_30354,N_31924);
nand U32046 (N_32046,N_30092,N_30073);
nand U32047 (N_32047,N_30344,N_30796);
xnor U32048 (N_32048,N_31145,N_30161);
xor U32049 (N_32049,N_30736,N_30257);
nor U32050 (N_32050,N_31959,N_31186);
xnor U32051 (N_32051,N_31376,N_30338);
and U32052 (N_32052,N_30729,N_31539);
or U32053 (N_32053,N_30935,N_31742);
xnor U32054 (N_32054,N_31255,N_30625);
nor U32055 (N_32055,N_31528,N_31856);
or U32056 (N_32056,N_30933,N_30724);
and U32057 (N_32057,N_30860,N_31581);
xor U32058 (N_32058,N_30088,N_31490);
nand U32059 (N_32059,N_31518,N_30016);
xor U32060 (N_32060,N_30938,N_31699);
or U32061 (N_32061,N_31181,N_31121);
nand U32062 (N_32062,N_31730,N_31401);
nand U32063 (N_32063,N_30632,N_30982);
xor U32064 (N_32064,N_30151,N_31393);
xnor U32065 (N_32065,N_31281,N_31236);
xor U32066 (N_32066,N_30447,N_30853);
nor U32067 (N_32067,N_30717,N_30352);
and U32068 (N_32068,N_30266,N_30702);
xor U32069 (N_32069,N_31814,N_31512);
xor U32070 (N_32070,N_31697,N_31992);
xnor U32071 (N_32071,N_30059,N_31233);
nor U32072 (N_32072,N_31615,N_31506);
xor U32073 (N_32073,N_31410,N_31143);
xor U32074 (N_32074,N_31865,N_31116);
nand U32075 (N_32075,N_31750,N_31883);
nor U32076 (N_32076,N_31250,N_30519);
and U32077 (N_32077,N_30744,N_30437);
nor U32078 (N_32078,N_30904,N_31030);
nand U32079 (N_32079,N_31107,N_30053);
nor U32080 (N_32080,N_31643,N_30004);
nand U32081 (N_32081,N_31449,N_31426);
or U32082 (N_32082,N_31874,N_31557);
xor U32083 (N_32083,N_31383,N_30765);
xnor U32084 (N_32084,N_30399,N_30347);
nand U32085 (N_32085,N_30044,N_30823);
nand U32086 (N_32086,N_30362,N_31405);
nand U32087 (N_32087,N_30355,N_30592);
or U32088 (N_32088,N_30500,N_31575);
or U32089 (N_32089,N_31523,N_30758);
and U32090 (N_32090,N_30855,N_31330);
nand U32091 (N_32091,N_30994,N_31673);
nand U32092 (N_32092,N_30143,N_31063);
nand U32093 (N_32093,N_31571,N_31602);
xnor U32094 (N_32094,N_31433,N_30971);
xnor U32095 (N_32095,N_31117,N_31827);
xnor U32096 (N_32096,N_30840,N_30996);
xor U32097 (N_32097,N_30430,N_31927);
xor U32098 (N_32098,N_30689,N_30115);
and U32099 (N_32099,N_30547,N_30630);
and U32100 (N_32100,N_30436,N_31911);
and U32101 (N_32101,N_30928,N_30969);
or U32102 (N_32102,N_30615,N_31029);
xor U32103 (N_32103,N_30556,N_31609);
or U32104 (N_32104,N_30041,N_30398);
nor U32105 (N_32105,N_31130,N_30948);
xnor U32106 (N_32106,N_30715,N_31316);
or U32107 (N_32107,N_30679,N_31810);
xor U32108 (N_32108,N_31682,N_31676);
nand U32109 (N_32109,N_30516,N_31944);
or U32110 (N_32110,N_31439,N_30423);
nor U32111 (N_32111,N_30414,N_31982);
and U32112 (N_32112,N_31765,N_30450);
nor U32113 (N_32113,N_31733,N_31066);
or U32114 (N_32114,N_30815,N_30907);
nor U32115 (N_32115,N_31495,N_31479);
xor U32116 (N_32116,N_30030,N_30506);
and U32117 (N_32117,N_31483,N_31890);
nor U32118 (N_32118,N_31237,N_30021);
and U32119 (N_32119,N_30951,N_30497);
or U32120 (N_32120,N_31341,N_30981);
nand U32121 (N_32121,N_31157,N_30181);
nand U32122 (N_32122,N_30007,N_30214);
nor U32123 (N_32123,N_30772,N_31205);
and U32124 (N_32124,N_30438,N_30140);
and U32125 (N_32125,N_30346,N_30018);
nor U32126 (N_32126,N_31525,N_30475);
and U32127 (N_32127,N_31104,N_30496);
and U32128 (N_32128,N_30569,N_30219);
and U32129 (N_32129,N_30080,N_30581);
nand U32130 (N_32130,N_30452,N_30263);
or U32131 (N_32131,N_31200,N_31652);
nor U32132 (N_32132,N_30017,N_31830);
nor U32133 (N_32133,N_30383,N_31511);
and U32134 (N_32134,N_31941,N_30977);
and U32135 (N_32135,N_31262,N_30393);
xnor U32136 (N_32136,N_30834,N_31139);
xor U32137 (N_32137,N_30427,N_31298);
nor U32138 (N_32138,N_30377,N_31432);
nor U32139 (N_32139,N_31731,N_30486);
and U32140 (N_32140,N_30645,N_30340);
or U32141 (N_32141,N_30463,N_31873);
xor U32142 (N_32142,N_30039,N_30609);
xnor U32143 (N_32143,N_31292,N_30696);
xor U32144 (N_32144,N_31429,N_30678);
and U32145 (N_32145,N_31753,N_31168);
and U32146 (N_32146,N_31215,N_30580);
and U32147 (N_32147,N_30617,N_30881);
and U32148 (N_32148,N_30731,N_31952);
nand U32149 (N_32149,N_31701,N_30976);
nand U32150 (N_32150,N_31335,N_31723);
and U32151 (N_32151,N_30210,N_30634);
or U32152 (N_32152,N_30799,N_30946);
xor U32153 (N_32153,N_31166,N_31118);
nor U32154 (N_32154,N_31305,N_31885);
xnor U32155 (N_32155,N_31520,N_30118);
or U32156 (N_32156,N_30136,N_30324);
xor U32157 (N_32157,N_30908,N_30224);
and U32158 (N_32158,N_31835,N_30009);
xor U32159 (N_32159,N_30160,N_30000);
xor U32160 (N_32160,N_30884,N_30903);
nor U32161 (N_32161,N_31208,N_31713);
or U32162 (N_32162,N_30601,N_30342);
xor U32163 (N_32163,N_31268,N_31880);
nand U32164 (N_32164,N_30809,N_31464);
nor U32165 (N_32165,N_30610,N_31582);
nand U32166 (N_32166,N_30428,N_30742);
and U32167 (N_32167,N_31407,N_31070);
xnor U32168 (N_32168,N_30723,N_30813);
or U32169 (N_32169,N_30199,N_31134);
or U32170 (N_32170,N_31092,N_31427);
nor U32171 (N_32171,N_31431,N_30985);
and U32172 (N_32172,N_30892,N_31576);
nor U32173 (N_32173,N_31350,N_31362);
nand U32174 (N_32174,N_30498,N_30591);
or U32175 (N_32175,N_31349,N_30852);
or U32176 (N_32176,N_31651,N_30856);
or U32177 (N_32177,N_31315,N_30562);
nand U32178 (N_32178,N_30783,N_31229);
or U32179 (N_32179,N_31372,N_31308);
and U32180 (N_32180,N_31780,N_31034);
nand U32181 (N_32181,N_31922,N_30924);
nand U32182 (N_32182,N_30068,N_31183);
xor U32183 (N_32183,N_30820,N_30201);
nor U32184 (N_32184,N_30487,N_31761);
and U32185 (N_32185,N_31684,N_30382);
xor U32186 (N_32186,N_30608,N_30267);
xnor U32187 (N_32187,N_30211,N_31562);
and U32188 (N_32188,N_31833,N_31360);
xor U32189 (N_32189,N_31995,N_31073);
nand U32190 (N_32190,N_31172,N_30781);
nor U32191 (N_32191,N_30114,N_31363);
nand U32192 (N_32192,N_30958,N_31419);
xor U32193 (N_32193,N_31715,N_30550);
and U32194 (N_32194,N_30560,N_31955);
nand U32195 (N_32195,N_30991,N_30682);
nor U32196 (N_32196,N_31103,N_30646);
and U32197 (N_32197,N_31743,N_31385);
or U32198 (N_32198,N_30275,N_30405);
nor U32199 (N_32199,N_30390,N_31365);
or U32200 (N_32200,N_30847,N_31267);
nor U32201 (N_32201,N_31832,N_30215);
nor U32202 (N_32202,N_30406,N_31558);
nor U32203 (N_32203,N_30006,N_31132);
nor U32204 (N_32204,N_31272,N_31003);
nor U32205 (N_32205,N_30345,N_30811);
nor U32206 (N_32206,N_31926,N_31792);
nand U32207 (N_32207,N_30013,N_31352);
nor U32208 (N_32208,N_30271,N_31958);
nand U32209 (N_32209,N_31553,N_30002);
and U32210 (N_32210,N_31996,N_31773);
or U32211 (N_32211,N_30337,N_31803);
nor U32212 (N_32212,N_30999,N_30313);
nand U32213 (N_32213,N_31402,N_30228);
nand U32214 (N_32214,N_31155,N_31224);
or U32215 (N_32215,N_31878,N_31194);
or U32216 (N_32216,N_30588,N_30426);
xnor U32217 (N_32217,N_31908,N_31093);
xnor U32218 (N_32218,N_30862,N_30328);
or U32219 (N_32219,N_31800,N_30599);
xnor U32220 (N_32220,N_30795,N_31983);
and U32221 (N_32221,N_31403,N_31095);
nand U32222 (N_32222,N_31189,N_31074);
and U32223 (N_32223,N_30240,N_30824);
nor U32224 (N_32224,N_30208,N_31202);
nor U32225 (N_32225,N_30768,N_30705);
and U32226 (N_32226,N_30070,N_30858);
nand U32227 (N_32227,N_31641,N_31437);
or U32228 (N_32228,N_30404,N_31864);
nor U32229 (N_32229,N_31062,N_31160);
xor U32230 (N_32230,N_30207,N_30621);
or U32231 (N_32231,N_31276,N_30917);
or U32232 (N_32232,N_31319,N_30034);
nor U32233 (N_32233,N_30864,N_30420);
and U32234 (N_32234,N_31120,N_31583);
or U32235 (N_32235,N_30553,N_31109);
nand U32236 (N_32236,N_31968,N_30358);
nor U32237 (N_32237,N_30507,N_31179);
nor U32238 (N_32238,N_31106,N_30415);
and U32239 (N_32239,N_31210,N_31804);
or U32240 (N_32240,N_31621,N_31223);
xor U32241 (N_32241,N_30727,N_31185);
nand U32242 (N_32242,N_31887,N_31416);
xnor U32243 (N_32243,N_31845,N_30670);
and U32244 (N_32244,N_31133,N_31559);
or U32245 (N_32245,N_30655,N_30687);
nor U32246 (N_32246,N_31633,N_31022);
or U32247 (N_32247,N_31717,N_31752);
or U32248 (N_32248,N_30076,N_30578);
nor U32249 (N_32249,N_30083,N_30418);
nor U32250 (N_32250,N_31057,N_30901);
xor U32251 (N_32251,N_31015,N_30356);
nor U32252 (N_32252,N_30410,N_31754);
or U32253 (N_32253,N_31026,N_31053);
nor U32254 (N_32254,N_30746,N_30294);
nand U32255 (N_32255,N_31445,N_31171);
nand U32256 (N_32256,N_31551,N_31076);
xnor U32257 (N_32257,N_30132,N_30960);
nand U32258 (N_32258,N_31078,N_30594);
xor U32259 (N_32259,N_31082,N_31328);
and U32260 (N_32260,N_30010,N_30432);
nor U32261 (N_32261,N_30077,N_30582);
or U32262 (N_32262,N_30019,N_30654);
nand U32263 (N_32263,N_30921,N_31114);
nand U32264 (N_32264,N_30079,N_30321);
nor U32265 (N_32265,N_31014,N_30025);
xnor U32266 (N_32266,N_31290,N_31893);
and U32267 (N_32267,N_31039,N_30798);
or U32268 (N_32268,N_31069,N_31028);
nand U32269 (N_32269,N_30116,N_31212);
xor U32270 (N_32270,N_31517,N_30467);
nor U32271 (N_32271,N_30492,N_30311);
or U32272 (N_32272,N_30698,N_31649);
or U32273 (N_32273,N_30198,N_30336);
or U32274 (N_32274,N_30407,N_31176);
nand U32275 (N_32275,N_31745,N_30431);
nor U32276 (N_32276,N_31550,N_30671);
nor U32277 (N_32277,N_31805,N_31936);
nor U32278 (N_32278,N_30932,N_30886);
nor U32279 (N_32279,N_31678,N_30193);
and U32280 (N_32280,N_30848,N_30005);
or U32281 (N_32281,N_31273,N_31438);
xor U32282 (N_32282,N_31987,N_31219);
xnor U32283 (N_32283,N_31627,N_31313);
and U32284 (N_32284,N_30082,N_31784);
or U32285 (N_32285,N_30966,N_30803);
and U32286 (N_32286,N_31694,N_31796);
nor U32287 (N_32287,N_30561,N_30446);
and U32288 (N_32288,N_30676,N_31879);
or U32289 (N_32289,N_30922,N_30995);
xnor U32290 (N_32290,N_30648,N_31625);
or U32291 (N_32291,N_31096,N_30205);
or U32292 (N_32292,N_30071,N_31954);
and U32293 (N_32293,N_30147,N_30288);
xor U32294 (N_32294,N_31683,N_31404);
xnor U32295 (N_32295,N_31221,N_31767);
nand U32296 (N_32296,N_30916,N_30064);
nor U32297 (N_32297,N_30156,N_30280);
nand U32298 (N_32298,N_30125,N_31881);
xor U32299 (N_32299,N_30883,N_30268);
nand U32300 (N_32300,N_30639,N_31976);
and U32301 (N_32301,N_31882,N_31795);
xnor U32302 (N_32302,N_30636,N_31012);
xnor U32303 (N_32303,N_30032,N_31367);
or U32304 (N_32304,N_31459,N_30704);
nor U32305 (N_32305,N_30052,N_31301);
and U32306 (N_32306,N_31147,N_30669);
or U32307 (N_32307,N_30048,N_31428);
and U32308 (N_32308,N_30135,N_30491);
xnor U32309 (N_32309,N_31953,N_31573);
nand U32310 (N_32310,N_30939,N_30332);
xor U32311 (N_32311,N_30392,N_30379);
nor U32312 (N_32312,N_30272,N_30534);
nand U32313 (N_32313,N_31671,N_31718);
or U32314 (N_32314,N_30528,N_30757);
xnor U32315 (N_32315,N_30229,N_31919);
and U32316 (N_32316,N_31857,N_31923);
nand U32317 (N_32317,N_30433,N_31720);
nor U32318 (N_32318,N_31465,N_31515);
nand U32319 (N_32319,N_30102,N_30289);
nand U32320 (N_32320,N_30627,N_30117);
xnor U32321 (N_32321,N_31333,N_30234);
nor U32322 (N_32322,N_31421,N_31749);
nor U32323 (N_32323,N_30902,N_30416);
and U32324 (N_32324,N_31309,N_30239);
nor U32325 (N_32325,N_31425,N_30973);
and U32326 (N_32326,N_30735,N_31819);
nand U32327 (N_32327,N_30369,N_30490);
or U32328 (N_32328,N_31928,N_30213);
nor U32329 (N_32329,N_30564,N_31868);
xor U32330 (N_32330,N_30168,N_30777);
and U32331 (N_32331,N_31307,N_30863);
nand U32332 (N_32332,N_31261,N_31161);
nor U32333 (N_32333,N_31534,N_31310);
xor U32334 (N_32334,N_31667,N_30179);
nand U32335 (N_32335,N_31605,N_31600);
nand U32336 (N_32336,N_31768,N_30106);
nor U32337 (N_32337,N_31642,N_31038);
nand U32338 (N_32338,N_30359,N_31248);
or U32339 (N_32339,N_31500,N_31314);
nor U32340 (N_32340,N_31794,N_31001);
nor U32341 (N_32341,N_31138,N_30605);
xor U32342 (N_32342,N_31843,N_30111);
or U32343 (N_32343,N_30489,N_30276);
and U32344 (N_32344,N_30633,N_31706);
nor U32345 (N_32345,N_31415,N_31760);
nand U32346 (N_32346,N_30067,N_30691);
or U32347 (N_32347,N_31691,N_30451);
nor U32348 (N_32348,N_30740,N_30058);
xnor U32349 (N_32349,N_31471,N_30297);
and U32350 (N_32350,N_30365,N_30714);
or U32351 (N_32351,N_30218,N_30846);
xnor U32352 (N_32352,N_30061,N_31702);
xor U32353 (N_32353,N_31379,N_31011);
or U32354 (N_32354,N_31005,N_30959);
nand U32355 (N_32355,N_31790,N_30441);
xor U32356 (N_32356,N_30527,N_31646);
and U32357 (N_32357,N_30885,N_31653);
nand U32358 (N_32358,N_31971,N_30770);
nor U32359 (N_32359,N_30069,N_31374);
and U32360 (N_32360,N_30330,N_30022);
or U32361 (N_32361,N_30699,N_30422);
nand U32362 (N_32362,N_31163,N_31888);
nor U32363 (N_32363,N_30372,N_31080);
xnor U32364 (N_32364,N_31182,N_30402);
or U32365 (N_32365,N_30797,N_30435);
nor U32366 (N_32366,N_30968,N_31339);
nor U32367 (N_32367,N_31277,N_31046);
nand U32368 (N_32368,N_31178,N_30137);
nor U32369 (N_32369,N_30529,N_30371);
nand U32370 (N_32370,N_30252,N_31430);
nand U32371 (N_32371,N_31640,N_31925);
nor U32372 (N_32372,N_30096,N_31608);
nand U32373 (N_32373,N_31844,N_30130);
nand U32374 (N_32374,N_30963,N_31806);
xor U32375 (N_32375,N_30949,N_31597);
xor U32376 (N_32376,N_31264,N_31388);
and U32377 (N_32377,N_30308,N_31595);
xor U32378 (N_32378,N_31981,N_30157);
nor U32379 (N_32379,N_31196,N_31962);
xnor U32380 (N_32380,N_31146,N_31808);
xor U32381 (N_32381,N_30003,N_31192);
xor U32382 (N_32382,N_31572,N_30539);
nor U32383 (N_32383,N_30987,N_30301);
and U32384 (N_32384,N_30587,N_31849);
or U32385 (N_32385,N_31209,N_30316);
nor U32386 (N_32386,N_30162,N_30386);
nand U32387 (N_32387,N_31173,N_30373);
or U32388 (N_32388,N_30790,N_30776);
xnor U32389 (N_32389,N_31661,N_30220);
and U32390 (N_32390,N_30827,N_31447);
xnor U32391 (N_32391,N_31351,N_30389);
nand U32392 (N_32392,N_31448,N_30876);
xnor U32393 (N_32393,N_31443,N_31793);
nor U32394 (N_32394,N_31510,N_31293);
nand U32395 (N_32395,N_31990,N_30360);
xnor U32396 (N_32396,N_31637,N_31492);
and U32397 (N_32397,N_30217,N_31984);
nand U32398 (N_32398,N_31809,N_30107);
or U32399 (N_32399,N_31318,N_30265);
xor U32400 (N_32400,N_31817,N_31675);
or U32401 (N_32401,N_31246,N_31541);
xor U32402 (N_32402,N_31774,N_31574);
and U32403 (N_32403,N_30442,N_30882);
nor U32404 (N_32404,N_31050,N_30417);
and U32405 (N_32405,N_30898,N_31917);
nor U32406 (N_32406,N_30997,N_30842);
xnor U32407 (N_32407,N_30826,N_30919);
xor U32408 (N_32408,N_30749,N_30155);
nand U32409 (N_32409,N_31366,N_30230);
nand U32410 (N_32410,N_31131,N_31037);
xnor U32411 (N_32411,N_30760,N_30484);
xor U32412 (N_32412,N_30753,N_31239);
xor U32413 (N_32413,N_30817,N_31782);
xnor U32414 (N_32414,N_31850,N_31253);
nor U32415 (N_32415,N_31934,N_31396);
xnor U32416 (N_32416,N_31662,N_31555);
xor U32417 (N_32417,N_31630,N_30533);
or U32418 (N_32418,N_31418,N_31538);
or U32419 (N_32419,N_30286,N_31587);
and U32420 (N_32420,N_30335,N_30703);
and U32421 (N_32421,N_30094,N_31125);
nor U32422 (N_32422,N_30602,N_30887);
nand U32423 (N_32423,N_31227,N_30557);
or U32424 (N_32424,N_31851,N_31537);
or U32425 (N_32425,N_30818,N_30176);
nand U32426 (N_32426,N_31670,N_31618);
xor U32427 (N_32427,N_30026,N_31054);
nand U32428 (N_32428,N_31741,N_30614);
nor U32429 (N_32429,N_30909,N_31386);
nor U32430 (N_32430,N_31122,N_31631);
nand U32431 (N_32431,N_31493,N_31665);
xor U32432 (N_32432,N_30148,N_31148);
and U32433 (N_32433,N_30401,N_31450);
and U32434 (N_32434,N_31611,N_30859);
nor U32435 (N_32435,N_30603,N_31484);
or U32436 (N_32436,N_30046,N_30967);
xnor U32437 (N_32437,N_31135,N_30895);
nor U32438 (N_32438,N_30711,N_30223);
nor U32439 (N_32439,N_31719,N_31007);
and U32440 (N_32440,N_30145,N_30712);
or U32441 (N_32441,N_31536,N_31929);
and U32442 (N_32442,N_31816,N_30351);
nand U32443 (N_32443,N_30694,N_31863);
and U32444 (N_32444,N_30105,N_31705);
and U32445 (N_32445,N_31610,N_30743);
xor U32446 (N_32446,N_30304,N_31469);
nor U32447 (N_32447,N_31889,N_30101);
nor U32448 (N_32448,N_30327,N_30734);
xnor U32449 (N_32449,N_31629,N_30443);
nor U32450 (N_32450,N_30957,N_31894);
xor U32451 (N_32451,N_30642,N_31972);
nand U32452 (N_32452,N_31762,N_31487);
nor U32453 (N_32453,N_31124,N_30965);
xor U32454 (N_32454,N_30501,N_30253);
nand U32455 (N_32455,N_30644,N_31025);
nor U32456 (N_32456,N_30381,N_31757);
xnor U32457 (N_32457,N_31554,N_31543);
nor U32458 (N_32458,N_30845,N_31547);
nand U32459 (N_32459,N_31306,N_30690);
or U32460 (N_32460,N_30387,N_31692);
nand U32461 (N_32461,N_30063,N_31409);
xor U32462 (N_32462,N_31855,N_30471);
nor U32463 (N_32463,N_31658,N_31902);
nand U32464 (N_32464,N_31280,N_31380);
xor U32465 (N_32465,N_30150,N_30260);
nor U32466 (N_32466,N_30334,N_30085);
nand U32467 (N_32467,N_31271,N_30649);
nand U32468 (N_32468,N_30835,N_30290);
or U32469 (N_32469,N_31823,N_30185);
or U32470 (N_32470,N_30659,N_30095);
xor U32471 (N_32471,N_30015,N_30343);
or U32472 (N_32472,N_30139,N_31847);
nor U32473 (N_32473,N_31771,N_31324);
nand U32474 (N_32474,N_31606,N_30978);
nor U32475 (N_32475,N_31156,N_30400);
or U32476 (N_32476,N_30200,N_31619);
and U32477 (N_32477,N_31100,N_30350);
xnor U32478 (N_32478,N_30169,N_30075);
xnor U32479 (N_32479,N_31140,N_31943);
and U32480 (N_32480,N_31175,N_30624);
nand U32481 (N_32481,N_31939,N_30133);
or U32482 (N_32482,N_31820,N_30412);
nand U32483 (N_32483,N_30322,N_31353);
xor U32484 (N_32484,N_30238,N_31297);
xor U32485 (N_32485,N_31866,N_30586);
nor U32486 (N_32486,N_30178,N_31094);
nor U32487 (N_32487,N_30555,N_31446);
nand U32488 (N_32488,N_31907,N_30091);
or U32489 (N_32489,N_30035,N_30585);
nand U32490 (N_32490,N_30593,N_30906);
xnor U32491 (N_32491,N_30459,N_30889);
and U32492 (N_32492,N_30453,N_31897);
nor U32493 (N_32493,N_30927,N_30040);
xnor U32494 (N_32494,N_30087,N_31993);
and U32495 (N_32495,N_30810,N_31737);
nor U32496 (N_32496,N_31516,N_31617);
nor U32497 (N_32497,N_31875,N_30598);
and U32498 (N_32498,N_30368,N_31337);
nor U32499 (N_32499,N_31291,N_31687);
nand U32500 (N_32500,N_30546,N_30525);
xor U32501 (N_32501,N_30623,N_30510);
and U32502 (N_32502,N_30914,N_30604);
or U32503 (N_32503,N_31681,N_31560);
or U32504 (N_32504,N_31287,N_30250);
and U32505 (N_32505,N_30197,N_30086);
nand U32506 (N_32506,N_30099,N_30024);
nand U32507 (N_32507,N_31532,N_30523);
xnor U32508 (N_32508,N_31785,N_31991);
nand U32509 (N_32509,N_30119,N_31604);
and U32510 (N_32510,N_30540,N_31535);
and U32511 (N_32511,N_30339,N_31499);
or U32512 (N_32512,N_31783,N_30620);
or U32513 (N_32513,N_31180,N_31861);
nand U32514 (N_32514,N_30395,N_31354);
nand U32515 (N_32515,N_30851,N_31312);
or U32516 (N_32516,N_30940,N_31193);
xor U32517 (N_32517,N_30650,N_30880);
and U32518 (N_32518,N_30050,N_30665);
nor U32519 (N_32519,N_31384,N_30923);
nor U32520 (N_32520,N_31399,N_30477);
nor U32521 (N_32521,N_30579,N_30606);
xnor U32522 (N_32522,N_31184,N_31481);
nand U32523 (N_32523,N_30074,N_31527);
nand U32524 (N_32524,N_31839,N_31158);
or U32525 (N_32525,N_31470,N_31657);
nor U32526 (N_32526,N_31542,N_30535);
or U32527 (N_32527,N_30188,N_31325);
nand U32528 (N_32528,N_31279,N_30023);
nand U32529 (N_32529,N_31585,N_31501);
nor U32530 (N_32530,N_31044,N_31296);
xor U32531 (N_32531,N_31975,N_31453);
nor U32532 (N_32532,N_30526,N_31747);
nand U32533 (N_32533,N_30033,N_31278);
xnor U32534 (N_32534,N_30710,N_31829);
nand U32535 (N_32535,N_31390,N_30936);
nor U32536 (N_32536,N_31540,N_31411);
and U32537 (N_32537,N_30993,N_30121);
or U32538 (N_32538,N_31931,N_31978);
xor U32539 (N_32539,N_30725,N_30370);
or U32540 (N_32540,N_30693,N_31381);
xor U32541 (N_32541,N_30066,N_31612);
and U32542 (N_32542,N_30911,N_30988);
or U32543 (N_32543,N_31243,N_30476);
xnor U32544 (N_32544,N_30396,N_31870);
nor U32545 (N_32545,N_30964,N_30584);
or U32546 (N_32546,N_31592,N_30618);
nor U32547 (N_32547,N_30930,N_30170);
nor U32548 (N_32548,N_31825,N_31340);
nor U32549 (N_32549,N_31513,N_30072);
nand U32550 (N_32550,N_30899,N_31440);
and U32551 (N_32551,N_31645,N_31323);
and U32552 (N_32552,N_31732,N_30262);
xor U32553 (N_32553,N_31586,N_31299);
nor U32554 (N_32554,N_31935,N_30411);
xnor U32555 (N_32555,N_31018,N_31801);
and U32556 (N_32556,N_30751,N_30242);
and U32557 (N_32557,N_31151,N_30986);
or U32558 (N_32558,N_31032,N_31589);
nor U32559 (N_32559,N_30172,N_30057);
and U32560 (N_32560,N_31444,N_30264);
or U32561 (N_32561,N_31332,N_30302);
or U32562 (N_32562,N_31150,N_30794);
or U32563 (N_32563,N_30122,N_31549);
nor U32564 (N_32564,N_30774,N_31932);
nand U32565 (N_32565,N_31454,N_30637);
nand U32566 (N_32566,N_31552,N_31077);
xor U32567 (N_32567,N_30246,N_30521);
xor U32568 (N_32568,N_31343,N_30954);
nand U32569 (N_32569,N_30349,N_31436);
nor U32570 (N_32570,N_30232,N_30577);
nor U32571 (N_32571,N_31040,N_30915);
xor U32572 (N_32572,N_30686,N_30950);
and U32573 (N_32573,N_30541,N_30684);
nand U32574 (N_32574,N_31813,N_30681);
or U32575 (N_32575,N_30869,N_31282);
or U32576 (N_32576,N_30189,N_30295);
xnor U32577 (N_32577,N_30098,N_30049);
nor U32578 (N_32578,N_30647,N_30329);
and U32579 (N_32579,N_30173,N_30544);
and U32580 (N_32580,N_31564,N_30695);
or U32581 (N_32581,N_30495,N_31509);
xnor U32582 (N_32582,N_30212,N_31578);
or U32583 (N_32583,N_30270,N_31957);
nand U32584 (N_32584,N_31748,N_30206);
nand U32585 (N_32585,N_30469,N_31327);
or U32586 (N_32586,N_30931,N_30187);
or U32587 (N_32587,N_30261,N_31989);
nor U32588 (N_32588,N_31854,N_30707);
xnor U32589 (N_32589,N_31626,N_30622);
nor U32590 (N_32590,N_31696,N_30713);
nand U32591 (N_32591,N_30912,N_30806);
xor U32592 (N_32592,N_30709,N_30031);
xnor U32593 (N_32593,N_31858,N_30472);
nor U32594 (N_32594,N_30741,N_31580);
nor U32595 (N_32595,N_30833,N_30728);
nand U32596 (N_32596,N_30298,N_30318);
nor U32597 (N_32597,N_31862,N_30112);
or U32598 (N_32598,N_31901,N_30551);
nor U32599 (N_32599,N_30658,N_31685);
xor U32600 (N_32600,N_30191,N_31254);
nand U32601 (N_32601,N_30512,N_31345);
xor U32602 (N_32602,N_31686,N_31004);
and U32603 (N_32603,N_30812,N_30520);
or U32604 (N_32604,N_30631,N_31714);
xnor U32605 (N_32605,N_30192,N_31199);
xnor U32606 (N_32606,N_31659,N_30391);
or U32607 (N_32607,N_30844,N_30661);
nor U32608 (N_32608,N_30755,N_30854);
or U32609 (N_32609,N_31422,N_31169);
or U32610 (N_32610,N_31548,N_30413);
or U32611 (N_32611,N_31905,N_30989);
and U32612 (N_32612,N_31036,N_31394);
or U32613 (N_32613,N_31295,N_31974);
xnor U32614 (N_32614,N_31979,N_31755);
or U32615 (N_32615,N_31999,N_31698);
and U32616 (N_32616,N_31111,N_30165);
or U32617 (N_32617,N_30905,N_30641);
xnor U32618 (N_32618,N_30805,N_31206);
xor U32619 (N_32619,N_31047,N_30748);
nor U32620 (N_32620,N_30237,N_31727);
nor U32621 (N_32621,N_30828,N_30154);
or U32622 (N_32622,N_31244,N_31442);
nor U32623 (N_32623,N_31474,N_30688);
nand U32624 (N_32624,N_31346,N_31256);
or U32625 (N_32625,N_31491,N_31607);
or U32626 (N_32626,N_31251,N_30677);
or U32627 (N_32627,N_31568,N_30804);
xnor U32628 (N_32628,N_31364,N_30182);
nor U32629 (N_32629,N_31203,N_30793);
nor U32630 (N_32630,N_30761,N_31556);
nor U32631 (N_32631,N_31530,N_30675);
and U32632 (N_32632,N_30508,N_31545);
nand U32633 (N_32633,N_31079,N_30269);
nand U32634 (N_32634,N_31406,N_31891);
xnor U32635 (N_32635,N_30062,N_30460);
or U32636 (N_32636,N_31217,N_30517);
nor U32637 (N_32637,N_31916,N_30177);
xnor U32638 (N_32638,N_31638,N_30282);
nand U32639 (N_32639,N_31624,N_31098);
or U32640 (N_32640,N_31956,N_30611);
xor U32641 (N_32641,N_30331,N_30708);
or U32642 (N_32642,N_31258,N_31700);
nand U32643 (N_32643,N_30054,N_31710);
xnor U32644 (N_32644,N_31915,N_30020);
and U32645 (N_32645,N_31846,N_31269);
nor U32646 (N_32646,N_31488,N_31377);
or U32647 (N_32647,N_31660,N_30448);
nand U32648 (N_32648,N_31086,N_30607);
nand U32649 (N_32649,N_31084,N_31918);
or U32650 (N_32650,N_30314,N_30129);
nand U32651 (N_32651,N_31480,N_30385);
nand U32652 (N_32652,N_31336,N_31724);
or U32653 (N_32653,N_30754,N_31744);
xnor U32654 (N_32654,N_30126,N_31049);
nand U32655 (N_32655,N_30281,N_30480);
or U32656 (N_32656,N_31842,N_30445);
nand U32657 (N_32657,N_31997,N_31942);
and U32658 (N_32658,N_31616,N_30638);
or U32659 (N_32659,N_30458,N_31174);
or U32660 (N_32660,N_30788,N_30277);
or U32661 (N_32661,N_30202,N_30008);
nand U32662 (N_32662,N_31188,N_30434);
nand U32663 (N_32663,N_30216,N_30745);
xor U32664 (N_32664,N_30771,N_31284);
nand U32665 (N_32665,N_31119,N_31791);
nand U32666 (N_32666,N_31232,N_31358);
xor U32667 (N_32667,N_31371,N_30733);
nor U32668 (N_32668,N_30065,N_30194);
and U32669 (N_32669,N_31059,N_31728);
xor U32670 (N_32670,N_30320,N_31473);
nand U32671 (N_32671,N_30522,N_30947);
nor U32672 (N_32672,N_30663,N_30424);
and U32673 (N_32673,N_31391,N_30097);
nand U32674 (N_32674,N_31772,N_31461);
or U32675 (N_32675,N_30583,N_31693);
nor U32676 (N_32676,N_31679,N_31906);
and U32677 (N_32677,N_31164,N_31725);
xnor U32678 (N_32678,N_30791,N_31204);
nor U32679 (N_32679,N_30530,N_31263);
nor U32680 (N_32680,N_30367,N_30047);
nand U32681 (N_32681,N_30038,N_30786);
and U32682 (N_32682,N_31563,N_31486);
or U32683 (N_32683,N_30056,N_31220);
and U32684 (N_32684,N_30186,N_30113);
xnor U32685 (N_32685,N_31836,N_30730);
nor U32686 (N_32686,N_30893,N_30952);
or U32687 (N_32687,N_31909,N_31656);
xor U32688 (N_32688,N_30027,N_31266);
nor U32689 (N_32689,N_30333,N_30425);
nand U32690 (N_32690,N_31304,N_31455);
nand U32691 (N_32691,N_31949,N_31920);
nand U32692 (N_32692,N_30700,N_31736);
or U32693 (N_32693,N_30683,N_31485);
nor U32694 (N_32694,N_30303,N_30180);
and U32695 (N_32695,N_30738,N_31758);
nand U32696 (N_32696,N_30051,N_30918);
and U32697 (N_32697,N_31435,N_30158);
or U32698 (N_32698,N_30474,N_31788);
nor U32699 (N_32699,N_31502,N_31588);
xnor U32700 (N_32700,N_30629,N_30766);
or U32701 (N_32701,N_30167,N_30673);
xor U32702 (N_32702,N_31751,N_31020);
nand U32703 (N_32703,N_31321,N_30666);
and U32704 (N_32704,N_31947,N_30756);
or U32705 (N_32705,N_30465,N_31408);
xnor U32706 (N_32706,N_31519,N_30299);
nor U32707 (N_32707,N_31677,N_31289);
or U32708 (N_32708,N_30849,N_31478);
nand U32709 (N_32709,N_31872,N_30287);
nand U32710 (N_32710,N_31721,N_31051);
and U32711 (N_32711,N_31023,N_31998);
nand U32712 (N_32712,N_31570,N_30462);
xnor U32713 (N_32713,N_31061,N_30226);
xnor U32714 (N_32714,N_30929,N_30662);
or U32715 (N_32715,N_30283,N_31060);
xnor U32716 (N_32716,N_30910,N_30894);
and U32717 (N_32717,N_30867,N_30296);
and U32718 (N_32718,N_31596,N_30831);
nor U32719 (N_32719,N_31400,N_30408);
and U32720 (N_32720,N_30478,N_31198);
or U32721 (N_32721,N_30247,N_31294);
xnor U32722 (N_32722,N_31187,N_30502);
or U32723 (N_32723,N_31565,N_30600);
or U32724 (N_32724,N_31505,N_31225);
nor U32725 (N_32725,N_30449,N_30861);
or U32726 (N_32726,N_31211,N_31948);
or U32727 (N_32727,N_31462,N_31822);
and U32728 (N_32728,N_31398,N_30870);
or U32729 (N_32729,N_31622,N_31900);
xor U32730 (N_32730,N_31740,N_30762);
and U32731 (N_32731,N_30175,N_30814);
nand U32732 (N_32732,N_31648,N_31242);
xor U32733 (N_32733,N_30706,N_31144);
nand U32734 (N_32734,N_30254,N_31871);
nand U32735 (N_32735,N_31265,N_31154);
nand U32736 (N_32736,N_31064,N_31722);
nor U32737 (N_32737,N_30536,N_30570);
nand U32738 (N_32738,N_31838,N_31933);
or U32739 (N_32739,N_31594,N_31170);
nand U32740 (N_32740,N_30542,N_31136);
or U32741 (N_32741,N_30868,N_31672);
nor U32742 (N_32742,N_31489,N_31821);
nand U32743 (N_32743,N_31359,N_30920);
or U32744 (N_32744,N_31746,N_31655);
nor U32745 (N_32745,N_30720,N_31964);
xnor U32746 (N_32746,N_30504,N_31218);
xnor U32747 (N_32747,N_30789,N_31356);
and U32748 (N_32748,N_31065,N_30612);
nand U32749 (N_32749,N_31620,N_30306);
xnor U32750 (N_32750,N_31071,N_30975);
nand U32751 (N_32751,N_31113,N_31397);
or U32752 (N_32752,N_30291,N_30759);
or U32753 (N_32753,N_30235,N_30956);
and U32754 (N_32754,N_31238,N_30955);
nor U32755 (N_32755,N_31370,N_30726);
or U32756 (N_32756,N_31241,N_31628);
nor U32757 (N_32757,N_30888,N_31815);
nand U32758 (N_32758,N_31392,N_30310);
nor U32759 (N_32759,N_31766,N_31708);
and U32760 (N_32760,N_30376,N_31898);
nor U32761 (N_32761,N_31650,N_30236);
nand U32762 (N_32762,N_30055,N_30875);
or U32763 (N_32763,N_31876,N_31834);
xor U32764 (N_32764,N_30925,N_31159);
or U32765 (N_32765,N_30752,N_31818);
and U32766 (N_32766,N_30384,N_31853);
and U32767 (N_32767,N_31496,N_30801);
nand U32768 (N_32768,N_30380,N_31288);
xnor U32769 (N_32769,N_31162,N_31912);
and U32770 (N_32770,N_30515,N_30357);
xnor U32771 (N_32771,N_31807,N_30983);
and U32772 (N_32772,N_31734,N_30227);
or U32773 (N_32773,N_30248,N_31674);
nor U32774 (N_32774,N_31689,N_31841);
nor U32775 (N_32775,N_31504,N_31778);
xor U32776 (N_32776,N_30596,N_30081);
and U32777 (N_32777,N_31460,N_30305);
nor U32778 (N_32778,N_31075,N_31577);
or U32779 (N_32779,N_31056,N_31300);
nor U32780 (N_32780,N_31195,N_30573);
and U32781 (N_32781,N_31331,N_30716);
or U32782 (N_32782,N_30361,N_31434);
xnor U32783 (N_32783,N_30171,N_30839);
xnor U32784 (N_32784,N_30374,N_30764);
or U32785 (N_32785,N_31895,N_30732);
nand U32786 (N_32786,N_31497,N_30378);
nand U32787 (N_32787,N_31190,N_31521);
xor U32788 (N_32788,N_31546,N_31177);
nor U32789 (N_32789,N_31382,N_30792);
xnor U32790 (N_32790,N_31735,N_31561);
and U32791 (N_32791,N_30364,N_31635);
and U32792 (N_32792,N_30037,N_30479);
nand U32793 (N_32793,N_31058,N_30866);
xor U32794 (N_32794,N_30874,N_31191);
xor U32795 (N_32795,N_31048,N_31378);
xor U32796 (N_32796,N_31087,N_30574);
nand U32797 (N_32797,N_30980,N_31127);
and U32798 (N_32798,N_30685,N_30865);
or U32799 (N_32799,N_30552,N_30292);
or U32800 (N_32800,N_30249,N_30787);
and U32801 (N_32801,N_30456,N_30123);
or U32802 (N_32802,N_31967,N_30499);
and U32803 (N_32803,N_31387,N_30127);
or U32804 (N_32804,N_31896,N_31463);
nor U32805 (N_32805,N_30972,N_30877);
and U32806 (N_32806,N_30773,N_31859);
nand U32807 (N_32807,N_31458,N_30667);
or U32808 (N_32808,N_31357,N_31013);
nand U32809 (N_32809,N_31342,N_30209);
xor U32810 (N_32810,N_31704,N_30174);
nand U32811 (N_32811,N_31102,N_31326);
or U32812 (N_32812,N_31214,N_30485);
or U32813 (N_32813,N_30589,N_30195);
or U32814 (N_32814,N_30944,N_31787);
nor U32815 (N_32815,N_31286,N_31375);
nor U32816 (N_32816,N_30871,N_30255);
xor U32817 (N_32817,N_31249,N_30273);
xnor U32818 (N_32818,N_30913,N_31973);
xnor U32819 (N_32819,N_31089,N_30619);
nor U32820 (N_32820,N_31599,N_31945);
nor U32821 (N_32821,N_30554,N_30873);
nor U32822 (N_32822,N_31475,N_31413);
or U32823 (N_32823,N_31980,N_30110);
nor U32824 (N_32824,N_31777,N_30464);
xor U32825 (N_32825,N_30293,N_30466);
and U32826 (N_32826,N_31252,N_31769);
xnor U32827 (N_32827,N_30737,N_31668);
xnor U32828 (N_32828,N_30348,N_31569);
or U32829 (N_32829,N_30131,N_31088);
and U32830 (N_32830,N_31508,N_30397);
and U32831 (N_32831,N_30233,N_30159);
and U32832 (N_32832,N_30829,N_31503);
xnor U32833 (N_32833,N_30183,N_30470);
xor U32834 (N_32834,N_31852,N_30613);
or U32835 (N_32835,N_30782,N_31529);
xnor U32836 (N_32836,N_30421,N_31634);
xnor U32837 (N_32837,N_31008,N_31016);
and U32838 (N_32838,N_30808,N_31903);
and U32839 (N_32839,N_30120,N_30830);
and U32840 (N_32840,N_31153,N_30979);
xnor U32841 (N_32841,N_31798,N_30984);
nor U32842 (N_32842,N_30481,N_31950);
nand U32843 (N_32843,N_30891,N_31664);
nand U32844 (N_32844,N_30653,N_31201);
xor U32845 (N_32845,N_31763,N_31128);
nand U32846 (N_32846,N_31348,N_31123);
nor U32847 (N_32847,N_31115,N_30942);
or U32848 (N_32848,N_30409,N_31786);
nand U32849 (N_32849,N_31904,N_30388);
xor U32850 (N_32850,N_31197,N_30656);
xnor U32851 (N_32851,N_30353,N_31303);
nand U32852 (N_32852,N_30493,N_31613);
xnor U32853 (N_32853,N_31270,N_31593);
or U32854 (N_32854,N_30309,N_31598);
nand U32855 (N_32855,N_30128,N_30900);
or U32856 (N_32856,N_31826,N_30256);
nand U32857 (N_32857,N_31302,N_31142);
nor U32858 (N_32858,N_30152,N_30545);
xor U32859 (N_32859,N_31245,N_31591);
xnor U32860 (N_32860,N_30974,N_31027);
or U32861 (N_32861,N_31877,N_31021);
xnor U32862 (N_32862,N_30775,N_30518);
or U32863 (N_32863,N_31963,N_31412);
and U32864 (N_32864,N_31068,N_30597);
nand U32865 (N_32865,N_30036,N_31322);
nand U32866 (N_32866,N_31680,N_31647);
nand U32867 (N_32867,N_31985,N_30802);
nand U32868 (N_32868,N_30537,N_31960);
nand U32869 (N_32869,N_31275,N_30643);
and U32870 (N_32870,N_30163,N_31797);
nor U32871 (N_32871,N_30146,N_30457);
xor U32872 (N_32872,N_31776,N_30836);
nand U32873 (N_32873,N_30440,N_31729);
nor U32874 (N_32874,N_30668,N_31417);
nand U32875 (N_32875,N_30012,N_30990);
nand U32876 (N_32876,N_31414,N_31526);
nor U32877 (N_32877,N_31072,N_31522);
nand U32878 (N_32878,N_30549,N_31494);
xnor U32879 (N_32879,N_31055,N_30785);
nor U32880 (N_32880,N_30274,N_31477);
nor U32881 (N_32881,N_30640,N_30635);
and U32882 (N_32882,N_30721,N_30559);
nor U32883 (N_32883,N_30872,N_31590);
nand U32884 (N_32884,N_31913,N_31467);
nand U32885 (N_32885,N_30576,N_30970);
nand U32886 (N_32886,N_30454,N_31108);
xnor U32887 (N_32887,N_31126,N_31456);
nand U32888 (N_32888,N_31006,N_31759);
and U32889 (N_32889,N_31031,N_30701);
nor U32890 (N_32890,N_30692,N_30807);
nand U32891 (N_32891,N_31476,N_30750);
nor U32892 (N_32892,N_31869,N_30800);
nor U32893 (N_32893,N_30153,N_30503);
xnor U32894 (N_32894,N_31584,N_31112);
and U32895 (N_32895,N_30674,N_30138);
nor U32896 (N_32896,N_30455,N_30483);
xor U32897 (N_32897,N_31152,N_30548);
nand U32898 (N_32898,N_31884,N_31165);
xnor U32899 (N_32899,N_30719,N_30444);
xor U32900 (N_32900,N_30251,N_31334);
and U32901 (N_32901,N_31614,N_30419);
or U32902 (N_32902,N_31260,N_30962);
and U32903 (N_32903,N_31756,N_31002);
xnor U32904 (N_32904,N_31091,N_31938);
or U32905 (N_32905,N_30680,N_31110);
nand U32906 (N_32906,N_30222,N_30822);
xor U32907 (N_32907,N_31423,N_30312);
or U32908 (N_32908,N_31468,N_30259);
nand U32909 (N_32909,N_30934,N_31961);
xor U32910 (N_32910,N_31860,N_31669);
or U32911 (N_32911,N_30341,N_30279);
or U32912 (N_32912,N_31101,N_30937);
or U32913 (N_32913,N_31988,N_30363);
nor U32914 (N_32914,N_30575,N_30657);
nand U32915 (N_32915,N_31566,N_31690);
and U32916 (N_32916,N_30144,N_30590);
and U32917 (N_32917,N_30109,N_30103);
nand U32918 (N_32918,N_31567,N_30494);
or U32919 (N_32919,N_30616,N_30300);
and U32920 (N_32920,N_30850,N_31052);
or U32921 (N_32921,N_31329,N_30992);
xor U32922 (N_32922,N_30093,N_31231);
nand U32923 (N_32923,N_30821,N_30325);
xnor U32924 (N_32924,N_31636,N_30780);
xnor U32925 (N_32925,N_31344,N_31899);
nor U32926 (N_32926,N_31274,N_30258);
xnor U32927 (N_32927,N_31081,N_31812);
or U32928 (N_32928,N_31977,N_31369);
xnor U32929 (N_32929,N_31498,N_30558);
nand U32930 (N_32930,N_30042,N_31285);
and U32931 (N_32931,N_31017,N_31361);
xor U32932 (N_32932,N_31951,N_30531);
and U32933 (N_32933,N_30945,N_30825);
xor U32934 (N_32934,N_31043,N_31524);
nor U32935 (N_32935,N_30078,N_30166);
xnor U32936 (N_32936,N_31688,N_31711);
nand U32937 (N_32937,N_31507,N_30543);
xor U32938 (N_32938,N_30953,N_30628);
and U32939 (N_32939,N_31848,N_30660);
nor U32940 (N_32940,N_30843,N_30513);
and U32941 (N_32941,N_31799,N_31910);
xor U32942 (N_32942,N_30090,N_30626);
nand U32943 (N_32943,N_30763,N_31639);
or U32944 (N_32944,N_31228,N_30568);
xnor U32945 (N_32945,N_31141,N_30366);
nand U32946 (N_32946,N_30532,N_31247);
or U32947 (N_32947,N_30284,N_31937);
or U32948 (N_32948,N_31041,N_30778);
nand U32949 (N_32949,N_31466,N_30672);
and U32950 (N_32950,N_31994,N_31531);
and U32951 (N_32951,N_31482,N_30897);
nor U32952 (N_32952,N_31097,N_31969);
and U32953 (N_32953,N_31514,N_31347);
or U32954 (N_32954,N_31317,N_30941);
or U32955 (N_32955,N_30429,N_30784);
xnor U32956 (N_32956,N_31235,N_31739);
nand U32957 (N_32957,N_30514,N_31867);
nand U32958 (N_32958,N_30089,N_30571);
or U32959 (N_32959,N_31010,N_30204);
or U32960 (N_32960,N_30565,N_31338);
nor U32961 (N_32961,N_30319,N_30243);
xor U32962 (N_32962,N_30014,N_30315);
or U32963 (N_32963,N_31886,N_30879);
xor U32964 (N_32964,N_30108,N_30231);
nor U32965 (N_32965,N_30567,N_31965);
xnor U32966 (N_32966,N_30245,N_31811);
nand U32967 (N_32967,N_30524,N_31424);
nor U32968 (N_32968,N_30838,N_30326);
xor U32969 (N_32969,N_31703,N_31726);
nand U32970 (N_32970,N_31921,N_30029);
nor U32971 (N_32971,N_30001,N_31213);
nand U32972 (N_32972,N_30045,N_30538);
and U32973 (N_32973,N_31035,N_31045);
nand U32974 (N_32974,N_31226,N_31234);
nor U32975 (N_32975,N_30141,N_30769);
nand U32976 (N_32976,N_30375,N_30857);
nor U32977 (N_32977,N_31623,N_31137);
nand U32978 (N_32978,N_31603,N_30394);
xnor U32979 (N_32979,N_31775,N_31019);
and U32980 (N_32980,N_31840,N_31764);
nor U32981 (N_32981,N_31632,N_31802);
or U32982 (N_32982,N_31695,N_31940);
nand U32983 (N_32983,N_31441,N_31738);
nand U32984 (N_32984,N_30509,N_31083);
and U32985 (N_32985,N_31129,N_31024);
nand U32986 (N_32986,N_30473,N_30011);
and U32987 (N_32987,N_30595,N_30043);
nor U32988 (N_32988,N_30505,N_31930);
and U32989 (N_32989,N_30317,N_30142);
nand U32990 (N_32990,N_31452,N_30461);
nand U32991 (N_32991,N_31533,N_31420);
nor U32992 (N_32992,N_31090,N_31986);
nor U32993 (N_32993,N_31770,N_31451);
nor U32994 (N_32994,N_31457,N_30060);
nor U32995 (N_32995,N_30124,N_31257);
nor U32996 (N_32996,N_31283,N_31837);
or U32997 (N_32997,N_30832,N_31892);
nand U32998 (N_32998,N_30890,N_31716);
nor U32999 (N_32999,N_31395,N_31666);
and U33000 (N_33000,N_31282,N_30750);
and U33001 (N_33001,N_30075,N_31262);
nor U33002 (N_33002,N_31724,N_30774);
nor U33003 (N_33003,N_30757,N_31065);
xor U33004 (N_33004,N_30530,N_31426);
nand U33005 (N_33005,N_30445,N_31385);
or U33006 (N_33006,N_30664,N_30986);
xor U33007 (N_33007,N_30999,N_31392);
nor U33008 (N_33008,N_30376,N_30521);
nand U33009 (N_33009,N_31802,N_30136);
nor U33010 (N_33010,N_31663,N_30370);
nand U33011 (N_33011,N_30120,N_31581);
nand U33012 (N_33012,N_30170,N_31462);
or U33013 (N_33013,N_30246,N_31825);
and U33014 (N_33014,N_31855,N_30104);
nor U33015 (N_33015,N_30419,N_30397);
or U33016 (N_33016,N_31552,N_30959);
xnor U33017 (N_33017,N_30913,N_31049);
and U33018 (N_33018,N_30121,N_31507);
or U33019 (N_33019,N_31413,N_30846);
and U33020 (N_33020,N_30144,N_30654);
xor U33021 (N_33021,N_31113,N_31413);
or U33022 (N_33022,N_31744,N_31453);
xor U33023 (N_33023,N_31295,N_31733);
nor U33024 (N_33024,N_30643,N_31574);
or U33025 (N_33025,N_30149,N_31213);
xor U33026 (N_33026,N_31696,N_30869);
and U33027 (N_33027,N_31085,N_31230);
nand U33028 (N_33028,N_31715,N_31084);
nand U33029 (N_33029,N_30352,N_30004);
or U33030 (N_33030,N_30162,N_31705);
nand U33031 (N_33031,N_30068,N_30658);
xnor U33032 (N_33032,N_31084,N_31640);
nand U33033 (N_33033,N_31752,N_31091);
or U33034 (N_33034,N_30594,N_31102);
and U33035 (N_33035,N_31527,N_30178);
nand U33036 (N_33036,N_31162,N_30013);
nor U33037 (N_33037,N_30446,N_31318);
nand U33038 (N_33038,N_30031,N_31739);
nand U33039 (N_33039,N_30827,N_30977);
xor U33040 (N_33040,N_31053,N_31066);
and U33041 (N_33041,N_30060,N_31070);
or U33042 (N_33042,N_31373,N_31385);
nor U33043 (N_33043,N_31687,N_31171);
nor U33044 (N_33044,N_31312,N_30045);
and U33045 (N_33045,N_30282,N_31498);
nor U33046 (N_33046,N_31137,N_30281);
or U33047 (N_33047,N_31898,N_30156);
or U33048 (N_33048,N_31850,N_30577);
nor U33049 (N_33049,N_30937,N_31561);
and U33050 (N_33050,N_30122,N_30402);
nor U33051 (N_33051,N_31410,N_31757);
nor U33052 (N_33052,N_30663,N_30645);
and U33053 (N_33053,N_30842,N_30836);
or U33054 (N_33054,N_30368,N_31751);
xor U33055 (N_33055,N_31421,N_31878);
nor U33056 (N_33056,N_31817,N_31400);
nor U33057 (N_33057,N_31870,N_31950);
nand U33058 (N_33058,N_31316,N_31414);
or U33059 (N_33059,N_30342,N_30285);
nor U33060 (N_33060,N_31397,N_31423);
xor U33061 (N_33061,N_31989,N_31791);
xnor U33062 (N_33062,N_31584,N_31005);
nor U33063 (N_33063,N_31340,N_30811);
xnor U33064 (N_33064,N_30038,N_31728);
nor U33065 (N_33065,N_30571,N_30527);
nor U33066 (N_33066,N_30686,N_30389);
and U33067 (N_33067,N_30449,N_31268);
nand U33068 (N_33068,N_31454,N_30365);
or U33069 (N_33069,N_31197,N_30178);
nor U33070 (N_33070,N_30025,N_31600);
xor U33071 (N_33071,N_31548,N_31306);
nand U33072 (N_33072,N_30845,N_31008);
and U33073 (N_33073,N_30821,N_30083);
nor U33074 (N_33074,N_31802,N_30053);
and U33075 (N_33075,N_31195,N_31395);
and U33076 (N_33076,N_31318,N_30734);
nor U33077 (N_33077,N_31293,N_31752);
xnor U33078 (N_33078,N_30323,N_30354);
nand U33079 (N_33079,N_30683,N_31793);
xnor U33080 (N_33080,N_31043,N_31911);
or U33081 (N_33081,N_30303,N_31329);
and U33082 (N_33082,N_30630,N_31551);
or U33083 (N_33083,N_30989,N_31516);
and U33084 (N_33084,N_30454,N_31311);
nor U33085 (N_33085,N_31743,N_30378);
nor U33086 (N_33086,N_30547,N_31592);
xnor U33087 (N_33087,N_30041,N_30884);
and U33088 (N_33088,N_31896,N_30002);
nand U33089 (N_33089,N_31314,N_31055);
xor U33090 (N_33090,N_30324,N_30424);
nand U33091 (N_33091,N_30893,N_30201);
xor U33092 (N_33092,N_30585,N_31806);
and U33093 (N_33093,N_31498,N_31591);
or U33094 (N_33094,N_30505,N_30794);
and U33095 (N_33095,N_30369,N_31642);
xnor U33096 (N_33096,N_30698,N_31000);
xor U33097 (N_33097,N_31001,N_30401);
xor U33098 (N_33098,N_30236,N_30628);
or U33099 (N_33099,N_30998,N_30729);
nand U33100 (N_33100,N_30181,N_30643);
and U33101 (N_33101,N_31749,N_31394);
xnor U33102 (N_33102,N_31625,N_30160);
and U33103 (N_33103,N_30665,N_31882);
nand U33104 (N_33104,N_30727,N_30551);
nand U33105 (N_33105,N_30740,N_31142);
nand U33106 (N_33106,N_30332,N_31931);
nor U33107 (N_33107,N_30385,N_30520);
nand U33108 (N_33108,N_30211,N_31018);
and U33109 (N_33109,N_30792,N_30670);
xor U33110 (N_33110,N_30490,N_31921);
xor U33111 (N_33111,N_30003,N_30378);
nand U33112 (N_33112,N_30272,N_31455);
or U33113 (N_33113,N_30661,N_30012);
nand U33114 (N_33114,N_31881,N_30482);
nand U33115 (N_33115,N_31790,N_31302);
nor U33116 (N_33116,N_31986,N_31475);
xnor U33117 (N_33117,N_30052,N_31880);
or U33118 (N_33118,N_30271,N_30495);
xor U33119 (N_33119,N_31222,N_30854);
nor U33120 (N_33120,N_30109,N_31509);
or U33121 (N_33121,N_30765,N_31102);
or U33122 (N_33122,N_30067,N_30657);
nor U33123 (N_33123,N_30682,N_31709);
xor U33124 (N_33124,N_30595,N_31852);
or U33125 (N_33125,N_30399,N_31831);
xnor U33126 (N_33126,N_30336,N_30252);
nor U33127 (N_33127,N_31712,N_31260);
xor U33128 (N_33128,N_30260,N_31330);
xor U33129 (N_33129,N_31280,N_31477);
and U33130 (N_33130,N_30213,N_30313);
and U33131 (N_33131,N_30135,N_30199);
nor U33132 (N_33132,N_31524,N_31087);
nand U33133 (N_33133,N_30008,N_31000);
and U33134 (N_33134,N_31763,N_30704);
nor U33135 (N_33135,N_31228,N_30182);
and U33136 (N_33136,N_30941,N_30226);
or U33137 (N_33137,N_31558,N_31956);
nor U33138 (N_33138,N_30466,N_30029);
nand U33139 (N_33139,N_31012,N_30490);
and U33140 (N_33140,N_30451,N_30912);
and U33141 (N_33141,N_30382,N_30916);
nor U33142 (N_33142,N_31403,N_31539);
nor U33143 (N_33143,N_31571,N_31163);
and U33144 (N_33144,N_30348,N_31418);
and U33145 (N_33145,N_30372,N_31949);
nand U33146 (N_33146,N_31828,N_30706);
nor U33147 (N_33147,N_30603,N_31288);
or U33148 (N_33148,N_30759,N_30638);
nor U33149 (N_33149,N_31929,N_31223);
and U33150 (N_33150,N_31574,N_31827);
nand U33151 (N_33151,N_30910,N_30995);
and U33152 (N_33152,N_31947,N_30115);
xor U33153 (N_33153,N_31173,N_30267);
nor U33154 (N_33154,N_30285,N_30663);
nor U33155 (N_33155,N_31086,N_31993);
nand U33156 (N_33156,N_31476,N_31484);
xnor U33157 (N_33157,N_31776,N_31366);
nand U33158 (N_33158,N_31569,N_30437);
or U33159 (N_33159,N_30781,N_30961);
xnor U33160 (N_33160,N_31660,N_30571);
nor U33161 (N_33161,N_31305,N_30718);
and U33162 (N_33162,N_31891,N_30311);
or U33163 (N_33163,N_31914,N_30234);
xor U33164 (N_33164,N_30413,N_30505);
or U33165 (N_33165,N_31837,N_31674);
and U33166 (N_33166,N_30286,N_30574);
or U33167 (N_33167,N_31255,N_31971);
or U33168 (N_33168,N_30779,N_31590);
and U33169 (N_33169,N_30916,N_31785);
nor U33170 (N_33170,N_31837,N_31415);
and U33171 (N_33171,N_31886,N_31315);
nor U33172 (N_33172,N_30202,N_31787);
nand U33173 (N_33173,N_30633,N_30376);
or U33174 (N_33174,N_30040,N_31183);
nor U33175 (N_33175,N_30414,N_30108);
xor U33176 (N_33176,N_31123,N_31224);
and U33177 (N_33177,N_30444,N_31440);
and U33178 (N_33178,N_30879,N_31132);
and U33179 (N_33179,N_31879,N_30860);
and U33180 (N_33180,N_31743,N_31383);
nand U33181 (N_33181,N_31558,N_31988);
nor U33182 (N_33182,N_30727,N_30499);
and U33183 (N_33183,N_30243,N_30218);
xnor U33184 (N_33184,N_31214,N_30512);
and U33185 (N_33185,N_30186,N_31698);
nand U33186 (N_33186,N_31857,N_31841);
xor U33187 (N_33187,N_31028,N_31245);
and U33188 (N_33188,N_30489,N_31820);
and U33189 (N_33189,N_30912,N_30151);
or U33190 (N_33190,N_31238,N_31029);
nand U33191 (N_33191,N_30426,N_31304);
and U33192 (N_33192,N_31940,N_30374);
or U33193 (N_33193,N_31330,N_31717);
and U33194 (N_33194,N_30204,N_31214);
or U33195 (N_33195,N_30993,N_31639);
xor U33196 (N_33196,N_31720,N_30605);
nor U33197 (N_33197,N_31805,N_30894);
nor U33198 (N_33198,N_30108,N_30627);
nor U33199 (N_33199,N_31686,N_30242);
xnor U33200 (N_33200,N_30416,N_30615);
or U33201 (N_33201,N_30283,N_31457);
or U33202 (N_33202,N_30964,N_31120);
and U33203 (N_33203,N_31267,N_31500);
xnor U33204 (N_33204,N_31503,N_30337);
nor U33205 (N_33205,N_31468,N_31913);
or U33206 (N_33206,N_31646,N_31668);
nor U33207 (N_33207,N_30025,N_31229);
or U33208 (N_33208,N_30258,N_31918);
and U33209 (N_33209,N_30187,N_30292);
nor U33210 (N_33210,N_30962,N_30250);
or U33211 (N_33211,N_30460,N_30227);
nand U33212 (N_33212,N_31670,N_30359);
nand U33213 (N_33213,N_31003,N_30798);
nand U33214 (N_33214,N_30250,N_31698);
and U33215 (N_33215,N_30671,N_30992);
nor U33216 (N_33216,N_30016,N_31770);
xor U33217 (N_33217,N_30292,N_30548);
nand U33218 (N_33218,N_31960,N_31477);
or U33219 (N_33219,N_31589,N_31904);
xor U33220 (N_33220,N_30108,N_31952);
or U33221 (N_33221,N_31020,N_31976);
nor U33222 (N_33222,N_30292,N_30099);
and U33223 (N_33223,N_31774,N_31470);
nand U33224 (N_33224,N_31986,N_30561);
or U33225 (N_33225,N_30866,N_31751);
nor U33226 (N_33226,N_30920,N_30522);
and U33227 (N_33227,N_31122,N_30082);
xor U33228 (N_33228,N_30455,N_31753);
nand U33229 (N_33229,N_30666,N_31029);
nor U33230 (N_33230,N_30774,N_30944);
nand U33231 (N_33231,N_30874,N_31271);
and U33232 (N_33232,N_30536,N_31162);
and U33233 (N_33233,N_30902,N_30825);
nand U33234 (N_33234,N_30670,N_31330);
and U33235 (N_33235,N_30422,N_31412);
or U33236 (N_33236,N_31053,N_31465);
nor U33237 (N_33237,N_31000,N_30763);
or U33238 (N_33238,N_31869,N_31235);
xnor U33239 (N_33239,N_30473,N_30637);
xor U33240 (N_33240,N_31579,N_30278);
and U33241 (N_33241,N_31234,N_31468);
and U33242 (N_33242,N_30013,N_30749);
and U33243 (N_33243,N_30846,N_30075);
and U33244 (N_33244,N_31503,N_30314);
and U33245 (N_33245,N_31993,N_30443);
xnor U33246 (N_33246,N_31178,N_31459);
and U33247 (N_33247,N_31356,N_31116);
nand U33248 (N_33248,N_30777,N_30417);
and U33249 (N_33249,N_30209,N_30487);
nand U33250 (N_33250,N_31609,N_30927);
or U33251 (N_33251,N_30860,N_31916);
or U33252 (N_33252,N_30088,N_30454);
or U33253 (N_33253,N_31493,N_31295);
xor U33254 (N_33254,N_31787,N_31640);
nor U33255 (N_33255,N_30033,N_30872);
or U33256 (N_33256,N_31145,N_30626);
nand U33257 (N_33257,N_31728,N_31840);
nand U33258 (N_33258,N_30308,N_31693);
xnor U33259 (N_33259,N_31124,N_31530);
nor U33260 (N_33260,N_30873,N_30075);
xnor U33261 (N_33261,N_31667,N_30533);
nand U33262 (N_33262,N_30751,N_31344);
nand U33263 (N_33263,N_30497,N_31400);
xor U33264 (N_33264,N_30987,N_31420);
or U33265 (N_33265,N_31781,N_30597);
or U33266 (N_33266,N_31672,N_30052);
nor U33267 (N_33267,N_31996,N_31906);
xnor U33268 (N_33268,N_31867,N_31488);
nor U33269 (N_33269,N_30577,N_30670);
xor U33270 (N_33270,N_30443,N_30868);
xnor U33271 (N_33271,N_30532,N_31264);
nand U33272 (N_33272,N_30078,N_30132);
nand U33273 (N_33273,N_30117,N_31670);
and U33274 (N_33274,N_31471,N_30981);
or U33275 (N_33275,N_30175,N_31847);
nand U33276 (N_33276,N_31978,N_31958);
xor U33277 (N_33277,N_30970,N_30967);
and U33278 (N_33278,N_30772,N_31013);
or U33279 (N_33279,N_30115,N_31405);
nand U33280 (N_33280,N_31646,N_31969);
or U33281 (N_33281,N_30583,N_31636);
or U33282 (N_33282,N_30764,N_31764);
or U33283 (N_33283,N_30779,N_31345);
xor U33284 (N_33284,N_31027,N_30032);
or U33285 (N_33285,N_30898,N_31689);
and U33286 (N_33286,N_31012,N_31258);
nor U33287 (N_33287,N_31788,N_31054);
nor U33288 (N_33288,N_31318,N_30979);
and U33289 (N_33289,N_31874,N_31829);
xnor U33290 (N_33290,N_30889,N_30042);
nor U33291 (N_33291,N_30560,N_31946);
and U33292 (N_33292,N_31087,N_31907);
or U33293 (N_33293,N_30920,N_31629);
nor U33294 (N_33294,N_31130,N_31477);
nor U33295 (N_33295,N_30229,N_30941);
or U33296 (N_33296,N_30926,N_31555);
and U33297 (N_33297,N_30134,N_31917);
xnor U33298 (N_33298,N_30426,N_31546);
xnor U33299 (N_33299,N_31931,N_30854);
nand U33300 (N_33300,N_31806,N_31666);
or U33301 (N_33301,N_31116,N_30536);
or U33302 (N_33302,N_31747,N_30500);
and U33303 (N_33303,N_30335,N_30450);
nor U33304 (N_33304,N_31489,N_31163);
and U33305 (N_33305,N_30510,N_31860);
nor U33306 (N_33306,N_31864,N_30220);
and U33307 (N_33307,N_31857,N_31352);
and U33308 (N_33308,N_31170,N_30355);
xor U33309 (N_33309,N_30308,N_30048);
and U33310 (N_33310,N_31868,N_30462);
or U33311 (N_33311,N_30452,N_30935);
and U33312 (N_33312,N_31560,N_30500);
or U33313 (N_33313,N_30975,N_31379);
or U33314 (N_33314,N_30487,N_30303);
or U33315 (N_33315,N_31644,N_31386);
nor U33316 (N_33316,N_31152,N_31291);
xor U33317 (N_33317,N_30526,N_31975);
or U33318 (N_33318,N_31227,N_31615);
nor U33319 (N_33319,N_30351,N_31317);
or U33320 (N_33320,N_30022,N_31960);
and U33321 (N_33321,N_30061,N_30703);
xnor U33322 (N_33322,N_30553,N_31515);
or U33323 (N_33323,N_31098,N_31541);
and U33324 (N_33324,N_30064,N_30338);
or U33325 (N_33325,N_31630,N_31976);
or U33326 (N_33326,N_30645,N_30004);
nand U33327 (N_33327,N_30274,N_30758);
nand U33328 (N_33328,N_31226,N_30045);
and U33329 (N_33329,N_31939,N_31737);
xnor U33330 (N_33330,N_31639,N_30651);
nand U33331 (N_33331,N_30838,N_31338);
nor U33332 (N_33332,N_30683,N_31061);
nor U33333 (N_33333,N_31912,N_31966);
or U33334 (N_33334,N_31284,N_31520);
or U33335 (N_33335,N_31990,N_31943);
and U33336 (N_33336,N_30322,N_30235);
nand U33337 (N_33337,N_30254,N_30463);
or U33338 (N_33338,N_31435,N_31449);
nand U33339 (N_33339,N_31549,N_31793);
xor U33340 (N_33340,N_30807,N_31906);
nor U33341 (N_33341,N_30681,N_31257);
and U33342 (N_33342,N_31786,N_30027);
nor U33343 (N_33343,N_31102,N_31261);
or U33344 (N_33344,N_31845,N_31606);
and U33345 (N_33345,N_31097,N_30085);
and U33346 (N_33346,N_31134,N_30213);
or U33347 (N_33347,N_30099,N_30597);
xnor U33348 (N_33348,N_31476,N_30815);
nor U33349 (N_33349,N_31227,N_31596);
nand U33350 (N_33350,N_31930,N_30351);
nand U33351 (N_33351,N_31462,N_30765);
nand U33352 (N_33352,N_31923,N_31985);
nor U33353 (N_33353,N_30824,N_30210);
and U33354 (N_33354,N_30322,N_30587);
and U33355 (N_33355,N_31056,N_31040);
or U33356 (N_33356,N_30918,N_31003);
xnor U33357 (N_33357,N_30209,N_30256);
xnor U33358 (N_33358,N_30962,N_31232);
nor U33359 (N_33359,N_30474,N_31283);
nand U33360 (N_33360,N_31505,N_31390);
and U33361 (N_33361,N_30009,N_31904);
or U33362 (N_33362,N_31405,N_31701);
nor U33363 (N_33363,N_30183,N_30934);
nor U33364 (N_33364,N_30332,N_31598);
or U33365 (N_33365,N_30126,N_30438);
or U33366 (N_33366,N_30155,N_30132);
nand U33367 (N_33367,N_31470,N_30550);
xor U33368 (N_33368,N_30740,N_31660);
and U33369 (N_33369,N_31346,N_31178);
and U33370 (N_33370,N_30396,N_30828);
nand U33371 (N_33371,N_31624,N_30438);
nand U33372 (N_33372,N_31270,N_30636);
and U33373 (N_33373,N_31198,N_30776);
nand U33374 (N_33374,N_31866,N_30741);
nand U33375 (N_33375,N_31986,N_30901);
xnor U33376 (N_33376,N_31701,N_31601);
xor U33377 (N_33377,N_30926,N_31892);
and U33378 (N_33378,N_30747,N_30000);
nand U33379 (N_33379,N_31642,N_31463);
nand U33380 (N_33380,N_30642,N_30628);
xor U33381 (N_33381,N_31856,N_31481);
xor U33382 (N_33382,N_30916,N_30413);
nand U33383 (N_33383,N_30999,N_31469);
xor U33384 (N_33384,N_31672,N_31719);
nor U33385 (N_33385,N_31144,N_30004);
nor U33386 (N_33386,N_31701,N_30214);
or U33387 (N_33387,N_31749,N_31685);
nor U33388 (N_33388,N_30620,N_30173);
xor U33389 (N_33389,N_30612,N_31172);
and U33390 (N_33390,N_31378,N_31508);
nor U33391 (N_33391,N_30605,N_30669);
nand U33392 (N_33392,N_30265,N_31478);
nand U33393 (N_33393,N_31784,N_31816);
xnor U33394 (N_33394,N_31533,N_31490);
and U33395 (N_33395,N_31180,N_30536);
and U33396 (N_33396,N_31014,N_30889);
nand U33397 (N_33397,N_30501,N_31284);
or U33398 (N_33398,N_31076,N_31688);
nand U33399 (N_33399,N_31613,N_30172);
xnor U33400 (N_33400,N_31678,N_31270);
nand U33401 (N_33401,N_31792,N_30767);
nor U33402 (N_33402,N_30091,N_31584);
xor U33403 (N_33403,N_30117,N_30239);
xnor U33404 (N_33404,N_30502,N_31575);
or U33405 (N_33405,N_31379,N_30839);
xnor U33406 (N_33406,N_31997,N_31545);
nor U33407 (N_33407,N_31835,N_30748);
nand U33408 (N_33408,N_31901,N_30494);
and U33409 (N_33409,N_30099,N_30287);
or U33410 (N_33410,N_31114,N_31591);
nor U33411 (N_33411,N_31284,N_31651);
nor U33412 (N_33412,N_31665,N_31877);
and U33413 (N_33413,N_31979,N_31531);
xor U33414 (N_33414,N_30014,N_31726);
nor U33415 (N_33415,N_30772,N_30153);
nor U33416 (N_33416,N_31030,N_31672);
or U33417 (N_33417,N_30084,N_30912);
xnor U33418 (N_33418,N_31653,N_31496);
nand U33419 (N_33419,N_30356,N_30518);
nand U33420 (N_33420,N_30518,N_30223);
nand U33421 (N_33421,N_31585,N_31219);
nor U33422 (N_33422,N_31786,N_30454);
xor U33423 (N_33423,N_31310,N_30789);
nand U33424 (N_33424,N_31513,N_31462);
nand U33425 (N_33425,N_30483,N_30029);
nand U33426 (N_33426,N_30862,N_30663);
and U33427 (N_33427,N_31837,N_30148);
xnor U33428 (N_33428,N_30753,N_30322);
nand U33429 (N_33429,N_30547,N_31401);
or U33430 (N_33430,N_31356,N_30622);
or U33431 (N_33431,N_31512,N_30652);
nand U33432 (N_33432,N_30468,N_30823);
nor U33433 (N_33433,N_31015,N_31509);
and U33434 (N_33434,N_30447,N_31700);
xnor U33435 (N_33435,N_31097,N_31254);
and U33436 (N_33436,N_31309,N_30488);
and U33437 (N_33437,N_30390,N_31016);
nor U33438 (N_33438,N_31872,N_30666);
nand U33439 (N_33439,N_30129,N_31266);
nand U33440 (N_33440,N_31713,N_30079);
or U33441 (N_33441,N_30112,N_30883);
or U33442 (N_33442,N_31836,N_31393);
or U33443 (N_33443,N_31852,N_31382);
and U33444 (N_33444,N_30087,N_31969);
nor U33445 (N_33445,N_31296,N_31531);
nor U33446 (N_33446,N_31945,N_31436);
nor U33447 (N_33447,N_31818,N_31690);
and U33448 (N_33448,N_31286,N_31178);
nor U33449 (N_33449,N_30764,N_31516);
and U33450 (N_33450,N_31069,N_30820);
and U33451 (N_33451,N_30903,N_30262);
xor U33452 (N_33452,N_31362,N_31996);
nor U33453 (N_33453,N_30497,N_31318);
xor U33454 (N_33454,N_30348,N_30361);
or U33455 (N_33455,N_31086,N_31483);
and U33456 (N_33456,N_31522,N_31915);
and U33457 (N_33457,N_31521,N_30728);
and U33458 (N_33458,N_30153,N_31569);
nand U33459 (N_33459,N_30365,N_30752);
nor U33460 (N_33460,N_31890,N_31476);
nor U33461 (N_33461,N_31616,N_30432);
nor U33462 (N_33462,N_30643,N_31009);
nand U33463 (N_33463,N_30237,N_31652);
and U33464 (N_33464,N_31473,N_30454);
xor U33465 (N_33465,N_31837,N_30582);
nand U33466 (N_33466,N_30558,N_30712);
xnor U33467 (N_33467,N_30287,N_30235);
and U33468 (N_33468,N_31345,N_31346);
and U33469 (N_33469,N_30773,N_30799);
and U33470 (N_33470,N_30899,N_31159);
nor U33471 (N_33471,N_31787,N_30757);
xor U33472 (N_33472,N_31531,N_31655);
xor U33473 (N_33473,N_30561,N_31008);
xnor U33474 (N_33474,N_31455,N_30716);
and U33475 (N_33475,N_30324,N_31960);
nand U33476 (N_33476,N_30053,N_30695);
xor U33477 (N_33477,N_31685,N_30349);
and U33478 (N_33478,N_31617,N_30176);
nor U33479 (N_33479,N_31268,N_30458);
nand U33480 (N_33480,N_30516,N_30255);
or U33481 (N_33481,N_31199,N_30489);
xnor U33482 (N_33482,N_30990,N_31062);
xor U33483 (N_33483,N_31200,N_30228);
and U33484 (N_33484,N_31476,N_30136);
or U33485 (N_33485,N_31096,N_30499);
and U33486 (N_33486,N_31807,N_30179);
or U33487 (N_33487,N_31702,N_31165);
xnor U33488 (N_33488,N_31030,N_30236);
nor U33489 (N_33489,N_31637,N_31470);
or U33490 (N_33490,N_31396,N_31020);
or U33491 (N_33491,N_30241,N_30242);
and U33492 (N_33492,N_30645,N_30944);
nand U33493 (N_33493,N_31146,N_31622);
or U33494 (N_33494,N_31208,N_31249);
xor U33495 (N_33495,N_30190,N_30389);
xor U33496 (N_33496,N_31953,N_31939);
or U33497 (N_33497,N_30004,N_30979);
nor U33498 (N_33498,N_30425,N_30854);
nor U33499 (N_33499,N_31605,N_31430);
or U33500 (N_33500,N_30140,N_30046);
nor U33501 (N_33501,N_31956,N_31120);
nor U33502 (N_33502,N_31142,N_30092);
or U33503 (N_33503,N_30302,N_30929);
xnor U33504 (N_33504,N_30144,N_30430);
nand U33505 (N_33505,N_31668,N_30400);
nor U33506 (N_33506,N_31401,N_30051);
nand U33507 (N_33507,N_31594,N_31593);
nand U33508 (N_33508,N_31859,N_30114);
or U33509 (N_33509,N_31557,N_31200);
nor U33510 (N_33510,N_30163,N_30735);
nand U33511 (N_33511,N_31405,N_31343);
or U33512 (N_33512,N_31549,N_30563);
xnor U33513 (N_33513,N_30598,N_31299);
or U33514 (N_33514,N_30067,N_31512);
nor U33515 (N_33515,N_30405,N_31651);
or U33516 (N_33516,N_31951,N_31187);
or U33517 (N_33517,N_31674,N_31118);
nor U33518 (N_33518,N_31940,N_31755);
and U33519 (N_33519,N_30275,N_30205);
xor U33520 (N_33520,N_30991,N_30036);
nor U33521 (N_33521,N_31883,N_30369);
nand U33522 (N_33522,N_30814,N_31296);
nand U33523 (N_33523,N_30672,N_30412);
xor U33524 (N_33524,N_31265,N_30477);
or U33525 (N_33525,N_30271,N_30618);
nand U33526 (N_33526,N_31621,N_30883);
or U33527 (N_33527,N_30672,N_30933);
nand U33528 (N_33528,N_31992,N_31592);
or U33529 (N_33529,N_30255,N_30738);
nor U33530 (N_33530,N_30803,N_31434);
and U33531 (N_33531,N_30585,N_31448);
or U33532 (N_33532,N_30501,N_31042);
nor U33533 (N_33533,N_30000,N_30309);
xor U33534 (N_33534,N_30013,N_30072);
nand U33535 (N_33535,N_31631,N_31825);
nor U33536 (N_33536,N_30973,N_30752);
and U33537 (N_33537,N_30383,N_30273);
or U33538 (N_33538,N_31081,N_30784);
and U33539 (N_33539,N_31369,N_30101);
or U33540 (N_33540,N_31120,N_30290);
and U33541 (N_33541,N_31297,N_31725);
and U33542 (N_33542,N_30722,N_30838);
xor U33543 (N_33543,N_31324,N_31061);
nor U33544 (N_33544,N_30968,N_31849);
nor U33545 (N_33545,N_30785,N_31071);
nand U33546 (N_33546,N_30687,N_31608);
nor U33547 (N_33547,N_30281,N_31206);
xnor U33548 (N_33548,N_30676,N_31711);
and U33549 (N_33549,N_30906,N_31148);
nor U33550 (N_33550,N_30014,N_31140);
and U33551 (N_33551,N_30714,N_31146);
nor U33552 (N_33552,N_31550,N_30510);
xnor U33553 (N_33553,N_30871,N_31605);
nand U33554 (N_33554,N_30401,N_30741);
and U33555 (N_33555,N_30301,N_31733);
xor U33556 (N_33556,N_30816,N_31415);
xor U33557 (N_33557,N_30069,N_30402);
and U33558 (N_33558,N_30603,N_30879);
nand U33559 (N_33559,N_31141,N_31629);
nor U33560 (N_33560,N_31698,N_31644);
xor U33561 (N_33561,N_30051,N_31477);
or U33562 (N_33562,N_30277,N_31038);
or U33563 (N_33563,N_30923,N_31491);
or U33564 (N_33564,N_31018,N_31681);
or U33565 (N_33565,N_31212,N_31160);
nand U33566 (N_33566,N_31169,N_30746);
nand U33567 (N_33567,N_31195,N_31893);
nor U33568 (N_33568,N_30977,N_30387);
and U33569 (N_33569,N_30462,N_30524);
xor U33570 (N_33570,N_31029,N_30842);
and U33571 (N_33571,N_31791,N_30177);
and U33572 (N_33572,N_30617,N_30809);
nand U33573 (N_33573,N_31322,N_31222);
xnor U33574 (N_33574,N_31648,N_31320);
and U33575 (N_33575,N_30823,N_31292);
nor U33576 (N_33576,N_31269,N_30658);
xnor U33577 (N_33577,N_31287,N_30228);
or U33578 (N_33578,N_31457,N_31296);
nand U33579 (N_33579,N_30994,N_30303);
nor U33580 (N_33580,N_30194,N_31093);
xnor U33581 (N_33581,N_31465,N_31888);
or U33582 (N_33582,N_31797,N_31551);
xor U33583 (N_33583,N_30706,N_31489);
or U33584 (N_33584,N_30517,N_30180);
or U33585 (N_33585,N_30214,N_30166);
and U33586 (N_33586,N_31992,N_30720);
nand U33587 (N_33587,N_31373,N_30469);
nand U33588 (N_33588,N_30542,N_30278);
and U33589 (N_33589,N_30202,N_30056);
or U33590 (N_33590,N_30943,N_30029);
xor U33591 (N_33591,N_31285,N_31085);
nand U33592 (N_33592,N_30831,N_30242);
nor U33593 (N_33593,N_30011,N_31915);
nand U33594 (N_33594,N_31715,N_31519);
xnor U33595 (N_33595,N_30017,N_31885);
nor U33596 (N_33596,N_31406,N_31512);
and U33597 (N_33597,N_30096,N_30223);
and U33598 (N_33598,N_30392,N_30622);
nand U33599 (N_33599,N_30119,N_31597);
nor U33600 (N_33600,N_30297,N_31282);
and U33601 (N_33601,N_30242,N_30445);
nand U33602 (N_33602,N_31699,N_30650);
xnor U33603 (N_33603,N_31850,N_30629);
and U33604 (N_33604,N_30419,N_30487);
nand U33605 (N_33605,N_30356,N_30884);
or U33606 (N_33606,N_30868,N_30787);
nand U33607 (N_33607,N_31493,N_30474);
nor U33608 (N_33608,N_30700,N_31862);
and U33609 (N_33609,N_31043,N_30627);
nor U33610 (N_33610,N_30137,N_30292);
xnor U33611 (N_33611,N_31167,N_31420);
nand U33612 (N_33612,N_30621,N_30396);
xor U33613 (N_33613,N_31557,N_30559);
nand U33614 (N_33614,N_31383,N_30389);
nor U33615 (N_33615,N_31427,N_31992);
or U33616 (N_33616,N_31104,N_31877);
nor U33617 (N_33617,N_31753,N_31697);
or U33618 (N_33618,N_30563,N_31510);
and U33619 (N_33619,N_31538,N_30434);
or U33620 (N_33620,N_31960,N_30140);
and U33621 (N_33621,N_31557,N_30155);
nand U33622 (N_33622,N_31301,N_31407);
nand U33623 (N_33623,N_31391,N_30130);
nor U33624 (N_33624,N_31956,N_31835);
nand U33625 (N_33625,N_31606,N_30253);
and U33626 (N_33626,N_31133,N_30820);
xor U33627 (N_33627,N_30301,N_31634);
and U33628 (N_33628,N_30877,N_31154);
xnor U33629 (N_33629,N_31834,N_31401);
xnor U33630 (N_33630,N_31268,N_31625);
and U33631 (N_33631,N_30020,N_30548);
nand U33632 (N_33632,N_31903,N_30488);
nand U33633 (N_33633,N_31132,N_30853);
or U33634 (N_33634,N_30091,N_31336);
xnor U33635 (N_33635,N_31959,N_30908);
xnor U33636 (N_33636,N_31153,N_31144);
and U33637 (N_33637,N_30055,N_30391);
nand U33638 (N_33638,N_31754,N_30615);
xor U33639 (N_33639,N_31204,N_31463);
and U33640 (N_33640,N_31001,N_31681);
or U33641 (N_33641,N_30758,N_30845);
nand U33642 (N_33642,N_31270,N_31784);
or U33643 (N_33643,N_30190,N_30604);
nor U33644 (N_33644,N_30597,N_30538);
nand U33645 (N_33645,N_30741,N_30047);
nand U33646 (N_33646,N_30341,N_30032);
or U33647 (N_33647,N_31041,N_30629);
xor U33648 (N_33648,N_31356,N_30589);
and U33649 (N_33649,N_30412,N_31961);
xor U33650 (N_33650,N_31815,N_30714);
nand U33651 (N_33651,N_31637,N_31553);
and U33652 (N_33652,N_30117,N_30307);
nand U33653 (N_33653,N_30345,N_31360);
nand U33654 (N_33654,N_30450,N_30713);
or U33655 (N_33655,N_31067,N_31772);
and U33656 (N_33656,N_30455,N_31036);
or U33657 (N_33657,N_30237,N_30736);
nor U33658 (N_33658,N_30982,N_30695);
nor U33659 (N_33659,N_31161,N_30764);
and U33660 (N_33660,N_30405,N_31131);
and U33661 (N_33661,N_30480,N_31532);
xnor U33662 (N_33662,N_30439,N_31289);
xnor U33663 (N_33663,N_30998,N_30960);
nand U33664 (N_33664,N_31996,N_30340);
nand U33665 (N_33665,N_31912,N_30513);
xnor U33666 (N_33666,N_31664,N_31984);
xnor U33667 (N_33667,N_31466,N_31372);
nand U33668 (N_33668,N_30779,N_31239);
nor U33669 (N_33669,N_31665,N_30242);
nor U33670 (N_33670,N_31696,N_31234);
nand U33671 (N_33671,N_31640,N_31008);
xnor U33672 (N_33672,N_31822,N_31692);
xor U33673 (N_33673,N_30441,N_31100);
nor U33674 (N_33674,N_31082,N_31917);
nor U33675 (N_33675,N_30350,N_30467);
or U33676 (N_33676,N_30584,N_31578);
nor U33677 (N_33677,N_30444,N_31546);
nor U33678 (N_33678,N_31972,N_30726);
nor U33679 (N_33679,N_31126,N_30496);
xnor U33680 (N_33680,N_31395,N_31054);
and U33681 (N_33681,N_31197,N_30376);
and U33682 (N_33682,N_30638,N_30010);
nand U33683 (N_33683,N_30276,N_30447);
nand U33684 (N_33684,N_31909,N_31509);
or U33685 (N_33685,N_30789,N_31704);
nor U33686 (N_33686,N_30308,N_30911);
xnor U33687 (N_33687,N_31565,N_31274);
and U33688 (N_33688,N_31192,N_31689);
and U33689 (N_33689,N_30835,N_31247);
nand U33690 (N_33690,N_30909,N_31879);
xnor U33691 (N_33691,N_30640,N_31810);
and U33692 (N_33692,N_31230,N_31986);
nor U33693 (N_33693,N_31858,N_30684);
xor U33694 (N_33694,N_30294,N_31494);
nor U33695 (N_33695,N_31665,N_30599);
nor U33696 (N_33696,N_30424,N_31292);
and U33697 (N_33697,N_30818,N_30701);
xnor U33698 (N_33698,N_30338,N_31622);
nor U33699 (N_33699,N_31258,N_30472);
xnor U33700 (N_33700,N_31058,N_31155);
nand U33701 (N_33701,N_31948,N_31801);
nor U33702 (N_33702,N_31105,N_30033);
and U33703 (N_33703,N_31805,N_30355);
nand U33704 (N_33704,N_30834,N_30630);
nand U33705 (N_33705,N_30249,N_30596);
or U33706 (N_33706,N_30490,N_30430);
xor U33707 (N_33707,N_31864,N_30059);
nand U33708 (N_33708,N_31899,N_31016);
nand U33709 (N_33709,N_30358,N_30351);
or U33710 (N_33710,N_30501,N_30768);
nand U33711 (N_33711,N_30540,N_31191);
and U33712 (N_33712,N_30038,N_30661);
nand U33713 (N_33713,N_31054,N_30899);
nor U33714 (N_33714,N_30541,N_31396);
xnor U33715 (N_33715,N_30791,N_31149);
xnor U33716 (N_33716,N_30229,N_31939);
nand U33717 (N_33717,N_31928,N_31290);
or U33718 (N_33718,N_30053,N_31525);
or U33719 (N_33719,N_30217,N_31888);
xor U33720 (N_33720,N_31665,N_31922);
nand U33721 (N_33721,N_31612,N_30818);
xnor U33722 (N_33722,N_31941,N_31141);
nor U33723 (N_33723,N_30902,N_31995);
or U33724 (N_33724,N_31257,N_31447);
and U33725 (N_33725,N_31256,N_31171);
nor U33726 (N_33726,N_31973,N_31404);
nor U33727 (N_33727,N_31562,N_31964);
nor U33728 (N_33728,N_30200,N_30624);
nand U33729 (N_33729,N_30633,N_30090);
and U33730 (N_33730,N_30943,N_30013);
nor U33731 (N_33731,N_31189,N_31941);
or U33732 (N_33732,N_30251,N_31928);
xor U33733 (N_33733,N_31751,N_31502);
nand U33734 (N_33734,N_31374,N_31898);
or U33735 (N_33735,N_30458,N_30175);
xor U33736 (N_33736,N_30934,N_31539);
xor U33737 (N_33737,N_30188,N_31115);
nor U33738 (N_33738,N_31198,N_31276);
nor U33739 (N_33739,N_31598,N_31139);
and U33740 (N_33740,N_30758,N_31775);
nor U33741 (N_33741,N_31396,N_30597);
or U33742 (N_33742,N_30044,N_31559);
or U33743 (N_33743,N_30874,N_30357);
nor U33744 (N_33744,N_31657,N_30770);
or U33745 (N_33745,N_30368,N_31816);
and U33746 (N_33746,N_31272,N_31706);
nor U33747 (N_33747,N_31272,N_30287);
or U33748 (N_33748,N_30281,N_31505);
or U33749 (N_33749,N_30703,N_31726);
nand U33750 (N_33750,N_30829,N_30096);
nor U33751 (N_33751,N_31866,N_31529);
or U33752 (N_33752,N_30853,N_30198);
nor U33753 (N_33753,N_31069,N_31999);
or U33754 (N_33754,N_31641,N_31049);
xnor U33755 (N_33755,N_31045,N_31512);
and U33756 (N_33756,N_31602,N_31046);
nand U33757 (N_33757,N_30200,N_30751);
or U33758 (N_33758,N_31011,N_31879);
or U33759 (N_33759,N_31059,N_31365);
nand U33760 (N_33760,N_31737,N_31611);
nor U33761 (N_33761,N_30961,N_31305);
or U33762 (N_33762,N_30793,N_31223);
nand U33763 (N_33763,N_31752,N_30876);
xor U33764 (N_33764,N_30991,N_30686);
nand U33765 (N_33765,N_31148,N_31953);
or U33766 (N_33766,N_30921,N_30683);
nand U33767 (N_33767,N_30479,N_30576);
xor U33768 (N_33768,N_30700,N_31295);
or U33769 (N_33769,N_30823,N_30760);
nand U33770 (N_33770,N_31267,N_31531);
nand U33771 (N_33771,N_30108,N_31403);
nor U33772 (N_33772,N_31322,N_31739);
nand U33773 (N_33773,N_30207,N_30490);
nand U33774 (N_33774,N_31057,N_30147);
xor U33775 (N_33775,N_30681,N_31776);
nand U33776 (N_33776,N_31358,N_30510);
nand U33777 (N_33777,N_30299,N_31080);
or U33778 (N_33778,N_30861,N_30037);
and U33779 (N_33779,N_31282,N_30192);
nor U33780 (N_33780,N_30100,N_31051);
xnor U33781 (N_33781,N_30164,N_31785);
nand U33782 (N_33782,N_30251,N_31513);
xnor U33783 (N_33783,N_30549,N_31435);
nand U33784 (N_33784,N_31910,N_30820);
xor U33785 (N_33785,N_31151,N_30508);
and U33786 (N_33786,N_30010,N_30263);
nand U33787 (N_33787,N_30319,N_31544);
nand U33788 (N_33788,N_30436,N_30869);
nor U33789 (N_33789,N_31377,N_31653);
nor U33790 (N_33790,N_30805,N_30324);
and U33791 (N_33791,N_30072,N_31928);
and U33792 (N_33792,N_31434,N_30362);
nand U33793 (N_33793,N_31210,N_31985);
nand U33794 (N_33794,N_31868,N_31227);
xor U33795 (N_33795,N_31574,N_30621);
and U33796 (N_33796,N_30326,N_30250);
xnor U33797 (N_33797,N_31982,N_31223);
nand U33798 (N_33798,N_31024,N_31552);
nand U33799 (N_33799,N_30826,N_31826);
and U33800 (N_33800,N_31685,N_31777);
nand U33801 (N_33801,N_31854,N_30843);
or U33802 (N_33802,N_30434,N_31614);
or U33803 (N_33803,N_30138,N_30012);
nand U33804 (N_33804,N_30026,N_30334);
nor U33805 (N_33805,N_31640,N_31286);
or U33806 (N_33806,N_30176,N_31685);
or U33807 (N_33807,N_31976,N_31295);
and U33808 (N_33808,N_31567,N_31858);
and U33809 (N_33809,N_31287,N_30599);
and U33810 (N_33810,N_31395,N_31057);
nand U33811 (N_33811,N_31075,N_31873);
or U33812 (N_33812,N_31161,N_30677);
nor U33813 (N_33813,N_31603,N_31734);
nor U33814 (N_33814,N_30955,N_31156);
and U33815 (N_33815,N_31927,N_30543);
xnor U33816 (N_33816,N_30655,N_31343);
and U33817 (N_33817,N_31947,N_31907);
or U33818 (N_33818,N_30152,N_30066);
nor U33819 (N_33819,N_31868,N_31265);
xnor U33820 (N_33820,N_30282,N_30441);
and U33821 (N_33821,N_30311,N_30957);
and U33822 (N_33822,N_30465,N_30865);
or U33823 (N_33823,N_31176,N_30516);
nand U33824 (N_33824,N_31714,N_30165);
nor U33825 (N_33825,N_30610,N_31586);
or U33826 (N_33826,N_31443,N_30422);
nand U33827 (N_33827,N_30728,N_30341);
nor U33828 (N_33828,N_31130,N_30864);
and U33829 (N_33829,N_30135,N_30866);
nor U33830 (N_33830,N_31728,N_31984);
or U33831 (N_33831,N_31162,N_30767);
or U33832 (N_33832,N_31678,N_31811);
or U33833 (N_33833,N_31509,N_30902);
nand U33834 (N_33834,N_30671,N_31207);
and U33835 (N_33835,N_31004,N_30555);
nor U33836 (N_33836,N_30354,N_31465);
nand U33837 (N_33837,N_31037,N_31644);
nand U33838 (N_33838,N_31173,N_30275);
xor U33839 (N_33839,N_31981,N_30051);
xor U33840 (N_33840,N_31077,N_30295);
nand U33841 (N_33841,N_30632,N_30343);
and U33842 (N_33842,N_31694,N_30941);
nand U33843 (N_33843,N_30081,N_30946);
or U33844 (N_33844,N_31058,N_31365);
xnor U33845 (N_33845,N_31948,N_30970);
or U33846 (N_33846,N_30899,N_31978);
and U33847 (N_33847,N_30336,N_30869);
or U33848 (N_33848,N_31801,N_31200);
and U33849 (N_33849,N_30564,N_31489);
or U33850 (N_33850,N_31721,N_31885);
nor U33851 (N_33851,N_30233,N_31265);
nand U33852 (N_33852,N_30555,N_31745);
nor U33853 (N_33853,N_30993,N_31491);
or U33854 (N_33854,N_30455,N_30044);
nand U33855 (N_33855,N_30374,N_31046);
or U33856 (N_33856,N_30322,N_31862);
nand U33857 (N_33857,N_31030,N_31306);
nor U33858 (N_33858,N_30270,N_31484);
nor U33859 (N_33859,N_31948,N_31411);
or U33860 (N_33860,N_30761,N_31533);
and U33861 (N_33861,N_31611,N_31128);
nor U33862 (N_33862,N_31047,N_30447);
and U33863 (N_33863,N_30742,N_31029);
and U33864 (N_33864,N_30513,N_31339);
nand U33865 (N_33865,N_31798,N_31103);
nand U33866 (N_33866,N_30777,N_30763);
and U33867 (N_33867,N_30230,N_30106);
nor U33868 (N_33868,N_31127,N_30447);
nand U33869 (N_33869,N_31172,N_30555);
nor U33870 (N_33870,N_31720,N_31988);
and U33871 (N_33871,N_31136,N_30734);
nor U33872 (N_33872,N_31420,N_30884);
or U33873 (N_33873,N_31054,N_30279);
or U33874 (N_33874,N_31685,N_31844);
and U33875 (N_33875,N_30478,N_30456);
and U33876 (N_33876,N_30650,N_30713);
nand U33877 (N_33877,N_31085,N_30545);
and U33878 (N_33878,N_30920,N_31747);
and U33879 (N_33879,N_31976,N_31934);
nor U33880 (N_33880,N_30508,N_31730);
nor U33881 (N_33881,N_30386,N_30856);
nand U33882 (N_33882,N_30357,N_31608);
and U33883 (N_33883,N_31696,N_30739);
nor U33884 (N_33884,N_31711,N_31296);
xnor U33885 (N_33885,N_30378,N_31182);
nor U33886 (N_33886,N_31921,N_31771);
and U33887 (N_33887,N_30464,N_31791);
or U33888 (N_33888,N_30460,N_31620);
nor U33889 (N_33889,N_31773,N_30523);
and U33890 (N_33890,N_31204,N_31099);
and U33891 (N_33891,N_30435,N_30981);
and U33892 (N_33892,N_30181,N_30388);
xnor U33893 (N_33893,N_30363,N_31102);
xnor U33894 (N_33894,N_31103,N_30381);
nor U33895 (N_33895,N_31094,N_31659);
xor U33896 (N_33896,N_30592,N_31240);
nor U33897 (N_33897,N_31899,N_30355);
nor U33898 (N_33898,N_31450,N_30636);
and U33899 (N_33899,N_31659,N_30780);
nor U33900 (N_33900,N_30563,N_31612);
nand U33901 (N_33901,N_30263,N_30633);
nand U33902 (N_33902,N_30025,N_31896);
and U33903 (N_33903,N_31596,N_31007);
and U33904 (N_33904,N_30544,N_30346);
or U33905 (N_33905,N_31007,N_31572);
xnor U33906 (N_33906,N_30858,N_31928);
xnor U33907 (N_33907,N_30080,N_30926);
and U33908 (N_33908,N_31895,N_31751);
nand U33909 (N_33909,N_31752,N_30126);
nand U33910 (N_33910,N_30900,N_30222);
and U33911 (N_33911,N_31390,N_31614);
xnor U33912 (N_33912,N_31946,N_30012);
nand U33913 (N_33913,N_31839,N_31213);
nor U33914 (N_33914,N_30014,N_31822);
nand U33915 (N_33915,N_31941,N_31696);
or U33916 (N_33916,N_31853,N_30086);
xnor U33917 (N_33917,N_31192,N_30854);
nor U33918 (N_33918,N_31947,N_31540);
nand U33919 (N_33919,N_31780,N_31816);
nor U33920 (N_33920,N_31095,N_31783);
and U33921 (N_33921,N_30011,N_30311);
nor U33922 (N_33922,N_30073,N_31524);
and U33923 (N_33923,N_31413,N_30530);
and U33924 (N_33924,N_30484,N_31356);
nor U33925 (N_33925,N_31362,N_31344);
and U33926 (N_33926,N_31260,N_30622);
or U33927 (N_33927,N_30903,N_30782);
nand U33928 (N_33928,N_31339,N_31359);
and U33929 (N_33929,N_30283,N_31000);
nand U33930 (N_33930,N_31457,N_31295);
nand U33931 (N_33931,N_31375,N_31714);
or U33932 (N_33932,N_30112,N_31950);
xnor U33933 (N_33933,N_31826,N_31494);
and U33934 (N_33934,N_31726,N_31728);
xor U33935 (N_33935,N_31923,N_31429);
or U33936 (N_33936,N_30727,N_30550);
or U33937 (N_33937,N_30908,N_31083);
nor U33938 (N_33938,N_31729,N_31945);
nand U33939 (N_33939,N_30143,N_31654);
or U33940 (N_33940,N_30105,N_31796);
or U33941 (N_33941,N_30534,N_30644);
nand U33942 (N_33942,N_30831,N_30139);
nor U33943 (N_33943,N_31083,N_30915);
xor U33944 (N_33944,N_31901,N_30505);
nand U33945 (N_33945,N_30112,N_30911);
nand U33946 (N_33946,N_30898,N_31524);
nand U33947 (N_33947,N_31847,N_31939);
and U33948 (N_33948,N_30995,N_30642);
or U33949 (N_33949,N_31992,N_31868);
or U33950 (N_33950,N_30861,N_31924);
nor U33951 (N_33951,N_31880,N_31246);
xor U33952 (N_33952,N_30378,N_30412);
and U33953 (N_33953,N_31352,N_31055);
and U33954 (N_33954,N_31366,N_30750);
xnor U33955 (N_33955,N_31487,N_30964);
nand U33956 (N_33956,N_30222,N_31784);
nor U33957 (N_33957,N_31744,N_30925);
and U33958 (N_33958,N_31191,N_30715);
nor U33959 (N_33959,N_31682,N_31844);
or U33960 (N_33960,N_30185,N_31820);
nor U33961 (N_33961,N_31939,N_31963);
xnor U33962 (N_33962,N_30472,N_30510);
or U33963 (N_33963,N_31835,N_30002);
nand U33964 (N_33964,N_30785,N_30534);
xor U33965 (N_33965,N_31622,N_31181);
or U33966 (N_33966,N_31568,N_31153);
xor U33967 (N_33967,N_30746,N_31117);
nor U33968 (N_33968,N_31789,N_30652);
and U33969 (N_33969,N_31619,N_31063);
nor U33970 (N_33970,N_30016,N_30019);
nand U33971 (N_33971,N_31807,N_30571);
and U33972 (N_33972,N_30669,N_31338);
nor U33973 (N_33973,N_30703,N_31507);
or U33974 (N_33974,N_31784,N_31081);
or U33975 (N_33975,N_31549,N_30014);
nor U33976 (N_33976,N_31541,N_30887);
or U33977 (N_33977,N_30390,N_31164);
nor U33978 (N_33978,N_30924,N_31024);
xnor U33979 (N_33979,N_31657,N_30427);
or U33980 (N_33980,N_31085,N_31183);
or U33981 (N_33981,N_31337,N_31406);
xor U33982 (N_33982,N_31169,N_30200);
nor U33983 (N_33983,N_31592,N_31948);
nand U33984 (N_33984,N_30650,N_30068);
nor U33985 (N_33985,N_31300,N_30547);
nor U33986 (N_33986,N_30491,N_31025);
nor U33987 (N_33987,N_30531,N_31804);
nor U33988 (N_33988,N_31443,N_30145);
xor U33989 (N_33989,N_30289,N_30480);
nand U33990 (N_33990,N_30038,N_30859);
and U33991 (N_33991,N_30501,N_30744);
xnor U33992 (N_33992,N_30737,N_30735);
xor U33993 (N_33993,N_31750,N_31077);
or U33994 (N_33994,N_30133,N_30682);
nor U33995 (N_33995,N_30994,N_30174);
nor U33996 (N_33996,N_30894,N_31278);
nor U33997 (N_33997,N_31459,N_31948);
and U33998 (N_33998,N_30484,N_31526);
xor U33999 (N_33999,N_30938,N_31558);
nand U34000 (N_34000,N_32871,N_33899);
or U34001 (N_34001,N_32318,N_32838);
nor U34002 (N_34002,N_32135,N_33693);
or U34003 (N_34003,N_33913,N_32757);
or U34004 (N_34004,N_33032,N_32881);
nor U34005 (N_34005,N_33858,N_33074);
or U34006 (N_34006,N_33796,N_33099);
and U34007 (N_34007,N_32493,N_32533);
nor U34008 (N_34008,N_33713,N_33878);
nand U34009 (N_34009,N_32197,N_32096);
nor U34010 (N_34010,N_33321,N_32547);
nand U34011 (N_34011,N_33272,N_32646);
xor U34012 (N_34012,N_33060,N_33153);
or U34013 (N_34013,N_33541,N_32637);
xor U34014 (N_34014,N_32216,N_33277);
nand U34015 (N_34015,N_33230,N_33786);
nor U34016 (N_34016,N_33160,N_32352);
or U34017 (N_34017,N_33577,N_33138);
nand U34018 (N_34018,N_32449,N_32589);
or U34019 (N_34019,N_32633,N_33283);
nor U34020 (N_34020,N_33871,N_32179);
and U34021 (N_34021,N_33753,N_32190);
or U34022 (N_34022,N_33891,N_33831);
or U34023 (N_34023,N_32319,N_32950);
or U34024 (N_34024,N_32685,N_33194);
or U34025 (N_34025,N_32000,N_32971);
nand U34026 (N_34026,N_33918,N_33555);
nor U34027 (N_34027,N_32123,N_32867);
and U34028 (N_34028,N_33680,N_33136);
nor U34029 (N_34029,N_32500,N_33872);
nand U34030 (N_34030,N_33788,N_32879);
nor U34031 (N_34031,N_33968,N_32453);
and U34032 (N_34032,N_33125,N_33288);
xor U34033 (N_34033,N_32237,N_33806);
or U34034 (N_34034,N_33925,N_33742);
xnor U34035 (N_34035,N_33972,N_33076);
nor U34036 (N_34036,N_32969,N_33839);
and U34037 (N_34037,N_32606,N_33107);
nand U34038 (N_34038,N_33428,N_33904);
nand U34039 (N_34039,N_32035,N_33824);
xor U34040 (N_34040,N_33111,N_33670);
nor U34041 (N_34041,N_33731,N_32566);
nor U34042 (N_34042,N_32718,N_32667);
nor U34043 (N_34043,N_32717,N_32555);
xnor U34044 (N_34044,N_33493,N_33148);
and U34045 (N_34045,N_33236,N_33095);
and U34046 (N_34046,N_32704,N_32465);
or U34047 (N_34047,N_32174,N_32306);
nor U34048 (N_34048,N_33479,N_32368);
nor U34049 (N_34049,N_33695,N_33237);
nand U34050 (N_34050,N_32726,N_32150);
or U34051 (N_34051,N_33619,N_33378);
nand U34052 (N_34052,N_32999,N_32719);
and U34053 (N_34053,N_32787,N_33804);
and U34054 (N_34054,N_33643,N_32145);
nand U34055 (N_34055,N_33291,N_33984);
nor U34056 (N_34056,N_32082,N_32599);
nor U34057 (N_34057,N_33710,N_33275);
nand U34058 (N_34058,N_32085,N_32665);
or U34059 (N_34059,N_32042,N_33654);
or U34060 (N_34060,N_33084,N_32673);
nand U34061 (N_34061,N_32182,N_32040);
nor U34062 (N_34062,N_33828,N_33309);
and U34063 (N_34063,N_33267,N_32399);
xnor U34064 (N_34064,N_32911,N_33652);
or U34065 (N_34065,N_32954,N_32086);
nor U34066 (N_34066,N_33343,N_32058);
xor U34067 (N_34067,N_33337,N_33265);
nor U34068 (N_34068,N_32217,N_32298);
and U34069 (N_34069,N_32476,N_33232);
nand U34070 (N_34070,N_32469,N_32025);
or U34071 (N_34071,N_32947,N_33108);
and U34072 (N_34072,N_33537,N_32391);
or U34073 (N_34073,N_32921,N_33412);
xnor U34074 (N_34074,N_32267,N_32546);
nand U34075 (N_34075,N_32367,N_32143);
xnor U34076 (N_34076,N_33874,N_32343);
or U34077 (N_34077,N_32048,N_32804);
xor U34078 (N_34078,N_33489,N_33519);
and U34079 (N_34079,N_33690,N_33249);
nor U34080 (N_34080,N_32608,N_32905);
or U34081 (N_34081,N_32842,N_33509);
nand U34082 (N_34082,N_33631,N_33386);
nor U34083 (N_34083,N_32003,N_33001);
nor U34084 (N_34084,N_32900,N_33761);
or U34085 (N_34085,N_32429,N_33988);
nor U34086 (N_34086,N_33305,N_33481);
or U34087 (N_34087,N_33186,N_32935);
or U34088 (N_34088,N_32055,N_33687);
nor U34089 (N_34089,N_32882,N_33764);
nor U34090 (N_34090,N_33461,N_32997);
and U34091 (N_34091,N_33682,N_32683);
xnor U34092 (N_34092,N_32419,N_33521);
nand U34093 (N_34093,N_33650,N_33420);
nand U34094 (N_34094,N_33030,N_32193);
or U34095 (N_34095,N_32266,N_33715);
xor U34096 (N_34096,N_33317,N_32528);
xnor U34097 (N_34097,N_32864,N_33864);
nand U34098 (N_34098,N_32295,N_32170);
and U34099 (N_34099,N_32962,N_33333);
xnor U34100 (N_34100,N_33532,N_32623);
and U34101 (N_34101,N_32617,N_33585);
nor U34102 (N_34102,N_32053,N_32549);
or U34103 (N_34103,N_32272,N_32264);
xor U34104 (N_34104,N_32274,N_32664);
nand U34105 (N_34105,N_33487,N_32551);
xnor U34106 (N_34106,N_32052,N_32092);
or U34107 (N_34107,N_32958,N_33868);
nand U34108 (N_34108,N_33953,N_32666);
nor U34109 (N_34109,N_33534,N_33402);
nor U34110 (N_34110,N_32990,N_33280);
or U34111 (N_34111,N_33573,N_33058);
nor U34112 (N_34112,N_32708,N_33971);
xor U34113 (N_34113,N_33188,N_32552);
or U34114 (N_34114,N_32998,N_32618);
nand U34115 (N_34115,N_33235,N_33331);
xor U34116 (N_34116,N_32894,N_33626);
or U34117 (N_34117,N_33314,N_32577);
xnor U34118 (N_34118,N_33934,N_33963);
nor U34119 (N_34119,N_33976,N_32723);
nand U34120 (N_34120,N_33370,N_33303);
xnor U34121 (N_34121,N_33007,N_32532);
nand U34122 (N_34122,N_33944,N_33444);
xnor U34123 (N_34123,N_32394,N_32627);
or U34124 (N_34124,N_32173,N_33967);
nand U34125 (N_34125,N_32927,N_32821);
or U34126 (N_34126,N_32372,N_32464);
xnor U34127 (N_34127,N_32856,N_32983);
or U34128 (N_34128,N_32545,N_33889);
or U34129 (N_34129,N_32426,N_33632);
or U34130 (N_34130,N_32575,N_33767);
or U34131 (N_34131,N_33085,N_32582);
nor U34132 (N_34132,N_32099,N_33132);
or U34133 (N_34133,N_33997,N_32460);
xnor U34134 (N_34134,N_33244,N_33008);
nor U34135 (N_34135,N_33578,N_32177);
nand U34136 (N_34136,N_32562,N_32258);
nor U34137 (N_34137,N_32303,N_33293);
and U34138 (N_34138,N_32713,N_33956);
nor U34139 (N_34139,N_33162,N_32231);
or U34140 (N_34140,N_32149,N_33676);
xor U34141 (N_34141,N_33596,N_32909);
or U34142 (N_34142,N_33453,N_32784);
or U34143 (N_34143,N_33109,N_32986);
xnor U34144 (N_34144,N_32317,N_32732);
and U34145 (N_34145,N_33214,N_32586);
xnor U34146 (N_34146,N_33310,N_32454);
nand U34147 (N_34147,N_33723,N_32014);
and U34148 (N_34148,N_32556,N_33430);
xor U34149 (N_34149,N_32915,N_32333);
xor U34150 (N_34150,N_32620,N_33141);
nand U34151 (N_34151,N_32913,N_32975);
nand U34152 (N_34152,N_32060,N_32591);
nor U34153 (N_34153,N_33556,N_33599);
nand U34154 (N_34154,N_33013,N_33339);
nand U34155 (N_34155,N_33510,N_33476);
or U34156 (N_34156,N_32166,N_33233);
nor U34157 (N_34157,N_33584,N_33583);
or U34158 (N_34158,N_32300,N_33165);
nand U34159 (N_34159,N_32679,N_32898);
nand U34160 (N_34160,N_33689,N_32373);
nand U34161 (N_34161,N_33175,N_32155);
and U34162 (N_34162,N_32697,N_32183);
xnor U34163 (N_34163,N_33221,N_33691);
nand U34164 (N_34164,N_32638,N_33973);
nor U34165 (N_34165,N_32891,N_32378);
and U34166 (N_34166,N_33135,N_32750);
or U34167 (N_34167,N_32428,N_32874);
or U34168 (N_34168,N_32758,N_33863);
or U34169 (N_34169,N_33250,N_32832);
or U34170 (N_34170,N_32824,N_32369);
and U34171 (N_34171,N_32316,N_32583);
or U34172 (N_34172,N_33524,N_33661);
xor U34173 (N_34173,N_32347,N_33762);
xnor U34174 (N_34174,N_32032,N_33719);
nor U34175 (N_34175,N_32105,N_32475);
or U34176 (N_34176,N_32111,N_33147);
nor U34177 (N_34177,N_33200,N_33876);
xor U34178 (N_34178,N_33717,N_32321);
nor U34179 (N_34179,N_33590,N_33780);
or U34180 (N_34180,N_32178,N_32030);
nand U34181 (N_34181,N_32939,N_32854);
nor U34182 (N_34182,N_33558,N_33102);
and U34183 (N_34183,N_32424,N_32213);
xnor U34184 (N_34184,N_33121,N_32201);
or U34185 (N_34185,N_33607,N_33993);
or U34186 (N_34186,N_33660,N_33455);
and U34187 (N_34187,N_33417,N_33808);
xor U34188 (N_34188,N_32792,N_33260);
or U34189 (N_34189,N_32595,N_33284);
or U34190 (N_34190,N_33618,N_33900);
or U34191 (N_34191,N_32108,N_33513);
or U34192 (N_34192,N_32341,N_33877);
nand U34193 (N_34193,N_33082,N_33729);
and U34194 (N_34194,N_32479,N_32794);
or U34195 (N_34195,N_33749,N_33087);
nand U34196 (N_34196,N_33127,N_33580);
nor U34197 (N_34197,N_32657,N_32271);
or U34198 (N_34198,N_33016,N_33543);
nor U34199 (N_34199,N_33367,N_33906);
nand U34200 (N_34200,N_33353,N_33002);
or U34201 (N_34201,N_32746,N_32406);
nand U34202 (N_34202,N_32539,N_32043);
nand U34203 (N_34203,N_32687,N_33166);
nor U34204 (N_34204,N_33300,N_33202);
or U34205 (N_34205,N_33189,N_33066);
nand U34206 (N_34206,N_33752,N_33604);
and U34207 (N_34207,N_33962,N_32840);
nand U34208 (N_34208,N_33168,N_32332);
nor U34209 (N_34209,N_33015,N_32379);
nand U34210 (N_34210,N_32561,N_33748);
xor U34211 (N_34211,N_32356,N_33301);
nor U34212 (N_34212,N_33021,N_33570);
or U34213 (N_34213,N_32313,N_33564);
xor U34214 (N_34214,N_32560,N_33139);
and U34215 (N_34215,N_32579,N_32634);
and U34216 (N_34216,N_32194,N_32045);
or U34217 (N_34217,N_32389,N_33491);
nor U34218 (N_34218,N_33949,N_33811);
nand U34219 (N_34219,N_33268,N_32243);
and U34220 (N_34220,N_33485,N_33329);
and U34221 (N_34221,N_33197,N_33348);
nor U34222 (N_34222,N_33671,N_33639);
xor U34223 (N_34223,N_33457,N_33061);
and U34224 (N_34224,N_32219,N_32176);
and U34225 (N_34225,N_33316,N_33451);
nor U34226 (N_34226,N_32448,N_33550);
nor U34227 (N_34227,N_32171,N_32596);
xor U34228 (N_34228,N_33649,N_32912);
or U34229 (N_34229,N_32180,N_32820);
xnor U34230 (N_34230,N_33696,N_33887);
nand U34231 (N_34231,N_33373,N_33145);
or U34232 (N_34232,N_33299,N_33199);
or U34233 (N_34233,N_32408,N_32208);
and U34234 (N_34234,N_33245,N_33156);
nand U34235 (N_34235,N_32335,N_33842);
xnor U34236 (N_34236,N_33937,N_33860);
and U34237 (N_34237,N_32214,N_33964);
xnor U34238 (N_34238,N_32284,N_33044);
and U34239 (N_34239,N_32594,N_33629);
or U34240 (N_34240,N_32896,N_33648);
and U34241 (N_34241,N_33033,N_33483);
nand U34242 (N_34242,N_33914,N_33473);
nor U34243 (N_34243,N_32498,N_32291);
nand U34244 (N_34244,N_33396,N_32028);
xnor U34245 (N_34245,N_33184,N_33700);
nand U34246 (N_34246,N_33129,N_32576);
xnor U34247 (N_34247,N_33651,N_32625);
nand U34248 (N_34248,N_32557,N_33264);
nor U34249 (N_34249,N_33722,N_33820);
and U34250 (N_34250,N_32049,N_32895);
nor U34251 (N_34251,N_33926,N_33813);
or U34252 (N_34252,N_32807,N_32270);
and U34253 (N_34253,N_33622,N_33776);
xor U34254 (N_34254,N_33759,N_32160);
xor U34255 (N_34255,N_33803,N_33969);
and U34256 (N_34256,N_33315,N_32908);
nand U34257 (N_34257,N_32810,N_32626);
nand U34258 (N_34258,N_33987,N_32433);
nand U34259 (N_34259,N_33845,N_33829);
nand U34260 (N_34260,N_32140,N_33432);
and U34261 (N_34261,N_32711,N_32525);
xor U34262 (N_34262,N_33330,N_32985);
nor U34263 (N_34263,N_32977,N_33207);
xnor U34264 (N_34264,N_33017,N_33641);
xor U34265 (N_34265,N_32862,N_32158);
nor U34266 (N_34266,N_32897,N_33581);
xnor U34267 (N_34267,N_33802,N_32061);
or U34268 (N_34268,N_32365,N_32302);
xnor U34269 (N_34269,N_33851,N_33932);
xnor U34270 (N_34270,N_32542,N_33227);
nand U34271 (N_34271,N_32327,N_32984);
and U34272 (N_34272,N_33328,N_32008);
and U34273 (N_34273,N_32438,N_33379);
and U34274 (N_34274,N_32868,N_32051);
xor U34275 (N_34275,N_33440,N_33196);
nand U34276 (N_34276,N_33371,N_32870);
or U34277 (N_34277,N_32507,N_32287);
and U34278 (N_34278,N_32121,N_32534);
and U34279 (N_34279,N_33124,N_33707);
nand U34280 (N_34280,N_33441,N_32506);
nand U34281 (N_34281,N_32315,N_32678);
or U34282 (N_34282,N_32255,N_32934);
nand U34283 (N_34283,N_33994,N_32037);
nand U34284 (N_34284,N_32353,N_32100);
xnor U34285 (N_34285,N_33867,N_33429);
and U34286 (N_34286,N_32865,N_32495);
and U34287 (N_34287,N_33486,N_32970);
nor U34288 (N_34288,N_32029,N_32355);
xor U34289 (N_34289,N_33357,N_33130);
nor U34290 (N_34290,N_32153,N_33431);
nand U34291 (N_34291,N_32730,N_33048);
nand U34292 (N_34292,N_32693,N_32662);
nor U34293 (N_34293,N_33818,N_32972);
xnor U34294 (N_34294,N_32437,N_32932);
or U34295 (N_34295,N_32484,N_33614);
nor U34296 (N_34296,N_33990,N_32244);
nor U34297 (N_34297,N_33688,N_33478);
or U34298 (N_34298,N_33665,N_33285);
nor U34299 (N_34299,N_32658,N_33816);
and U34300 (N_34300,N_33122,N_33815);
nor U34301 (N_34301,N_32567,N_33365);
nor U34302 (N_34302,N_33664,N_33388);
and U34303 (N_34303,N_33902,N_33387);
nand U34304 (N_34304,N_32925,N_32828);
nand U34305 (N_34305,N_32128,N_33472);
nand U34306 (N_34306,N_32541,N_33452);
nor U34307 (N_34307,N_33390,N_33185);
and U34308 (N_34308,N_32462,N_32098);
or U34309 (N_34309,N_33292,N_33039);
nor U34310 (N_34310,N_33137,N_32322);
and U34311 (N_34311,N_33374,N_32141);
and U34312 (N_34312,N_32529,N_32818);
and U34313 (N_34313,N_33494,N_33078);
nor U34314 (N_34314,N_33736,N_32743);
xor U34315 (N_34315,N_33907,N_32366);
nor U34316 (N_34316,N_33525,N_32712);
and U34317 (N_34317,N_33854,N_33928);
and U34318 (N_34318,N_32783,N_33888);
or U34319 (N_34319,N_33411,N_33324);
xnor U34320 (N_34320,N_32521,N_33336);
nor U34321 (N_34321,N_33024,N_33552);
or U34322 (N_34322,N_32152,N_32122);
nor U34323 (N_34323,N_33855,N_32548);
xor U34324 (N_34324,N_32349,N_33208);
nor U34325 (N_34325,N_33248,N_32069);
or U34326 (N_34326,N_33045,N_33623);
and U34327 (N_34327,N_33086,N_32587);
xor U34328 (N_34328,N_32022,N_33603);
and U34329 (N_34329,N_33012,N_33959);
or U34330 (N_34330,N_32621,N_32699);
or U34331 (N_34331,N_32585,N_32848);
nand U34332 (N_34332,N_33612,N_32346);
nand U34333 (N_34333,N_32919,N_32375);
nor U34334 (N_34334,N_32961,N_32457);
xor U34335 (N_34335,N_32860,N_32559);
or U34336 (N_34336,N_32817,N_32508);
nor U34337 (N_34337,N_32436,N_33598);
nand U34338 (N_34338,N_33311,N_32979);
and U34339 (N_34339,N_33458,N_32427);
nor U34340 (N_34340,N_32756,N_33068);
xor U34341 (N_34341,N_32130,N_33426);
nor U34342 (N_34342,N_33110,N_32224);
or U34343 (N_34343,N_33724,N_32851);
and U34344 (N_34344,N_32852,N_33150);
and U34345 (N_34345,N_33825,N_32641);
or U34346 (N_34346,N_32796,N_33031);
nor U34347 (N_34347,N_32101,N_33970);
or U34348 (N_34348,N_33703,N_32799);
xnor U34349 (N_34349,N_33446,N_33117);
nor U34350 (N_34350,N_33875,N_33289);
xor U34351 (N_34351,N_32572,N_33659);
and U34352 (N_34352,N_32210,N_32899);
and U34353 (N_34353,N_33609,N_32707);
and U34354 (N_34354,N_32188,N_33296);
xor U34355 (N_34355,N_32826,N_32450);
or U34356 (N_34356,N_33879,N_33701);
and U34357 (N_34357,N_33850,N_33011);
or U34358 (N_34358,N_33146,N_32727);
nor U34359 (N_34359,N_32885,N_32764);
and U34360 (N_34360,N_32443,N_33097);
xor U34361 (N_34361,N_33053,N_32946);
nor U34362 (N_34362,N_32422,N_32413);
nor U34363 (N_34363,N_32706,N_33253);
or U34364 (N_34364,N_32200,N_33869);
nand U34365 (N_34365,N_32729,N_32689);
nand U34366 (N_34366,N_32220,N_32502);
nor U34367 (N_34367,N_33338,N_33929);
nor U34368 (N_34368,N_32949,N_33433);
and U34369 (N_34369,N_32063,N_32139);
xnor U34370 (N_34370,N_33256,N_32263);
nor U34371 (N_34371,N_32285,N_33363);
nor U34372 (N_34372,N_33025,N_33051);
nand U34373 (N_34373,N_32277,N_33258);
nor U34374 (N_34374,N_33203,N_33018);
and U34375 (N_34375,N_33528,N_32923);
xor U34376 (N_34376,N_33587,N_32994);
nor U34377 (N_34377,N_33615,N_33500);
nand U34378 (N_34378,N_32425,N_33038);
nand U34379 (N_34379,N_32113,N_33950);
nand U34380 (N_34380,N_33754,N_32661);
nor U34381 (N_34381,N_32609,N_33627);
and U34382 (N_34382,N_32941,N_33490);
nor U34383 (N_34383,N_33133,N_32650);
nand U34384 (N_34384,N_32814,N_33134);
xor U34385 (N_34385,N_32054,N_33931);
nand U34386 (N_34386,N_32550,N_33728);
xnor U34387 (N_34387,N_32248,N_32876);
or U34388 (N_34388,N_33437,N_33104);
and U34389 (N_34389,N_32038,N_32524);
nor U34390 (N_34390,N_32074,N_33171);
or U34391 (N_34391,N_32701,N_32613);
xor U34392 (N_34392,N_32581,N_33840);
or U34393 (N_34393,N_32418,N_32268);
xor U34394 (N_34394,N_33636,N_32081);
or U34395 (N_34395,N_32036,N_33940);
or U34396 (N_34396,N_33985,N_33775);
or U34397 (N_34397,N_32488,N_32047);
xnor U34398 (N_34398,N_33154,N_33407);
nor U34399 (N_34399,N_32802,N_32386);
xor U34400 (N_34400,N_32884,N_33376);
or U34401 (N_34401,N_33617,N_33702);
or U34402 (N_34402,N_33434,N_33128);
nor U34403 (N_34403,N_33957,N_32376);
or U34404 (N_34404,N_32512,N_33569);
nand U34405 (N_34405,N_33774,N_32736);
or U34406 (N_34406,N_33463,N_32033);
or U34407 (N_34407,N_32866,N_33091);
and U34408 (N_34408,N_33276,N_33572);
xor U34409 (N_34409,N_32013,N_33389);
xnor U34410 (N_34410,N_32602,N_32354);
nand U34411 (N_34411,N_32195,N_32039);
nand U34412 (N_34412,N_32527,N_33354);
or U34413 (N_34413,N_33958,N_33766);
nand U34414 (N_34414,N_32936,N_32112);
nor U34415 (N_34415,N_32959,N_32075);
and U34416 (N_34416,N_33594,N_32070);
nand U34417 (N_34417,N_33394,N_33859);
or U34418 (N_34418,N_32722,N_33611);
xor U34419 (N_34419,N_33255,N_32404);
and U34420 (N_34420,N_33533,N_32903);
and U34421 (N_34421,N_32326,N_33861);
nor U34422 (N_34422,N_32239,N_32215);
nor U34423 (N_34423,N_32423,N_32250);
or U34424 (N_34424,N_33055,N_33894);
or U34425 (N_34425,N_32181,N_32643);
nor U34426 (N_34426,N_33647,N_32138);
and U34427 (N_34427,N_32083,N_33467);
or U34428 (N_34428,N_32831,N_32275);
xor U34429 (N_34429,N_33010,N_32698);
and U34430 (N_34430,N_33229,N_33919);
or U34431 (N_34431,N_32593,N_33356);
nor U34432 (N_34432,N_33404,N_33482);
nor U34433 (N_34433,N_33542,N_33637);
nand U34434 (N_34434,N_32445,N_33941);
nand U34435 (N_34435,N_32104,N_32668);
and U34436 (N_34436,N_32119,N_33908);
nand U34437 (N_34437,N_33224,N_33995);
or U34438 (N_34438,N_32742,N_33730);
nand U34439 (N_34439,N_32918,N_33795);
nor U34440 (N_34440,N_33006,N_33819);
nor U34441 (N_34441,N_32755,N_32242);
or U34442 (N_34442,N_32509,N_32775);
or U34443 (N_34443,N_32522,N_32716);
nand U34444 (N_34444,N_33507,N_32702);
or U34445 (N_34445,N_32888,N_33727);
nand U34446 (N_34446,N_32077,N_33096);
nor U34447 (N_34447,N_32050,N_32293);
xor U34448 (N_34448,N_33241,N_33335);
xor U34449 (N_34449,N_32580,N_33418);
and U34450 (N_34450,N_32440,N_32393);
or U34451 (N_34451,N_32691,N_33903);
or U34452 (N_34452,N_32948,N_32021);
or U34453 (N_34453,N_33408,N_32308);
nor U34454 (N_34454,N_33955,N_33050);
and U34455 (N_34455,N_32117,N_32257);
nand U34456 (N_34456,N_33259,N_32499);
or U34457 (N_34457,N_32165,N_33307);
nor U34458 (N_34458,N_33409,N_33901);
nor U34459 (N_34459,N_32084,N_33989);
and U34460 (N_34460,N_32012,N_33847);
nor U34461 (N_34461,N_33635,N_32636);
nand U34462 (N_34462,N_32385,N_33327);
xor U34463 (N_34463,N_32490,N_33566);
nand U34464 (N_34464,N_33741,N_32487);
nand U34465 (N_34465,N_33527,N_33571);
nor U34466 (N_34466,N_33880,N_32630);
and U34467 (N_34467,N_33239,N_33415);
nand U34468 (N_34468,N_33529,N_33905);
xnor U34469 (N_34469,N_32805,N_32312);
nor U34470 (N_34470,N_33518,N_32186);
or U34471 (N_34471,N_33821,N_32955);
xor U34472 (N_34472,N_33274,N_33760);
nand U34473 (N_34473,N_33747,N_33377);
nand U34474 (N_34474,N_33169,N_32872);
xnor U34475 (N_34475,N_33801,N_32001);
nand U34476 (N_34476,N_33746,N_33923);
or U34477 (N_34477,N_32125,N_32516);
xor U34478 (N_34478,N_32763,N_32497);
and U34479 (N_34479,N_33195,N_32218);
and U34480 (N_34480,N_33368,N_32654);
nand U34481 (N_34481,N_32095,N_33666);
xor U34482 (N_34482,N_32403,N_33205);
or U34483 (N_34483,N_33504,N_33098);
or U34484 (N_34484,N_32980,N_33948);
xnor U34485 (N_34485,N_33574,N_33346);
or U34486 (N_34486,N_33088,N_32780);
or U34487 (N_34487,N_33270,N_33771);
and U34488 (N_34488,N_33982,N_33545);
xnor U34489 (N_34489,N_32079,N_33251);
nand U34490 (N_34490,N_32733,N_33273);
xor U34491 (N_34491,N_33553,N_32543);
and U34492 (N_34492,N_32611,N_32471);
nand U34493 (N_34493,N_33886,N_32340);
and U34494 (N_34494,N_33805,N_32696);
and U34495 (N_34495,N_33716,N_33263);
and U34496 (N_34496,N_32635,N_32670);
and U34497 (N_34497,N_33706,N_32836);
nand U34498 (N_34498,N_32523,N_33502);
and U34499 (N_34499,N_32314,N_32292);
and U34500 (N_34500,N_33506,N_32720);
nor U34501 (N_34501,N_32960,N_33744);
nand U34502 (N_34502,N_33447,N_33658);
nand U34503 (N_34503,N_32952,N_32451);
and U34504 (N_34504,N_33213,N_33159);
xnor U34505 (N_34505,N_32622,N_33836);
xor U34506 (N_34506,N_32459,N_33980);
or U34507 (N_34507,N_32320,N_32768);
nand U34508 (N_34508,N_32816,N_33306);
xnor U34509 (N_34509,N_32574,N_33708);
and U34510 (N_34510,N_33442,N_32265);
nor U34511 (N_34511,N_32930,N_33436);
nor U34512 (N_34512,N_33743,N_32494);
or U34513 (N_34513,N_32325,N_33403);
nand U34514 (N_34514,N_33699,N_33077);
or U34515 (N_34515,N_32823,N_32446);
and U34516 (N_34516,N_32377,N_33966);
or U34517 (N_34517,N_32294,N_33677);
nor U34518 (N_34518,N_33254,N_33810);
or U34519 (N_34519,N_33465,N_33385);
and U34520 (N_34520,N_33857,N_32067);
and U34521 (N_34521,N_32071,N_32956);
or U34522 (N_34522,N_32765,N_33909);
and U34523 (N_34523,N_32311,N_32380);
and U34524 (N_34524,N_33466,N_32410);
nor U34525 (N_34525,N_32570,N_32184);
xnor U34526 (N_34526,N_32144,N_32843);
or U34527 (N_34527,N_32290,N_33977);
nand U34528 (N_34528,N_32452,N_32769);
xor U34529 (N_34529,N_32859,N_33391);
nand U34530 (N_34530,N_32466,N_32411);
nor U34531 (N_34531,N_32519,N_32520);
nand U34532 (N_34532,N_32234,N_32922);
and U34533 (N_34533,N_32841,N_32834);
xnor U34534 (N_34534,N_33522,N_33628);
nand U34535 (N_34535,N_33067,N_32558);
and U34536 (N_34536,N_32211,N_32597);
and U34537 (N_34537,N_32914,N_32695);
xnor U34538 (N_34538,N_33003,N_32359);
nand U34539 (N_34539,N_32917,N_33470);
or U34540 (N_34540,N_32400,N_33380);
nand U34541 (N_34541,N_32118,N_33784);
nand U34542 (N_34542,N_33341,N_33005);
or U34543 (N_34543,N_33610,N_32120);
nand U34544 (N_34544,N_33332,N_32788);
or U34545 (N_34545,N_32041,N_33974);
nor U34546 (N_34546,N_33520,N_33172);
or U34547 (N_34547,N_32342,N_32605);
or U34548 (N_34548,N_32847,N_32288);
nand U34549 (N_34549,N_32115,N_32191);
nor U34550 (N_34550,N_33539,N_33414);
xor U34551 (N_34551,N_33123,N_33720);
xor U34552 (N_34552,N_33488,N_32415);
or U34553 (N_34553,N_33644,N_33662);
and U34554 (N_34554,N_32639,N_33181);
and U34555 (N_34555,N_33935,N_32660);
or U34556 (N_34556,N_33999,N_32987);
nand U34557 (N_34557,N_33568,N_32849);
nor U34558 (N_34558,N_32228,N_32782);
nand U34559 (N_34559,N_32222,N_33495);
nor U34560 (N_34560,N_33459,N_32857);
and U34561 (N_34561,N_32439,N_33595);
and U34562 (N_34562,N_32205,N_32904);
and U34563 (N_34563,N_33884,N_32944);
xor U34564 (N_34564,N_33290,N_32924);
xnor U34565 (N_34565,N_33355,N_32677);
and U34566 (N_34566,N_33591,N_33262);
and U34567 (N_34567,N_32348,N_32486);
nor U34568 (N_34568,N_33075,N_32822);
and U34569 (N_34569,N_33120,N_32221);
xor U34570 (N_34570,N_32571,N_33427);
nor U34571 (N_34571,N_32926,N_33226);
nor U34572 (N_34572,N_33020,N_32811);
nor U34573 (N_34573,N_32825,N_33745);
nor U34574 (N_34574,N_33785,N_33733);
nor U34575 (N_34575,N_33834,N_33751);
and U34576 (N_34576,N_33930,N_32444);
nor U34577 (N_34577,N_33261,N_33893);
nor U34578 (N_34578,N_33456,N_32790);
or U34579 (N_34579,N_33375,N_33115);
nor U34580 (N_34580,N_33369,N_32094);
nand U34581 (N_34581,N_32056,N_33601);
nor U34582 (N_34582,N_33673,N_33755);
nand U34583 (N_34583,N_33549,N_32744);
xor U34584 (N_34584,N_33800,N_33342);
or U34585 (N_34585,N_33526,N_32198);
nor U34586 (N_34586,N_32940,N_33352);
nand U34587 (N_34587,N_33484,N_32324);
xor U34588 (N_34588,N_33849,N_33308);
and U34589 (N_34589,N_32240,N_32203);
nor U34590 (N_34590,N_32280,N_33735);
xor U34591 (N_34591,N_32953,N_32624);
nand U34592 (N_34592,N_33846,N_33606);
nor U34593 (N_34593,N_33517,N_33978);
xnor U34594 (N_34594,N_33624,N_32362);
and U34595 (N_34595,N_32771,N_32162);
nor U34596 (N_34596,N_32136,N_32126);
nor U34597 (N_34597,N_32080,N_32875);
xnor U34598 (N_34598,N_32207,N_33826);
nor U34599 (N_34599,N_33435,N_33157);
xnor U34600 (N_34600,N_33892,N_33358);
or U34601 (N_34601,N_32015,N_33885);
nor U34602 (N_34602,N_32204,N_32776);
and U34603 (N_34603,N_33638,N_33789);
or U34604 (N_34604,N_33960,N_32563);
and U34605 (N_34605,N_33113,N_32749);
xor U34606 (N_34606,N_32345,N_32642);
nand U34607 (N_34607,N_32674,N_33079);
or U34608 (N_34608,N_32978,N_32007);
and U34609 (N_34609,N_32421,N_33726);
or U34610 (N_34610,N_33142,N_33242);
xnor U34611 (N_34611,N_32910,N_32107);
nor U34612 (N_34612,N_32034,N_33642);
and U34613 (N_34613,N_33621,N_32441);
nor U34614 (N_34614,N_33419,N_33936);
or U34615 (N_34615,N_32059,N_33187);
nand U34616 (N_34616,N_33781,N_33344);
or U34617 (N_34617,N_32336,N_32785);
xor U34618 (N_34618,N_33757,N_33062);
xor U34619 (N_34619,N_33616,N_32901);
or U34620 (N_34620,N_32078,N_32323);
nand U34621 (N_34621,N_33439,N_33799);
xor U34622 (N_34622,N_32024,N_33946);
and U34623 (N_34623,N_33588,N_32131);
or U34624 (N_34624,N_32779,N_33350);
and U34625 (N_34625,N_32518,N_32089);
and U34626 (N_34626,N_33257,N_32458);
nor U34627 (N_34627,N_33103,N_32133);
nand U34628 (N_34628,N_33852,N_33711);
and U34629 (N_34629,N_32127,N_32645);
and U34630 (N_34630,N_32644,N_33562);
nand U34631 (N_34631,N_32772,N_33209);
nor U34632 (N_34632,N_33856,N_33511);
or U34633 (N_34633,N_33634,N_33681);
nor U34634 (N_34634,N_32943,N_32600);
nor U34635 (N_34635,N_32501,N_33837);
nor U34636 (N_34636,N_32588,N_33675);
xor U34637 (N_34637,N_33514,N_32728);
xnor U34638 (N_34638,N_33646,N_33471);
and U34639 (N_34639,N_32553,N_33996);
and U34640 (N_34640,N_33883,N_32991);
and U34641 (N_34641,N_33933,N_33054);
or U34642 (N_34642,N_33916,N_33992);
or U34643 (N_34643,N_32745,N_33464);
and U34644 (N_34644,N_33896,N_32361);
nand U34645 (N_34645,N_32407,N_32819);
and U34646 (N_34646,N_33943,N_32467);
and U34647 (N_34647,N_32233,N_32601);
nor U34648 (N_34648,N_33072,N_33787);
xnor U34649 (N_34649,N_32371,N_33945);
or U34650 (N_34650,N_32212,N_32504);
and U34651 (N_34651,N_32002,N_33178);
xnor U34652 (N_34652,N_32072,N_32019);
or U34653 (N_34653,N_33398,N_32786);
or U34654 (N_34654,N_33100,N_33049);
nand U34655 (N_34655,N_32388,N_33155);
xor U34656 (N_34656,N_33176,N_32442);
nor U34657 (N_34657,N_32417,N_32741);
or U34658 (N_34658,N_32245,N_32766);
nand U34659 (N_34659,N_32880,N_32829);
or U34660 (N_34660,N_32714,N_32262);
xnor U34661 (N_34661,N_32846,N_33597);
xor U34662 (N_34662,N_32777,N_33092);
nand U34663 (N_34663,N_32676,N_33536);
xnor U34664 (N_34664,N_33340,N_33756);
nor U34665 (N_34665,N_33772,N_32483);
or U34666 (N_34666,N_32725,N_32773);
nand U34667 (N_34667,N_33835,N_33180);
nor U34668 (N_34668,N_33070,N_32102);
and U34669 (N_34669,N_32296,N_33961);
or U34670 (N_34670,N_32513,N_32996);
or U34671 (N_34671,N_32740,N_33423);
and U34672 (N_34672,N_33921,N_32526);
nand U34673 (N_34673,N_32068,N_32480);
and U34674 (N_34674,N_32995,N_32907);
and U34675 (N_34675,N_33223,N_33600);
and U34676 (N_34676,N_33401,N_33037);
or U34677 (N_34677,N_32967,N_32966);
nor U34678 (N_34678,N_33559,N_33046);
nor U34679 (N_34679,N_32514,N_33204);
or U34680 (N_34680,N_32199,N_32185);
nand U34681 (N_34681,N_33593,N_33704);
and U34682 (N_34682,N_33809,N_33938);
or U34683 (N_34683,N_33535,N_33922);
nor U34684 (N_34684,N_33215,N_32159);
or U34685 (N_34685,N_32256,N_33384);
and U34686 (N_34686,N_33823,N_33870);
nor U34687 (N_34687,N_33531,N_33023);
nand U34688 (N_34688,N_33843,N_33848);
nor U34689 (N_34689,N_32360,N_33983);
nand U34690 (N_34690,N_33832,N_32616);
nand U34691 (N_34691,N_33895,N_32238);
xnor U34692 (N_34692,N_33939,N_32383);
and U34693 (N_34693,N_33106,N_32226);
or U34694 (N_34694,N_32206,N_32093);
nand U34695 (N_34695,N_32103,N_33694);
nor U34696 (N_34696,N_33167,N_33718);
and U34697 (N_34697,N_32850,N_32815);
or U34698 (N_34698,N_33173,N_33438);
and U34699 (N_34699,N_32812,N_33684);
xnor U34700 (N_34700,N_33313,N_33679);
xnor U34701 (N_34701,N_33882,N_32496);
nor U34702 (N_34702,N_33240,N_32861);
nor U34703 (N_34703,N_32964,N_32350);
and U34704 (N_34704,N_33360,N_32844);
nor U34705 (N_34705,N_32269,N_32304);
and U34706 (N_34706,N_33225,N_32503);
nand U34707 (N_34707,N_33004,N_32748);
or U34708 (N_34708,N_32564,N_33792);
nor U34709 (N_34709,N_32331,N_32878);
nand U34710 (N_34710,N_32974,N_33496);
and U34711 (N_34711,N_33965,N_32931);
nor U34712 (N_34712,N_33243,N_33059);
nor U34713 (N_34713,N_33445,N_32023);
xnor U34714 (N_34714,N_32663,N_33035);
xor U34715 (N_34715,N_33625,N_33238);
nand U34716 (N_34716,N_33219,N_33910);
and U34717 (N_34717,N_33475,N_33247);
and U34718 (N_34718,N_33105,N_33416);
or U34719 (N_34719,N_33986,N_32142);
xor U34720 (N_34720,N_33252,N_33318);
and U34721 (N_34721,N_33783,N_32795);
and U34722 (N_34722,N_33131,N_32992);
nor U34723 (N_34723,N_33029,N_32202);
nand U34724 (N_34724,N_32339,N_32813);
xor U34725 (N_34725,N_32057,N_32760);
or U34726 (N_34726,N_32737,N_33790);
nor U34727 (N_34727,N_33981,N_32690);
nand U34728 (N_34728,N_33116,N_32688);
xnor U34729 (N_34729,N_32235,N_33334);
nor U34730 (N_34730,N_33319,N_33177);
nor U34731 (N_34731,N_32489,N_32278);
xnor U34732 (N_34732,N_32470,N_32187);
or U34733 (N_34733,N_33322,N_33143);
or U34734 (N_34734,N_33667,N_32455);
xor U34735 (N_34735,N_32011,N_32531);
nand U34736 (N_34736,N_32610,N_33234);
nand U34737 (N_34737,N_32797,N_32808);
nor U34738 (N_34738,N_32612,N_32281);
or U34739 (N_34739,N_33063,N_33605);
and U34740 (N_34740,N_33118,N_33516);
and U34741 (N_34741,N_32517,N_32164);
nand U34742 (N_34742,N_32590,N_32189);
xor U34743 (N_34743,N_33589,N_33738);
and U34744 (N_34744,N_33312,N_32398);
or U34745 (N_34745,N_32409,N_33608);
or U34746 (N_34746,N_32491,N_32686);
and U34747 (N_34747,N_32088,N_32481);
or U34748 (N_34748,N_32957,N_32632);
nand U34749 (N_34749,N_32330,N_33216);
or U34750 (N_34750,N_32087,N_33381);
nor U34751 (N_34751,N_33294,N_33083);
or U34752 (N_34752,N_33565,N_32137);
nor U34753 (N_34753,N_32124,N_33112);
nand U34754 (N_34754,N_33763,N_32752);
nor U34755 (N_34755,N_33830,N_33286);
or U34756 (N_34756,N_33170,N_33047);
nand U34757 (N_34757,N_33383,N_32853);
nor U34758 (N_34758,N_32603,N_33304);
or U34759 (N_34759,N_32669,N_32565);
and U34760 (N_34760,N_32598,N_33499);
or U34761 (N_34761,N_32161,N_32592);
nand U34762 (N_34762,N_32097,N_33501);
nand U34763 (N_34763,N_33791,N_32482);
nor U34764 (N_34764,N_33927,N_32928);
or U34765 (N_34765,N_33393,N_33480);
xnor U34766 (N_34766,N_32845,N_32309);
and U34767 (N_34767,N_32578,N_32090);
xor U34768 (N_34768,N_33797,N_33161);
or U34769 (N_34769,N_33477,N_33602);
xnor U34770 (N_34770,N_33019,N_33523);
nor U34771 (N_34771,N_32151,N_32759);
xor U34772 (N_34772,N_33952,N_32929);
nand U34773 (N_34773,N_32246,N_33325);
nand U34774 (N_34774,N_33560,N_33201);
or U34775 (N_34775,N_32937,N_33561);
and U34776 (N_34776,N_32010,N_32619);
xor U34777 (N_34777,N_32252,N_33114);
or U34778 (N_34778,N_32259,N_32282);
xnor U34779 (N_34779,N_32942,N_32329);
nor U34780 (N_34780,N_32781,N_33217);
or U34781 (N_34781,N_32196,N_32738);
or U34782 (N_34782,N_33320,N_33548);
nor U34783 (N_34783,N_32430,N_32301);
or U34784 (N_34784,N_32492,N_32276);
nand U34785 (N_34785,N_32753,N_33043);
nor U34786 (N_34786,N_33685,N_32798);
nand U34787 (N_34787,N_32631,N_32344);
xnor U34788 (N_34788,N_33119,N_32073);
xor U34789 (N_34789,N_32363,N_32005);
xnor U34790 (N_34790,N_33163,N_32307);
nand U34791 (N_34791,N_33663,N_33302);
nand U34792 (N_34792,N_32016,N_32261);
xnor U34793 (N_34793,N_33297,N_33640);
nor U34794 (N_34794,N_32279,N_32260);
or U34795 (N_34795,N_33424,N_32993);
xnor U34796 (N_34796,N_33620,N_33954);
nor U34797 (N_34797,N_33052,N_32146);
or U34798 (N_34798,N_33406,N_32692);
nor U34799 (N_34799,N_33770,N_32735);
and U34800 (N_34800,N_33975,N_33630);
nand U34801 (N_34801,N_33399,N_32886);
and U34802 (N_34802,N_33281,N_32017);
xnor U34803 (N_34803,N_32584,N_33094);
nand U34804 (N_34804,N_32283,N_33814);
nor U34805 (N_34805,N_33269,N_32384);
and U34806 (N_34806,N_32132,N_33397);
xnor U34807 (N_34807,N_33866,N_32739);
nand U34808 (N_34808,N_32474,N_33151);
nor U34809 (N_34809,N_33474,N_32305);
and U34810 (N_34810,N_32109,N_33210);
nand U34811 (N_34811,N_33998,N_33911);
or U34812 (N_34812,N_33022,N_32869);
and U34813 (N_34813,N_32447,N_33503);
nor U34814 (N_34814,N_32065,N_32569);
or U34815 (N_34815,N_32156,N_32134);
nor U34816 (N_34816,N_33266,N_33833);
or U34817 (N_34817,N_32653,N_32681);
xnor U34818 (N_34818,N_32530,N_33206);
and U34819 (N_34819,N_32299,N_33697);
nand U34820 (N_34820,N_32175,N_33323);
nor U34821 (N_34821,N_33725,N_33395);
and U34822 (N_34822,N_33282,N_32839);
nor U34823 (N_34823,N_32297,N_32110);
xor U34824 (N_34824,N_32420,N_32963);
xor U34825 (N_34825,N_32709,N_33222);
nor U34826 (N_34826,N_33028,N_33582);
xnor U34827 (N_34827,N_33400,N_33182);
nor U34828 (N_34828,N_33073,N_32945);
and U34829 (N_34829,N_32538,N_32392);
xor U34830 (N_34830,N_33164,N_33000);
or U34831 (N_34831,N_32289,N_33920);
and U34832 (N_34832,N_32672,N_33326);
or U34833 (N_34833,N_32855,N_33807);
nand U34834 (N_34834,N_33881,N_33817);
and U34835 (N_34835,N_32835,N_32154);
nor U34836 (N_34836,N_32472,N_32705);
or U34837 (N_34837,N_33101,N_32762);
and U34838 (N_34838,N_33812,N_33705);
and U34839 (N_34839,N_33827,N_32731);
xnor U34840 (N_34840,N_32511,N_32981);
or U34841 (N_34841,N_32968,N_33359);
or U34842 (N_34842,N_33765,N_32951);
nor U34843 (N_34843,N_32310,N_32114);
xor U34844 (N_34844,N_32247,N_33287);
and U34845 (N_34845,N_33351,N_33822);
nor U34846 (N_34846,N_32715,N_32456);
and U34847 (N_34847,N_32833,N_33613);
xnor U34848 (N_34848,N_32973,N_33750);
or U34849 (N_34849,N_32241,N_32965);
xor U34850 (N_34850,N_33448,N_32044);
xnor U34851 (N_34851,N_32830,N_33579);
and U34852 (N_34852,N_33873,N_32982);
nand U34853 (N_34853,N_32734,N_33645);
and U34854 (N_34854,N_33027,N_33793);
or U34855 (N_34855,N_32387,N_33152);
and U34856 (N_34856,N_32382,N_32537);
nand U34857 (N_34857,N_32671,N_32434);
and U34858 (N_34858,N_33686,N_33449);
nand U34859 (N_34859,N_32535,N_33065);
nor U34860 (N_34860,N_32648,N_33190);
or U34861 (N_34861,N_33469,N_33853);
and U34862 (N_34862,N_32890,N_32806);
xnor U34863 (N_34863,N_32227,N_32232);
nor U34864 (N_34864,N_32976,N_32629);
nand U34865 (N_34865,N_33512,N_32236);
and U34866 (N_34866,N_33382,N_33898);
or U34867 (N_34867,N_32076,N_33071);
and U34868 (N_34868,N_33498,N_32147);
and U34869 (N_34869,N_33492,N_33798);
and U34870 (N_34870,N_33779,N_33405);
nand U34871 (N_34871,N_33714,N_33674);
nor U34872 (N_34872,N_33505,N_32554);
and U34873 (N_34873,N_32431,N_33844);
nor U34874 (N_34874,N_32091,N_32223);
and U34875 (N_34875,N_32651,N_32468);
or U34876 (N_34876,N_33158,N_32004);
nand U34877 (N_34877,N_33777,N_33392);
nor U34878 (N_34878,N_32477,N_33721);
or U34879 (N_34879,N_33547,N_33657);
or U34880 (N_34880,N_32338,N_33069);
nor U34881 (N_34881,N_33212,N_33193);
xnor U34882 (N_34882,N_32381,N_33557);
nor U34883 (N_34883,N_32390,N_33009);
nand U34884 (N_34884,N_32432,N_33014);
nand U34885 (N_34885,N_32920,N_32026);
nor U34886 (N_34886,N_32774,N_32167);
xor U34887 (N_34887,N_32416,N_33144);
xnor U34888 (N_34888,N_32229,N_33361);
xnor U34889 (N_34889,N_32837,N_33586);
nand U34890 (N_34890,N_32544,N_32751);
or U34891 (N_34891,N_32515,N_33546);
nand U34892 (N_34892,N_32682,N_32801);
and U34893 (N_34893,N_33174,N_32253);
nor U34894 (N_34894,N_32827,N_33683);
xor U34895 (N_34895,N_32652,N_33231);
nor U34896 (N_34896,N_32573,N_32761);
and U34897 (N_34897,N_33041,N_33080);
and U34898 (N_34898,N_33364,N_32412);
xnor U34899 (N_34899,N_32066,N_33951);
and U34900 (N_34900,N_33042,N_32724);
xor U34901 (N_34901,N_33218,N_32461);
and U34902 (N_34902,N_33246,N_33540);
or U34903 (N_34903,N_32397,N_32863);
xor U34904 (N_34904,N_33567,N_33712);
and U34905 (N_34905,N_33890,N_33592);
nor U34906 (N_34906,N_32249,N_33345);
and U34907 (N_34907,N_33093,N_32027);
nand U34908 (N_34908,N_33942,N_32675);
xnor U34909 (N_34909,N_33554,N_32789);
or U34910 (N_34910,N_33198,N_33422);
nor U34911 (N_34911,N_32062,N_33734);
xor U34912 (N_34912,N_32754,N_32402);
or U34913 (N_34913,N_33530,N_32793);
nor U34914 (N_34914,N_32374,N_33672);
nand U34915 (N_34915,N_33057,N_33081);
nor U34916 (N_34916,N_32906,N_32169);
and U34917 (N_34917,N_32364,N_33064);
nand U34918 (N_34918,N_33026,N_32902);
xnor U34919 (N_34919,N_33413,N_33497);
and U34920 (N_34920,N_32568,N_32989);
xor U34921 (N_34921,N_33372,N_33179);
nor U34922 (N_34922,N_32659,N_33656);
and U34923 (N_34923,N_33034,N_33347);
nand U34924 (N_34924,N_32649,N_33841);
or U34925 (N_34925,N_33758,N_33576);
xor U34926 (N_34926,N_33443,N_32463);
nand U34927 (N_34927,N_33538,N_32889);
nor U34928 (N_34928,N_32006,N_33633);
or U34929 (N_34929,N_32647,N_33183);
nand U34930 (N_34930,N_32615,N_32933);
or U34931 (N_34931,N_33515,N_32230);
nor U34932 (N_34932,N_33454,N_33563);
nand U34933 (N_34933,N_33668,N_32018);
or U34934 (N_34934,N_32628,N_32655);
nor U34935 (N_34935,N_33410,N_33421);
or U34936 (N_34936,N_33460,N_32251);
xor U34937 (N_34937,N_32273,N_33090);
or U34938 (N_34938,N_33655,N_32887);
and U34939 (N_34939,N_33739,N_33036);
and U34940 (N_34940,N_33991,N_33915);
xnor U34941 (N_34941,N_32401,N_32192);
nand U34942 (N_34942,N_32747,N_32064);
nand U34943 (N_34943,N_32473,N_33056);
nor U34944 (N_34944,N_32046,N_32163);
nor U34945 (N_34945,N_33740,N_33450);
xnor U34946 (N_34946,N_33737,N_33149);
and U34947 (N_34947,N_32607,N_32328);
xor U34948 (N_34948,N_33947,N_33295);
or U34949 (N_34949,N_32791,N_32873);
nor U34950 (N_34950,N_32800,N_33228);
xor U34951 (N_34951,N_32803,N_33508);
and U34952 (N_34952,N_32684,N_33192);
nand U34953 (N_34953,N_33211,N_32536);
and U34954 (N_34954,N_32148,N_33279);
or U34955 (N_34955,N_32020,N_32485);
nor U34956 (N_34956,N_32505,N_32337);
or U34957 (N_34957,N_33917,N_33773);
or U34958 (N_34958,N_32414,N_33191);
or U34959 (N_34959,N_32009,N_32157);
nand U34960 (N_34960,N_32710,N_32916);
nor U34961 (N_34961,N_33709,N_33425);
or U34962 (N_34962,N_33865,N_33271);
xor U34963 (N_34963,N_32938,N_33140);
nor U34964 (N_34964,N_32129,N_32680);
xnor U34965 (N_34965,N_33040,N_33912);
or U34966 (N_34966,N_32858,N_33462);
and U34967 (N_34967,N_33278,N_32640);
or U34968 (N_34968,N_33468,N_32478);
nand U34969 (N_34969,N_33769,N_32435);
xor U34970 (N_34970,N_33669,N_33220);
and U34971 (N_34971,N_33575,N_32209);
xor U34972 (N_34972,N_32770,N_33897);
or U34973 (N_34973,N_32334,N_32656);
and U34974 (N_34974,N_32767,N_33782);
nor U34975 (N_34975,N_32604,N_32351);
nor U34976 (N_34976,N_32510,N_32778);
xor U34977 (N_34977,N_33862,N_32877);
xor U34978 (N_34978,N_33653,N_32396);
and U34979 (N_34979,N_32357,N_32106);
and U34980 (N_34980,N_32172,N_32405);
nand U34981 (N_34981,N_32809,N_33979);
or U34982 (N_34982,N_32721,N_33366);
or U34983 (N_34983,N_33778,N_33838);
xnor U34984 (N_34984,N_32225,N_32116);
and U34985 (N_34985,N_32031,N_33794);
or U34986 (N_34986,N_32286,N_32694);
and U34987 (N_34987,N_32883,N_32358);
nor U34988 (N_34988,N_33692,N_32703);
nand U34989 (N_34989,N_33362,N_32892);
and U34990 (N_34990,N_33768,N_32988);
nor U34991 (N_34991,N_32254,N_32700);
xor U34992 (N_34992,N_33089,N_32395);
nor U34993 (N_34993,N_33678,N_33349);
xor U34994 (N_34994,N_32614,N_33732);
nand U34995 (N_34995,N_33551,N_33298);
xnor U34996 (N_34996,N_32540,N_32370);
nand U34997 (N_34997,N_33924,N_32893);
nor U34998 (N_34998,N_33698,N_33544);
and U34999 (N_34999,N_32168,N_33126);
nand U35000 (N_35000,N_33013,N_33416);
nand U35001 (N_35001,N_32327,N_32541);
or U35002 (N_35002,N_33924,N_33848);
nor U35003 (N_35003,N_32679,N_33876);
xor U35004 (N_35004,N_32981,N_33497);
nor U35005 (N_35005,N_33963,N_32527);
nor U35006 (N_35006,N_33541,N_33542);
or U35007 (N_35007,N_33279,N_32255);
or U35008 (N_35008,N_32142,N_33912);
nor U35009 (N_35009,N_33923,N_33214);
and U35010 (N_35010,N_33683,N_33485);
or U35011 (N_35011,N_32026,N_32494);
or U35012 (N_35012,N_33591,N_33198);
nor U35013 (N_35013,N_32303,N_33380);
and U35014 (N_35014,N_32856,N_32804);
xor U35015 (N_35015,N_33784,N_33465);
xor U35016 (N_35016,N_33903,N_33932);
or U35017 (N_35017,N_32212,N_32491);
and U35018 (N_35018,N_33986,N_33319);
nor U35019 (N_35019,N_33633,N_32043);
nor U35020 (N_35020,N_32460,N_33688);
and U35021 (N_35021,N_33816,N_32823);
or U35022 (N_35022,N_33052,N_32935);
nor U35023 (N_35023,N_33357,N_32053);
nand U35024 (N_35024,N_33482,N_32807);
or U35025 (N_35025,N_32225,N_33636);
nor U35026 (N_35026,N_32368,N_33734);
nor U35027 (N_35027,N_33860,N_33805);
nor U35028 (N_35028,N_32710,N_32432);
or U35029 (N_35029,N_33292,N_32893);
nor U35030 (N_35030,N_33911,N_32195);
nand U35031 (N_35031,N_33256,N_32705);
xnor U35032 (N_35032,N_33466,N_33770);
and U35033 (N_35033,N_32245,N_33320);
and U35034 (N_35034,N_32555,N_32501);
and U35035 (N_35035,N_32698,N_33580);
and U35036 (N_35036,N_32812,N_32661);
nand U35037 (N_35037,N_33426,N_33273);
or U35038 (N_35038,N_32745,N_33748);
and U35039 (N_35039,N_32395,N_33943);
xor U35040 (N_35040,N_33999,N_33640);
or U35041 (N_35041,N_33378,N_32268);
xor U35042 (N_35042,N_33468,N_33236);
and U35043 (N_35043,N_32647,N_33993);
nand U35044 (N_35044,N_32663,N_32108);
or U35045 (N_35045,N_33258,N_33328);
xnor U35046 (N_35046,N_32261,N_32444);
nand U35047 (N_35047,N_33139,N_32269);
xnor U35048 (N_35048,N_33084,N_33498);
and U35049 (N_35049,N_33345,N_32688);
nor U35050 (N_35050,N_33733,N_32859);
and U35051 (N_35051,N_32085,N_33238);
and U35052 (N_35052,N_32732,N_32048);
nor U35053 (N_35053,N_33332,N_33626);
xnor U35054 (N_35054,N_33689,N_33602);
nor U35055 (N_35055,N_33514,N_33492);
and U35056 (N_35056,N_33100,N_33065);
or U35057 (N_35057,N_32157,N_32469);
xor U35058 (N_35058,N_33757,N_32656);
and U35059 (N_35059,N_32588,N_33791);
xor U35060 (N_35060,N_32180,N_33927);
and U35061 (N_35061,N_32189,N_33346);
xnor U35062 (N_35062,N_33496,N_33781);
xor U35063 (N_35063,N_33031,N_32579);
and U35064 (N_35064,N_33886,N_33802);
nor U35065 (N_35065,N_33771,N_32718);
and U35066 (N_35066,N_32370,N_32899);
nor U35067 (N_35067,N_32084,N_33203);
xor U35068 (N_35068,N_32440,N_32439);
xnor U35069 (N_35069,N_32094,N_32146);
nor U35070 (N_35070,N_32046,N_32054);
or U35071 (N_35071,N_32775,N_33463);
nand U35072 (N_35072,N_32813,N_33993);
xnor U35073 (N_35073,N_32922,N_32830);
or U35074 (N_35074,N_32306,N_33415);
and U35075 (N_35075,N_32641,N_33780);
or U35076 (N_35076,N_33629,N_32032);
or U35077 (N_35077,N_33711,N_33786);
and U35078 (N_35078,N_33631,N_33470);
and U35079 (N_35079,N_32281,N_33454);
and U35080 (N_35080,N_32032,N_32487);
nor U35081 (N_35081,N_32986,N_32397);
nand U35082 (N_35082,N_32502,N_33731);
nand U35083 (N_35083,N_33762,N_33595);
nand U35084 (N_35084,N_33295,N_32535);
nor U35085 (N_35085,N_32968,N_32999);
and U35086 (N_35086,N_32753,N_33080);
or U35087 (N_35087,N_33314,N_33558);
nand U35088 (N_35088,N_32353,N_33912);
xor U35089 (N_35089,N_33021,N_32283);
nor U35090 (N_35090,N_32694,N_32372);
nand U35091 (N_35091,N_33223,N_32538);
and U35092 (N_35092,N_32604,N_33815);
nor U35093 (N_35093,N_33029,N_33572);
nor U35094 (N_35094,N_32703,N_32602);
and U35095 (N_35095,N_32007,N_32220);
xor U35096 (N_35096,N_33314,N_33453);
nand U35097 (N_35097,N_32521,N_32349);
xnor U35098 (N_35098,N_32266,N_32903);
nand U35099 (N_35099,N_32914,N_32950);
or U35100 (N_35100,N_32530,N_33668);
nor U35101 (N_35101,N_32705,N_32234);
or U35102 (N_35102,N_33127,N_33436);
xor U35103 (N_35103,N_32415,N_32346);
xor U35104 (N_35104,N_32271,N_32242);
or U35105 (N_35105,N_32158,N_33860);
or U35106 (N_35106,N_33984,N_32195);
nand U35107 (N_35107,N_33532,N_33434);
nor U35108 (N_35108,N_32668,N_32144);
and U35109 (N_35109,N_32899,N_33521);
nor U35110 (N_35110,N_32829,N_32765);
nand U35111 (N_35111,N_33900,N_33202);
or U35112 (N_35112,N_33967,N_33016);
nor U35113 (N_35113,N_33248,N_33000);
nor U35114 (N_35114,N_33330,N_32992);
and U35115 (N_35115,N_32137,N_33787);
and U35116 (N_35116,N_32736,N_33035);
and U35117 (N_35117,N_32227,N_33959);
and U35118 (N_35118,N_33255,N_33931);
or U35119 (N_35119,N_32780,N_33744);
xor U35120 (N_35120,N_32035,N_32542);
nand U35121 (N_35121,N_32576,N_32883);
nand U35122 (N_35122,N_32894,N_33054);
nand U35123 (N_35123,N_32502,N_33323);
xor U35124 (N_35124,N_33299,N_32400);
and U35125 (N_35125,N_32353,N_33061);
or U35126 (N_35126,N_33141,N_32473);
nand U35127 (N_35127,N_32143,N_32211);
or U35128 (N_35128,N_32665,N_32044);
xnor U35129 (N_35129,N_32995,N_33259);
xnor U35130 (N_35130,N_33757,N_33673);
or U35131 (N_35131,N_33754,N_32611);
or U35132 (N_35132,N_33234,N_33103);
nand U35133 (N_35133,N_33272,N_33069);
nand U35134 (N_35134,N_33546,N_33218);
or U35135 (N_35135,N_33659,N_32427);
or U35136 (N_35136,N_32815,N_33714);
nand U35137 (N_35137,N_33723,N_33394);
nand U35138 (N_35138,N_32586,N_33965);
or U35139 (N_35139,N_32820,N_33805);
or U35140 (N_35140,N_33400,N_33944);
and U35141 (N_35141,N_33287,N_33464);
xor U35142 (N_35142,N_32787,N_32343);
xnor U35143 (N_35143,N_32012,N_32095);
nand U35144 (N_35144,N_32732,N_32559);
or U35145 (N_35145,N_33318,N_33988);
or U35146 (N_35146,N_33909,N_33133);
and U35147 (N_35147,N_33490,N_33302);
nor U35148 (N_35148,N_32317,N_33492);
xor U35149 (N_35149,N_33509,N_32527);
nand U35150 (N_35150,N_33901,N_32137);
nor U35151 (N_35151,N_33188,N_32348);
nor U35152 (N_35152,N_33306,N_33777);
nand U35153 (N_35153,N_32180,N_33268);
nor U35154 (N_35154,N_33331,N_32999);
and U35155 (N_35155,N_32214,N_32350);
xnor U35156 (N_35156,N_33929,N_33117);
or U35157 (N_35157,N_32810,N_33192);
or U35158 (N_35158,N_32936,N_32293);
nand U35159 (N_35159,N_33945,N_32494);
nand U35160 (N_35160,N_32592,N_33364);
or U35161 (N_35161,N_32629,N_33577);
nand U35162 (N_35162,N_32750,N_32030);
nor U35163 (N_35163,N_32957,N_33236);
nand U35164 (N_35164,N_33880,N_32045);
or U35165 (N_35165,N_32762,N_33179);
nor U35166 (N_35166,N_32966,N_32373);
nand U35167 (N_35167,N_32536,N_33426);
nor U35168 (N_35168,N_32080,N_32567);
nor U35169 (N_35169,N_33047,N_32851);
xnor U35170 (N_35170,N_32198,N_32717);
or U35171 (N_35171,N_33937,N_32136);
nor U35172 (N_35172,N_32412,N_32546);
and U35173 (N_35173,N_33138,N_33505);
nand U35174 (N_35174,N_33248,N_32453);
xor U35175 (N_35175,N_33988,N_32238);
xnor U35176 (N_35176,N_33569,N_32832);
or U35177 (N_35177,N_33932,N_33369);
nor U35178 (N_35178,N_32520,N_33552);
nor U35179 (N_35179,N_32754,N_33645);
or U35180 (N_35180,N_33578,N_33856);
nand U35181 (N_35181,N_33652,N_33407);
or U35182 (N_35182,N_32788,N_33355);
or U35183 (N_35183,N_32563,N_32666);
or U35184 (N_35184,N_32763,N_33784);
nor U35185 (N_35185,N_33013,N_33885);
or U35186 (N_35186,N_32446,N_32588);
and U35187 (N_35187,N_32034,N_33755);
nand U35188 (N_35188,N_32915,N_33396);
xor U35189 (N_35189,N_33547,N_32041);
xor U35190 (N_35190,N_32341,N_32178);
or U35191 (N_35191,N_32092,N_33772);
and U35192 (N_35192,N_33664,N_33630);
and U35193 (N_35193,N_33779,N_32503);
nand U35194 (N_35194,N_32822,N_33321);
nand U35195 (N_35195,N_32737,N_32575);
and U35196 (N_35196,N_32194,N_33789);
or U35197 (N_35197,N_33113,N_33833);
nor U35198 (N_35198,N_33111,N_32403);
xor U35199 (N_35199,N_33765,N_32922);
nand U35200 (N_35200,N_32278,N_33962);
nor U35201 (N_35201,N_32183,N_32341);
xnor U35202 (N_35202,N_33702,N_33283);
nor U35203 (N_35203,N_32144,N_32801);
xnor U35204 (N_35204,N_32645,N_33950);
xnor U35205 (N_35205,N_32606,N_33794);
nor U35206 (N_35206,N_32690,N_32101);
nand U35207 (N_35207,N_33211,N_32338);
and U35208 (N_35208,N_33346,N_33613);
nor U35209 (N_35209,N_33986,N_32325);
and U35210 (N_35210,N_32511,N_32712);
xor U35211 (N_35211,N_33770,N_33117);
nor U35212 (N_35212,N_32585,N_33461);
nand U35213 (N_35213,N_33974,N_32978);
nor U35214 (N_35214,N_33088,N_33806);
and U35215 (N_35215,N_32035,N_32618);
xnor U35216 (N_35216,N_33595,N_33887);
xor U35217 (N_35217,N_33649,N_33788);
nor U35218 (N_35218,N_33406,N_33905);
xor U35219 (N_35219,N_32451,N_33382);
nor U35220 (N_35220,N_33337,N_33125);
or U35221 (N_35221,N_33618,N_32697);
or U35222 (N_35222,N_32061,N_32666);
or U35223 (N_35223,N_33678,N_33895);
nand U35224 (N_35224,N_33353,N_33506);
nand U35225 (N_35225,N_33689,N_32628);
xnor U35226 (N_35226,N_33811,N_33529);
or U35227 (N_35227,N_33568,N_33033);
xnor U35228 (N_35228,N_33827,N_33600);
nor U35229 (N_35229,N_32250,N_32418);
nor U35230 (N_35230,N_32705,N_33160);
xnor U35231 (N_35231,N_33171,N_32217);
nand U35232 (N_35232,N_33918,N_33668);
and U35233 (N_35233,N_32318,N_33049);
xor U35234 (N_35234,N_32917,N_32008);
xor U35235 (N_35235,N_32270,N_32124);
xnor U35236 (N_35236,N_33588,N_33140);
xnor U35237 (N_35237,N_32324,N_32384);
nor U35238 (N_35238,N_32322,N_33845);
xnor U35239 (N_35239,N_33333,N_32314);
or U35240 (N_35240,N_32578,N_32537);
nand U35241 (N_35241,N_32960,N_32170);
nor U35242 (N_35242,N_33010,N_32080);
nand U35243 (N_35243,N_33515,N_32094);
xnor U35244 (N_35244,N_32904,N_32892);
nor U35245 (N_35245,N_33723,N_32276);
nor U35246 (N_35246,N_33389,N_32908);
xnor U35247 (N_35247,N_32995,N_33904);
and U35248 (N_35248,N_33635,N_32935);
nor U35249 (N_35249,N_32011,N_33524);
and U35250 (N_35250,N_33119,N_33028);
nor U35251 (N_35251,N_33609,N_32854);
nand U35252 (N_35252,N_33717,N_32590);
nor U35253 (N_35253,N_33481,N_32100);
and U35254 (N_35254,N_32163,N_32940);
and U35255 (N_35255,N_33195,N_33612);
nand U35256 (N_35256,N_32582,N_33023);
xor U35257 (N_35257,N_33094,N_32346);
xor U35258 (N_35258,N_33952,N_33006);
and U35259 (N_35259,N_33659,N_33743);
xnor U35260 (N_35260,N_32553,N_33521);
nor U35261 (N_35261,N_33016,N_33025);
or U35262 (N_35262,N_32353,N_32365);
xor U35263 (N_35263,N_33801,N_32463);
nor U35264 (N_35264,N_33071,N_32852);
nor U35265 (N_35265,N_33171,N_33126);
or U35266 (N_35266,N_32351,N_33160);
and U35267 (N_35267,N_32288,N_32240);
nor U35268 (N_35268,N_33811,N_33751);
xnor U35269 (N_35269,N_32143,N_33528);
and U35270 (N_35270,N_33956,N_32728);
xnor U35271 (N_35271,N_33852,N_32513);
nor U35272 (N_35272,N_33527,N_32366);
or U35273 (N_35273,N_33694,N_32366);
or U35274 (N_35274,N_32940,N_33669);
nand U35275 (N_35275,N_33618,N_33111);
or U35276 (N_35276,N_33686,N_32919);
xor U35277 (N_35277,N_33570,N_33068);
nand U35278 (N_35278,N_32275,N_33956);
or U35279 (N_35279,N_32774,N_32242);
and U35280 (N_35280,N_32786,N_32842);
and U35281 (N_35281,N_32853,N_33380);
nand U35282 (N_35282,N_32064,N_32878);
nor U35283 (N_35283,N_32342,N_32823);
nor U35284 (N_35284,N_32653,N_32889);
nand U35285 (N_35285,N_32248,N_32677);
and U35286 (N_35286,N_32757,N_33369);
or U35287 (N_35287,N_33093,N_32064);
or U35288 (N_35288,N_32179,N_32914);
or U35289 (N_35289,N_33861,N_33746);
and U35290 (N_35290,N_33723,N_32210);
or U35291 (N_35291,N_33303,N_33474);
and U35292 (N_35292,N_33869,N_32263);
xnor U35293 (N_35293,N_32088,N_33117);
or U35294 (N_35294,N_32518,N_32525);
xnor U35295 (N_35295,N_32928,N_33717);
and U35296 (N_35296,N_32137,N_33390);
xnor U35297 (N_35297,N_32072,N_33640);
nand U35298 (N_35298,N_32415,N_32635);
nand U35299 (N_35299,N_33554,N_33157);
or U35300 (N_35300,N_33106,N_32036);
or U35301 (N_35301,N_33350,N_33979);
nor U35302 (N_35302,N_32104,N_33884);
and U35303 (N_35303,N_32519,N_33829);
or U35304 (N_35304,N_33493,N_32116);
xnor U35305 (N_35305,N_33762,N_33056);
xor U35306 (N_35306,N_33182,N_33141);
or U35307 (N_35307,N_32574,N_33310);
xor U35308 (N_35308,N_32057,N_33283);
nor U35309 (N_35309,N_33684,N_33271);
and U35310 (N_35310,N_32605,N_33040);
nand U35311 (N_35311,N_33660,N_32102);
or U35312 (N_35312,N_32952,N_32813);
or U35313 (N_35313,N_33779,N_33392);
and U35314 (N_35314,N_32755,N_32008);
nand U35315 (N_35315,N_32724,N_32177);
xor U35316 (N_35316,N_33964,N_33955);
or U35317 (N_35317,N_33921,N_32226);
nor U35318 (N_35318,N_32009,N_33303);
nand U35319 (N_35319,N_33887,N_33578);
nor U35320 (N_35320,N_33353,N_32415);
or U35321 (N_35321,N_32397,N_32586);
nor U35322 (N_35322,N_32951,N_32357);
nor U35323 (N_35323,N_32703,N_32151);
and U35324 (N_35324,N_33473,N_32300);
nor U35325 (N_35325,N_33620,N_33140);
nand U35326 (N_35326,N_33538,N_32300);
or U35327 (N_35327,N_32502,N_33907);
xnor U35328 (N_35328,N_33245,N_33367);
or U35329 (N_35329,N_32695,N_32097);
nor U35330 (N_35330,N_32869,N_32157);
xor U35331 (N_35331,N_32858,N_32893);
and U35332 (N_35332,N_32969,N_32463);
xor U35333 (N_35333,N_32833,N_33337);
nor U35334 (N_35334,N_33750,N_33061);
nand U35335 (N_35335,N_32900,N_32244);
xor U35336 (N_35336,N_33794,N_32840);
nor U35337 (N_35337,N_33622,N_33186);
and U35338 (N_35338,N_32687,N_33289);
nand U35339 (N_35339,N_32229,N_33650);
and U35340 (N_35340,N_33230,N_33103);
nor U35341 (N_35341,N_32822,N_33028);
nand U35342 (N_35342,N_33541,N_33476);
or U35343 (N_35343,N_33049,N_32851);
nand U35344 (N_35344,N_33736,N_32658);
nand U35345 (N_35345,N_33426,N_32436);
nand U35346 (N_35346,N_33756,N_33277);
nor U35347 (N_35347,N_32191,N_32494);
xnor U35348 (N_35348,N_32670,N_32031);
nand U35349 (N_35349,N_32502,N_33557);
nand U35350 (N_35350,N_32260,N_32376);
nor U35351 (N_35351,N_32554,N_32856);
nor U35352 (N_35352,N_32154,N_33002);
nand U35353 (N_35353,N_33443,N_32777);
nand U35354 (N_35354,N_33118,N_32727);
nand U35355 (N_35355,N_32315,N_33881);
xor U35356 (N_35356,N_32831,N_32555);
and U35357 (N_35357,N_33061,N_33366);
and U35358 (N_35358,N_32464,N_32346);
or U35359 (N_35359,N_33268,N_32510);
nor U35360 (N_35360,N_32701,N_32776);
xor U35361 (N_35361,N_33825,N_33855);
or U35362 (N_35362,N_33953,N_33695);
nand U35363 (N_35363,N_33063,N_33856);
and U35364 (N_35364,N_33596,N_33695);
nand U35365 (N_35365,N_33503,N_33625);
nand U35366 (N_35366,N_32735,N_33923);
and U35367 (N_35367,N_32648,N_32102);
xor U35368 (N_35368,N_32778,N_33792);
and U35369 (N_35369,N_33096,N_32306);
and U35370 (N_35370,N_32547,N_32577);
xor U35371 (N_35371,N_32511,N_33979);
or U35372 (N_35372,N_33531,N_33640);
nand U35373 (N_35373,N_32592,N_32804);
nor U35374 (N_35374,N_32630,N_32751);
nor U35375 (N_35375,N_32963,N_33159);
nor U35376 (N_35376,N_33380,N_33763);
and U35377 (N_35377,N_33809,N_33433);
xor U35378 (N_35378,N_32020,N_32372);
or U35379 (N_35379,N_32356,N_32581);
or U35380 (N_35380,N_32826,N_32684);
nand U35381 (N_35381,N_33031,N_32041);
nand U35382 (N_35382,N_32554,N_33500);
and U35383 (N_35383,N_32893,N_33412);
nand U35384 (N_35384,N_33895,N_33169);
and U35385 (N_35385,N_33309,N_32850);
or U35386 (N_35386,N_33320,N_33078);
or U35387 (N_35387,N_33725,N_33256);
or U35388 (N_35388,N_33139,N_32952);
and U35389 (N_35389,N_33661,N_33507);
nor U35390 (N_35390,N_33841,N_33495);
and U35391 (N_35391,N_33806,N_32671);
nand U35392 (N_35392,N_33279,N_33205);
nand U35393 (N_35393,N_33470,N_33794);
and U35394 (N_35394,N_33708,N_32129);
nor U35395 (N_35395,N_32235,N_33035);
xor U35396 (N_35396,N_32389,N_33969);
or U35397 (N_35397,N_33161,N_33067);
nor U35398 (N_35398,N_33548,N_32596);
xnor U35399 (N_35399,N_33698,N_33953);
xnor U35400 (N_35400,N_33148,N_33267);
and U35401 (N_35401,N_33240,N_32469);
xnor U35402 (N_35402,N_32030,N_32339);
xnor U35403 (N_35403,N_33625,N_33867);
and U35404 (N_35404,N_33220,N_32581);
xor U35405 (N_35405,N_33338,N_33225);
nand U35406 (N_35406,N_33935,N_33964);
xnor U35407 (N_35407,N_33275,N_32583);
or U35408 (N_35408,N_33188,N_33635);
xnor U35409 (N_35409,N_33183,N_33875);
xor U35410 (N_35410,N_32032,N_33087);
nand U35411 (N_35411,N_33007,N_33317);
nor U35412 (N_35412,N_33177,N_33853);
nor U35413 (N_35413,N_32547,N_33623);
xnor U35414 (N_35414,N_33532,N_33935);
and U35415 (N_35415,N_33925,N_32521);
and U35416 (N_35416,N_33687,N_32252);
nor U35417 (N_35417,N_32615,N_33699);
xnor U35418 (N_35418,N_32065,N_32727);
and U35419 (N_35419,N_33846,N_32255);
or U35420 (N_35420,N_32961,N_32916);
nor U35421 (N_35421,N_32432,N_32427);
nor U35422 (N_35422,N_33927,N_32764);
nand U35423 (N_35423,N_32718,N_32646);
nand U35424 (N_35424,N_32252,N_32027);
and U35425 (N_35425,N_33167,N_32766);
or U35426 (N_35426,N_33394,N_33923);
nor U35427 (N_35427,N_33023,N_33803);
nand U35428 (N_35428,N_32996,N_32596);
nand U35429 (N_35429,N_32383,N_32641);
and U35430 (N_35430,N_32032,N_32235);
or U35431 (N_35431,N_33522,N_32081);
nor U35432 (N_35432,N_33608,N_33906);
and U35433 (N_35433,N_33239,N_32886);
and U35434 (N_35434,N_32686,N_32875);
xnor U35435 (N_35435,N_33080,N_32978);
or U35436 (N_35436,N_33449,N_32218);
nand U35437 (N_35437,N_33143,N_32583);
and U35438 (N_35438,N_32116,N_33880);
nor U35439 (N_35439,N_33765,N_32834);
nor U35440 (N_35440,N_33641,N_32514);
nor U35441 (N_35441,N_33995,N_32238);
nor U35442 (N_35442,N_32185,N_33502);
nor U35443 (N_35443,N_32158,N_33750);
and U35444 (N_35444,N_32793,N_33321);
nor U35445 (N_35445,N_33444,N_32475);
and U35446 (N_35446,N_33957,N_32501);
and U35447 (N_35447,N_32718,N_33951);
nand U35448 (N_35448,N_33683,N_32971);
or U35449 (N_35449,N_32653,N_33837);
or U35450 (N_35450,N_32774,N_33096);
xnor U35451 (N_35451,N_32152,N_33898);
and U35452 (N_35452,N_33602,N_32509);
xnor U35453 (N_35453,N_33062,N_33668);
or U35454 (N_35454,N_32631,N_32464);
nor U35455 (N_35455,N_33630,N_32699);
nand U35456 (N_35456,N_33497,N_33899);
and U35457 (N_35457,N_32260,N_33768);
nor U35458 (N_35458,N_33175,N_33560);
and U35459 (N_35459,N_32679,N_32900);
nand U35460 (N_35460,N_33001,N_32044);
xnor U35461 (N_35461,N_33990,N_32330);
nor U35462 (N_35462,N_33269,N_33724);
nand U35463 (N_35463,N_33148,N_33597);
nor U35464 (N_35464,N_33951,N_33527);
and U35465 (N_35465,N_33407,N_33243);
xor U35466 (N_35466,N_33041,N_33620);
nor U35467 (N_35467,N_33542,N_33729);
nor U35468 (N_35468,N_33039,N_33146);
nor U35469 (N_35469,N_33798,N_32734);
and U35470 (N_35470,N_32310,N_32308);
nand U35471 (N_35471,N_32566,N_33158);
and U35472 (N_35472,N_32716,N_32007);
and U35473 (N_35473,N_32684,N_33322);
xor U35474 (N_35474,N_32192,N_33991);
nor U35475 (N_35475,N_33752,N_33086);
nor U35476 (N_35476,N_32676,N_33748);
or U35477 (N_35477,N_32147,N_33032);
nand U35478 (N_35478,N_33103,N_32449);
nand U35479 (N_35479,N_32270,N_33193);
xnor U35480 (N_35480,N_33833,N_33467);
nor U35481 (N_35481,N_32395,N_33104);
and U35482 (N_35482,N_32842,N_33471);
nand U35483 (N_35483,N_33249,N_32119);
nand U35484 (N_35484,N_33681,N_32816);
nand U35485 (N_35485,N_32799,N_33612);
and U35486 (N_35486,N_32120,N_33795);
nor U35487 (N_35487,N_33854,N_32572);
xor U35488 (N_35488,N_32872,N_32926);
nand U35489 (N_35489,N_32211,N_32984);
nor U35490 (N_35490,N_33463,N_33799);
nand U35491 (N_35491,N_33205,N_32030);
nand U35492 (N_35492,N_33121,N_32139);
and U35493 (N_35493,N_32624,N_33660);
or U35494 (N_35494,N_33804,N_33012);
or U35495 (N_35495,N_33547,N_32017);
nand U35496 (N_35496,N_32593,N_33086);
or U35497 (N_35497,N_33851,N_33746);
and U35498 (N_35498,N_32785,N_33752);
xnor U35499 (N_35499,N_33550,N_33670);
xnor U35500 (N_35500,N_33070,N_33720);
and U35501 (N_35501,N_32771,N_33852);
xor U35502 (N_35502,N_33981,N_32250);
nor U35503 (N_35503,N_32073,N_33683);
nand U35504 (N_35504,N_33259,N_33963);
or U35505 (N_35505,N_32086,N_32006);
and U35506 (N_35506,N_33109,N_32045);
nand U35507 (N_35507,N_33806,N_32200);
and U35508 (N_35508,N_32576,N_33817);
nor U35509 (N_35509,N_33483,N_32830);
or U35510 (N_35510,N_33243,N_32525);
nor U35511 (N_35511,N_33173,N_32131);
or U35512 (N_35512,N_33250,N_32786);
nor U35513 (N_35513,N_32836,N_33745);
nand U35514 (N_35514,N_33719,N_32960);
nand U35515 (N_35515,N_33624,N_32889);
and U35516 (N_35516,N_33114,N_33922);
or U35517 (N_35517,N_33751,N_33020);
nand U35518 (N_35518,N_33546,N_32406);
or U35519 (N_35519,N_33795,N_32703);
nor U35520 (N_35520,N_32675,N_33813);
nor U35521 (N_35521,N_33649,N_33941);
and U35522 (N_35522,N_32879,N_33322);
xnor U35523 (N_35523,N_32552,N_33633);
xnor U35524 (N_35524,N_33606,N_32617);
or U35525 (N_35525,N_32145,N_33881);
or U35526 (N_35526,N_32663,N_32883);
and U35527 (N_35527,N_33416,N_32029);
xnor U35528 (N_35528,N_32295,N_32823);
or U35529 (N_35529,N_33655,N_32653);
and U35530 (N_35530,N_33458,N_33431);
or U35531 (N_35531,N_33359,N_32242);
and U35532 (N_35532,N_32377,N_32443);
nand U35533 (N_35533,N_32191,N_32359);
and U35534 (N_35534,N_33963,N_33595);
or U35535 (N_35535,N_32752,N_33663);
nand U35536 (N_35536,N_33421,N_32643);
or U35537 (N_35537,N_33600,N_32353);
and U35538 (N_35538,N_33798,N_32349);
or U35539 (N_35539,N_32327,N_32825);
or U35540 (N_35540,N_33681,N_33385);
nor U35541 (N_35541,N_32134,N_33701);
and U35542 (N_35542,N_33129,N_33187);
nor U35543 (N_35543,N_32143,N_32263);
nand U35544 (N_35544,N_33512,N_33418);
or U35545 (N_35545,N_32359,N_33348);
nor U35546 (N_35546,N_33973,N_33247);
and U35547 (N_35547,N_33232,N_32336);
nor U35548 (N_35548,N_32679,N_32515);
nand U35549 (N_35549,N_33210,N_32339);
or U35550 (N_35550,N_33735,N_33909);
nor U35551 (N_35551,N_32915,N_33779);
or U35552 (N_35552,N_33632,N_32703);
xor U35553 (N_35553,N_33537,N_32396);
or U35554 (N_35554,N_33398,N_32337);
or U35555 (N_35555,N_33580,N_32662);
nor U35556 (N_35556,N_33373,N_33363);
nor U35557 (N_35557,N_32430,N_33585);
nor U35558 (N_35558,N_33761,N_32534);
nor U35559 (N_35559,N_32688,N_32480);
or U35560 (N_35560,N_33941,N_33052);
nand U35561 (N_35561,N_33025,N_32522);
xnor U35562 (N_35562,N_32699,N_32244);
nand U35563 (N_35563,N_33350,N_32877);
and U35564 (N_35564,N_32434,N_32729);
and U35565 (N_35565,N_33342,N_33219);
or U35566 (N_35566,N_33816,N_32221);
and U35567 (N_35567,N_32642,N_32484);
nor U35568 (N_35568,N_32718,N_32811);
nor U35569 (N_35569,N_32286,N_33223);
and U35570 (N_35570,N_33142,N_32745);
or U35571 (N_35571,N_32384,N_33093);
nand U35572 (N_35572,N_33860,N_33892);
xnor U35573 (N_35573,N_32127,N_32797);
nand U35574 (N_35574,N_32750,N_33287);
or U35575 (N_35575,N_33993,N_33039);
or U35576 (N_35576,N_33712,N_32685);
nor U35577 (N_35577,N_33929,N_32242);
nand U35578 (N_35578,N_33519,N_32204);
nor U35579 (N_35579,N_33825,N_33018);
nor U35580 (N_35580,N_32593,N_33744);
nor U35581 (N_35581,N_33063,N_33793);
nand U35582 (N_35582,N_32408,N_32029);
nand U35583 (N_35583,N_33725,N_33114);
or U35584 (N_35584,N_33568,N_33588);
nand U35585 (N_35585,N_33370,N_32759);
and U35586 (N_35586,N_32316,N_33495);
and U35587 (N_35587,N_32826,N_32121);
nand U35588 (N_35588,N_32877,N_33436);
nor U35589 (N_35589,N_33861,N_33708);
and U35590 (N_35590,N_33659,N_33587);
xor U35591 (N_35591,N_32850,N_32939);
and U35592 (N_35592,N_33461,N_33313);
or U35593 (N_35593,N_32005,N_32310);
nand U35594 (N_35594,N_32818,N_33220);
xnor U35595 (N_35595,N_32407,N_32893);
nand U35596 (N_35596,N_32336,N_33001);
xor U35597 (N_35597,N_32022,N_33351);
nand U35598 (N_35598,N_33109,N_32545);
xnor U35599 (N_35599,N_32472,N_32232);
nor U35600 (N_35600,N_33377,N_33096);
xnor U35601 (N_35601,N_32400,N_32563);
nor U35602 (N_35602,N_33735,N_32160);
nor U35603 (N_35603,N_32484,N_33893);
or U35604 (N_35604,N_32975,N_32844);
nand U35605 (N_35605,N_33611,N_32526);
xnor U35606 (N_35606,N_32112,N_33485);
xnor U35607 (N_35607,N_32834,N_33772);
nor U35608 (N_35608,N_33970,N_32640);
or U35609 (N_35609,N_33107,N_33405);
nand U35610 (N_35610,N_32361,N_32867);
nand U35611 (N_35611,N_33954,N_33974);
nor U35612 (N_35612,N_32065,N_33670);
xnor U35613 (N_35613,N_33873,N_33302);
or U35614 (N_35614,N_32092,N_32058);
nand U35615 (N_35615,N_33072,N_33294);
xnor U35616 (N_35616,N_33593,N_33990);
nand U35617 (N_35617,N_33893,N_32907);
nand U35618 (N_35618,N_32941,N_32692);
xor U35619 (N_35619,N_32192,N_32525);
and U35620 (N_35620,N_33152,N_32578);
nand U35621 (N_35621,N_32211,N_33405);
and U35622 (N_35622,N_32182,N_33326);
xor U35623 (N_35623,N_32703,N_33819);
or U35624 (N_35624,N_33597,N_32070);
and U35625 (N_35625,N_33507,N_32784);
xnor U35626 (N_35626,N_32787,N_32962);
or U35627 (N_35627,N_32737,N_32063);
or U35628 (N_35628,N_32318,N_33118);
nand U35629 (N_35629,N_32269,N_32858);
xnor U35630 (N_35630,N_32730,N_33841);
or U35631 (N_35631,N_33227,N_33457);
or U35632 (N_35632,N_33784,N_32452);
xnor U35633 (N_35633,N_33014,N_33965);
and U35634 (N_35634,N_33285,N_33876);
or U35635 (N_35635,N_32693,N_33932);
xnor U35636 (N_35636,N_33248,N_33771);
and U35637 (N_35637,N_33871,N_33949);
or U35638 (N_35638,N_33330,N_32210);
nand U35639 (N_35639,N_32999,N_33532);
xor U35640 (N_35640,N_32502,N_33976);
and U35641 (N_35641,N_33985,N_33093);
or U35642 (N_35642,N_32543,N_32383);
xor U35643 (N_35643,N_33415,N_32497);
nor U35644 (N_35644,N_32702,N_32690);
nor U35645 (N_35645,N_33845,N_33529);
or U35646 (N_35646,N_33304,N_33661);
and U35647 (N_35647,N_32797,N_32111);
nor U35648 (N_35648,N_32641,N_32842);
and U35649 (N_35649,N_33000,N_32077);
nor U35650 (N_35650,N_32516,N_33199);
nor U35651 (N_35651,N_33422,N_33337);
or U35652 (N_35652,N_32711,N_32060);
nand U35653 (N_35653,N_32752,N_32032);
xor U35654 (N_35654,N_32877,N_32441);
or U35655 (N_35655,N_32172,N_33488);
or U35656 (N_35656,N_32722,N_33419);
nand U35657 (N_35657,N_33731,N_32002);
nor U35658 (N_35658,N_33692,N_32554);
nor U35659 (N_35659,N_32423,N_33649);
xnor U35660 (N_35660,N_32232,N_33568);
nand U35661 (N_35661,N_32781,N_33493);
nor U35662 (N_35662,N_33618,N_32487);
nor U35663 (N_35663,N_32448,N_33604);
and U35664 (N_35664,N_33366,N_33510);
nor U35665 (N_35665,N_32543,N_33905);
and U35666 (N_35666,N_32819,N_33418);
nor U35667 (N_35667,N_33867,N_33400);
and U35668 (N_35668,N_32639,N_33238);
or U35669 (N_35669,N_32362,N_32288);
or U35670 (N_35670,N_33086,N_32784);
xor U35671 (N_35671,N_33368,N_33421);
nor U35672 (N_35672,N_33210,N_33997);
nand U35673 (N_35673,N_32587,N_33523);
nor U35674 (N_35674,N_33647,N_32150);
nand U35675 (N_35675,N_33490,N_33716);
or U35676 (N_35676,N_33622,N_32040);
nand U35677 (N_35677,N_32044,N_33911);
xor U35678 (N_35678,N_32373,N_32034);
nand U35679 (N_35679,N_33554,N_32180);
or U35680 (N_35680,N_33678,N_32739);
nor U35681 (N_35681,N_32900,N_32475);
nor U35682 (N_35682,N_32538,N_33678);
xor U35683 (N_35683,N_33193,N_33575);
nor U35684 (N_35684,N_33410,N_32999);
nor U35685 (N_35685,N_32111,N_33940);
nand U35686 (N_35686,N_33452,N_33196);
and U35687 (N_35687,N_32543,N_33590);
nand U35688 (N_35688,N_33881,N_32760);
xor U35689 (N_35689,N_33847,N_32513);
or U35690 (N_35690,N_33352,N_33923);
nand U35691 (N_35691,N_32819,N_32985);
and U35692 (N_35692,N_32678,N_32711);
nor U35693 (N_35693,N_33971,N_33419);
xor U35694 (N_35694,N_32894,N_33707);
or U35695 (N_35695,N_32184,N_32446);
or U35696 (N_35696,N_32052,N_33505);
nor U35697 (N_35697,N_33087,N_33953);
nor U35698 (N_35698,N_32079,N_33150);
and U35699 (N_35699,N_32800,N_32985);
xor U35700 (N_35700,N_33656,N_33871);
or U35701 (N_35701,N_32120,N_33775);
and U35702 (N_35702,N_32720,N_32058);
or U35703 (N_35703,N_33919,N_32628);
xor U35704 (N_35704,N_32203,N_33986);
xnor U35705 (N_35705,N_32605,N_32047);
nor U35706 (N_35706,N_32807,N_32055);
nand U35707 (N_35707,N_32419,N_33875);
nor U35708 (N_35708,N_33100,N_33115);
nor U35709 (N_35709,N_32747,N_33323);
nor U35710 (N_35710,N_32703,N_32072);
nor U35711 (N_35711,N_32263,N_33261);
or U35712 (N_35712,N_32267,N_32998);
or U35713 (N_35713,N_32744,N_32507);
and U35714 (N_35714,N_33895,N_32883);
or U35715 (N_35715,N_32544,N_33298);
or U35716 (N_35716,N_32470,N_32549);
nand U35717 (N_35717,N_33904,N_33880);
and U35718 (N_35718,N_32938,N_33382);
or U35719 (N_35719,N_33519,N_32356);
nand U35720 (N_35720,N_32146,N_32737);
and U35721 (N_35721,N_32009,N_32383);
or U35722 (N_35722,N_33663,N_32506);
or U35723 (N_35723,N_32827,N_32962);
and U35724 (N_35724,N_32587,N_33300);
nor U35725 (N_35725,N_33269,N_32807);
and U35726 (N_35726,N_32267,N_33495);
nand U35727 (N_35727,N_32652,N_33971);
nand U35728 (N_35728,N_33874,N_33237);
or U35729 (N_35729,N_32943,N_33710);
and U35730 (N_35730,N_33102,N_32686);
and U35731 (N_35731,N_33746,N_33888);
xor U35732 (N_35732,N_32837,N_33973);
nor U35733 (N_35733,N_33462,N_33556);
xor U35734 (N_35734,N_33326,N_33095);
nand U35735 (N_35735,N_32129,N_32986);
and U35736 (N_35736,N_32587,N_33222);
xnor U35737 (N_35737,N_32271,N_33582);
and U35738 (N_35738,N_33853,N_32332);
nor U35739 (N_35739,N_33741,N_33383);
and U35740 (N_35740,N_32918,N_33938);
xnor U35741 (N_35741,N_32943,N_32677);
nand U35742 (N_35742,N_32728,N_33096);
nor U35743 (N_35743,N_32248,N_32892);
nor U35744 (N_35744,N_33566,N_32372);
nor U35745 (N_35745,N_33080,N_33893);
xnor U35746 (N_35746,N_33251,N_33970);
or U35747 (N_35747,N_32541,N_33662);
nor U35748 (N_35748,N_33937,N_32330);
nor U35749 (N_35749,N_33668,N_32039);
or U35750 (N_35750,N_32054,N_33284);
xnor U35751 (N_35751,N_32081,N_33852);
xnor U35752 (N_35752,N_33100,N_32058);
nand U35753 (N_35753,N_33052,N_33503);
nand U35754 (N_35754,N_32103,N_32096);
nor U35755 (N_35755,N_33283,N_32873);
xor U35756 (N_35756,N_33482,N_32270);
nor U35757 (N_35757,N_32893,N_32589);
or U35758 (N_35758,N_33271,N_33235);
xor U35759 (N_35759,N_33331,N_33741);
and U35760 (N_35760,N_33877,N_32326);
nor U35761 (N_35761,N_32872,N_33255);
nand U35762 (N_35762,N_32623,N_32915);
nor U35763 (N_35763,N_32101,N_33100);
or U35764 (N_35764,N_33194,N_33597);
or U35765 (N_35765,N_32186,N_32753);
or U35766 (N_35766,N_32835,N_32076);
and U35767 (N_35767,N_32514,N_33078);
and U35768 (N_35768,N_33514,N_33858);
nor U35769 (N_35769,N_32566,N_32800);
and U35770 (N_35770,N_32548,N_32260);
and U35771 (N_35771,N_33184,N_33535);
nor U35772 (N_35772,N_33092,N_32734);
or U35773 (N_35773,N_33163,N_32057);
and U35774 (N_35774,N_32540,N_32230);
xnor U35775 (N_35775,N_33877,N_32584);
and U35776 (N_35776,N_33648,N_32393);
xor U35777 (N_35777,N_32063,N_32950);
nand U35778 (N_35778,N_32152,N_32290);
xnor U35779 (N_35779,N_33815,N_32877);
nor U35780 (N_35780,N_33299,N_32830);
xnor U35781 (N_35781,N_32953,N_33755);
and U35782 (N_35782,N_33469,N_32304);
and U35783 (N_35783,N_33533,N_33112);
nand U35784 (N_35784,N_33675,N_32284);
xnor U35785 (N_35785,N_33018,N_33543);
nand U35786 (N_35786,N_32587,N_33376);
nor U35787 (N_35787,N_32685,N_33847);
nor U35788 (N_35788,N_33120,N_33482);
and U35789 (N_35789,N_32599,N_32582);
xor U35790 (N_35790,N_33549,N_33990);
xnor U35791 (N_35791,N_32028,N_33601);
nor U35792 (N_35792,N_33111,N_33848);
nand U35793 (N_35793,N_33722,N_33997);
or U35794 (N_35794,N_32688,N_32087);
xor U35795 (N_35795,N_32136,N_32796);
nand U35796 (N_35796,N_32251,N_32793);
and U35797 (N_35797,N_33809,N_33237);
and U35798 (N_35798,N_32442,N_33193);
xnor U35799 (N_35799,N_33754,N_33616);
and U35800 (N_35800,N_33354,N_32845);
xor U35801 (N_35801,N_32331,N_33481);
nor U35802 (N_35802,N_32142,N_33809);
or U35803 (N_35803,N_32956,N_33578);
xor U35804 (N_35804,N_32554,N_33784);
and U35805 (N_35805,N_32726,N_32277);
or U35806 (N_35806,N_33751,N_33890);
nand U35807 (N_35807,N_33543,N_33166);
and U35808 (N_35808,N_32927,N_32172);
or U35809 (N_35809,N_33851,N_32741);
nand U35810 (N_35810,N_33784,N_32577);
nand U35811 (N_35811,N_32227,N_33230);
xnor U35812 (N_35812,N_33465,N_33649);
xor U35813 (N_35813,N_33054,N_32644);
and U35814 (N_35814,N_33312,N_32876);
and U35815 (N_35815,N_32322,N_32688);
and U35816 (N_35816,N_33707,N_33591);
nand U35817 (N_35817,N_32061,N_32898);
xnor U35818 (N_35818,N_33773,N_33939);
and U35819 (N_35819,N_33453,N_33158);
and U35820 (N_35820,N_33649,N_32068);
or U35821 (N_35821,N_32953,N_32922);
xor U35822 (N_35822,N_32855,N_32934);
or U35823 (N_35823,N_32127,N_32487);
nor U35824 (N_35824,N_32575,N_32104);
or U35825 (N_35825,N_33524,N_33377);
nand U35826 (N_35826,N_32570,N_33328);
nor U35827 (N_35827,N_32229,N_33401);
or U35828 (N_35828,N_33747,N_33787);
nor U35829 (N_35829,N_32077,N_33118);
and U35830 (N_35830,N_32482,N_33729);
and U35831 (N_35831,N_32636,N_32170);
nand U35832 (N_35832,N_33991,N_32523);
nand U35833 (N_35833,N_33118,N_33408);
nand U35834 (N_35834,N_32317,N_32687);
nand U35835 (N_35835,N_33574,N_32277);
and U35836 (N_35836,N_32678,N_32242);
nor U35837 (N_35837,N_32002,N_32603);
xnor U35838 (N_35838,N_32996,N_32665);
nand U35839 (N_35839,N_32525,N_33567);
xnor U35840 (N_35840,N_32428,N_33138);
nand U35841 (N_35841,N_33413,N_32101);
or U35842 (N_35842,N_33224,N_33160);
xnor U35843 (N_35843,N_33551,N_32026);
or U35844 (N_35844,N_32968,N_33695);
and U35845 (N_35845,N_33580,N_32864);
nor U35846 (N_35846,N_33301,N_32549);
xor U35847 (N_35847,N_32574,N_32018);
and U35848 (N_35848,N_32672,N_33927);
nand U35849 (N_35849,N_32423,N_33981);
xnor U35850 (N_35850,N_32399,N_32961);
or U35851 (N_35851,N_32850,N_33881);
and U35852 (N_35852,N_32368,N_33981);
xor U35853 (N_35853,N_33080,N_33757);
and U35854 (N_35854,N_32691,N_32213);
nor U35855 (N_35855,N_32394,N_33352);
xor U35856 (N_35856,N_33445,N_32444);
or U35857 (N_35857,N_32634,N_33119);
or U35858 (N_35858,N_32561,N_32949);
xnor U35859 (N_35859,N_32514,N_33085);
or U35860 (N_35860,N_32863,N_33368);
or U35861 (N_35861,N_33598,N_32468);
or U35862 (N_35862,N_32296,N_33489);
nand U35863 (N_35863,N_33294,N_33809);
xor U35864 (N_35864,N_33993,N_32844);
nor U35865 (N_35865,N_33232,N_32351);
nor U35866 (N_35866,N_33323,N_33636);
nor U35867 (N_35867,N_33193,N_33999);
nor U35868 (N_35868,N_32605,N_33087);
nor U35869 (N_35869,N_33817,N_33544);
xor U35870 (N_35870,N_32252,N_32706);
nor U35871 (N_35871,N_32914,N_33381);
nor U35872 (N_35872,N_33263,N_33692);
nor U35873 (N_35873,N_32715,N_32290);
nand U35874 (N_35874,N_33610,N_33041);
or U35875 (N_35875,N_32210,N_33729);
nand U35876 (N_35876,N_32051,N_33020);
nor U35877 (N_35877,N_33224,N_33078);
xor U35878 (N_35878,N_32224,N_33973);
xnor U35879 (N_35879,N_33143,N_33576);
nand U35880 (N_35880,N_32277,N_33660);
or U35881 (N_35881,N_32108,N_32467);
and U35882 (N_35882,N_32366,N_33668);
or U35883 (N_35883,N_33485,N_33007);
nand U35884 (N_35884,N_32107,N_32666);
xor U35885 (N_35885,N_32965,N_32922);
or U35886 (N_35886,N_33909,N_33540);
and U35887 (N_35887,N_32014,N_33534);
or U35888 (N_35888,N_33905,N_32157);
xnor U35889 (N_35889,N_32542,N_32524);
nand U35890 (N_35890,N_33606,N_33506);
nor U35891 (N_35891,N_33774,N_32703);
xnor U35892 (N_35892,N_32629,N_33863);
or U35893 (N_35893,N_32214,N_33601);
xor U35894 (N_35894,N_32883,N_33556);
and U35895 (N_35895,N_32758,N_33766);
nor U35896 (N_35896,N_33285,N_32787);
nand U35897 (N_35897,N_33266,N_33857);
or U35898 (N_35898,N_32810,N_33660);
or U35899 (N_35899,N_33924,N_33361);
nor U35900 (N_35900,N_32400,N_32187);
or U35901 (N_35901,N_32390,N_33638);
xnor U35902 (N_35902,N_32229,N_33584);
xnor U35903 (N_35903,N_33554,N_32758);
xor U35904 (N_35904,N_33299,N_33322);
nor U35905 (N_35905,N_33598,N_32726);
nor U35906 (N_35906,N_33389,N_33877);
nand U35907 (N_35907,N_32816,N_32143);
or U35908 (N_35908,N_32622,N_33059);
or U35909 (N_35909,N_33214,N_32730);
nand U35910 (N_35910,N_33767,N_33257);
and U35911 (N_35911,N_32665,N_32414);
xor U35912 (N_35912,N_32794,N_32156);
nand U35913 (N_35913,N_32878,N_33582);
nor U35914 (N_35914,N_32919,N_32479);
nor U35915 (N_35915,N_33888,N_32580);
xor U35916 (N_35916,N_33331,N_32056);
nor U35917 (N_35917,N_33040,N_32887);
xnor U35918 (N_35918,N_32142,N_32611);
xor U35919 (N_35919,N_33190,N_33152);
xor U35920 (N_35920,N_33430,N_32847);
xor U35921 (N_35921,N_33644,N_33610);
nand U35922 (N_35922,N_32316,N_32815);
nand U35923 (N_35923,N_33556,N_32298);
or U35924 (N_35924,N_32014,N_32199);
xnor U35925 (N_35925,N_32648,N_33607);
nand U35926 (N_35926,N_33245,N_32883);
or U35927 (N_35927,N_32460,N_32006);
nor U35928 (N_35928,N_32359,N_33238);
nand U35929 (N_35929,N_32926,N_33981);
nand U35930 (N_35930,N_33027,N_33852);
and U35931 (N_35931,N_33156,N_33468);
nand U35932 (N_35932,N_33819,N_32266);
nor U35933 (N_35933,N_33938,N_32231);
nor U35934 (N_35934,N_32466,N_32011);
xnor U35935 (N_35935,N_32321,N_33716);
nand U35936 (N_35936,N_32934,N_32491);
xnor U35937 (N_35937,N_33847,N_33463);
nor U35938 (N_35938,N_32902,N_33010);
xor U35939 (N_35939,N_33694,N_32714);
nand U35940 (N_35940,N_32899,N_33272);
or U35941 (N_35941,N_32463,N_32335);
or U35942 (N_35942,N_33378,N_32017);
or U35943 (N_35943,N_33832,N_33643);
nand U35944 (N_35944,N_32349,N_33603);
nor U35945 (N_35945,N_32000,N_32794);
and U35946 (N_35946,N_33143,N_32329);
or U35947 (N_35947,N_33397,N_33763);
nand U35948 (N_35948,N_32931,N_33031);
xor U35949 (N_35949,N_32839,N_32587);
nand U35950 (N_35950,N_32883,N_32626);
and U35951 (N_35951,N_33981,N_33627);
nor U35952 (N_35952,N_33015,N_33039);
xor U35953 (N_35953,N_32567,N_32890);
nor U35954 (N_35954,N_33059,N_33385);
and U35955 (N_35955,N_32590,N_32648);
or U35956 (N_35956,N_32963,N_33875);
or U35957 (N_35957,N_32672,N_33579);
and U35958 (N_35958,N_33447,N_33718);
xor U35959 (N_35959,N_33256,N_32125);
and U35960 (N_35960,N_33408,N_32776);
nand U35961 (N_35961,N_32669,N_32018);
xor U35962 (N_35962,N_32801,N_32616);
nand U35963 (N_35963,N_32888,N_32906);
or U35964 (N_35964,N_33199,N_33878);
and U35965 (N_35965,N_33368,N_32349);
and U35966 (N_35966,N_32071,N_32622);
nand U35967 (N_35967,N_32626,N_33583);
xnor U35968 (N_35968,N_32578,N_33566);
or U35969 (N_35969,N_33889,N_32681);
nor U35970 (N_35970,N_32346,N_33789);
and U35971 (N_35971,N_33660,N_32446);
nor U35972 (N_35972,N_32294,N_33489);
nor U35973 (N_35973,N_32104,N_32325);
and U35974 (N_35974,N_33880,N_32842);
or U35975 (N_35975,N_32641,N_32220);
or U35976 (N_35976,N_32980,N_32562);
and U35977 (N_35977,N_33085,N_32460);
nand U35978 (N_35978,N_32290,N_33451);
and U35979 (N_35979,N_32695,N_32982);
or U35980 (N_35980,N_33123,N_32164);
xnor U35981 (N_35981,N_33212,N_33906);
xnor U35982 (N_35982,N_33907,N_33294);
and U35983 (N_35983,N_33716,N_33801);
and U35984 (N_35984,N_33713,N_33896);
nand U35985 (N_35985,N_32037,N_32501);
nor U35986 (N_35986,N_33649,N_32997);
or U35987 (N_35987,N_32175,N_33949);
or U35988 (N_35988,N_33593,N_33367);
or U35989 (N_35989,N_33619,N_32774);
xnor U35990 (N_35990,N_32705,N_33149);
xor U35991 (N_35991,N_33339,N_32765);
nor U35992 (N_35992,N_32851,N_32119);
nor U35993 (N_35993,N_33977,N_32901);
xnor U35994 (N_35994,N_33380,N_32152);
xnor U35995 (N_35995,N_32198,N_32875);
or U35996 (N_35996,N_32624,N_32291);
or U35997 (N_35997,N_33442,N_32627);
nand U35998 (N_35998,N_33153,N_32229);
nand U35999 (N_35999,N_32174,N_32087);
nor U36000 (N_36000,N_34677,N_34950);
and U36001 (N_36001,N_35721,N_35935);
nand U36002 (N_36002,N_35951,N_34893);
or U36003 (N_36003,N_34493,N_34113);
xor U36004 (N_36004,N_34654,N_34690);
and U36005 (N_36005,N_34014,N_35858);
or U36006 (N_36006,N_34152,N_34625);
nor U36007 (N_36007,N_35647,N_35225);
or U36008 (N_36008,N_35822,N_35749);
nand U36009 (N_36009,N_34088,N_34849);
and U36010 (N_36010,N_34208,N_35844);
or U36011 (N_36011,N_34560,N_35271);
xnor U36012 (N_36012,N_35881,N_35253);
and U36013 (N_36013,N_34920,N_35702);
xor U36014 (N_36014,N_35382,N_35366);
xnor U36015 (N_36015,N_34610,N_34706);
nand U36016 (N_36016,N_34639,N_34028);
and U36017 (N_36017,N_35354,N_34843);
or U36018 (N_36018,N_34636,N_35661);
nand U36019 (N_36019,N_34653,N_35226);
xor U36020 (N_36020,N_34987,N_34705);
nand U36021 (N_36021,N_34886,N_35241);
nor U36022 (N_36022,N_35758,N_35407);
nor U36023 (N_36023,N_35638,N_34575);
or U36024 (N_36024,N_35133,N_35415);
or U36025 (N_36025,N_35047,N_34070);
and U36026 (N_36026,N_35768,N_34366);
nand U36027 (N_36027,N_34289,N_35350);
and U36028 (N_36028,N_35213,N_35677);
or U36029 (N_36029,N_34368,N_34490);
nand U36030 (N_36030,N_35479,N_35869);
or U36031 (N_36031,N_35641,N_35900);
nand U36032 (N_36032,N_34558,N_34206);
or U36033 (N_36033,N_34561,N_34486);
nand U36034 (N_36034,N_34295,N_34091);
nand U36035 (N_36035,N_35733,N_34660);
nand U36036 (N_36036,N_35142,N_34500);
nand U36037 (N_36037,N_34124,N_34433);
xor U36038 (N_36038,N_35052,N_35372);
and U36039 (N_36039,N_35176,N_35347);
or U36040 (N_36040,N_34032,N_35195);
and U36041 (N_36041,N_35705,N_35989);
nand U36042 (N_36042,N_34202,N_35408);
nor U36043 (N_36043,N_34929,N_34156);
xnor U36044 (N_36044,N_34995,N_35897);
nand U36045 (N_36045,N_35919,N_34195);
and U36046 (N_36046,N_34443,N_34543);
or U36047 (N_36047,N_34919,N_35077);
nor U36048 (N_36048,N_34780,N_35614);
nand U36049 (N_36049,N_34082,N_34530);
and U36050 (N_36050,N_34686,N_34376);
xnor U36051 (N_36051,N_35853,N_34139);
nand U36052 (N_36052,N_34890,N_35363);
xor U36053 (N_36053,N_34421,N_35006);
and U36054 (N_36054,N_34205,N_35492);
xnor U36055 (N_36055,N_34744,N_34984);
nand U36056 (N_36056,N_34297,N_35083);
nor U36057 (N_36057,N_34661,N_34906);
nor U36058 (N_36058,N_35927,N_34727);
and U36059 (N_36059,N_35055,N_35180);
nor U36060 (N_36060,N_34072,N_34630);
or U36061 (N_36061,N_35068,N_34483);
nor U36062 (N_36062,N_35623,N_34916);
xnor U36063 (N_36063,N_35802,N_34436);
or U36064 (N_36064,N_35866,N_34798);
and U36065 (N_36065,N_35712,N_34467);
xnor U36066 (N_36066,N_34214,N_35544);
xnor U36067 (N_36067,N_35940,N_34182);
xor U36068 (N_36068,N_34027,N_35442);
nor U36069 (N_36069,N_35400,N_35526);
nand U36070 (N_36070,N_35154,N_34932);
or U36071 (N_36071,N_34374,N_35141);
or U36072 (N_36072,N_34167,N_35737);
xnor U36073 (N_36073,N_34823,N_34528);
nand U36074 (N_36074,N_35509,N_34790);
xor U36075 (N_36075,N_34311,N_35459);
nor U36076 (N_36076,N_35717,N_34682);
xor U36077 (N_36077,N_35558,N_35275);
or U36078 (N_36078,N_34952,N_35973);
nor U36079 (N_36079,N_35748,N_34701);
and U36080 (N_36080,N_34938,N_35388);
and U36081 (N_36081,N_34512,N_34855);
xor U36082 (N_36082,N_34328,N_34544);
xnor U36083 (N_36083,N_35863,N_34618);
xnor U36084 (N_36084,N_34187,N_35918);
nor U36085 (N_36085,N_34656,N_35824);
or U36086 (N_36086,N_34079,N_34393);
xor U36087 (N_36087,N_34990,N_35430);
nand U36088 (N_36088,N_34840,N_35106);
nor U36089 (N_36089,N_34506,N_34410);
or U36090 (N_36090,N_34779,N_34522);
and U36091 (N_36091,N_34137,N_34339);
xor U36092 (N_36092,N_35123,N_35530);
xnor U36093 (N_36093,N_34818,N_34135);
and U36094 (N_36094,N_35199,N_35126);
and U36095 (N_36095,N_34239,N_35117);
or U36096 (N_36096,N_34708,N_34737);
and U36097 (N_36097,N_34684,N_34336);
or U36098 (N_36098,N_35628,N_35567);
nand U36099 (N_36099,N_34250,N_34056);
nand U36100 (N_36100,N_34478,N_34674);
xnor U36101 (N_36101,N_34894,N_34900);
nand U36102 (N_36102,N_34590,N_34983);
or U36103 (N_36103,N_35483,N_35284);
or U36104 (N_36104,N_34658,N_34060);
nand U36105 (N_36105,N_35140,N_34918);
nor U36106 (N_36106,N_35086,N_35913);
xnor U36107 (N_36107,N_34911,N_35860);
nand U36108 (N_36108,N_34848,N_35198);
nor U36109 (N_36109,N_34564,N_35865);
or U36110 (N_36110,N_35118,N_35809);
nand U36111 (N_36111,N_35839,N_35320);
and U36112 (N_36112,N_35091,N_35619);
or U36113 (N_36113,N_35201,N_34691);
nor U36114 (N_36114,N_34363,N_34271);
nor U36115 (N_36115,N_35132,N_35773);
and U36116 (N_36116,N_35481,N_34966);
or U36117 (N_36117,N_35626,N_34043);
or U36118 (N_36118,N_35044,N_34021);
nor U36119 (N_36119,N_35398,N_35110);
xor U36120 (N_36120,N_35362,N_34872);
and U36121 (N_36121,N_35827,N_35531);
xnor U36122 (N_36122,N_35690,N_34867);
nor U36123 (N_36123,N_35533,N_34634);
or U36124 (N_36124,N_35963,N_34449);
nand U36125 (N_36125,N_35143,N_34411);
nand U36126 (N_36126,N_34216,N_35668);
nand U36127 (N_36127,N_35490,N_35672);
nor U36128 (N_36128,N_35801,N_35013);
or U36129 (N_36129,N_34972,N_35611);
or U36130 (N_36130,N_35975,N_34059);
xor U36131 (N_36131,N_34494,N_35417);
or U36132 (N_36132,N_34108,N_34819);
xor U36133 (N_36133,N_35129,N_34054);
or U36134 (N_36134,N_34314,N_34240);
nand U36135 (N_36135,N_35682,N_34852);
or U36136 (N_36136,N_34540,N_34954);
nor U36137 (N_36137,N_35293,N_35826);
nor U36138 (N_36138,N_34412,N_34310);
and U36139 (N_36139,N_34621,N_34236);
nand U36140 (N_36140,N_34683,N_35834);
or U36141 (N_36141,N_35580,N_34902);
xnor U36142 (N_36142,N_34342,N_35755);
or U36143 (N_36143,N_35200,N_34642);
xor U36144 (N_36144,N_35384,N_35561);
nand U36145 (N_36145,N_35263,N_35878);
or U36146 (N_36146,N_35676,N_34169);
nor U36147 (N_36147,N_35122,N_34773);
xnor U36148 (N_36148,N_34833,N_35740);
nand U36149 (N_36149,N_35174,N_35114);
nor U36150 (N_36150,N_34510,N_35447);
and U36151 (N_36151,N_35903,N_35757);
nor U36152 (N_36152,N_34860,N_35080);
nor U36153 (N_36153,N_34158,N_35317);
nor U36154 (N_36154,N_34948,N_35152);
nor U36155 (N_36155,N_35179,N_34270);
nor U36156 (N_36156,N_35039,N_34107);
nor U36157 (N_36157,N_34042,N_34749);
nor U36158 (N_36158,N_35852,N_34365);
xnor U36159 (N_36159,N_35026,N_35663);
nand U36160 (N_36160,N_35011,N_35723);
or U36161 (N_36161,N_34509,N_35751);
nand U36162 (N_36162,N_34098,N_34907);
or U36163 (N_36163,N_35867,N_35589);
or U36164 (N_36164,N_35000,N_35428);
nand U36165 (N_36165,N_35437,N_35028);
or U36166 (N_36166,N_34742,N_34864);
nand U36167 (N_36167,N_34178,N_34055);
xnor U36168 (N_36168,N_35246,N_35703);
nand U36169 (N_36169,N_34981,N_35770);
or U36170 (N_36170,N_35019,N_34891);
nor U36171 (N_36171,N_35351,N_35411);
nand U36172 (N_36172,N_35798,N_35596);
nor U36173 (N_36173,N_35244,N_34430);
and U36174 (N_36174,N_35454,N_34184);
and U36175 (N_36175,N_34259,N_34445);
or U36176 (N_36176,N_35082,N_34896);
nor U36177 (N_36177,N_34306,N_35169);
and U36178 (N_36178,N_35714,N_34804);
nor U36179 (N_36179,N_35393,N_34740);
xnor U36180 (N_36180,N_34587,N_35840);
or U36181 (N_36181,N_34163,N_34909);
nand U36182 (N_36182,N_35762,N_35831);
and U36183 (N_36183,N_34541,N_35707);
and U36184 (N_36184,N_34360,N_34667);
nor U36185 (N_36185,N_34053,N_34065);
and U36186 (N_36186,N_35559,N_34130);
nor U36187 (N_36187,N_34504,N_35528);
nor U36188 (N_36188,N_34067,N_35220);
nor U36189 (N_36189,N_34024,N_34762);
or U36190 (N_36190,N_35054,N_34772);
and U36191 (N_36191,N_35997,N_34317);
or U36192 (N_36192,N_34877,N_34707);
xor U36193 (N_36193,N_34887,N_34956);
xnor U36194 (N_36194,N_34424,N_35609);
or U36195 (N_36195,N_35806,N_35074);
or U36196 (N_36196,N_35352,N_34034);
nand U36197 (N_36197,N_34148,N_34489);
xnor U36198 (N_36198,N_35273,N_34322);
xor U36199 (N_36199,N_35189,N_35261);
nand U36200 (N_36200,N_35353,N_34928);
or U36201 (N_36201,N_34598,N_35945);
xnor U36202 (N_36202,N_34614,N_35958);
and U36203 (N_36203,N_34892,N_35786);
nor U36204 (N_36204,N_34232,N_35207);
nor U36205 (N_36205,N_35204,N_34331);
xnor U36206 (N_36206,N_34930,N_35929);
or U36207 (N_36207,N_35608,N_35099);
nand U36208 (N_36208,N_34353,N_35771);
xor U36209 (N_36209,N_34479,N_34570);
xnor U36210 (N_36210,N_35370,N_34793);
nand U36211 (N_36211,N_35256,N_35949);
nand U36212 (N_36212,N_34738,N_34764);
or U36213 (N_36213,N_34334,N_35078);
nor U36214 (N_36214,N_35440,N_35984);
and U36215 (N_36215,N_35633,N_34097);
and U36216 (N_36216,N_35874,N_34300);
nor U36217 (N_36217,N_34038,N_34235);
nor U36218 (N_36218,N_34125,N_34358);
or U36219 (N_36219,N_34454,N_35727);
xnor U36220 (N_36220,N_35891,N_34718);
or U36221 (N_36221,N_35178,N_34809);
nor U36222 (N_36222,N_34471,N_34037);
and U36223 (N_36223,N_34689,N_35349);
nor U36224 (N_36224,N_35911,N_35513);
or U36225 (N_36225,N_34562,N_34626);
and U36226 (N_36226,N_34709,N_35412);
nor U36227 (N_36227,N_35257,N_35267);
xnor U36228 (N_36228,N_35519,N_34402);
and U36229 (N_36229,N_34847,N_35542);
or U36230 (N_36230,N_34023,N_35890);
and U36231 (N_36231,N_35644,N_34347);
and U36232 (N_36232,N_35240,N_35171);
and U36233 (N_36233,N_34251,N_35337);
or U36234 (N_36234,N_34255,N_35796);
xor U36235 (N_36235,N_35566,N_34061);
or U36236 (N_36236,N_35998,N_35165);
and U36237 (N_36237,N_34190,N_35836);
nor U36238 (N_36238,N_34497,N_34815);
nand U36239 (N_36239,N_35683,N_35694);
xor U36240 (N_36240,N_35007,N_34794);
nand U36241 (N_36241,N_34778,N_34947);
nand U36242 (N_36242,N_34977,N_34588);
nand U36243 (N_36243,N_34549,N_35475);
nor U36244 (N_36244,N_34666,N_34371);
or U36245 (N_36245,N_34595,N_35194);
nor U36246 (N_36246,N_34465,N_35265);
xnor U36247 (N_36247,N_35805,N_34796);
and U36248 (N_36248,N_35675,N_34219);
nand U36249 (N_36249,N_35322,N_35323);
nand U36250 (N_36250,N_35234,N_35906);
xnor U36251 (N_36251,N_34939,N_34631);
nand U36252 (N_36252,N_34172,N_35395);
nand U36253 (N_36253,N_35954,N_34143);
and U36254 (N_36254,N_35286,N_35760);
and U36255 (N_36255,N_35653,N_35312);
xor U36256 (N_36256,N_34370,N_34451);
and U36257 (N_36257,N_35334,N_35095);
nor U36258 (N_36258,N_34761,N_35765);
and U36259 (N_36259,N_35879,N_35811);
and U36260 (N_36260,N_35947,N_35208);
nor U36261 (N_36261,N_35423,N_34385);
xor U36262 (N_36262,N_35445,N_35134);
xor U36263 (N_36263,N_35792,N_35472);
and U36264 (N_36264,N_35688,N_34730);
and U36265 (N_36265,N_34234,N_34559);
and U36266 (N_36266,N_35974,N_34352);
nand U36267 (N_36267,N_35851,N_34924);
nor U36268 (N_36268,N_34556,N_35387);
or U36269 (N_36269,N_34523,N_34937);
nand U36270 (N_36270,N_35752,N_35592);
xor U36271 (N_36271,N_34294,N_35983);
nand U36272 (N_36272,N_35987,N_35642);
nor U36273 (N_36273,N_34222,N_34080);
nor U36274 (N_36274,N_34777,N_34462);
or U36275 (N_36275,N_34601,N_34285);
nor U36276 (N_36276,N_34111,N_34927);
or U36277 (N_36277,N_35767,N_35730);
or U36278 (N_36278,N_34752,N_35184);
xnor U36279 (N_36279,N_34011,N_35885);
xnor U36280 (N_36280,N_34399,N_34694);
or U36281 (N_36281,N_35462,N_34305);
nand U36282 (N_36282,N_34046,N_35789);
or U36283 (N_36283,N_34498,N_35441);
or U36284 (N_36284,N_35264,N_34333);
or U36285 (N_36285,N_35465,N_34717);
xnor U36286 (N_36286,N_34142,N_35986);
or U36287 (N_36287,N_35590,N_34254);
xor U36288 (N_36288,N_34505,N_35237);
nand U36289 (N_36289,N_34600,N_35988);
and U36290 (N_36290,N_35904,N_34212);
nor U36291 (N_36291,N_35072,N_34612);
or U36292 (N_36292,N_35438,N_34982);
or U36293 (N_36293,N_34678,N_35955);
nor U36294 (N_36294,N_34280,N_35894);
xnor U36295 (N_36295,N_34484,N_35346);
or U36296 (N_36296,N_35923,N_35329);
xor U36297 (N_36297,N_34101,N_35845);
and U36298 (N_36298,N_34378,N_34406);
and U36299 (N_36299,N_35009,N_34791);
and U36300 (N_36300,N_34058,N_34233);
or U36301 (N_36301,N_35260,N_35431);
or U36302 (N_36302,N_35756,N_34400);
nand U36303 (N_36303,N_34487,N_34367);
xor U36304 (N_36304,N_34585,N_34403);
xnor U36305 (N_36305,N_34116,N_34957);
xnor U36306 (N_36306,N_35124,N_34469);
xor U36307 (N_36307,N_34105,N_35120);
nor U36308 (N_36308,N_34078,N_35478);
and U36309 (N_36309,N_35004,N_35364);
nor U36310 (N_36310,N_35485,N_34258);
and U36311 (N_36311,N_34873,N_34743);
nor U36312 (N_36312,N_35279,N_34934);
nor U36313 (N_36313,N_34463,N_35338);
nand U36314 (N_36314,N_34940,N_34472);
nor U36315 (N_36315,N_34751,N_35854);
nor U36316 (N_36316,N_35270,N_35288);
nand U36317 (N_36317,N_34850,N_35131);
xor U36318 (N_36318,N_34087,N_35548);
xnor U36319 (N_36319,N_35578,N_35278);
xnor U36320 (N_36320,N_35404,N_35046);
xor U36321 (N_36321,N_35630,N_34180);
nand U36322 (N_36322,N_34668,N_34470);
nor U36323 (N_36323,N_35464,N_35800);
and U36324 (N_36324,N_35090,N_34820);
nor U36325 (N_36325,N_34753,N_35223);
nand U36326 (N_36326,N_35813,N_35144);
or U36327 (N_36327,N_35425,N_34834);
nand U36328 (N_36328,N_34325,N_35302);
and U36329 (N_36329,N_35754,N_35146);
nand U36330 (N_36330,N_34052,N_34515);
nor U36331 (N_36331,N_34286,N_34335);
and U36332 (N_36332,N_34964,N_34359);
xor U36333 (N_36333,N_34801,N_34186);
and U36334 (N_36334,N_34252,N_35274);
nand U36335 (N_36335,N_35383,N_34611);
nand U36336 (N_36336,N_35300,N_34218);
xnor U36337 (N_36337,N_34949,N_34501);
nor U36338 (N_36338,N_35324,N_34533);
or U36339 (N_36339,N_35570,N_35409);
xnor U36340 (N_36340,N_34797,N_34879);
xnor U36341 (N_36341,N_34571,N_35238);
xnor U36342 (N_36342,N_35173,N_34320);
xnor U36343 (N_36343,N_34349,N_35138);
xnor U36344 (N_36344,N_34375,N_35342);
xnor U36345 (N_36345,N_35228,N_35344);
and U36346 (N_36346,N_34593,N_35062);
nand U36347 (N_36347,N_34516,N_34104);
and U36348 (N_36348,N_35687,N_35307);
and U36349 (N_36349,N_34453,N_35125);
and U36350 (N_36350,N_34003,N_35219);
or U36351 (N_36351,N_34344,N_35048);
and U36352 (N_36352,N_35027,N_34131);
nor U36353 (N_36353,N_35368,N_35549);
or U36354 (N_36354,N_34207,N_34389);
and U36355 (N_36355,N_34569,N_34237);
xnor U36356 (N_36356,N_34438,N_35977);
nand U36357 (N_36357,N_34974,N_34200);
or U36358 (N_36358,N_34446,N_34404);
nand U36359 (N_36359,N_35015,N_34348);
and U36360 (N_36360,N_35227,N_35799);
xor U36361 (N_36361,N_35001,N_34044);
or U36362 (N_36362,N_35634,N_35883);
nand U36363 (N_36363,N_35598,N_35410);
nand U36364 (N_36364,N_35982,N_34276);
and U36365 (N_36365,N_34304,N_35031);
and U36366 (N_36366,N_35139,N_34031);
xnor U36367 (N_36367,N_34998,N_35588);
xnor U36368 (N_36368,N_34788,N_35726);
and U36369 (N_36369,N_35876,N_34632);
or U36370 (N_36370,N_35632,N_34269);
and U36371 (N_36371,N_35862,N_35658);
and U36372 (N_36372,N_34785,N_35795);
nand U36373 (N_36373,N_34464,N_35565);
or U36374 (N_36374,N_34576,N_34159);
or U36375 (N_36375,N_35691,N_34263);
and U36376 (N_36376,N_34461,N_35163);
and U36377 (N_36377,N_35825,N_35772);
nand U36378 (N_36378,N_35816,N_35024);
nor U36379 (N_36379,N_34532,N_34926);
and U36380 (N_36380,N_34117,N_35685);
and U36381 (N_36381,N_35369,N_34083);
xnor U36382 (N_36382,N_34969,N_35128);
nor U36383 (N_36383,N_35092,N_35991);
nor U36384 (N_36384,N_34589,N_34605);
nor U36385 (N_36385,N_35820,N_35418);
nor U36386 (N_36386,N_35343,N_34468);
nand U36387 (N_36387,N_35656,N_34480);
xnor U36388 (N_36388,N_35003,N_34965);
nor U36389 (N_36389,N_34203,N_35280);
and U36390 (N_36390,N_35787,N_34002);
nand U36391 (N_36391,N_35692,N_34529);
xor U36392 (N_36392,N_35665,N_35882);
nor U36393 (N_36393,N_34329,N_34888);
and U36394 (N_36394,N_34805,N_35094);
nand U36395 (N_36395,N_35980,N_35849);
or U36396 (N_36396,N_35901,N_34275);
and U36397 (N_36397,N_34917,N_34923);
or U36398 (N_36398,N_34419,N_34007);
xnor U36399 (N_36399,N_35791,N_34715);
nand U36400 (N_36400,N_35190,N_34481);
and U36401 (N_36401,N_34782,N_35328);
nor U36402 (N_36402,N_34685,N_35210);
nand U36403 (N_36403,N_35058,N_35311);
or U36404 (N_36404,N_35164,N_34337);
or U36405 (N_36405,N_35042,N_35401);
nor U36406 (N_36406,N_35871,N_35487);
xnor U36407 (N_36407,N_35291,N_35783);
nand U36408 (N_36408,N_35645,N_34866);
or U36409 (N_36409,N_35616,N_34748);
nand U36410 (N_36410,N_34971,N_35309);
nor U36411 (N_36411,N_35075,N_35474);
and U36412 (N_36412,N_35814,N_35893);
nand U36413 (N_36413,N_34085,N_34524);
or U36414 (N_36414,N_35167,N_34637);
nor U36415 (N_36415,N_34553,N_34695);
nor U36416 (N_36416,N_35486,N_35319);
or U36417 (N_36417,N_35230,N_34089);
nand U36418 (N_36418,N_34765,N_34832);
or U36419 (N_36419,N_35379,N_35175);
xnor U36420 (N_36420,N_34151,N_34093);
or U36421 (N_36421,N_35872,N_34408);
nand U36422 (N_36422,N_34578,N_34792);
xnor U36423 (N_36423,N_35108,N_34013);
and U36424 (N_36424,N_35833,N_34381);
and U36425 (N_36425,N_35736,N_35403);
nor U36426 (N_36426,N_35930,N_34508);
or U36427 (N_36427,N_34176,N_34517);
xnor U36428 (N_36428,N_34670,N_35941);
or U36429 (N_36429,N_35635,N_34664);
nor U36430 (N_36430,N_34960,N_35107);
nor U36431 (N_36431,N_35211,N_34299);
or U36432 (N_36432,N_34821,N_35022);
nor U36433 (N_36433,N_35506,N_34750);
and U36434 (N_36434,N_35061,N_34811);
xnor U36435 (N_36435,N_35336,N_34865);
nor U36436 (N_36436,N_34787,N_35602);
nor U36437 (N_36437,N_34473,N_35356);
nand U36438 (N_36438,N_34420,N_34746);
or U36439 (N_36439,N_35892,N_35788);
xor U36440 (N_36440,N_35448,N_34247);
nand U36441 (N_36441,N_34745,N_34635);
nand U36442 (N_36442,N_34565,N_34580);
nand U36443 (N_36443,N_34096,N_35569);
or U36444 (N_36444,N_35166,N_35766);
and U36445 (N_36445,N_35574,N_35381);
and U36446 (N_36446,N_35426,N_34362);
nor U36447 (N_36447,N_34573,N_35249);
xnor U36448 (N_36448,N_34671,N_34262);
and U36449 (N_36449,N_35841,N_34531);
or U36450 (N_36450,N_35064,N_34416);
or U36451 (N_36451,N_35266,N_35386);
and U36452 (N_36452,N_34026,N_35763);
nand U36453 (N_36453,N_35057,N_34768);
xnor U36454 (N_36454,N_34351,N_34165);
or U36455 (N_36455,N_35563,N_34040);
or U36456 (N_36456,N_35625,N_34659);
nand U36457 (N_36457,N_35020,N_35696);
xor U36458 (N_36458,N_35908,N_35520);
and U36459 (N_36459,N_34068,N_34795);
nor U36460 (N_36460,N_34377,N_34380);
or U36461 (N_36461,N_34599,N_34883);
nand U36462 (N_36462,N_35301,N_34292);
nor U36463 (N_36463,N_34265,N_34164);
nor U36464 (N_36464,N_34301,N_35053);
nor U36465 (N_36465,N_35670,N_35637);
and U36466 (N_36466,N_34364,N_35148);
nor U36467 (N_36467,N_34597,N_34126);
nand U36468 (N_36468,N_34608,N_35367);
nand U36469 (N_36469,N_35781,N_35910);
or U36470 (N_36470,N_35750,N_34931);
or U36471 (N_36471,N_34963,N_35699);
and U36472 (N_36472,N_34112,N_34474);
nand U36473 (N_36473,N_35303,N_34133);
nor U36474 (N_36474,N_35926,N_34168);
nand U36475 (N_36475,N_34179,N_35944);
nor U36476 (N_36476,N_35584,N_34343);
and U36477 (N_36477,N_34741,N_34012);
nand U36478 (N_36478,N_35536,N_35021);
or U36479 (N_36479,N_35579,N_34141);
nor U36480 (N_36480,N_35081,N_34488);
and U36481 (N_36481,N_35896,N_34617);
or U36482 (N_36482,N_34211,N_34283);
and U36483 (N_36483,N_34273,N_34298);
nand U36484 (N_36484,N_35582,N_35332);
or U36485 (N_36485,N_34210,N_35613);
nand U36486 (N_36486,N_34413,N_35522);
xor U36487 (N_36487,N_34946,N_35355);
or U36488 (N_36488,N_34502,N_35151);
and U36489 (N_36489,N_34303,N_34628);
xor U36490 (N_36490,N_34392,N_34759);
nand U36491 (N_36491,N_35116,N_34279);
or U36492 (N_36492,N_35577,N_34763);
xnor U36493 (N_36493,N_35420,N_34574);
nand U36494 (N_36494,N_35087,N_35032);
and U36495 (N_36495,N_34001,N_35861);
nor U36496 (N_36496,N_35188,N_35215);
or U36497 (N_36497,N_35231,N_34885);
and U36498 (N_36498,N_35056,N_35725);
nor U36499 (N_36499,N_35203,N_34188);
nor U36500 (N_36500,N_34288,N_35547);
and U36501 (N_36501,N_35170,N_35468);
and U36502 (N_36502,N_34147,N_35212);
xor U36503 (N_36503,N_35427,N_35546);
nand U36504 (N_36504,N_35205,N_34491);
xnor U36505 (N_36505,N_35761,N_35731);
xnor U36506 (N_36506,N_35976,N_35664);
or U36507 (N_36507,N_35823,N_35667);
xor U36508 (N_36508,N_34324,N_34062);
nand U36509 (N_36509,N_35243,N_35600);
and U36510 (N_36510,N_35654,N_34010);
or U36511 (N_36511,N_34084,N_35202);
xor U36512 (N_36512,N_35794,N_35285);
xnor U36513 (N_36513,N_35599,N_34858);
nor U36514 (N_36514,N_34227,N_35217);
or U36515 (N_36515,N_35995,N_35277);
and U36516 (N_36516,N_35540,N_35875);
or U36517 (N_36517,N_35491,N_34898);
or U36518 (N_36518,N_35097,N_34967);
nor U36519 (N_36519,N_35990,N_35551);
xnor U36520 (N_36520,N_35585,N_34997);
or U36521 (N_36521,N_35887,N_34991);
and U36522 (N_36522,N_35961,N_35535);
or U36523 (N_36523,N_35432,N_35943);
xor U36524 (N_36524,N_34213,N_34734);
nand U36525 (N_36525,N_35847,N_35130);
nor U36526 (N_36526,N_35934,N_34278);
or U36527 (N_36527,N_34889,N_34248);
nor U36528 (N_36528,N_34914,N_35708);
and U36529 (N_36529,N_35103,N_34581);
and U36530 (N_36530,N_34193,N_34657);
and U36531 (N_36531,N_35242,N_34241);
and U36532 (N_36532,N_34030,N_35119);
or U36533 (N_36533,N_34739,N_35837);
nand U36534 (N_36534,N_34397,N_34017);
nor U36535 (N_36535,N_35538,N_34092);
nor U36536 (N_36536,N_34577,N_34958);
nor U36537 (N_36537,N_34895,N_34231);
xor U36538 (N_36538,N_34459,N_34713);
and U36539 (N_36539,N_35523,N_34194);
nor U36540 (N_36540,N_34627,N_35880);
or U36541 (N_36541,N_35895,N_34857);
or U36542 (N_36542,N_34477,N_34287);
nor U36543 (N_36543,N_35245,N_35070);
and U36544 (N_36544,N_34448,N_34548);
xor U36545 (N_36545,N_35575,N_35686);
and U36546 (N_36546,N_35100,N_34881);
nor U36547 (N_36547,N_34161,N_35631);
or U36548 (N_36548,N_35937,N_34988);
and U36549 (N_36549,N_34048,N_34757);
and U36550 (N_36550,N_34645,N_35994);
nand U36551 (N_36551,N_34567,N_34692);
nor U36552 (N_36552,N_35594,N_34874);
nand U36553 (N_36553,N_34846,N_34992);
and U36554 (N_36554,N_35917,N_35159);
nand U36555 (N_36555,N_34973,N_34527);
nor U36556 (N_36556,N_35127,N_35534);
xor U36557 (N_36557,N_34290,N_35374);
and U36558 (N_36558,N_35191,N_35251);
and U36559 (N_36559,N_35453,N_34910);
and U36560 (N_36560,N_34466,N_35907);
nor U36561 (N_36561,N_34826,N_35711);
and U36562 (N_36562,N_34099,N_34394);
nor U36563 (N_36563,N_34854,N_34274);
nand U36564 (N_36564,N_34844,N_35510);
or U36565 (N_36565,N_35950,N_35790);
and U36566 (N_36566,N_34830,N_34475);
nor U36567 (N_36567,N_35466,N_34189);
or U36568 (N_36568,N_35394,N_35689);
and U36569 (N_36569,N_35697,N_35255);
xor U36570 (N_36570,N_35463,N_35079);
nand U36571 (N_36571,N_34733,N_35380);
nand U36572 (N_36572,N_34868,N_34253);
nand U36573 (N_36573,N_34676,N_35469);
nor U36574 (N_36574,N_34035,N_34405);
nor U36575 (N_36575,N_35743,N_35568);
nor U36576 (N_36576,N_35564,N_35450);
xnor U36577 (N_36577,N_34434,N_35158);
xnor U36578 (N_36578,N_34361,N_34555);
xor U36579 (N_36579,N_34018,N_34812);
or U36580 (N_36580,N_34050,N_34357);
or U36581 (N_36581,N_34521,N_34029);
nand U36582 (N_36582,N_35636,N_34884);
nand U36583 (N_36583,N_34284,N_35679);
or U36584 (N_36584,N_34526,N_35218);
and U36585 (N_36585,N_34086,N_34485);
and U36586 (N_36586,N_35089,N_35915);
and U36587 (N_36587,N_35718,N_35573);
nand U36588 (N_36588,N_35605,N_34444);
or U36589 (N_36589,N_35516,N_34675);
and U36590 (N_36590,N_34839,N_34882);
nor U36591 (N_36591,N_34153,N_35499);
and U36592 (N_36592,N_35292,N_35392);
nor U36593 (N_36593,N_35268,N_35610);
and U36594 (N_36594,N_35359,N_34615);
and U36595 (N_36595,N_35229,N_34729);
nor U36596 (N_36596,N_34842,N_35993);
nor U36597 (N_36597,N_34662,N_35345);
and U36598 (N_36598,N_35615,N_34383);
xor U36599 (N_36599,N_34513,N_35715);
xor U36600 (N_36600,N_34170,N_34936);
nor U36601 (N_36601,N_34201,N_34223);
xnor U36602 (N_36602,N_34316,N_34633);
nor U36603 (N_36603,N_35870,N_35258);
and U36604 (N_36604,N_35315,N_35063);
or U36605 (N_36605,N_35406,N_34022);
xor U36606 (N_36606,N_35545,N_34755);
and U36607 (N_36607,N_35804,N_35254);
nand U36608 (N_36608,N_35477,N_34330);
nand U36609 (N_36609,N_34648,N_34204);
or U36610 (N_36610,N_35093,N_35886);
and U36611 (N_36611,N_35348,N_34697);
or U36612 (N_36612,N_35484,N_35957);
nor U36613 (N_36613,N_35742,N_34075);
nand U36614 (N_36614,N_34073,N_34452);
or U36615 (N_36615,N_34875,N_35051);
or U36616 (N_36616,N_34712,N_34702);
xor U36617 (N_36617,N_35527,N_35856);
nand U36618 (N_36618,N_35050,N_34878);
nor U36619 (N_36619,N_35624,N_35192);
nand U36620 (N_36620,N_35422,N_34827);
xnor U36621 (N_36621,N_34257,N_34572);
and U36622 (N_36622,N_34945,N_35289);
nor U36623 (N_36623,N_34953,N_34767);
and U36624 (N_36624,N_34825,N_34735);
or U36625 (N_36625,N_34398,N_34326);
or U36626 (N_36626,N_35357,N_34064);
nor U36627 (N_36627,N_35135,N_35701);
nor U36628 (N_36628,N_35553,N_35150);
or U36629 (N_36629,N_35467,N_35706);
or U36630 (N_36630,N_34579,N_34220);
xnor U36631 (N_36631,N_35999,N_35295);
nor U36632 (N_36632,N_35038,N_35700);
xnor U36633 (N_36633,N_34837,N_35298);
xnor U36634 (N_36634,N_35331,N_34722);
and U36635 (N_36635,N_34817,N_35539);
and U36636 (N_36636,N_34863,N_34177);
or U36637 (N_36637,N_35648,N_35784);
nor U36638 (N_36638,N_34609,N_34495);
xnor U36639 (N_36639,N_35532,N_35076);
and U36640 (N_36640,N_35060,N_34756);
nand U36641 (N_36641,N_35716,N_35197);
nor U36642 (N_36642,N_35684,N_35931);
or U36643 (N_36643,N_35873,N_35209);
xor U36644 (N_36644,N_34120,N_35657);
nor U36645 (N_36645,N_35898,N_35177);
or U36646 (N_36646,N_34025,N_35017);
and U36647 (N_36647,N_35497,N_35376);
xnor U36648 (N_36648,N_35314,N_35720);
or U36649 (N_36649,N_35807,N_34036);
nand U36650 (N_36650,N_35928,N_34217);
xor U36651 (N_36651,N_35970,N_34941);
nor U36652 (N_36652,N_34197,N_34700);
and U36653 (N_36653,N_35502,N_34229);
and U36654 (N_36654,N_34810,N_34861);
and U36655 (N_36655,N_35912,N_34816);
nand U36656 (N_36656,N_35495,N_34315);
and U36657 (N_36657,N_35713,N_35236);
xor U36658 (N_36658,N_35932,N_35511);
or U36659 (N_36659,N_34432,N_35972);
xor U36660 (N_36660,N_35358,N_35489);
nor U36661 (N_36661,N_34803,N_35719);
xor U36662 (N_36662,N_34557,N_35734);
or U36663 (N_36663,N_35618,N_35433);
xnor U36664 (N_36664,N_35439,N_35517);
or U36665 (N_36665,N_34192,N_34725);
xnor U36666 (N_36666,N_34760,N_34019);
nor U36667 (N_36667,N_34431,N_35843);
and U36668 (N_36668,N_34118,N_34731);
nand U36669 (N_36669,N_35399,N_34592);
and U36670 (N_36670,N_35316,N_35693);
and U36671 (N_36671,N_34975,N_34869);
nor U36672 (N_36672,N_35145,N_34616);
and U36673 (N_36673,N_34968,N_35341);
xnor U36674 (N_36674,N_35330,N_34994);
or U36675 (N_36675,N_35507,N_34566);
or U36676 (N_36676,N_34758,N_35846);
and U36677 (N_36677,N_34492,N_34687);
or U36678 (N_36678,N_34439,N_35008);
nor U36679 (N_36679,N_34033,N_35782);
nand U36680 (N_36680,N_35889,N_34423);
nand U36681 (N_36681,N_34249,N_34921);
or U36682 (N_36682,N_34268,N_34196);
and U36683 (N_36683,N_35043,N_34856);
nand U36684 (N_36684,N_34629,N_34396);
and U36685 (N_36685,N_35327,N_35552);
or U36686 (N_36686,N_34649,N_35617);
nand U36687 (N_36687,N_35010,N_35828);
nand U36688 (N_36688,N_34644,N_35325);
nand U36689 (N_36689,N_34261,N_34129);
xnor U36690 (N_36690,N_35451,N_34415);
nand U36691 (N_36691,N_34904,N_34157);
or U36692 (N_36692,N_35030,N_35810);
nand U36693 (N_36693,N_35112,N_34519);
nor U36694 (N_36694,N_35952,N_35842);
nor U36695 (N_36695,N_34536,N_35034);
nor U36696 (N_36696,N_34647,N_35962);
or U36697 (N_36697,N_34020,N_34450);
or U36698 (N_36698,N_34808,N_34836);
or U36699 (N_36699,N_34943,N_35971);
and U36700 (N_36700,N_35537,N_35333);
nand U36701 (N_36701,N_34006,N_35924);
xor U36702 (N_36702,N_35040,N_34198);
nor U36703 (N_36703,N_34905,N_34455);
xor U36704 (N_36704,N_35710,N_34244);
nand U36705 (N_36705,N_34736,N_34267);
xnor U36706 (N_36706,N_34000,N_35262);
xor U36707 (N_36707,N_35365,N_34063);
nand U36708 (N_36708,N_34672,N_34824);
xnor U36709 (N_36709,N_34132,N_35493);
or U36710 (N_36710,N_34308,N_34728);
nand U36711 (N_36711,N_35709,N_34191);
or U36712 (N_36712,N_34312,N_35666);
xor U36713 (N_36713,N_35543,N_35777);
or U36714 (N_36714,N_35396,N_35916);
xor U36715 (N_36715,N_35942,N_35235);
nor U36716 (N_36716,N_34876,N_35390);
nand U36717 (N_36717,N_35818,N_34862);
or U36718 (N_36718,N_35819,N_34665);
and U36719 (N_36719,N_35593,N_35601);
nor U36720 (N_36720,N_35434,N_35680);
and U36721 (N_36721,N_35059,N_34221);
or U36722 (N_36722,N_35555,N_34638);
nand U36723 (N_36723,N_34802,N_34770);
and U36724 (N_36724,N_35371,N_34183);
or U36725 (N_36725,N_34228,N_34518);
xnor U36726 (N_36726,N_34390,N_35969);
or U36727 (N_36727,N_34766,N_34109);
nor U36728 (N_36728,N_35978,N_34422);
nand U36729 (N_36729,N_34095,N_35018);
xor U36730 (N_36730,N_35501,N_35992);
xor U36731 (N_36731,N_34673,N_34710);
nor U36732 (N_36732,N_35728,N_34807);
nand U36733 (N_36733,N_35023,N_35581);
nand U36734 (N_36734,N_35361,N_34174);
nor U36735 (N_36735,N_34978,N_34103);
and U36736 (N_36736,N_34245,N_34441);
nand U36737 (N_36737,N_34623,N_34373);
or U36738 (N_36738,N_35554,N_34386);
and U36739 (N_36739,N_34679,N_35524);
nand U36740 (N_36740,N_35429,N_35877);
or U36741 (N_36741,N_34134,N_34071);
and U36742 (N_36742,N_34915,N_34838);
xnor U36743 (N_36743,N_34514,N_35294);
nor U36744 (N_36744,N_34822,N_34901);
or U36745 (N_36745,N_35216,N_35113);
nor U36746 (N_36746,N_34640,N_34345);
nand U36747 (N_36747,N_35933,N_35471);
nand U36748 (N_36748,N_35424,N_35629);
nor U36749 (N_36749,N_35049,N_35829);
and U36750 (N_36750,N_34372,N_35282);
and U36751 (N_36751,N_35753,N_34903);
or U36752 (N_36752,N_34696,N_34594);
or U36753 (N_36753,N_35488,N_34922);
nand U36754 (N_36754,N_34425,N_35247);
nor U36755 (N_36755,N_35360,N_35457);
nor U36756 (N_36756,N_34538,N_35678);
or U36757 (N_36757,N_34976,N_34355);
xor U36758 (N_36758,N_34090,N_34009);
xor U36759 (N_36759,N_35735,N_35835);
nor U36760 (N_36760,N_34149,N_35595);
xor U36761 (N_36761,N_35224,N_34238);
nand U36762 (N_36762,N_35925,N_34591);
nand U36763 (N_36763,N_34789,N_34979);
nor U36764 (N_36764,N_35157,N_34754);
and U36765 (N_36765,N_35659,N_34851);
nor U36766 (N_36766,N_35421,N_34049);
and U36767 (N_36767,N_34145,N_34369);
nand U36768 (N_36768,N_34784,N_34401);
or U36769 (N_36769,N_35161,N_34534);
and U36770 (N_36770,N_35456,N_34016);
or U36771 (N_36771,N_34871,N_35452);
xor U36772 (N_36772,N_35340,N_35029);
nand U36773 (N_36773,N_34256,N_34102);
or U36774 (N_36774,N_35868,N_34442);
and U36775 (N_36775,N_35162,N_34272);
or U36776 (N_36776,N_34719,N_34853);
nor U36777 (N_36777,N_35458,N_35673);
or U36778 (N_36778,N_34094,N_34899);
nand U36779 (N_36779,N_34996,N_35948);
nand U36780 (N_36780,N_35669,N_34309);
nor U36781 (N_36781,N_35096,N_35102);
xnor U36782 (N_36782,N_34379,N_34277);
nor U36783 (N_36783,N_35156,N_35821);
xnor U36784 (N_36784,N_35620,N_35414);
or U36785 (N_36785,N_34296,N_34507);
nor U36786 (N_36786,N_34015,N_35780);
xnor U36787 (N_36787,N_34732,N_34800);
xnor U36788 (N_36788,N_35073,N_34136);
nor U36789 (N_36789,N_35759,N_34613);
or U36790 (N_36790,N_35681,N_35416);
and U36791 (N_36791,N_34716,N_35639);
nor U36792 (N_36792,N_35402,N_35640);
or U36793 (N_36793,N_34427,N_34260);
nor U36794 (N_36794,N_34115,N_35375);
or U36795 (N_36795,N_35308,N_34039);
and U36796 (N_36796,N_34230,N_35541);
nor U36797 (N_36797,N_35012,N_35239);
and U36798 (N_36798,N_35652,N_34699);
xor U36799 (N_36799,N_34171,N_35461);
xnor U36800 (N_36800,N_34535,N_34652);
or U36801 (N_36801,N_35252,N_34704);
or U36802 (N_36802,N_35739,N_34327);
nor U36803 (N_36803,N_34511,N_34747);
or U36804 (N_36804,N_35698,N_35111);
and U36805 (N_36805,N_34781,N_35967);
xnor U36806 (N_36806,N_35649,N_34418);
nor U36807 (N_36807,N_34323,N_35606);
and U36808 (N_36808,N_34607,N_34582);
nor U36809 (N_36809,N_35088,N_34776);
xnor U36810 (N_36810,N_34908,N_35014);
nand U36811 (N_36811,N_35722,N_34155);
nor U36812 (N_36812,N_34774,N_35505);
and U36813 (N_36813,N_35321,N_34127);
nor U36814 (N_36814,N_35529,N_34332);
or U36815 (N_36815,N_35774,N_35436);
nand U36816 (N_36816,N_35147,N_35470);
xnor U36817 (N_36817,N_34547,N_35938);
nand U36818 (N_36818,N_35936,N_34989);
xnor U36819 (N_36819,N_34980,N_35848);
xnor U36820 (N_36820,N_35996,N_34313);
and U36821 (N_36821,N_35914,N_35660);
nor U36822 (N_36822,N_35504,N_34458);
and U36823 (N_36823,N_34650,N_34651);
and U36824 (N_36824,N_35515,N_34688);
or U36825 (N_36825,N_35830,N_34457);
nand U36826 (N_36826,N_35172,N_35981);
nor U36827 (N_36827,N_34429,N_34551);
or U36828 (N_36828,N_35815,N_34769);
and U36829 (N_36829,N_35494,N_35248);
xnor U36830 (N_36830,N_34880,N_34199);
xor U36831 (N_36831,N_34835,N_35084);
nor U36832 (N_36832,N_34913,N_35729);
or U36833 (N_36833,N_35136,N_35153);
xor U36834 (N_36834,N_34081,N_34338);
nor U36835 (N_36835,N_35446,N_34643);
nand U36836 (N_36836,N_35627,N_34291);
and U36837 (N_36837,N_35069,N_34356);
or U36838 (N_36838,N_34264,N_35480);
nand U36839 (N_36839,N_35793,N_35778);
xor U36840 (N_36840,N_34714,N_35299);
xnor U36841 (N_36841,N_35036,N_34384);
xor U36842 (N_36842,N_35193,N_34724);
xnor U36843 (N_36843,N_35576,N_35769);
nand U36844 (N_36844,N_34786,N_35745);
and U36845 (N_36845,N_35738,N_35503);
and U36846 (N_36846,N_34140,N_34282);
or U36847 (N_36847,N_34166,N_34870);
xor U36848 (N_36848,N_34437,N_35621);
nor U36849 (N_36849,N_35067,N_35281);
or U36850 (N_36850,N_34110,N_34925);
nand U36851 (N_36851,N_34783,N_34606);
nand U36852 (N_36852,N_34912,N_34537);
and U36853 (N_36853,N_35373,N_35306);
or U36854 (N_36854,N_35905,N_34409);
xnor U36855 (N_36855,N_34962,N_35222);
nand U36856 (N_36856,N_35521,N_35155);
nor U36857 (N_36857,N_34545,N_34041);
and U36858 (N_36858,N_35586,N_35785);
nor U36859 (N_36859,N_35378,N_35909);
nand U36860 (N_36860,N_34970,N_35808);
or U36861 (N_36861,N_34391,N_34447);
nor U36862 (N_36862,N_34814,N_35979);
or U36863 (N_36863,N_34482,N_34663);
nand U36864 (N_36864,N_34496,N_35603);
or U36865 (N_36865,N_34603,N_34622);
nand U36866 (N_36866,N_34944,N_35105);
xnor U36867 (N_36867,N_34122,N_34321);
nand U36868 (N_36868,N_35168,N_34726);
and U36869 (N_36869,N_35607,N_34242);
or U36870 (N_36870,N_35662,N_35115);
xnor U36871 (N_36871,N_34942,N_34681);
nand U36872 (N_36872,N_34539,N_34499);
nor U36873 (N_36873,N_35196,N_34341);
and U36874 (N_36874,N_35587,N_35518);
nand U36875 (N_36875,N_34005,N_35250);
and U36876 (N_36876,N_34138,N_34051);
xor U36877 (N_36877,N_35305,N_35276);
xnor U36878 (N_36878,N_34004,N_34568);
and U36879 (N_36879,N_34723,N_34354);
nor U36880 (N_36880,N_35956,N_35137);
nor U36881 (N_36881,N_35182,N_34698);
or U36882 (N_36882,N_34144,N_35747);
nand U36883 (N_36883,N_34119,N_34897);
nor U36884 (N_36884,N_35435,N_35695);
and U36885 (N_36885,N_34428,N_34307);
nor U36886 (N_36886,N_35413,N_34520);
xor U36887 (N_36887,N_35121,N_35855);
nand U36888 (N_36888,N_34121,N_34806);
nor U36889 (N_36889,N_34175,N_35233);
or U36890 (N_36890,N_35965,N_34999);
nor U36891 (N_36891,N_35109,N_35183);
and U36892 (N_36892,N_35591,N_35339);
or U36893 (N_36893,N_34951,N_34525);
or U36894 (N_36894,N_34933,N_35922);
nor U36895 (N_36895,N_34646,N_35562);
nand U36896 (N_36896,N_34185,N_34703);
nand U36897 (N_36897,N_34993,N_34456);
and U36898 (N_36898,N_34243,N_34106);
nand U36899 (N_36899,N_35326,N_35397);
nor U36900 (N_36900,N_34828,N_34959);
and U36901 (N_36901,N_35597,N_35296);
xor U36902 (N_36902,N_35385,N_35604);
xnor U36903 (N_36903,N_35443,N_34620);
nand U36904 (N_36904,N_35498,N_34246);
or U36905 (N_36905,N_35612,N_34173);
nor U36906 (N_36906,N_35310,N_35732);
nor U36907 (N_36907,N_35186,N_34224);
or U36908 (N_36908,N_34074,N_34721);
and U36909 (N_36909,N_35496,N_35959);
or U36910 (N_36910,N_35313,N_34293);
and U36911 (N_36911,N_35572,N_34641);
nand U36912 (N_36912,N_35964,N_35016);
nand U36913 (N_36913,N_34417,N_34154);
or U36914 (N_36914,N_34720,N_35335);
nand U36915 (N_36915,N_35920,N_34388);
and U36916 (N_36916,N_35966,N_34318);
nor U36917 (N_36917,N_35939,N_34711);
nor U36918 (N_36918,N_34319,N_34845);
and U36919 (N_36919,N_35045,N_34476);
xor U36920 (N_36920,N_35884,N_35449);
nor U36921 (N_36921,N_35921,N_35005);
and U36922 (N_36922,N_35746,N_34302);
nor U36923 (N_36923,N_34604,N_35377);
nor U36924 (N_36924,N_35779,N_34619);
nand U36925 (N_36925,N_34146,N_34008);
nor U36926 (N_36926,N_35101,N_35838);
nand U36927 (N_36927,N_34669,N_34387);
xnor U36928 (N_36928,N_34550,N_35985);
and U36929 (N_36929,N_34047,N_35556);
nand U36930 (N_36930,N_34563,N_35514);
xor U36931 (N_36931,N_34057,N_34069);
nor U36932 (N_36932,N_35283,N_34552);
xor U36933 (N_36933,N_35455,N_34584);
and U36934 (N_36934,N_34123,N_35444);
xnor U36935 (N_36935,N_35864,N_34655);
or U36936 (N_36936,N_34546,N_34225);
xnor U36937 (N_36937,N_35651,N_35269);
xor U36938 (N_36938,N_34829,N_35646);
nand U36939 (N_36939,N_34775,N_35622);
nand U36940 (N_36940,N_35560,N_35033);
and U36941 (N_36941,N_34503,N_34346);
nor U36942 (N_36942,N_35187,N_35304);
and U36943 (N_36943,N_35968,N_35185);
and U36944 (N_36944,N_34077,N_35583);
nor U36945 (N_36945,N_35259,N_35297);
or U36946 (N_36946,N_34100,N_34266);
and U36947 (N_36947,N_34128,N_35857);
or U36948 (N_36948,N_35287,N_34076);
and U36949 (N_36949,N_35272,N_34440);
xnor U36950 (N_36950,N_35389,N_35724);
or U36951 (N_36951,N_35671,N_35419);
and U36952 (N_36952,N_34281,N_35817);
and U36953 (N_36953,N_34460,N_35797);
xnor U36954 (N_36954,N_34831,N_35803);
nor U36955 (N_36955,N_35960,N_34935);
xnor U36956 (N_36956,N_34340,N_35655);
and U36957 (N_36957,N_34586,N_34414);
nor U36958 (N_36958,N_35674,N_34209);
xor U36959 (N_36959,N_35946,N_34583);
nand U36960 (N_36960,N_34407,N_34554);
or U36961 (N_36961,N_34066,N_35460);
xor U36962 (N_36962,N_35650,N_34961);
xor U36963 (N_36963,N_35037,N_35041);
and U36964 (N_36964,N_35859,N_35232);
or U36965 (N_36965,N_34435,N_34426);
xnor U36966 (N_36966,N_34350,N_35149);
or U36967 (N_36967,N_34045,N_35214);
xnor U36968 (N_36968,N_34680,N_34859);
nor U36969 (N_36969,N_35221,N_35104);
xnor U36970 (N_36970,N_35025,N_35318);
nand U36971 (N_36971,N_35482,N_35775);
or U36972 (N_36972,N_35741,N_34382);
nand U36973 (N_36973,N_34150,N_35098);
or U36974 (N_36974,N_35500,N_34596);
and U36975 (N_36975,N_35512,N_35206);
or U36976 (N_36976,N_35832,N_35899);
or U36977 (N_36977,N_35391,N_34841);
nand U36978 (N_36978,N_35290,N_35888);
and U36979 (N_36979,N_35065,N_35181);
or U36980 (N_36980,N_34181,N_35508);
and U36981 (N_36981,N_35850,N_34602);
nor U36982 (N_36982,N_34162,N_35764);
or U36983 (N_36983,N_34226,N_35776);
nor U36984 (N_36984,N_34955,N_34114);
nor U36985 (N_36985,N_35085,N_35071);
xnor U36986 (N_36986,N_35704,N_35473);
and U36987 (N_36987,N_34624,N_35160);
nor U36988 (N_36988,N_34799,N_35812);
and U36989 (N_36989,N_34985,N_35066);
and U36990 (N_36990,N_35571,N_34986);
nor U36991 (N_36991,N_35902,N_34160);
nor U36992 (N_36992,N_35002,N_35525);
and U36993 (N_36993,N_35550,N_35643);
nor U36994 (N_36994,N_34771,N_34395);
xor U36995 (N_36995,N_35405,N_35476);
or U36996 (N_36996,N_34813,N_34215);
and U36997 (N_36997,N_35035,N_35557);
xnor U36998 (N_36998,N_35744,N_35953);
nor U36999 (N_36999,N_34542,N_34693);
nor U37000 (N_37000,N_34141,N_35420);
or U37001 (N_37001,N_34246,N_34543);
nand U37002 (N_37002,N_35924,N_35049);
or U37003 (N_37003,N_35881,N_35133);
nand U37004 (N_37004,N_34538,N_35227);
nand U37005 (N_37005,N_34112,N_35208);
xnor U37006 (N_37006,N_35255,N_35915);
and U37007 (N_37007,N_34023,N_34017);
xor U37008 (N_37008,N_35552,N_35240);
xor U37009 (N_37009,N_35819,N_35934);
nor U37010 (N_37010,N_34348,N_35708);
nand U37011 (N_37011,N_35318,N_34807);
nand U37012 (N_37012,N_34609,N_35934);
xnor U37013 (N_37013,N_34569,N_34880);
nor U37014 (N_37014,N_34852,N_34681);
xor U37015 (N_37015,N_35140,N_34257);
nor U37016 (N_37016,N_35171,N_35631);
nand U37017 (N_37017,N_35237,N_34993);
or U37018 (N_37018,N_34831,N_35031);
xnor U37019 (N_37019,N_34035,N_34624);
and U37020 (N_37020,N_34181,N_34948);
or U37021 (N_37021,N_35862,N_35071);
xnor U37022 (N_37022,N_35051,N_35602);
and U37023 (N_37023,N_34645,N_35988);
nand U37024 (N_37024,N_34219,N_34982);
or U37025 (N_37025,N_34463,N_34789);
xnor U37026 (N_37026,N_35620,N_34268);
nand U37027 (N_37027,N_34029,N_35685);
xor U37028 (N_37028,N_35562,N_35051);
nor U37029 (N_37029,N_34609,N_34341);
and U37030 (N_37030,N_34615,N_35658);
xnor U37031 (N_37031,N_35048,N_35882);
xor U37032 (N_37032,N_35134,N_34596);
or U37033 (N_37033,N_35803,N_34580);
nand U37034 (N_37034,N_35258,N_35445);
nand U37035 (N_37035,N_34194,N_35731);
xor U37036 (N_37036,N_34928,N_35153);
and U37037 (N_37037,N_35659,N_34746);
or U37038 (N_37038,N_35167,N_35605);
and U37039 (N_37039,N_35712,N_34991);
nor U37040 (N_37040,N_35544,N_35483);
xor U37041 (N_37041,N_34704,N_35706);
and U37042 (N_37042,N_35508,N_34967);
nand U37043 (N_37043,N_35364,N_35147);
and U37044 (N_37044,N_34363,N_35406);
nor U37045 (N_37045,N_35640,N_34248);
and U37046 (N_37046,N_35897,N_34498);
nor U37047 (N_37047,N_34088,N_34917);
or U37048 (N_37048,N_35203,N_35578);
or U37049 (N_37049,N_35553,N_35817);
nor U37050 (N_37050,N_34182,N_34070);
xnor U37051 (N_37051,N_34882,N_35878);
nor U37052 (N_37052,N_34551,N_35580);
nor U37053 (N_37053,N_34774,N_35534);
or U37054 (N_37054,N_35977,N_35210);
xor U37055 (N_37055,N_35318,N_35226);
or U37056 (N_37056,N_35282,N_34821);
nand U37057 (N_37057,N_34968,N_34205);
nor U37058 (N_37058,N_35423,N_34298);
xor U37059 (N_37059,N_35384,N_34906);
nand U37060 (N_37060,N_35045,N_34027);
nand U37061 (N_37061,N_34511,N_34609);
nor U37062 (N_37062,N_34216,N_34168);
xnor U37063 (N_37063,N_35884,N_34863);
xor U37064 (N_37064,N_34230,N_35912);
xor U37065 (N_37065,N_35354,N_34113);
xnor U37066 (N_37066,N_34369,N_34499);
and U37067 (N_37067,N_35138,N_35145);
nor U37068 (N_37068,N_34557,N_34299);
and U37069 (N_37069,N_34497,N_34177);
xor U37070 (N_37070,N_34366,N_35909);
xor U37071 (N_37071,N_34713,N_35181);
and U37072 (N_37072,N_35017,N_35172);
or U37073 (N_37073,N_34424,N_34023);
or U37074 (N_37074,N_35604,N_34146);
and U37075 (N_37075,N_35316,N_34095);
xor U37076 (N_37076,N_34660,N_34428);
xor U37077 (N_37077,N_35727,N_34846);
nor U37078 (N_37078,N_34155,N_35972);
nand U37079 (N_37079,N_34807,N_35086);
xnor U37080 (N_37080,N_35539,N_34883);
and U37081 (N_37081,N_34968,N_34851);
and U37082 (N_37082,N_35001,N_35179);
or U37083 (N_37083,N_35542,N_34997);
nand U37084 (N_37084,N_34956,N_35445);
or U37085 (N_37085,N_35896,N_35296);
nand U37086 (N_37086,N_34522,N_34311);
nor U37087 (N_37087,N_34052,N_34835);
xor U37088 (N_37088,N_34113,N_35314);
xor U37089 (N_37089,N_34612,N_34576);
nand U37090 (N_37090,N_35109,N_35140);
nor U37091 (N_37091,N_35607,N_34156);
or U37092 (N_37092,N_34109,N_35459);
nor U37093 (N_37093,N_35210,N_34497);
xnor U37094 (N_37094,N_34642,N_35344);
and U37095 (N_37095,N_34563,N_35208);
xnor U37096 (N_37096,N_35455,N_34627);
xor U37097 (N_37097,N_35109,N_35394);
xnor U37098 (N_37098,N_35766,N_34019);
xnor U37099 (N_37099,N_35234,N_35841);
or U37100 (N_37100,N_34883,N_34989);
nor U37101 (N_37101,N_35567,N_35029);
and U37102 (N_37102,N_35886,N_34819);
nand U37103 (N_37103,N_34366,N_34220);
xor U37104 (N_37104,N_35277,N_34815);
or U37105 (N_37105,N_35968,N_35538);
nor U37106 (N_37106,N_35078,N_34859);
xor U37107 (N_37107,N_35398,N_34563);
or U37108 (N_37108,N_34913,N_35462);
and U37109 (N_37109,N_35747,N_34283);
nor U37110 (N_37110,N_35734,N_35549);
and U37111 (N_37111,N_35995,N_34825);
nor U37112 (N_37112,N_35138,N_35158);
and U37113 (N_37113,N_35380,N_34639);
xnor U37114 (N_37114,N_35419,N_34722);
nand U37115 (N_37115,N_35300,N_35033);
xnor U37116 (N_37116,N_34447,N_34367);
xnor U37117 (N_37117,N_35410,N_35311);
xnor U37118 (N_37118,N_34579,N_34557);
nand U37119 (N_37119,N_35826,N_35918);
or U37120 (N_37120,N_35432,N_34070);
nor U37121 (N_37121,N_34870,N_35921);
nor U37122 (N_37122,N_35360,N_35647);
or U37123 (N_37123,N_35113,N_35646);
nor U37124 (N_37124,N_34063,N_35318);
nor U37125 (N_37125,N_34671,N_34935);
xnor U37126 (N_37126,N_35488,N_34769);
xor U37127 (N_37127,N_35855,N_35818);
nand U37128 (N_37128,N_35507,N_35488);
nor U37129 (N_37129,N_35592,N_34698);
xnor U37130 (N_37130,N_35365,N_35504);
nor U37131 (N_37131,N_35584,N_34239);
nor U37132 (N_37132,N_35041,N_35021);
nand U37133 (N_37133,N_35091,N_35411);
nor U37134 (N_37134,N_35113,N_34449);
or U37135 (N_37135,N_34984,N_34781);
or U37136 (N_37136,N_34870,N_35507);
nor U37137 (N_37137,N_35183,N_35483);
or U37138 (N_37138,N_34515,N_34913);
and U37139 (N_37139,N_35524,N_35317);
or U37140 (N_37140,N_34069,N_34298);
xor U37141 (N_37141,N_34488,N_35501);
xnor U37142 (N_37142,N_35799,N_35623);
xor U37143 (N_37143,N_35570,N_34238);
and U37144 (N_37144,N_34427,N_35665);
nand U37145 (N_37145,N_34439,N_35006);
xnor U37146 (N_37146,N_35749,N_35018);
xnor U37147 (N_37147,N_35754,N_35455);
and U37148 (N_37148,N_34775,N_34045);
and U37149 (N_37149,N_34507,N_34771);
nor U37150 (N_37150,N_35416,N_35893);
xor U37151 (N_37151,N_34934,N_35510);
or U37152 (N_37152,N_35757,N_34125);
and U37153 (N_37153,N_35956,N_35646);
nand U37154 (N_37154,N_34054,N_35604);
or U37155 (N_37155,N_35105,N_35016);
and U37156 (N_37156,N_35796,N_35517);
nand U37157 (N_37157,N_35480,N_35611);
and U37158 (N_37158,N_34607,N_35970);
nand U37159 (N_37159,N_34761,N_34910);
nand U37160 (N_37160,N_35157,N_34969);
and U37161 (N_37161,N_34472,N_34667);
and U37162 (N_37162,N_35216,N_35500);
or U37163 (N_37163,N_34115,N_34556);
nand U37164 (N_37164,N_35663,N_35441);
nand U37165 (N_37165,N_34214,N_34268);
nand U37166 (N_37166,N_34558,N_34962);
and U37167 (N_37167,N_34373,N_35425);
xor U37168 (N_37168,N_35544,N_35717);
or U37169 (N_37169,N_34947,N_34941);
nor U37170 (N_37170,N_34081,N_35753);
or U37171 (N_37171,N_34555,N_34059);
and U37172 (N_37172,N_35380,N_34571);
nor U37173 (N_37173,N_34290,N_34090);
and U37174 (N_37174,N_35327,N_35911);
and U37175 (N_37175,N_35024,N_34159);
nand U37176 (N_37176,N_34581,N_35649);
nand U37177 (N_37177,N_35876,N_34622);
xor U37178 (N_37178,N_34857,N_35406);
nand U37179 (N_37179,N_34970,N_35819);
or U37180 (N_37180,N_34376,N_35086);
xor U37181 (N_37181,N_35859,N_34408);
or U37182 (N_37182,N_35703,N_35736);
and U37183 (N_37183,N_34875,N_34309);
and U37184 (N_37184,N_35137,N_35310);
or U37185 (N_37185,N_34475,N_35729);
xnor U37186 (N_37186,N_34904,N_34713);
or U37187 (N_37187,N_35547,N_35229);
nand U37188 (N_37188,N_35616,N_35946);
or U37189 (N_37189,N_34683,N_35971);
and U37190 (N_37190,N_34089,N_35389);
and U37191 (N_37191,N_34983,N_35758);
or U37192 (N_37192,N_34112,N_34027);
or U37193 (N_37193,N_34644,N_35048);
or U37194 (N_37194,N_35658,N_34704);
nand U37195 (N_37195,N_34048,N_35454);
and U37196 (N_37196,N_34226,N_34797);
nor U37197 (N_37197,N_35914,N_35471);
and U37198 (N_37198,N_34614,N_34714);
and U37199 (N_37199,N_34522,N_35590);
or U37200 (N_37200,N_35813,N_34888);
and U37201 (N_37201,N_35772,N_34130);
or U37202 (N_37202,N_35232,N_34245);
xor U37203 (N_37203,N_34161,N_35718);
and U37204 (N_37204,N_35355,N_35074);
and U37205 (N_37205,N_34325,N_35238);
nor U37206 (N_37206,N_34252,N_35289);
and U37207 (N_37207,N_35170,N_35350);
nand U37208 (N_37208,N_34715,N_35194);
nor U37209 (N_37209,N_34332,N_35168);
and U37210 (N_37210,N_35720,N_34584);
nor U37211 (N_37211,N_35157,N_35741);
and U37212 (N_37212,N_34467,N_35941);
nand U37213 (N_37213,N_35029,N_34274);
or U37214 (N_37214,N_35376,N_35846);
nor U37215 (N_37215,N_35495,N_34784);
or U37216 (N_37216,N_35721,N_34026);
xor U37217 (N_37217,N_35331,N_34117);
nor U37218 (N_37218,N_34255,N_35622);
and U37219 (N_37219,N_35483,N_35446);
xnor U37220 (N_37220,N_35848,N_35567);
xnor U37221 (N_37221,N_34653,N_34119);
and U37222 (N_37222,N_35331,N_35233);
or U37223 (N_37223,N_34008,N_35174);
nor U37224 (N_37224,N_34500,N_35309);
and U37225 (N_37225,N_34518,N_34945);
and U37226 (N_37226,N_34010,N_34331);
and U37227 (N_37227,N_34522,N_34202);
xor U37228 (N_37228,N_35797,N_34576);
or U37229 (N_37229,N_34197,N_35155);
xor U37230 (N_37230,N_35495,N_35919);
nor U37231 (N_37231,N_35994,N_34521);
nand U37232 (N_37232,N_35368,N_35441);
and U37233 (N_37233,N_35998,N_34006);
nand U37234 (N_37234,N_34234,N_35262);
xor U37235 (N_37235,N_34130,N_34148);
xor U37236 (N_37236,N_35122,N_35667);
or U37237 (N_37237,N_34522,N_34682);
and U37238 (N_37238,N_35781,N_35695);
xor U37239 (N_37239,N_34733,N_34546);
nand U37240 (N_37240,N_35100,N_34500);
and U37241 (N_37241,N_35944,N_34373);
or U37242 (N_37242,N_35148,N_35840);
nand U37243 (N_37243,N_34426,N_35404);
nor U37244 (N_37244,N_35198,N_34482);
and U37245 (N_37245,N_35851,N_35556);
xnor U37246 (N_37246,N_35646,N_35814);
xor U37247 (N_37247,N_35937,N_34297);
nand U37248 (N_37248,N_34871,N_35115);
or U37249 (N_37249,N_35652,N_34613);
or U37250 (N_37250,N_35874,N_35837);
nor U37251 (N_37251,N_35101,N_34063);
nor U37252 (N_37252,N_35024,N_34966);
and U37253 (N_37253,N_34256,N_34379);
or U37254 (N_37254,N_34758,N_34971);
nor U37255 (N_37255,N_35432,N_34677);
and U37256 (N_37256,N_34530,N_34103);
xnor U37257 (N_37257,N_35038,N_34922);
nand U37258 (N_37258,N_35844,N_34878);
nand U37259 (N_37259,N_35315,N_35678);
or U37260 (N_37260,N_34184,N_35274);
or U37261 (N_37261,N_34902,N_34182);
or U37262 (N_37262,N_34340,N_34613);
nand U37263 (N_37263,N_35559,N_35253);
nor U37264 (N_37264,N_35706,N_35090);
nand U37265 (N_37265,N_35315,N_35571);
and U37266 (N_37266,N_34573,N_34040);
nor U37267 (N_37267,N_35599,N_35940);
xnor U37268 (N_37268,N_35603,N_34681);
or U37269 (N_37269,N_34611,N_34762);
nor U37270 (N_37270,N_35115,N_35207);
nand U37271 (N_37271,N_34466,N_34704);
nand U37272 (N_37272,N_35408,N_35236);
nand U37273 (N_37273,N_35182,N_34102);
and U37274 (N_37274,N_35166,N_35591);
nor U37275 (N_37275,N_34496,N_34867);
nand U37276 (N_37276,N_35490,N_35550);
nor U37277 (N_37277,N_34008,N_34666);
or U37278 (N_37278,N_34936,N_34091);
nand U37279 (N_37279,N_35309,N_35580);
nand U37280 (N_37280,N_35760,N_34965);
nand U37281 (N_37281,N_35929,N_35607);
or U37282 (N_37282,N_34113,N_34246);
nor U37283 (N_37283,N_34989,N_34027);
nand U37284 (N_37284,N_35356,N_34308);
nand U37285 (N_37285,N_35175,N_35656);
or U37286 (N_37286,N_34904,N_34170);
xnor U37287 (N_37287,N_34360,N_35254);
or U37288 (N_37288,N_35440,N_35426);
and U37289 (N_37289,N_35588,N_35825);
xor U37290 (N_37290,N_34939,N_35071);
nor U37291 (N_37291,N_34686,N_35577);
nor U37292 (N_37292,N_35702,N_35118);
or U37293 (N_37293,N_34284,N_35449);
nor U37294 (N_37294,N_34731,N_35383);
xor U37295 (N_37295,N_34646,N_34521);
xor U37296 (N_37296,N_35013,N_34738);
nor U37297 (N_37297,N_35291,N_35199);
nor U37298 (N_37298,N_34472,N_35745);
and U37299 (N_37299,N_35769,N_34307);
and U37300 (N_37300,N_35591,N_34052);
and U37301 (N_37301,N_35028,N_35754);
xnor U37302 (N_37302,N_35806,N_34316);
xor U37303 (N_37303,N_35277,N_35044);
and U37304 (N_37304,N_35251,N_34431);
nor U37305 (N_37305,N_34474,N_35418);
xor U37306 (N_37306,N_35077,N_34419);
nor U37307 (N_37307,N_34489,N_35434);
or U37308 (N_37308,N_35468,N_35632);
nand U37309 (N_37309,N_34419,N_34727);
xnor U37310 (N_37310,N_35391,N_34332);
nor U37311 (N_37311,N_35102,N_35397);
and U37312 (N_37312,N_34137,N_34397);
or U37313 (N_37313,N_35285,N_34203);
xor U37314 (N_37314,N_35559,N_34982);
nor U37315 (N_37315,N_34358,N_34373);
nor U37316 (N_37316,N_34050,N_34039);
and U37317 (N_37317,N_34510,N_34436);
nor U37318 (N_37318,N_35680,N_34045);
or U37319 (N_37319,N_34719,N_34087);
and U37320 (N_37320,N_35198,N_35680);
xor U37321 (N_37321,N_35381,N_35463);
nor U37322 (N_37322,N_35154,N_34415);
xor U37323 (N_37323,N_35945,N_35838);
or U37324 (N_37324,N_34779,N_35592);
nor U37325 (N_37325,N_34402,N_34448);
and U37326 (N_37326,N_34010,N_35050);
and U37327 (N_37327,N_34556,N_35675);
nor U37328 (N_37328,N_34132,N_35333);
or U37329 (N_37329,N_34620,N_34656);
nor U37330 (N_37330,N_35103,N_35928);
nand U37331 (N_37331,N_35889,N_34191);
nor U37332 (N_37332,N_34052,N_34976);
xnor U37333 (N_37333,N_35910,N_34707);
nor U37334 (N_37334,N_35159,N_35459);
nor U37335 (N_37335,N_34883,N_35113);
and U37336 (N_37336,N_35582,N_35952);
xor U37337 (N_37337,N_35697,N_34427);
and U37338 (N_37338,N_35206,N_35269);
and U37339 (N_37339,N_34358,N_35570);
nor U37340 (N_37340,N_35096,N_35285);
nor U37341 (N_37341,N_35368,N_35394);
nand U37342 (N_37342,N_34110,N_34327);
nor U37343 (N_37343,N_35295,N_35003);
nand U37344 (N_37344,N_34506,N_34578);
nand U37345 (N_37345,N_34521,N_35007);
nand U37346 (N_37346,N_34608,N_34857);
or U37347 (N_37347,N_35752,N_35129);
nand U37348 (N_37348,N_35891,N_35350);
nand U37349 (N_37349,N_35789,N_34865);
and U37350 (N_37350,N_34779,N_35651);
nor U37351 (N_37351,N_35917,N_34642);
and U37352 (N_37352,N_35663,N_35528);
and U37353 (N_37353,N_34044,N_35056);
and U37354 (N_37354,N_35638,N_34991);
xor U37355 (N_37355,N_35882,N_35092);
xor U37356 (N_37356,N_34630,N_35754);
and U37357 (N_37357,N_34758,N_34415);
and U37358 (N_37358,N_35641,N_35352);
nor U37359 (N_37359,N_34556,N_35595);
nand U37360 (N_37360,N_35403,N_34773);
nor U37361 (N_37361,N_34274,N_34386);
and U37362 (N_37362,N_35500,N_35498);
nor U37363 (N_37363,N_35570,N_35932);
nor U37364 (N_37364,N_34143,N_35372);
nand U37365 (N_37365,N_34399,N_35614);
nor U37366 (N_37366,N_35961,N_34096);
nand U37367 (N_37367,N_35741,N_35233);
nor U37368 (N_37368,N_35079,N_35298);
or U37369 (N_37369,N_35622,N_35234);
or U37370 (N_37370,N_35767,N_35569);
and U37371 (N_37371,N_35701,N_34150);
nand U37372 (N_37372,N_35389,N_34451);
and U37373 (N_37373,N_34382,N_35277);
or U37374 (N_37374,N_34065,N_34548);
xor U37375 (N_37375,N_34771,N_35194);
xnor U37376 (N_37376,N_34468,N_35952);
and U37377 (N_37377,N_34310,N_34743);
xnor U37378 (N_37378,N_35979,N_34411);
nor U37379 (N_37379,N_35056,N_34120);
nand U37380 (N_37380,N_34788,N_35672);
and U37381 (N_37381,N_34962,N_35981);
nand U37382 (N_37382,N_34574,N_34595);
nand U37383 (N_37383,N_35320,N_34766);
nor U37384 (N_37384,N_34869,N_34437);
xor U37385 (N_37385,N_34778,N_35409);
and U37386 (N_37386,N_35959,N_35999);
nand U37387 (N_37387,N_34468,N_35533);
nand U37388 (N_37388,N_35547,N_35279);
nand U37389 (N_37389,N_34940,N_34075);
and U37390 (N_37390,N_34178,N_34213);
nor U37391 (N_37391,N_35476,N_34643);
nand U37392 (N_37392,N_34436,N_34894);
xor U37393 (N_37393,N_35724,N_34891);
and U37394 (N_37394,N_35125,N_35902);
nand U37395 (N_37395,N_34236,N_35603);
xor U37396 (N_37396,N_34812,N_35697);
nor U37397 (N_37397,N_35128,N_34944);
and U37398 (N_37398,N_34071,N_35268);
or U37399 (N_37399,N_35448,N_34558);
or U37400 (N_37400,N_34910,N_35660);
or U37401 (N_37401,N_35187,N_35101);
or U37402 (N_37402,N_34622,N_35108);
and U37403 (N_37403,N_35257,N_35420);
nor U37404 (N_37404,N_34687,N_35544);
and U37405 (N_37405,N_35522,N_35648);
and U37406 (N_37406,N_34228,N_34772);
xnor U37407 (N_37407,N_35754,N_35760);
and U37408 (N_37408,N_35923,N_34813);
or U37409 (N_37409,N_35811,N_35016);
and U37410 (N_37410,N_34494,N_35171);
xnor U37411 (N_37411,N_35723,N_34406);
xor U37412 (N_37412,N_34133,N_34552);
nor U37413 (N_37413,N_34554,N_34593);
xnor U37414 (N_37414,N_34150,N_34370);
nor U37415 (N_37415,N_35774,N_34193);
nand U37416 (N_37416,N_35511,N_35300);
and U37417 (N_37417,N_35376,N_35436);
nand U37418 (N_37418,N_35173,N_35319);
nand U37419 (N_37419,N_35943,N_34976);
and U37420 (N_37420,N_34093,N_34976);
nand U37421 (N_37421,N_35089,N_35709);
xor U37422 (N_37422,N_34408,N_34450);
and U37423 (N_37423,N_34769,N_35031);
nand U37424 (N_37424,N_35906,N_35981);
or U37425 (N_37425,N_35939,N_35751);
nor U37426 (N_37426,N_35061,N_34641);
or U37427 (N_37427,N_35082,N_34169);
or U37428 (N_37428,N_35541,N_35809);
xnor U37429 (N_37429,N_34453,N_34315);
nand U37430 (N_37430,N_34173,N_35677);
xnor U37431 (N_37431,N_34530,N_34556);
nand U37432 (N_37432,N_35932,N_35298);
and U37433 (N_37433,N_35769,N_34908);
nand U37434 (N_37434,N_34228,N_34382);
nor U37435 (N_37435,N_35997,N_34445);
and U37436 (N_37436,N_34355,N_34820);
nand U37437 (N_37437,N_34601,N_35328);
xor U37438 (N_37438,N_35550,N_34160);
xnor U37439 (N_37439,N_35076,N_34270);
or U37440 (N_37440,N_34264,N_34424);
xor U37441 (N_37441,N_34224,N_34798);
xnor U37442 (N_37442,N_35988,N_35759);
nand U37443 (N_37443,N_34934,N_35480);
xnor U37444 (N_37444,N_35933,N_35661);
xnor U37445 (N_37445,N_34707,N_34088);
or U37446 (N_37446,N_34073,N_35492);
or U37447 (N_37447,N_35373,N_35274);
nor U37448 (N_37448,N_34677,N_34330);
nand U37449 (N_37449,N_34272,N_35837);
nand U37450 (N_37450,N_35625,N_34916);
and U37451 (N_37451,N_35835,N_34729);
nor U37452 (N_37452,N_35213,N_35823);
xnor U37453 (N_37453,N_34331,N_35674);
and U37454 (N_37454,N_35096,N_35153);
nand U37455 (N_37455,N_34508,N_34672);
or U37456 (N_37456,N_34866,N_34597);
xor U37457 (N_37457,N_34401,N_34275);
nand U37458 (N_37458,N_34779,N_35677);
nand U37459 (N_37459,N_35829,N_34807);
and U37460 (N_37460,N_35399,N_34746);
xor U37461 (N_37461,N_35250,N_34599);
and U37462 (N_37462,N_35578,N_35101);
xnor U37463 (N_37463,N_35597,N_35623);
nand U37464 (N_37464,N_34230,N_35718);
nand U37465 (N_37465,N_34166,N_34564);
or U37466 (N_37466,N_34190,N_34532);
and U37467 (N_37467,N_34901,N_35088);
and U37468 (N_37468,N_34371,N_35736);
nor U37469 (N_37469,N_35358,N_35722);
and U37470 (N_37470,N_34580,N_34262);
nand U37471 (N_37471,N_35406,N_34585);
xnor U37472 (N_37472,N_34447,N_34613);
xor U37473 (N_37473,N_35526,N_35396);
xor U37474 (N_37474,N_35698,N_34413);
xnor U37475 (N_37475,N_35204,N_35089);
xnor U37476 (N_37476,N_35868,N_34826);
or U37477 (N_37477,N_34124,N_34058);
xnor U37478 (N_37478,N_34045,N_35554);
nor U37479 (N_37479,N_34850,N_34901);
nand U37480 (N_37480,N_34359,N_34175);
and U37481 (N_37481,N_34479,N_34702);
and U37482 (N_37482,N_34291,N_35938);
nor U37483 (N_37483,N_34324,N_34336);
nor U37484 (N_37484,N_34562,N_35254);
nor U37485 (N_37485,N_35062,N_35648);
or U37486 (N_37486,N_34920,N_34582);
or U37487 (N_37487,N_35545,N_35811);
nor U37488 (N_37488,N_34291,N_35715);
nor U37489 (N_37489,N_34207,N_35997);
nor U37490 (N_37490,N_35614,N_35554);
nand U37491 (N_37491,N_34507,N_34969);
nand U37492 (N_37492,N_35605,N_34933);
and U37493 (N_37493,N_35271,N_34106);
xor U37494 (N_37494,N_35489,N_34541);
nor U37495 (N_37495,N_34812,N_35483);
xnor U37496 (N_37496,N_34081,N_35693);
and U37497 (N_37497,N_35526,N_34841);
nor U37498 (N_37498,N_34180,N_34722);
nor U37499 (N_37499,N_35847,N_34372);
xnor U37500 (N_37500,N_34414,N_35000);
nor U37501 (N_37501,N_35817,N_35670);
or U37502 (N_37502,N_34977,N_35242);
or U37503 (N_37503,N_35362,N_35829);
xnor U37504 (N_37504,N_35848,N_34788);
and U37505 (N_37505,N_35284,N_35185);
and U37506 (N_37506,N_34925,N_34873);
nand U37507 (N_37507,N_35396,N_35762);
nor U37508 (N_37508,N_35439,N_35974);
and U37509 (N_37509,N_35566,N_34703);
or U37510 (N_37510,N_34150,N_35714);
nand U37511 (N_37511,N_35297,N_34955);
nor U37512 (N_37512,N_35189,N_35033);
and U37513 (N_37513,N_35906,N_35320);
nor U37514 (N_37514,N_35689,N_34553);
xor U37515 (N_37515,N_34204,N_34531);
nor U37516 (N_37516,N_35773,N_34111);
and U37517 (N_37517,N_34355,N_34255);
or U37518 (N_37518,N_35677,N_34532);
nor U37519 (N_37519,N_34945,N_35895);
nor U37520 (N_37520,N_35860,N_34008);
xor U37521 (N_37521,N_34176,N_34057);
and U37522 (N_37522,N_35229,N_34613);
or U37523 (N_37523,N_35320,N_34165);
nand U37524 (N_37524,N_35801,N_35378);
and U37525 (N_37525,N_34820,N_34408);
and U37526 (N_37526,N_34360,N_34165);
nand U37527 (N_37527,N_35169,N_35853);
xor U37528 (N_37528,N_35798,N_34685);
and U37529 (N_37529,N_35716,N_35732);
nor U37530 (N_37530,N_34253,N_34790);
nand U37531 (N_37531,N_34476,N_35020);
or U37532 (N_37532,N_35498,N_34807);
and U37533 (N_37533,N_35475,N_35814);
nand U37534 (N_37534,N_35122,N_34271);
nand U37535 (N_37535,N_35754,N_35438);
xor U37536 (N_37536,N_34017,N_35942);
or U37537 (N_37537,N_35643,N_34990);
xnor U37538 (N_37538,N_34584,N_35492);
or U37539 (N_37539,N_34609,N_35204);
and U37540 (N_37540,N_34693,N_35782);
nor U37541 (N_37541,N_34422,N_35360);
nand U37542 (N_37542,N_34955,N_34253);
or U37543 (N_37543,N_34601,N_34015);
nor U37544 (N_37544,N_34471,N_35121);
nor U37545 (N_37545,N_34006,N_34642);
and U37546 (N_37546,N_34546,N_34952);
nor U37547 (N_37547,N_34941,N_34739);
nor U37548 (N_37548,N_34725,N_34145);
nand U37549 (N_37549,N_35097,N_34245);
and U37550 (N_37550,N_35885,N_34598);
or U37551 (N_37551,N_34026,N_34372);
nand U37552 (N_37552,N_34649,N_34459);
xor U37553 (N_37553,N_34124,N_34368);
or U37554 (N_37554,N_35818,N_35049);
or U37555 (N_37555,N_34292,N_34386);
xnor U37556 (N_37556,N_34935,N_34389);
and U37557 (N_37557,N_35996,N_34601);
or U37558 (N_37558,N_35250,N_34018);
nor U37559 (N_37559,N_35099,N_34150);
nor U37560 (N_37560,N_35108,N_34651);
or U37561 (N_37561,N_34336,N_34656);
or U37562 (N_37562,N_34875,N_35714);
and U37563 (N_37563,N_34980,N_35202);
or U37564 (N_37564,N_35444,N_35697);
or U37565 (N_37565,N_34891,N_35891);
xnor U37566 (N_37566,N_35948,N_34132);
nor U37567 (N_37567,N_35488,N_35257);
or U37568 (N_37568,N_34789,N_35946);
or U37569 (N_37569,N_35083,N_35194);
or U37570 (N_37570,N_35293,N_34688);
and U37571 (N_37571,N_34124,N_35264);
nor U37572 (N_37572,N_35143,N_34091);
or U37573 (N_37573,N_34554,N_34590);
xnor U37574 (N_37574,N_34654,N_34569);
nand U37575 (N_37575,N_34725,N_35580);
or U37576 (N_37576,N_34994,N_35872);
and U37577 (N_37577,N_35209,N_35778);
nor U37578 (N_37578,N_34435,N_34935);
and U37579 (N_37579,N_35900,N_34268);
nand U37580 (N_37580,N_35056,N_35676);
or U37581 (N_37581,N_34142,N_35561);
xnor U37582 (N_37582,N_35744,N_34286);
xor U37583 (N_37583,N_34055,N_35519);
or U37584 (N_37584,N_34779,N_35567);
nand U37585 (N_37585,N_35569,N_34265);
nand U37586 (N_37586,N_34984,N_35574);
or U37587 (N_37587,N_35590,N_35103);
and U37588 (N_37588,N_34360,N_35167);
nor U37589 (N_37589,N_35823,N_34463);
and U37590 (N_37590,N_35648,N_35759);
nor U37591 (N_37591,N_35773,N_34609);
nand U37592 (N_37592,N_35605,N_35851);
and U37593 (N_37593,N_35334,N_34605);
nor U37594 (N_37594,N_34120,N_35023);
and U37595 (N_37595,N_35846,N_35975);
nand U37596 (N_37596,N_35635,N_34088);
nor U37597 (N_37597,N_35280,N_35080);
and U37598 (N_37598,N_35377,N_34921);
nand U37599 (N_37599,N_34196,N_34153);
xor U37600 (N_37600,N_34704,N_35113);
nor U37601 (N_37601,N_35356,N_34924);
or U37602 (N_37602,N_35393,N_35084);
and U37603 (N_37603,N_35792,N_34065);
and U37604 (N_37604,N_35681,N_35174);
nor U37605 (N_37605,N_34279,N_34265);
nand U37606 (N_37606,N_35817,N_34600);
nor U37607 (N_37607,N_34746,N_34135);
and U37608 (N_37608,N_35965,N_34420);
or U37609 (N_37609,N_35616,N_35092);
and U37610 (N_37610,N_34458,N_34686);
nand U37611 (N_37611,N_34173,N_34336);
nor U37612 (N_37612,N_35953,N_35288);
nand U37613 (N_37613,N_34192,N_34118);
nand U37614 (N_37614,N_34974,N_35878);
or U37615 (N_37615,N_34290,N_35387);
and U37616 (N_37616,N_35763,N_35686);
or U37617 (N_37617,N_34554,N_34905);
and U37618 (N_37618,N_34321,N_34395);
nor U37619 (N_37619,N_34446,N_35509);
or U37620 (N_37620,N_35753,N_35389);
nor U37621 (N_37621,N_34652,N_35908);
and U37622 (N_37622,N_34084,N_35056);
and U37623 (N_37623,N_35556,N_35874);
nor U37624 (N_37624,N_34189,N_34320);
xnor U37625 (N_37625,N_34747,N_35687);
or U37626 (N_37626,N_35737,N_34598);
nand U37627 (N_37627,N_35167,N_35182);
and U37628 (N_37628,N_35619,N_35341);
or U37629 (N_37629,N_34038,N_34752);
xor U37630 (N_37630,N_35031,N_34417);
nor U37631 (N_37631,N_34861,N_35877);
or U37632 (N_37632,N_35585,N_35675);
or U37633 (N_37633,N_35832,N_34558);
xnor U37634 (N_37634,N_35126,N_34367);
and U37635 (N_37635,N_34663,N_34521);
nor U37636 (N_37636,N_35484,N_34581);
nor U37637 (N_37637,N_34666,N_35906);
nand U37638 (N_37638,N_34162,N_35402);
xnor U37639 (N_37639,N_35737,N_34500);
xor U37640 (N_37640,N_34376,N_34217);
or U37641 (N_37641,N_35837,N_35102);
nor U37642 (N_37642,N_35754,N_34464);
and U37643 (N_37643,N_35927,N_34137);
nor U37644 (N_37644,N_34530,N_34994);
xor U37645 (N_37645,N_35994,N_34874);
nor U37646 (N_37646,N_34330,N_35326);
or U37647 (N_37647,N_35268,N_35207);
and U37648 (N_37648,N_34126,N_35724);
nand U37649 (N_37649,N_34999,N_34574);
nor U37650 (N_37650,N_35421,N_34885);
nand U37651 (N_37651,N_34854,N_35779);
nand U37652 (N_37652,N_35759,N_35003);
or U37653 (N_37653,N_34159,N_35637);
nor U37654 (N_37654,N_35346,N_34577);
xnor U37655 (N_37655,N_35017,N_35679);
nand U37656 (N_37656,N_34507,N_35761);
xor U37657 (N_37657,N_35683,N_35720);
and U37658 (N_37658,N_35247,N_35913);
nor U37659 (N_37659,N_34661,N_35763);
xor U37660 (N_37660,N_35161,N_34908);
and U37661 (N_37661,N_34479,N_35630);
nor U37662 (N_37662,N_35464,N_34987);
nand U37663 (N_37663,N_34532,N_35647);
and U37664 (N_37664,N_34238,N_35783);
and U37665 (N_37665,N_34945,N_34887);
nand U37666 (N_37666,N_34037,N_35357);
and U37667 (N_37667,N_34246,N_34534);
or U37668 (N_37668,N_34061,N_34266);
xnor U37669 (N_37669,N_35108,N_35621);
and U37670 (N_37670,N_35537,N_35593);
nand U37671 (N_37671,N_34010,N_34695);
nand U37672 (N_37672,N_34876,N_35514);
or U37673 (N_37673,N_35138,N_35801);
xnor U37674 (N_37674,N_35678,N_34815);
nor U37675 (N_37675,N_35477,N_34195);
or U37676 (N_37676,N_35212,N_35573);
or U37677 (N_37677,N_35699,N_35895);
nand U37678 (N_37678,N_34050,N_35456);
nand U37679 (N_37679,N_34092,N_34417);
and U37680 (N_37680,N_35106,N_35066);
nor U37681 (N_37681,N_35194,N_35965);
nor U37682 (N_37682,N_34946,N_35605);
and U37683 (N_37683,N_35110,N_35232);
nor U37684 (N_37684,N_35388,N_34137);
xor U37685 (N_37685,N_34575,N_34901);
nand U37686 (N_37686,N_35921,N_34722);
and U37687 (N_37687,N_34913,N_34035);
or U37688 (N_37688,N_34764,N_35016);
xor U37689 (N_37689,N_34027,N_35524);
or U37690 (N_37690,N_35634,N_35016);
or U37691 (N_37691,N_35470,N_34832);
or U37692 (N_37692,N_35237,N_35394);
or U37693 (N_37693,N_34349,N_34934);
or U37694 (N_37694,N_35086,N_34191);
nor U37695 (N_37695,N_34646,N_34183);
and U37696 (N_37696,N_34823,N_35154);
and U37697 (N_37697,N_35830,N_35473);
nor U37698 (N_37698,N_34289,N_34797);
and U37699 (N_37699,N_35611,N_35417);
nand U37700 (N_37700,N_34641,N_34446);
and U37701 (N_37701,N_34654,N_35935);
nand U37702 (N_37702,N_34161,N_35908);
nor U37703 (N_37703,N_34062,N_34369);
nor U37704 (N_37704,N_34416,N_34224);
nand U37705 (N_37705,N_34808,N_34825);
and U37706 (N_37706,N_35549,N_34398);
or U37707 (N_37707,N_35874,N_34332);
nand U37708 (N_37708,N_35255,N_34919);
nand U37709 (N_37709,N_34670,N_35737);
nor U37710 (N_37710,N_35569,N_35085);
xor U37711 (N_37711,N_34154,N_35551);
xor U37712 (N_37712,N_35924,N_35154);
or U37713 (N_37713,N_35714,N_35914);
nand U37714 (N_37714,N_34709,N_34213);
nand U37715 (N_37715,N_34496,N_35074);
or U37716 (N_37716,N_35442,N_35772);
nor U37717 (N_37717,N_34978,N_35994);
or U37718 (N_37718,N_34805,N_35107);
nor U37719 (N_37719,N_34776,N_35696);
xor U37720 (N_37720,N_35612,N_34392);
or U37721 (N_37721,N_34964,N_35701);
xnor U37722 (N_37722,N_34529,N_35555);
or U37723 (N_37723,N_35953,N_34745);
and U37724 (N_37724,N_35280,N_34955);
nor U37725 (N_37725,N_34511,N_34784);
nor U37726 (N_37726,N_34145,N_34179);
xnor U37727 (N_37727,N_34759,N_34776);
or U37728 (N_37728,N_34018,N_35088);
nand U37729 (N_37729,N_34926,N_35739);
or U37730 (N_37730,N_34614,N_34511);
nand U37731 (N_37731,N_35990,N_34800);
or U37732 (N_37732,N_35482,N_35451);
or U37733 (N_37733,N_35281,N_35479);
nor U37734 (N_37734,N_35914,N_35492);
and U37735 (N_37735,N_35868,N_35001);
nand U37736 (N_37736,N_35083,N_35710);
nand U37737 (N_37737,N_35089,N_35131);
or U37738 (N_37738,N_35412,N_34876);
nand U37739 (N_37739,N_34515,N_35824);
or U37740 (N_37740,N_35815,N_34832);
nor U37741 (N_37741,N_35071,N_35235);
and U37742 (N_37742,N_35451,N_35352);
or U37743 (N_37743,N_34480,N_35831);
nand U37744 (N_37744,N_35638,N_35681);
nand U37745 (N_37745,N_34299,N_35979);
or U37746 (N_37746,N_34393,N_35249);
nand U37747 (N_37747,N_34953,N_34863);
and U37748 (N_37748,N_34850,N_34191);
nand U37749 (N_37749,N_35517,N_34421);
or U37750 (N_37750,N_34079,N_34476);
or U37751 (N_37751,N_35633,N_34044);
xnor U37752 (N_37752,N_34895,N_35166);
or U37753 (N_37753,N_34500,N_34734);
and U37754 (N_37754,N_35986,N_35463);
and U37755 (N_37755,N_34845,N_35015);
or U37756 (N_37756,N_34753,N_35151);
nand U37757 (N_37757,N_35479,N_34922);
xnor U37758 (N_37758,N_35183,N_34705);
nor U37759 (N_37759,N_35628,N_34954);
nor U37760 (N_37760,N_35921,N_34078);
or U37761 (N_37761,N_35141,N_35438);
and U37762 (N_37762,N_34142,N_34097);
nor U37763 (N_37763,N_34078,N_35525);
and U37764 (N_37764,N_34478,N_35631);
and U37765 (N_37765,N_34275,N_35920);
nand U37766 (N_37766,N_34986,N_35801);
or U37767 (N_37767,N_34599,N_34183);
nand U37768 (N_37768,N_35149,N_35801);
nand U37769 (N_37769,N_35373,N_34218);
or U37770 (N_37770,N_34169,N_34994);
and U37771 (N_37771,N_34083,N_34816);
nand U37772 (N_37772,N_34221,N_34867);
or U37773 (N_37773,N_35251,N_34620);
or U37774 (N_37774,N_34409,N_34526);
xnor U37775 (N_37775,N_35701,N_35605);
nand U37776 (N_37776,N_34396,N_35126);
nor U37777 (N_37777,N_35258,N_35273);
xnor U37778 (N_37778,N_34268,N_35656);
nand U37779 (N_37779,N_35461,N_35336);
nand U37780 (N_37780,N_34508,N_35008);
and U37781 (N_37781,N_34766,N_34187);
nor U37782 (N_37782,N_35196,N_34311);
nor U37783 (N_37783,N_35506,N_34777);
nor U37784 (N_37784,N_35647,N_34213);
and U37785 (N_37785,N_35004,N_34568);
xor U37786 (N_37786,N_34920,N_35935);
or U37787 (N_37787,N_34294,N_35350);
and U37788 (N_37788,N_34605,N_35956);
xor U37789 (N_37789,N_34644,N_34699);
xnor U37790 (N_37790,N_34517,N_35664);
nand U37791 (N_37791,N_35922,N_34459);
nor U37792 (N_37792,N_34103,N_35044);
or U37793 (N_37793,N_34641,N_34666);
and U37794 (N_37794,N_34149,N_34174);
nand U37795 (N_37795,N_34692,N_35501);
and U37796 (N_37796,N_35872,N_34150);
and U37797 (N_37797,N_34571,N_35591);
or U37798 (N_37798,N_35579,N_34298);
xnor U37799 (N_37799,N_34405,N_35421);
and U37800 (N_37800,N_34620,N_35078);
nor U37801 (N_37801,N_35094,N_34635);
nand U37802 (N_37802,N_35092,N_34097);
and U37803 (N_37803,N_35195,N_34326);
or U37804 (N_37804,N_34837,N_34678);
xnor U37805 (N_37805,N_35989,N_35189);
or U37806 (N_37806,N_34606,N_35978);
nand U37807 (N_37807,N_34882,N_34450);
nor U37808 (N_37808,N_35705,N_34832);
or U37809 (N_37809,N_35429,N_34604);
xor U37810 (N_37810,N_35204,N_35499);
and U37811 (N_37811,N_35356,N_34609);
nor U37812 (N_37812,N_35442,N_34398);
and U37813 (N_37813,N_34985,N_34020);
nor U37814 (N_37814,N_35196,N_34711);
nand U37815 (N_37815,N_34852,N_34585);
xor U37816 (N_37816,N_34346,N_34506);
nor U37817 (N_37817,N_34535,N_34028);
or U37818 (N_37818,N_34041,N_35741);
nor U37819 (N_37819,N_34769,N_34065);
xor U37820 (N_37820,N_34550,N_34318);
nor U37821 (N_37821,N_35336,N_35760);
xor U37822 (N_37822,N_35581,N_35213);
xnor U37823 (N_37823,N_35332,N_34924);
xnor U37824 (N_37824,N_35995,N_34421);
nor U37825 (N_37825,N_35883,N_35990);
or U37826 (N_37826,N_34044,N_34598);
xor U37827 (N_37827,N_34149,N_34450);
or U37828 (N_37828,N_34634,N_34346);
or U37829 (N_37829,N_35599,N_35679);
or U37830 (N_37830,N_34655,N_34000);
and U37831 (N_37831,N_35707,N_35123);
nor U37832 (N_37832,N_34964,N_35312);
nor U37833 (N_37833,N_35443,N_35308);
xnor U37834 (N_37834,N_35629,N_35613);
and U37835 (N_37835,N_34360,N_35337);
nand U37836 (N_37836,N_34165,N_35350);
nor U37837 (N_37837,N_34873,N_35466);
and U37838 (N_37838,N_35921,N_35191);
nand U37839 (N_37839,N_35895,N_35231);
nand U37840 (N_37840,N_34833,N_35375);
and U37841 (N_37841,N_34083,N_35022);
nand U37842 (N_37842,N_35115,N_35097);
nor U37843 (N_37843,N_35430,N_34725);
xor U37844 (N_37844,N_35677,N_34703);
and U37845 (N_37845,N_34211,N_34994);
nand U37846 (N_37846,N_35063,N_35188);
nand U37847 (N_37847,N_35559,N_35738);
xor U37848 (N_37848,N_35680,N_34279);
nand U37849 (N_37849,N_34870,N_34142);
xnor U37850 (N_37850,N_34306,N_34533);
nor U37851 (N_37851,N_34632,N_34805);
or U37852 (N_37852,N_35231,N_35768);
nor U37853 (N_37853,N_34780,N_34682);
or U37854 (N_37854,N_35571,N_35325);
and U37855 (N_37855,N_35808,N_34168);
xnor U37856 (N_37856,N_35068,N_35240);
nand U37857 (N_37857,N_35777,N_35316);
nand U37858 (N_37858,N_34768,N_35910);
or U37859 (N_37859,N_35128,N_35792);
xnor U37860 (N_37860,N_35045,N_34695);
nand U37861 (N_37861,N_35218,N_34559);
nor U37862 (N_37862,N_35769,N_35444);
nor U37863 (N_37863,N_35543,N_35164);
nor U37864 (N_37864,N_34228,N_35109);
xnor U37865 (N_37865,N_34607,N_34320);
and U37866 (N_37866,N_35439,N_34222);
and U37867 (N_37867,N_34526,N_35958);
and U37868 (N_37868,N_35075,N_34600);
and U37869 (N_37869,N_35173,N_34036);
nor U37870 (N_37870,N_35575,N_34561);
xnor U37871 (N_37871,N_34017,N_34709);
nor U37872 (N_37872,N_34616,N_35993);
and U37873 (N_37873,N_35461,N_35076);
xnor U37874 (N_37874,N_34682,N_34126);
nand U37875 (N_37875,N_34574,N_35294);
nand U37876 (N_37876,N_34121,N_35345);
or U37877 (N_37877,N_35393,N_35682);
xor U37878 (N_37878,N_35569,N_34429);
and U37879 (N_37879,N_34852,N_35334);
xnor U37880 (N_37880,N_34504,N_35126);
xnor U37881 (N_37881,N_34666,N_34012);
xnor U37882 (N_37882,N_35664,N_35203);
or U37883 (N_37883,N_34354,N_35702);
and U37884 (N_37884,N_35349,N_34200);
and U37885 (N_37885,N_34350,N_34402);
nor U37886 (N_37886,N_34355,N_35775);
and U37887 (N_37887,N_35433,N_35812);
xor U37888 (N_37888,N_35156,N_35263);
or U37889 (N_37889,N_34501,N_34681);
or U37890 (N_37890,N_35508,N_35140);
xnor U37891 (N_37891,N_34987,N_35853);
nand U37892 (N_37892,N_34914,N_35566);
nor U37893 (N_37893,N_35770,N_34841);
xor U37894 (N_37894,N_35891,N_35125);
and U37895 (N_37895,N_34048,N_34748);
and U37896 (N_37896,N_35848,N_35198);
xnor U37897 (N_37897,N_34904,N_35741);
and U37898 (N_37898,N_34947,N_35037);
nor U37899 (N_37899,N_34846,N_35364);
or U37900 (N_37900,N_34695,N_34404);
or U37901 (N_37901,N_35579,N_35943);
and U37902 (N_37902,N_34771,N_35686);
nor U37903 (N_37903,N_35195,N_35337);
nor U37904 (N_37904,N_35587,N_35806);
xor U37905 (N_37905,N_35828,N_34992);
xnor U37906 (N_37906,N_34526,N_35090);
xor U37907 (N_37907,N_35231,N_35518);
nor U37908 (N_37908,N_34688,N_35497);
and U37909 (N_37909,N_34096,N_35775);
xor U37910 (N_37910,N_34186,N_34178);
or U37911 (N_37911,N_35174,N_34350);
and U37912 (N_37912,N_34592,N_34315);
nand U37913 (N_37913,N_34054,N_34626);
xor U37914 (N_37914,N_35070,N_35633);
or U37915 (N_37915,N_35706,N_35769);
nor U37916 (N_37916,N_35989,N_34992);
or U37917 (N_37917,N_35388,N_34221);
nor U37918 (N_37918,N_34764,N_34428);
nor U37919 (N_37919,N_34590,N_34595);
or U37920 (N_37920,N_34663,N_35386);
or U37921 (N_37921,N_34640,N_35920);
nor U37922 (N_37922,N_34741,N_35754);
nand U37923 (N_37923,N_34248,N_34222);
nand U37924 (N_37924,N_35152,N_34706);
xor U37925 (N_37925,N_34962,N_34037);
xor U37926 (N_37926,N_34872,N_34777);
nor U37927 (N_37927,N_35894,N_35154);
xnor U37928 (N_37928,N_34716,N_34384);
xor U37929 (N_37929,N_35537,N_35254);
and U37930 (N_37930,N_35752,N_35587);
and U37931 (N_37931,N_35891,N_35226);
and U37932 (N_37932,N_35317,N_35933);
nor U37933 (N_37933,N_35709,N_35326);
xor U37934 (N_37934,N_34795,N_35694);
and U37935 (N_37935,N_34157,N_34214);
xor U37936 (N_37936,N_35234,N_35837);
and U37937 (N_37937,N_34271,N_34605);
xnor U37938 (N_37938,N_34032,N_34653);
and U37939 (N_37939,N_35667,N_34667);
and U37940 (N_37940,N_35287,N_35579);
and U37941 (N_37941,N_34662,N_34800);
and U37942 (N_37942,N_35818,N_34247);
nand U37943 (N_37943,N_35829,N_35498);
or U37944 (N_37944,N_35398,N_34031);
xnor U37945 (N_37945,N_35872,N_34409);
and U37946 (N_37946,N_35358,N_34468);
and U37947 (N_37947,N_35899,N_34661);
xnor U37948 (N_37948,N_34899,N_35531);
nand U37949 (N_37949,N_34898,N_34409);
nor U37950 (N_37950,N_35171,N_34853);
nor U37951 (N_37951,N_35734,N_35827);
xor U37952 (N_37952,N_35967,N_35668);
xnor U37953 (N_37953,N_35339,N_34749);
nand U37954 (N_37954,N_35499,N_34067);
or U37955 (N_37955,N_34585,N_34611);
xor U37956 (N_37956,N_35697,N_34291);
and U37957 (N_37957,N_35671,N_34341);
xor U37958 (N_37958,N_35663,N_34394);
nor U37959 (N_37959,N_34659,N_35336);
or U37960 (N_37960,N_34062,N_34946);
nor U37961 (N_37961,N_34199,N_35292);
or U37962 (N_37962,N_35961,N_34023);
or U37963 (N_37963,N_35101,N_34878);
nor U37964 (N_37964,N_35668,N_35998);
and U37965 (N_37965,N_35503,N_35039);
nor U37966 (N_37966,N_34062,N_35586);
nor U37967 (N_37967,N_34217,N_35429);
nand U37968 (N_37968,N_34402,N_35717);
nand U37969 (N_37969,N_35406,N_34653);
and U37970 (N_37970,N_35376,N_35051);
xnor U37971 (N_37971,N_35681,N_35034);
or U37972 (N_37972,N_34127,N_35060);
nor U37973 (N_37973,N_35769,N_35868);
nand U37974 (N_37974,N_35098,N_35236);
nor U37975 (N_37975,N_35498,N_35051);
and U37976 (N_37976,N_34710,N_34810);
and U37977 (N_37977,N_34374,N_35805);
xor U37978 (N_37978,N_35106,N_34987);
or U37979 (N_37979,N_35355,N_35689);
xnor U37980 (N_37980,N_35761,N_35019);
nor U37981 (N_37981,N_34632,N_35681);
or U37982 (N_37982,N_35494,N_34233);
or U37983 (N_37983,N_34766,N_35191);
nor U37984 (N_37984,N_34416,N_35864);
nor U37985 (N_37985,N_34754,N_34700);
or U37986 (N_37986,N_35773,N_34755);
and U37987 (N_37987,N_35911,N_35854);
and U37988 (N_37988,N_35201,N_34807);
xor U37989 (N_37989,N_34803,N_34276);
nand U37990 (N_37990,N_35460,N_35269);
and U37991 (N_37991,N_34284,N_35383);
and U37992 (N_37992,N_35296,N_35509);
and U37993 (N_37993,N_35777,N_35025);
or U37994 (N_37994,N_35918,N_34781);
nor U37995 (N_37995,N_35878,N_35512);
or U37996 (N_37996,N_34347,N_35832);
xnor U37997 (N_37997,N_34147,N_35934);
xnor U37998 (N_37998,N_35448,N_34977);
nand U37999 (N_37999,N_35068,N_35925);
nand U38000 (N_38000,N_37083,N_36187);
and U38001 (N_38001,N_37359,N_37935);
or U38002 (N_38002,N_36244,N_36095);
or U38003 (N_38003,N_37126,N_36333);
xnor U38004 (N_38004,N_36625,N_36119);
nor U38005 (N_38005,N_36078,N_37467);
and U38006 (N_38006,N_36050,N_36978);
xnor U38007 (N_38007,N_36169,N_37193);
nand U38008 (N_38008,N_36336,N_37893);
xor U38009 (N_38009,N_36765,N_36622);
nand U38010 (N_38010,N_37332,N_36670);
and U38011 (N_38011,N_37377,N_37975);
and U38012 (N_38012,N_37044,N_37026);
or U38013 (N_38013,N_36129,N_36366);
and U38014 (N_38014,N_36355,N_36111);
nor U38015 (N_38015,N_36387,N_36498);
or U38016 (N_38016,N_37391,N_37829);
nor U38017 (N_38017,N_37498,N_37197);
or U38018 (N_38018,N_37149,N_36928);
nand U38019 (N_38019,N_37061,N_36947);
nand U38020 (N_38020,N_37246,N_36974);
and U38021 (N_38021,N_36584,N_37213);
nand U38022 (N_38022,N_37964,N_36686);
nand U38023 (N_38023,N_36878,N_37606);
or U38024 (N_38024,N_37580,N_37618);
nor U38025 (N_38025,N_37748,N_37469);
nand U38026 (N_38026,N_36077,N_36870);
xor U38027 (N_38027,N_36609,N_36190);
xnor U38028 (N_38028,N_37667,N_36661);
nand U38029 (N_38029,N_37593,N_36473);
nor U38030 (N_38030,N_37774,N_36036);
xnor U38031 (N_38031,N_37992,N_36549);
nor U38032 (N_38032,N_36553,N_37943);
xor U38033 (N_38033,N_36478,N_36486);
nand U38034 (N_38034,N_36463,N_37030);
or U38035 (N_38035,N_36933,N_36304);
nand U38036 (N_38036,N_36967,N_37620);
nor U38037 (N_38037,N_36042,N_37368);
and U38038 (N_38038,N_36955,N_37301);
and U38039 (N_38039,N_36108,N_36721);
and U38040 (N_38040,N_36737,N_36591);
nand U38041 (N_38041,N_36165,N_37437);
nor U38042 (N_38042,N_37412,N_36511);
xnor U38043 (N_38043,N_36127,N_36016);
nor U38044 (N_38044,N_36521,N_37429);
nand U38045 (N_38045,N_37688,N_37942);
or U38046 (N_38046,N_37600,N_36821);
nor U38047 (N_38047,N_37830,N_37940);
and U38048 (N_38048,N_36277,N_36259);
or U38049 (N_38049,N_36262,N_36960);
nand U38050 (N_38050,N_36707,N_37554);
xor U38051 (N_38051,N_37521,N_36233);
nor U38052 (N_38052,N_37537,N_36443);
nand U38053 (N_38053,N_36340,N_37298);
and U38054 (N_38054,N_36230,N_36196);
and U38055 (N_38055,N_37937,N_37608);
and U38056 (N_38056,N_36317,N_36899);
and U38057 (N_38057,N_37109,N_36102);
and U38058 (N_38058,N_37400,N_37591);
or U38059 (N_38059,N_36097,N_36538);
xor U38060 (N_38060,N_37435,N_36871);
xnor U38061 (N_38061,N_36448,N_36866);
nand U38062 (N_38062,N_36432,N_36041);
nand U38063 (N_38063,N_36306,N_36323);
xor U38064 (N_38064,N_37509,N_36717);
nand U38065 (N_38065,N_36950,N_37569);
or U38066 (N_38066,N_37990,N_37443);
and U38067 (N_38067,N_37663,N_36272);
and U38068 (N_38068,N_37764,N_37331);
xor U38069 (N_38069,N_36382,N_36930);
and U38070 (N_38070,N_36483,N_36923);
nand U38071 (N_38071,N_37224,N_37707);
nor U38072 (N_38072,N_36434,N_37392);
and U38073 (N_38073,N_37386,N_37594);
nand U38074 (N_38074,N_37456,N_36994);
or U38075 (N_38075,N_36738,N_36364);
or U38076 (N_38076,N_37320,N_36972);
xor U38077 (N_38077,N_36416,N_37573);
xor U38078 (N_38078,N_36653,N_37635);
or U38079 (N_38079,N_37533,N_37231);
and U38080 (N_38080,N_36384,N_37210);
and U38081 (N_38081,N_37676,N_37963);
nand U38082 (N_38082,N_36959,N_37179);
and U38083 (N_38083,N_37070,N_36507);
nand U38084 (N_38084,N_36912,N_37114);
nand U38085 (N_38085,N_37513,N_37328);
xor U38086 (N_38086,N_36424,N_37903);
or U38087 (N_38087,N_36567,N_37441);
or U38088 (N_38088,N_36598,N_37343);
or U38089 (N_38089,N_36999,N_36203);
nor U38090 (N_38090,N_37334,N_36254);
or U38091 (N_38091,N_36564,N_36793);
nand U38092 (N_38092,N_37326,N_36435);
and U38093 (N_38093,N_37217,N_37819);
xnor U38094 (N_38094,N_37872,N_36734);
and U38095 (N_38095,N_37708,N_36880);
xnor U38096 (N_38096,N_36638,N_36318);
nor U38097 (N_38097,N_36087,N_37852);
xnor U38098 (N_38098,N_36715,N_37712);
xor U38099 (N_38099,N_37578,N_36552);
and U38100 (N_38100,N_36997,N_37789);
xnor U38101 (N_38101,N_37928,N_37455);
nor U38102 (N_38102,N_37877,N_36437);
and U38103 (N_38103,N_36517,N_36695);
and U38104 (N_38104,N_37395,N_36904);
and U38105 (N_38105,N_37837,N_37093);
or U38106 (N_38106,N_36634,N_36338);
and U38107 (N_38107,N_37308,N_37505);
and U38108 (N_38108,N_37751,N_36080);
and U38109 (N_38109,N_36070,N_37589);
nand U38110 (N_38110,N_37651,N_36942);
and U38111 (N_38111,N_37831,N_37011);
and U38112 (N_38112,N_36869,N_37726);
and U38113 (N_38113,N_36520,N_37432);
nor U38114 (N_38114,N_37303,N_37247);
nand U38115 (N_38115,N_37373,N_37120);
nor U38116 (N_38116,N_36966,N_36874);
xor U38117 (N_38117,N_37015,N_37004);
xnor U38118 (N_38118,N_36454,N_36688);
and U38119 (N_38119,N_37727,N_37347);
or U38120 (N_38120,N_37705,N_37849);
nor U38121 (N_38121,N_36969,N_36245);
xnor U38122 (N_38122,N_37188,N_37010);
or U38123 (N_38123,N_36587,N_37183);
and U38124 (N_38124,N_36404,N_36510);
xor U38125 (N_38125,N_37911,N_37826);
or U38126 (N_38126,N_36133,N_36479);
or U38127 (N_38127,N_37507,N_37912);
or U38128 (N_38128,N_36680,N_36894);
xnor U38129 (N_38129,N_37960,N_37613);
or U38130 (N_38130,N_36815,N_36291);
nor U38131 (N_38131,N_37192,N_37427);
nand U38132 (N_38132,N_37257,N_36065);
nor U38133 (N_38133,N_36181,N_36716);
or U38134 (N_38134,N_36768,N_36832);
nand U38135 (N_38135,N_36032,N_37158);
or U38136 (N_38136,N_36692,N_36147);
nand U38137 (N_38137,N_37581,N_37187);
nor U38138 (N_38138,N_37460,N_36615);
xnor U38139 (N_38139,N_37348,N_37772);
xnor U38140 (N_38140,N_36548,N_37746);
and U38141 (N_38141,N_36683,N_36410);
or U38142 (N_38142,N_37218,N_36005);
nand U38143 (N_38143,N_37492,N_37865);
nand U38144 (N_38144,N_36423,N_36412);
nand U38145 (N_38145,N_37627,N_36140);
and U38146 (N_38146,N_36013,N_37756);
and U38147 (N_38147,N_37933,N_37622);
nand U38148 (N_38148,N_37290,N_37049);
nor U38149 (N_38149,N_37922,N_37761);
nor U38150 (N_38150,N_36636,N_37067);
nand U38151 (N_38151,N_37814,N_36892);
xnor U38152 (N_38152,N_37272,N_37662);
and U38153 (N_38153,N_37861,N_37486);
xor U38154 (N_38154,N_37110,N_37833);
and U38155 (N_38155,N_36698,N_36575);
or U38156 (N_38156,N_37767,N_37987);
or U38157 (N_38157,N_36009,N_37869);
and U38158 (N_38158,N_36319,N_36544);
nand U38159 (N_38159,N_36195,N_36727);
or U38160 (N_38160,N_36945,N_36038);
and U38161 (N_38161,N_37967,N_37068);
nand U38162 (N_38162,N_36913,N_36864);
or U38163 (N_38163,N_36808,N_36503);
and U38164 (N_38164,N_37932,N_36565);
nand U38165 (N_38165,N_37019,N_37677);
or U38166 (N_38166,N_36986,N_36153);
xor U38167 (N_38167,N_37471,N_37512);
or U38168 (N_38168,N_37804,N_37057);
xnor U38169 (N_38169,N_37559,N_37151);
xor U38170 (N_38170,N_37838,N_36497);
and U38171 (N_38171,N_37240,N_36281);
nor U38172 (N_38172,N_36058,N_36215);
or U38173 (N_38173,N_37071,N_37478);
nand U38174 (N_38174,N_36266,N_37549);
xor U38175 (N_38175,N_37802,N_36173);
nor U38176 (N_38176,N_36441,N_37863);
and U38177 (N_38177,N_36535,N_36946);
or U38178 (N_38178,N_37292,N_36392);
and U38179 (N_38179,N_36916,N_37371);
nor U38180 (N_38180,N_37502,N_36977);
nor U38181 (N_38181,N_37884,N_37982);
xnor U38182 (N_38182,N_37695,N_37939);
and U38183 (N_38183,N_36436,N_36818);
nand U38184 (N_38184,N_37989,N_36360);
nand U38185 (N_38185,N_37646,N_36971);
nor U38186 (N_38186,N_37132,N_36571);
or U38187 (N_38187,N_37853,N_37166);
xor U38188 (N_38188,N_37462,N_37641);
nand U38189 (N_38189,N_37858,N_37379);
nand U38190 (N_38190,N_36865,N_37031);
and U38191 (N_38191,N_37144,N_37546);
nand U38192 (N_38192,N_37557,N_37261);
or U38193 (N_38193,N_37353,N_37730);
nand U38194 (N_38194,N_36543,N_36143);
and U38195 (N_38195,N_36027,N_36430);
xnor U38196 (N_38196,N_37882,N_37946);
nor U38197 (N_38197,N_37545,N_36561);
xor U38198 (N_38198,N_36607,N_36170);
xor U38199 (N_38199,N_36316,N_37765);
or U38200 (N_38200,N_36491,N_36643);
xnor U38201 (N_38201,N_36624,N_37121);
nor U38202 (N_38202,N_37785,N_37307);
or U38203 (N_38203,N_37464,N_37983);
nor U38204 (N_38204,N_36773,N_36938);
or U38205 (N_38205,N_37895,N_37926);
nand U38206 (N_38206,N_37856,N_36784);
or U38207 (N_38207,N_36646,N_36590);
xor U38208 (N_38208,N_36176,N_36677);
nor U38209 (N_38209,N_36699,N_37344);
nor U38210 (N_38210,N_36458,N_36171);
nor U38211 (N_38211,N_37384,N_36779);
nor U38212 (N_38212,N_37526,N_36370);
or U38213 (N_38213,N_36008,N_36706);
xor U38214 (N_38214,N_37040,N_37354);
or U38215 (N_38215,N_37757,N_37609);
nand U38216 (N_38216,N_37104,N_37283);
nor U38217 (N_38217,N_36332,N_37191);
or U38218 (N_38218,N_36081,N_36834);
and U38219 (N_38219,N_37686,N_36246);
or U38220 (N_38220,N_36123,N_37419);
or U38221 (N_38221,N_36684,N_36903);
nand U38222 (N_38222,N_36307,N_36858);
or U38223 (N_38223,N_36121,N_36528);
xor U38224 (N_38224,N_36885,N_37080);
nand U38225 (N_38225,N_36512,N_36192);
nand U38226 (N_38226,N_37571,N_37153);
nor U38227 (N_38227,N_36714,N_37342);
xnor U38228 (N_38228,N_37986,N_36341);
and U38229 (N_38229,N_37938,N_37793);
or U38230 (N_38230,N_36264,N_36073);
nor U38231 (N_38231,N_36461,N_36194);
or U38232 (N_38232,N_37434,N_37178);
and U38233 (N_38233,N_36944,N_36700);
xor U38234 (N_38234,N_37491,N_37143);
and U38235 (N_38235,N_37925,N_36848);
xor U38236 (N_38236,N_36372,N_37945);
nand U38237 (N_38237,N_37703,N_36618);
nand U38238 (N_38238,N_36172,N_36481);
nor U38239 (N_38239,N_36248,N_37115);
and U38240 (N_38240,N_36285,N_37020);
xnor U38241 (N_38241,N_36130,N_36149);
and U38242 (N_38242,N_37604,N_36592);
nand U38243 (N_38243,N_37993,N_37484);
and U38244 (N_38244,N_36811,N_37846);
and U38245 (N_38245,N_37776,N_37979);
nand U38246 (N_38246,N_36347,N_37485);
xnor U38247 (N_38247,N_36787,N_37225);
xor U38248 (N_38248,N_37198,N_37710);
and U38249 (N_38249,N_36827,N_36019);
or U38250 (N_38250,N_37250,N_36952);
nand U38251 (N_38251,N_37397,N_36676);
nor U38252 (N_38252,N_37661,N_37184);
nand U38253 (N_38253,N_36740,N_37605);
xor U38254 (N_38254,N_37452,N_37162);
xnor U38255 (N_38255,N_36791,N_37066);
and U38256 (N_38256,N_37901,N_36589);
and U38257 (N_38257,N_37466,N_36105);
and U38258 (N_38258,N_36061,N_36506);
and U38259 (N_38259,N_36996,N_36284);
or U38260 (N_38260,N_36722,N_36305);
nand U38261 (N_38261,N_36515,N_37001);
xnor U38262 (N_38262,N_37823,N_37547);
or U38263 (N_38263,N_36949,N_36600);
xnor U38264 (N_38264,N_37836,N_36413);
nor U38265 (N_38265,N_37269,N_36447);
nor U38266 (N_38266,N_36719,N_37064);
or U38267 (N_38267,N_37273,N_36691);
xor U38268 (N_38268,N_37442,N_36909);
nor U38269 (N_38269,N_37255,N_37540);
nor U38270 (N_38270,N_37750,N_36359);
xor U38271 (N_38271,N_36045,N_36369);
and U38272 (N_38272,N_36539,N_36229);
or U38273 (N_38273,N_37039,N_37025);
nand U38274 (N_38274,N_37725,N_37116);
or U38275 (N_38275,N_37382,N_36362);
nor U38276 (N_38276,N_36635,N_36872);
or U38277 (N_38277,N_37014,N_37806);
nor U38278 (N_38278,N_37470,N_36242);
or U38279 (N_38279,N_37024,N_36154);
or U38280 (N_38280,N_36380,N_36725);
or U38281 (N_38281,N_37504,N_37367);
or U38282 (N_38282,N_36802,N_36099);
xnor U38283 (N_38283,N_36139,N_36315);
and U38284 (N_38284,N_36729,N_36752);
or U38285 (N_38285,N_36619,N_37062);
nor U38286 (N_38286,N_37032,N_36024);
or U38287 (N_38287,N_36429,N_37438);
nand U38288 (N_38288,N_36534,N_37917);
nand U38289 (N_38289,N_36975,N_36137);
nand U38290 (N_38290,N_36720,N_36496);
xnor U38291 (N_38291,N_36225,N_37864);
and U38292 (N_38292,N_36251,N_36325);
or U38293 (N_38293,N_36274,N_36446);
nor U38294 (N_38294,N_37998,N_37668);
xnor U38295 (N_38295,N_37468,N_37200);
and U38296 (N_38296,N_36605,N_37490);
and U38297 (N_38297,N_37634,N_36217);
xor U38298 (N_38298,N_36993,N_37848);
xnor U38299 (N_38299,N_36043,N_37127);
nor U38300 (N_38300,N_37684,N_37295);
nor U38301 (N_38301,N_37820,N_36354);
nor U38302 (N_38302,N_37189,N_37795);
nand U38303 (N_38303,N_36182,N_37107);
nor U38304 (N_38304,N_36125,N_37665);
and U38305 (N_38305,N_37131,N_37159);
and U38306 (N_38306,N_36457,N_37897);
xor U38307 (N_38307,N_37532,N_36569);
nand U38308 (N_38308,N_36898,N_36141);
nor U38309 (N_38309,N_36351,N_36184);
xor U38310 (N_38310,N_37284,N_37916);
xnor U38311 (N_38311,N_37601,N_37422);
or U38312 (N_38312,N_36557,N_36376);
nand U38313 (N_38313,N_37561,N_37313);
xor U38314 (N_38314,N_37381,N_36365);
xnor U38315 (N_38315,N_37799,N_36921);
or U38316 (N_38316,N_36985,N_36260);
nor U38317 (N_38317,N_37421,N_36053);
xnor U38318 (N_38318,N_36201,N_37973);
nand U38319 (N_38319,N_37161,N_37568);
nor U38320 (N_38320,N_36335,N_36326);
nand U38321 (N_38321,N_36243,N_37670);
xnor U38322 (N_38322,N_37517,N_37102);
and U38323 (N_38323,N_37645,N_36951);
xnor U38324 (N_38324,N_36389,N_36179);
xor U38325 (N_38325,N_37649,N_37385);
nand U38326 (N_38326,N_37275,N_36614);
nand U38327 (N_38327,N_36218,N_37553);
xor U38328 (N_38328,N_36420,N_36263);
nand U38329 (N_38329,N_36357,N_37274);
xor U38330 (N_38330,N_36442,N_37245);
xnor U38331 (N_38331,N_37163,N_37000);
nor U38332 (N_38332,N_36532,N_37124);
nand U38333 (N_38333,N_36499,N_37418);
nor U38334 (N_38334,N_36748,N_36232);
nand U38335 (N_38335,N_36428,N_36956);
nor U38336 (N_38336,N_36227,N_37828);
nand U38337 (N_38337,N_37075,N_37660);
nor U38338 (N_38338,N_36112,N_36785);
nor U38339 (N_38339,N_37253,N_36749);
nand U38340 (N_38340,N_36018,N_37630);
or U38341 (N_38341,N_37914,N_37415);
nor U38342 (N_38342,N_36675,N_36597);
nor U38343 (N_38343,N_36156,N_37278);
xnor U38344 (N_38344,N_37542,N_36488);
xor U38345 (N_38345,N_36900,N_37248);
nand U38346 (N_38346,N_36550,N_37790);
nor U38347 (N_38347,N_37244,N_36697);
or U38348 (N_38348,N_36069,N_37094);
nand U38349 (N_38349,N_37207,N_37874);
xor U38350 (N_38350,N_37216,N_37675);
or U38351 (N_38351,N_36519,N_36378);
xor U38352 (N_38352,N_36085,N_37165);
or U38353 (N_38353,N_37722,N_36665);
and U38354 (N_38354,N_36200,N_36160);
nand U38355 (N_38355,N_37324,N_37862);
nand U38356 (N_38356,N_37461,N_36462);
nand U38357 (N_38357,N_37739,N_36982);
xor U38358 (N_38358,N_36186,N_36627);
nand U38359 (N_38359,N_37402,N_36732);
or U38360 (N_38360,N_37205,N_37597);
xnor U38361 (N_38361,N_37779,N_37735);
xnor U38362 (N_38362,N_37088,N_37868);
nor U38363 (N_38363,N_37185,N_37976);
or U38364 (N_38364,N_37694,N_36470);
nand U38365 (N_38365,N_37626,N_36300);
and U38366 (N_38366,N_36604,N_36480);
nor U38367 (N_38367,N_37232,N_37807);
or U38368 (N_38368,N_37560,N_37587);
and U38369 (N_38369,N_36792,N_37749);
xnor U38370 (N_38370,N_37747,N_36261);
or U38371 (N_38371,N_36219,N_36174);
nor U38372 (N_38372,N_37832,N_37439);
nor U38373 (N_38373,N_36493,N_36025);
or U38374 (N_38374,N_36958,N_36014);
nor U38375 (N_38375,N_36303,N_37296);
xor U38376 (N_38376,N_36422,N_37805);
or U38377 (N_38377,N_37566,N_37514);
xor U38378 (N_38378,N_37155,N_36175);
xor U38379 (N_38379,N_36066,N_36690);
nand U38380 (N_38380,N_36595,N_36155);
or U38381 (N_38381,N_36456,N_37376);
nor U38382 (N_38382,N_36757,N_36213);
and U38383 (N_38383,N_36823,N_37564);
nor U38384 (N_38384,N_36761,N_36556);
nand U38385 (N_38385,N_37936,N_36396);
or U38386 (N_38386,N_36957,N_36011);
nor U38387 (N_38387,N_37584,N_37523);
and U38388 (N_38388,N_37425,N_37125);
or U38389 (N_38389,N_36852,N_37101);
nor U38390 (N_38390,N_37175,N_36295);
nor U38391 (N_38391,N_36199,N_36208);
nand U38392 (N_38392,N_36373,N_36702);
and U38393 (N_38393,N_36650,N_36588);
xor U38394 (N_38394,N_37366,N_36726);
or U38395 (N_38395,N_37007,N_37129);
nand U38396 (N_38396,N_37798,N_37238);
or U38397 (N_38397,N_36735,N_37628);
nor U38398 (N_38398,N_36703,N_36875);
or U38399 (N_38399,N_36788,N_36193);
nor U38400 (N_38400,N_36953,N_36256);
nor U38401 (N_38401,N_37731,N_37906);
or U38402 (N_38402,N_37632,N_37815);
nor U38403 (N_38403,N_36574,N_37276);
nor U38404 (N_38404,N_37704,N_36599);
or U38405 (N_38405,N_36881,N_37022);
nand U38406 (N_38406,N_36161,N_37541);
or U38407 (N_38407,N_37154,N_36640);
nand U38408 (N_38408,N_37528,N_36980);
nand U38409 (N_38409,N_37265,N_36158);
nand U38410 (N_38410,N_37590,N_36585);
nand U38411 (N_38411,N_36390,N_36508);
and U38412 (N_38412,N_37291,N_37433);
nand U38413 (N_38413,N_37881,N_37350);
and U38414 (N_38414,N_36465,N_36891);
nor U38415 (N_38415,N_36288,N_36138);
xnor U38416 (N_38416,N_37664,N_37956);
nor U38417 (N_38417,N_36144,N_37574);
nor U38418 (N_38418,N_37562,N_36466);
xnor U38419 (N_38419,N_36122,N_36253);
and U38420 (N_38420,N_37235,N_36915);
nand U38421 (N_38421,N_36501,N_37357);
nor U38422 (N_38422,N_37319,N_36596);
xnor U38423 (N_38423,N_36067,N_36107);
or U38424 (N_38424,N_37902,N_37745);
nor U38425 (N_38425,N_37317,N_37219);
or U38426 (N_38426,N_37074,N_37171);
or U38427 (N_38427,N_37929,N_36083);
xor U38428 (N_38428,N_37968,N_36271);
or U38429 (N_38429,N_37648,N_37034);
or U38430 (N_38430,N_37413,N_37279);
and U38431 (N_38431,N_37136,N_36135);
or U38432 (N_38432,N_37592,N_37984);
or U38433 (N_38433,N_37369,N_36555);
xnor U38434 (N_38434,N_37714,N_36022);
and U38435 (N_38435,N_36838,N_36003);
xor U38436 (N_38436,N_37612,N_37302);
and U38437 (N_38437,N_37122,N_37787);
and U38438 (N_38438,N_37174,N_37777);
nor U38439 (N_38439,N_36418,N_36252);
and U38440 (N_38440,N_37991,N_36001);
nor U38441 (N_38441,N_37203,N_36642);
or U38442 (N_38442,N_36131,N_37408);
nand U38443 (N_38443,N_36940,N_37969);
or U38444 (N_38444,N_36770,N_37729);
nor U38445 (N_38445,N_36536,N_36082);
nand U38446 (N_38446,N_37380,N_36055);
nand U38447 (N_38447,N_36917,N_37519);
nand U38448 (N_38448,N_36835,N_37794);
or U38449 (N_38449,N_36983,N_37293);
and U38450 (N_38450,N_37647,N_36659);
and U38451 (N_38451,N_36270,N_37315);
nor U38452 (N_38452,N_37222,N_36710);
nor U38453 (N_38453,N_36918,N_37840);
or U38454 (N_38454,N_37653,N_36603);
or U38455 (N_38455,N_37337,N_37268);
nand U38456 (N_38456,N_36103,N_37891);
or U38457 (N_38457,N_37176,N_37899);
xnor U38458 (N_38458,N_36731,N_36492);
and U38459 (N_38459,N_37711,N_37643);
xor U38460 (N_38460,N_36017,N_36746);
nor U38461 (N_38461,N_36920,N_36455);
and U38462 (N_38462,N_37199,N_36494);
or U38463 (N_38463,N_37781,N_36398);
or U38464 (N_38464,N_36267,N_36623);
xor U38465 (N_38465,N_36612,N_36469);
nand U38466 (N_38466,N_37954,N_37017);
nor U38467 (N_38467,N_36568,N_36693);
and U38468 (N_38468,N_37409,N_36778);
xor U38469 (N_38469,N_37878,N_37078);
nand U38470 (N_38470,N_37538,N_37550);
or U38471 (N_38471,N_36766,N_36216);
nand U38472 (N_38472,N_37423,N_37842);
nand U38473 (N_38473,N_36400,N_36884);
xor U38474 (N_38474,N_37894,N_36157);
nand U38475 (N_38475,N_36651,N_37416);
or U38476 (N_38476,N_37041,N_37281);
or U38477 (N_38477,N_36268,N_37812);
nand U38478 (N_38478,N_36617,N_36177);
or U38479 (N_38479,N_37038,N_36393);
xnor U38480 (N_38480,N_36411,N_36724);
and U38481 (N_38481,N_37841,N_37732);
nand U38482 (N_38482,N_36628,N_36460);
nor U38483 (N_38483,N_37363,N_36468);
and U38484 (N_38484,N_36180,N_37195);
xor U38485 (N_38485,N_36391,N_36763);
nand U38486 (N_38486,N_36386,N_36113);
xnor U38487 (N_38487,N_36321,N_37754);
nand U38488 (N_38488,N_36124,N_37843);
nor U38489 (N_38489,N_37839,N_36514);
xnor U38490 (N_38490,N_37476,N_36361);
or U38491 (N_38491,N_36901,N_37500);
xor U38492 (N_38492,N_37631,N_36010);
nand U38493 (N_38493,N_37113,N_36753);
nand U38494 (N_38494,N_36126,N_36367);
nand U38495 (N_38495,N_36128,N_37005);
and U38496 (N_38496,N_36862,N_37702);
and U38497 (N_38497,N_36795,N_36664);
xnor U38498 (N_38498,N_37771,N_37866);
or U38499 (N_38499,N_36718,N_36836);
nand U38500 (N_38500,N_37105,N_37316);
nor U38501 (N_38501,N_36562,N_37339);
nand U38502 (N_38502,N_36527,N_36150);
nand U38503 (N_38503,N_37403,N_37170);
or U38504 (N_38504,N_36772,N_36089);
and U38505 (N_38505,N_37314,N_37027);
nor U38506 (N_38506,N_36762,N_37322);
or U38507 (N_38507,N_36712,N_36035);
nand U38508 (N_38508,N_36101,N_37006);
nor U38509 (N_38509,N_37106,N_37908);
xor U38510 (N_38510,N_37152,N_36526);
and U38511 (N_38511,N_37055,N_36758);
nand U38512 (N_38512,N_37249,N_37698);
and U38513 (N_38513,N_37778,N_37050);
and U38514 (N_38514,N_37800,N_36188);
and U38515 (N_38515,N_36626,N_36805);
xor U38516 (N_38516,N_36037,N_36908);
and U38517 (N_38517,N_36343,N_37012);
nand U38518 (N_38518,N_37305,N_36681);
and U38519 (N_38519,N_36976,N_36610);
nand U38520 (N_38520,N_36385,N_37097);
and U38521 (N_38521,N_36547,N_36641);
xnor U38522 (N_38522,N_37090,N_37657);
nand U38523 (N_38523,N_37845,N_36110);
xnor U38524 (N_38524,N_37388,N_37548);
nor U38525 (N_38525,N_37565,N_36166);
nor U38526 (N_38526,N_37228,N_37060);
nor U38527 (N_38527,N_37780,N_37607);
nand U38528 (N_38528,N_37576,N_36839);
nor U38529 (N_38529,N_37023,N_36667);
nor U38530 (N_38530,N_37970,N_36408);
xnor U38531 (N_38531,N_37980,N_37924);
nor U38532 (N_38532,N_37073,N_37365);
xor U38533 (N_38533,N_36476,N_37656);
and U38534 (N_38534,N_37134,N_37048);
and U38535 (N_38535,N_36583,N_36941);
and U38536 (N_38536,N_36563,N_36397);
nor U38537 (N_38537,N_36849,N_37720);
and U38538 (N_38538,N_37742,N_37818);
nand U38539 (N_38539,N_36450,N_36100);
nor U38540 (N_38540,N_37687,N_37614);
nor U38541 (N_38541,N_36647,N_36666);
nand U38542 (N_38542,N_36525,N_36352);
nor U38543 (N_38543,N_36383,N_36231);
nor U38544 (N_38544,N_37312,N_36705);
or U38545 (N_38545,N_36669,N_37602);
nand U38546 (N_38546,N_36308,N_36220);
nand U38547 (N_38547,N_37959,N_37997);
nand U38548 (N_38548,N_36649,N_37016);
or U38549 (N_38549,N_37139,N_37721);
xnor U38550 (N_38550,N_37516,N_36132);
or U38551 (N_38551,N_36006,N_37428);
nor U38552 (N_38552,N_37280,N_37529);
nor U38553 (N_38553,N_36897,N_37890);
and U38554 (N_38554,N_37510,N_36485);
or U38555 (N_38555,N_36629,N_36353);
xor U38556 (N_38556,N_37563,N_37743);
or U38557 (N_38557,N_36048,N_37518);
nor U38558 (N_38558,N_37511,N_36541);
nand U38559 (N_38559,N_36970,N_37208);
and U38560 (N_38560,N_36687,N_36283);
or U38561 (N_38561,N_36730,N_36205);
or U38562 (N_38562,N_37503,N_37458);
and U38563 (N_38563,N_37681,N_37311);
nand U38564 (N_38564,N_36368,N_36222);
xor U38565 (N_38565,N_37595,N_37002);
nor U38566 (N_38566,N_37850,N_37262);
nand U38567 (N_38567,N_37059,N_36639);
and U38568 (N_38568,N_37029,N_36350);
xnor U38569 (N_38569,N_37362,N_37133);
or U38570 (N_38570,N_37459,N_36533);
nor U38571 (N_38571,N_36831,N_36068);
nand U38572 (N_38572,N_37543,N_36433);
and U38573 (N_38573,N_37209,N_36118);
and U38574 (N_38574,N_36755,N_36342);
and U38575 (N_38575,N_36459,N_36302);
or U38576 (N_38576,N_37069,N_37372);
or U38577 (N_38577,N_37333,N_37915);
xor U38578 (N_38578,N_36586,N_37449);
and U38579 (N_38579,N_37552,N_37880);
or U38580 (N_38580,N_36374,N_36671);
xnor U38581 (N_38581,N_36346,N_36210);
or U38582 (N_38582,N_36747,N_36109);
and U38583 (N_38583,N_37555,N_37671);
nand U38584 (N_38584,N_36882,N_37259);
and U38585 (N_38585,N_37375,N_36551);
nand U38586 (N_38586,N_36240,N_37446);
and U38587 (N_38587,N_37360,N_36804);
xnor U38588 (N_38588,N_36577,N_36250);
nor U38589 (N_38589,N_37346,N_37451);
xnor U38590 (N_38590,N_36120,N_36086);
or U38591 (N_38591,N_37962,N_36255);
nand U38592 (N_38592,N_36324,N_37762);
nand U38593 (N_38593,N_36637,N_36988);
and U38594 (N_38594,N_37018,N_37483);
or U38595 (N_38595,N_37824,N_36701);
xor U38596 (N_38596,N_36911,N_37407);
or U38597 (N_38597,N_36782,N_37625);
nor U38598 (N_38598,N_37410,N_37585);
nor U38599 (N_38599,N_37855,N_36464);
or U38600 (N_38600,N_37196,N_37264);
xor U38601 (N_38601,N_36769,N_37411);
xor U38602 (N_38602,N_36294,N_37300);
xnor U38603 (N_38603,N_37957,N_37194);
nand U38604 (N_38604,N_37474,N_37118);
nor U38605 (N_38605,N_37616,N_37639);
nand U38606 (N_38606,N_36846,N_37642);
or U38607 (N_38607,N_36445,N_37907);
xnor U38608 (N_38608,N_37782,N_37770);
and U38609 (N_38609,N_37629,N_37190);
xnor U38610 (N_38610,N_36924,N_36363);
or U38611 (N_38611,N_37898,N_37436);
xnor U38612 (N_38612,N_37242,N_36523);
or U38613 (N_38613,N_37008,N_37572);
xnor U38614 (N_38614,N_36876,N_36906);
and U38615 (N_38615,N_36709,N_36269);
or U38616 (N_38616,N_36033,N_36414);
nand U38617 (N_38617,N_37733,N_36672);
xnor U38618 (N_38618,N_36685,N_36682);
or U38619 (N_38619,N_37146,N_36399);
nand U38620 (N_38620,N_36968,N_37691);
nand U38621 (N_38621,N_36580,N_37389);
xor U38622 (N_38622,N_36075,N_36910);
or U38623 (N_38623,N_36490,N_37558);
nor U38624 (N_38624,N_37496,N_37028);
and U38625 (N_38625,N_36853,N_37239);
nor U38626 (N_38626,N_37336,N_36301);
or U38627 (N_38627,N_36883,N_37145);
xor U38628 (N_38628,N_36799,N_37965);
nor U38629 (N_38629,N_37150,N_37230);
and U38630 (N_38630,N_37501,N_37482);
and U38631 (N_38631,N_36237,N_37130);
nand U38632 (N_38632,N_36039,N_36998);
or U38633 (N_38633,N_36152,N_36789);
xor U38634 (N_38634,N_36062,N_37909);
or U38635 (N_38635,N_37755,N_37450);
or U38636 (N_38636,N_36334,N_37556);
nand U38637 (N_38637,N_36648,N_37457);
and U38638 (N_38638,N_37052,N_36760);
nor U38639 (N_38639,N_36888,N_36057);
xor U38640 (N_38640,N_37644,N_37141);
and U38641 (N_38641,N_36890,N_37974);
and U38642 (N_38642,N_37495,N_36224);
nand U38643 (N_38643,N_36954,N_37904);
nor U38644 (N_38644,N_36847,N_37065);
xnor U38645 (N_38645,N_36987,N_37215);
and U38646 (N_38646,N_36658,N_36026);
or U38647 (N_38647,N_36403,N_37816);
nand U38648 (N_38648,N_37575,N_36265);
nor U38649 (N_38649,N_37766,N_37111);
xnor U38650 (N_38650,N_36516,N_37157);
and U38651 (N_38651,N_37267,N_37091);
xor U38652 (N_38652,N_36020,N_36504);
and U38653 (N_38653,N_36209,N_36178);
xnor U38654 (N_38654,N_37857,N_37696);
or U38655 (N_38655,N_36495,N_37669);
or U38656 (N_38656,N_37988,N_37844);
xor U38657 (N_38657,N_36886,N_37237);
xnor U38658 (N_38658,N_37534,N_36239);
nor U38659 (N_38659,N_37092,N_36965);
and U38660 (N_38660,N_37737,N_36674);
xnor U38661 (N_38661,N_36046,N_37393);
and U38662 (N_38662,N_37325,N_36092);
nor U38663 (N_38663,N_36711,N_36162);
and U38664 (N_38664,N_36223,N_36708);
or U38665 (N_38665,N_37256,N_37035);
and U38666 (N_38666,N_37678,N_37889);
xnor U38667 (N_38667,N_36837,N_36631);
and U38668 (N_38668,N_37081,N_36927);
nand U38669 (N_38669,N_36925,N_37481);
nand U38670 (N_38670,N_37769,N_37426);
nor U38671 (N_38671,N_36198,N_37900);
nor U38672 (N_38672,N_37586,N_37356);
nand U38673 (N_38673,N_37021,N_37921);
and U38674 (N_38674,N_36863,N_37148);
or U38675 (N_38675,N_36893,N_36328);
and U38676 (N_38676,N_37420,N_37709);
xnor U38677 (N_38677,N_37086,N_37716);
nand U38678 (N_38678,N_36601,N_37699);
xor U38679 (N_38679,N_37615,N_37637);
or U38680 (N_38680,N_37531,N_37489);
nand U38681 (N_38681,N_36273,N_36134);
nand U38682 (N_38682,N_36421,N_37285);
xor U38683 (N_38683,N_37827,N_36820);
xor U38684 (N_38684,N_37119,N_36961);
nand U38685 (N_38685,N_36299,N_36207);
nor U38686 (N_38686,N_37251,N_36992);
nand U38687 (N_38687,N_36312,N_37655);
nor U38688 (N_38688,N_36331,N_36657);
xor U38689 (N_38689,N_37431,N_36214);
or U38690 (N_38690,N_36047,N_36051);
xor U38691 (N_38691,N_37221,N_37045);
and U38692 (N_38692,N_37335,N_37596);
or U38693 (N_38693,N_36513,N_37544);
nor U38694 (N_38694,N_37768,N_36091);
or U38695 (N_38695,N_36015,N_36750);
or U38696 (N_38696,N_37142,N_36206);
xnor U38697 (N_38697,N_37042,N_36375);
or U38698 (N_38698,N_36475,N_37744);
xnor U38699 (N_38699,N_36696,N_37477);
nand U38700 (N_38700,N_37896,N_37211);
xor U38701 (N_38701,N_37784,N_36522);
and U38702 (N_38702,N_36293,N_37650);
or U38703 (N_38703,N_36867,N_37673);
or U38704 (N_38704,N_37652,N_36228);
and U38705 (N_38705,N_36877,N_36191);
and U38706 (N_38706,N_36425,N_37994);
xnor U38707 (N_38707,N_37349,N_37463);
and U38708 (N_38708,N_36939,N_37736);
nand U38709 (N_38709,N_36402,N_36406);
nand U38710 (N_38710,N_36236,N_37289);
nor U38711 (N_38711,N_37610,N_37404);
xor U38712 (N_38712,N_36775,N_36327);
and U38713 (N_38713,N_37445,N_36136);
or U38714 (N_38714,N_36477,N_37266);
or U38715 (N_38715,N_36645,N_36907);
nand U38716 (N_38716,N_37233,N_36056);
xnor U38717 (N_38717,N_36573,N_36142);
and U38718 (N_38718,N_36286,N_36502);
xor U38719 (N_38719,N_36345,N_36467);
nor U38720 (N_38720,N_37082,N_37697);
nor U38721 (N_38721,N_37524,N_36474);
and U38722 (N_38722,N_36790,N_37103);
xnor U38723 (N_38723,N_36440,N_37520);
xnor U38724 (N_38724,N_37417,N_37879);
or U38725 (N_38725,N_36509,N_37582);
and U38726 (N_38726,N_37883,N_37085);
nor U38727 (N_38727,N_37623,N_36545);
nand U38728 (N_38728,N_36800,N_36887);
xnor U38729 (N_38729,N_37345,N_36146);
nand U38730 (N_38730,N_37394,N_37223);
and U38731 (N_38731,N_36531,N_37260);
nand U38732 (N_38732,N_36819,N_36829);
nor U38733 (N_38733,N_37341,N_37297);
or U38734 (N_38734,N_36540,N_37058);
nand U38735 (N_38735,N_37941,N_37598);
xnor U38736 (N_38736,N_36654,N_37723);
or U38737 (N_38737,N_36662,N_36310);
xor U38738 (N_38738,N_37947,N_36290);
and U38739 (N_38739,N_37084,N_37488);
and U38740 (N_38740,N_36560,N_37801);
or U38741 (N_38741,N_37287,N_37870);
or U38742 (N_38742,N_36922,N_36159);
nor U38743 (N_38743,N_36028,N_37934);
or U38744 (N_38744,N_36023,N_36419);
or U38745 (N_38745,N_36007,N_37791);
and U38746 (N_38746,N_37728,N_37783);
nor U38747 (N_38747,N_36409,N_37658);
xor U38748 (N_38748,N_36322,N_37603);
nand U38749 (N_38749,N_37633,N_37168);
nor U38750 (N_38750,N_36164,N_36962);
nand U38751 (N_38751,N_37810,N_36744);
xnor U38752 (N_38752,N_37885,N_36741);
xor U38753 (N_38753,N_36489,N_36660);
nor U38754 (N_38754,N_37920,N_37961);
xor U38755 (N_38755,N_36449,N_37398);
or U38756 (N_38756,N_36349,N_36090);
or U38757 (N_38757,N_37330,N_36487);
or U38758 (N_38758,N_37876,N_37690);
and U38759 (N_38759,N_37822,N_36850);
or U38760 (N_38760,N_36163,N_36117);
nand U38761 (N_38761,N_36578,N_37719);
nor U38762 (N_38762,N_36825,N_37679);
nor U38763 (N_38763,N_37715,N_37977);
xnor U38764 (N_38764,N_36739,N_37046);
xnor U38765 (N_38765,N_36049,N_36311);
or U38766 (N_38766,N_37948,N_36937);
nand U38767 (N_38767,N_37304,N_37072);
nand U38768 (N_38768,N_36963,N_37919);
nor U38769 (N_38769,N_37972,N_36767);
nor U38770 (N_38770,N_37364,N_36797);
xnor U38771 (N_38771,N_37910,N_36751);
nand U38772 (N_38772,N_37995,N_36742);
xor U38773 (N_38773,N_37813,N_36777);
or U38774 (N_38774,N_36873,N_36990);
xnor U38775 (N_38775,N_37424,N_37033);
or U38776 (N_38776,N_37738,N_36379);
xor U38777 (N_38777,N_37351,N_36071);
or U38778 (N_38778,N_37201,N_37212);
nor U38779 (N_38779,N_37243,N_36500);
or U38780 (N_38780,N_36063,N_37525);
nor U38781 (N_38781,N_37009,N_37137);
nor U38782 (N_38782,N_36822,N_36774);
nor U38783 (N_38783,N_36611,N_37619);
xnor U38784 (N_38784,N_37172,N_37108);
or U38785 (N_38785,N_36842,N_36570);
or U38786 (N_38786,N_37204,N_36830);
nor U38787 (N_38787,N_37138,N_36934);
nand U38788 (N_38788,N_37636,N_36401);
nor U38789 (N_38789,N_36620,N_36258);
and U38790 (N_38790,N_37803,N_37825);
and U38791 (N_38791,N_36358,N_37047);
and U38792 (N_38792,N_36084,N_36926);
nand U38793 (N_38793,N_36096,N_37788);
nor U38794 (N_38794,N_36914,N_37966);
and U38795 (N_38795,N_36796,N_37487);
and U38796 (N_38796,N_37128,N_37123);
or U38797 (N_38797,N_37399,N_37506);
or U38798 (N_38798,N_36803,N_36104);
or U38799 (N_38799,N_36764,N_37792);
nand U38800 (N_38800,N_37234,N_37753);
or U38801 (N_38801,N_37054,N_37508);
and U38802 (N_38802,N_36613,N_37288);
and U38803 (N_38803,N_36896,N_36833);
xnor U38804 (N_38804,N_36844,N_37773);
nor U38805 (N_38805,N_37430,N_36320);
nor U38806 (N_38806,N_37286,N_36012);
or U38807 (N_38807,N_37051,N_37087);
and U38808 (N_38808,N_36518,N_37227);
or U38809 (N_38809,N_37775,N_36608);
nand U38810 (N_38810,N_36197,N_36115);
or U38811 (N_38811,N_37321,N_37270);
or U38812 (N_38812,N_36948,N_36030);
xnor U38813 (N_38813,N_36652,N_36581);
nand U38814 (N_38814,N_37859,N_36812);
and U38815 (N_38815,N_36807,N_36704);
and U38816 (N_38816,N_37808,N_37953);
nand U38817 (N_38817,N_36407,N_36344);
or U38818 (N_38818,N_37454,N_36816);
nor U38819 (N_38819,N_37583,N_36857);
nand U38820 (N_38820,N_37978,N_37527);
xor U38821 (N_38821,N_36247,N_36226);
xor U38822 (N_38822,N_37672,N_36943);
nand U38823 (N_38823,N_37310,N_36004);
and U38824 (N_38824,N_36052,N_36776);
and U38825 (N_38825,N_36021,N_37741);
and U38826 (N_38826,N_36029,N_36713);
nor U38827 (N_38827,N_37043,N_36621);
nand U38828 (N_38828,N_37156,N_36616);
xnor U38829 (N_38829,N_36330,N_36204);
nor U38830 (N_38830,N_37579,N_37999);
nand U38831 (N_38831,N_37692,N_37241);
nor U38832 (N_38832,N_37140,N_37169);
nor U38833 (N_38833,N_36929,N_37930);
and U38834 (N_38834,N_36630,N_36754);
xor U38835 (N_38835,N_37355,N_37327);
xor U38836 (N_38836,N_37713,N_37611);
or U38837 (N_38837,N_36861,N_36348);
xor U38838 (N_38838,N_37306,N_37821);
or U38839 (N_38839,N_36289,N_37383);
nor U38840 (N_38840,N_36484,N_37220);
nand U38841 (N_38841,N_37475,N_36116);
nor U38842 (N_38842,N_36279,N_36098);
nand U38843 (N_38843,N_37100,N_36780);
xor U38844 (N_38844,N_37147,N_36183);
or U38845 (N_38845,N_36995,N_36211);
nand U38846 (N_38846,N_37659,N_37202);
and U38847 (N_38847,N_37796,N_37887);
or U38848 (N_38848,N_36854,N_36524);
and U38849 (N_38849,N_36801,N_37996);
or U38850 (N_38850,N_36377,N_37263);
nand U38851 (N_38851,N_36076,N_36297);
xnor U38852 (N_38852,N_36329,N_36189);
nor U38853 (N_38853,N_36668,N_36451);
nand U38854 (N_38854,N_37229,N_37638);
xnor U38855 (N_38855,N_37180,N_37640);
and U38856 (N_38856,N_37759,N_37522);
xnor U38857 (N_38857,N_36093,N_37095);
nand U38858 (N_38858,N_37621,N_36813);
xnor U38859 (N_38859,N_37338,N_36298);
xnor U38860 (N_38860,N_37063,N_36935);
xnor U38861 (N_38861,N_36221,N_36973);
nand U38862 (N_38862,N_36902,N_37949);
nand U38863 (N_38863,N_37440,N_37361);
or U38864 (N_38864,N_36845,N_36202);
and U38865 (N_38865,N_37036,N_36759);
nand U38866 (N_38866,N_37479,N_37077);
nor U38867 (N_38867,N_36733,N_36452);
nor U38868 (N_38868,N_37617,N_37493);
and U38869 (N_38869,N_36798,N_37099);
nor U38870 (N_38870,N_37577,N_37530);
or U38871 (N_38871,N_37160,N_37851);
and U38872 (N_38872,N_36919,N_37277);
xor U38873 (N_38873,N_37206,N_36554);
nor U38874 (N_38874,N_36694,N_36817);
xor U38875 (N_38875,N_37499,N_36794);
nand U38876 (N_38876,N_37835,N_37186);
and U38877 (N_38877,N_37258,N_37056);
nand U38878 (N_38878,N_36060,N_36632);
xor U38879 (N_38879,N_37680,N_37567);
xnor U38880 (N_38880,N_36040,N_36728);
nand U38881 (N_38881,N_37236,N_36235);
and U38882 (N_38882,N_37860,N_36931);
nor U38883 (N_38883,N_37717,N_36559);
nor U38884 (N_38884,N_37958,N_37888);
nand U38885 (N_38885,N_36151,N_36044);
or U38886 (N_38886,N_37182,N_36723);
xor U38887 (N_38887,N_36868,N_36031);
xor U38888 (N_38888,N_36633,N_37370);
nor U38889 (N_38889,N_36238,N_37971);
nor U38890 (N_38890,N_36530,N_37654);
xnor U38891 (N_38891,N_37494,N_36826);
xnor U38892 (N_38892,N_37682,N_36936);
xor U38893 (N_38893,N_37760,N_36212);
and U38894 (N_38894,N_37177,N_37685);
xnor U38895 (N_38895,N_37390,N_37406);
nor U38896 (N_38896,N_36472,N_37817);
or U38897 (N_38897,N_36002,N_37952);
or U38898 (N_38898,N_37447,N_37847);
nand U38899 (N_38899,N_36088,N_36879);
or U38900 (N_38900,N_36417,N_37329);
or U38901 (N_38901,N_37683,N_36895);
or U38902 (N_38902,N_37112,N_37666);
xor U38903 (N_38903,N_36851,N_37955);
or U38904 (N_38904,N_36579,N_37309);
or U38905 (N_38905,N_36431,N_36679);
nor U38906 (N_38906,N_36932,N_37927);
xnor U38907 (N_38907,N_36114,N_37096);
nand U38908 (N_38908,N_36981,N_36736);
nand U38909 (N_38909,N_36745,N_36287);
and U38910 (N_38910,N_36859,N_37079);
nand U38911 (N_38911,N_37340,N_36034);
xor U38912 (N_38912,N_36395,N_37854);
nor U38913 (N_38913,N_36145,N_36276);
xnor U38914 (N_38914,N_36371,N_36989);
xor U38915 (N_38915,N_37226,N_36529);
nor U38916 (N_38916,N_37515,N_37472);
nor U38917 (N_38917,N_36905,N_37951);
and U38918 (N_38918,N_36743,N_36280);
nor U38919 (N_38919,N_36079,N_37918);
xnor U38920 (N_38920,N_37892,N_36558);
or U38921 (N_38921,N_37873,N_36979);
nor U38922 (N_38922,N_37181,N_37480);
or U38923 (N_38923,N_37448,N_37913);
nand U38924 (N_38924,N_37465,N_37535);
and U38925 (N_38925,N_36106,N_37378);
or U38926 (N_38926,N_36394,N_37981);
nor U38927 (N_38927,N_36809,N_37405);
and U38928 (N_38928,N_36582,N_36094);
or U38929 (N_38929,N_36282,N_37473);
and U38930 (N_38930,N_37536,N_36576);
xnor U38931 (N_38931,N_37689,N_37570);
nor U38932 (N_38932,N_37740,N_37706);
or U38933 (N_38933,N_36257,N_37254);
nand U38934 (N_38934,N_36168,N_36292);
nand U38935 (N_38935,N_36405,N_36278);
or U38936 (N_38936,N_37352,N_36810);
nor U38937 (N_38937,N_36296,N_36656);
or U38938 (N_38938,N_37299,N_37539);
or U38939 (N_38939,N_36482,N_37786);
nor U38940 (N_38940,N_36426,N_36249);
nor U38941 (N_38941,N_36673,N_37588);
xor U38942 (N_38942,N_37076,N_37950);
nor U38943 (N_38943,N_37167,N_36241);
and U38944 (N_38944,N_37117,N_37374);
or U38945 (N_38945,N_36339,N_36546);
and U38946 (N_38946,N_37271,N_37752);
nand U38947 (N_38947,N_36806,N_36678);
nor U38948 (N_38948,N_36593,N_36655);
nor U38949 (N_38949,N_36313,N_37003);
xor U38950 (N_38950,N_37724,N_36644);
nor U38951 (N_38951,N_37396,N_36537);
or U38952 (N_38952,N_36309,N_36064);
nand U38953 (N_38953,N_36964,N_36054);
xor U38954 (N_38954,N_36381,N_36606);
xnor U38955 (N_38955,N_36572,N_36781);
and U38956 (N_38956,N_36356,N_36337);
xor U38957 (N_38957,N_36072,N_36602);
and U38958 (N_38958,N_37734,N_36814);
or U38959 (N_38959,N_36756,N_37013);
or U38960 (N_38960,N_37444,N_37252);
xor U38961 (N_38961,N_37173,N_37700);
nand U38962 (N_38962,N_37797,N_36453);
xnor U38963 (N_38963,N_36860,N_37867);
nand U38964 (N_38964,N_37497,N_36771);
and U38965 (N_38965,N_36148,N_37358);
nand U38966 (N_38966,N_37693,N_37985);
nor U38967 (N_38967,N_37135,N_36783);
xnor U38968 (N_38968,N_37624,N_36167);
xor U38969 (N_38969,N_36856,N_36275);
or U38970 (N_38970,N_37674,N_36444);
and U38971 (N_38971,N_37758,N_36786);
or U38972 (N_38972,N_37811,N_37089);
nand U38973 (N_38973,N_37763,N_36427);
xor U38974 (N_38974,N_36828,N_36840);
nor U38975 (N_38975,N_37875,N_36841);
nor U38976 (N_38976,N_36074,N_36984);
nand U38977 (N_38977,N_36991,N_37387);
nor U38978 (N_38978,N_36388,N_37453);
xor U38979 (N_38979,N_37701,N_36542);
xor U38980 (N_38980,N_37809,N_37923);
and U38981 (N_38981,N_37931,N_37905);
nand U38982 (N_38982,N_36000,N_36314);
or U38983 (N_38983,N_37401,N_37294);
nand U38984 (N_38984,N_37323,N_36059);
xnor U38985 (N_38985,N_37318,N_36689);
nand U38986 (N_38986,N_37718,N_37886);
nand U38987 (N_38987,N_36594,N_37414);
xor U38988 (N_38988,N_36843,N_37037);
nand U38989 (N_38989,N_36824,N_36185);
nand U38990 (N_38990,N_37098,N_37599);
nor U38991 (N_38991,N_36855,N_36438);
nand U38992 (N_38992,N_36471,N_36505);
nor U38993 (N_38993,N_37551,N_36889);
or U38994 (N_38994,N_37164,N_37834);
nor U38995 (N_38995,N_36566,N_36234);
and U38996 (N_38996,N_36663,N_37282);
and U38997 (N_38997,N_37871,N_36415);
or U38998 (N_38998,N_36439,N_37214);
or U38999 (N_38999,N_37944,N_37053);
xor U39000 (N_39000,N_36992,N_36351);
nor U39001 (N_39001,N_37862,N_36251);
xor U39002 (N_39002,N_37384,N_36318);
xor U39003 (N_39003,N_36358,N_36225);
xor U39004 (N_39004,N_36437,N_36539);
and U39005 (N_39005,N_36557,N_37733);
nor U39006 (N_39006,N_37569,N_36234);
or U39007 (N_39007,N_36795,N_37914);
nor U39008 (N_39008,N_37116,N_36352);
nor U39009 (N_39009,N_37534,N_37398);
and U39010 (N_39010,N_37500,N_37097);
or U39011 (N_39011,N_36725,N_36516);
nor U39012 (N_39012,N_36639,N_37695);
or U39013 (N_39013,N_37526,N_36121);
nor U39014 (N_39014,N_36684,N_37610);
nand U39015 (N_39015,N_37654,N_37125);
nor U39016 (N_39016,N_37747,N_37493);
nor U39017 (N_39017,N_37746,N_37577);
or U39018 (N_39018,N_37648,N_37974);
or U39019 (N_39019,N_36974,N_37635);
or U39020 (N_39020,N_36587,N_37604);
and U39021 (N_39021,N_36427,N_37363);
and U39022 (N_39022,N_36565,N_37312);
nor U39023 (N_39023,N_36107,N_37727);
nor U39024 (N_39024,N_36225,N_36600);
nor U39025 (N_39025,N_36428,N_36454);
nor U39026 (N_39026,N_37183,N_36452);
or U39027 (N_39027,N_36856,N_36418);
nor U39028 (N_39028,N_37096,N_36171);
nand U39029 (N_39029,N_37746,N_37819);
xnor U39030 (N_39030,N_37171,N_37718);
nor U39031 (N_39031,N_37482,N_37791);
nor U39032 (N_39032,N_37054,N_36179);
or U39033 (N_39033,N_37892,N_37275);
and U39034 (N_39034,N_36450,N_37337);
and U39035 (N_39035,N_37087,N_36950);
and U39036 (N_39036,N_37849,N_37217);
nor U39037 (N_39037,N_37379,N_37873);
nand U39038 (N_39038,N_37812,N_37490);
nand U39039 (N_39039,N_36769,N_36423);
nor U39040 (N_39040,N_37092,N_37575);
and U39041 (N_39041,N_36944,N_37042);
nand U39042 (N_39042,N_37058,N_36814);
xor U39043 (N_39043,N_37467,N_37516);
nor U39044 (N_39044,N_37923,N_37140);
and U39045 (N_39045,N_36324,N_37309);
xnor U39046 (N_39046,N_36613,N_36970);
and U39047 (N_39047,N_36302,N_37455);
and U39048 (N_39048,N_36561,N_37568);
nand U39049 (N_39049,N_36750,N_36579);
nor U39050 (N_39050,N_37100,N_36061);
nand U39051 (N_39051,N_36283,N_37419);
and U39052 (N_39052,N_36368,N_36601);
or U39053 (N_39053,N_37911,N_36234);
xnor U39054 (N_39054,N_36182,N_37745);
and U39055 (N_39055,N_36832,N_37657);
or U39056 (N_39056,N_37616,N_37508);
or U39057 (N_39057,N_36769,N_37952);
nor U39058 (N_39058,N_36404,N_37986);
nor U39059 (N_39059,N_37649,N_36070);
nand U39060 (N_39060,N_36499,N_36658);
nor U39061 (N_39061,N_36277,N_37655);
nand U39062 (N_39062,N_36599,N_37972);
nor U39063 (N_39063,N_37425,N_37286);
and U39064 (N_39064,N_37912,N_37496);
nand U39065 (N_39065,N_37392,N_36507);
nor U39066 (N_39066,N_37524,N_36867);
and U39067 (N_39067,N_37196,N_36100);
nor U39068 (N_39068,N_37161,N_37460);
and U39069 (N_39069,N_37155,N_36242);
nor U39070 (N_39070,N_36782,N_36934);
nor U39071 (N_39071,N_37073,N_37337);
nand U39072 (N_39072,N_36037,N_37090);
nand U39073 (N_39073,N_36864,N_36630);
nand U39074 (N_39074,N_36280,N_37922);
xnor U39075 (N_39075,N_37462,N_37309);
nand U39076 (N_39076,N_37264,N_36789);
or U39077 (N_39077,N_36756,N_36039);
and U39078 (N_39078,N_36976,N_37090);
nand U39079 (N_39079,N_36419,N_36957);
xnor U39080 (N_39080,N_37826,N_36565);
xnor U39081 (N_39081,N_36285,N_37612);
nand U39082 (N_39082,N_36970,N_36330);
nand U39083 (N_39083,N_36991,N_37863);
nand U39084 (N_39084,N_37377,N_36794);
or U39085 (N_39085,N_36584,N_36720);
and U39086 (N_39086,N_36388,N_36384);
nand U39087 (N_39087,N_37930,N_37755);
nor U39088 (N_39088,N_36144,N_37471);
nand U39089 (N_39089,N_36171,N_36473);
or U39090 (N_39090,N_37525,N_37038);
or U39091 (N_39091,N_36836,N_37119);
xor U39092 (N_39092,N_36771,N_37236);
nand U39093 (N_39093,N_37898,N_36146);
and U39094 (N_39094,N_37944,N_36265);
and U39095 (N_39095,N_37771,N_36531);
nor U39096 (N_39096,N_37567,N_36354);
or U39097 (N_39097,N_36209,N_37688);
xnor U39098 (N_39098,N_36618,N_36977);
and U39099 (N_39099,N_36099,N_36594);
xor U39100 (N_39100,N_36863,N_37920);
and U39101 (N_39101,N_36368,N_36738);
xnor U39102 (N_39102,N_36144,N_36985);
nor U39103 (N_39103,N_36175,N_37619);
or U39104 (N_39104,N_37733,N_37281);
nand U39105 (N_39105,N_36061,N_37099);
nor U39106 (N_39106,N_37078,N_37903);
nor U39107 (N_39107,N_37034,N_36050);
or U39108 (N_39108,N_37585,N_36572);
nor U39109 (N_39109,N_36385,N_36188);
nand U39110 (N_39110,N_36189,N_37768);
nand U39111 (N_39111,N_36355,N_36722);
xnor U39112 (N_39112,N_37115,N_37193);
nand U39113 (N_39113,N_36595,N_37198);
and U39114 (N_39114,N_36479,N_36917);
and U39115 (N_39115,N_36257,N_36627);
or U39116 (N_39116,N_36601,N_36086);
and U39117 (N_39117,N_37130,N_37802);
and U39118 (N_39118,N_37751,N_37154);
nor U39119 (N_39119,N_36664,N_36029);
and U39120 (N_39120,N_36747,N_36927);
nor U39121 (N_39121,N_37571,N_36414);
nand U39122 (N_39122,N_36914,N_36101);
nor U39123 (N_39123,N_37514,N_37293);
nor U39124 (N_39124,N_36607,N_37536);
xnor U39125 (N_39125,N_36959,N_37404);
or U39126 (N_39126,N_37541,N_36806);
nand U39127 (N_39127,N_37631,N_37350);
and U39128 (N_39128,N_36059,N_37436);
or U39129 (N_39129,N_36740,N_37682);
xor U39130 (N_39130,N_36257,N_36511);
nand U39131 (N_39131,N_37368,N_37058);
xor U39132 (N_39132,N_37231,N_36697);
or U39133 (N_39133,N_37956,N_37355);
xnor U39134 (N_39134,N_37304,N_36651);
or U39135 (N_39135,N_36009,N_36629);
and U39136 (N_39136,N_36182,N_37350);
and U39137 (N_39137,N_36777,N_37565);
xor U39138 (N_39138,N_37726,N_37602);
xor U39139 (N_39139,N_36784,N_37404);
or U39140 (N_39140,N_36743,N_37812);
nand U39141 (N_39141,N_37435,N_36332);
and U39142 (N_39142,N_36972,N_36466);
nor U39143 (N_39143,N_37149,N_37230);
nand U39144 (N_39144,N_37692,N_36430);
or U39145 (N_39145,N_36894,N_37641);
or U39146 (N_39146,N_36520,N_37913);
and U39147 (N_39147,N_36515,N_37798);
nand U39148 (N_39148,N_37806,N_37172);
or U39149 (N_39149,N_37645,N_37689);
nand U39150 (N_39150,N_37299,N_37003);
and U39151 (N_39151,N_37159,N_37390);
and U39152 (N_39152,N_37046,N_36643);
nand U39153 (N_39153,N_37138,N_37482);
and U39154 (N_39154,N_37156,N_36619);
or U39155 (N_39155,N_37447,N_36293);
or U39156 (N_39156,N_37387,N_36795);
and U39157 (N_39157,N_36649,N_36030);
xor U39158 (N_39158,N_37954,N_36931);
nor U39159 (N_39159,N_36051,N_36921);
and U39160 (N_39160,N_37673,N_37665);
or U39161 (N_39161,N_37518,N_36306);
or U39162 (N_39162,N_37262,N_37936);
and U39163 (N_39163,N_36422,N_36838);
or U39164 (N_39164,N_37460,N_36274);
and U39165 (N_39165,N_36546,N_36526);
nand U39166 (N_39166,N_37752,N_37158);
or U39167 (N_39167,N_36773,N_37761);
nor U39168 (N_39168,N_36914,N_36123);
and U39169 (N_39169,N_37079,N_36630);
nand U39170 (N_39170,N_36958,N_37369);
xor U39171 (N_39171,N_36826,N_37531);
xnor U39172 (N_39172,N_36034,N_37762);
or U39173 (N_39173,N_36316,N_37654);
nand U39174 (N_39174,N_37498,N_36432);
or U39175 (N_39175,N_37405,N_37198);
nand U39176 (N_39176,N_36929,N_36040);
or U39177 (N_39177,N_36520,N_37349);
or U39178 (N_39178,N_37915,N_36769);
nor U39179 (N_39179,N_36562,N_37615);
and U39180 (N_39180,N_36255,N_36741);
nand U39181 (N_39181,N_36615,N_36948);
or U39182 (N_39182,N_36294,N_36638);
nor U39183 (N_39183,N_37264,N_37806);
nor U39184 (N_39184,N_36322,N_37935);
nand U39185 (N_39185,N_36022,N_36952);
nand U39186 (N_39186,N_36320,N_36823);
xor U39187 (N_39187,N_37063,N_36732);
and U39188 (N_39188,N_37752,N_36475);
nor U39189 (N_39189,N_36724,N_36554);
nand U39190 (N_39190,N_37737,N_37133);
nor U39191 (N_39191,N_36500,N_36975);
and U39192 (N_39192,N_37753,N_37646);
or U39193 (N_39193,N_37358,N_36366);
xnor U39194 (N_39194,N_37827,N_37651);
or U39195 (N_39195,N_37606,N_36762);
xor U39196 (N_39196,N_37253,N_36933);
xnor U39197 (N_39197,N_37465,N_36924);
xor U39198 (N_39198,N_36332,N_36182);
or U39199 (N_39199,N_36867,N_36885);
or U39200 (N_39200,N_36230,N_36921);
or U39201 (N_39201,N_36595,N_37583);
nand U39202 (N_39202,N_36208,N_37369);
xor U39203 (N_39203,N_36511,N_36108);
xnor U39204 (N_39204,N_36616,N_37124);
or U39205 (N_39205,N_37868,N_37213);
nor U39206 (N_39206,N_37105,N_37036);
xnor U39207 (N_39207,N_37055,N_36909);
and U39208 (N_39208,N_36778,N_36383);
nor U39209 (N_39209,N_37756,N_36809);
xor U39210 (N_39210,N_37748,N_36026);
and U39211 (N_39211,N_37807,N_37059);
or U39212 (N_39212,N_36252,N_36584);
or U39213 (N_39213,N_37919,N_36268);
and U39214 (N_39214,N_36326,N_36069);
or U39215 (N_39215,N_37779,N_37949);
xnor U39216 (N_39216,N_37228,N_36990);
nand U39217 (N_39217,N_37528,N_36204);
xnor U39218 (N_39218,N_36695,N_36464);
and U39219 (N_39219,N_37684,N_37710);
nor U39220 (N_39220,N_37614,N_36196);
and U39221 (N_39221,N_37439,N_37740);
nand U39222 (N_39222,N_36928,N_36539);
xnor U39223 (N_39223,N_36487,N_37072);
nor U39224 (N_39224,N_36967,N_36313);
nor U39225 (N_39225,N_36166,N_36078);
nand U39226 (N_39226,N_37068,N_37473);
nand U39227 (N_39227,N_37105,N_36206);
nand U39228 (N_39228,N_37132,N_36175);
xnor U39229 (N_39229,N_37671,N_36537);
or U39230 (N_39230,N_37709,N_36295);
or U39231 (N_39231,N_36920,N_37187);
nor U39232 (N_39232,N_36539,N_36865);
xor U39233 (N_39233,N_36343,N_36622);
xor U39234 (N_39234,N_37909,N_36002);
and U39235 (N_39235,N_36897,N_37583);
nand U39236 (N_39236,N_36977,N_36240);
and U39237 (N_39237,N_37144,N_36827);
or U39238 (N_39238,N_37933,N_36185);
or U39239 (N_39239,N_36246,N_36610);
or U39240 (N_39240,N_36944,N_36097);
xor U39241 (N_39241,N_37343,N_37338);
and U39242 (N_39242,N_37719,N_37866);
xor U39243 (N_39243,N_36216,N_36928);
xor U39244 (N_39244,N_37470,N_36047);
xor U39245 (N_39245,N_36450,N_36120);
nand U39246 (N_39246,N_37318,N_37976);
or U39247 (N_39247,N_37928,N_36386);
nor U39248 (N_39248,N_37613,N_37779);
nand U39249 (N_39249,N_36357,N_37941);
nor U39250 (N_39250,N_36400,N_36695);
xor U39251 (N_39251,N_37434,N_36704);
or U39252 (N_39252,N_37527,N_36588);
and U39253 (N_39253,N_36715,N_37256);
nand U39254 (N_39254,N_36875,N_36034);
or U39255 (N_39255,N_37779,N_36103);
and U39256 (N_39256,N_37387,N_37418);
or U39257 (N_39257,N_36361,N_37361);
or U39258 (N_39258,N_36681,N_37431);
xor U39259 (N_39259,N_36739,N_36948);
or U39260 (N_39260,N_37289,N_37207);
xor U39261 (N_39261,N_36199,N_37163);
and U39262 (N_39262,N_36381,N_36976);
xor U39263 (N_39263,N_37248,N_36369);
or U39264 (N_39264,N_36733,N_37738);
and U39265 (N_39265,N_36931,N_37737);
nor U39266 (N_39266,N_36585,N_37585);
and U39267 (N_39267,N_36749,N_36527);
or U39268 (N_39268,N_36709,N_37236);
nor U39269 (N_39269,N_36063,N_36605);
xor U39270 (N_39270,N_36126,N_37221);
xnor U39271 (N_39271,N_37583,N_36416);
nand U39272 (N_39272,N_37298,N_36630);
or U39273 (N_39273,N_36988,N_36686);
nand U39274 (N_39274,N_37115,N_36448);
or U39275 (N_39275,N_37125,N_36918);
and U39276 (N_39276,N_36728,N_37524);
nor U39277 (N_39277,N_37139,N_37062);
nand U39278 (N_39278,N_36963,N_36407);
and U39279 (N_39279,N_36741,N_37272);
xor U39280 (N_39280,N_36356,N_36898);
xor U39281 (N_39281,N_37797,N_36253);
nor U39282 (N_39282,N_36370,N_36000);
nand U39283 (N_39283,N_36053,N_36789);
or U39284 (N_39284,N_37801,N_37633);
nor U39285 (N_39285,N_37728,N_36093);
or U39286 (N_39286,N_37037,N_37381);
and U39287 (N_39287,N_37553,N_36711);
nand U39288 (N_39288,N_37641,N_37295);
nor U39289 (N_39289,N_36501,N_36555);
xnor U39290 (N_39290,N_37230,N_37647);
nor U39291 (N_39291,N_37595,N_36690);
nand U39292 (N_39292,N_37236,N_37947);
and U39293 (N_39293,N_37525,N_36853);
nor U39294 (N_39294,N_36210,N_37831);
nand U39295 (N_39295,N_36148,N_37211);
or U39296 (N_39296,N_36622,N_36833);
or U39297 (N_39297,N_36898,N_36908);
and U39298 (N_39298,N_36380,N_37489);
or U39299 (N_39299,N_36996,N_36900);
nor U39300 (N_39300,N_37108,N_36227);
nand U39301 (N_39301,N_37956,N_37551);
nor U39302 (N_39302,N_37699,N_37394);
or U39303 (N_39303,N_37494,N_36147);
xnor U39304 (N_39304,N_37819,N_36819);
and U39305 (N_39305,N_37822,N_37369);
nand U39306 (N_39306,N_36375,N_37745);
nor U39307 (N_39307,N_37199,N_37553);
nor U39308 (N_39308,N_36094,N_36996);
xnor U39309 (N_39309,N_37853,N_37526);
and U39310 (N_39310,N_36453,N_37066);
nor U39311 (N_39311,N_37686,N_36257);
xor U39312 (N_39312,N_37869,N_37612);
nor U39313 (N_39313,N_37517,N_36835);
nand U39314 (N_39314,N_37980,N_36652);
xor U39315 (N_39315,N_36271,N_36474);
or U39316 (N_39316,N_37897,N_37435);
or U39317 (N_39317,N_36032,N_36883);
nor U39318 (N_39318,N_36982,N_36334);
or U39319 (N_39319,N_36170,N_36868);
nor U39320 (N_39320,N_37535,N_37499);
nor U39321 (N_39321,N_37728,N_37814);
xor U39322 (N_39322,N_37125,N_37021);
nand U39323 (N_39323,N_37760,N_37400);
or U39324 (N_39324,N_37688,N_36292);
or U39325 (N_39325,N_36493,N_36153);
nor U39326 (N_39326,N_37077,N_36873);
and U39327 (N_39327,N_37401,N_36153);
or U39328 (N_39328,N_36345,N_37231);
or U39329 (N_39329,N_37922,N_36815);
or U39330 (N_39330,N_37302,N_36890);
xnor U39331 (N_39331,N_36398,N_36638);
nand U39332 (N_39332,N_37623,N_36067);
nor U39333 (N_39333,N_36541,N_36533);
nor U39334 (N_39334,N_36001,N_36643);
nor U39335 (N_39335,N_36384,N_36806);
and U39336 (N_39336,N_37456,N_36995);
nand U39337 (N_39337,N_37482,N_37818);
xnor U39338 (N_39338,N_37500,N_37017);
or U39339 (N_39339,N_36474,N_37597);
nor U39340 (N_39340,N_36795,N_36213);
or U39341 (N_39341,N_37122,N_37063);
xnor U39342 (N_39342,N_37372,N_36120);
or U39343 (N_39343,N_37203,N_36027);
or U39344 (N_39344,N_36447,N_37598);
or U39345 (N_39345,N_37959,N_37302);
nand U39346 (N_39346,N_37302,N_36883);
or U39347 (N_39347,N_36645,N_36253);
xor U39348 (N_39348,N_36405,N_37674);
and U39349 (N_39349,N_36687,N_37442);
xor U39350 (N_39350,N_36481,N_36515);
xor U39351 (N_39351,N_37416,N_36125);
nor U39352 (N_39352,N_36626,N_36144);
xnor U39353 (N_39353,N_36075,N_36468);
or U39354 (N_39354,N_37658,N_36711);
nand U39355 (N_39355,N_37256,N_37452);
and U39356 (N_39356,N_36603,N_37236);
nor U39357 (N_39357,N_37330,N_36276);
and U39358 (N_39358,N_36867,N_36650);
nand U39359 (N_39359,N_36301,N_36453);
nand U39360 (N_39360,N_36553,N_37727);
or U39361 (N_39361,N_36512,N_37350);
or U39362 (N_39362,N_37957,N_36920);
nor U39363 (N_39363,N_36504,N_36670);
nor U39364 (N_39364,N_37927,N_36626);
or U39365 (N_39365,N_36783,N_36134);
nor U39366 (N_39366,N_37971,N_37617);
nand U39367 (N_39367,N_36016,N_36751);
nor U39368 (N_39368,N_37281,N_37337);
nand U39369 (N_39369,N_36256,N_36264);
or U39370 (N_39370,N_36271,N_37526);
nand U39371 (N_39371,N_36714,N_37979);
nor U39372 (N_39372,N_36601,N_36732);
nand U39373 (N_39373,N_37424,N_37873);
xnor U39374 (N_39374,N_37563,N_36515);
or U39375 (N_39375,N_36820,N_37118);
nand U39376 (N_39376,N_37020,N_36660);
nand U39377 (N_39377,N_36908,N_36414);
xor U39378 (N_39378,N_37107,N_36445);
or U39379 (N_39379,N_36053,N_37734);
nor U39380 (N_39380,N_37580,N_37323);
nor U39381 (N_39381,N_36758,N_36845);
xor U39382 (N_39382,N_36939,N_36322);
nand U39383 (N_39383,N_36568,N_37054);
or U39384 (N_39384,N_36724,N_37048);
or U39385 (N_39385,N_37299,N_37577);
nand U39386 (N_39386,N_36224,N_36115);
or U39387 (N_39387,N_36269,N_36077);
and U39388 (N_39388,N_36598,N_36421);
xnor U39389 (N_39389,N_36801,N_37623);
nand U39390 (N_39390,N_37579,N_36289);
or U39391 (N_39391,N_37088,N_36145);
nor U39392 (N_39392,N_36938,N_36072);
xor U39393 (N_39393,N_37643,N_37499);
xor U39394 (N_39394,N_37535,N_37076);
xor U39395 (N_39395,N_37607,N_37151);
nor U39396 (N_39396,N_36021,N_37211);
and U39397 (N_39397,N_37187,N_37508);
and U39398 (N_39398,N_37079,N_37199);
and U39399 (N_39399,N_37957,N_37664);
and U39400 (N_39400,N_36398,N_36890);
nand U39401 (N_39401,N_36290,N_36414);
and U39402 (N_39402,N_36363,N_36102);
nor U39403 (N_39403,N_36920,N_37136);
or U39404 (N_39404,N_36497,N_37977);
or U39405 (N_39405,N_36022,N_36230);
nand U39406 (N_39406,N_36136,N_36915);
xnor U39407 (N_39407,N_37837,N_37650);
nand U39408 (N_39408,N_36783,N_36922);
and U39409 (N_39409,N_36668,N_36093);
xor U39410 (N_39410,N_36681,N_36666);
xor U39411 (N_39411,N_36943,N_36799);
nand U39412 (N_39412,N_37330,N_36901);
nand U39413 (N_39413,N_36116,N_37944);
nand U39414 (N_39414,N_36041,N_36446);
and U39415 (N_39415,N_36381,N_36942);
or U39416 (N_39416,N_36994,N_36591);
or U39417 (N_39417,N_36988,N_37125);
and U39418 (N_39418,N_37203,N_37831);
and U39419 (N_39419,N_36003,N_37880);
or U39420 (N_39420,N_36876,N_36312);
nand U39421 (N_39421,N_37228,N_36134);
nor U39422 (N_39422,N_37129,N_36233);
nand U39423 (N_39423,N_37724,N_36105);
nor U39424 (N_39424,N_37851,N_36432);
nand U39425 (N_39425,N_36398,N_36718);
and U39426 (N_39426,N_36576,N_37946);
nor U39427 (N_39427,N_36381,N_37092);
nor U39428 (N_39428,N_37940,N_37492);
and U39429 (N_39429,N_36541,N_37359);
nand U39430 (N_39430,N_36291,N_36790);
xnor U39431 (N_39431,N_37341,N_36118);
and U39432 (N_39432,N_37836,N_36697);
and U39433 (N_39433,N_37591,N_37224);
nand U39434 (N_39434,N_37999,N_37881);
or U39435 (N_39435,N_36617,N_36249);
or U39436 (N_39436,N_36365,N_36513);
nor U39437 (N_39437,N_37426,N_36475);
or U39438 (N_39438,N_37761,N_37435);
xnor U39439 (N_39439,N_37595,N_36221);
nand U39440 (N_39440,N_36527,N_37455);
or U39441 (N_39441,N_36767,N_37050);
xor U39442 (N_39442,N_37445,N_36026);
and U39443 (N_39443,N_37261,N_37568);
nand U39444 (N_39444,N_37020,N_37179);
nor U39445 (N_39445,N_36981,N_36733);
nor U39446 (N_39446,N_37095,N_37900);
xor U39447 (N_39447,N_37620,N_36540);
nand U39448 (N_39448,N_37199,N_36031);
or U39449 (N_39449,N_36267,N_36350);
or U39450 (N_39450,N_36116,N_36242);
xor U39451 (N_39451,N_36016,N_36384);
nor U39452 (N_39452,N_37940,N_37194);
xor U39453 (N_39453,N_37713,N_37965);
nor U39454 (N_39454,N_37746,N_37180);
nand U39455 (N_39455,N_37182,N_36396);
nand U39456 (N_39456,N_36818,N_36513);
xnor U39457 (N_39457,N_36711,N_36627);
nand U39458 (N_39458,N_36894,N_36994);
or U39459 (N_39459,N_37527,N_37163);
nor U39460 (N_39460,N_36720,N_36016);
or U39461 (N_39461,N_36630,N_37627);
nand U39462 (N_39462,N_36253,N_37050);
or U39463 (N_39463,N_36791,N_37197);
xor U39464 (N_39464,N_36304,N_37984);
nor U39465 (N_39465,N_36710,N_37377);
and U39466 (N_39466,N_37418,N_37488);
nand U39467 (N_39467,N_36465,N_36462);
xor U39468 (N_39468,N_37514,N_36414);
or U39469 (N_39469,N_37864,N_37571);
nand U39470 (N_39470,N_36877,N_36994);
nand U39471 (N_39471,N_36042,N_36429);
or U39472 (N_39472,N_36338,N_37995);
or U39473 (N_39473,N_36369,N_36415);
or U39474 (N_39474,N_36430,N_37580);
or U39475 (N_39475,N_36905,N_37146);
and U39476 (N_39476,N_36206,N_36082);
nor U39477 (N_39477,N_36462,N_36480);
xnor U39478 (N_39478,N_36192,N_36430);
or U39479 (N_39479,N_36981,N_36099);
and U39480 (N_39480,N_37212,N_37957);
nand U39481 (N_39481,N_36744,N_36366);
xor U39482 (N_39482,N_36847,N_36091);
or U39483 (N_39483,N_36504,N_36756);
nor U39484 (N_39484,N_36610,N_36411);
xnor U39485 (N_39485,N_37578,N_36415);
and U39486 (N_39486,N_36190,N_36294);
and U39487 (N_39487,N_36563,N_36153);
and U39488 (N_39488,N_37580,N_36569);
and U39489 (N_39489,N_37773,N_37758);
and U39490 (N_39490,N_37976,N_36335);
or U39491 (N_39491,N_36452,N_36289);
nand U39492 (N_39492,N_36976,N_36592);
nor U39493 (N_39493,N_36549,N_37993);
and U39494 (N_39494,N_37007,N_37605);
or U39495 (N_39495,N_36513,N_37456);
xnor U39496 (N_39496,N_36871,N_37928);
nand U39497 (N_39497,N_37263,N_36811);
or U39498 (N_39498,N_37062,N_36726);
nor U39499 (N_39499,N_37322,N_36140);
nor U39500 (N_39500,N_36707,N_36697);
nor U39501 (N_39501,N_36350,N_36452);
and U39502 (N_39502,N_36542,N_37128);
nand U39503 (N_39503,N_37193,N_36885);
nor U39504 (N_39504,N_37497,N_36919);
and U39505 (N_39505,N_36023,N_36412);
nand U39506 (N_39506,N_36291,N_37762);
xnor U39507 (N_39507,N_37814,N_37481);
nor U39508 (N_39508,N_36729,N_37769);
and U39509 (N_39509,N_37281,N_36015);
xor U39510 (N_39510,N_36365,N_37150);
xnor U39511 (N_39511,N_36520,N_36037);
or U39512 (N_39512,N_37728,N_37118);
and U39513 (N_39513,N_37484,N_37628);
nor U39514 (N_39514,N_36560,N_36970);
and U39515 (N_39515,N_37121,N_37552);
and U39516 (N_39516,N_36256,N_36535);
xor U39517 (N_39517,N_37308,N_36310);
or U39518 (N_39518,N_36895,N_37249);
and U39519 (N_39519,N_37980,N_37703);
nor U39520 (N_39520,N_36695,N_37125);
or U39521 (N_39521,N_37271,N_37896);
xor U39522 (N_39522,N_37395,N_36040);
xnor U39523 (N_39523,N_37550,N_37523);
or U39524 (N_39524,N_36991,N_36809);
nor U39525 (N_39525,N_37965,N_37871);
xnor U39526 (N_39526,N_37872,N_37613);
or U39527 (N_39527,N_36465,N_36484);
or U39528 (N_39528,N_37931,N_36366);
and U39529 (N_39529,N_37719,N_37072);
nor U39530 (N_39530,N_37559,N_36631);
xor U39531 (N_39531,N_37005,N_36428);
xor U39532 (N_39532,N_36196,N_36173);
nor U39533 (N_39533,N_37340,N_37521);
xnor U39534 (N_39534,N_37837,N_36611);
nand U39535 (N_39535,N_37298,N_37014);
nor U39536 (N_39536,N_37331,N_37943);
nand U39537 (N_39537,N_37089,N_37915);
and U39538 (N_39538,N_37536,N_36433);
xnor U39539 (N_39539,N_37494,N_37374);
xor U39540 (N_39540,N_36827,N_37677);
and U39541 (N_39541,N_37337,N_36070);
xor U39542 (N_39542,N_37220,N_37655);
and U39543 (N_39543,N_37023,N_36897);
xor U39544 (N_39544,N_36714,N_36790);
and U39545 (N_39545,N_36475,N_37891);
nor U39546 (N_39546,N_37221,N_36166);
nor U39547 (N_39547,N_36585,N_36503);
and U39548 (N_39548,N_36741,N_36856);
and U39549 (N_39549,N_36574,N_36349);
xnor U39550 (N_39550,N_37892,N_36040);
nor U39551 (N_39551,N_36711,N_36607);
xnor U39552 (N_39552,N_36065,N_36249);
and U39553 (N_39553,N_37011,N_36152);
or U39554 (N_39554,N_37158,N_37804);
or U39555 (N_39555,N_36090,N_37704);
xnor U39556 (N_39556,N_36985,N_37598);
xor U39557 (N_39557,N_37613,N_37931);
or U39558 (N_39558,N_36662,N_37925);
nor U39559 (N_39559,N_37615,N_37328);
and U39560 (N_39560,N_36694,N_37749);
nand U39561 (N_39561,N_37493,N_37082);
nand U39562 (N_39562,N_37887,N_37693);
or U39563 (N_39563,N_37711,N_37660);
and U39564 (N_39564,N_36449,N_36804);
xor U39565 (N_39565,N_37310,N_36598);
and U39566 (N_39566,N_36570,N_36248);
nor U39567 (N_39567,N_36053,N_37252);
or U39568 (N_39568,N_36405,N_37451);
or U39569 (N_39569,N_36762,N_37798);
nor U39570 (N_39570,N_36102,N_37251);
and U39571 (N_39571,N_37233,N_37424);
nor U39572 (N_39572,N_36140,N_36359);
or U39573 (N_39573,N_36566,N_37843);
xnor U39574 (N_39574,N_36029,N_36829);
and U39575 (N_39575,N_36607,N_37730);
nor U39576 (N_39576,N_37726,N_36403);
or U39577 (N_39577,N_37746,N_37890);
or U39578 (N_39578,N_37929,N_37389);
nand U39579 (N_39579,N_36683,N_37460);
nor U39580 (N_39580,N_36801,N_37715);
and U39581 (N_39581,N_36609,N_36521);
nor U39582 (N_39582,N_36683,N_37571);
xor U39583 (N_39583,N_37440,N_36971);
nand U39584 (N_39584,N_36043,N_36181);
nor U39585 (N_39585,N_37452,N_36028);
nand U39586 (N_39586,N_36236,N_37213);
xor U39587 (N_39587,N_37300,N_36468);
or U39588 (N_39588,N_37060,N_37200);
nand U39589 (N_39589,N_36452,N_37697);
nor U39590 (N_39590,N_36396,N_37254);
or U39591 (N_39591,N_37067,N_36362);
xor U39592 (N_39592,N_36669,N_37051);
xnor U39593 (N_39593,N_37624,N_37763);
or U39594 (N_39594,N_37404,N_37808);
or U39595 (N_39595,N_36937,N_36110);
nand U39596 (N_39596,N_37731,N_37101);
nand U39597 (N_39597,N_36513,N_37084);
and U39598 (N_39598,N_36162,N_37479);
xor U39599 (N_39599,N_36980,N_37052);
nor U39600 (N_39600,N_36435,N_37502);
nor U39601 (N_39601,N_36065,N_37445);
and U39602 (N_39602,N_36148,N_37525);
and U39603 (N_39603,N_37731,N_37096);
xnor U39604 (N_39604,N_37479,N_37093);
or U39605 (N_39605,N_37356,N_36489);
nand U39606 (N_39606,N_36775,N_37986);
xnor U39607 (N_39607,N_36528,N_37848);
and U39608 (N_39608,N_36352,N_36013);
nand U39609 (N_39609,N_37327,N_36869);
nand U39610 (N_39610,N_36094,N_36879);
xor U39611 (N_39611,N_37319,N_37372);
nand U39612 (N_39612,N_37034,N_36489);
nor U39613 (N_39613,N_36380,N_37183);
xor U39614 (N_39614,N_37432,N_36426);
nand U39615 (N_39615,N_36486,N_36891);
xor U39616 (N_39616,N_36654,N_36507);
xnor U39617 (N_39617,N_37130,N_36943);
xnor U39618 (N_39618,N_36574,N_37038);
or U39619 (N_39619,N_36924,N_36595);
nand U39620 (N_39620,N_36555,N_37465);
xor U39621 (N_39621,N_36071,N_36626);
and U39622 (N_39622,N_36617,N_36800);
xor U39623 (N_39623,N_37962,N_36633);
or U39624 (N_39624,N_36597,N_36739);
nor U39625 (N_39625,N_36344,N_37614);
nor U39626 (N_39626,N_37911,N_37863);
nand U39627 (N_39627,N_36474,N_36629);
nand U39628 (N_39628,N_37122,N_36886);
nor U39629 (N_39629,N_36108,N_36700);
and U39630 (N_39630,N_36900,N_36224);
or U39631 (N_39631,N_37256,N_37804);
nor U39632 (N_39632,N_37041,N_37939);
xor U39633 (N_39633,N_36083,N_37696);
nand U39634 (N_39634,N_37259,N_37103);
nor U39635 (N_39635,N_36770,N_36415);
xnor U39636 (N_39636,N_36110,N_36966);
nor U39637 (N_39637,N_36321,N_36822);
nor U39638 (N_39638,N_37831,N_36987);
nand U39639 (N_39639,N_36006,N_37473);
nand U39640 (N_39640,N_37966,N_36944);
nor U39641 (N_39641,N_36848,N_36708);
and U39642 (N_39642,N_37737,N_37021);
xnor U39643 (N_39643,N_36302,N_36781);
nor U39644 (N_39644,N_36948,N_36765);
xnor U39645 (N_39645,N_36658,N_36296);
and U39646 (N_39646,N_37754,N_37327);
or U39647 (N_39647,N_36522,N_37498);
nor U39648 (N_39648,N_36750,N_36543);
nor U39649 (N_39649,N_36816,N_37272);
xnor U39650 (N_39650,N_36447,N_36692);
and U39651 (N_39651,N_36543,N_37190);
xor U39652 (N_39652,N_37844,N_36251);
nand U39653 (N_39653,N_36953,N_36434);
or U39654 (N_39654,N_37344,N_37870);
xnor U39655 (N_39655,N_36161,N_36242);
or U39656 (N_39656,N_36066,N_37234);
or U39657 (N_39657,N_36998,N_37812);
nand U39658 (N_39658,N_37467,N_36186);
and U39659 (N_39659,N_37108,N_37568);
or U39660 (N_39660,N_37075,N_37593);
or U39661 (N_39661,N_36422,N_37353);
and U39662 (N_39662,N_37581,N_37997);
nor U39663 (N_39663,N_37763,N_36717);
and U39664 (N_39664,N_37089,N_37504);
or U39665 (N_39665,N_36798,N_37873);
and U39666 (N_39666,N_37879,N_36527);
and U39667 (N_39667,N_36815,N_36704);
xnor U39668 (N_39668,N_37409,N_36518);
xnor U39669 (N_39669,N_36091,N_36467);
or U39670 (N_39670,N_36706,N_37245);
nand U39671 (N_39671,N_36089,N_37452);
and U39672 (N_39672,N_36949,N_37720);
or U39673 (N_39673,N_36629,N_37717);
xor U39674 (N_39674,N_37628,N_36838);
nand U39675 (N_39675,N_36494,N_36300);
xnor U39676 (N_39676,N_37754,N_36395);
nor U39677 (N_39677,N_36906,N_37104);
xnor U39678 (N_39678,N_37193,N_36632);
nor U39679 (N_39679,N_37178,N_37851);
and U39680 (N_39680,N_36829,N_36307);
xor U39681 (N_39681,N_37933,N_36826);
or U39682 (N_39682,N_36996,N_36139);
and U39683 (N_39683,N_36699,N_36614);
nor U39684 (N_39684,N_37050,N_36270);
or U39685 (N_39685,N_37571,N_37965);
nor U39686 (N_39686,N_37931,N_37658);
or U39687 (N_39687,N_36034,N_36303);
nor U39688 (N_39688,N_36907,N_37587);
and U39689 (N_39689,N_37642,N_37323);
or U39690 (N_39690,N_36633,N_36392);
or U39691 (N_39691,N_37422,N_37898);
nor U39692 (N_39692,N_37083,N_36970);
or U39693 (N_39693,N_36572,N_36934);
or U39694 (N_39694,N_36633,N_37600);
xor U39695 (N_39695,N_37707,N_37075);
and U39696 (N_39696,N_36789,N_37208);
nor U39697 (N_39697,N_37559,N_36132);
nand U39698 (N_39698,N_37939,N_36192);
or U39699 (N_39699,N_36042,N_36734);
nand U39700 (N_39700,N_36436,N_36690);
nor U39701 (N_39701,N_36680,N_37435);
and U39702 (N_39702,N_36075,N_37424);
or U39703 (N_39703,N_37568,N_37901);
xor U39704 (N_39704,N_36840,N_36566);
nand U39705 (N_39705,N_37804,N_37314);
nand U39706 (N_39706,N_36349,N_37655);
nor U39707 (N_39707,N_37290,N_36735);
nand U39708 (N_39708,N_37034,N_37767);
nor U39709 (N_39709,N_36725,N_36198);
nand U39710 (N_39710,N_36895,N_36653);
xnor U39711 (N_39711,N_37549,N_37788);
nor U39712 (N_39712,N_37864,N_36164);
or U39713 (N_39713,N_36376,N_36514);
or U39714 (N_39714,N_36581,N_36272);
and U39715 (N_39715,N_37542,N_36957);
nand U39716 (N_39716,N_36520,N_37099);
nor U39717 (N_39717,N_36763,N_37541);
nor U39718 (N_39718,N_37147,N_37938);
or U39719 (N_39719,N_37387,N_37500);
xor U39720 (N_39720,N_37364,N_36551);
or U39721 (N_39721,N_36655,N_36797);
nand U39722 (N_39722,N_36414,N_36807);
xnor U39723 (N_39723,N_36782,N_36794);
nor U39724 (N_39724,N_37207,N_37673);
xnor U39725 (N_39725,N_37873,N_37008);
or U39726 (N_39726,N_37153,N_36603);
xnor U39727 (N_39727,N_36972,N_37628);
and U39728 (N_39728,N_37880,N_36902);
xor U39729 (N_39729,N_37738,N_37508);
xnor U39730 (N_39730,N_37970,N_37901);
nand U39731 (N_39731,N_37645,N_37063);
and U39732 (N_39732,N_36668,N_36810);
nand U39733 (N_39733,N_37728,N_37850);
and U39734 (N_39734,N_37190,N_37296);
xor U39735 (N_39735,N_36949,N_37499);
or U39736 (N_39736,N_36428,N_36726);
nor U39737 (N_39737,N_37543,N_36898);
nor U39738 (N_39738,N_36950,N_37683);
and U39739 (N_39739,N_37541,N_36756);
nor U39740 (N_39740,N_37807,N_37569);
nand U39741 (N_39741,N_37088,N_36502);
nor U39742 (N_39742,N_37767,N_37306);
or U39743 (N_39743,N_37646,N_37020);
nor U39744 (N_39744,N_37847,N_37007);
nor U39745 (N_39745,N_36976,N_36788);
xnor U39746 (N_39746,N_37405,N_36962);
or U39747 (N_39747,N_37347,N_37965);
nand U39748 (N_39748,N_37829,N_37217);
or U39749 (N_39749,N_37799,N_36025);
and U39750 (N_39750,N_36125,N_36472);
nor U39751 (N_39751,N_36585,N_37382);
nand U39752 (N_39752,N_37882,N_37905);
and U39753 (N_39753,N_37242,N_36134);
nand U39754 (N_39754,N_36603,N_36822);
or U39755 (N_39755,N_37938,N_37055);
nor U39756 (N_39756,N_37561,N_37871);
nand U39757 (N_39757,N_37045,N_37835);
and U39758 (N_39758,N_37261,N_37306);
nor U39759 (N_39759,N_36069,N_36663);
and U39760 (N_39760,N_37148,N_36219);
xnor U39761 (N_39761,N_36477,N_37363);
nor U39762 (N_39762,N_36913,N_37197);
nor U39763 (N_39763,N_37586,N_36666);
nand U39764 (N_39764,N_36256,N_37213);
nand U39765 (N_39765,N_37266,N_36399);
xnor U39766 (N_39766,N_36073,N_36717);
and U39767 (N_39767,N_36731,N_36192);
and U39768 (N_39768,N_37350,N_37859);
xnor U39769 (N_39769,N_36978,N_36479);
nor U39770 (N_39770,N_37157,N_37138);
and U39771 (N_39771,N_37218,N_37930);
and U39772 (N_39772,N_37453,N_36046);
and U39773 (N_39773,N_36572,N_36048);
nand U39774 (N_39774,N_37847,N_37126);
nand U39775 (N_39775,N_37642,N_36022);
or U39776 (N_39776,N_36401,N_36468);
and U39777 (N_39777,N_36554,N_37631);
and U39778 (N_39778,N_37856,N_37711);
and U39779 (N_39779,N_37034,N_37662);
and U39780 (N_39780,N_37198,N_37010);
and U39781 (N_39781,N_36143,N_36875);
xor U39782 (N_39782,N_36129,N_37708);
and U39783 (N_39783,N_37020,N_36603);
and U39784 (N_39784,N_37006,N_36156);
xor U39785 (N_39785,N_37230,N_36497);
nor U39786 (N_39786,N_37765,N_36438);
nand U39787 (N_39787,N_37458,N_37659);
nand U39788 (N_39788,N_37705,N_36609);
nand U39789 (N_39789,N_36469,N_36040);
nor U39790 (N_39790,N_36803,N_37467);
nand U39791 (N_39791,N_37189,N_36352);
nand U39792 (N_39792,N_37785,N_36157);
xor U39793 (N_39793,N_36305,N_36469);
and U39794 (N_39794,N_36534,N_36865);
and U39795 (N_39795,N_36032,N_36659);
or U39796 (N_39796,N_36204,N_37773);
nand U39797 (N_39797,N_37815,N_37772);
or U39798 (N_39798,N_37473,N_37804);
and U39799 (N_39799,N_36046,N_36047);
nor U39800 (N_39800,N_36921,N_36915);
and U39801 (N_39801,N_36360,N_36537);
nor U39802 (N_39802,N_37952,N_36718);
or U39803 (N_39803,N_37445,N_36737);
and U39804 (N_39804,N_37663,N_37617);
xnor U39805 (N_39805,N_37544,N_36970);
or U39806 (N_39806,N_37817,N_37411);
xor U39807 (N_39807,N_36157,N_37796);
nor U39808 (N_39808,N_37410,N_37664);
and U39809 (N_39809,N_36721,N_37436);
xor U39810 (N_39810,N_36014,N_36075);
nor U39811 (N_39811,N_37464,N_37716);
nor U39812 (N_39812,N_37037,N_37405);
or U39813 (N_39813,N_36722,N_37616);
nand U39814 (N_39814,N_37449,N_36449);
nand U39815 (N_39815,N_36322,N_37704);
and U39816 (N_39816,N_36896,N_37852);
and U39817 (N_39817,N_36852,N_37413);
nand U39818 (N_39818,N_36076,N_36628);
xor U39819 (N_39819,N_37870,N_37636);
xor U39820 (N_39820,N_36907,N_37531);
xnor U39821 (N_39821,N_37008,N_37964);
nor U39822 (N_39822,N_36279,N_36353);
nor U39823 (N_39823,N_37295,N_36243);
nand U39824 (N_39824,N_36258,N_36748);
xor U39825 (N_39825,N_37558,N_36676);
or U39826 (N_39826,N_37150,N_37417);
nand U39827 (N_39827,N_37597,N_36089);
nor U39828 (N_39828,N_36207,N_37474);
and U39829 (N_39829,N_37939,N_37699);
nand U39830 (N_39830,N_36301,N_37455);
nand U39831 (N_39831,N_37414,N_37459);
or U39832 (N_39832,N_36836,N_36100);
or U39833 (N_39833,N_36846,N_36587);
nor U39834 (N_39834,N_36855,N_37620);
and U39835 (N_39835,N_36654,N_36802);
xor U39836 (N_39836,N_36366,N_37896);
and U39837 (N_39837,N_36626,N_37260);
and U39838 (N_39838,N_36171,N_37270);
xnor U39839 (N_39839,N_36794,N_36662);
xor U39840 (N_39840,N_36280,N_36813);
nand U39841 (N_39841,N_36935,N_36823);
nor U39842 (N_39842,N_37773,N_36197);
nor U39843 (N_39843,N_37222,N_36022);
and U39844 (N_39844,N_36486,N_36190);
and U39845 (N_39845,N_36689,N_37547);
or U39846 (N_39846,N_36814,N_36841);
nand U39847 (N_39847,N_36982,N_37187);
or U39848 (N_39848,N_37143,N_36801);
or U39849 (N_39849,N_36504,N_36498);
xnor U39850 (N_39850,N_36718,N_36749);
and U39851 (N_39851,N_36173,N_36413);
nor U39852 (N_39852,N_36692,N_37416);
nand U39853 (N_39853,N_37671,N_37612);
nor U39854 (N_39854,N_37031,N_36703);
nand U39855 (N_39855,N_37300,N_36057);
xnor U39856 (N_39856,N_37520,N_36828);
xnor U39857 (N_39857,N_36366,N_36160);
xor U39858 (N_39858,N_36170,N_36580);
or U39859 (N_39859,N_36552,N_36744);
and U39860 (N_39860,N_36812,N_37756);
nor U39861 (N_39861,N_36503,N_37911);
nor U39862 (N_39862,N_36859,N_37397);
and U39863 (N_39863,N_37819,N_36935);
xnor U39864 (N_39864,N_37701,N_37396);
nand U39865 (N_39865,N_36702,N_36687);
nand U39866 (N_39866,N_37764,N_36325);
and U39867 (N_39867,N_36056,N_36231);
xnor U39868 (N_39868,N_36986,N_37220);
xnor U39869 (N_39869,N_36964,N_36358);
nand U39870 (N_39870,N_37063,N_36063);
xor U39871 (N_39871,N_36850,N_36089);
or U39872 (N_39872,N_36640,N_37501);
nor U39873 (N_39873,N_37570,N_37187);
or U39874 (N_39874,N_36497,N_36786);
and U39875 (N_39875,N_36356,N_37776);
or U39876 (N_39876,N_36278,N_37937);
or U39877 (N_39877,N_36963,N_37973);
nand U39878 (N_39878,N_37685,N_36497);
nand U39879 (N_39879,N_36302,N_37932);
or U39880 (N_39880,N_37393,N_37436);
or U39881 (N_39881,N_36716,N_36257);
xor U39882 (N_39882,N_37731,N_37942);
and U39883 (N_39883,N_37729,N_37168);
nor U39884 (N_39884,N_37777,N_37534);
and U39885 (N_39885,N_37986,N_36413);
nor U39886 (N_39886,N_36018,N_37823);
nand U39887 (N_39887,N_37089,N_37126);
or U39888 (N_39888,N_36649,N_36447);
nor U39889 (N_39889,N_37061,N_37541);
and U39890 (N_39890,N_37579,N_36799);
and U39891 (N_39891,N_37820,N_36282);
and U39892 (N_39892,N_36786,N_37386);
xnor U39893 (N_39893,N_36338,N_36268);
nand U39894 (N_39894,N_37922,N_36526);
xnor U39895 (N_39895,N_37893,N_36914);
xnor U39896 (N_39896,N_36209,N_37621);
nor U39897 (N_39897,N_37931,N_37487);
nor U39898 (N_39898,N_36618,N_37881);
nor U39899 (N_39899,N_37334,N_37944);
and U39900 (N_39900,N_36806,N_37780);
and U39901 (N_39901,N_36571,N_37078);
xor U39902 (N_39902,N_36592,N_36607);
or U39903 (N_39903,N_37965,N_36176);
xnor U39904 (N_39904,N_36112,N_37302);
and U39905 (N_39905,N_37645,N_36386);
xnor U39906 (N_39906,N_37455,N_36863);
nand U39907 (N_39907,N_37720,N_37138);
nand U39908 (N_39908,N_37877,N_37644);
xnor U39909 (N_39909,N_37402,N_36385);
xor U39910 (N_39910,N_37799,N_36210);
and U39911 (N_39911,N_36460,N_37938);
and U39912 (N_39912,N_37168,N_36646);
xnor U39913 (N_39913,N_37370,N_36654);
nand U39914 (N_39914,N_36575,N_36477);
nor U39915 (N_39915,N_36680,N_36665);
nand U39916 (N_39916,N_36807,N_36099);
xnor U39917 (N_39917,N_36214,N_37961);
or U39918 (N_39918,N_37328,N_36187);
xnor U39919 (N_39919,N_36758,N_36588);
xor U39920 (N_39920,N_36669,N_36638);
nand U39921 (N_39921,N_36989,N_36880);
nand U39922 (N_39922,N_37576,N_37710);
nand U39923 (N_39923,N_37687,N_36742);
and U39924 (N_39924,N_37662,N_36218);
or U39925 (N_39925,N_36409,N_36595);
nand U39926 (N_39926,N_37304,N_36247);
xor U39927 (N_39927,N_36669,N_36189);
xnor U39928 (N_39928,N_37163,N_36737);
xnor U39929 (N_39929,N_36635,N_36076);
xor U39930 (N_39930,N_37503,N_37478);
xnor U39931 (N_39931,N_36458,N_36601);
and U39932 (N_39932,N_37496,N_37595);
nor U39933 (N_39933,N_37786,N_37722);
nor U39934 (N_39934,N_37276,N_36535);
nor U39935 (N_39935,N_37799,N_36760);
xor U39936 (N_39936,N_37130,N_37825);
and U39937 (N_39937,N_37318,N_37552);
or U39938 (N_39938,N_37582,N_37836);
and U39939 (N_39939,N_36709,N_37171);
xor U39940 (N_39940,N_36726,N_36366);
nor U39941 (N_39941,N_36686,N_37403);
or U39942 (N_39942,N_36159,N_37793);
nor U39943 (N_39943,N_36523,N_37504);
xor U39944 (N_39944,N_36467,N_36584);
or U39945 (N_39945,N_36282,N_36470);
nor U39946 (N_39946,N_36151,N_37642);
and U39947 (N_39947,N_36759,N_37569);
nor U39948 (N_39948,N_36887,N_37662);
or U39949 (N_39949,N_37241,N_37563);
or U39950 (N_39950,N_36392,N_37646);
or U39951 (N_39951,N_36494,N_37575);
or U39952 (N_39952,N_37271,N_36024);
nand U39953 (N_39953,N_36209,N_36469);
nand U39954 (N_39954,N_37982,N_37966);
nand U39955 (N_39955,N_37990,N_36979);
nor U39956 (N_39956,N_37076,N_37780);
and U39957 (N_39957,N_36611,N_36702);
nand U39958 (N_39958,N_37372,N_36463);
and U39959 (N_39959,N_36422,N_36484);
or U39960 (N_39960,N_36210,N_36293);
or U39961 (N_39961,N_36185,N_37792);
and U39962 (N_39962,N_36430,N_37850);
xor U39963 (N_39963,N_36561,N_37217);
and U39964 (N_39964,N_37126,N_36005);
and U39965 (N_39965,N_37968,N_36867);
xor U39966 (N_39966,N_37688,N_36941);
or U39967 (N_39967,N_36413,N_36725);
nand U39968 (N_39968,N_36276,N_36222);
nand U39969 (N_39969,N_37520,N_36146);
and U39970 (N_39970,N_37136,N_36571);
nor U39971 (N_39971,N_37298,N_37751);
or U39972 (N_39972,N_36136,N_37224);
and U39973 (N_39973,N_37595,N_36059);
nor U39974 (N_39974,N_36602,N_37466);
and U39975 (N_39975,N_36657,N_37698);
and U39976 (N_39976,N_36140,N_36608);
and U39977 (N_39977,N_37474,N_36153);
nand U39978 (N_39978,N_36491,N_37208);
nand U39979 (N_39979,N_36495,N_36535);
nor U39980 (N_39980,N_37440,N_37072);
xor U39981 (N_39981,N_37411,N_36847);
and U39982 (N_39982,N_37011,N_37168);
nor U39983 (N_39983,N_36214,N_36423);
xnor U39984 (N_39984,N_36118,N_37890);
and U39985 (N_39985,N_37986,N_36874);
and U39986 (N_39986,N_36260,N_36793);
xor U39987 (N_39987,N_36973,N_36602);
nor U39988 (N_39988,N_37442,N_36265);
or U39989 (N_39989,N_36622,N_37697);
nand U39990 (N_39990,N_36882,N_36459);
nand U39991 (N_39991,N_36383,N_36313);
and U39992 (N_39992,N_36500,N_36214);
or U39993 (N_39993,N_37273,N_36644);
and U39994 (N_39994,N_36238,N_36358);
xnor U39995 (N_39995,N_36641,N_36225);
xor U39996 (N_39996,N_37117,N_37259);
nand U39997 (N_39997,N_36526,N_37574);
nand U39998 (N_39998,N_37743,N_36174);
xnor U39999 (N_39999,N_36424,N_37228);
nor U40000 (N_40000,N_39285,N_39949);
and U40001 (N_40001,N_39268,N_38862);
nor U40002 (N_40002,N_38953,N_38001);
and U40003 (N_40003,N_38639,N_39388);
or U40004 (N_40004,N_38514,N_38722);
nor U40005 (N_40005,N_38534,N_39620);
nor U40006 (N_40006,N_38602,N_38334);
xnor U40007 (N_40007,N_39514,N_39551);
nand U40008 (N_40008,N_38116,N_39505);
or U40009 (N_40009,N_38033,N_38053);
nand U40010 (N_40010,N_38621,N_38336);
or U40011 (N_40011,N_39115,N_39701);
nand U40012 (N_40012,N_38876,N_39069);
nor U40013 (N_40013,N_39729,N_39479);
and U40014 (N_40014,N_38966,N_39908);
nor U40015 (N_40015,N_39386,N_39537);
nor U40016 (N_40016,N_39400,N_38441);
and U40017 (N_40017,N_39453,N_39432);
nand U40018 (N_40018,N_38932,N_39234);
and U40019 (N_40019,N_38279,N_39936);
and U40020 (N_40020,N_38617,N_39473);
nor U40021 (N_40021,N_38111,N_39890);
or U40022 (N_40022,N_38578,N_38773);
nor U40023 (N_40023,N_38775,N_39506);
xnor U40024 (N_40024,N_38102,N_38415);
or U40025 (N_40025,N_38086,N_39630);
nand U40026 (N_40026,N_38819,N_38791);
and U40027 (N_40027,N_38962,N_39963);
and U40028 (N_40028,N_39844,N_38297);
nor U40029 (N_40029,N_39112,N_38287);
and U40030 (N_40030,N_39725,N_38869);
nor U40031 (N_40031,N_38409,N_39222);
xnor U40032 (N_40032,N_38337,N_39328);
nor U40033 (N_40033,N_39539,N_39674);
nand U40034 (N_40034,N_39612,N_38364);
or U40035 (N_40035,N_39988,N_38741);
xnor U40036 (N_40036,N_39044,N_38531);
nand U40037 (N_40037,N_38906,N_39290);
nand U40038 (N_40038,N_38206,N_38315);
xor U40039 (N_40039,N_39102,N_38044);
nand U40040 (N_40040,N_38007,N_39028);
nor U40041 (N_40041,N_39590,N_38525);
xor U40042 (N_40042,N_39089,N_38668);
or U40043 (N_40043,N_39640,N_39039);
xnor U40044 (N_40044,N_39792,N_38834);
or U40045 (N_40045,N_38731,N_39848);
xor U40046 (N_40046,N_39648,N_38547);
and U40047 (N_40047,N_38931,N_39944);
or U40048 (N_40048,N_39957,N_38255);
nand U40049 (N_40049,N_38324,N_39472);
nand U40050 (N_40050,N_38625,N_38783);
nand U40051 (N_40051,N_39727,N_38307);
nor U40052 (N_40052,N_39356,N_39430);
xor U40053 (N_40053,N_38199,N_38978);
xnor U40054 (N_40054,N_38513,N_38339);
or U40055 (N_40055,N_38763,N_38034);
nor U40056 (N_40056,N_38943,N_38915);
nor U40057 (N_40057,N_38040,N_38855);
and U40058 (N_40058,N_38887,N_38490);
and U40059 (N_40059,N_39969,N_38495);
xnor U40060 (N_40060,N_38976,N_39993);
xnor U40061 (N_40061,N_38167,N_39183);
or U40062 (N_40062,N_39859,N_38839);
and U40063 (N_40063,N_39558,N_39423);
or U40064 (N_40064,N_39906,N_38325);
xnor U40065 (N_40065,N_38888,N_38186);
xnor U40066 (N_40066,N_39520,N_39713);
nand U40067 (N_40067,N_39035,N_38394);
xor U40068 (N_40068,N_39878,N_39835);
and U40069 (N_40069,N_38121,N_38142);
and U40070 (N_40070,N_39099,N_38784);
xor U40071 (N_40071,N_39469,N_39278);
nand U40072 (N_40072,N_38759,N_38940);
or U40073 (N_40073,N_38450,N_38429);
nand U40074 (N_40074,N_39735,N_38311);
xor U40075 (N_40075,N_38359,N_38354);
or U40076 (N_40076,N_39308,N_38042);
nand U40077 (N_40077,N_38821,N_38192);
and U40078 (N_40078,N_39580,N_38859);
or U40079 (N_40079,N_39646,N_38812);
or U40080 (N_40080,N_39962,N_38865);
nand U40081 (N_40081,N_39402,N_39641);
xor U40082 (N_40082,N_38463,N_38335);
nor U40083 (N_40083,N_39446,N_38210);
xnor U40084 (N_40084,N_38628,N_38293);
or U40085 (N_40085,N_38390,N_39912);
or U40086 (N_40086,N_39139,N_39953);
and U40087 (N_40087,N_39935,N_38381);
and U40088 (N_40088,N_38348,N_39360);
nand U40089 (N_40089,N_38250,N_39510);
nor U40090 (N_40090,N_39952,N_39869);
nand U40091 (N_40091,N_38949,N_39632);
nor U40092 (N_40092,N_39318,N_39773);
nor U40093 (N_40093,N_39030,N_38267);
nor U40094 (N_40094,N_39608,N_38332);
nand U40095 (N_40095,N_39536,N_39354);
nor U40096 (N_40096,N_39732,N_38938);
nand U40097 (N_40097,N_39972,N_38119);
nor U40098 (N_40098,N_38070,N_39829);
nor U40099 (N_40099,N_39097,N_38384);
or U40100 (N_40100,N_39160,N_39081);
xor U40101 (N_40101,N_38961,N_39295);
or U40102 (N_40102,N_39678,N_38930);
and U40103 (N_40103,N_38201,N_38769);
and U40104 (N_40104,N_39165,N_38360);
xnor U40105 (N_40105,N_38643,N_38471);
nor U40106 (N_40106,N_39574,N_39049);
or U40107 (N_40107,N_38678,N_39748);
nand U40108 (N_40108,N_39372,N_38137);
or U40109 (N_40109,N_38144,N_39696);
and U40110 (N_40110,N_39843,N_39679);
nand U40111 (N_40111,N_39794,N_39344);
or U40112 (N_40112,N_39670,N_39982);
nor U40113 (N_40113,N_39553,N_39872);
xor U40114 (N_40114,N_39359,N_38350);
xnor U40115 (N_40115,N_39105,N_39597);
or U40116 (N_40116,N_38130,N_39519);
xnor U40117 (N_40117,N_39206,N_38136);
nand U40118 (N_40118,N_39444,N_39243);
nor U40119 (N_40119,N_38713,N_38357);
and U40120 (N_40120,N_39304,N_39686);
nor U40121 (N_40121,N_39577,N_39650);
xnor U40122 (N_40122,N_39380,N_38173);
xor U40123 (N_40123,N_39016,N_38992);
xnor U40124 (N_40124,N_39639,N_38528);
nand U40125 (N_40125,N_38328,N_39364);
and U40126 (N_40126,N_38899,N_38893);
or U40127 (N_40127,N_38951,N_39482);
nor U40128 (N_40128,N_38470,N_38813);
nor U40129 (N_40129,N_38959,N_38043);
and U40130 (N_40130,N_39762,N_39722);
nor U40131 (N_40131,N_39447,N_39591);
xnor U40132 (N_40132,N_38372,N_39256);
or U40133 (N_40133,N_38977,N_39187);
and U40134 (N_40134,N_39275,N_38377);
nand U40135 (N_40135,N_39699,N_39156);
nor U40136 (N_40136,N_38836,N_38541);
nor U40137 (N_40137,N_38714,N_38113);
and U40138 (N_40138,N_38687,N_39778);
and U40139 (N_40139,N_39951,N_38934);
xor U40140 (N_40140,N_39260,N_38736);
or U40141 (N_40141,N_39994,N_39258);
nor U40142 (N_40142,N_38818,N_38724);
nor U40143 (N_40143,N_38342,N_38219);
nor U40144 (N_40144,N_38706,N_39368);
nand U40145 (N_40145,N_39079,N_39436);
and U40146 (N_40146,N_39034,N_38046);
and U40147 (N_40147,N_38669,N_38999);
nor U40148 (N_40148,N_39152,N_38543);
nand U40149 (N_40149,N_39512,N_38413);
or U40150 (N_40150,N_38389,N_39917);
xor U40151 (N_40151,N_39731,N_39253);
nor U40152 (N_40152,N_38875,N_39871);
or U40153 (N_40153,N_39642,N_39876);
xnor U40154 (N_40154,N_39895,N_39784);
nor U40155 (N_40155,N_38964,N_38952);
nor U40156 (N_40156,N_38627,N_38442);
and U40157 (N_40157,N_38268,N_39130);
or U40158 (N_40158,N_39978,N_39932);
or U40159 (N_40159,N_38633,N_39022);
xor U40160 (N_40160,N_39687,N_38764);
xnor U40161 (N_40161,N_39411,N_38634);
or U40162 (N_40162,N_39307,N_38516);
and U40163 (N_40163,N_38803,N_39154);
and U40164 (N_40164,N_38274,N_39006);
nand U40165 (N_40165,N_38971,N_38935);
and U40166 (N_40166,N_39570,N_39269);
xor U40167 (N_40167,N_39974,N_38527);
and U40168 (N_40168,N_38025,N_38011);
nand U40169 (N_40169,N_39730,N_39343);
or U40170 (N_40170,N_39733,N_39420);
or U40171 (N_40171,N_38449,N_38766);
or U40172 (N_40172,N_38807,N_38707);
nand U40173 (N_40173,N_38472,N_38697);
nand U40174 (N_40174,N_39144,N_39922);
xor U40175 (N_40175,N_38896,N_39149);
and U40176 (N_40176,N_39804,N_39349);
or U40177 (N_40177,N_39490,N_39973);
and U40178 (N_40178,N_39645,N_38781);
or U40179 (N_40179,N_38510,N_39476);
xor U40180 (N_40180,N_39567,N_38169);
xor U40181 (N_40181,N_38521,N_38092);
or U40182 (N_40182,N_38631,N_38462);
nand U40183 (N_40183,N_38566,N_39373);
nand U40184 (N_40184,N_39726,N_38588);
xor U40185 (N_40185,N_39720,N_38619);
nor U40186 (N_40186,N_39717,N_38770);
xor U40187 (N_40187,N_39823,N_39413);
nor U40188 (N_40188,N_38878,N_39709);
xnor U40189 (N_40189,N_38217,N_39799);
and U40190 (N_40190,N_39695,N_39104);
xor U40191 (N_40191,N_39262,N_39090);
xnor U40192 (N_40192,N_38845,N_38605);
and U40193 (N_40193,N_39058,N_38872);
nor U40194 (N_40194,N_38782,N_38558);
and U40195 (N_40195,N_39867,N_38738);
and U40196 (N_40196,N_38361,N_39404);
xnor U40197 (N_40197,N_39239,N_39885);
nand U40198 (N_40198,N_38141,N_38079);
nor U40199 (N_40199,N_38258,N_38433);
xnor U40200 (N_40200,N_39460,N_39854);
nand U40201 (N_40201,N_38316,N_39884);
and U40202 (N_40202,N_39497,N_38810);
and U40203 (N_40203,N_39427,N_38114);
nor U40204 (N_40204,N_38860,N_38115);
nor U40205 (N_40205,N_39579,N_39273);
xor U40206 (N_40206,N_38642,N_38582);
xor U40207 (N_40207,N_39348,N_38680);
and U40208 (N_40208,N_39248,N_39896);
xnor U40209 (N_40209,N_39389,N_38066);
and U40210 (N_40210,N_38160,N_38446);
or U40211 (N_40211,N_38383,N_38022);
nand U40212 (N_40212,N_38914,N_38685);
nand U40213 (N_40213,N_38800,N_38587);
nand U40214 (N_40214,N_39029,N_39394);
nand U40215 (N_40215,N_38660,N_38499);
and U40216 (N_40216,N_38264,N_39441);
and U40217 (N_40217,N_38254,N_39055);
and U40218 (N_40218,N_38211,N_38956);
xor U40219 (N_40219,N_39213,N_39439);
nor U40220 (N_40220,N_39673,N_38006);
nand U40221 (N_40221,N_39184,N_38132);
xor U40222 (N_40222,N_38289,N_38973);
or U40223 (N_40223,N_38322,N_38380);
nand U40224 (N_40224,N_39337,N_38607);
and U40225 (N_40225,N_39527,N_38234);
xnor U40226 (N_40226,N_39877,N_38576);
nand U40227 (N_40227,N_38400,N_39397);
or U40228 (N_40228,N_38581,N_39970);
and U40229 (N_40229,N_39740,N_39244);
and U40230 (N_40230,N_38184,N_38411);
or U40231 (N_40231,N_39488,N_38494);
nand U40232 (N_40232,N_38873,N_38776);
nand U40233 (N_40233,N_38879,N_38849);
and U40234 (N_40234,N_39150,N_39875);
xor U40235 (N_40235,N_38843,N_39301);
or U40236 (N_40236,N_38712,N_38670);
nor U40237 (N_40237,N_38591,N_39818);
nand U40238 (N_40238,N_39326,N_38134);
nor U40239 (N_40239,N_38138,N_38950);
and U40240 (N_40240,N_39571,N_39466);
or U40241 (N_40241,N_38280,N_38650);
and U40242 (N_40242,N_39496,N_39874);
xor U40243 (N_40243,N_39279,N_38095);
and U40244 (N_40244,N_39606,N_38064);
nor U40245 (N_40245,N_39137,N_39605);
nor U40246 (N_40246,N_39667,N_38735);
xnor U40247 (N_40247,N_39904,N_39452);
or U40248 (N_40248,N_39363,N_39398);
nand U40249 (N_40249,N_39220,N_39849);
xor U40250 (N_40250,N_39371,N_39418);
and U40251 (N_40251,N_38557,N_39437);
and U40252 (N_40252,N_39161,N_39199);
and U40253 (N_40253,N_39937,N_39544);
nand U40254 (N_40254,N_38031,N_39414);
and U40255 (N_40255,N_39950,N_39508);
and U40256 (N_40256,N_38886,N_38601);
or U40257 (N_40257,N_38148,N_38907);
or U40258 (N_40258,N_38209,N_38191);
or U40259 (N_40259,N_38594,N_38029);
and U40260 (N_40260,N_38434,N_39095);
or U40261 (N_40261,N_38613,N_38507);
and U40262 (N_40262,N_38427,N_39143);
nor U40263 (N_40263,N_38985,N_38272);
nor U40264 (N_40264,N_38406,N_39485);
xor U40265 (N_40265,N_39500,N_38754);
nand U40266 (N_40266,N_38676,N_38816);
or U40267 (N_40267,N_39048,N_38479);
xnor U40268 (N_40268,N_38901,N_39647);
nand U40269 (N_40269,N_38146,N_39535);
or U40270 (N_40270,N_39332,N_39955);
nor U40271 (N_40271,N_38397,N_38238);
nor U40272 (N_40272,N_38767,N_39123);
and U40273 (N_40273,N_38986,N_38969);
nand U40274 (N_40274,N_39942,N_39353);
and U40275 (N_40275,N_38889,N_39880);
and U40276 (N_40276,N_39438,N_38058);
and U40277 (N_40277,N_39663,N_39925);
or U40278 (N_40278,N_38057,N_39791);
nor U40279 (N_40279,N_38363,N_39769);
and U40280 (N_40280,N_39153,N_39031);
and U40281 (N_40281,N_38379,N_39565);
or U40282 (N_40282,N_38653,N_38532);
xnor U40283 (N_40283,N_38981,N_38681);
nand U40284 (N_40284,N_39627,N_39036);
nor U40285 (N_40285,N_39111,N_39756);
or U40286 (N_40286,N_39546,N_39440);
nor U40287 (N_40287,N_38538,N_39464);
xnor U40288 (N_40288,N_38651,N_38671);
nand U40289 (N_40289,N_38298,N_39201);
or U40290 (N_40290,N_39550,N_39008);
or U40291 (N_40291,N_39093,N_38161);
or U40292 (N_40292,N_38202,N_39074);
and U40293 (N_40293,N_39077,N_39327);
nand U40294 (N_40294,N_39812,N_39212);
or U40295 (N_40295,N_39666,N_39879);
nand U40296 (N_40296,N_38672,N_38301);
xnor U40297 (N_40297,N_38624,N_38028);
xor U40298 (N_40298,N_38103,N_39826);
nor U40299 (N_40299,N_39596,N_39007);
xnor U40300 (N_40300,N_38850,N_39738);
xor U40301 (N_40301,N_39832,N_38502);
nand U40302 (N_40302,N_38019,N_39379);
nand U40303 (N_40303,N_39797,N_39277);
nor U40304 (N_40304,N_38485,N_39080);
nor U40305 (N_40305,N_38285,N_39001);
nor U40306 (N_40306,N_39698,N_38644);
and U40307 (N_40307,N_39292,N_39893);
xnor U40308 (N_40308,N_38038,N_39405);
nor U40309 (N_40309,N_38047,N_39498);
xor U40310 (N_40310,N_39185,N_39624);
xnor U40311 (N_40311,N_38895,N_39208);
and U40312 (N_40312,N_39889,N_38259);
nor U40313 (N_40313,N_38151,N_39693);
and U40314 (N_40314,N_38108,N_38078);
or U40315 (N_40315,N_38590,N_39233);
xor U40316 (N_40316,N_39316,N_39158);
nor U40317 (N_40317,N_39902,N_39059);
nor U40318 (N_40318,N_39860,N_39822);
nand U40319 (N_40319,N_39559,N_39254);
xor U40320 (N_40320,N_38154,N_38798);
nand U40321 (N_40321,N_39324,N_38864);
nand U40322 (N_40322,N_38375,N_39845);
nand U40323 (N_40323,N_38744,N_38330);
or U40324 (N_40324,N_38743,N_38778);
or U40325 (N_40325,N_39930,N_39956);
nor U40326 (N_40326,N_38240,N_38693);
and U40327 (N_40327,N_39480,N_38858);
nor U40328 (N_40328,N_38002,N_39032);
and U40329 (N_40329,N_38245,N_39734);
and U40330 (N_40330,N_39120,N_39263);
or U40331 (N_40331,N_39406,N_39494);
and U40332 (N_40332,N_39065,N_39232);
xor U40333 (N_40333,N_38493,N_39305);
or U40334 (N_40334,N_39655,N_39689);
or U40335 (N_40335,N_38270,N_38623);
nor U40336 (N_40336,N_39657,N_38674);
or U40337 (N_40337,N_39037,N_38975);
and U40338 (N_40338,N_39317,N_39023);
xnor U40339 (N_40339,N_39331,N_39294);
or U40340 (N_40340,N_38995,N_38739);
xor U40341 (N_40341,N_39217,N_38478);
nor U40342 (N_40342,N_39366,N_39227);
and U40343 (N_40343,N_38861,N_38117);
xnor U40344 (N_40344,N_38524,N_39786);
nand U40345 (N_40345,N_38517,N_39827);
nand U40346 (N_40346,N_39330,N_39600);
nor U40347 (N_40347,N_39881,N_39598);
and U40348 (N_40348,N_38451,N_39766);
nand U40349 (N_40349,N_39374,N_39919);
xor U40350 (N_40350,N_39395,N_39259);
or U40351 (N_40351,N_39795,N_38970);
nand U40352 (N_40352,N_39928,N_38753);
nand U40353 (N_40353,N_38720,N_39126);
xnor U40354 (N_40354,N_38376,N_38804);
nand U40355 (N_40355,N_38395,N_39564);
or U40356 (N_40356,N_38501,N_38868);
xor U40357 (N_40357,N_38159,N_38829);
xor U40358 (N_40358,N_39736,N_38438);
nor U40359 (N_40359,N_38455,N_38750);
or U40360 (N_40360,N_39214,N_38640);
xnor U40361 (N_40361,N_39399,N_39475);
nand U40362 (N_40362,N_39357,N_38902);
or U40363 (N_40363,N_39724,N_38329);
nand U40364 (N_40364,N_39041,N_38948);
or U40365 (N_40365,N_39462,N_38247);
xnor U40366 (N_40366,N_39671,N_38133);
nor U40367 (N_40367,N_38326,N_38378);
nor U40368 (N_40368,N_39096,N_39189);
and U40369 (N_40369,N_38487,N_38425);
nand U40370 (N_40370,N_39749,N_38123);
nand U40371 (N_40371,N_39060,N_38874);
nand U40372 (N_40372,N_39387,N_39816);
or U40373 (N_40373,N_39581,N_38283);
or U40374 (N_40374,N_38120,N_38215);
and U40375 (N_40375,N_39367,N_39470);
or U40376 (N_40376,N_39716,N_38393);
xnor U40377 (N_40377,N_39021,N_39803);
and U40378 (N_40378,N_39604,N_39834);
or U40379 (N_40379,N_39790,N_38016);
and U40380 (N_40380,N_39654,N_39517);
nor U40381 (N_40381,N_38333,N_39163);
or U40382 (N_40382,N_38128,N_38341);
nor U40383 (N_40383,N_39168,N_38165);
or U40384 (N_40384,N_38994,N_38924);
or U40385 (N_40385,N_39776,N_38984);
nand U40386 (N_40386,N_39613,N_39133);
xnor U40387 (N_40387,N_38577,N_38012);
and U40388 (N_40388,N_39000,N_38796);
nor U40389 (N_40389,N_39659,N_38068);
or U40390 (N_40390,N_39824,N_38340);
or U40391 (N_40391,N_39455,N_39562);
xnor U40392 (N_40392,N_39057,N_39499);
xor U40393 (N_40393,N_39677,N_39429);
or U40394 (N_40394,N_39151,N_39311);
xor U40395 (N_40395,N_39718,N_38936);
xnor U40396 (N_40396,N_38831,N_38508);
or U40397 (N_40397,N_39690,N_39381);
nor U40398 (N_40398,N_39511,N_39252);
nand U40399 (N_40399,N_39628,N_38657);
and U40400 (N_40400,N_39898,N_38917);
or U40401 (N_40401,N_39410,N_38539);
or U40402 (N_40402,N_39013,N_38912);
nand U40403 (N_40403,N_38570,N_39665);
and U40404 (N_40404,N_38916,N_39779);
and U40405 (N_40405,N_38545,N_38909);
xnor U40406 (N_40406,N_38407,N_38903);
and U40407 (N_40407,N_39382,N_39393);
or U40408 (N_40408,N_38062,N_38905);
or U40409 (N_40409,N_38371,N_39159);
and U40410 (N_40410,N_38152,N_39342);
xnor U40411 (N_40411,N_39662,N_38846);
nand U40412 (N_40412,N_38841,N_38039);
nand U40413 (N_40413,N_39319,N_39107);
nor U40414 (N_40414,N_38466,N_39523);
or U40415 (N_40415,N_39723,N_38468);
nand U40416 (N_40416,N_39618,N_38820);
or U40417 (N_40417,N_38749,N_38511);
nor U40418 (N_40418,N_38880,N_39235);
xor U40419 (N_40419,N_39180,N_39284);
and U40420 (N_40420,N_38913,N_39421);
nand U40421 (N_40421,N_39968,N_38178);
and U40422 (N_40422,N_39224,N_39538);
and U40423 (N_40423,N_38465,N_38638);
xor U40424 (N_40424,N_39043,N_38540);
or U40425 (N_40425,N_38554,N_39954);
nor U40426 (N_40426,N_39179,N_38691);
nor U40427 (N_40427,N_38368,N_39484);
xor U40428 (N_40428,N_38195,N_39417);
nor U40429 (N_40429,N_38645,N_38811);
nor U40430 (N_40430,N_38049,N_39010);
nor U40431 (N_40431,N_38248,N_38760);
and U40432 (N_40432,N_39811,N_39383);
or U40433 (N_40433,N_39793,N_39114);
or U40434 (N_40434,N_38980,N_38310);
or U40435 (N_40435,N_38282,N_39191);
and U40436 (N_40436,N_38945,N_38097);
xor U40437 (N_40437,N_38428,N_39599);
and U40438 (N_40438,N_39578,N_38147);
or U40439 (N_40439,N_39664,N_38614);
and U40440 (N_40440,N_39549,N_39063);
nor U40441 (N_40441,N_38193,N_39743);
or U40442 (N_40442,N_39467,N_39231);
and U40443 (N_40443,N_39422,N_39245);
nand U40444 (N_40444,N_39712,N_39503);
or U40445 (N_40445,N_38610,N_39901);
nor U40446 (N_40446,N_39487,N_39471);
nand U40447 (N_40447,N_39219,N_38233);
or U40448 (N_40448,N_39370,N_38535);
nor U40449 (N_40449,N_39109,N_38606);
and U40450 (N_40450,N_38126,N_38740);
nor U40451 (N_40451,N_39335,N_38317);
xnor U40452 (N_40452,N_38942,N_38491);
nor U40453 (N_40453,N_39548,N_38923);
nor U40454 (N_40454,N_39346,N_38983);
or U40455 (N_40455,N_38871,N_38220);
and U40456 (N_40456,N_38157,N_38974);
nand U40457 (N_40457,N_38496,N_38822);
nand U40458 (N_40458,N_39146,N_39250);
nand U40459 (N_40459,N_38608,N_39171);
and U40460 (N_40460,N_38515,N_39148);
nand U40461 (N_40461,N_38960,N_38399);
nor U40462 (N_40462,N_38051,N_38222);
and U40463 (N_40463,N_38085,N_38338);
and U40464 (N_40464,N_39333,N_38682);
and U40465 (N_40465,N_39173,N_38140);
or U40466 (N_40466,N_38221,N_39113);
and U40467 (N_40467,N_38904,N_38504);
nor U40468 (N_40468,N_38814,N_38698);
or U40469 (N_40469,N_38344,N_39967);
xor U40470 (N_40470,N_38799,N_38615);
xor U40471 (N_40471,N_38703,N_38098);
nand U40472 (N_40472,N_38562,N_38198);
or U40473 (N_40473,N_39325,N_39237);
xor U40474 (N_40474,N_38089,N_39061);
and U40475 (N_40475,N_38063,N_39323);
or U40476 (N_40476,N_38305,N_38537);
nor U40477 (N_40477,N_38592,N_38990);
and U40478 (N_40478,N_39905,N_39862);
nor U40479 (N_40479,N_38278,N_38244);
nor U40480 (N_40480,N_38690,N_38398);
and U40481 (N_40481,N_39086,N_38852);
nor U40482 (N_40482,N_39450,N_38055);
and U40483 (N_40483,N_38241,N_38786);
nand U40484 (N_40484,N_38461,N_39443);
and U40485 (N_40485,N_38143,N_39991);
and U40486 (N_40486,N_39226,N_38838);
nor U40487 (N_40487,N_39170,N_38667);
nand U40488 (N_40488,N_38734,N_39981);
xnor U40489 (N_40489,N_39434,N_38401);
or U40490 (N_40490,N_39339,N_38452);
nor U40491 (N_40491,N_39755,N_38729);
nor U40492 (N_40492,N_39300,N_39513);
and U40493 (N_40493,N_38751,N_38069);
nor U40494 (N_40494,N_38701,N_38505);
nor U40495 (N_40495,N_38937,N_39412);
or U40496 (N_40496,N_38027,N_39110);
nand U40497 (N_40497,N_38373,N_39176);
nor U40498 (N_40498,N_38200,N_39817);
nand U40499 (N_40499,N_38780,N_39986);
nand U40500 (N_40500,N_38454,N_38742);
nand U40501 (N_40501,N_38844,N_39236);
or U40502 (N_40502,N_38024,N_39918);
nand U40503 (N_40503,N_39005,N_39660);
nand U40504 (N_40504,N_38149,N_38794);
nand U40505 (N_40505,N_39873,N_38403);
nand U40506 (N_40506,N_39045,N_39836);
nand U40507 (N_40507,N_39280,N_39744);
nand U40508 (N_40508,N_39561,N_39758);
or U40509 (N_40509,N_39251,N_39644);
nor U40510 (N_40510,N_38444,N_39965);
xnor U40511 (N_40511,N_38396,N_39341);
or U40512 (N_40512,N_39672,N_38806);
xor U40513 (N_40513,N_39933,N_38700);
or U40514 (N_40514,N_38519,N_38789);
nand U40515 (N_40515,N_39938,N_38544);
or U40516 (N_40516,N_38498,N_39092);
xnor U40517 (N_40517,N_38300,N_39197);
nor U40518 (N_40518,N_38883,N_39478);
xor U40519 (N_40519,N_38431,N_39853);
or U40520 (N_40520,N_39491,N_38559);
or U40521 (N_40521,N_39589,N_38177);
nor U40522 (N_40522,N_38237,N_38072);
nand U40523 (N_40523,N_38797,N_38979);
and U40524 (N_40524,N_39637,N_38677);
nor U40525 (N_40525,N_38929,N_39653);
nor U40526 (N_40526,N_39416,N_38847);
or U40527 (N_40527,N_38367,N_38546);
nand U40528 (N_40528,N_38223,N_38721);
and U40529 (N_40529,N_39392,N_39507);
xor U40530 (N_40530,N_38166,N_38302);
nand U40531 (N_40531,N_38856,N_39456);
nor U40532 (N_40532,N_39706,N_38885);
xnor U40533 (N_40533,N_38652,N_39775);
nand U40534 (N_40534,N_39682,N_38374);
xor U40535 (N_40535,N_38281,N_38972);
nor U40536 (N_40536,N_38648,N_39495);
and U40537 (N_40537,N_38686,N_39566);
and U40538 (N_40538,N_39155,N_38620);
nor U40539 (N_40539,N_39085,N_39091);
or U40540 (N_40540,N_38392,N_39136);
nand U40541 (N_40541,N_39692,N_38589);
nor U40542 (N_40542,N_39961,N_38164);
xor U40543 (N_40543,N_39934,N_38629);
or U40544 (N_40544,N_38026,N_38925);
nor U40545 (N_40545,N_38104,N_39891);
and U40546 (N_40546,N_38414,N_38197);
nand U40547 (N_40547,N_38509,N_38500);
or U40548 (N_40548,N_38107,N_38084);
and U40549 (N_40549,N_39246,N_38318);
or U40550 (N_40550,N_38075,N_39229);
or U40551 (N_40551,N_39582,N_39622);
nand U40552 (N_40552,N_39594,N_39602);
or U40553 (N_40553,N_39721,N_38356);
and U40554 (N_40554,N_38218,N_39532);
or U40555 (N_40555,N_38430,N_38189);
and U40556 (N_40556,N_39106,N_39866);
nand U40557 (N_40557,N_38649,N_38110);
nor U40558 (N_40558,N_38153,N_39593);
and U40559 (N_40559,N_38655,N_39675);
or U40560 (N_40560,N_39131,N_38939);
and U40561 (N_40561,N_39760,N_38225);
nor U40562 (N_40562,N_38658,N_38269);
xnor U40563 (N_40563,N_39850,N_39801);
xnor U40564 (N_40564,N_39752,N_38216);
nand U40565 (N_40565,N_38599,N_39068);
nor U40566 (N_40566,N_39924,N_39225);
nor U40567 (N_40567,N_39272,N_38035);
nor U40568 (N_40568,N_38569,N_39509);
and U40569 (N_40569,N_39819,N_39166);
nand U40570 (N_40570,N_38056,N_39449);
or U40571 (N_40571,N_38892,N_39528);
nand U40572 (N_40572,N_38530,N_38196);
nand U40573 (N_40573,N_38659,N_39557);
and U40574 (N_40574,N_39783,N_38512);
and U40575 (N_40575,N_39003,N_39502);
nor U40576 (N_40576,N_39157,N_38867);
or U40577 (N_40577,N_38235,N_39894);
or U40578 (N_40578,N_39631,N_39595);
xnor U40579 (N_40579,N_38911,N_39771);
nand U40580 (N_40580,N_39715,N_39182);
or U40581 (N_40581,N_38074,N_39601);
nor U40582 (N_40582,N_38564,N_38239);
nand U40583 (N_40583,N_39261,N_39680);
nand U40584 (N_40584,N_39768,N_39274);
and U40585 (N_40585,N_39424,N_38277);
xor U40586 (N_40586,N_39193,N_38275);
nand U40587 (N_40587,N_39322,N_39555);
xor U40588 (N_40588,N_38266,N_38884);
nor U40589 (N_40589,N_38603,N_38158);
xor U40590 (N_40590,N_39825,N_38405);
nor U40591 (N_40591,N_38276,N_38314);
xor U40592 (N_40592,N_38612,N_38723);
nor U40593 (N_40593,N_38853,N_39289);
or U40594 (N_40594,N_38118,N_38683);
nand U40595 (N_40595,N_39098,N_39868);
nand U40596 (N_40596,N_38477,N_39907);
nor U40597 (N_40597,N_38071,N_38857);
nand U40598 (N_40598,N_38553,N_38037);
nand U40599 (N_40599,N_38561,N_39765);
and U40600 (N_40600,N_38637,N_38163);
xnor U40601 (N_40601,N_39062,N_38632);
or U40602 (N_40602,N_38101,N_39078);
nand U40603 (N_40603,N_38369,N_38998);
or U40604 (N_40604,N_39350,N_39838);
or U40605 (N_40605,N_39587,N_39737);
or U40606 (N_40606,N_38421,N_39892);
xnor U40607 (N_40607,N_39124,N_39711);
or U40608 (N_40608,N_38257,N_38774);
or U40609 (N_40609,N_38747,N_39704);
nand U40610 (N_40610,N_38702,N_39865);
or U40611 (N_40611,N_39926,N_38646);
nor U40612 (N_40612,N_39888,N_39073);
xnor U40613 (N_40613,N_38792,N_39851);
nand U40614 (N_40614,N_38286,N_39636);
xor U40615 (N_40615,N_38982,N_39616);
xor U40616 (N_40616,N_39128,N_38437);
nand U40617 (N_40617,N_39863,N_38474);
xnor U40618 (N_40618,N_39837,N_38150);
or U40619 (N_40619,N_38746,N_39287);
nor U40620 (N_40620,N_39563,N_39805);
xnor U40621 (N_40621,N_39056,N_38256);
or U40622 (N_40622,N_38017,N_39521);
or U40623 (N_40623,N_38968,N_38492);
xor U40624 (N_40624,N_38162,N_38208);
nor U40625 (N_40625,N_39800,N_38227);
nand U40626 (N_40626,N_39188,N_39789);
xnor U40627 (N_40627,N_39267,N_39847);
or U40628 (N_40628,N_38226,N_39603);
xnor U40629 (N_40629,N_39929,N_39700);
or U40630 (N_40630,N_38520,N_38600);
nor U40631 (N_40631,N_39998,N_39483);
nor U40632 (N_40632,N_39223,N_39014);
and U40633 (N_40633,N_39831,N_39746);
xor U40634 (N_40634,N_38647,N_39534);
or U40635 (N_40635,N_39489,N_39230);
and U40636 (N_40636,N_38190,N_38963);
and U40637 (N_40637,N_39807,N_38106);
and U40638 (N_40638,N_38611,N_38699);
xnor U40639 (N_40639,N_39409,N_38684);
and U40640 (N_40640,N_39821,N_38730);
and U40641 (N_40641,N_38469,N_38583);
nor U40642 (N_40642,N_39707,N_38023);
or U40643 (N_40643,N_39377,N_39046);
nand U40644 (N_40644,N_38497,N_38726);
xor U40645 (N_40645,N_39345,N_39780);
xor U40646 (N_40646,N_38518,N_39310);
and U40647 (N_40647,N_39117,N_38788);
xnor U40648 (N_40648,N_38488,N_39750);
and U40649 (N_40649,N_38476,N_39025);
nand U40650 (N_40650,N_39669,N_39203);
and U40651 (N_40651,N_38253,N_39314);
or U40652 (N_40652,N_38382,N_39530);
nor U40653 (N_40653,N_39075,N_38848);
or U40654 (N_40654,N_38480,N_39340);
or U40655 (N_40655,N_39939,N_38758);
and U40656 (N_40656,N_38596,N_38529);
and U40657 (N_40657,N_39668,N_39913);
nor U40658 (N_40658,N_38231,N_39072);
or U40659 (N_40659,N_38288,N_39649);
xnor U40660 (N_40660,N_38921,N_39384);
xor U40661 (N_40661,N_39923,N_39419);
and U40662 (N_40662,N_38252,N_39619);
and U40663 (N_40663,N_39634,N_39378);
nand U40664 (N_40664,N_38355,N_39198);
nand U40665 (N_40665,N_39592,N_38018);
and U40666 (N_40666,N_38548,N_39369);
or U40667 (N_40667,N_39445,N_38168);
nand U40668 (N_40668,N_39282,N_39067);
xnor U40669 (N_40669,N_38087,N_39545);
nor U40670 (N_40670,N_39238,N_38188);
xnor U40671 (N_40671,N_38320,N_38926);
nor U40672 (N_40672,N_38793,N_38571);
xnor U40673 (N_40673,N_38122,N_39702);
nor U40674 (N_40674,N_39897,N_38432);
or U40675 (N_40675,N_39815,N_38593);
and U40676 (N_40676,N_39569,N_39012);
xnor U40677 (N_40677,N_38439,N_39358);
and U40678 (N_40678,N_39264,N_38447);
nor U40679 (N_40679,N_38284,N_38299);
or U40680 (N_40680,N_39611,N_38145);
xor U40681 (N_40681,N_39742,N_38170);
nand U40682 (N_40682,N_39615,N_38506);
and U40683 (N_40683,N_38958,N_38306);
or U40684 (N_40684,N_38251,N_39852);
nand U40685 (N_40685,N_38584,N_38061);
nand U40686 (N_40686,N_38362,N_38036);
and U40687 (N_40687,N_38156,N_38954);
or U40688 (N_40688,N_38933,N_38125);
nor U40689 (N_40689,N_39757,N_38719);
and U40690 (N_40690,N_39216,N_39018);
nand U40691 (N_40691,N_39984,N_38656);
nor U40692 (N_40692,N_38194,N_38618);
nor U40693 (N_40693,N_39298,N_39542);
or U40694 (N_40694,N_39297,N_39610);
or U40695 (N_40695,N_38989,N_38898);
and U40696 (N_40696,N_38174,N_38386);
xnor U40697 (N_40697,N_38331,N_39051);
nand U40698 (N_40698,N_39255,N_39145);
nor U40699 (N_40699,N_38290,N_39299);
xor U40700 (N_40700,N_38572,N_39172);
nor U40701 (N_40701,N_38303,N_39053);
nor U40702 (N_40702,N_39966,N_38464);
and U40703 (N_40703,N_39833,N_38408);
nand U40704 (N_40704,N_39504,N_38131);
xor U40705 (N_40705,N_38265,N_39283);
or U40706 (N_40706,N_39362,N_39428);
nor U40707 (N_40707,N_39609,N_39992);
xnor U40708 (N_40708,N_39276,N_39458);
and U40709 (N_40709,N_39996,N_38580);
nand U40710 (N_40710,N_39943,N_39754);
or U40711 (N_40711,N_39915,N_38567);
xnor U40712 (N_40712,N_38426,N_38732);
nor U40713 (N_40713,N_39017,N_39625);
or U40714 (N_40714,N_38630,N_39719);
nor U40715 (N_40715,N_38366,N_38636);
or U40716 (N_40716,N_39767,N_39809);
nor U40717 (N_40717,N_39813,N_39958);
xor U40718 (N_40718,N_39524,N_38030);
nor U40719 (N_40719,N_38319,N_38768);
or U40720 (N_40720,N_38922,N_38533);
nor U40721 (N_40721,N_39989,N_39741);
nand U40722 (N_40722,N_39178,N_38560);
nor U40723 (N_40723,N_39312,N_39802);
and U40724 (N_40724,N_38854,N_39840);
and U40725 (N_40725,N_38345,N_38967);
nor U40726 (N_40726,N_38067,N_38065);
and U40727 (N_40727,N_38790,N_38663);
xnor U40728 (N_40728,N_39525,N_39215);
or U40729 (N_40729,N_38015,N_38388);
and U40730 (N_40730,N_39228,N_39560);
and U40731 (N_40731,N_39964,N_39142);
xor U40732 (N_40732,N_39635,N_38021);
and U40733 (N_40733,N_39408,N_38755);
xnor U40734 (N_40734,N_39959,N_38109);
or U40735 (N_40735,N_39431,N_38263);
nor U40736 (N_40736,N_38100,N_39676);
and U40737 (N_40737,N_38661,N_39218);
nor U40738 (N_40738,N_39909,N_38597);
and U40739 (N_40739,N_38212,N_38716);
nor U40740 (N_40740,N_38484,N_38664);
xnor U40741 (N_40741,N_38708,N_39522);
or U40742 (N_40742,N_38271,N_38694);
nand U40743 (N_40743,N_39195,N_38833);
nor U40744 (N_40744,N_39985,N_38832);
and U40745 (N_40745,N_38483,N_39798);
nand U40746 (N_40746,N_38242,N_38077);
and U40747 (N_40747,N_39940,N_39390);
nand U40748 (N_40748,N_39027,N_39477);
or U40749 (N_40749,N_39336,N_38851);
xor U40750 (N_40750,N_39688,N_38052);
or U40751 (N_40751,N_38091,N_38261);
and U40752 (N_40752,N_39995,N_39119);
or U40753 (N_40753,N_39529,N_39772);
xnor U40754 (N_40754,N_39306,N_38081);
nor U40755 (N_40755,N_39787,N_38882);
or U40756 (N_40756,N_39820,N_39753);
or U40757 (N_40757,N_39247,N_38787);
nand U40758 (N_40758,N_39303,N_39814);
nor U40759 (N_40759,N_39518,N_39334);
and U40760 (N_40760,N_38877,N_39916);
nor U40761 (N_40761,N_38622,N_39396);
nand U40762 (N_40762,N_38947,N_39977);
or U40763 (N_40763,N_38551,N_38236);
nand U40764 (N_40764,N_38771,N_38991);
nor U40765 (N_40765,N_39240,N_39052);
and U40766 (N_40766,N_38013,N_39026);
nand U40767 (N_40767,N_39806,N_38988);
nand U40768 (N_40768,N_39747,N_38801);
nor U40769 (N_40769,N_38777,N_39175);
and U40770 (N_40770,N_38752,N_38004);
nor U40771 (N_40771,N_38232,N_39658);
and U40772 (N_40772,N_38352,N_39856);
nand U40773 (N_40773,N_38919,N_38323);
and U40774 (N_40774,N_38457,N_39584);
and U40775 (N_40775,N_39882,N_39286);
nor U40776 (N_40776,N_38410,N_38987);
and U40777 (N_40777,N_39211,N_38957);
nand U40778 (N_40778,N_38555,N_38779);
and U40779 (N_40779,N_39947,N_39088);
xnor U40780 (N_40780,N_38422,N_38387);
nor U40781 (N_40781,N_38175,N_39975);
or U40782 (N_40782,N_39501,N_38347);
nand U40783 (N_40783,N_39777,N_38997);
nand U40784 (N_40784,N_39361,N_38900);
and U40785 (N_40785,N_38503,N_38946);
nor U40786 (N_40786,N_39751,N_38417);
and U40787 (N_40787,N_39899,N_38891);
and U40788 (N_40788,N_39375,N_39415);
or U40789 (N_40789,N_38054,N_39543);
xnor U40790 (N_40790,N_38840,N_38835);
nor U40791 (N_40791,N_38666,N_39691);
nand U40792 (N_40792,N_39315,N_39921);
nand U40793 (N_40793,N_38418,N_38795);
or U40794 (N_40794,N_39281,N_39781);
and U40795 (N_40795,N_39320,N_39064);
xor U40796 (N_40796,N_39533,N_39204);
nor U40797 (N_40797,N_38308,N_38733);
nor U40798 (N_40798,N_39774,N_38842);
nand U40799 (N_40799,N_39047,N_39705);
and U40800 (N_40800,N_39376,N_39576);
or U40801 (N_40801,N_38662,N_39291);
nor U40802 (N_40802,N_39714,N_38294);
or U40803 (N_40803,N_39135,N_39900);
nand U40804 (N_40804,N_39125,N_38689);
xor U40805 (N_40805,N_39572,N_38176);
nor U40806 (N_40806,N_38180,N_39910);
or U40807 (N_40807,N_39083,N_38765);
nand U40808 (N_40808,N_39857,N_39903);
nand U40809 (N_40809,N_39999,N_38041);
or U40810 (N_40810,N_38010,N_38704);
nor U40811 (N_40811,N_38014,N_39054);
nor U40812 (N_40812,N_39554,N_39683);
and U40813 (N_40813,N_39626,N_39087);
or U40814 (N_40814,N_38928,N_39547);
or U40815 (N_40815,N_39190,N_38045);
nand U40816 (N_40816,N_38112,N_39960);
and U40817 (N_40817,N_39020,N_39782);
nor U40818 (N_40818,N_39181,N_38709);
and U40819 (N_40819,N_39858,N_38343);
nor U40820 (N_40820,N_38420,N_39162);
and U40821 (N_40821,N_38181,N_39103);
nand U40822 (N_40822,N_38927,N_39459);
and U40823 (N_40823,N_38090,N_39976);
nand U40824 (N_40824,N_39710,N_39071);
nor U40825 (N_40825,N_39886,N_39810);
xnor U40826 (N_40826,N_39242,N_39745);
and U40827 (N_40827,N_39192,N_39870);
or U40828 (N_40828,N_38486,N_38443);
or U40829 (N_40829,N_38688,N_38445);
nor U40830 (N_40830,N_38105,N_39633);
and U40831 (N_40831,N_39763,N_38641);
and U40832 (N_40832,N_39703,N_38718);
nor U40833 (N_40833,N_38837,N_39481);
xnor U40834 (N_40834,N_38183,N_38595);
xnor U40835 (N_40835,N_39169,N_39573);
nor U40836 (N_40836,N_39129,N_38351);
and U40837 (N_40837,N_38556,N_39941);
xnor U40838 (N_40838,N_38881,N_38550);
xnor U40839 (N_40839,N_38635,N_39614);
and U40840 (N_40840,N_38996,N_38440);
and U40841 (N_40841,N_38965,N_38828);
nand U40842 (N_40842,N_39401,N_38805);
xor U40843 (N_40843,N_38585,N_39697);
or U40844 (N_40844,N_39321,N_39583);
nor U40845 (N_40845,N_38757,N_39196);
xnor U40846 (N_40846,N_39040,N_39209);
xnor U40847 (N_40847,N_38412,N_38815);
nor U40848 (N_40848,N_38675,N_39127);
xor U40849 (N_40849,N_38453,N_39066);
xnor U40850 (N_40850,N_38920,N_39329);
and U40851 (N_40851,N_38358,N_39887);
nor U40852 (N_40852,N_38944,N_39914);
nand U40853 (N_40853,N_38416,N_38565);
or U40854 (N_40854,N_39147,N_39241);
nor U40855 (N_40855,N_38096,N_38574);
nor U40856 (N_40856,N_38083,N_38321);
or U40857 (N_40857,N_39945,N_38008);
or U40858 (N_40858,N_38552,N_38908);
and U40859 (N_40859,N_39351,N_39365);
xnor U40860 (N_40860,N_38032,N_39288);
and U40861 (N_40861,N_39019,N_39980);
xor U40862 (N_40862,N_39461,N_38817);
and U40863 (N_40863,N_39629,N_39177);
and U40864 (N_40864,N_39841,N_38481);
nor U40865 (N_40865,N_38402,N_38579);
xor U40866 (N_40866,N_39552,N_39403);
nor U40867 (N_40867,N_38424,N_38955);
xnor U40868 (N_40868,N_38482,N_38745);
and U40869 (N_40869,N_39761,N_39407);
xor U40870 (N_40870,N_38456,N_38295);
nand U40871 (N_40871,N_39186,N_38762);
xnor U40872 (N_40872,N_39728,N_39861);
nand U40873 (N_40873,N_39621,N_38260);
or U40874 (N_40874,N_39138,N_39516);
or U40875 (N_40875,N_39015,N_39076);
and U40876 (N_40876,N_39911,N_39568);
or U40877 (N_40877,N_38172,N_38460);
xor U40878 (N_40878,N_38458,N_38291);
or U40879 (N_40879,N_38073,N_38313);
xnor U40880 (N_40880,N_39313,N_38727);
nor U40881 (N_40881,N_39468,N_38609);
or U40882 (N_40882,N_38941,N_39271);
and U40883 (N_40883,N_39042,N_39492);
nand U40884 (N_40884,N_38224,N_39442);
and U40885 (N_40885,N_39426,N_39205);
xnor U40886 (N_40886,N_38099,N_38568);
and U40887 (N_40887,N_39652,N_39221);
xnor U40888 (N_40888,N_38207,N_39971);
nand U40889 (N_40889,N_39617,N_39210);
nor U40890 (N_40890,N_38296,N_38870);
or U40891 (N_40891,N_39457,N_39118);
and U40892 (N_40892,N_38213,N_38910);
nor U40893 (N_40893,N_39448,N_39997);
and U40894 (N_40894,N_39681,N_38863);
xnor U40895 (N_40895,N_39694,N_39270);
nor U40896 (N_40896,N_38673,N_39108);
and U40897 (N_40897,N_39983,N_39855);
and U40898 (N_40898,N_39739,N_38756);
nor U40899 (N_40899,N_39033,N_39990);
or U40900 (N_40900,N_39556,N_38273);
and U40901 (N_40901,N_39249,N_39293);
or U40902 (N_40902,N_38243,N_38918);
nor U40903 (N_40903,N_38182,N_39134);
nor U40904 (N_40904,N_38094,N_38205);
nand U40905 (N_40905,N_39309,N_38761);
nor U40906 (N_40906,N_38246,N_39164);
nor U40907 (N_40907,N_39764,N_38050);
and U40908 (N_40908,N_38522,N_38467);
xor U40909 (N_40909,N_38772,N_39708);
xor U40910 (N_40910,N_39454,N_39540);
nand U40911 (N_40911,N_38711,N_39385);
nor U40912 (N_40912,N_38728,N_39656);
and U40913 (N_40913,N_38076,N_39515);
or U40914 (N_40914,N_39770,N_39101);
and U40915 (N_40915,N_39391,N_38080);
and U40916 (N_40916,N_38009,N_38228);
or U40917 (N_40917,N_38292,N_39194);
or U40918 (N_40918,N_38000,N_39946);
nand U40919 (N_40919,N_39931,N_39140);
xnor U40920 (N_40920,N_38785,N_38185);
nor U40921 (N_40921,N_38135,N_39433);
or U40922 (N_40922,N_39927,N_39463);
nor U40923 (N_40923,N_38824,N_39684);
and U40924 (N_40924,N_38542,N_38309);
and U40925 (N_40925,N_39493,N_38262);
nor U40926 (N_40926,N_39338,N_38436);
or U40927 (N_40927,N_39207,N_39200);
nand U40928 (N_40928,N_39100,N_38604);
nand U40929 (N_40929,N_39685,N_39541);
nand U40930 (N_40930,N_38353,N_39588);
nand U40931 (N_40931,N_38489,N_39132);
xor U40932 (N_40932,N_39347,N_39302);
xor U40933 (N_40933,N_38830,N_39759);
or U40934 (N_40934,N_38124,N_39864);
nand U40935 (N_40935,N_38346,N_38696);
or U40936 (N_40936,N_38705,N_38715);
xnor U40937 (N_40937,N_39141,N_39355);
xnor U40938 (N_40938,N_38809,N_38129);
or U40939 (N_40939,N_39070,N_39257);
nand U40940 (N_40940,N_38894,N_39167);
nor U40941 (N_40941,N_38575,N_39352);
xor U40942 (N_40942,N_38679,N_38127);
nor U40943 (N_40943,N_38005,N_38692);
xor U40944 (N_40944,N_38808,N_39828);
or U40945 (N_40945,N_38155,N_38312);
xor U40946 (N_40946,N_38391,N_39842);
nand U40947 (N_40947,N_39174,N_38825);
nor U40948 (N_40948,N_39585,N_38419);
xnor U40949 (N_40949,N_38060,N_38654);
or U40950 (N_40950,N_39425,N_38526);
nor U40951 (N_40951,N_38890,N_39202);
nand U40952 (N_40952,N_38897,N_38826);
xor U40953 (N_40953,N_38048,N_38187);
nor U40954 (N_40954,N_39024,N_38059);
or U40955 (N_40955,N_38349,N_38523);
nand U40956 (N_40956,N_39788,N_39987);
and U40957 (N_40957,N_39116,N_39531);
and U40958 (N_40958,N_38214,N_39084);
nor U40959 (N_40959,N_39121,N_38866);
nor U40960 (N_40960,N_39638,N_38020);
nor U40961 (N_40961,N_39526,N_38179);
nand U40962 (N_40962,N_38370,N_39808);
nor U40963 (N_40963,N_38385,N_39265);
xnor U40964 (N_40964,N_39094,N_38327);
nand U40965 (N_40965,N_38710,N_39002);
and U40966 (N_40966,N_38725,N_39296);
and U40967 (N_40967,N_38536,N_38171);
nor U40968 (N_40968,N_39474,N_38665);
nand U40969 (N_40969,N_39785,N_39050);
nor U40970 (N_40970,N_39586,N_39796);
nor U40971 (N_40971,N_38204,N_38304);
or U40972 (N_40972,N_39038,N_39948);
nor U40973 (N_40973,N_38626,N_38827);
xor U40974 (N_40974,N_38459,N_38139);
or U40975 (N_40975,N_38435,N_38003);
nor U40976 (N_40976,N_38695,N_39651);
xor U40977 (N_40977,N_39979,N_38616);
or U40978 (N_40978,N_38802,N_38737);
nand U40979 (N_40979,N_38249,N_38230);
xor U40980 (N_40980,N_38082,N_39465);
and U40981 (N_40981,N_38717,N_39011);
xor U40982 (N_40982,N_38203,N_38448);
and U40983 (N_40983,N_39575,N_39266);
and U40984 (N_40984,N_38473,N_39082);
xnor U40985 (N_40985,N_38088,N_38993);
xor U40986 (N_40986,N_39661,N_39643);
nor U40987 (N_40987,N_38586,N_38823);
xnor U40988 (N_40988,N_39451,N_39486);
nand U40989 (N_40989,N_39883,N_39920);
or U40990 (N_40990,N_39623,N_39830);
nand U40991 (N_40991,N_39846,N_38365);
and U40992 (N_40992,N_39009,N_38229);
xnor U40993 (N_40993,N_38475,N_38404);
xor U40994 (N_40994,N_38598,N_39004);
nand U40995 (N_40995,N_38093,N_38549);
nand U40996 (N_40996,N_39607,N_39122);
xnor U40997 (N_40997,N_38573,N_39435);
and U40998 (N_40998,N_39839,N_38423);
and U40999 (N_40999,N_38748,N_38563);
xnor U41000 (N_41000,N_38086,N_38455);
or U41001 (N_41001,N_38776,N_39802);
and U41002 (N_41002,N_38247,N_39942);
xor U41003 (N_41003,N_38411,N_39448);
and U41004 (N_41004,N_39651,N_38083);
or U41005 (N_41005,N_39530,N_38917);
nor U41006 (N_41006,N_39458,N_39047);
and U41007 (N_41007,N_38577,N_39829);
nand U41008 (N_41008,N_39442,N_39526);
or U41009 (N_41009,N_39990,N_39386);
or U41010 (N_41010,N_38624,N_38490);
xnor U41011 (N_41011,N_38539,N_39761);
xnor U41012 (N_41012,N_38909,N_38499);
or U41013 (N_41013,N_38431,N_39877);
nor U41014 (N_41014,N_38508,N_39950);
xor U41015 (N_41015,N_38298,N_39348);
nand U41016 (N_41016,N_38474,N_39873);
xnor U41017 (N_41017,N_38726,N_38560);
and U41018 (N_41018,N_38641,N_38636);
xor U41019 (N_41019,N_38104,N_38774);
nand U41020 (N_41020,N_38718,N_39141);
nand U41021 (N_41021,N_38371,N_39476);
or U41022 (N_41022,N_39436,N_38803);
nor U41023 (N_41023,N_38258,N_38699);
and U41024 (N_41024,N_38733,N_39653);
xor U41025 (N_41025,N_39751,N_39516);
and U41026 (N_41026,N_38287,N_38061);
xor U41027 (N_41027,N_38236,N_38129);
and U41028 (N_41028,N_38014,N_39675);
xnor U41029 (N_41029,N_39621,N_39691);
xor U41030 (N_41030,N_39830,N_38420);
nor U41031 (N_41031,N_38041,N_38160);
xor U41032 (N_41032,N_38495,N_38467);
nand U41033 (N_41033,N_38352,N_39140);
or U41034 (N_41034,N_38181,N_38786);
xnor U41035 (N_41035,N_39678,N_38957);
xor U41036 (N_41036,N_39856,N_38883);
nor U41037 (N_41037,N_39450,N_38101);
or U41038 (N_41038,N_38175,N_38846);
nor U41039 (N_41039,N_38934,N_39649);
or U41040 (N_41040,N_38475,N_38804);
nand U41041 (N_41041,N_39654,N_38164);
or U41042 (N_41042,N_38758,N_38843);
nand U41043 (N_41043,N_39600,N_38088);
and U41044 (N_41044,N_38609,N_38804);
nor U41045 (N_41045,N_38559,N_38703);
or U41046 (N_41046,N_39513,N_38607);
and U41047 (N_41047,N_38264,N_39826);
xor U41048 (N_41048,N_39186,N_39429);
and U41049 (N_41049,N_38502,N_38803);
nand U41050 (N_41050,N_39807,N_38345);
xnor U41051 (N_41051,N_38121,N_39381);
or U41052 (N_41052,N_39620,N_38822);
and U41053 (N_41053,N_38294,N_39131);
xor U41054 (N_41054,N_38646,N_38345);
nand U41055 (N_41055,N_38206,N_38740);
nand U41056 (N_41056,N_39200,N_39760);
nor U41057 (N_41057,N_39854,N_39255);
or U41058 (N_41058,N_38373,N_39161);
nand U41059 (N_41059,N_38961,N_39159);
or U41060 (N_41060,N_38382,N_39650);
nand U41061 (N_41061,N_38540,N_38689);
nor U41062 (N_41062,N_39953,N_38101);
or U41063 (N_41063,N_38557,N_39427);
nand U41064 (N_41064,N_39050,N_38919);
nor U41065 (N_41065,N_39172,N_39389);
and U41066 (N_41066,N_38318,N_38358);
and U41067 (N_41067,N_38240,N_39737);
nor U41068 (N_41068,N_39787,N_39728);
nand U41069 (N_41069,N_38201,N_38718);
nor U41070 (N_41070,N_38123,N_39039);
or U41071 (N_41071,N_38805,N_39665);
xor U41072 (N_41072,N_39122,N_39367);
nor U41073 (N_41073,N_38998,N_38640);
or U41074 (N_41074,N_39094,N_38625);
nor U41075 (N_41075,N_38975,N_38522);
and U41076 (N_41076,N_38024,N_39616);
xnor U41077 (N_41077,N_39437,N_39724);
nor U41078 (N_41078,N_39825,N_38961);
nand U41079 (N_41079,N_39656,N_38310);
nand U41080 (N_41080,N_38608,N_38450);
or U41081 (N_41081,N_38218,N_39830);
and U41082 (N_41082,N_39262,N_39489);
nand U41083 (N_41083,N_39246,N_39320);
nor U41084 (N_41084,N_39209,N_38406);
or U41085 (N_41085,N_39546,N_39357);
nand U41086 (N_41086,N_39682,N_38997);
or U41087 (N_41087,N_38281,N_38300);
or U41088 (N_41088,N_38906,N_38747);
and U41089 (N_41089,N_38117,N_38587);
and U41090 (N_41090,N_38670,N_38164);
nor U41091 (N_41091,N_38728,N_38731);
nor U41092 (N_41092,N_38961,N_38294);
nand U41093 (N_41093,N_38333,N_39999);
nor U41094 (N_41094,N_39793,N_39020);
and U41095 (N_41095,N_39886,N_38122);
nor U41096 (N_41096,N_39973,N_39750);
or U41097 (N_41097,N_38788,N_38536);
nor U41098 (N_41098,N_38824,N_39530);
nand U41099 (N_41099,N_38895,N_39296);
nand U41100 (N_41100,N_39195,N_38830);
and U41101 (N_41101,N_38026,N_39067);
or U41102 (N_41102,N_39705,N_38839);
or U41103 (N_41103,N_39732,N_39640);
nand U41104 (N_41104,N_38715,N_38637);
xor U41105 (N_41105,N_39375,N_39007);
nor U41106 (N_41106,N_38416,N_38928);
xor U41107 (N_41107,N_39055,N_38199);
and U41108 (N_41108,N_39495,N_38722);
or U41109 (N_41109,N_38217,N_38335);
and U41110 (N_41110,N_38165,N_39268);
nand U41111 (N_41111,N_39408,N_38852);
and U41112 (N_41112,N_38416,N_38142);
and U41113 (N_41113,N_38763,N_38427);
xnor U41114 (N_41114,N_39529,N_38879);
nand U41115 (N_41115,N_38055,N_38382);
nor U41116 (N_41116,N_39672,N_38765);
nor U41117 (N_41117,N_39078,N_39559);
xnor U41118 (N_41118,N_38444,N_38895);
and U41119 (N_41119,N_39132,N_38622);
nor U41120 (N_41120,N_38125,N_39744);
and U41121 (N_41121,N_39713,N_39455);
and U41122 (N_41122,N_38582,N_38303);
nor U41123 (N_41123,N_38730,N_38638);
and U41124 (N_41124,N_39611,N_39069);
nor U41125 (N_41125,N_38632,N_38977);
and U41126 (N_41126,N_38603,N_38845);
or U41127 (N_41127,N_38651,N_39591);
nand U41128 (N_41128,N_38539,N_38992);
nor U41129 (N_41129,N_39723,N_38216);
or U41130 (N_41130,N_39371,N_39907);
nor U41131 (N_41131,N_39774,N_39020);
nor U41132 (N_41132,N_39845,N_39222);
xor U41133 (N_41133,N_38245,N_39467);
nor U41134 (N_41134,N_38573,N_39495);
and U41135 (N_41135,N_38736,N_38892);
xnor U41136 (N_41136,N_38454,N_39773);
or U41137 (N_41137,N_38939,N_38837);
nor U41138 (N_41138,N_39534,N_38243);
xnor U41139 (N_41139,N_38052,N_39884);
nor U41140 (N_41140,N_38717,N_38073);
nor U41141 (N_41141,N_38231,N_38612);
and U41142 (N_41142,N_39092,N_39419);
or U41143 (N_41143,N_38167,N_39037);
nor U41144 (N_41144,N_39817,N_39928);
and U41145 (N_41145,N_39818,N_39037);
xnor U41146 (N_41146,N_38009,N_39468);
nor U41147 (N_41147,N_38960,N_39139);
or U41148 (N_41148,N_38304,N_39976);
nand U41149 (N_41149,N_39613,N_38327);
and U41150 (N_41150,N_39119,N_38913);
and U41151 (N_41151,N_38290,N_39777);
or U41152 (N_41152,N_38262,N_39263);
and U41153 (N_41153,N_38120,N_38429);
nand U41154 (N_41154,N_39157,N_39748);
nand U41155 (N_41155,N_39239,N_38292);
and U41156 (N_41156,N_38565,N_38832);
xnor U41157 (N_41157,N_38309,N_39074);
and U41158 (N_41158,N_38150,N_39836);
xnor U41159 (N_41159,N_38446,N_38187);
and U41160 (N_41160,N_39220,N_39576);
or U41161 (N_41161,N_38927,N_38707);
or U41162 (N_41162,N_39082,N_38144);
or U41163 (N_41163,N_39230,N_38179);
xnor U41164 (N_41164,N_39082,N_39064);
xnor U41165 (N_41165,N_39808,N_39666);
or U41166 (N_41166,N_39596,N_38489);
nor U41167 (N_41167,N_38825,N_39872);
xnor U41168 (N_41168,N_39370,N_38077);
or U41169 (N_41169,N_39022,N_38734);
or U41170 (N_41170,N_39886,N_38659);
and U41171 (N_41171,N_38058,N_39109);
and U41172 (N_41172,N_38142,N_38841);
xnor U41173 (N_41173,N_38426,N_39370);
or U41174 (N_41174,N_38711,N_39370);
xor U41175 (N_41175,N_39784,N_39003);
or U41176 (N_41176,N_39884,N_38668);
nand U41177 (N_41177,N_39035,N_38741);
nor U41178 (N_41178,N_39355,N_39291);
nand U41179 (N_41179,N_39256,N_39731);
or U41180 (N_41180,N_39356,N_39389);
nand U41181 (N_41181,N_38387,N_38053);
nand U41182 (N_41182,N_39876,N_39854);
nor U41183 (N_41183,N_38701,N_38939);
xnor U41184 (N_41184,N_38957,N_38953);
or U41185 (N_41185,N_39027,N_38613);
and U41186 (N_41186,N_38700,N_39747);
nor U41187 (N_41187,N_39079,N_38034);
nand U41188 (N_41188,N_38140,N_39458);
or U41189 (N_41189,N_39448,N_39820);
nand U41190 (N_41190,N_38369,N_38890);
or U41191 (N_41191,N_38396,N_39575);
nor U41192 (N_41192,N_39493,N_38384);
or U41193 (N_41193,N_38548,N_38250);
nor U41194 (N_41194,N_38514,N_38587);
xor U41195 (N_41195,N_39381,N_38531);
and U41196 (N_41196,N_38992,N_38185);
nand U41197 (N_41197,N_38707,N_39097);
nor U41198 (N_41198,N_39263,N_38324);
nand U41199 (N_41199,N_38155,N_39907);
and U41200 (N_41200,N_38005,N_39186);
xnor U41201 (N_41201,N_38742,N_39179);
and U41202 (N_41202,N_38136,N_38671);
nor U41203 (N_41203,N_39409,N_38317);
and U41204 (N_41204,N_38199,N_38279);
or U41205 (N_41205,N_38269,N_38425);
and U41206 (N_41206,N_38113,N_38808);
nand U41207 (N_41207,N_39700,N_39825);
xor U41208 (N_41208,N_38673,N_38857);
nand U41209 (N_41209,N_38937,N_39746);
and U41210 (N_41210,N_39810,N_39076);
nor U41211 (N_41211,N_39163,N_39125);
or U41212 (N_41212,N_39193,N_39709);
or U41213 (N_41213,N_38315,N_38087);
nand U41214 (N_41214,N_38112,N_39814);
and U41215 (N_41215,N_38353,N_38549);
or U41216 (N_41216,N_39724,N_39985);
xor U41217 (N_41217,N_39656,N_38820);
and U41218 (N_41218,N_38962,N_39399);
or U41219 (N_41219,N_38969,N_39688);
nand U41220 (N_41220,N_38178,N_38338);
xnor U41221 (N_41221,N_38522,N_39192);
and U41222 (N_41222,N_39967,N_38456);
xnor U41223 (N_41223,N_38931,N_39318);
nor U41224 (N_41224,N_39457,N_38422);
nand U41225 (N_41225,N_38336,N_39246);
nor U41226 (N_41226,N_38299,N_39689);
and U41227 (N_41227,N_39447,N_38036);
or U41228 (N_41228,N_39838,N_39720);
and U41229 (N_41229,N_39365,N_38557);
and U41230 (N_41230,N_38380,N_39884);
and U41231 (N_41231,N_39309,N_39438);
and U41232 (N_41232,N_39993,N_39581);
xnor U41233 (N_41233,N_39772,N_38992);
xor U41234 (N_41234,N_38942,N_38755);
xnor U41235 (N_41235,N_38218,N_38986);
and U41236 (N_41236,N_38224,N_38225);
nand U41237 (N_41237,N_39617,N_38279);
xnor U41238 (N_41238,N_38877,N_39248);
and U41239 (N_41239,N_39651,N_39363);
nor U41240 (N_41240,N_38764,N_38402);
nor U41241 (N_41241,N_39416,N_38615);
and U41242 (N_41242,N_38614,N_39489);
and U41243 (N_41243,N_39910,N_39883);
nand U41244 (N_41244,N_38319,N_38460);
nor U41245 (N_41245,N_39266,N_38870);
nor U41246 (N_41246,N_38512,N_38173);
nor U41247 (N_41247,N_39654,N_39834);
nor U41248 (N_41248,N_39525,N_38346);
or U41249 (N_41249,N_38676,N_39053);
nor U41250 (N_41250,N_38664,N_39392);
or U41251 (N_41251,N_39185,N_39689);
nor U41252 (N_41252,N_39508,N_38379);
and U41253 (N_41253,N_39430,N_39537);
xnor U41254 (N_41254,N_39542,N_39639);
nand U41255 (N_41255,N_39098,N_39386);
xor U41256 (N_41256,N_38491,N_38261);
xor U41257 (N_41257,N_38619,N_39208);
nor U41258 (N_41258,N_39117,N_39409);
or U41259 (N_41259,N_39204,N_39452);
or U41260 (N_41260,N_38627,N_38775);
xnor U41261 (N_41261,N_38669,N_39710);
xnor U41262 (N_41262,N_39114,N_39419);
or U41263 (N_41263,N_39640,N_38455);
and U41264 (N_41264,N_39557,N_38211);
and U41265 (N_41265,N_39414,N_38495);
nand U41266 (N_41266,N_38805,N_38175);
and U41267 (N_41267,N_38881,N_38803);
and U41268 (N_41268,N_39853,N_38463);
nand U41269 (N_41269,N_38529,N_39877);
xor U41270 (N_41270,N_38805,N_38661);
or U41271 (N_41271,N_39055,N_38997);
nand U41272 (N_41272,N_39166,N_39316);
or U41273 (N_41273,N_39881,N_38900);
nor U41274 (N_41274,N_39195,N_39016);
xnor U41275 (N_41275,N_38417,N_38394);
nor U41276 (N_41276,N_38177,N_38765);
nand U41277 (N_41277,N_39293,N_39153);
nor U41278 (N_41278,N_38232,N_39150);
and U41279 (N_41279,N_38993,N_39810);
and U41280 (N_41280,N_38378,N_39780);
and U41281 (N_41281,N_39658,N_38117);
or U41282 (N_41282,N_38625,N_39373);
nor U41283 (N_41283,N_38106,N_38525);
nor U41284 (N_41284,N_39486,N_39106);
xor U41285 (N_41285,N_39158,N_38993);
or U41286 (N_41286,N_38295,N_38985);
or U41287 (N_41287,N_38070,N_39718);
and U41288 (N_41288,N_38321,N_39541);
and U41289 (N_41289,N_39969,N_38035);
and U41290 (N_41290,N_38547,N_38500);
nor U41291 (N_41291,N_39995,N_38888);
xnor U41292 (N_41292,N_38842,N_38682);
or U41293 (N_41293,N_38826,N_38238);
or U41294 (N_41294,N_38497,N_39948);
xor U41295 (N_41295,N_38823,N_39296);
xnor U41296 (N_41296,N_39919,N_39154);
and U41297 (N_41297,N_38359,N_39364);
xor U41298 (N_41298,N_39423,N_38220);
nand U41299 (N_41299,N_39795,N_38321);
or U41300 (N_41300,N_38552,N_38255);
or U41301 (N_41301,N_39888,N_39151);
nor U41302 (N_41302,N_38426,N_39758);
nor U41303 (N_41303,N_38113,N_39259);
nand U41304 (N_41304,N_38878,N_39035);
or U41305 (N_41305,N_38273,N_39290);
xor U41306 (N_41306,N_38062,N_39382);
nor U41307 (N_41307,N_39414,N_38887);
nand U41308 (N_41308,N_38697,N_39868);
nor U41309 (N_41309,N_39471,N_39135);
xnor U41310 (N_41310,N_38741,N_39998);
nor U41311 (N_41311,N_38687,N_38135);
xnor U41312 (N_41312,N_38113,N_39960);
nand U41313 (N_41313,N_38717,N_39336);
and U41314 (N_41314,N_38731,N_39920);
and U41315 (N_41315,N_38565,N_39329);
and U41316 (N_41316,N_39277,N_38609);
xnor U41317 (N_41317,N_39152,N_38042);
nor U41318 (N_41318,N_38514,N_39285);
nand U41319 (N_41319,N_38693,N_39264);
nand U41320 (N_41320,N_39091,N_38207);
or U41321 (N_41321,N_38291,N_38852);
nor U41322 (N_41322,N_38153,N_38610);
nor U41323 (N_41323,N_38764,N_39738);
nor U41324 (N_41324,N_39275,N_38206);
nand U41325 (N_41325,N_38880,N_38428);
or U41326 (N_41326,N_38513,N_39868);
xnor U41327 (N_41327,N_39128,N_39992);
xor U41328 (N_41328,N_39025,N_38239);
xor U41329 (N_41329,N_39016,N_39344);
nor U41330 (N_41330,N_39909,N_39634);
nand U41331 (N_41331,N_39319,N_39088);
or U41332 (N_41332,N_39085,N_39484);
and U41333 (N_41333,N_38351,N_39676);
or U41334 (N_41334,N_38470,N_39898);
xnor U41335 (N_41335,N_39925,N_39174);
xor U41336 (N_41336,N_38666,N_39932);
nand U41337 (N_41337,N_39344,N_39392);
or U41338 (N_41338,N_38175,N_38747);
xnor U41339 (N_41339,N_39973,N_38261);
xnor U41340 (N_41340,N_38917,N_39284);
and U41341 (N_41341,N_39915,N_38768);
xor U41342 (N_41342,N_38305,N_39127);
or U41343 (N_41343,N_38628,N_38418);
nand U41344 (N_41344,N_38481,N_39058);
or U41345 (N_41345,N_38153,N_39828);
xor U41346 (N_41346,N_38184,N_38253);
nand U41347 (N_41347,N_38065,N_38159);
and U41348 (N_41348,N_38731,N_38448);
nor U41349 (N_41349,N_39184,N_38900);
or U41350 (N_41350,N_39155,N_38201);
nand U41351 (N_41351,N_38881,N_39631);
and U41352 (N_41352,N_38587,N_38627);
or U41353 (N_41353,N_39638,N_39111);
nand U41354 (N_41354,N_38007,N_39510);
or U41355 (N_41355,N_38527,N_38630);
xnor U41356 (N_41356,N_39539,N_38003);
or U41357 (N_41357,N_39875,N_39765);
xnor U41358 (N_41358,N_39365,N_39003);
nor U41359 (N_41359,N_39759,N_39150);
nor U41360 (N_41360,N_38197,N_38676);
or U41361 (N_41361,N_38772,N_38036);
xnor U41362 (N_41362,N_38463,N_38022);
or U41363 (N_41363,N_38526,N_38396);
xor U41364 (N_41364,N_39451,N_39664);
and U41365 (N_41365,N_39278,N_39397);
xnor U41366 (N_41366,N_38899,N_38441);
nand U41367 (N_41367,N_39777,N_38085);
or U41368 (N_41368,N_39215,N_39961);
nor U41369 (N_41369,N_38378,N_38540);
nor U41370 (N_41370,N_38754,N_38909);
nand U41371 (N_41371,N_39082,N_39173);
or U41372 (N_41372,N_38810,N_38699);
and U41373 (N_41373,N_38551,N_38629);
and U41374 (N_41374,N_38014,N_39548);
nand U41375 (N_41375,N_38221,N_39037);
nand U41376 (N_41376,N_38713,N_39265);
xor U41377 (N_41377,N_39177,N_38962);
xor U41378 (N_41378,N_39765,N_39323);
xnor U41379 (N_41379,N_39765,N_38105);
xor U41380 (N_41380,N_38063,N_39775);
or U41381 (N_41381,N_39509,N_38523);
nand U41382 (N_41382,N_38313,N_39331);
and U41383 (N_41383,N_38481,N_39332);
or U41384 (N_41384,N_39862,N_38222);
xor U41385 (N_41385,N_39003,N_38105);
nand U41386 (N_41386,N_38130,N_38897);
or U41387 (N_41387,N_38661,N_38413);
nand U41388 (N_41388,N_38863,N_38781);
and U41389 (N_41389,N_38775,N_38237);
and U41390 (N_41390,N_39011,N_39464);
nor U41391 (N_41391,N_38727,N_38306);
nand U41392 (N_41392,N_39860,N_39394);
or U41393 (N_41393,N_38786,N_38794);
nand U41394 (N_41394,N_38848,N_39165);
or U41395 (N_41395,N_39288,N_38424);
nand U41396 (N_41396,N_39089,N_39513);
xor U41397 (N_41397,N_39664,N_38428);
xor U41398 (N_41398,N_38153,N_39677);
and U41399 (N_41399,N_38079,N_39998);
or U41400 (N_41400,N_39670,N_38472);
and U41401 (N_41401,N_39677,N_38778);
nor U41402 (N_41402,N_38059,N_39516);
or U41403 (N_41403,N_38995,N_39108);
and U41404 (N_41404,N_38702,N_39696);
nor U41405 (N_41405,N_38649,N_39191);
and U41406 (N_41406,N_38153,N_38770);
nor U41407 (N_41407,N_38155,N_38246);
and U41408 (N_41408,N_38179,N_39486);
or U41409 (N_41409,N_39714,N_39485);
and U41410 (N_41410,N_39606,N_39574);
xnor U41411 (N_41411,N_38501,N_39567);
nor U41412 (N_41412,N_38517,N_38749);
xnor U41413 (N_41413,N_38784,N_39439);
and U41414 (N_41414,N_39253,N_39335);
xor U41415 (N_41415,N_38999,N_38695);
nand U41416 (N_41416,N_39152,N_39100);
nand U41417 (N_41417,N_39394,N_38635);
xor U41418 (N_41418,N_39940,N_39699);
and U41419 (N_41419,N_39073,N_38391);
xor U41420 (N_41420,N_39041,N_38551);
or U41421 (N_41421,N_39954,N_38011);
and U41422 (N_41422,N_39149,N_38523);
or U41423 (N_41423,N_38406,N_39614);
and U41424 (N_41424,N_39853,N_38012);
nor U41425 (N_41425,N_38615,N_38127);
nand U41426 (N_41426,N_39535,N_39522);
xnor U41427 (N_41427,N_38436,N_38473);
xor U41428 (N_41428,N_39157,N_39177);
and U41429 (N_41429,N_39761,N_39236);
xnor U41430 (N_41430,N_39120,N_39275);
xnor U41431 (N_41431,N_39044,N_38936);
nor U41432 (N_41432,N_39571,N_39390);
nand U41433 (N_41433,N_39342,N_38571);
xnor U41434 (N_41434,N_39539,N_39118);
xnor U41435 (N_41435,N_39491,N_38237);
or U41436 (N_41436,N_38227,N_39574);
nand U41437 (N_41437,N_38780,N_39428);
and U41438 (N_41438,N_38109,N_38189);
nor U41439 (N_41439,N_39093,N_38232);
nor U41440 (N_41440,N_38650,N_39877);
nor U41441 (N_41441,N_39509,N_38696);
or U41442 (N_41442,N_38482,N_39712);
nor U41443 (N_41443,N_38734,N_39696);
xor U41444 (N_41444,N_39800,N_39855);
nand U41445 (N_41445,N_39815,N_39245);
or U41446 (N_41446,N_39396,N_39576);
nor U41447 (N_41447,N_38045,N_38911);
or U41448 (N_41448,N_39645,N_39629);
nand U41449 (N_41449,N_38348,N_39472);
and U41450 (N_41450,N_39548,N_38605);
nand U41451 (N_41451,N_39039,N_39292);
nor U41452 (N_41452,N_38475,N_38930);
or U41453 (N_41453,N_38658,N_39112);
and U41454 (N_41454,N_38378,N_39144);
or U41455 (N_41455,N_39865,N_39760);
xor U41456 (N_41456,N_39445,N_39968);
xnor U41457 (N_41457,N_38181,N_39583);
nand U41458 (N_41458,N_38860,N_39534);
nand U41459 (N_41459,N_38573,N_38158);
and U41460 (N_41460,N_38396,N_38727);
xor U41461 (N_41461,N_38916,N_39158);
and U41462 (N_41462,N_39426,N_38902);
nor U41463 (N_41463,N_39109,N_39480);
or U41464 (N_41464,N_38292,N_39501);
or U41465 (N_41465,N_38220,N_38903);
and U41466 (N_41466,N_38147,N_39538);
or U41467 (N_41467,N_38512,N_39614);
nor U41468 (N_41468,N_38134,N_38961);
nand U41469 (N_41469,N_39713,N_39847);
and U41470 (N_41470,N_39155,N_39973);
or U41471 (N_41471,N_39639,N_38677);
and U41472 (N_41472,N_38879,N_38298);
xor U41473 (N_41473,N_38597,N_38695);
or U41474 (N_41474,N_39170,N_38443);
or U41475 (N_41475,N_39549,N_39170);
nand U41476 (N_41476,N_39233,N_39088);
nor U41477 (N_41477,N_38782,N_38867);
nor U41478 (N_41478,N_39468,N_39180);
or U41479 (N_41479,N_38067,N_39581);
nor U41480 (N_41480,N_38946,N_39834);
nor U41481 (N_41481,N_38529,N_39386);
nor U41482 (N_41482,N_39687,N_39455);
nor U41483 (N_41483,N_39663,N_38063);
nor U41484 (N_41484,N_38330,N_39931);
nor U41485 (N_41485,N_39224,N_38279);
or U41486 (N_41486,N_39131,N_39302);
nor U41487 (N_41487,N_39238,N_39327);
nand U41488 (N_41488,N_39879,N_39004);
or U41489 (N_41489,N_39280,N_39083);
or U41490 (N_41490,N_39354,N_38088);
nand U41491 (N_41491,N_39958,N_38081);
or U41492 (N_41492,N_38483,N_39440);
nor U41493 (N_41493,N_39620,N_39143);
xnor U41494 (N_41494,N_39964,N_39971);
and U41495 (N_41495,N_39335,N_39057);
xor U41496 (N_41496,N_39916,N_39920);
or U41497 (N_41497,N_39667,N_38640);
nor U41498 (N_41498,N_38408,N_38949);
and U41499 (N_41499,N_39136,N_39301);
nand U41500 (N_41500,N_38549,N_39076);
or U41501 (N_41501,N_39631,N_39131);
or U41502 (N_41502,N_38558,N_38696);
and U41503 (N_41503,N_38825,N_38466);
and U41504 (N_41504,N_39929,N_39077);
nor U41505 (N_41505,N_38316,N_38242);
xnor U41506 (N_41506,N_38042,N_39026);
or U41507 (N_41507,N_39300,N_38526);
nand U41508 (N_41508,N_39050,N_39721);
or U41509 (N_41509,N_38372,N_38783);
nor U41510 (N_41510,N_38504,N_39014);
nor U41511 (N_41511,N_38812,N_39959);
nand U41512 (N_41512,N_38872,N_38148);
nor U41513 (N_41513,N_38367,N_38731);
or U41514 (N_41514,N_39458,N_39497);
nor U41515 (N_41515,N_38497,N_38409);
or U41516 (N_41516,N_38627,N_39310);
or U41517 (N_41517,N_38301,N_38679);
nor U41518 (N_41518,N_38092,N_38334);
nand U41519 (N_41519,N_38754,N_38367);
nor U41520 (N_41520,N_38900,N_39930);
nand U41521 (N_41521,N_38792,N_39233);
and U41522 (N_41522,N_39822,N_39793);
or U41523 (N_41523,N_39932,N_38471);
nand U41524 (N_41524,N_38132,N_38776);
xnor U41525 (N_41525,N_38592,N_38383);
and U41526 (N_41526,N_38569,N_39682);
or U41527 (N_41527,N_38442,N_39047);
or U41528 (N_41528,N_38196,N_38566);
nor U41529 (N_41529,N_38603,N_38901);
xnor U41530 (N_41530,N_38003,N_38771);
xnor U41531 (N_41531,N_38213,N_39595);
or U41532 (N_41532,N_38452,N_38877);
xor U41533 (N_41533,N_39613,N_39868);
and U41534 (N_41534,N_39167,N_38842);
and U41535 (N_41535,N_39631,N_38154);
and U41536 (N_41536,N_38363,N_39760);
xor U41537 (N_41537,N_38058,N_38229);
xor U41538 (N_41538,N_39600,N_39154);
or U41539 (N_41539,N_38529,N_38309);
nor U41540 (N_41540,N_39955,N_39996);
nor U41541 (N_41541,N_39313,N_38965);
nand U41542 (N_41542,N_39078,N_39964);
nor U41543 (N_41543,N_38532,N_39559);
nor U41544 (N_41544,N_38410,N_39995);
or U41545 (N_41545,N_39235,N_39899);
nor U41546 (N_41546,N_39478,N_38144);
or U41547 (N_41547,N_38309,N_38249);
nor U41548 (N_41548,N_39438,N_38095);
nand U41549 (N_41549,N_38690,N_38554);
nor U41550 (N_41550,N_38107,N_38689);
or U41551 (N_41551,N_39730,N_39439);
nor U41552 (N_41552,N_39169,N_38712);
nand U41553 (N_41553,N_39672,N_38230);
nand U41554 (N_41554,N_39514,N_39299);
nand U41555 (N_41555,N_38635,N_38393);
xnor U41556 (N_41556,N_38972,N_39723);
xor U41557 (N_41557,N_38039,N_38508);
nand U41558 (N_41558,N_38115,N_38748);
nand U41559 (N_41559,N_38298,N_39485);
nor U41560 (N_41560,N_38606,N_38013);
nor U41561 (N_41561,N_38050,N_38462);
nand U41562 (N_41562,N_38746,N_39344);
xor U41563 (N_41563,N_38120,N_38013);
and U41564 (N_41564,N_39200,N_38814);
nor U41565 (N_41565,N_38630,N_38468);
xnor U41566 (N_41566,N_38249,N_39262);
nor U41567 (N_41567,N_39803,N_39849);
xnor U41568 (N_41568,N_38764,N_38912);
and U41569 (N_41569,N_38551,N_38305);
and U41570 (N_41570,N_39356,N_38673);
and U41571 (N_41571,N_38704,N_38398);
nand U41572 (N_41572,N_39485,N_38829);
and U41573 (N_41573,N_38144,N_38287);
nand U41574 (N_41574,N_38095,N_39293);
xor U41575 (N_41575,N_38074,N_38354);
nor U41576 (N_41576,N_39851,N_38124);
nand U41577 (N_41577,N_38799,N_39815);
nor U41578 (N_41578,N_38746,N_38397);
xnor U41579 (N_41579,N_38217,N_38056);
and U41580 (N_41580,N_38795,N_38241);
xnor U41581 (N_41581,N_39685,N_39225);
and U41582 (N_41582,N_38722,N_39367);
nor U41583 (N_41583,N_39109,N_38381);
nor U41584 (N_41584,N_39765,N_39796);
nor U41585 (N_41585,N_39562,N_39737);
and U41586 (N_41586,N_39088,N_39622);
xor U41587 (N_41587,N_39719,N_39495);
xnor U41588 (N_41588,N_38163,N_38412);
or U41589 (N_41589,N_38215,N_39071);
nand U41590 (N_41590,N_38750,N_38650);
nor U41591 (N_41591,N_38600,N_39758);
and U41592 (N_41592,N_39935,N_39442);
or U41593 (N_41593,N_39045,N_39022);
nand U41594 (N_41594,N_38925,N_38817);
and U41595 (N_41595,N_39651,N_39453);
or U41596 (N_41596,N_38370,N_39881);
and U41597 (N_41597,N_39012,N_38225);
and U41598 (N_41598,N_39151,N_38645);
and U41599 (N_41599,N_38922,N_38422);
nor U41600 (N_41600,N_39647,N_38638);
xnor U41601 (N_41601,N_38972,N_39197);
and U41602 (N_41602,N_39446,N_38175);
xor U41603 (N_41603,N_38151,N_38202);
nor U41604 (N_41604,N_38571,N_39424);
or U41605 (N_41605,N_38130,N_39298);
or U41606 (N_41606,N_38064,N_38753);
or U41607 (N_41607,N_39586,N_38243);
nor U41608 (N_41608,N_38364,N_38802);
and U41609 (N_41609,N_39772,N_38712);
nand U41610 (N_41610,N_39137,N_39133);
or U41611 (N_41611,N_38263,N_39438);
nand U41612 (N_41612,N_38995,N_38421);
nor U41613 (N_41613,N_38014,N_39670);
nor U41614 (N_41614,N_39049,N_38817);
nand U41615 (N_41615,N_39750,N_38757);
xnor U41616 (N_41616,N_38467,N_38243);
xor U41617 (N_41617,N_38033,N_38699);
nor U41618 (N_41618,N_38668,N_39599);
and U41619 (N_41619,N_39178,N_39741);
nand U41620 (N_41620,N_38323,N_38613);
and U41621 (N_41621,N_38188,N_39281);
xnor U41622 (N_41622,N_39182,N_39506);
and U41623 (N_41623,N_38350,N_38994);
xnor U41624 (N_41624,N_38550,N_39590);
and U41625 (N_41625,N_38922,N_38920);
or U41626 (N_41626,N_39455,N_39294);
or U41627 (N_41627,N_39972,N_39615);
and U41628 (N_41628,N_38106,N_38167);
xor U41629 (N_41629,N_38180,N_39216);
xnor U41630 (N_41630,N_39771,N_38666);
xor U41631 (N_41631,N_39037,N_39331);
or U41632 (N_41632,N_39288,N_39874);
xnor U41633 (N_41633,N_39015,N_39867);
or U41634 (N_41634,N_39628,N_39805);
nand U41635 (N_41635,N_39727,N_39595);
nand U41636 (N_41636,N_38388,N_38526);
nor U41637 (N_41637,N_38849,N_38606);
and U41638 (N_41638,N_39648,N_39549);
and U41639 (N_41639,N_38657,N_38732);
nand U41640 (N_41640,N_38548,N_38144);
nor U41641 (N_41641,N_39985,N_39590);
nor U41642 (N_41642,N_39837,N_38176);
or U41643 (N_41643,N_38768,N_39747);
nor U41644 (N_41644,N_39547,N_38540);
nand U41645 (N_41645,N_39704,N_39537);
or U41646 (N_41646,N_39132,N_39778);
nor U41647 (N_41647,N_39773,N_39367);
or U41648 (N_41648,N_39782,N_39521);
and U41649 (N_41649,N_39104,N_38423);
and U41650 (N_41650,N_39253,N_39165);
nand U41651 (N_41651,N_38548,N_39507);
nand U41652 (N_41652,N_38335,N_39964);
nand U41653 (N_41653,N_39563,N_39875);
nor U41654 (N_41654,N_39423,N_38721);
or U41655 (N_41655,N_38442,N_38859);
or U41656 (N_41656,N_38208,N_38236);
or U41657 (N_41657,N_38029,N_39038);
or U41658 (N_41658,N_38616,N_39134);
nand U41659 (N_41659,N_39704,N_38443);
and U41660 (N_41660,N_38480,N_39127);
xnor U41661 (N_41661,N_39448,N_38888);
and U41662 (N_41662,N_38683,N_39183);
nand U41663 (N_41663,N_39798,N_39856);
and U41664 (N_41664,N_39324,N_39088);
nand U41665 (N_41665,N_39611,N_38165);
nand U41666 (N_41666,N_38037,N_38775);
xnor U41667 (N_41667,N_38746,N_38446);
xor U41668 (N_41668,N_39654,N_39472);
nor U41669 (N_41669,N_38068,N_39352);
xor U41670 (N_41670,N_38532,N_38395);
xor U41671 (N_41671,N_39147,N_38704);
xnor U41672 (N_41672,N_38415,N_39086);
xor U41673 (N_41673,N_39763,N_38055);
nor U41674 (N_41674,N_39389,N_39864);
and U41675 (N_41675,N_39603,N_38410);
or U41676 (N_41676,N_38238,N_39600);
and U41677 (N_41677,N_38685,N_39972);
or U41678 (N_41678,N_39445,N_39200);
or U41679 (N_41679,N_39333,N_38366);
xor U41680 (N_41680,N_39961,N_39473);
and U41681 (N_41681,N_39182,N_38859);
xor U41682 (N_41682,N_39015,N_39071);
nand U41683 (N_41683,N_39783,N_39673);
xnor U41684 (N_41684,N_38358,N_38347);
nand U41685 (N_41685,N_38044,N_38356);
and U41686 (N_41686,N_38704,N_38968);
or U41687 (N_41687,N_39844,N_38525);
or U41688 (N_41688,N_39756,N_39075);
or U41689 (N_41689,N_38616,N_38458);
and U41690 (N_41690,N_38426,N_38903);
nor U41691 (N_41691,N_38137,N_38935);
xor U41692 (N_41692,N_38875,N_38307);
nor U41693 (N_41693,N_39014,N_38634);
nand U41694 (N_41694,N_38133,N_39936);
or U41695 (N_41695,N_38576,N_38224);
and U41696 (N_41696,N_39562,N_38889);
xnor U41697 (N_41697,N_39362,N_38666);
nand U41698 (N_41698,N_38232,N_39013);
and U41699 (N_41699,N_39921,N_38341);
nand U41700 (N_41700,N_38835,N_39898);
or U41701 (N_41701,N_39935,N_38917);
xnor U41702 (N_41702,N_39544,N_39895);
nor U41703 (N_41703,N_39311,N_39767);
and U41704 (N_41704,N_38935,N_38725);
and U41705 (N_41705,N_39494,N_38829);
xnor U41706 (N_41706,N_39637,N_39163);
and U41707 (N_41707,N_38906,N_38338);
xor U41708 (N_41708,N_39797,N_39521);
nand U41709 (N_41709,N_39360,N_39558);
nand U41710 (N_41710,N_38498,N_38613);
nor U41711 (N_41711,N_39747,N_38602);
nor U41712 (N_41712,N_39988,N_39012);
nor U41713 (N_41713,N_39696,N_38295);
or U41714 (N_41714,N_38601,N_38485);
and U41715 (N_41715,N_39161,N_38244);
nand U41716 (N_41716,N_39005,N_39996);
and U41717 (N_41717,N_39937,N_38287);
and U41718 (N_41718,N_39467,N_38128);
and U41719 (N_41719,N_38835,N_38519);
or U41720 (N_41720,N_39290,N_39552);
nand U41721 (N_41721,N_39193,N_38987);
xor U41722 (N_41722,N_38900,N_39140);
and U41723 (N_41723,N_39222,N_38182);
and U41724 (N_41724,N_38063,N_39735);
or U41725 (N_41725,N_39450,N_39172);
xor U41726 (N_41726,N_38201,N_38628);
and U41727 (N_41727,N_39000,N_38568);
and U41728 (N_41728,N_38228,N_38676);
nand U41729 (N_41729,N_39321,N_39850);
or U41730 (N_41730,N_38905,N_39977);
and U41731 (N_41731,N_39018,N_38605);
nand U41732 (N_41732,N_39005,N_38333);
and U41733 (N_41733,N_39048,N_39301);
and U41734 (N_41734,N_38469,N_38391);
nand U41735 (N_41735,N_39435,N_39610);
and U41736 (N_41736,N_39942,N_38135);
xor U41737 (N_41737,N_38976,N_39381);
or U41738 (N_41738,N_38052,N_38489);
xor U41739 (N_41739,N_38491,N_38316);
xnor U41740 (N_41740,N_39065,N_39380);
nand U41741 (N_41741,N_38190,N_38462);
nor U41742 (N_41742,N_38674,N_38227);
nor U41743 (N_41743,N_39013,N_39226);
xor U41744 (N_41744,N_38579,N_39223);
nand U41745 (N_41745,N_38754,N_39415);
nand U41746 (N_41746,N_39165,N_38285);
or U41747 (N_41747,N_38306,N_38405);
and U41748 (N_41748,N_39948,N_38844);
nand U41749 (N_41749,N_39839,N_39366);
nand U41750 (N_41750,N_39398,N_38636);
nand U41751 (N_41751,N_39445,N_38771);
and U41752 (N_41752,N_38674,N_39056);
or U41753 (N_41753,N_39452,N_38709);
or U41754 (N_41754,N_38255,N_39460);
and U41755 (N_41755,N_39530,N_38228);
nand U41756 (N_41756,N_38269,N_39687);
and U41757 (N_41757,N_38138,N_38618);
xnor U41758 (N_41758,N_38165,N_38176);
nor U41759 (N_41759,N_39642,N_38628);
nor U41760 (N_41760,N_39049,N_39961);
nor U41761 (N_41761,N_39165,N_39961);
or U41762 (N_41762,N_38874,N_39045);
nand U41763 (N_41763,N_38514,N_39578);
nor U41764 (N_41764,N_39734,N_39248);
nor U41765 (N_41765,N_38122,N_38884);
xor U41766 (N_41766,N_39634,N_39709);
and U41767 (N_41767,N_38376,N_38030);
and U41768 (N_41768,N_39605,N_38279);
nand U41769 (N_41769,N_38949,N_39652);
xnor U41770 (N_41770,N_38346,N_38580);
or U41771 (N_41771,N_38722,N_38587);
nand U41772 (N_41772,N_38374,N_38223);
and U41773 (N_41773,N_39417,N_38763);
xor U41774 (N_41774,N_38850,N_39430);
nor U41775 (N_41775,N_38777,N_38480);
nor U41776 (N_41776,N_39926,N_39364);
xnor U41777 (N_41777,N_38026,N_38035);
and U41778 (N_41778,N_39553,N_39514);
xor U41779 (N_41779,N_38593,N_39887);
xor U41780 (N_41780,N_39165,N_39339);
nand U41781 (N_41781,N_39604,N_39611);
xnor U41782 (N_41782,N_39838,N_38214);
nor U41783 (N_41783,N_38022,N_39434);
and U41784 (N_41784,N_38536,N_38356);
xnor U41785 (N_41785,N_38482,N_39991);
and U41786 (N_41786,N_38931,N_39575);
xor U41787 (N_41787,N_38075,N_38788);
xor U41788 (N_41788,N_38432,N_38347);
nand U41789 (N_41789,N_38436,N_38347);
and U41790 (N_41790,N_39728,N_39057);
nand U41791 (N_41791,N_38379,N_39923);
nand U41792 (N_41792,N_38506,N_38189);
or U41793 (N_41793,N_38856,N_39184);
xor U41794 (N_41794,N_39749,N_38435);
or U41795 (N_41795,N_38004,N_38692);
and U41796 (N_41796,N_39184,N_39246);
and U41797 (N_41797,N_38234,N_39380);
or U41798 (N_41798,N_39315,N_39706);
nor U41799 (N_41799,N_39168,N_39709);
or U41800 (N_41800,N_39032,N_38217);
xnor U41801 (N_41801,N_39491,N_39752);
or U41802 (N_41802,N_38160,N_38110);
xor U41803 (N_41803,N_39999,N_39453);
xor U41804 (N_41804,N_38569,N_38181);
and U41805 (N_41805,N_39191,N_39384);
or U41806 (N_41806,N_38525,N_38485);
xnor U41807 (N_41807,N_38710,N_39596);
xor U41808 (N_41808,N_38535,N_38471);
or U41809 (N_41809,N_39517,N_39734);
nand U41810 (N_41810,N_38532,N_39368);
nor U41811 (N_41811,N_38156,N_39113);
and U41812 (N_41812,N_39793,N_38805);
or U41813 (N_41813,N_38731,N_38341);
nand U41814 (N_41814,N_38452,N_38930);
nor U41815 (N_41815,N_39715,N_38426);
nor U41816 (N_41816,N_38747,N_38467);
or U41817 (N_41817,N_38042,N_38938);
and U41818 (N_41818,N_39301,N_38354);
nor U41819 (N_41819,N_38982,N_39875);
nand U41820 (N_41820,N_39951,N_39446);
xor U41821 (N_41821,N_39534,N_39770);
nand U41822 (N_41822,N_38643,N_38719);
or U41823 (N_41823,N_39939,N_39944);
nand U41824 (N_41824,N_39705,N_38746);
nor U41825 (N_41825,N_39903,N_39848);
nand U41826 (N_41826,N_38997,N_39784);
or U41827 (N_41827,N_38080,N_38039);
nand U41828 (N_41828,N_39333,N_39978);
or U41829 (N_41829,N_38268,N_39825);
nand U41830 (N_41830,N_39105,N_38026);
and U41831 (N_41831,N_38766,N_38861);
xnor U41832 (N_41832,N_38658,N_39186);
nand U41833 (N_41833,N_38154,N_38676);
nor U41834 (N_41834,N_38068,N_38297);
and U41835 (N_41835,N_39065,N_38262);
nor U41836 (N_41836,N_38183,N_38179);
or U41837 (N_41837,N_39819,N_39775);
nand U41838 (N_41838,N_38487,N_38345);
xnor U41839 (N_41839,N_38691,N_38001);
or U41840 (N_41840,N_38973,N_39338);
nor U41841 (N_41841,N_39994,N_39478);
and U41842 (N_41842,N_39386,N_39757);
and U41843 (N_41843,N_39070,N_39827);
and U41844 (N_41844,N_38691,N_38805);
nor U41845 (N_41845,N_38286,N_38926);
xor U41846 (N_41846,N_39367,N_38714);
nor U41847 (N_41847,N_39668,N_39806);
nor U41848 (N_41848,N_39710,N_39999);
or U41849 (N_41849,N_39823,N_38791);
nand U41850 (N_41850,N_39576,N_39721);
and U41851 (N_41851,N_38801,N_38143);
or U41852 (N_41852,N_38970,N_38148);
nor U41853 (N_41853,N_39102,N_39862);
and U41854 (N_41854,N_39023,N_39597);
xnor U41855 (N_41855,N_39556,N_39771);
nor U41856 (N_41856,N_38678,N_39276);
nand U41857 (N_41857,N_39703,N_39661);
or U41858 (N_41858,N_38318,N_39132);
nand U41859 (N_41859,N_39709,N_39879);
nand U41860 (N_41860,N_39026,N_39504);
and U41861 (N_41861,N_39158,N_38059);
and U41862 (N_41862,N_39421,N_39449);
and U41863 (N_41863,N_38740,N_38924);
xnor U41864 (N_41864,N_38281,N_38975);
xnor U41865 (N_41865,N_39609,N_39389);
and U41866 (N_41866,N_38864,N_39719);
and U41867 (N_41867,N_39804,N_39051);
xnor U41868 (N_41868,N_39258,N_39576);
or U41869 (N_41869,N_39986,N_38347);
and U41870 (N_41870,N_38500,N_38070);
nand U41871 (N_41871,N_38049,N_38645);
nor U41872 (N_41872,N_39896,N_39044);
xnor U41873 (N_41873,N_38218,N_39011);
xnor U41874 (N_41874,N_39278,N_39199);
and U41875 (N_41875,N_39447,N_38760);
nor U41876 (N_41876,N_39204,N_39885);
xor U41877 (N_41877,N_39432,N_39565);
nor U41878 (N_41878,N_38307,N_38969);
nor U41879 (N_41879,N_38043,N_39855);
and U41880 (N_41880,N_38723,N_39970);
nor U41881 (N_41881,N_38917,N_38144);
xnor U41882 (N_41882,N_38306,N_39292);
nor U41883 (N_41883,N_38706,N_38378);
nand U41884 (N_41884,N_38015,N_39332);
and U41885 (N_41885,N_39815,N_38226);
and U41886 (N_41886,N_38116,N_39993);
and U41887 (N_41887,N_38125,N_39101);
or U41888 (N_41888,N_39588,N_39338);
nand U41889 (N_41889,N_39477,N_39871);
nor U41890 (N_41890,N_39858,N_38682);
nand U41891 (N_41891,N_39407,N_38474);
or U41892 (N_41892,N_39514,N_38795);
nand U41893 (N_41893,N_39506,N_38785);
xor U41894 (N_41894,N_39232,N_38376);
and U41895 (N_41895,N_39429,N_39899);
nand U41896 (N_41896,N_39254,N_38176);
and U41897 (N_41897,N_39112,N_38106);
or U41898 (N_41898,N_38997,N_39315);
or U41899 (N_41899,N_38673,N_38820);
nand U41900 (N_41900,N_39277,N_39822);
xnor U41901 (N_41901,N_39745,N_39121);
xor U41902 (N_41902,N_38208,N_39396);
nand U41903 (N_41903,N_39436,N_39724);
nor U41904 (N_41904,N_38466,N_38863);
nor U41905 (N_41905,N_39847,N_39767);
and U41906 (N_41906,N_39160,N_39016);
nor U41907 (N_41907,N_38823,N_38484);
and U41908 (N_41908,N_39653,N_39216);
and U41909 (N_41909,N_38839,N_38329);
and U41910 (N_41910,N_39255,N_38107);
and U41911 (N_41911,N_39431,N_38825);
and U41912 (N_41912,N_39069,N_39331);
xnor U41913 (N_41913,N_38175,N_39493);
or U41914 (N_41914,N_39398,N_39158);
nand U41915 (N_41915,N_38497,N_38356);
xnor U41916 (N_41916,N_39954,N_39162);
nand U41917 (N_41917,N_39243,N_38476);
xnor U41918 (N_41918,N_38626,N_38694);
nand U41919 (N_41919,N_38336,N_38082);
or U41920 (N_41920,N_38177,N_39495);
nand U41921 (N_41921,N_38251,N_38318);
xnor U41922 (N_41922,N_38132,N_39588);
nand U41923 (N_41923,N_38744,N_38110);
xnor U41924 (N_41924,N_39169,N_38063);
nor U41925 (N_41925,N_38844,N_38149);
xor U41926 (N_41926,N_39577,N_39799);
or U41927 (N_41927,N_39100,N_38767);
and U41928 (N_41928,N_38202,N_38567);
or U41929 (N_41929,N_38899,N_39883);
nor U41930 (N_41930,N_39977,N_39150);
or U41931 (N_41931,N_38976,N_38812);
nand U41932 (N_41932,N_39112,N_39074);
nor U41933 (N_41933,N_39793,N_38012);
and U41934 (N_41934,N_38572,N_39208);
and U41935 (N_41935,N_38418,N_39760);
nand U41936 (N_41936,N_39828,N_38780);
and U41937 (N_41937,N_38529,N_39319);
xor U41938 (N_41938,N_38467,N_38788);
and U41939 (N_41939,N_38306,N_38475);
xor U41940 (N_41940,N_38954,N_38360);
or U41941 (N_41941,N_38513,N_39747);
nor U41942 (N_41942,N_39069,N_38314);
or U41943 (N_41943,N_39169,N_39417);
or U41944 (N_41944,N_38805,N_38977);
and U41945 (N_41945,N_39199,N_38264);
xor U41946 (N_41946,N_38860,N_38519);
xor U41947 (N_41947,N_38418,N_39355);
nor U41948 (N_41948,N_38638,N_39088);
xor U41949 (N_41949,N_38253,N_39913);
or U41950 (N_41950,N_38204,N_39152);
and U41951 (N_41951,N_39938,N_38603);
and U41952 (N_41952,N_38273,N_38478);
xnor U41953 (N_41953,N_39040,N_38845);
or U41954 (N_41954,N_39011,N_39378);
nor U41955 (N_41955,N_39965,N_38091);
xnor U41956 (N_41956,N_39873,N_39405);
and U41957 (N_41957,N_38927,N_38365);
or U41958 (N_41958,N_38117,N_38149);
or U41959 (N_41959,N_38756,N_39546);
xnor U41960 (N_41960,N_38282,N_39696);
or U41961 (N_41961,N_39716,N_39259);
xor U41962 (N_41962,N_39475,N_39914);
xor U41963 (N_41963,N_38586,N_38659);
or U41964 (N_41964,N_38958,N_39250);
nand U41965 (N_41965,N_39707,N_39913);
nand U41966 (N_41966,N_39922,N_39694);
or U41967 (N_41967,N_39433,N_38144);
xnor U41968 (N_41968,N_39793,N_39499);
and U41969 (N_41969,N_39060,N_38499);
and U41970 (N_41970,N_39960,N_38711);
xor U41971 (N_41971,N_38610,N_39583);
nor U41972 (N_41972,N_39858,N_38281);
xor U41973 (N_41973,N_38539,N_39349);
nor U41974 (N_41974,N_38051,N_38202);
and U41975 (N_41975,N_38652,N_39767);
or U41976 (N_41976,N_38521,N_38000);
or U41977 (N_41977,N_39841,N_39257);
and U41978 (N_41978,N_39823,N_39844);
nor U41979 (N_41979,N_39732,N_39053);
xor U41980 (N_41980,N_39160,N_39404);
and U41981 (N_41981,N_39270,N_39460);
or U41982 (N_41982,N_38654,N_38258);
nor U41983 (N_41983,N_38572,N_39675);
or U41984 (N_41984,N_38891,N_38009);
or U41985 (N_41985,N_38477,N_39690);
nor U41986 (N_41986,N_38766,N_39791);
xor U41987 (N_41987,N_39201,N_38251);
nand U41988 (N_41988,N_39929,N_39068);
and U41989 (N_41989,N_38611,N_38688);
nand U41990 (N_41990,N_39341,N_38952);
nand U41991 (N_41991,N_39396,N_39491);
xor U41992 (N_41992,N_38426,N_39046);
or U41993 (N_41993,N_38274,N_39596);
nor U41994 (N_41994,N_39202,N_38448);
nand U41995 (N_41995,N_39238,N_39330);
nor U41996 (N_41996,N_39300,N_38270);
nor U41997 (N_41997,N_39172,N_39516);
and U41998 (N_41998,N_39185,N_38858);
or U41999 (N_41999,N_38277,N_39040);
nor U42000 (N_42000,N_40490,N_40171);
xnor U42001 (N_42001,N_40140,N_40448);
and U42002 (N_42002,N_40526,N_40762);
or U42003 (N_42003,N_41127,N_41190);
and U42004 (N_42004,N_41722,N_40331);
or U42005 (N_42005,N_41430,N_41147);
or U42006 (N_42006,N_40091,N_40803);
or U42007 (N_42007,N_40181,N_41259);
and U42008 (N_42008,N_40728,N_41058);
or U42009 (N_42009,N_41726,N_41186);
xnor U42010 (N_42010,N_41841,N_41605);
nand U42011 (N_42011,N_40115,N_41923);
nand U42012 (N_42012,N_41702,N_41176);
xor U42013 (N_42013,N_41326,N_41482);
or U42014 (N_42014,N_41325,N_41636);
or U42015 (N_42015,N_41477,N_40363);
nor U42016 (N_42016,N_40040,N_40218);
xnor U42017 (N_42017,N_41341,N_41081);
xnor U42018 (N_42018,N_41836,N_40816);
or U42019 (N_42019,N_40642,N_40824);
xnor U42020 (N_42020,N_41216,N_41301);
nor U42021 (N_42021,N_40174,N_40295);
nor U42022 (N_42022,N_41932,N_41268);
nor U42023 (N_42023,N_40608,N_40794);
nor U42024 (N_42024,N_40279,N_40635);
xor U42025 (N_42025,N_40423,N_40583);
nand U42026 (N_42026,N_40383,N_40597);
xor U42027 (N_42027,N_41600,N_41908);
and U42028 (N_42028,N_40437,N_40001);
xor U42029 (N_42029,N_41876,N_41562);
or U42030 (N_42030,N_40334,N_40875);
or U42031 (N_42031,N_41360,N_40492);
or U42032 (N_42032,N_41742,N_41468);
nor U42033 (N_42033,N_41161,N_40850);
or U42034 (N_42034,N_41311,N_41135);
nor U42035 (N_42035,N_40791,N_40451);
and U42036 (N_42036,N_40516,N_41116);
xor U42037 (N_42037,N_40907,N_40258);
xor U42038 (N_42038,N_40746,N_40256);
and U42039 (N_42039,N_40864,N_40060);
and U42040 (N_42040,N_40111,N_41957);
and U42041 (N_42041,N_40679,N_41038);
nor U42042 (N_42042,N_40846,N_41180);
or U42043 (N_42043,N_41055,N_40053);
xor U42044 (N_42044,N_41099,N_40231);
nand U42045 (N_42045,N_41552,N_40827);
or U42046 (N_42046,N_41648,N_41453);
nand U42047 (N_42047,N_40872,N_41500);
nor U42048 (N_42048,N_41663,N_40800);
xnor U42049 (N_42049,N_41888,N_40068);
nor U42050 (N_42050,N_40687,N_41304);
nor U42051 (N_42051,N_40579,N_41461);
nor U42052 (N_42052,N_40806,N_40229);
and U42053 (N_42053,N_40325,N_41434);
or U42054 (N_42054,N_40236,N_41222);
or U42055 (N_42055,N_41357,N_41654);
nor U42056 (N_42056,N_41917,N_40403);
nor U42057 (N_42057,N_41043,N_40213);
nor U42058 (N_42058,N_40613,N_40012);
xnor U42059 (N_42059,N_41194,N_40688);
nor U42060 (N_42060,N_41983,N_41735);
or U42061 (N_42061,N_40386,N_40998);
nand U42062 (N_42062,N_40939,N_40961);
nand U42063 (N_42063,N_41313,N_41721);
and U42064 (N_42064,N_41064,N_40949);
nor U42065 (N_42065,N_41681,N_40049);
xor U42066 (N_42066,N_41246,N_40967);
nor U42067 (N_42067,N_41181,N_40191);
xnor U42068 (N_42068,N_41741,N_40641);
or U42069 (N_42069,N_40653,N_40724);
and U42070 (N_42070,N_40350,N_40539);
nand U42071 (N_42071,N_40960,N_41974);
nor U42072 (N_42072,N_40376,N_40156);
and U42073 (N_42073,N_41238,N_40739);
or U42074 (N_42074,N_41228,N_41336);
nor U42075 (N_42075,N_40695,N_40084);
xor U42076 (N_42076,N_41329,N_40668);
nor U42077 (N_42077,N_40149,N_41077);
nor U42078 (N_42078,N_40254,N_41340);
and U42079 (N_42079,N_41850,N_41130);
and U42080 (N_42080,N_41272,N_40249);
xor U42081 (N_42081,N_41240,N_40102);
and U42082 (N_42082,N_40931,N_41730);
nor U42083 (N_42083,N_41380,N_40580);
or U42084 (N_42084,N_40896,N_41182);
nor U42085 (N_42085,N_41188,N_40116);
nand U42086 (N_42086,N_41635,N_41203);
and U42087 (N_42087,N_40372,N_41758);
or U42088 (N_42088,N_41886,N_41124);
xnor U42089 (N_42089,N_41369,N_41003);
xnor U42090 (N_42090,N_41433,N_40065);
nand U42091 (N_42091,N_40133,N_40203);
or U42092 (N_42092,N_40158,N_40639);
nor U42093 (N_42093,N_41112,N_41693);
xnor U42094 (N_42094,N_41596,N_40211);
and U42095 (N_42095,N_40388,N_40222);
nor U42096 (N_42096,N_41437,N_40311);
xnor U42097 (N_42097,N_41348,N_41354);
or U42098 (N_42098,N_40333,N_40019);
nand U42099 (N_42099,N_41084,N_40301);
xnor U42100 (N_42100,N_40245,N_41017);
and U42101 (N_42101,N_40699,N_40953);
and U42102 (N_42102,N_41986,N_41746);
nor U42103 (N_42103,N_41457,N_40031);
nand U42104 (N_42104,N_40702,N_41144);
nor U42105 (N_42105,N_40066,N_40811);
nor U42106 (N_42106,N_40856,N_41717);
nand U42107 (N_42107,N_41108,N_41901);
nor U42108 (N_42108,N_40889,N_40082);
or U42109 (N_42109,N_41692,N_40131);
or U42110 (N_42110,N_41294,N_41981);
and U42111 (N_42111,N_41873,N_40129);
nand U42112 (N_42112,N_41868,N_40230);
or U42113 (N_42113,N_41364,N_41193);
and U42114 (N_42114,N_41456,N_41395);
nand U42115 (N_42115,N_40566,N_41015);
and U42116 (N_42116,N_41418,N_41470);
xnor U42117 (N_42117,N_41572,N_41443);
nor U42118 (N_42118,N_41624,N_41544);
xnor U42119 (N_42119,N_41531,N_40975);
nand U42120 (N_42120,N_41211,N_40757);
and U42121 (N_42121,N_40795,N_40667);
or U42122 (N_42122,N_40654,N_41813);
and U42123 (N_42123,N_40424,N_40602);
and U42124 (N_42124,N_40523,N_41292);
nand U42125 (N_42125,N_40081,N_40737);
xor U42126 (N_42126,N_41997,N_41761);
or U42127 (N_42127,N_41706,N_41258);
xor U42128 (N_42128,N_41031,N_41881);
xor U42129 (N_42129,N_41783,N_40652);
nand U42130 (N_42130,N_41109,N_41241);
or U42131 (N_42131,N_41314,N_41494);
or U42132 (N_42132,N_40464,N_40938);
or U42133 (N_42133,N_40479,N_41802);
xnor U42134 (N_42134,N_40705,N_41811);
xor U42135 (N_42135,N_40310,N_40810);
and U42136 (N_42136,N_41484,N_41611);
or U42137 (N_42137,N_41963,N_40585);
xnor U42138 (N_42138,N_41858,N_41764);
or U42139 (N_42139,N_40221,N_40360);
nand U42140 (N_42140,N_40833,N_41065);
or U42141 (N_42141,N_41283,N_41990);
nor U42142 (N_42142,N_40849,N_41736);
nor U42143 (N_42143,N_40521,N_41964);
and U42144 (N_42144,N_41256,N_40582);
or U42145 (N_42145,N_40290,N_40003);
nand U42146 (N_42146,N_40027,N_41392);
nor U42147 (N_42147,N_41709,N_40493);
xor U42148 (N_42148,N_41248,N_41793);
or U42149 (N_42149,N_41271,N_40793);
nand U42150 (N_42150,N_40441,N_41198);
nor U42151 (N_42151,N_40101,N_40267);
nand U42152 (N_42152,N_41138,N_41310);
xnor U42153 (N_42153,N_40789,N_41425);
or U42154 (N_42154,N_40948,N_41195);
and U42155 (N_42155,N_41607,N_41987);
or U42156 (N_42156,N_40572,N_41541);
nand U42157 (N_42157,N_40586,N_40745);
and U42158 (N_42158,N_40165,N_40125);
xnor U42159 (N_42159,N_40603,N_41106);
nand U42160 (N_42160,N_41522,N_40512);
and U42161 (N_42161,N_40275,N_41447);
nor U42162 (N_42162,N_41865,N_40765);
or U42163 (N_42163,N_41778,N_40238);
or U42164 (N_42164,N_40039,N_40505);
xnor U42165 (N_42165,N_40721,N_41724);
or U42166 (N_42166,N_40911,N_41011);
or U42167 (N_42167,N_41739,N_41141);
and U42168 (N_42168,N_40294,N_41414);
xor U42169 (N_42169,N_41556,N_41894);
or U42170 (N_42170,N_40204,N_41975);
nand U42171 (N_42171,N_40573,N_41202);
xnor U42172 (N_42172,N_40237,N_41496);
and U42173 (N_42173,N_41563,N_41929);
xnor U42174 (N_42174,N_40227,N_41087);
nand U42175 (N_42175,N_41966,N_40624);
or U42176 (N_42176,N_41740,N_40255);
nor U42177 (N_42177,N_40543,N_41543);
and U42178 (N_42178,N_41651,N_41179);
xnor U42179 (N_42179,N_41826,N_40339);
nor U42180 (N_42180,N_41570,N_40137);
xor U42181 (N_42181,N_40515,N_40980);
nand U42182 (N_42182,N_40893,N_41703);
nand U42183 (N_42183,N_40822,N_40250);
xor U42184 (N_42184,N_41105,N_40062);
nor U42185 (N_42185,N_40020,N_40665);
xnor U42186 (N_42186,N_41845,N_41375);
xor U42187 (N_42187,N_40844,N_40392);
and U42188 (N_42188,N_41864,N_40917);
nand U42189 (N_42189,N_40957,N_41690);
nand U42190 (N_42190,N_40244,N_40405);
xor U42191 (N_42191,N_41595,N_41688);
nand U42192 (N_42192,N_41132,N_40010);
nor U42193 (N_42193,N_40243,N_41689);
xnor U42194 (N_42194,N_41455,N_40324);
nand U42195 (N_42195,N_41766,N_40536);
xnor U42196 (N_42196,N_40368,N_40271);
and U42197 (N_42197,N_40365,N_40086);
nand U42198 (N_42198,N_41503,N_41435);
xor U42199 (N_42199,N_40106,N_40418);
nand U42200 (N_42200,N_41946,N_41860);
nand U42201 (N_42201,N_40742,N_41091);
xnor U42202 (N_42202,N_40600,N_41097);
nand U42203 (N_42203,N_40735,N_40345);
or U42204 (N_42204,N_40943,N_40873);
nor U42205 (N_42205,N_41576,N_40529);
or U42206 (N_42206,N_40432,N_40183);
xnor U42207 (N_42207,N_41041,N_41660);
and U42208 (N_42208,N_40925,N_40495);
xnor U42209 (N_42209,N_40828,N_41386);
nand U42210 (N_42210,N_41781,N_40918);
nand U42211 (N_42211,N_41927,N_41823);
xor U42212 (N_42212,N_40192,N_41442);
nand U42213 (N_42213,N_41679,N_40775);
or U42214 (N_42214,N_40663,N_40172);
and U42215 (N_42215,N_40933,N_40449);
or U42216 (N_42216,N_40371,N_41048);
nand U42217 (N_42217,N_41027,N_41977);
and U42218 (N_42218,N_41073,N_40825);
xnor U42219 (N_42219,N_41286,N_41320);
nor U42220 (N_42220,N_40196,N_40971);
nor U42221 (N_42221,N_41396,N_40314);
nand U42222 (N_42222,N_40942,N_41535);
xor U42223 (N_42223,N_41363,N_40160);
nor U42224 (N_42224,N_41010,N_41005);
nor U42225 (N_42225,N_41903,N_41490);
or U42226 (N_42226,N_40814,N_40812);
or U42227 (N_42227,N_41670,N_41972);
nand U42228 (N_42228,N_41851,N_41644);
nor U42229 (N_42229,N_40879,N_41322);
or U42230 (N_42230,N_40093,N_40182);
xnor U42231 (N_42231,N_40344,N_40234);
nor U42232 (N_42232,N_40138,N_41224);
or U42233 (N_42233,N_40364,N_41574);
and U42234 (N_42234,N_40459,N_41473);
xnor U42235 (N_42235,N_41206,N_41843);
nor U42236 (N_42236,N_40269,N_40621);
nor U42237 (N_42237,N_40660,N_41497);
and U42238 (N_42238,N_41047,N_41007);
or U42239 (N_42239,N_40940,N_40103);
or U42240 (N_42240,N_40853,N_41847);
and U42241 (N_42241,N_40693,N_40581);
or U42242 (N_42242,N_40513,N_40951);
and U42243 (N_42243,N_41002,N_40709);
and U42244 (N_42244,N_40753,N_41356);
and U42245 (N_42245,N_40589,N_40527);
nand U42246 (N_42246,N_40443,N_41581);
nor U42247 (N_42247,N_40578,N_41267);
nand U42248 (N_42248,N_40535,N_40494);
or U42249 (N_42249,N_41316,N_40385);
nand U42250 (N_42250,N_41111,N_41936);
nor U42251 (N_42251,N_41829,N_40335);
nand U42252 (N_42252,N_41790,N_40916);
xnor U42253 (N_42253,N_41683,N_41131);
nand U42254 (N_42254,N_41520,N_40177);
nor U42255 (N_42255,N_41485,N_41968);
xor U42256 (N_42256,N_40570,N_41287);
nor U42257 (N_42257,N_41819,N_40764);
nand U42258 (N_42258,N_40591,N_41221);
xor U42259 (N_42259,N_41390,N_41217);
and U42260 (N_42260,N_40650,N_40926);
nand U42261 (N_42261,N_40422,N_40359);
and U42262 (N_42262,N_41393,N_40538);
xor U42263 (N_42263,N_40818,N_41650);
nor U42264 (N_42264,N_40646,N_40743);
xnor U42265 (N_42265,N_41512,N_40223);
or U42266 (N_42266,N_41962,N_41906);
xor U42267 (N_42267,N_40966,N_40870);
xnor U42268 (N_42268,N_41625,N_41852);
nor U42269 (N_42269,N_40763,N_41093);
xor U42270 (N_42270,N_41634,N_40104);
xnor U42271 (N_42271,N_40122,N_41063);
nor U42272 (N_42272,N_40018,N_41712);
nor U42273 (N_42273,N_40077,N_41402);
nor U42274 (N_42274,N_41980,N_41428);
or U42275 (N_42275,N_40601,N_41912);
and U42276 (N_42276,N_41776,N_40829);
nand U42277 (N_42277,N_40124,N_40910);
nor U42278 (N_42278,N_40291,N_41508);
nand U42279 (N_42279,N_41158,N_40734);
nor U42280 (N_42280,N_40740,N_40657);
and U42281 (N_42281,N_41426,N_40528);
nand U42282 (N_42282,N_41372,N_41044);
xor U42283 (N_42283,N_41582,N_40683);
nand U42284 (N_42284,N_41649,N_40799);
or U42285 (N_42285,N_40067,N_40792);
xor U42286 (N_42286,N_41952,N_40970);
xor U42287 (N_42287,N_41374,N_41284);
or U42288 (N_42288,N_41505,N_40461);
nor U42289 (N_42289,N_41818,N_41958);
or U42290 (N_42290,N_41924,N_40456);
and U42291 (N_42291,N_41377,N_40035);
xnor U42292 (N_42292,N_40047,N_40399);
or U42293 (N_42293,N_40554,N_41480);
or U42294 (N_42294,N_40913,N_40075);
nor U42295 (N_42295,N_41633,N_40785);
and U42296 (N_42296,N_41026,N_40598);
nor U42297 (N_42297,N_41998,N_41359);
nand U42298 (N_42298,N_41604,N_40747);
xor U42299 (N_42299,N_40944,N_40315);
nor U42300 (N_42300,N_41707,N_40831);
nor U42301 (N_42301,N_40779,N_41299);
nor U42302 (N_42302,N_40074,N_41708);
or U42303 (N_42303,N_40120,N_40712);
or U42304 (N_42304,N_41884,N_41245);
or U42305 (N_42305,N_40014,N_41028);
nor U42306 (N_42306,N_41796,N_41115);
or U42307 (N_42307,N_40248,N_40397);
xor U42308 (N_42308,N_40777,N_41511);
xnor U42309 (N_42309,N_40008,N_40590);
nor U42310 (N_42310,N_41810,N_40848);
and U42311 (N_42311,N_41687,N_40072);
nor U42312 (N_42312,N_40078,N_41351);
xnor U42313 (N_42313,N_40752,N_40952);
or U42314 (N_42314,N_40552,N_41928);
nand U42315 (N_42315,N_41558,N_41092);
and U42316 (N_42316,N_40083,N_41768);
nand U42317 (N_42317,N_41459,N_41538);
nand U42318 (N_42318,N_41784,N_40316);
nor U42319 (N_42319,N_40684,N_41728);
or U42320 (N_42320,N_40395,N_40332);
nand U42321 (N_42321,N_40013,N_41458);
and U42322 (N_42322,N_40587,N_41332);
and U42323 (N_42323,N_41514,N_41891);
nand U42324 (N_42324,N_40284,N_41820);
or U42325 (N_42325,N_40381,N_41815);
and U42326 (N_42326,N_40080,N_40867);
or U42327 (N_42327,N_41502,N_41639);
and U42328 (N_42328,N_41139,N_40408);
or U42329 (N_42329,N_41244,N_40313);
and U42330 (N_42330,N_41344,N_41406);
nor U42331 (N_42331,N_40146,N_41382);
and U42332 (N_42332,N_41830,N_40599);
nand U42333 (N_42333,N_40773,N_41573);
nand U42334 (N_42334,N_41792,N_41715);
and U42335 (N_42335,N_41166,N_40268);
and U42336 (N_42336,N_41300,N_40030);
and U42337 (N_42337,N_40715,N_40736);
xnor U42338 (N_42338,N_40166,N_41530);
and U42339 (N_42339,N_41879,N_41817);
nand U42340 (N_42340,N_41282,N_41309);
nor U42341 (N_42341,N_40860,N_41018);
or U42342 (N_42342,N_41874,N_40945);
nor U42343 (N_42343,N_40935,N_41070);
nand U42344 (N_42344,N_41451,N_41014);
and U42345 (N_42345,N_41812,N_41212);
xnor U42346 (N_42346,N_40780,N_40438);
or U42347 (N_42347,N_40404,N_40261);
xnor U42348 (N_42348,N_41822,N_40520);
or U42349 (N_42349,N_41226,N_41699);
or U42350 (N_42350,N_40225,N_41469);
nor U42351 (N_42351,N_41909,N_40052);
nor U42352 (N_42352,N_41350,N_41523);
and U42353 (N_42353,N_41960,N_41905);
or U42354 (N_42354,N_41780,N_40787);
or U42355 (N_42355,N_40946,N_41398);
nand U42356 (N_42356,N_41916,N_41436);
nand U42357 (N_42357,N_41675,N_41760);
nor U42358 (N_42358,N_40710,N_41030);
nor U42359 (N_42359,N_40436,N_40769);
and U42360 (N_42360,N_41237,N_40379);
nand U42361 (N_42361,N_40700,N_41861);
and U42362 (N_42362,N_41101,N_41976);
nand U42363 (N_42363,N_40126,N_40760);
and U42364 (N_42364,N_40341,N_41857);
and U42365 (N_42365,N_40612,N_40409);
nor U42366 (N_42366,N_41612,N_40092);
and U42367 (N_42367,N_40299,N_40420);
and U42368 (N_42368,N_41452,N_41013);
or U42369 (N_42369,N_41247,N_40978);
nor U42370 (N_42370,N_41201,N_40377);
nand U42371 (N_42371,N_40499,N_40750);
xor U42372 (N_42372,N_41995,N_41545);
nor U42373 (N_42373,N_41765,N_41463);
or U42374 (N_42374,N_40309,N_40452);
nand U42375 (N_42375,N_41889,N_41799);
xnor U42376 (N_42376,N_40055,N_40038);
or U42377 (N_42377,N_41384,N_41560);
nand U42378 (N_42378,N_41527,N_41913);
or U42379 (N_42379,N_40026,N_40997);
or U42380 (N_42380,N_40119,N_40929);
or U42381 (N_42381,N_40167,N_41704);
and U42382 (N_42382,N_41673,N_40164);
xor U42383 (N_42383,N_40645,N_41462);
or U42384 (N_42384,N_41755,N_40962);
nand U42385 (N_42385,N_41775,N_41590);
and U42386 (N_42386,N_41536,N_41239);
nor U42387 (N_42387,N_41791,N_41930);
nand U42388 (N_42388,N_40009,N_40882);
xor U42389 (N_42389,N_41233,N_41183);
nor U42390 (N_42390,N_40704,N_40776);
nand U42391 (N_42391,N_41750,N_40046);
nand U42392 (N_42392,N_41123,N_40903);
nor U42393 (N_42393,N_40274,N_41056);
nor U42394 (N_42394,N_40406,N_41561);
nand U42395 (N_42395,N_41526,N_40079);
xnor U42396 (N_42396,N_40865,N_41568);
xor U42397 (N_42397,N_40974,N_41723);
xnor U42398 (N_42398,N_41478,N_41037);
and U42399 (N_42399,N_41479,N_41645);
xor U42400 (N_42400,N_41991,N_40169);
xor U42401 (N_42401,N_41528,N_40987);
or U42402 (N_42402,N_40037,N_41674);
nand U42403 (N_42403,N_40936,N_40061);
and U42404 (N_42404,N_41516,N_40427);
nand U42405 (N_42405,N_40934,N_40890);
or U42406 (N_42406,N_40293,N_41095);
xnor U42407 (N_42407,N_40994,N_40134);
nor U42408 (N_42408,N_41165,N_41609);
and U42409 (N_42409,N_40729,N_40537);
and U42410 (N_42410,N_40841,N_40932);
nor U42411 (N_42411,N_41994,N_41236);
and U42412 (N_42412,N_41564,N_40625);
nor U42413 (N_42413,N_40006,N_40207);
and U42414 (N_42414,N_40280,N_41794);
or U42415 (N_42415,N_40193,N_40755);
or U42416 (N_42416,N_41278,N_41883);
and U42417 (N_42417,N_41464,N_41854);
nand U42418 (N_42418,N_40281,N_41078);
or U42419 (N_42419,N_40412,N_41880);
or U42420 (N_42420,N_40575,N_40189);
or U42421 (N_42421,N_41427,N_41506);
xnor U42422 (N_42422,N_40902,N_41501);
xor U42423 (N_42423,N_41410,N_41695);
nor U42424 (N_42424,N_40996,N_40723);
xor U42425 (N_42425,N_41066,N_40210);
nor U42426 (N_42426,N_41965,N_40050);
xnor U42427 (N_42427,N_40549,N_40253);
xor U42428 (N_42428,N_40797,N_41255);
xnor U42429 (N_42429,N_41155,N_41825);
or U42430 (N_42430,N_40476,N_40462);
and U42431 (N_42431,N_40626,N_41806);
xor U42432 (N_42432,N_41697,N_41659);
xor U42433 (N_42433,N_40500,N_41737);
xor U42434 (N_42434,N_41057,N_40298);
nor U42435 (N_42435,N_40112,N_41515);
nor U42436 (N_42436,N_41488,N_40897);
nor U42437 (N_42437,N_40842,N_40766);
nor U42438 (N_42438,N_41075,N_41417);
or U42439 (N_42439,N_41999,N_41266);
or U42440 (N_42440,N_40632,N_41150);
or U42441 (N_42441,N_41591,N_41725);
and U42442 (N_42442,N_41339,N_41257);
and U42443 (N_42443,N_41349,N_41415);
xor U42444 (N_42444,N_40370,N_40215);
nand U42445 (N_42445,N_40450,N_41982);
nand U42446 (N_42446,N_41751,N_41303);
nand U42447 (N_42447,N_41487,N_40655);
xor U42448 (N_42448,N_40878,N_40670);
xnor U42449 (N_42449,N_40501,N_41647);
or U42450 (N_42450,N_41638,N_40358);
xnor U42451 (N_42451,N_41085,N_41956);
nor U42452 (N_42452,N_40353,N_40021);
and U42453 (N_42453,N_40048,N_41931);
nand U42454 (N_42454,N_40201,N_41853);
xor U42455 (N_42455,N_40384,N_41404);
xor U42456 (N_42456,N_41992,N_40110);
nor U42457 (N_42457,N_40886,N_40387);
nor U42458 (N_42458,N_40312,N_41666);
xor U42459 (N_42459,N_41872,N_41738);
and U42460 (N_42460,N_41009,N_41513);
nand U42461 (N_42461,N_41366,N_41342);
and U42462 (N_42462,N_40781,N_41347);
xor U42463 (N_42463,N_41291,N_40919);
nand U42464 (N_42464,N_40468,N_40265);
or U42465 (N_42465,N_41173,N_40958);
and U42466 (N_42466,N_40063,N_40680);
nor U42467 (N_42467,N_40540,N_40330);
nor U42468 (N_42468,N_40562,N_40348);
nand U42469 (N_42469,N_41481,N_41448);
nand U42470 (N_42470,N_41499,N_41337);
or U42471 (N_42471,N_41554,N_41907);
nand U42472 (N_42472,N_40057,N_40984);
xor U42473 (N_42473,N_40927,N_40731);
nand U42474 (N_42474,N_40871,N_41012);
or U42475 (N_42475,N_40402,N_40532);
nand U42476 (N_42476,N_40444,N_41678);
and U42477 (N_42477,N_41029,N_40969);
and U42478 (N_42478,N_41388,N_41323);
xor U42479 (N_42479,N_41330,N_41920);
nand U42480 (N_42480,N_41749,N_40005);
nor U42481 (N_42481,N_41602,N_40714);
nand U42482 (N_42482,N_41537,N_40751);
nor U42483 (N_42483,N_41493,N_40504);
nor U42484 (N_42484,N_41532,N_40163);
and U42485 (N_42485,N_41383,N_40272);
and U42486 (N_42486,N_40446,N_40622);
and U42487 (N_42487,N_40161,N_41385);
and U42488 (N_42488,N_41207,N_41269);
and U42489 (N_42489,N_41779,N_41664);
xor U42490 (N_42490,N_40908,N_41331);
nand U42491 (N_42491,N_40346,N_41205);
nand U42492 (N_42492,N_40246,N_40148);
nor U42493 (N_42493,N_41785,N_41023);
nand U42494 (N_42494,N_40283,N_41389);
and U42495 (N_42495,N_40858,N_41782);
xor U42496 (N_42496,N_40992,N_41599);
or U42497 (N_42497,N_40130,N_41904);
nand U42498 (N_42498,N_41900,N_40142);
nor U42499 (N_42499,N_40440,N_41899);
nor U42500 (N_42500,N_40707,N_41412);
nand U42501 (N_42501,N_40428,N_41571);
nand U42502 (N_42502,N_40717,N_40843);
and U42503 (N_42503,N_40617,N_41996);
and U42504 (N_42504,N_40954,N_41475);
and U42505 (N_42505,N_41379,N_40719);
xnor U42506 (N_42506,N_41052,N_40155);
nand U42507 (N_42507,N_41080,N_41720);
and U42508 (N_42508,N_40226,N_41682);
nor U42509 (N_42509,N_40664,N_41376);
nand U42510 (N_42510,N_40894,N_40389);
nor U42511 (N_42511,N_41137,N_41343);
and U42512 (N_42512,N_40491,N_40885);
or U42513 (N_42513,N_41275,N_41204);
xnor U42514 (N_42514,N_41555,N_41795);
nor U42515 (N_42515,N_40524,N_40568);
xnor U42516 (N_42516,N_41973,N_41837);
xnor U42517 (N_42517,N_40692,N_40349);
or U42518 (N_42518,N_40088,N_41731);
and U42519 (N_42519,N_40178,N_40198);
nor U42520 (N_42520,N_41333,N_40676);
or U42521 (N_42521,N_41807,N_40964);
and U42522 (N_42522,N_40071,N_40347);
nand U42523 (N_42523,N_40584,N_41338);
and U42524 (N_42524,N_41926,N_40445);
xnor U42525 (N_42525,N_40087,N_41446);
and U42526 (N_42526,N_40718,N_40442);
nand U42527 (N_42527,N_40877,N_41594);
nor U42528 (N_42528,N_40732,N_41285);
xnor U42529 (N_42529,N_41399,N_41071);
nor U42530 (N_42530,N_40567,N_40197);
nor U42531 (N_42531,N_40202,N_40533);
or U42532 (N_42532,N_40786,N_40393);
or U42533 (N_42533,N_40553,N_41062);
nor U42534 (N_42534,N_40028,N_41662);
and U42535 (N_42535,N_41915,N_40713);
nor U42536 (N_42536,N_40145,N_40696);
nor U42537 (N_42537,N_40675,N_41307);
nor U42538 (N_42538,N_40308,N_41597);
and U42539 (N_42539,N_41652,N_41117);
or U42540 (N_42540,N_40011,N_40986);
nand U42541 (N_42541,N_41824,N_40132);
or U42542 (N_42542,N_40117,N_41569);
xnor U42543 (N_42543,N_40465,N_41801);
nor U42544 (N_42544,N_40059,N_41618);
or U42545 (N_42545,N_41686,N_40296);
and U42546 (N_42546,N_40478,N_40629);
or U42547 (N_42547,N_41431,N_40139);
or U42548 (N_42548,N_41621,N_41762);
or U42549 (N_42549,N_41321,N_40135);
or U42550 (N_42550,N_41557,N_40637);
nand U42551 (N_42551,N_40895,N_40042);
xnor U42552 (N_42552,N_41978,N_41169);
and U42553 (N_42553,N_41352,N_41629);
and U42554 (N_42554,N_40905,N_41100);
and U42555 (N_42555,N_41828,N_41967);
and U42556 (N_42556,N_41051,N_40840);
and U42557 (N_42557,N_40289,N_41407);
nand U42558 (N_42558,N_40830,N_41786);
xor U42559 (N_42559,N_40593,N_41580);
xor U42560 (N_42560,N_40686,N_41752);
or U42561 (N_42561,N_41185,N_41870);
nor U42562 (N_42562,N_40089,N_40056);
nand U42563 (N_42563,N_41989,N_40123);
nor U42564 (N_42564,N_41578,N_41090);
and U42565 (N_42565,N_41250,N_40391);
and U42566 (N_42566,N_41753,N_40002);
or U42567 (N_42567,N_40200,N_41684);
or U42568 (N_42568,N_40143,N_40260);
xor U42569 (N_42569,N_41942,N_40220);
or U42570 (N_42570,N_41069,N_41263);
nand U42571 (N_42571,N_40774,N_40433);
xor U42572 (N_42572,N_41076,N_41685);
nand U42573 (N_42573,N_40460,N_40681);
or U42574 (N_42574,N_40336,N_41432);
nor U42575 (N_42575,N_41146,N_40472);
and U42576 (N_42576,N_40716,N_41642);
nand U42577 (N_42577,N_40338,N_41606);
nand U42578 (N_42578,N_40690,N_41068);
or U42579 (N_42579,N_40288,N_41588);
xor U42580 (N_42580,N_40790,N_41118);
xor U42581 (N_42581,N_40525,N_41276);
nand U42582 (N_42582,N_40252,N_41743);
and U42583 (N_42583,N_41419,N_41000);
or U42584 (N_42584,N_41640,N_40069);
xnor U42585 (N_42585,N_40851,N_41334);
nand U42586 (N_42586,N_41914,N_40741);
nor U42587 (N_42587,N_41700,N_41004);
or U42588 (N_42588,N_41797,N_40113);
nand U42589 (N_42589,N_41358,N_41264);
or U42590 (N_42590,N_41489,N_40807);
or U42591 (N_42591,N_40674,N_41519);
xnor U42592 (N_42592,N_40195,N_40242);
nor U42593 (N_42593,N_40209,N_41584);
nor U42594 (N_42594,N_41655,N_41948);
nand U42595 (N_42595,N_41833,N_40141);
and U42596 (N_42596,N_41371,N_40556);
or U42597 (N_42597,N_41305,N_40150);
or U42598 (N_42598,N_40214,N_41420);
or U42599 (N_42599,N_40151,N_41669);
and U42600 (N_42600,N_40983,N_40947);
or U42601 (N_42601,N_40749,N_40121);
or U42602 (N_42602,N_40264,N_40819);
xnor U42603 (N_42603,N_41122,N_40396);
xor U42604 (N_42604,N_41951,N_41719);
and U42605 (N_42605,N_41317,N_40235);
nand U42606 (N_42606,N_41656,N_40228);
nand U42607 (N_42607,N_41630,N_40619);
xor U42608 (N_42608,N_41328,N_41733);
xnor U42609 (N_42609,N_41219,N_40482);
nand U42610 (N_42610,N_41757,N_40173);
and U42611 (N_42611,N_40489,N_40551);
or U42612 (N_42612,N_41466,N_41495);
nand U42613 (N_42613,N_41770,N_40023);
nor U42614 (N_42614,N_40475,N_41610);
xnor U42615 (N_42615,N_41082,N_40628);
nor U42616 (N_42616,N_41626,N_40502);
and U42617 (N_42617,N_40506,N_40486);
nor U42618 (N_42618,N_41460,N_40434);
or U42619 (N_42619,N_41559,N_40514);
and U42620 (N_42620,N_40995,N_41444);
or U42621 (N_42621,N_40891,N_41113);
and U42622 (N_42622,N_40569,N_41943);
xor U42623 (N_42623,N_40128,N_41034);
or U42624 (N_42624,N_41110,N_41315);
xnor U42625 (N_42625,N_40796,N_41054);
nor U42626 (N_42626,N_40956,N_41401);
xnor U42627 (N_42627,N_41229,N_40206);
nor U42628 (N_42628,N_41890,N_41445);
or U42629 (N_42629,N_41747,N_40862);
nor U42630 (N_42630,N_40029,N_41643);
or U42631 (N_42631,N_41397,N_41298);
nor U42632 (N_42632,N_41279,N_40778);
nor U42633 (N_42633,N_40147,N_40767);
nor U42634 (N_42634,N_40708,N_41676);
xnor U42635 (N_42635,N_41295,N_41696);
nand U42636 (N_42636,N_41498,N_40899);
nand U42637 (N_42637,N_41391,N_41429);
and U42638 (N_42638,N_40880,N_40847);
and U42639 (N_42639,N_41641,N_41945);
nor U42640 (N_42640,N_41805,N_41156);
and U42641 (N_42641,N_41368,N_41694);
nor U42642 (N_42642,N_41970,N_41575);
or U42643 (N_42643,N_40698,N_40638);
xor U42644 (N_42644,N_41454,N_41157);
xor U42645 (N_42645,N_41955,N_40901);
nand U42646 (N_42646,N_40484,N_40319);
nand U42647 (N_42647,N_40682,N_40627);
nand U42648 (N_42648,N_40378,N_40928);
and U42649 (N_42649,N_40884,N_40044);
nor U42650 (N_42650,N_40754,N_41953);
nor U42651 (N_42651,N_40297,N_40179);
or U42652 (N_42652,N_40342,N_40233);
and U42653 (N_42653,N_41627,N_41152);
nor U42654 (N_42654,N_41361,N_41657);
and U42655 (N_42655,N_40070,N_41006);
nor U42656 (N_42656,N_40701,N_40623);
nor U42657 (N_42657,N_40411,N_40922);
xor U42658 (N_42658,N_40303,N_40328);
nand U42659 (N_42659,N_40320,N_40955);
xnor U42660 (N_42660,N_41804,N_40374);
nor U42661 (N_42661,N_40355,N_40835);
xnor U42662 (N_42662,N_41672,N_41667);
nand U42663 (N_42663,N_41270,N_40454);
nand U42664 (N_42664,N_41387,N_41698);
nor U42665 (N_42665,N_40407,N_41362);
xor U42666 (N_42666,N_40496,N_40634);
nand U42667 (N_42667,N_41378,N_41021);
nor U42668 (N_42668,N_40205,N_40838);
xor U42669 (N_42669,N_41260,N_40609);
nand U42670 (N_42670,N_40898,N_41882);
nand U42671 (N_42671,N_41798,N_40278);
nand U42672 (N_42672,N_40507,N_41308);
nand U42673 (N_42673,N_41547,N_41631);
nor U42674 (N_42674,N_40431,N_41518);
or U42675 (N_42675,N_40326,N_40118);
or U42676 (N_42676,N_41661,N_40577);
nor U42677 (N_42677,N_40988,N_40127);
and U42678 (N_42678,N_41231,N_40881);
nand U42679 (N_42679,N_40759,N_41859);
or U42680 (N_42680,N_40644,N_41885);
xor U42681 (N_42681,N_41653,N_40109);
nor U42682 (N_42682,N_41318,N_41614);
and U42683 (N_42683,N_41492,N_40307);
nand U42684 (N_42684,N_40869,N_40318);
nor U42685 (N_42685,N_40285,N_41324);
xor U42686 (N_42686,N_40772,N_40691);
nor U42687 (N_42687,N_40592,N_40522);
or U42688 (N_42688,N_41918,N_40633);
and U42689 (N_42689,N_40394,N_40545);
and U42690 (N_42690,N_41834,N_41919);
xnor U42691 (N_42691,N_40240,N_41128);
or U42692 (N_42692,N_40921,N_40287);
xnor U42693 (N_42693,N_40176,N_40788);
xor U42694 (N_42694,N_40631,N_41411);
or U42695 (N_42695,N_41744,N_40090);
and U42696 (N_42696,N_40854,N_40805);
nand U42697 (N_42697,N_40357,N_40321);
or U42698 (N_42698,N_40993,N_41421);
and U42699 (N_42699,N_41200,N_40534);
and U42700 (N_42700,N_40511,N_40892);
xnor U42701 (N_42701,N_40305,N_40977);
nor U42702 (N_42702,N_41705,N_41046);
or U42703 (N_42703,N_40439,N_40722);
or U42704 (N_42704,N_40000,N_40876);
xnor U42705 (N_42705,N_40263,N_41032);
or U42706 (N_42706,N_41668,N_41234);
nand U42707 (N_42707,N_40923,N_41148);
nand U42708 (N_42708,N_41842,N_40426);
nand U42709 (N_42709,N_40366,N_41277);
xnor U42710 (N_42710,N_40930,N_40257);
and U42711 (N_42711,N_40159,N_40085);
xor U42712 (N_42712,N_41658,N_40466);
nor U42713 (N_42713,N_40720,N_40036);
nand U42714 (N_42714,N_41542,N_41290);
or U42715 (N_42715,N_40808,N_40051);
xor U42716 (N_42716,N_40888,N_40813);
nor U42717 (N_42717,N_40247,N_41774);
or U42718 (N_42718,N_41094,N_41126);
and U42719 (N_42719,N_40706,N_41922);
or U42720 (N_42720,N_41413,N_40783);
or U42721 (N_42721,N_41213,N_41210);
and U42722 (N_42722,N_40277,N_41718);
nor U42723 (N_42723,N_41476,N_40004);
nand U42724 (N_42724,N_41759,N_41424);
or U42725 (N_42725,N_40604,N_40017);
or U42726 (N_42726,N_41840,N_41623);
and U42727 (N_42727,N_41808,N_41039);
and U42728 (N_42728,N_41230,N_40306);
nand U42729 (N_42729,N_40186,N_41988);
nor U42730 (N_42730,N_40180,N_41486);
nor U42731 (N_42731,N_41035,N_40541);
xor U42732 (N_42732,N_40615,N_40973);
nand U42733 (N_42733,N_40924,N_40007);
nor U42734 (N_42734,N_41306,N_41367);
or U42735 (N_42735,N_41565,N_40162);
nor U42736 (N_42736,N_41353,N_41297);
xor U42737 (N_42737,N_41939,N_41252);
xnor U42738 (N_42738,N_41423,N_41971);
nor U42739 (N_42739,N_41691,N_41844);
nand U42740 (N_42740,N_40744,N_41249);
or U42741 (N_42741,N_41566,N_41855);
and U42742 (N_42742,N_41151,N_40022);
and U42743 (N_42743,N_40868,N_41969);
or U42744 (N_42744,N_41984,N_41716);
xnor U42745 (N_42745,N_40859,N_41539);
xnor U42746 (N_42746,N_41134,N_41355);
nand U42747 (N_42747,N_40563,N_40470);
xor U42748 (N_42748,N_40758,N_41677);
nor U42749 (N_42749,N_40697,N_41507);
nand U42750 (N_42750,N_40611,N_40547);
nor U42751 (N_42751,N_41671,N_40194);
nor U42752 (N_42752,N_41045,N_41835);
and U42753 (N_42753,N_41440,N_41763);
nor U42754 (N_42754,N_40034,N_41472);
nand U42755 (N_42755,N_41335,N_40447);
and U42756 (N_42756,N_40576,N_40414);
nand U42757 (N_42757,N_40845,N_40292);
xnor U42758 (N_42758,N_41265,N_40154);
xor U42759 (N_42759,N_41756,N_41098);
nor U42760 (N_42760,N_40530,N_40463);
and U42761 (N_42761,N_41892,N_41074);
nand U42762 (N_42762,N_40662,N_41754);
nand U42763 (N_42763,N_40669,N_40025);
xor U42764 (N_42764,N_41405,N_40519);
or U42765 (N_42765,N_40152,N_40855);
and U42766 (N_42766,N_40282,N_41251);
or U42767 (N_42767,N_41839,N_40595);
nand U42768 (N_42768,N_40485,N_40574);
nand U42769 (N_42769,N_41040,N_40912);
nand U42770 (N_42770,N_41871,N_41060);
nand U42771 (N_42771,N_40170,N_40982);
or U42772 (N_42772,N_41898,N_40322);
or U42773 (N_42773,N_40457,N_40144);
or U42774 (N_42774,N_40666,N_41125);
nor U42775 (N_42775,N_40390,N_41061);
nor U42776 (N_42776,N_41866,N_40756);
xor U42777 (N_42777,N_41102,N_41450);
nor U42778 (N_42778,N_41400,N_40588);
xor U42779 (N_42779,N_41273,N_40689);
nor U42780 (N_42780,N_41281,N_40887);
nor U42781 (N_42781,N_40771,N_41587);
nor U42782 (N_42782,N_40656,N_41465);
nand U42783 (N_42783,N_41589,N_40616);
nand U42784 (N_42784,N_40809,N_40487);
nand U42785 (N_42785,N_41941,N_40909);
and U42786 (N_42786,N_40999,N_40094);
nor U42787 (N_42787,N_41713,N_41777);
xnor U42788 (N_42788,N_40480,N_41171);
or U42789 (N_42789,N_40531,N_41167);
xnor U42790 (N_42790,N_40510,N_40981);
nor U42791 (N_42791,N_41160,N_40823);
nand U42792 (N_42792,N_40477,N_41209);
nor U42793 (N_42793,N_41745,N_41187);
or U42794 (N_42794,N_40904,N_40658);
or U42795 (N_42795,N_40677,N_40738);
nor U42796 (N_42796,N_41510,N_40618);
nor U42797 (N_42797,N_41072,N_41214);
nor U42798 (N_42798,N_41579,N_40509);
xnor U42799 (N_42799,N_40561,N_41827);
xor U42800 (N_42800,N_41529,N_40607);
and U42801 (N_42801,N_41616,N_41875);
or U42802 (N_42802,N_41937,N_40659);
nand U42803 (N_42803,N_40991,N_40356);
and U42804 (N_42804,N_41769,N_40651);
nor U42805 (N_42805,N_41049,N_40685);
xor U42806 (N_42806,N_41985,N_40605);
and U42807 (N_42807,N_41789,N_41129);
nor U42808 (N_42808,N_40016,N_40251);
or U42809 (N_42809,N_41549,N_41832);
nor U42810 (N_42810,N_41114,N_41196);
nand U42811 (N_42811,N_41911,N_40099);
xor U42812 (N_42812,N_40471,N_41504);
xnor U42813 (N_42813,N_41439,N_40972);
nand U42814 (N_42814,N_41154,N_40286);
nor U42815 (N_42815,N_41586,N_41254);
nor U42816 (N_42816,N_41954,N_41525);
xnor U42817 (N_42817,N_41665,N_40175);
and U42818 (N_42818,N_40354,N_41862);
xor U42819 (N_42819,N_40419,N_40730);
nand U42820 (N_42820,N_40337,N_40906);
nor U42821 (N_42821,N_41893,N_40435);
or U42822 (N_42822,N_41059,N_40558);
or U42823 (N_42823,N_41613,N_40073);
or U42824 (N_42824,N_40550,N_40989);
or U42825 (N_42825,N_40976,N_41615);
and U42826 (N_42826,N_40430,N_40136);
xnor U42827 (N_42827,N_40481,N_40212);
or U42828 (N_42828,N_40802,N_41816);
nand U42829 (N_42829,N_41274,N_40064);
or U42830 (N_42830,N_40815,N_40097);
nand U42831 (N_42831,N_40606,N_40821);
nand U42832 (N_42832,N_40990,N_40874);
or U42833 (N_42833,N_41849,N_41593);
xnor U42834 (N_42834,N_40362,N_40473);
xor U42835 (N_42835,N_40024,N_41235);
and U42836 (N_42836,N_41949,N_41617);
xor U42837 (N_42837,N_41096,N_40273);
nor U42838 (N_42838,N_40770,N_40232);
or U42839 (N_42839,N_40453,N_40400);
nand U42840 (N_42840,N_41585,N_40560);
nand U42841 (N_42841,N_40304,N_40076);
or U42842 (N_42842,N_41598,N_41042);
or U42843 (N_42843,N_41809,N_41053);
nor U42844 (N_42844,N_41192,N_41897);
and U42845 (N_42845,N_40784,N_40748);
nand U42846 (N_42846,N_41771,N_40959);
xor U42847 (N_42847,N_41869,N_40914);
and U42848 (N_42848,N_40672,N_40266);
or U42849 (N_42849,N_40647,N_41178);
xor U42850 (N_42850,N_40834,N_40559);
or U42851 (N_42851,N_40614,N_41577);
and U42852 (N_42852,N_40413,N_41394);
or U42853 (N_42853,N_40557,N_40937);
nor U42854 (N_42854,N_41993,N_40153);
nor U42855 (N_42855,N_41020,N_41483);
and U42856 (N_42856,N_40361,N_40866);
xnor U42857 (N_42857,N_41191,N_41521);
xor U42858 (N_42858,N_41933,N_41628);
nor U42859 (N_42859,N_41938,N_41517);
and U42860 (N_42860,N_41121,N_40863);
nand U42861 (N_42861,N_41831,N_41727);
xor U42862 (N_42862,N_41787,N_41408);
nand U42863 (N_42863,N_41218,N_40542);
xnor U42864 (N_42864,N_40733,N_41959);
xnor U42865 (N_42865,N_40640,N_41863);
and U42866 (N_42866,N_41944,N_40596);
or U42867 (N_42867,N_40190,N_41159);
and U42868 (N_42868,N_40401,N_41136);
and U42869 (N_42869,N_40985,N_40483);
or U42870 (N_42870,N_41293,N_41199);
nor U42871 (N_42871,N_41083,N_40900);
xor U42872 (N_42872,N_41961,N_41145);
nor U42873 (N_42873,N_40649,N_41262);
nand U42874 (N_42874,N_41153,N_40262);
xnor U42875 (N_42875,N_40219,N_40711);
or U42876 (N_42876,N_40782,N_41189);
nand U42877 (N_42877,N_40648,N_41925);
nor U42878 (N_42878,N_41540,N_40239);
nor U42879 (N_42879,N_41261,N_41280);
or U42880 (N_42880,N_40270,N_41921);
xnor U42881 (N_42881,N_41422,N_40184);
nand U42882 (N_42882,N_41381,N_40826);
nor U42883 (N_42883,N_40883,N_41373);
xor U42884 (N_42884,N_40302,N_40343);
or U42885 (N_42885,N_40340,N_40518);
xor U42886 (N_42886,N_40015,N_41534);
xor U42887 (N_42887,N_41067,N_41172);
and U42888 (N_42888,N_40369,N_40224);
or U42889 (N_42889,N_41940,N_41365);
nor U42890 (N_42890,N_41646,N_40610);
and U42891 (N_42891,N_40416,N_41856);
or U42892 (N_42892,N_41143,N_40185);
or U42893 (N_42893,N_40837,N_41509);
or U42894 (N_42894,N_40276,N_40861);
and U42895 (N_42895,N_40630,N_41935);
xnor U42896 (N_42896,N_40661,N_40373);
nor U42897 (N_42897,N_40798,N_40839);
nand U42898 (N_42898,N_40503,N_41133);
nor U42899 (N_42899,N_40725,N_40458);
xor U42900 (N_42900,N_41184,N_40375);
or U42901 (N_42901,N_40474,N_40367);
or U42902 (N_42902,N_41312,N_41474);
nor U42903 (N_42903,N_40703,N_41140);
nand U42904 (N_42904,N_40768,N_40300);
xnor U42905 (N_42905,N_40979,N_41232);
xnor U42906 (N_42906,N_41370,N_41734);
and U42907 (N_42907,N_41979,N_40836);
and U42908 (N_42908,N_41632,N_41603);
and U42909 (N_42909,N_41619,N_40832);
and U42910 (N_42910,N_41319,N_40852);
xor U42911 (N_42911,N_40678,N_40673);
and U42912 (N_42912,N_41220,N_40259);
nand U42913 (N_42913,N_40950,N_40098);
and U42914 (N_42914,N_41164,N_41773);
xnor U42915 (N_42915,N_41001,N_41223);
nand U42916 (N_42916,N_40571,N_41567);
and U42917 (N_42917,N_41848,N_40429);
nand U42918 (N_42918,N_41767,N_40187);
xor U42919 (N_42919,N_40380,N_40915);
and U42920 (N_42920,N_41467,N_41168);
and U42921 (N_42921,N_40565,N_41910);
nor U42922 (N_42922,N_40801,N_41409);
nand U42923 (N_42923,N_41289,N_41583);
and U42924 (N_42924,N_40058,N_41950);
nand U42925 (N_42925,N_41788,N_41016);
and U42926 (N_42926,N_40941,N_40694);
or U42927 (N_42927,N_41471,N_40105);
xor U42928 (N_42928,N_40643,N_41327);
or U42929 (N_42929,N_41896,N_41895);
nor U42930 (N_42930,N_41710,N_41553);
and U42931 (N_42931,N_41208,N_41024);
nor U42932 (N_42932,N_41416,N_40216);
xor U42933 (N_42933,N_40965,N_40327);
xor U42934 (N_42934,N_40157,N_41592);
nand U42935 (N_42935,N_41902,N_41838);
nor U42936 (N_42936,N_41524,N_41177);
or U42937 (N_42937,N_41548,N_41107);
and U42938 (N_42938,N_40594,N_41546);
nand U42939 (N_42939,N_40425,N_41403);
nor U42940 (N_42940,N_40382,N_41814);
or U42941 (N_42941,N_41120,N_41050);
and U42942 (N_42942,N_41175,N_40820);
or U42943 (N_42943,N_41772,N_41846);
or U42944 (N_42944,N_41441,N_41302);
and U42945 (N_42945,N_41019,N_41104);
nor U42946 (N_42946,N_40488,N_41288);
or U42947 (N_42947,N_40498,N_41821);
nand U42948 (N_42948,N_41867,N_40467);
nand U42949 (N_42949,N_40096,N_41036);
nand U42950 (N_42950,N_40168,N_41748);
xor U42951 (N_42951,N_41637,N_41033);
xnor U42952 (N_42952,N_41551,N_40352);
or U42953 (N_42953,N_40671,N_41163);
and U42954 (N_42954,N_40546,N_40199);
xor U42955 (N_42955,N_40726,N_40415);
nor U42956 (N_42956,N_40963,N_41533);
nor U42957 (N_42957,N_40421,N_41887);
nor U42958 (N_42958,N_40817,N_41022);
nor U42959 (N_42959,N_41119,N_41079);
and U42960 (N_42960,N_41253,N_40041);
or U42961 (N_42961,N_40761,N_41296);
or U42962 (N_42962,N_41346,N_41877);
nand U42963 (N_42963,N_41934,N_40033);
nand U42964 (N_42964,N_40410,N_41550);
or U42965 (N_42965,N_40323,N_41197);
or U42966 (N_42966,N_40857,N_40217);
and U42967 (N_42967,N_40398,N_40188);
xor U42968 (N_42968,N_41025,N_41729);
or U42969 (N_42969,N_41608,N_41345);
xor U42970 (N_42970,N_41491,N_40045);
and U42971 (N_42971,N_40508,N_41225);
and U42972 (N_42972,N_41008,N_41438);
or U42973 (N_42973,N_40114,N_41711);
nand U42974 (N_42974,N_41089,N_40497);
and U42975 (N_42975,N_41449,N_41803);
xor U42976 (N_42976,N_40548,N_41162);
and U42977 (N_42977,N_40920,N_41149);
nor U42978 (N_42978,N_40317,N_40968);
or U42979 (N_42979,N_40469,N_40241);
xor U42980 (N_42980,N_40417,N_40727);
or U42981 (N_42981,N_40054,N_41601);
and U42982 (N_42982,N_41086,N_40108);
and U42983 (N_42983,N_41714,N_41088);
or U42984 (N_42984,N_40095,N_40100);
xnor U42985 (N_42985,N_41800,N_40544);
or U42986 (N_42986,N_40620,N_41142);
xnor U42987 (N_42987,N_40208,N_40564);
nor U42988 (N_42988,N_41620,N_40351);
xnor U42989 (N_42989,N_40043,N_40517);
nand U42990 (N_42990,N_41680,N_41174);
and U42991 (N_42991,N_41243,N_41227);
or U42992 (N_42992,N_41622,N_41732);
and U42993 (N_42993,N_41103,N_41242);
xor U42994 (N_42994,N_40804,N_40455);
xnor U42995 (N_42995,N_41947,N_40555);
and U42996 (N_42996,N_41878,N_40636);
and U42997 (N_42997,N_41701,N_40329);
and U42998 (N_42998,N_40032,N_40107);
nand U42999 (N_42999,N_41170,N_41215);
or U43000 (N_43000,N_40825,N_41198);
nor U43001 (N_43001,N_40234,N_40861);
and U43002 (N_43002,N_41396,N_41046);
and U43003 (N_43003,N_40370,N_41155);
and U43004 (N_43004,N_41084,N_40246);
or U43005 (N_43005,N_41456,N_40994);
nand U43006 (N_43006,N_40057,N_41440);
and U43007 (N_43007,N_40198,N_41466);
nand U43008 (N_43008,N_40491,N_40657);
xor U43009 (N_43009,N_41391,N_41244);
nand U43010 (N_43010,N_40448,N_40479);
and U43011 (N_43011,N_41175,N_40313);
xor U43012 (N_43012,N_40058,N_41255);
or U43013 (N_43013,N_41313,N_41532);
xnor U43014 (N_43014,N_40979,N_40372);
nand U43015 (N_43015,N_40576,N_40755);
xor U43016 (N_43016,N_41117,N_41063);
nand U43017 (N_43017,N_41415,N_41284);
nor U43018 (N_43018,N_41982,N_40878);
nand U43019 (N_43019,N_40123,N_40335);
nor U43020 (N_43020,N_41323,N_41745);
and U43021 (N_43021,N_40073,N_41534);
xnor U43022 (N_43022,N_41027,N_41485);
xor U43023 (N_43023,N_40961,N_41665);
nor U43024 (N_43024,N_41616,N_41361);
and U43025 (N_43025,N_41159,N_40407);
and U43026 (N_43026,N_41800,N_41249);
xnor U43027 (N_43027,N_41835,N_40925);
and U43028 (N_43028,N_41656,N_40616);
xor U43029 (N_43029,N_40627,N_40713);
nand U43030 (N_43030,N_40971,N_40241);
nor U43031 (N_43031,N_40028,N_41407);
nand U43032 (N_43032,N_40369,N_41171);
or U43033 (N_43033,N_40590,N_41726);
or U43034 (N_43034,N_40414,N_41842);
and U43035 (N_43035,N_41124,N_41967);
nand U43036 (N_43036,N_41232,N_40001);
and U43037 (N_43037,N_40016,N_40657);
nor U43038 (N_43038,N_40686,N_40293);
nor U43039 (N_43039,N_40540,N_40285);
nor U43040 (N_43040,N_40307,N_41794);
or U43041 (N_43041,N_41511,N_40647);
xor U43042 (N_43042,N_41872,N_41704);
nand U43043 (N_43043,N_41309,N_41050);
xnor U43044 (N_43044,N_40575,N_41796);
nor U43045 (N_43045,N_41258,N_40861);
or U43046 (N_43046,N_41593,N_41690);
nand U43047 (N_43047,N_40294,N_41409);
or U43048 (N_43048,N_40385,N_40951);
nor U43049 (N_43049,N_40836,N_41690);
or U43050 (N_43050,N_40798,N_40343);
and U43051 (N_43051,N_40279,N_41759);
nor U43052 (N_43052,N_40639,N_40519);
nor U43053 (N_43053,N_41044,N_41377);
nor U43054 (N_43054,N_41630,N_40494);
and U43055 (N_43055,N_40000,N_40172);
nand U43056 (N_43056,N_40085,N_41034);
and U43057 (N_43057,N_40116,N_41550);
nand U43058 (N_43058,N_41569,N_40576);
and U43059 (N_43059,N_40531,N_41236);
nand U43060 (N_43060,N_40477,N_41557);
and U43061 (N_43061,N_41352,N_40295);
or U43062 (N_43062,N_41562,N_40228);
or U43063 (N_43063,N_40561,N_41677);
or U43064 (N_43064,N_41138,N_41122);
and U43065 (N_43065,N_41484,N_40178);
nand U43066 (N_43066,N_40719,N_41607);
nor U43067 (N_43067,N_40446,N_41230);
and U43068 (N_43068,N_40692,N_41808);
or U43069 (N_43069,N_40004,N_40472);
nor U43070 (N_43070,N_41295,N_41561);
nor U43071 (N_43071,N_40897,N_41741);
and U43072 (N_43072,N_41531,N_41252);
nor U43073 (N_43073,N_41161,N_41866);
xnor U43074 (N_43074,N_41863,N_41987);
nand U43075 (N_43075,N_40851,N_40237);
nor U43076 (N_43076,N_40763,N_40488);
nor U43077 (N_43077,N_40489,N_41352);
nand U43078 (N_43078,N_41217,N_41730);
xor U43079 (N_43079,N_40409,N_41473);
nand U43080 (N_43080,N_41712,N_41919);
xnor U43081 (N_43081,N_41629,N_41386);
nand U43082 (N_43082,N_40468,N_41883);
nor U43083 (N_43083,N_40782,N_41770);
nand U43084 (N_43084,N_41580,N_40530);
nand U43085 (N_43085,N_40628,N_41206);
or U43086 (N_43086,N_40374,N_40649);
or U43087 (N_43087,N_40373,N_40348);
xor U43088 (N_43088,N_41892,N_41676);
nor U43089 (N_43089,N_41960,N_41605);
or U43090 (N_43090,N_41546,N_41297);
or U43091 (N_43091,N_41891,N_40813);
nand U43092 (N_43092,N_41054,N_41630);
nor U43093 (N_43093,N_40646,N_41051);
xnor U43094 (N_43094,N_40333,N_40913);
xor U43095 (N_43095,N_40989,N_40875);
xnor U43096 (N_43096,N_41335,N_41256);
nor U43097 (N_43097,N_41344,N_40502);
or U43098 (N_43098,N_40773,N_41352);
xnor U43099 (N_43099,N_41590,N_40686);
and U43100 (N_43100,N_40726,N_40023);
and U43101 (N_43101,N_41123,N_40519);
nor U43102 (N_43102,N_41348,N_40500);
or U43103 (N_43103,N_41013,N_41371);
nor U43104 (N_43104,N_41893,N_40067);
or U43105 (N_43105,N_40308,N_40218);
or U43106 (N_43106,N_40678,N_41837);
nor U43107 (N_43107,N_40820,N_40741);
or U43108 (N_43108,N_41539,N_40984);
and U43109 (N_43109,N_41626,N_40913);
or U43110 (N_43110,N_41977,N_40263);
nand U43111 (N_43111,N_41454,N_40885);
nand U43112 (N_43112,N_40102,N_41349);
nor U43113 (N_43113,N_40665,N_40007);
or U43114 (N_43114,N_41459,N_40075);
xnor U43115 (N_43115,N_40732,N_41556);
or U43116 (N_43116,N_41469,N_41891);
and U43117 (N_43117,N_41324,N_40766);
nor U43118 (N_43118,N_41799,N_40666);
xor U43119 (N_43119,N_41165,N_40615);
nor U43120 (N_43120,N_40884,N_41070);
nand U43121 (N_43121,N_40636,N_41654);
and U43122 (N_43122,N_41648,N_40268);
xor U43123 (N_43123,N_40655,N_41074);
and U43124 (N_43124,N_40141,N_40094);
xnor U43125 (N_43125,N_40261,N_41713);
nor U43126 (N_43126,N_40259,N_40352);
and U43127 (N_43127,N_40506,N_41954);
nand U43128 (N_43128,N_41916,N_40196);
xor U43129 (N_43129,N_40773,N_40069);
or U43130 (N_43130,N_40048,N_41601);
nor U43131 (N_43131,N_40933,N_40132);
or U43132 (N_43132,N_41819,N_41592);
and U43133 (N_43133,N_41981,N_40256);
and U43134 (N_43134,N_41798,N_41575);
xnor U43135 (N_43135,N_40040,N_40937);
nand U43136 (N_43136,N_41979,N_41602);
nand U43137 (N_43137,N_41444,N_40259);
nand U43138 (N_43138,N_41713,N_41528);
or U43139 (N_43139,N_41901,N_40538);
nand U43140 (N_43140,N_41569,N_41549);
xnor U43141 (N_43141,N_41085,N_41431);
xor U43142 (N_43142,N_41962,N_40571);
and U43143 (N_43143,N_40423,N_41368);
or U43144 (N_43144,N_40038,N_41503);
nand U43145 (N_43145,N_41321,N_40857);
or U43146 (N_43146,N_41218,N_40696);
xnor U43147 (N_43147,N_40120,N_41214);
xor U43148 (N_43148,N_41744,N_41153);
xnor U43149 (N_43149,N_41279,N_40886);
nand U43150 (N_43150,N_41578,N_41504);
nor U43151 (N_43151,N_40211,N_41505);
or U43152 (N_43152,N_41619,N_40470);
xor U43153 (N_43153,N_40472,N_40026);
and U43154 (N_43154,N_40632,N_41799);
and U43155 (N_43155,N_40817,N_41586);
xnor U43156 (N_43156,N_41301,N_40773);
nor U43157 (N_43157,N_41620,N_41109);
and U43158 (N_43158,N_40306,N_40376);
nand U43159 (N_43159,N_41894,N_41419);
nor U43160 (N_43160,N_41131,N_40161);
nand U43161 (N_43161,N_40272,N_40370);
or U43162 (N_43162,N_41682,N_40978);
nand U43163 (N_43163,N_40440,N_41783);
nor U43164 (N_43164,N_41858,N_40997);
nor U43165 (N_43165,N_41745,N_40213);
and U43166 (N_43166,N_41877,N_41305);
xnor U43167 (N_43167,N_41805,N_41303);
and U43168 (N_43168,N_40222,N_41787);
and U43169 (N_43169,N_41620,N_41092);
nor U43170 (N_43170,N_41853,N_40416);
or U43171 (N_43171,N_40004,N_40100);
and U43172 (N_43172,N_40534,N_40457);
or U43173 (N_43173,N_41174,N_40543);
and U43174 (N_43174,N_41570,N_40036);
or U43175 (N_43175,N_40812,N_40157);
nand U43176 (N_43176,N_40319,N_41796);
and U43177 (N_43177,N_41276,N_41560);
and U43178 (N_43178,N_41712,N_41529);
and U43179 (N_43179,N_41337,N_40096);
and U43180 (N_43180,N_40916,N_40443);
nor U43181 (N_43181,N_41808,N_41724);
or U43182 (N_43182,N_41089,N_40004);
and U43183 (N_43183,N_40548,N_40241);
nand U43184 (N_43184,N_40451,N_41389);
and U43185 (N_43185,N_41931,N_41537);
xnor U43186 (N_43186,N_41294,N_41064);
and U43187 (N_43187,N_40571,N_40237);
or U43188 (N_43188,N_41193,N_41771);
or U43189 (N_43189,N_41205,N_40188);
or U43190 (N_43190,N_41062,N_41382);
or U43191 (N_43191,N_41456,N_41106);
or U43192 (N_43192,N_41129,N_41100);
nor U43193 (N_43193,N_41435,N_41077);
nor U43194 (N_43194,N_40090,N_41571);
or U43195 (N_43195,N_40765,N_40836);
and U43196 (N_43196,N_41855,N_40289);
nor U43197 (N_43197,N_40940,N_40245);
and U43198 (N_43198,N_40169,N_41634);
xnor U43199 (N_43199,N_40473,N_41657);
xor U43200 (N_43200,N_40042,N_40198);
nand U43201 (N_43201,N_40284,N_40922);
nor U43202 (N_43202,N_41086,N_41432);
xor U43203 (N_43203,N_40209,N_40597);
nand U43204 (N_43204,N_40395,N_41745);
xnor U43205 (N_43205,N_41131,N_41722);
xnor U43206 (N_43206,N_40713,N_40691);
nor U43207 (N_43207,N_41077,N_40741);
nor U43208 (N_43208,N_41501,N_40687);
or U43209 (N_43209,N_40580,N_41060);
or U43210 (N_43210,N_40762,N_40230);
xor U43211 (N_43211,N_40524,N_41392);
and U43212 (N_43212,N_41940,N_41033);
nor U43213 (N_43213,N_40801,N_40620);
or U43214 (N_43214,N_41382,N_41114);
xnor U43215 (N_43215,N_40551,N_40826);
or U43216 (N_43216,N_40219,N_40170);
and U43217 (N_43217,N_40255,N_41841);
xnor U43218 (N_43218,N_40494,N_41774);
nand U43219 (N_43219,N_41118,N_40669);
and U43220 (N_43220,N_41059,N_41944);
xor U43221 (N_43221,N_41642,N_40286);
or U43222 (N_43222,N_41122,N_41340);
and U43223 (N_43223,N_41971,N_41497);
nand U43224 (N_43224,N_40802,N_41851);
or U43225 (N_43225,N_40366,N_40893);
xnor U43226 (N_43226,N_41691,N_40074);
nand U43227 (N_43227,N_41294,N_40113);
and U43228 (N_43228,N_41794,N_40398);
and U43229 (N_43229,N_40363,N_41374);
nand U43230 (N_43230,N_40216,N_41203);
and U43231 (N_43231,N_41935,N_40691);
or U43232 (N_43232,N_40417,N_41855);
nand U43233 (N_43233,N_40645,N_41690);
xnor U43234 (N_43234,N_40031,N_41515);
xnor U43235 (N_43235,N_40481,N_41135);
and U43236 (N_43236,N_40929,N_41582);
nor U43237 (N_43237,N_40693,N_41687);
and U43238 (N_43238,N_40652,N_41030);
nand U43239 (N_43239,N_41333,N_40237);
xnor U43240 (N_43240,N_40119,N_41178);
xnor U43241 (N_43241,N_41154,N_40372);
nor U43242 (N_43242,N_40605,N_40977);
nor U43243 (N_43243,N_40353,N_41189);
nor U43244 (N_43244,N_41214,N_41933);
nand U43245 (N_43245,N_41472,N_40311);
xor U43246 (N_43246,N_40445,N_41082);
nand U43247 (N_43247,N_41847,N_41261);
nor U43248 (N_43248,N_41875,N_40615);
and U43249 (N_43249,N_41832,N_41664);
xor U43250 (N_43250,N_40838,N_40499);
xor U43251 (N_43251,N_40007,N_41974);
xor U43252 (N_43252,N_41373,N_41620);
xnor U43253 (N_43253,N_41485,N_40138);
xor U43254 (N_43254,N_41739,N_40960);
nor U43255 (N_43255,N_40385,N_40437);
or U43256 (N_43256,N_41856,N_41674);
and U43257 (N_43257,N_41732,N_41730);
xor U43258 (N_43258,N_41107,N_40689);
xor U43259 (N_43259,N_41891,N_41473);
xor U43260 (N_43260,N_41904,N_41210);
xor U43261 (N_43261,N_41164,N_40160);
and U43262 (N_43262,N_40012,N_41853);
xnor U43263 (N_43263,N_40523,N_40317);
nand U43264 (N_43264,N_41821,N_41596);
or U43265 (N_43265,N_41299,N_40187);
nor U43266 (N_43266,N_40265,N_40942);
nor U43267 (N_43267,N_40187,N_41940);
and U43268 (N_43268,N_41750,N_41416);
or U43269 (N_43269,N_40296,N_40952);
xor U43270 (N_43270,N_41941,N_40096);
nor U43271 (N_43271,N_40841,N_41734);
nand U43272 (N_43272,N_41698,N_40602);
or U43273 (N_43273,N_41672,N_41811);
and U43274 (N_43274,N_40190,N_41572);
or U43275 (N_43275,N_40522,N_40093);
or U43276 (N_43276,N_40788,N_40655);
and U43277 (N_43277,N_40887,N_41122);
xnor U43278 (N_43278,N_41398,N_41438);
nor U43279 (N_43279,N_41786,N_40613);
and U43280 (N_43280,N_40507,N_41276);
nand U43281 (N_43281,N_41043,N_40644);
nor U43282 (N_43282,N_40043,N_40166);
nor U43283 (N_43283,N_41410,N_41119);
xor U43284 (N_43284,N_41421,N_41956);
or U43285 (N_43285,N_40503,N_40741);
xor U43286 (N_43286,N_41782,N_40021);
xnor U43287 (N_43287,N_41899,N_40136);
or U43288 (N_43288,N_41229,N_40062);
and U43289 (N_43289,N_41060,N_40314);
nand U43290 (N_43290,N_40431,N_40542);
xnor U43291 (N_43291,N_40976,N_41838);
nor U43292 (N_43292,N_41505,N_40839);
nor U43293 (N_43293,N_41016,N_40883);
nor U43294 (N_43294,N_41346,N_40347);
nand U43295 (N_43295,N_41422,N_41194);
nor U43296 (N_43296,N_40147,N_41016);
and U43297 (N_43297,N_40726,N_40938);
nor U43298 (N_43298,N_41260,N_41138);
and U43299 (N_43299,N_40220,N_40298);
nor U43300 (N_43300,N_41268,N_40728);
nor U43301 (N_43301,N_41712,N_41490);
nor U43302 (N_43302,N_40800,N_40416);
nand U43303 (N_43303,N_40488,N_40910);
nand U43304 (N_43304,N_41232,N_41923);
nor U43305 (N_43305,N_41693,N_41919);
or U43306 (N_43306,N_41646,N_41201);
or U43307 (N_43307,N_40240,N_41470);
xnor U43308 (N_43308,N_41214,N_40799);
nand U43309 (N_43309,N_41306,N_41189);
nand U43310 (N_43310,N_41322,N_41239);
nand U43311 (N_43311,N_41776,N_41636);
nand U43312 (N_43312,N_41309,N_41882);
and U43313 (N_43313,N_40034,N_40820);
and U43314 (N_43314,N_41682,N_41521);
xnor U43315 (N_43315,N_40099,N_40426);
nor U43316 (N_43316,N_40545,N_40533);
xnor U43317 (N_43317,N_41746,N_40802);
and U43318 (N_43318,N_41256,N_40257);
nand U43319 (N_43319,N_41816,N_40367);
or U43320 (N_43320,N_41695,N_41878);
xnor U43321 (N_43321,N_40173,N_41582);
nand U43322 (N_43322,N_40434,N_40766);
or U43323 (N_43323,N_41454,N_40823);
nand U43324 (N_43324,N_40300,N_40974);
xnor U43325 (N_43325,N_41218,N_41846);
and U43326 (N_43326,N_41563,N_41622);
nand U43327 (N_43327,N_41424,N_41907);
xnor U43328 (N_43328,N_41074,N_41799);
nand U43329 (N_43329,N_40588,N_41561);
nor U43330 (N_43330,N_40417,N_40237);
and U43331 (N_43331,N_41298,N_40206);
nand U43332 (N_43332,N_40599,N_40393);
nand U43333 (N_43333,N_40195,N_41844);
nor U43334 (N_43334,N_40293,N_41150);
and U43335 (N_43335,N_41021,N_40087);
nand U43336 (N_43336,N_40520,N_40712);
nor U43337 (N_43337,N_41194,N_41474);
xnor U43338 (N_43338,N_40775,N_40056);
and U43339 (N_43339,N_41361,N_41775);
nand U43340 (N_43340,N_40920,N_41201);
nand U43341 (N_43341,N_40583,N_40295);
xor U43342 (N_43342,N_41599,N_40910);
and U43343 (N_43343,N_40142,N_41135);
and U43344 (N_43344,N_40815,N_40095);
nor U43345 (N_43345,N_40521,N_41678);
nor U43346 (N_43346,N_41364,N_41591);
xnor U43347 (N_43347,N_40251,N_40044);
xor U43348 (N_43348,N_40999,N_40735);
or U43349 (N_43349,N_40268,N_40759);
xnor U43350 (N_43350,N_41393,N_41302);
or U43351 (N_43351,N_41701,N_41626);
nand U43352 (N_43352,N_40000,N_41707);
nand U43353 (N_43353,N_41029,N_41269);
or U43354 (N_43354,N_40843,N_40890);
xor U43355 (N_43355,N_41650,N_40613);
xnor U43356 (N_43356,N_41079,N_41914);
nor U43357 (N_43357,N_41098,N_41234);
xor U43358 (N_43358,N_41607,N_40142);
nor U43359 (N_43359,N_41318,N_40534);
or U43360 (N_43360,N_41350,N_40408);
xnor U43361 (N_43361,N_41090,N_40509);
nand U43362 (N_43362,N_41824,N_41927);
nand U43363 (N_43363,N_41496,N_40488);
nor U43364 (N_43364,N_40521,N_40504);
xor U43365 (N_43365,N_41070,N_41652);
nor U43366 (N_43366,N_41011,N_40987);
and U43367 (N_43367,N_41729,N_40176);
nand U43368 (N_43368,N_40890,N_40540);
nor U43369 (N_43369,N_40282,N_41618);
and U43370 (N_43370,N_41414,N_41194);
xnor U43371 (N_43371,N_41875,N_40606);
or U43372 (N_43372,N_41552,N_40831);
nand U43373 (N_43373,N_41171,N_40387);
nand U43374 (N_43374,N_41080,N_40424);
nand U43375 (N_43375,N_40154,N_41629);
xnor U43376 (N_43376,N_40559,N_40478);
nor U43377 (N_43377,N_40822,N_41154);
xor U43378 (N_43378,N_41961,N_40635);
xnor U43379 (N_43379,N_41198,N_40435);
xor U43380 (N_43380,N_41561,N_40564);
nor U43381 (N_43381,N_40301,N_41160);
xnor U43382 (N_43382,N_41600,N_41274);
xor U43383 (N_43383,N_40028,N_41268);
nand U43384 (N_43384,N_41206,N_41328);
or U43385 (N_43385,N_41478,N_40810);
nor U43386 (N_43386,N_40787,N_40838);
and U43387 (N_43387,N_41777,N_41222);
and U43388 (N_43388,N_40348,N_41082);
or U43389 (N_43389,N_41506,N_40320);
xnor U43390 (N_43390,N_41374,N_40391);
nand U43391 (N_43391,N_40127,N_41194);
xor U43392 (N_43392,N_40836,N_40874);
nand U43393 (N_43393,N_41539,N_40617);
nor U43394 (N_43394,N_40607,N_41433);
nor U43395 (N_43395,N_41199,N_40761);
xnor U43396 (N_43396,N_41425,N_41686);
or U43397 (N_43397,N_41036,N_40653);
xnor U43398 (N_43398,N_40941,N_40051);
nor U43399 (N_43399,N_41645,N_40192);
and U43400 (N_43400,N_41955,N_41284);
xnor U43401 (N_43401,N_41497,N_40219);
nor U43402 (N_43402,N_41501,N_40532);
xnor U43403 (N_43403,N_40144,N_41384);
and U43404 (N_43404,N_41313,N_40721);
and U43405 (N_43405,N_40014,N_40698);
nor U43406 (N_43406,N_40117,N_41355);
xor U43407 (N_43407,N_40605,N_41552);
nand U43408 (N_43408,N_40935,N_40983);
and U43409 (N_43409,N_40240,N_41900);
nor U43410 (N_43410,N_41361,N_40577);
nor U43411 (N_43411,N_40956,N_41512);
xnor U43412 (N_43412,N_41815,N_41885);
or U43413 (N_43413,N_40316,N_41061);
or U43414 (N_43414,N_41933,N_40035);
xnor U43415 (N_43415,N_41662,N_40953);
nor U43416 (N_43416,N_41611,N_41116);
and U43417 (N_43417,N_40112,N_40428);
and U43418 (N_43418,N_40114,N_41005);
xnor U43419 (N_43419,N_40633,N_41745);
nor U43420 (N_43420,N_41926,N_41533);
nand U43421 (N_43421,N_41838,N_40173);
or U43422 (N_43422,N_40312,N_40009);
nand U43423 (N_43423,N_41510,N_40863);
xor U43424 (N_43424,N_41548,N_40969);
or U43425 (N_43425,N_40905,N_40528);
xor U43426 (N_43426,N_41694,N_41258);
or U43427 (N_43427,N_41620,N_41786);
nand U43428 (N_43428,N_41608,N_41358);
xnor U43429 (N_43429,N_40470,N_40397);
nor U43430 (N_43430,N_40848,N_41177);
or U43431 (N_43431,N_40773,N_40212);
and U43432 (N_43432,N_41596,N_41692);
nand U43433 (N_43433,N_41799,N_40432);
nand U43434 (N_43434,N_40507,N_41088);
xnor U43435 (N_43435,N_41273,N_41803);
xor U43436 (N_43436,N_40623,N_41125);
xor U43437 (N_43437,N_40786,N_40367);
nand U43438 (N_43438,N_41422,N_41734);
nand U43439 (N_43439,N_40649,N_40158);
nor U43440 (N_43440,N_41972,N_41756);
and U43441 (N_43441,N_40120,N_40153);
xnor U43442 (N_43442,N_41269,N_40060);
and U43443 (N_43443,N_40799,N_41481);
or U43444 (N_43444,N_40055,N_40561);
nand U43445 (N_43445,N_40324,N_41593);
nand U43446 (N_43446,N_40477,N_41702);
nor U43447 (N_43447,N_41338,N_41462);
nand U43448 (N_43448,N_41160,N_40394);
nor U43449 (N_43449,N_41696,N_41927);
or U43450 (N_43450,N_40236,N_41387);
nor U43451 (N_43451,N_40404,N_40355);
xor U43452 (N_43452,N_40587,N_41364);
and U43453 (N_43453,N_41786,N_40664);
xor U43454 (N_43454,N_40930,N_40811);
xor U43455 (N_43455,N_41655,N_40144);
or U43456 (N_43456,N_40021,N_40681);
or U43457 (N_43457,N_40494,N_40299);
nand U43458 (N_43458,N_40303,N_41275);
and U43459 (N_43459,N_41373,N_41155);
and U43460 (N_43460,N_40278,N_40178);
or U43461 (N_43461,N_40693,N_41841);
or U43462 (N_43462,N_41395,N_41784);
xnor U43463 (N_43463,N_41244,N_40640);
or U43464 (N_43464,N_40699,N_41622);
nand U43465 (N_43465,N_40283,N_40872);
or U43466 (N_43466,N_40425,N_40915);
xnor U43467 (N_43467,N_40533,N_40155);
nand U43468 (N_43468,N_41474,N_40762);
nand U43469 (N_43469,N_40496,N_40190);
and U43470 (N_43470,N_40986,N_41711);
nor U43471 (N_43471,N_41506,N_41041);
and U43472 (N_43472,N_41983,N_41154);
xor U43473 (N_43473,N_41765,N_40047);
or U43474 (N_43474,N_40482,N_40611);
or U43475 (N_43475,N_40566,N_40570);
or U43476 (N_43476,N_41401,N_40198);
xnor U43477 (N_43477,N_40206,N_41795);
nor U43478 (N_43478,N_40023,N_41448);
xnor U43479 (N_43479,N_41039,N_40147);
xnor U43480 (N_43480,N_41868,N_41750);
xnor U43481 (N_43481,N_41587,N_40665);
nand U43482 (N_43482,N_41466,N_40828);
or U43483 (N_43483,N_40444,N_41847);
nand U43484 (N_43484,N_40788,N_41515);
nor U43485 (N_43485,N_40697,N_40604);
nand U43486 (N_43486,N_40887,N_41732);
xor U43487 (N_43487,N_41291,N_41533);
and U43488 (N_43488,N_40607,N_41776);
nand U43489 (N_43489,N_41304,N_41425);
xor U43490 (N_43490,N_41536,N_40344);
xor U43491 (N_43491,N_41488,N_40083);
nand U43492 (N_43492,N_41009,N_41519);
xor U43493 (N_43493,N_41415,N_41788);
and U43494 (N_43494,N_40765,N_40436);
and U43495 (N_43495,N_41841,N_40143);
and U43496 (N_43496,N_40688,N_41826);
and U43497 (N_43497,N_40868,N_41572);
xor U43498 (N_43498,N_40831,N_40172);
nand U43499 (N_43499,N_40275,N_40752);
nand U43500 (N_43500,N_41772,N_41473);
or U43501 (N_43501,N_41759,N_40506);
and U43502 (N_43502,N_41134,N_40944);
or U43503 (N_43503,N_41792,N_41106);
or U43504 (N_43504,N_41368,N_40886);
xnor U43505 (N_43505,N_41900,N_41095);
or U43506 (N_43506,N_41908,N_41596);
or U43507 (N_43507,N_40075,N_41096);
and U43508 (N_43508,N_40912,N_40462);
and U43509 (N_43509,N_41016,N_40148);
and U43510 (N_43510,N_41410,N_40467);
nor U43511 (N_43511,N_41936,N_40720);
nand U43512 (N_43512,N_40681,N_40756);
nand U43513 (N_43513,N_41976,N_41273);
and U43514 (N_43514,N_40498,N_40631);
and U43515 (N_43515,N_41238,N_40293);
and U43516 (N_43516,N_40675,N_40568);
xor U43517 (N_43517,N_41775,N_40608);
or U43518 (N_43518,N_41157,N_40799);
xor U43519 (N_43519,N_40804,N_41985);
xnor U43520 (N_43520,N_41925,N_41092);
nor U43521 (N_43521,N_40565,N_41651);
or U43522 (N_43522,N_40771,N_41724);
or U43523 (N_43523,N_41283,N_41687);
and U43524 (N_43524,N_40561,N_40360);
or U43525 (N_43525,N_40490,N_40850);
or U43526 (N_43526,N_40097,N_40183);
nor U43527 (N_43527,N_40897,N_40356);
or U43528 (N_43528,N_40046,N_40674);
and U43529 (N_43529,N_40886,N_40530);
xor U43530 (N_43530,N_41066,N_41449);
nor U43531 (N_43531,N_40455,N_40003);
or U43532 (N_43532,N_40492,N_40292);
nand U43533 (N_43533,N_41825,N_40104);
nor U43534 (N_43534,N_40264,N_41806);
nor U43535 (N_43535,N_41046,N_40673);
or U43536 (N_43536,N_41944,N_40515);
xnor U43537 (N_43537,N_40868,N_40920);
nor U43538 (N_43538,N_41468,N_41727);
xor U43539 (N_43539,N_41960,N_41880);
nor U43540 (N_43540,N_40680,N_40110);
nor U43541 (N_43541,N_41761,N_41413);
xor U43542 (N_43542,N_40339,N_41308);
xor U43543 (N_43543,N_40040,N_40451);
nor U43544 (N_43544,N_40965,N_41639);
or U43545 (N_43545,N_41542,N_41273);
xnor U43546 (N_43546,N_40396,N_40518);
nor U43547 (N_43547,N_40550,N_40363);
xnor U43548 (N_43548,N_40377,N_41673);
nand U43549 (N_43549,N_40053,N_40919);
or U43550 (N_43550,N_41984,N_41886);
nand U43551 (N_43551,N_40617,N_40683);
nor U43552 (N_43552,N_40588,N_40920);
nand U43553 (N_43553,N_40085,N_40318);
xor U43554 (N_43554,N_41596,N_41516);
nor U43555 (N_43555,N_40056,N_41960);
and U43556 (N_43556,N_40121,N_41251);
nor U43557 (N_43557,N_41514,N_41431);
and U43558 (N_43558,N_40797,N_41938);
and U43559 (N_43559,N_40645,N_40218);
nand U43560 (N_43560,N_40489,N_40786);
nor U43561 (N_43561,N_41502,N_41962);
nor U43562 (N_43562,N_41315,N_40554);
nand U43563 (N_43563,N_40256,N_41896);
nand U43564 (N_43564,N_41303,N_40168);
or U43565 (N_43565,N_40289,N_41330);
nor U43566 (N_43566,N_41142,N_40284);
nand U43567 (N_43567,N_40555,N_40629);
and U43568 (N_43568,N_40804,N_40545);
nor U43569 (N_43569,N_40678,N_40282);
xnor U43570 (N_43570,N_41272,N_41325);
and U43571 (N_43571,N_40649,N_41126);
xnor U43572 (N_43572,N_41204,N_40363);
nand U43573 (N_43573,N_41311,N_40533);
xor U43574 (N_43574,N_40598,N_41706);
nor U43575 (N_43575,N_40377,N_40661);
nor U43576 (N_43576,N_40276,N_41777);
nor U43577 (N_43577,N_41355,N_40526);
nand U43578 (N_43578,N_41214,N_40855);
and U43579 (N_43579,N_40246,N_40973);
nor U43580 (N_43580,N_41334,N_41365);
nor U43581 (N_43581,N_40287,N_40630);
xnor U43582 (N_43582,N_41448,N_40730);
and U43583 (N_43583,N_40708,N_40852);
nand U43584 (N_43584,N_41991,N_41216);
nand U43585 (N_43585,N_40765,N_40622);
and U43586 (N_43586,N_41703,N_41100);
nand U43587 (N_43587,N_41749,N_41761);
xor U43588 (N_43588,N_41989,N_41413);
nor U43589 (N_43589,N_41155,N_41061);
xnor U43590 (N_43590,N_41215,N_41565);
nor U43591 (N_43591,N_40197,N_40466);
and U43592 (N_43592,N_40500,N_41188);
nand U43593 (N_43593,N_40834,N_40182);
and U43594 (N_43594,N_40098,N_40495);
or U43595 (N_43595,N_40237,N_41719);
nor U43596 (N_43596,N_40512,N_41479);
xor U43597 (N_43597,N_40164,N_40586);
nand U43598 (N_43598,N_41360,N_41991);
nand U43599 (N_43599,N_40093,N_40207);
or U43600 (N_43600,N_41185,N_40227);
or U43601 (N_43601,N_41894,N_40855);
nand U43602 (N_43602,N_40543,N_41036);
nor U43603 (N_43603,N_41026,N_41264);
nand U43604 (N_43604,N_40657,N_41149);
xnor U43605 (N_43605,N_40481,N_40422);
nor U43606 (N_43606,N_40147,N_41903);
xnor U43607 (N_43607,N_40256,N_40638);
nand U43608 (N_43608,N_40669,N_41771);
nand U43609 (N_43609,N_40130,N_41679);
or U43610 (N_43610,N_40710,N_40375);
and U43611 (N_43611,N_41029,N_41368);
or U43612 (N_43612,N_40628,N_40116);
or U43613 (N_43613,N_41270,N_40662);
nor U43614 (N_43614,N_41894,N_41239);
nor U43615 (N_43615,N_40372,N_41300);
nand U43616 (N_43616,N_40948,N_40490);
and U43617 (N_43617,N_41908,N_40835);
xor U43618 (N_43618,N_40385,N_41182);
nor U43619 (N_43619,N_41554,N_40438);
nand U43620 (N_43620,N_41900,N_40323);
or U43621 (N_43621,N_41643,N_40847);
xor U43622 (N_43622,N_41494,N_40174);
or U43623 (N_43623,N_41966,N_41386);
or U43624 (N_43624,N_40422,N_40971);
nor U43625 (N_43625,N_41920,N_41779);
and U43626 (N_43626,N_41927,N_40742);
or U43627 (N_43627,N_41889,N_40394);
and U43628 (N_43628,N_41598,N_40712);
nand U43629 (N_43629,N_41420,N_40599);
and U43630 (N_43630,N_40345,N_41306);
or U43631 (N_43631,N_41457,N_40010);
and U43632 (N_43632,N_40535,N_40401);
nor U43633 (N_43633,N_40202,N_40174);
xnor U43634 (N_43634,N_40644,N_41449);
xnor U43635 (N_43635,N_40200,N_40882);
and U43636 (N_43636,N_41117,N_40602);
nand U43637 (N_43637,N_40828,N_40146);
nand U43638 (N_43638,N_40975,N_41747);
or U43639 (N_43639,N_40322,N_41553);
nor U43640 (N_43640,N_40486,N_41197);
xnor U43641 (N_43641,N_41532,N_41419);
nor U43642 (N_43642,N_41481,N_40152);
nand U43643 (N_43643,N_41830,N_41384);
nor U43644 (N_43644,N_41259,N_40027);
or U43645 (N_43645,N_40732,N_40844);
nand U43646 (N_43646,N_40055,N_41059);
and U43647 (N_43647,N_41956,N_41716);
xnor U43648 (N_43648,N_40053,N_41126);
xnor U43649 (N_43649,N_41937,N_40756);
nand U43650 (N_43650,N_41582,N_41109);
xor U43651 (N_43651,N_41201,N_41656);
or U43652 (N_43652,N_40707,N_40847);
nor U43653 (N_43653,N_41587,N_40157);
or U43654 (N_43654,N_41244,N_40190);
or U43655 (N_43655,N_40777,N_41090);
and U43656 (N_43656,N_40677,N_40384);
or U43657 (N_43657,N_41838,N_41626);
nand U43658 (N_43658,N_40174,N_40241);
nor U43659 (N_43659,N_40258,N_41125);
xor U43660 (N_43660,N_41229,N_40698);
or U43661 (N_43661,N_40044,N_40321);
or U43662 (N_43662,N_40221,N_40336);
or U43663 (N_43663,N_40863,N_41723);
or U43664 (N_43664,N_41254,N_40388);
or U43665 (N_43665,N_41161,N_41368);
nand U43666 (N_43666,N_40256,N_41750);
xor U43667 (N_43667,N_41512,N_41528);
or U43668 (N_43668,N_40944,N_41271);
xnor U43669 (N_43669,N_41448,N_40293);
or U43670 (N_43670,N_41788,N_40860);
nand U43671 (N_43671,N_40035,N_41636);
and U43672 (N_43672,N_40928,N_40899);
nor U43673 (N_43673,N_40202,N_41053);
or U43674 (N_43674,N_40457,N_40423);
and U43675 (N_43675,N_40839,N_41347);
or U43676 (N_43676,N_41844,N_41221);
or U43677 (N_43677,N_40372,N_41041);
xor U43678 (N_43678,N_41986,N_41835);
xnor U43679 (N_43679,N_41626,N_41850);
xor U43680 (N_43680,N_41846,N_41489);
or U43681 (N_43681,N_40525,N_40087);
xnor U43682 (N_43682,N_40667,N_41482);
nand U43683 (N_43683,N_40336,N_41829);
xor U43684 (N_43684,N_41357,N_40480);
nor U43685 (N_43685,N_41431,N_41860);
nand U43686 (N_43686,N_41766,N_40104);
nand U43687 (N_43687,N_41677,N_41200);
and U43688 (N_43688,N_41677,N_41777);
nand U43689 (N_43689,N_40173,N_41302);
or U43690 (N_43690,N_41821,N_41894);
nor U43691 (N_43691,N_40755,N_41970);
nor U43692 (N_43692,N_40038,N_41642);
xor U43693 (N_43693,N_41603,N_41860);
nand U43694 (N_43694,N_40960,N_40844);
and U43695 (N_43695,N_41891,N_41857);
or U43696 (N_43696,N_40242,N_40783);
nand U43697 (N_43697,N_41136,N_40222);
nand U43698 (N_43698,N_40193,N_40557);
or U43699 (N_43699,N_41262,N_41177);
and U43700 (N_43700,N_41518,N_41954);
nor U43701 (N_43701,N_40281,N_40487);
and U43702 (N_43702,N_41114,N_41726);
or U43703 (N_43703,N_41500,N_40043);
or U43704 (N_43704,N_40870,N_41540);
nor U43705 (N_43705,N_41036,N_41928);
or U43706 (N_43706,N_41256,N_40361);
or U43707 (N_43707,N_40265,N_41008);
xnor U43708 (N_43708,N_40172,N_41765);
and U43709 (N_43709,N_40476,N_41112);
and U43710 (N_43710,N_41856,N_41608);
and U43711 (N_43711,N_41903,N_41857);
xnor U43712 (N_43712,N_40016,N_40878);
nand U43713 (N_43713,N_41955,N_41279);
or U43714 (N_43714,N_40957,N_40669);
xnor U43715 (N_43715,N_41795,N_41750);
nor U43716 (N_43716,N_40512,N_40358);
nand U43717 (N_43717,N_40368,N_41556);
nor U43718 (N_43718,N_40042,N_40591);
or U43719 (N_43719,N_41861,N_40057);
nor U43720 (N_43720,N_40538,N_40301);
nor U43721 (N_43721,N_41587,N_41053);
and U43722 (N_43722,N_40365,N_40800);
xor U43723 (N_43723,N_41489,N_40557);
and U43724 (N_43724,N_40141,N_40619);
or U43725 (N_43725,N_40420,N_40596);
or U43726 (N_43726,N_40763,N_41139);
xor U43727 (N_43727,N_40990,N_40404);
or U43728 (N_43728,N_40796,N_40476);
nand U43729 (N_43729,N_41796,N_41412);
xor U43730 (N_43730,N_41381,N_40231);
or U43731 (N_43731,N_41123,N_40953);
nor U43732 (N_43732,N_40643,N_41321);
and U43733 (N_43733,N_40714,N_41924);
nand U43734 (N_43734,N_40031,N_41990);
nand U43735 (N_43735,N_40361,N_40488);
xor U43736 (N_43736,N_40603,N_40495);
and U43737 (N_43737,N_40713,N_41350);
or U43738 (N_43738,N_41309,N_41062);
nand U43739 (N_43739,N_41776,N_40988);
nor U43740 (N_43740,N_40713,N_40682);
and U43741 (N_43741,N_41224,N_40964);
nor U43742 (N_43742,N_40163,N_41556);
xnor U43743 (N_43743,N_40763,N_41484);
or U43744 (N_43744,N_41380,N_40820);
or U43745 (N_43745,N_41313,N_41432);
and U43746 (N_43746,N_40940,N_40451);
and U43747 (N_43747,N_40409,N_41347);
nand U43748 (N_43748,N_40494,N_41470);
nand U43749 (N_43749,N_41340,N_41597);
xor U43750 (N_43750,N_40231,N_40843);
nand U43751 (N_43751,N_40954,N_40894);
xor U43752 (N_43752,N_40251,N_41367);
nor U43753 (N_43753,N_41349,N_40930);
or U43754 (N_43754,N_41979,N_40280);
or U43755 (N_43755,N_41065,N_40324);
nor U43756 (N_43756,N_40231,N_41743);
xnor U43757 (N_43757,N_40593,N_40689);
or U43758 (N_43758,N_41639,N_40961);
xnor U43759 (N_43759,N_40579,N_40424);
or U43760 (N_43760,N_40513,N_41226);
nand U43761 (N_43761,N_40939,N_40881);
nand U43762 (N_43762,N_41458,N_41056);
xnor U43763 (N_43763,N_41472,N_41438);
xnor U43764 (N_43764,N_40118,N_41450);
xor U43765 (N_43765,N_40612,N_40476);
xor U43766 (N_43766,N_41301,N_40202);
and U43767 (N_43767,N_40858,N_40681);
and U43768 (N_43768,N_41092,N_40780);
xnor U43769 (N_43769,N_40311,N_40575);
xor U43770 (N_43770,N_41677,N_40040);
or U43771 (N_43771,N_40653,N_41366);
and U43772 (N_43772,N_41365,N_40538);
and U43773 (N_43773,N_41780,N_41591);
and U43774 (N_43774,N_41965,N_40731);
xor U43775 (N_43775,N_41119,N_41273);
nor U43776 (N_43776,N_40721,N_40580);
nand U43777 (N_43777,N_41024,N_41774);
or U43778 (N_43778,N_41907,N_41596);
or U43779 (N_43779,N_41770,N_40985);
xor U43780 (N_43780,N_41250,N_41799);
nor U43781 (N_43781,N_41439,N_41686);
or U43782 (N_43782,N_40276,N_40542);
or U43783 (N_43783,N_41902,N_41653);
and U43784 (N_43784,N_40674,N_40578);
xnor U43785 (N_43785,N_41558,N_40830);
and U43786 (N_43786,N_41585,N_41801);
or U43787 (N_43787,N_40759,N_41086);
nand U43788 (N_43788,N_41953,N_40047);
xor U43789 (N_43789,N_40444,N_40183);
and U43790 (N_43790,N_40294,N_40747);
and U43791 (N_43791,N_41929,N_40099);
xor U43792 (N_43792,N_41139,N_40994);
nand U43793 (N_43793,N_40580,N_40343);
nand U43794 (N_43794,N_41436,N_40781);
nor U43795 (N_43795,N_41518,N_41177);
or U43796 (N_43796,N_41405,N_40508);
or U43797 (N_43797,N_41084,N_41895);
or U43798 (N_43798,N_41393,N_40960);
and U43799 (N_43799,N_41331,N_41286);
nor U43800 (N_43800,N_41126,N_40962);
nand U43801 (N_43801,N_41866,N_40811);
xnor U43802 (N_43802,N_40679,N_41413);
and U43803 (N_43803,N_40044,N_40418);
nand U43804 (N_43804,N_40037,N_41121);
or U43805 (N_43805,N_41738,N_41600);
nor U43806 (N_43806,N_41416,N_40245);
xnor U43807 (N_43807,N_40929,N_40825);
or U43808 (N_43808,N_40062,N_40393);
nor U43809 (N_43809,N_40240,N_40979);
nor U43810 (N_43810,N_40391,N_41639);
or U43811 (N_43811,N_40133,N_41431);
and U43812 (N_43812,N_41187,N_40011);
and U43813 (N_43813,N_40106,N_41790);
and U43814 (N_43814,N_41032,N_40198);
xnor U43815 (N_43815,N_41965,N_40412);
nor U43816 (N_43816,N_40340,N_41176);
nand U43817 (N_43817,N_41918,N_40660);
nand U43818 (N_43818,N_41823,N_41123);
xnor U43819 (N_43819,N_41171,N_40342);
or U43820 (N_43820,N_40652,N_40625);
nor U43821 (N_43821,N_41912,N_41941);
nand U43822 (N_43822,N_40648,N_41613);
nor U43823 (N_43823,N_41755,N_41417);
and U43824 (N_43824,N_40407,N_41320);
xnor U43825 (N_43825,N_41655,N_40114);
xor U43826 (N_43826,N_40793,N_40051);
or U43827 (N_43827,N_41372,N_41011);
and U43828 (N_43828,N_41508,N_41407);
and U43829 (N_43829,N_40136,N_40176);
nand U43830 (N_43830,N_41404,N_40826);
or U43831 (N_43831,N_40923,N_41026);
nor U43832 (N_43832,N_41826,N_41693);
nor U43833 (N_43833,N_40170,N_41502);
and U43834 (N_43834,N_40530,N_40368);
and U43835 (N_43835,N_40939,N_41418);
nand U43836 (N_43836,N_41619,N_40186);
or U43837 (N_43837,N_40223,N_41991);
nor U43838 (N_43838,N_41237,N_40898);
nor U43839 (N_43839,N_41491,N_41741);
and U43840 (N_43840,N_41911,N_40839);
and U43841 (N_43841,N_40411,N_40431);
xnor U43842 (N_43842,N_41474,N_40341);
nand U43843 (N_43843,N_41496,N_40377);
nor U43844 (N_43844,N_41486,N_40465);
nand U43845 (N_43845,N_41478,N_40430);
or U43846 (N_43846,N_40490,N_40886);
or U43847 (N_43847,N_40873,N_41787);
or U43848 (N_43848,N_40734,N_40045);
or U43849 (N_43849,N_40525,N_41264);
nor U43850 (N_43850,N_40959,N_41877);
nor U43851 (N_43851,N_40281,N_40812);
nand U43852 (N_43852,N_40879,N_41876);
and U43853 (N_43853,N_41306,N_40107);
nor U43854 (N_43854,N_41837,N_40590);
xor U43855 (N_43855,N_40631,N_41549);
xor U43856 (N_43856,N_41287,N_40718);
nand U43857 (N_43857,N_40133,N_41475);
and U43858 (N_43858,N_41510,N_40733);
nand U43859 (N_43859,N_41248,N_41240);
xor U43860 (N_43860,N_40358,N_41078);
xnor U43861 (N_43861,N_41133,N_41035);
and U43862 (N_43862,N_40653,N_41488);
and U43863 (N_43863,N_41949,N_41195);
xnor U43864 (N_43864,N_41638,N_41823);
nor U43865 (N_43865,N_40819,N_40507);
xnor U43866 (N_43866,N_40478,N_41619);
xnor U43867 (N_43867,N_41122,N_41319);
nor U43868 (N_43868,N_40288,N_40109);
or U43869 (N_43869,N_40838,N_41860);
and U43870 (N_43870,N_41516,N_40779);
nand U43871 (N_43871,N_41814,N_40931);
nor U43872 (N_43872,N_40140,N_40765);
and U43873 (N_43873,N_41812,N_40806);
nand U43874 (N_43874,N_41461,N_41264);
nand U43875 (N_43875,N_40816,N_40906);
xnor U43876 (N_43876,N_41777,N_40396);
nand U43877 (N_43877,N_40712,N_40907);
or U43878 (N_43878,N_40702,N_41191);
or U43879 (N_43879,N_40477,N_41564);
and U43880 (N_43880,N_40722,N_40099);
and U43881 (N_43881,N_40834,N_40214);
xnor U43882 (N_43882,N_40069,N_41219);
nand U43883 (N_43883,N_40928,N_40587);
nand U43884 (N_43884,N_41383,N_41955);
xor U43885 (N_43885,N_41888,N_41821);
or U43886 (N_43886,N_41701,N_40686);
and U43887 (N_43887,N_41719,N_40114);
nand U43888 (N_43888,N_41609,N_41051);
nand U43889 (N_43889,N_41255,N_41944);
xnor U43890 (N_43890,N_41280,N_40361);
or U43891 (N_43891,N_40743,N_40571);
and U43892 (N_43892,N_41632,N_40402);
xor U43893 (N_43893,N_41746,N_40257);
or U43894 (N_43894,N_40010,N_40745);
nand U43895 (N_43895,N_40900,N_41870);
or U43896 (N_43896,N_41264,N_41705);
nand U43897 (N_43897,N_41233,N_41333);
nand U43898 (N_43898,N_41134,N_40954);
and U43899 (N_43899,N_41822,N_41954);
nand U43900 (N_43900,N_41122,N_40554);
or U43901 (N_43901,N_40706,N_41919);
nand U43902 (N_43902,N_40549,N_41861);
and U43903 (N_43903,N_40341,N_40617);
xor U43904 (N_43904,N_40760,N_40494);
nor U43905 (N_43905,N_40916,N_41989);
or U43906 (N_43906,N_40671,N_40838);
nand U43907 (N_43907,N_41489,N_41046);
nor U43908 (N_43908,N_40526,N_41653);
nand U43909 (N_43909,N_40587,N_41949);
or U43910 (N_43910,N_41272,N_40268);
or U43911 (N_43911,N_41075,N_41550);
nor U43912 (N_43912,N_41111,N_40195);
nand U43913 (N_43913,N_40034,N_41747);
nand U43914 (N_43914,N_41083,N_40972);
xor U43915 (N_43915,N_40510,N_40967);
or U43916 (N_43916,N_41045,N_41998);
nor U43917 (N_43917,N_40951,N_41257);
and U43918 (N_43918,N_40883,N_40107);
or U43919 (N_43919,N_41724,N_41889);
or U43920 (N_43920,N_41238,N_40796);
or U43921 (N_43921,N_41234,N_40164);
and U43922 (N_43922,N_41258,N_40059);
xor U43923 (N_43923,N_41698,N_41991);
nand U43924 (N_43924,N_41930,N_41750);
nor U43925 (N_43925,N_41984,N_40327);
xnor U43926 (N_43926,N_41626,N_41000);
and U43927 (N_43927,N_40589,N_41233);
and U43928 (N_43928,N_40776,N_41684);
nand U43929 (N_43929,N_40730,N_41203);
and U43930 (N_43930,N_41535,N_40158);
nor U43931 (N_43931,N_40970,N_41921);
nand U43932 (N_43932,N_40541,N_41925);
and U43933 (N_43933,N_41015,N_40350);
or U43934 (N_43934,N_40521,N_40877);
or U43935 (N_43935,N_41011,N_40392);
and U43936 (N_43936,N_41418,N_40180);
and U43937 (N_43937,N_41377,N_41259);
nand U43938 (N_43938,N_40526,N_40769);
xnor U43939 (N_43939,N_40143,N_40234);
nor U43940 (N_43940,N_40769,N_40253);
xor U43941 (N_43941,N_41253,N_40511);
and U43942 (N_43942,N_41896,N_41422);
and U43943 (N_43943,N_40174,N_41776);
and U43944 (N_43944,N_40506,N_41889);
nor U43945 (N_43945,N_40545,N_40760);
xor U43946 (N_43946,N_40705,N_40725);
xnor U43947 (N_43947,N_41233,N_40167);
nor U43948 (N_43948,N_41025,N_40944);
nand U43949 (N_43949,N_41202,N_40722);
nor U43950 (N_43950,N_40679,N_40085);
nor U43951 (N_43951,N_41782,N_40475);
or U43952 (N_43952,N_40529,N_40050);
and U43953 (N_43953,N_41542,N_41000);
or U43954 (N_43954,N_40840,N_41544);
nor U43955 (N_43955,N_41797,N_41543);
nor U43956 (N_43956,N_40501,N_40312);
nand U43957 (N_43957,N_40506,N_40090);
or U43958 (N_43958,N_40872,N_40423);
and U43959 (N_43959,N_40670,N_41087);
xnor U43960 (N_43960,N_41809,N_41817);
or U43961 (N_43961,N_40572,N_41102);
or U43962 (N_43962,N_41306,N_40503);
nor U43963 (N_43963,N_40472,N_40429);
nand U43964 (N_43964,N_41478,N_40241);
nor U43965 (N_43965,N_40180,N_40812);
nand U43966 (N_43966,N_41396,N_40211);
or U43967 (N_43967,N_40498,N_40053);
nor U43968 (N_43968,N_40548,N_40941);
nand U43969 (N_43969,N_40477,N_41603);
xnor U43970 (N_43970,N_40217,N_40580);
nor U43971 (N_43971,N_40088,N_41658);
nor U43972 (N_43972,N_40494,N_41337);
nand U43973 (N_43973,N_40773,N_40995);
nand U43974 (N_43974,N_41883,N_40250);
nor U43975 (N_43975,N_40811,N_40698);
nor U43976 (N_43976,N_40146,N_40472);
and U43977 (N_43977,N_40836,N_40248);
xnor U43978 (N_43978,N_41970,N_41636);
xnor U43979 (N_43979,N_41464,N_41661);
xor U43980 (N_43980,N_40893,N_40543);
nand U43981 (N_43981,N_41206,N_41581);
and U43982 (N_43982,N_41479,N_41852);
and U43983 (N_43983,N_40763,N_40016);
or U43984 (N_43984,N_41103,N_40941);
xor U43985 (N_43985,N_40062,N_41323);
nand U43986 (N_43986,N_40960,N_41747);
xor U43987 (N_43987,N_40839,N_41709);
xnor U43988 (N_43988,N_41900,N_41227);
xnor U43989 (N_43989,N_40648,N_41307);
nor U43990 (N_43990,N_40069,N_41076);
nor U43991 (N_43991,N_41981,N_40602);
and U43992 (N_43992,N_40514,N_41321);
or U43993 (N_43993,N_40735,N_40482);
and U43994 (N_43994,N_40381,N_40146);
nor U43995 (N_43995,N_41826,N_40225);
and U43996 (N_43996,N_41346,N_40387);
xnor U43997 (N_43997,N_41583,N_40978);
xor U43998 (N_43998,N_41090,N_41022);
and U43999 (N_43999,N_40203,N_40602);
nand U44000 (N_44000,N_43695,N_43370);
nand U44001 (N_44001,N_42295,N_43259);
and U44002 (N_44002,N_43077,N_43288);
nand U44003 (N_44003,N_43844,N_43228);
nor U44004 (N_44004,N_42769,N_42373);
xnor U44005 (N_44005,N_43810,N_42882);
or U44006 (N_44006,N_43216,N_42068);
and U44007 (N_44007,N_43504,N_42365);
nor U44008 (N_44008,N_43709,N_42687);
xor U44009 (N_44009,N_42027,N_42437);
nor U44010 (N_44010,N_43722,N_42553);
or U44011 (N_44011,N_43892,N_43962);
nand U44012 (N_44012,N_42860,N_43053);
nand U44013 (N_44013,N_42163,N_43935);
xnor U44014 (N_44014,N_43424,N_42511);
nor U44015 (N_44015,N_42085,N_43969);
nand U44016 (N_44016,N_43867,N_42035);
xnor U44017 (N_44017,N_42794,N_42904);
and U44018 (N_44018,N_42870,N_42773);
nor U44019 (N_44019,N_43586,N_42734);
or U44020 (N_44020,N_42240,N_43774);
and U44021 (N_44021,N_42722,N_43912);
and U44022 (N_44022,N_42417,N_42227);
nor U44023 (N_44023,N_42940,N_43669);
nand U44024 (N_44024,N_43219,N_43283);
nand U44025 (N_44025,N_42237,N_43515);
and U44026 (N_44026,N_42479,N_43990);
nand U44027 (N_44027,N_42966,N_42728);
xnor U44028 (N_44028,N_43580,N_43750);
xor U44029 (N_44029,N_42592,N_43270);
nor U44030 (N_44030,N_42761,N_42402);
nor U44031 (N_44031,N_42810,N_42421);
nand U44032 (N_44032,N_43206,N_42918);
or U44033 (N_44033,N_42989,N_42106);
nand U44034 (N_44034,N_43401,N_42880);
nand U44035 (N_44035,N_43018,N_43576);
nor U44036 (N_44036,N_42132,N_42403);
nand U44037 (N_44037,N_43532,N_43347);
xnor U44038 (N_44038,N_42384,N_42610);
xnor U44039 (N_44039,N_42385,N_43595);
xnor U44040 (N_44040,N_42919,N_43970);
and U44041 (N_44041,N_42429,N_42122);
xnor U44042 (N_44042,N_43826,N_42829);
nor U44043 (N_44043,N_43394,N_42501);
xnor U44044 (N_44044,N_42816,N_42454);
nor U44045 (N_44045,N_43457,N_42790);
or U44046 (N_44046,N_43195,N_43254);
and U44047 (N_44047,N_42236,N_42216);
xor U44048 (N_44048,N_43146,N_43732);
nand U44049 (N_44049,N_42518,N_43545);
and U44050 (N_44050,N_43608,N_42928);
nor U44051 (N_44051,N_42674,N_43325);
and U44052 (N_44052,N_42475,N_43764);
nor U44053 (N_44053,N_42672,N_42493);
and U44054 (N_44054,N_42895,N_42289);
nand U44055 (N_44055,N_42241,N_42766);
xnor U44056 (N_44056,N_43852,N_43498);
and U44057 (N_44057,N_42225,N_43908);
xor U44058 (N_44058,N_42709,N_43904);
nand U44059 (N_44059,N_43964,N_43518);
nand U44060 (N_44060,N_43085,N_42815);
nand U44061 (N_44061,N_42753,N_42509);
xnor U44062 (N_44062,N_43909,N_43056);
nand U44063 (N_44063,N_42375,N_43869);
nor U44064 (N_44064,N_43539,N_43827);
or U44065 (N_44065,N_42695,N_42108);
nor U44066 (N_44066,N_42037,N_42626);
and U44067 (N_44067,N_42821,N_42540);
nand U44068 (N_44068,N_43658,N_43020);
and U44069 (N_44069,N_43585,N_43327);
or U44070 (N_44070,N_43763,N_42303);
nor U44071 (N_44071,N_42982,N_43080);
nor U44072 (N_44072,N_43530,N_43096);
and U44073 (N_44073,N_42066,N_43256);
nor U44074 (N_44074,N_43286,N_42332);
and U44075 (N_44075,N_43147,N_42044);
nor U44076 (N_44076,N_43741,N_43637);
xor U44077 (N_44077,N_43311,N_43355);
or U44078 (N_44078,N_42148,N_42909);
nor U44079 (N_44079,N_42294,N_43492);
or U44080 (N_44080,N_42595,N_42472);
or U44081 (N_44081,N_43662,N_42731);
nand U44082 (N_44082,N_43297,N_42577);
and U44083 (N_44083,N_43363,N_43136);
xor U44084 (N_44084,N_43600,N_43204);
or U44085 (N_44085,N_42388,N_42207);
and U44086 (N_44086,N_42206,N_43734);
nand U44087 (N_44087,N_43007,N_43108);
and U44088 (N_44088,N_43373,N_43850);
nand U44089 (N_44089,N_43198,N_43239);
nand U44090 (N_44090,N_43451,N_43686);
xnor U44091 (N_44091,N_43873,N_43026);
nand U44092 (N_44092,N_42308,N_43169);
xor U44093 (N_44093,N_42845,N_43824);
nand U44094 (N_44094,N_42483,N_43454);
nand U44095 (N_44095,N_43302,N_43588);
nand U44096 (N_44096,N_42017,N_43197);
xnor U44097 (N_44097,N_43379,N_43409);
nor U44098 (N_44098,N_42350,N_42278);
and U44099 (N_44099,N_43482,N_43183);
and U44100 (N_44100,N_42746,N_43716);
nor U44101 (N_44101,N_42155,N_43092);
nand U44102 (N_44102,N_42410,N_43821);
nand U44103 (N_44103,N_43618,N_43107);
or U44104 (N_44104,N_43229,N_42224);
and U44105 (N_44105,N_42458,N_42946);
nor U44106 (N_44106,N_43898,N_43663);
nor U44107 (N_44107,N_43322,N_43341);
nand U44108 (N_44108,N_43926,N_43809);
and U44109 (N_44109,N_43677,N_43052);
nor U44110 (N_44110,N_43778,N_43913);
nand U44111 (N_44111,N_43729,N_43996);
or U44112 (N_44112,N_43856,N_42061);
nor U44113 (N_44113,N_42651,N_42187);
nand U44114 (N_44114,N_43217,N_43364);
and U44115 (N_44115,N_43737,N_43337);
nand U44116 (N_44116,N_43340,N_43562);
or U44117 (N_44117,N_42331,N_43049);
nand U44118 (N_44118,N_42670,N_42496);
nand U44119 (N_44119,N_42611,N_43615);
or U44120 (N_44120,N_42287,N_42751);
nor U44121 (N_44121,N_43865,N_43657);
and U44122 (N_44122,N_43782,N_42789);
nor U44123 (N_44123,N_42513,N_43034);
or U44124 (N_44124,N_43446,N_43621);
nor U44125 (N_44125,N_42129,N_42811);
nand U44126 (N_44126,N_42555,N_42414);
nand U44127 (N_44127,N_43649,N_42266);
and U44128 (N_44128,N_42014,N_42183);
nor U44129 (N_44129,N_42901,N_42352);
xor U44130 (N_44130,N_42271,N_42964);
xor U44131 (N_44131,N_43071,N_43383);
xor U44132 (N_44132,N_42416,N_42917);
and U44133 (N_44133,N_43829,N_42806);
or U44134 (N_44134,N_42981,N_43345);
nor U44135 (N_44135,N_42680,N_43119);
xor U44136 (N_44136,N_43911,N_43441);
and U44137 (N_44137,N_43845,N_43592);
and U44138 (N_44138,N_43287,N_43321);
nor U44139 (N_44139,N_42643,N_42074);
xor U44140 (N_44140,N_43491,N_43210);
nand U44141 (N_44141,N_43252,N_43805);
xnor U44142 (N_44142,N_42091,N_42443);
nor U44143 (N_44143,N_43786,N_43486);
nor U44144 (N_44144,N_42608,N_43074);
and U44145 (N_44145,N_42973,N_43481);
nor U44146 (N_44146,N_42311,N_43992);
xnor U44147 (N_44147,N_43211,N_43298);
nor U44148 (N_44148,N_42263,N_43509);
xor U44149 (N_44149,N_43106,N_42057);
or U44150 (N_44150,N_42320,N_43762);
or U44151 (N_44151,N_42329,N_43180);
or U44152 (N_44152,N_43253,N_42358);
xor U44153 (N_44153,N_42342,N_42046);
nor U44154 (N_44154,N_42433,N_43471);
and U44155 (N_44155,N_42599,N_43958);
nand U44156 (N_44156,N_43109,N_43613);
xor U44157 (N_44157,N_42005,N_42052);
or U44158 (N_44158,N_43468,N_43124);
nand U44159 (N_44159,N_42393,N_43267);
xnor U44160 (N_44160,N_42843,N_42879);
and U44161 (N_44161,N_42231,N_43861);
or U44162 (N_44162,N_42137,N_42465);
and U44163 (N_44163,N_42010,N_43334);
nor U44164 (N_44164,N_43469,N_43921);
nor U44165 (N_44165,N_42103,N_43555);
xor U44166 (N_44166,N_42777,N_43245);
nand U44167 (N_44167,N_42162,N_43652);
nand U44168 (N_44168,N_43569,N_43848);
xor U44169 (N_44169,N_43366,N_43301);
xor U44170 (N_44170,N_42424,N_43430);
nor U44171 (N_44171,N_42796,N_42988);
or U44172 (N_44172,N_43214,N_43384);
or U44173 (N_44173,N_43354,N_42243);
nand U44174 (N_44174,N_42684,N_42693);
and U44175 (N_44175,N_42211,N_43917);
or U44176 (N_44176,N_43015,N_43342);
or U44177 (N_44177,N_42253,N_43416);
or U44178 (N_44178,N_43715,N_43113);
xor U44179 (N_44179,N_42671,N_43041);
or U44180 (N_44180,N_43171,N_43771);
nand U44181 (N_44181,N_42723,N_42788);
xor U44182 (N_44182,N_43360,N_43307);
and U44183 (N_44183,N_43859,N_43014);
or U44184 (N_44184,N_43993,N_42093);
and U44185 (N_44185,N_43292,N_43436);
nand U44186 (N_44186,N_43227,N_43804);
or U44187 (N_44187,N_42400,N_43619);
xnor U44188 (N_44188,N_42087,N_43756);
and U44189 (N_44189,N_42830,N_43439);
xor U44190 (N_44190,N_42560,N_43985);
or U44191 (N_44191,N_42043,N_43220);
and U44192 (N_44192,N_43522,N_43099);
nor U44193 (N_44193,N_42778,N_42374);
nor U44194 (N_44194,N_42118,N_42242);
or U44195 (N_44195,N_43487,N_42854);
nor U44196 (N_44196,N_43808,N_42404);
nand U44197 (N_44197,N_42954,N_42482);
xnor U44198 (N_44198,N_43224,N_43023);
and U44199 (N_44199,N_43403,N_43419);
xnor U44200 (N_44200,N_42967,N_42564);
nand U44201 (N_44201,N_43378,N_43701);
nor U44202 (N_44202,N_43513,N_42025);
nor U44203 (N_44203,N_43058,N_43453);
nand U44204 (N_44204,N_42034,N_42545);
nor U44205 (N_44205,N_43931,N_43694);
nand U44206 (N_44206,N_43117,N_43676);
and U44207 (N_44207,N_43777,N_42318);
or U44208 (N_44208,N_43779,N_43192);
xor U44209 (N_44209,N_42543,N_42857);
xor U44210 (N_44210,N_42239,N_42488);
xor U44211 (N_44211,N_42182,N_42171);
nand U44212 (N_44212,N_43488,N_43900);
and U44213 (N_44213,N_43775,N_42411);
nand U44214 (N_44214,N_42547,N_42609);
and U44215 (N_44215,N_42473,N_43554);
and U44216 (N_44216,N_42196,N_42570);
and U44217 (N_44217,N_43170,N_43063);
xnor U44218 (N_44218,N_43101,N_43280);
and U44219 (N_44219,N_42996,N_42268);
xor U44220 (N_44220,N_43235,N_43590);
nand U44221 (N_44221,N_42624,N_43942);
nor U44222 (N_44222,N_43402,N_42346);
xor U44223 (N_44223,N_42568,N_43371);
nand U44224 (N_44224,N_42924,N_43202);
nand U44225 (N_44225,N_43262,N_42667);
or U44226 (N_44226,N_42498,N_43382);
nor U44227 (N_44227,N_42556,N_43306);
and U44228 (N_44228,N_42313,N_42164);
and U44229 (N_44229,N_43651,N_42081);
xor U44230 (N_44230,N_42640,N_42689);
or U44231 (N_44231,N_42180,N_43673);
or U44232 (N_44232,N_42152,N_43250);
and U44233 (N_44233,N_42158,N_42461);
nor U44234 (N_44234,N_42665,N_42076);
or U44235 (N_44235,N_42480,N_43995);
or U44236 (N_44236,N_43027,N_42885);
or U44237 (N_44237,N_42732,N_42519);
and U44238 (N_44238,N_42307,N_43690);
nor U44239 (N_44239,N_42112,N_43244);
xnor U44240 (N_44240,N_42219,N_43547);
nand U44241 (N_44241,N_43104,N_43294);
nand U44242 (N_44242,N_43698,N_42551);
or U44243 (N_44243,N_42584,N_43391);
xor U44244 (N_44244,N_43485,N_43659);
and U44245 (N_44245,N_43418,N_42676);
or U44246 (N_44246,N_42745,N_42386);
or U44247 (N_44247,N_42250,N_43500);
or U44248 (N_44248,N_42537,N_42150);
and U44249 (N_44249,N_42698,N_42997);
nand U44250 (N_44250,N_43794,N_43123);
or U44251 (N_44251,N_42062,N_43664);
nor U44252 (N_44252,N_43427,N_42985);
and U44253 (N_44253,N_43291,N_42541);
and U44254 (N_44254,N_43024,N_42869);
and U44255 (N_44255,N_43512,N_43377);
xnor U44256 (N_44256,N_42256,N_42455);
or U44257 (N_44257,N_42507,N_42705);
nand U44258 (N_44258,N_43495,N_42628);
nand U44259 (N_44259,N_42944,N_42492);
or U44260 (N_44260,N_42515,N_42644);
or U44261 (N_44261,N_42317,N_42856);
nand U44262 (N_44262,N_43447,N_43178);
and U44263 (N_44263,N_42549,N_43514);
nor U44264 (N_44264,N_43066,N_42450);
nor U44265 (N_44265,N_43432,N_43986);
xor U44266 (N_44266,N_43744,N_42774);
xor U44267 (N_44267,N_43784,N_42649);
xor U44268 (N_44268,N_42340,N_42284);
nand U44269 (N_44269,N_42097,N_43184);
xnor U44270 (N_44270,N_42032,N_43857);
nor U44271 (N_44271,N_42696,N_42657);
and U44272 (N_44272,N_42726,N_42362);
or U44273 (N_44273,N_42001,N_43628);
xor U44274 (N_44274,N_43893,N_42781);
or U44275 (N_44275,N_42664,N_42491);
or U44276 (N_44276,N_42136,N_42855);
nor U44277 (N_44277,N_42893,N_43017);
nand U44278 (N_44278,N_42446,N_42502);
nand U44279 (N_44279,N_43589,N_42073);
nand U44280 (N_44280,N_43933,N_43271);
nor U44281 (N_44281,N_43497,N_42953);
nor U44282 (N_44282,N_42528,N_43002);
xnor U44283 (N_44283,N_42286,N_43974);
xor U44284 (N_44284,N_42166,N_42396);
and U44285 (N_44285,N_43200,N_42272);
xnor U44286 (N_44286,N_42026,N_42399);
nor U44287 (N_44287,N_42487,N_43067);
nor U44288 (N_44288,N_43381,N_43352);
xnor U44289 (N_44289,N_43179,N_43526);
xor U44290 (N_44290,N_42531,N_42316);
nor U44291 (N_44291,N_42526,N_43790);
xor U44292 (N_44292,N_42712,N_43255);
nand U44293 (N_44293,N_43632,N_42762);
or U44294 (N_44294,N_42096,N_42356);
and U44295 (N_44295,N_42435,N_42058);
xnor U44296 (N_44296,N_43475,N_42601);
and U44297 (N_44297,N_42120,N_43710);
or U44298 (N_44298,N_43639,N_43733);
xnor U44299 (N_44299,N_43043,N_42558);
or U44300 (N_44300,N_42776,N_43112);
xor U44301 (N_44301,N_43838,N_42823);
and U44302 (N_44302,N_42629,N_43358);
xor U44303 (N_44303,N_42425,N_42474);
xnor U44304 (N_44304,N_42993,N_43506);
xor U44305 (N_44305,N_42191,N_42138);
xnor U44306 (N_44306,N_43479,N_43781);
and U44307 (N_44307,N_43279,N_42792);
nand U44308 (N_44308,N_43039,N_43937);
or U44309 (N_44309,N_43718,N_42517);
or U44310 (N_44310,N_42963,N_43187);
and U44311 (N_44311,N_42758,N_43830);
nor U44312 (N_44312,N_43415,N_42775);
xnor U44313 (N_44313,N_42153,N_43152);
xor U44314 (N_44314,N_43455,N_43438);
nor U44315 (N_44315,N_42983,N_42991);
xor U44316 (N_44316,N_42970,N_43413);
or U44317 (N_44317,N_43646,N_42791);
nand U44318 (N_44318,N_42839,N_43584);
nor U44319 (N_44319,N_43444,N_42754);
nand U44320 (N_44320,N_42619,N_42139);
and U44321 (N_44321,N_42865,N_43233);
nand U44322 (N_44322,N_43703,N_42064);
nand U44323 (N_44323,N_43702,N_42102);
and U44324 (N_44324,N_42932,N_43412);
xor U44325 (N_44325,N_42960,N_42500);
nor U44326 (N_44326,N_43385,N_42593);
and U44327 (N_44327,N_43330,N_42617);
or U44328 (N_44328,N_43496,N_43994);
or U44329 (N_44329,N_43470,N_42189);
nor U44330 (N_44330,N_42589,N_43392);
xor U44331 (N_44331,N_42451,N_42955);
or U44332 (N_44332,N_43797,N_42548);
nand U44333 (N_44333,N_43213,N_43671);
and U44334 (N_44334,N_43816,N_43094);
and U44335 (N_44335,N_43625,N_43563);
nand U44336 (N_44336,N_42975,N_42801);
nand U44337 (N_44337,N_43837,N_42008);
nor U44338 (N_44338,N_43435,N_42992);
and U44339 (N_44339,N_42221,N_43407);
nand U44340 (N_44340,N_42562,N_42656);
and U44341 (N_44341,N_42477,N_43230);
or U44342 (N_44342,N_43886,N_42020);
and U44343 (N_44343,N_42710,N_43815);
and U44344 (N_44344,N_43174,N_42004);
nand U44345 (N_44345,N_42625,N_42898);
xnor U44346 (N_44346,N_43802,N_43343);
nand U44347 (N_44347,N_43967,N_42929);
or U44348 (N_44348,N_43708,N_42795);
xnor U44349 (N_44349,N_43743,N_43350);
xor U44350 (N_44350,N_42117,N_43299);
or U44351 (N_44351,N_43054,N_42161);
and U44352 (N_44352,N_42002,N_43987);
nand U44353 (N_44353,N_43564,N_42718);
xnor U44354 (N_44354,N_42510,N_43687);
xor U44355 (N_44355,N_43949,N_42038);
or U44356 (N_44356,N_42372,N_43818);
or U44357 (N_44357,N_43194,N_42700);
xor U44358 (N_44358,N_42169,N_43654);
or U44359 (N_44359,N_42438,N_43776);
nor U44360 (N_44360,N_43285,N_42395);
or U44361 (N_44361,N_43141,N_43983);
xnor U44362 (N_44362,N_42867,N_42021);
nand U44363 (N_44363,N_42273,N_43568);
and U44364 (N_44364,N_42916,N_43059);
or U44365 (N_44365,N_43357,N_42456);
xnor U44366 (N_44366,N_42614,N_43329);
xnor U44367 (N_44367,N_43275,N_42522);
nand U44368 (N_44368,N_43605,N_42304);
or U44369 (N_44369,N_43519,N_42323);
xnor U44370 (N_44370,N_42333,N_43847);
or U44371 (N_44371,N_43550,N_43612);
or U44372 (N_44372,N_43901,N_43713);
and U44373 (N_44373,N_43839,N_43616);
and U44374 (N_44374,N_42943,N_43855);
and U44375 (N_44375,N_42602,N_43156);
nor U44376 (N_44376,N_43507,N_42974);
or U44377 (N_44377,N_42381,N_42029);
nor U44378 (N_44378,N_42508,N_43305);
and U44379 (N_44379,N_43951,N_42623);
or U44380 (N_44380,N_42581,N_42367);
xnor U44381 (N_44381,N_43450,N_42053);
nor U44382 (N_44382,N_42279,N_42125);
xnor U44383 (N_44383,N_42244,N_42188);
xor U44384 (N_44384,N_42725,N_43158);
and U44385 (N_44385,N_42334,N_42178);
nor U44386 (N_44386,N_43751,N_43667);
nor U44387 (N_44387,N_43780,N_43560);
or U44388 (N_44388,N_42322,N_42530);
or U44389 (N_44389,N_43989,N_42663);
nand U44390 (N_44390,N_42337,N_43164);
nor U44391 (N_44391,N_42747,N_42047);
xor U44392 (N_44392,N_42486,N_42588);
and U44393 (N_44393,N_42878,N_42765);
nor U44394 (N_44394,N_42220,N_43546);
nand U44395 (N_44395,N_42195,N_42165);
nand U44396 (N_44396,N_42605,N_42921);
nor U44397 (N_44397,N_43396,N_43249);
and U44398 (N_44398,N_42230,N_43796);
nor U44399 (N_44399,N_43927,N_42172);
or U44400 (N_44400,N_43361,N_43871);
nor U44401 (N_44401,N_42694,N_43793);
nor U44402 (N_44402,N_43312,N_42704);
or U44403 (N_44403,N_42658,N_43541);
or U44404 (N_44404,N_42084,N_43408);
nor U44405 (N_44405,N_43160,N_43903);
nand U44406 (N_44406,N_43966,N_42086);
nor U44407 (N_44407,N_42301,N_42679);
nand U44408 (N_44408,N_42742,N_42802);
nor U44409 (N_44409,N_43095,N_42730);
and U44410 (N_44410,N_43005,N_42756);
nor U44411 (N_44411,N_43699,N_43760);
or U44412 (N_44412,N_43785,N_43072);
nand U44413 (N_44413,N_42524,N_43073);
xnor U44414 (N_44414,N_42685,N_42354);
xnor U44415 (N_44415,N_42585,N_43878);
nor U44416 (N_44416,N_42706,N_43190);
nand U44417 (N_44417,N_43222,N_43707);
nand U44418 (N_44418,N_42627,N_43902);
xor U44419 (N_44419,N_42262,N_42699);
or U44420 (N_44420,N_42719,N_43528);
nor U44421 (N_44421,N_42210,N_43304);
nor U44422 (N_44422,N_43689,N_43772);
nand U44423 (N_44423,N_42222,N_42807);
nor U44424 (N_44424,N_42941,N_43248);
or U44425 (N_44425,N_42145,N_42361);
nand U44426 (N_44426,N_43320,N_43314);
and U44427 (N_44427,N_42054,N_43883);
and U44428 (N_44428,N_43181,N_43945);
nor U44429 (N_44429,N_43484,N_43051);
or U44430 (N_44430,N_42914,N_43088);
nor U44431 (N_44431,N_43380,N_42060);
or U44432 (N_44432,N_43142,N_42597);
and U44433 (N_44433,N_42525,N_43128);
or U44434 (N_44434,N_42088,N_43581);
nand U44435 (N_44435,N_42969,N_43971);
xor U44436 (N_44436,N_43422,N_43650);
xnor U44437 (N_44437,N_43728,N_42896);
xor U44438 (N_44438,N_43807,N_42780);
or U44439 (N_44439,N_43736,N_43310);
and U44440 (N_44440,N_42767,N_42750);
nand U44441 (N_44441,N_43251,N_43918);
or U44442 (N_44442,N_42538,N_43161);
or U44443 (N_44443,N_43362,N_43932);
nand U44444 (N_44444,N_43114,N_42319);
or U44445 (N_44445,N_43452,N_42119);
and U44446 (N_44446,N_43692,N_42306);
or U44447 (N_44447,N_43278,N_42290);
or U44448 (N_44448,N_42124,N_42246);
nand U44449 (N_44449,N_43185,N_43876);
or U44450 (N_44450,N_42291,N_42205);
or U44451 (N_44451,N_43753,N_42234);
nor U44452 (N_44452,N_42883,N_43463);
nor U44453 (N_44453,N_43603,N_42764);
nand U44454 (N_44454,N_42380,N_42652);
nand U44455 (N_44455,N_42089,N_43511);
or U44456 (N_44456,N_42615,N_42849);
nor U44457 (N_44457,N_43565,N_43458);
nor U44458 (N_44458,N_43536,N_42407);
and U44459 (N_44459,N_43799,N_42134);
or U44460 (N_44460,N_42567,N_42907);
nand U44461 (N_44461,N_42733,N_42078);
or U44462 (N_44462,N_42714,N_43749);
nand U44463 (N_44463,N_43551,N_42877);
nand U44464 (N_44464,N_42460,N_42170);
nand U44465 (N_44465,N_42748,N_43100);
and U44466 (N_44466,N_43393,N_42258);
nor U44467 (N_44467,N_42420,N_42848);
nand U44468 (N_44468,N_43201,N_42606);
nand U44469 (N_44469,N_43765,N_42871);
or U44470 (N_44470,N_42464,N_43405);
xor U44471 (N_44471,N_42641,N_42419);
nand U44472 (N_44472,N_42655,N_43336);
and U44473 (N_44473,N_42797,N_42961);
xnor U44474 (N_44474,N_43188,N_42654);
nor U44475 (N_44475,N_43843,N_42912);
or U44476 (N_44476,N_42864,N_42804);
nor U44477 (N_44477,N_43527,N_43523);
and U44478 (N_44478,N_43466,N_42889);
xor U44479 (N_44479,N_43577,N_42554);
or U44480 (N_44480,N_43868,N_43397);
and U44481 (N_44481,N_43503,N_43905);
nor U44482 (N_44482,N_43508,N_43313);
nor U44483 (N_44483,N_43636,N_43315);
nand U44484 (N_44484,N_43448,N_43353);
nor U44485 (N_44485,N_42123,N_43277);
nor U44486 (N_44486,N_43236,N_43110);
xor U44487 (N_44487,N_42648,N_43060);
nand U44488 (N_44488,N_42413,N_43269);
xnor U44489 (N_44489,N_42031,N_42900);
and U44490 (N_44490,N_43831,N_42957);
or U44491 (N_44491,N_42862,N_43028);
or U44492 (N_44492,N_42484,N_43570);
and U44493 (N_44493,N_43189,N_43120);
xnor U44494 (N_44494,N_42666,N_42987);
and U44495 (N_44495,N_43062,N_43571);
nand U44496 (N_44496,N_42264,N_42434);
xor U44497 (N_44497,N_42927,N_42939);
nor U44498 (N_44498,N_42401,N_42343);
nand U44499 (N_44499,N_43610,N_43812);
and U44500 (N_44500,N_42637,N_42669);
xor U44501 (N_44501,N_43919,N_43151);
nand U44502 (N_44502,N_43691,N_43597);
nand U44503 (N_44503,N_42355,N_42280);
nand U44504 (N_44504,N_42270,N_42620);
and U44505 (N_44505,N_42906,N_43944);
or U44506 (N_44506,N_42716,N_43963);
or U44507 (N_44507,N_42514,N_43031);
nand U44508 (N_44508,N_42310,N_43638);
or U44509 (N_44509,N_42092,N_42398);
nand U44510 (N_44510,N_42378,N_42559);
nor U44511 (N_44511,N_42956,N_42978);
nor U44512 (N_44512,N_42986,N_42544);
nor U44513 (N_44513,N_43331,N_42126);
nor U44514 (N_44514,N_42977,N_42288);
and U44515 (N_44515,N_42905,N_43975);
and U44516 (N_44516,N_43356,N_42535);
and U44517 (N_44517,N_43787,N_43714);
and U44518 (N_44518,N_42837,N_43317);
nor U44519 (N_44519,N_43226,N_43042);
xor U44520 (N_44520,N_42505,N_42574);
and U44521 (N_44521,N_42633,N_42269);
nand U44522 (N_44522,N_43681,N_42759);
nor U44523 (N_44523,N_42635,N_42469);
nor U44524 (N_44524,N_42033,N_43449);
and U44525 (N_44525,N_43129,N_42740);
and U44526 (N_44526,N_43138,N_42768);
nand U44527 (N_44527,N_43711,N_43144);
or U44528 (N_44528,N_42937,N_42850);
xor U44529 (N_44529,N_42859,N_43629);
nor U44530 (N_44530,N_42049,N_42107);
and U44531 (N_44531,N_43719,N_43726);
or U44532 (N_44532,N_43425,N_43332);
or U44533 (N_44533,N_42866,N_43670);
xnor U44534 (N_44534,N_43293,N_42353);
xor U44535 (N_44535,N_43761,N_42293);
nor U44536 (N_44536,N_42703,N_42024);
or U44537 (N_44537,N_42377,N_42209);
xnor U44538 (N_44538,N_43602,N_43238);
nand U44539 (N_44539,N_42949,N_43961);
and U44540 (N_44540,N_43521,N_43344);
nor U44541 (N_44541,N_42887,N_43817);
nor U44542 (N_44542,N_42007,N_43084);
and U44543 (N_44543,N_43208,N_42818);
nand U44544 (N_44544,N_43437,N_43860);
xor U44545 (N_44545,N_43842,N_42412);
nor U44546 (N_44546,N_42415,N_42546);
or U44547 (N_44547,N_42405,N_43968);
nand U44548 (N_44548,N_42082,N_42813);
xor U44549 (N_44549,N_43135,N_43623);
nor U44550 (N_44550,N_43429,N_43607);
nand U44551 (N_44551,N_43578,N_42506);
xor U44552 (N_44552,N_42111,N_42051);
and U44553 (N_44553,N_42881,N_42952);
nor U44554 (N_44554,N_43205,N_42604);
nor U44555 (N_44555,N_43895,N_42143);
and U44556 (N_44556,N_43168,N_43770);
nand U44557 (N_44557,N_42387,N_42721);
and U44558 (N_44558,N_42841,N_43102);
and U44559 (N_44559,N_42245,N_42199);
and U44560 (N_44560,N_42891,N_43583);
nor U44561 (N_44561,N_42861,N_43599);
and U44562 (N_44562,N_42281,N_42995);
and U44563 (N_44563,N_42779,N_42520);
and U44564 (N_44564,N_43833,N_42444);
and U44565 (N_44565,N_43009,N_43624);
or U44566 (N_44566,N_42418,N_42448);
and U44567 (N_44567,N_43093,N_43849);
nor U44568 (N_44568,N_43960,N_42561);
nand U44569 (N_44569,N_43376,N_43685);
nand U44570 (N_44570,N_42233,N_42922);
nor U44571 (N_44571,N_42067,N_43001);
nor U44572 (N_44572,N_43853,N_42382);
nor U44573 (N_44573,N_43127,N_43572);
or U44574 (N_44574,N_42432,N_42140);
and U44575 (N_44575,N_43081,N_43851);
xnor U44576 (N_44576,N_43955,N_42527);
xnor U44577 (N_44577,N_43609,N_43411);
nor U44578 (N_44578,N_43389,N_42575);
and U44579 (N_44579,N_42232,N_43011);
nor U44580 (N_44580,N_42392,N_42471);
nand U44581 (N_44581,N_43648,N_42594);
nor U44582 (N_44582,N_43981,N_43622);
and U44583 (N_44583,N_43423,N_43899);
or U44584 (N_44584,N_43553,N_42799);
nor U44585 (N_44585,N_43630,N_42782);
nand U44586 (N_44586,N_42336,N_42744);
nor U44587 (N_44587,N_42638,N_42890);
nand U44588 (N_44588,N_43035,N_42908);
nor U44589 (N_44589,N_43055,N_43083);
and U44590 (N_44590,N_42330,N_42133);
xor U44591 (N_44591,N_42098,N_43678);
xnor U44592 (N_44592,N_42351,N_43490);
and U44593 (N_44593,N_42447,N_43494);
or U44594 (N_44594,N_42834,N_43272);
nand U44595 (N_44595,N_43791,N_43957);
nand U44596 (N_44596,N_43505,N_43395);
or U44597 (N_44597,N_43999,N_43727);
and U44598 (N_44598,N_42204,N_43929);
xnor U44599 (N_44599,N_42100,N_43349);
nand U44600 (N_44600,N_42565,N_43406);
nor U44601 (N_44601,N_43617,N_43973);
xor U44602 (N_44602,N_43032,N_43019);
xor U44603 (N_44603,N_42176,N_43165);
and U44604 (N_44604,N_43587,N_43982);
and U44605 (N_44605,N_42065,N_43745);
nand U44606 (N_44606,N_42736,N_42179);
or U44607 (N_44607,N_43643,N_43367);
and U44608 (N_44608,N_42613,N_42639);
or U44609 (N_44609,N_43295,N_42426);
nand U44610 (N_44610,N_42453,N_43155);
nor U44611 (N_44611,N_43875,N_42192);
nand U44612 (N_44612,N_43400,N_42662);
nand U44613 (N_44613,N_43910,N_43950);
and U44614 (N_44614,N_43724,N_43390);
nand U44615 (N_44615,N_42926,N_42772);
or U44616 (N_44616,N_43064,N_43757);
or U44617 (N_44617,N_42872,N_43025);
or U44618 (N_44618,N_43207,N_43149);
nand U44619 (N_44619,N_43533,N_43328);
or U44620 (N_44620,N_43467,N_43567);
nand U44621 (N_44621,N_42851,N_43754);
nor U44622 (N_44622,N_43348,N_42072);
nor U44623 (N_44623,N_42177,N_43087);
and U44624 (N_44624,N_43076,N_42452);
and U44625 (N_44625,N_43022,N_43697);
or U44626 (N_44626,N_43282,N_43215);
nand U44627 (N_44627,N_43037,N_43811);
nor U44628 (N_44628,N_43140,N_43656);
and U44629 (N_44629,N_42128,N_43006);
nand U44630 (N_44630,N_43510,N_43596);
and U44631 (N_44631,N_43008,N_42299);
or U44632 (N_44632,N_43889,N_42490);
and U44633 (N_44633,N_43887,N_42587);
and U44634 (N_44634,N_43517,N_42724);
nand U44635 (N_44635,N_42571,N_43978);
xor U44636 (N_44636,N_43021,N_43132);
and U44637 (N_44637,N_43237,N_42884);
or U44638 (N_44638,N_42406,N_43626);
or U44639 (N_44639,N_43767,N_42022);
nand U44640 (N_44640,N_43862,N_43044);
nand U44641 (N_44641,N_42499,N_43029);
nor U44642 (N_44642,N_42142,N_42990);
nand U44643 (N_44643,N_43257,N_43137);
and U44644 (N_44644,N_42713,N_43604);
or U44645 (N_44645,N_42314,N_42532);
or U44646 (N_44646,N_42300,N_42852);
nand U44647 (N_44647,N_42784,N_42678);
xor U44648 (N_44648,N_43126,N_42292);
and U44649 (N_44649,N_42853,N_43679);
or U44650 (N_44650,N_42603,N_43046);
xor U44651 (N_44651,N_42586,N_43688);
nor U44652 (N_44652,N_43445,N_42173);
nor U44653 (N_44653,N_42113,N_42121);
and U44654 (N_44654,N_43665,N_43428);
xnor U44655 (N_44655,N_42550,N_42994);
and U44656 (N_44656,N_42394,N_42440);
or U44657 (N_44657,N_42247,N_42533);
and U44658 (N_44658,N_42181,N_43696);
or U44659 (N_44659,N_42563,N_42436);
xor U44660 (N_44660,N_43976,N_43426);
or U44661 (N_44661,N_42110,N_42911);
nand U44662 (N_44662,N_42831,N_42449);
and U44663 (N_44663,N_42370,N_42529);
nor U44664 (N_44664,N_43880,N_43977);
nand U44665 (N_44665,N_42494,N_42557);
and U44666 (N_44666,N_43247,N_42979);
or U44667 (N_44667,N_43801,N_42154);
xnor U44668 (N_44668,N_43048,N_43388);
xor U44669 (N_44669,N_43125,N_43943);
xnor U44670 (N_44670,N_42298,N_42105);
or U44671 (N_44671,N_42793,N_42735);
xor U44672 (N_44672,N_42214,N_42820);
xor U44673 (N_44673,N_43460,N_43456);
nand U44674 (N_44674,N_42833,N_42379);
or U44675 (N_44675,N_43813,N_42503);
xor U44676 (N_44676,N_42160,N_43525);
and U44677 (N_44677,N_43930,N_43800);
nor U44678 (N_44678,N_42368,N_43706);
nand U44679 (N_44679,N_43863,N_43433);
nand U44680 (N_44680,N_42836,N_42681);
or U44681 (N_44681,N_42030,N_42569);
or U44682 (N_44682,N_42276,N_42677);
nand U44683 (N_44683,N_42079,N_43274);
nor U44684 (N_44684,N_42015,N_42439);
nor U44685 (N_44685,N_43680,N_43134);
xor U44686 (N_44686,N_42376,N_42616);
or U44687 (N_44687,N_42069,N_43068);
xor U44688 (N_44688,N_43221,N_43891);
or U44689 (N_44689,N_43374,N_43065);
or U44690 (N_44690,N_43266,N_43683);
or U44691 (N_44691,N_43281,N_42003);
and U44692 (N_44692,N_42215,N_43948);
nand U44693 (N_44693,N_42094,N_42383);
or U44694 (N_44694,N_42325,N_42095);
or U44695 (N_44695,N_43877,N_43462);
nand U44696 (N_44696,N_42803,N_43309);
xor U44697 (N_44697,N_42156,N_43828);
or U44698 (N_44698,N_43300,N_43264);
nor U44699 (N_44699,N_43705,N_43846);
and U44700 (N_44700,N_42738,N_43674);
and U44701 (N_44701,N_43520,N_43725);
or U44702 (N_44702,N_42023,N_43644);
xor U44703 (N_44703,N_43882,N_43284);
nand U44704 (N_44704,N_42194,N_42431);
and U44705 (N_44705,N_43196,N_43789);
xnor U44706 (N_44706,N_42115,N_42200);
nand U44707 (N_44707,N_42326,N_43558);
or U44708 (N_44708,N_43258,N_42573);
nor U44709 (N_44709,N_42489,N_42013);
nand U44710 (N_44710,N_43231,N_42621);
and U44711 (N_44711,N_43182,N_42457);
xnor U44712 (N_44712,N_42168,N_42131);
or U44713 (N_44713,N_43410,N_42042);
xnor U44714 (N_44714,N_43593,N_42267);
or U44715 (N_44715,N_42213,N_42817);
nand U44716 (N_44716,N_42642,N_43537);
xnor U44717 (N_44717,N_43404,N_42265);
or U44718 (N_44718,N_42692,N_43038);
and U44719 (N_44719,N_42339,N_42958);
and U44720 (N_44720,N_42827,N_42868);
nand U44721 (N_44721,N_42968,N_42886);
nor U44722 (N_44722,N_43387,N_42835);
nand U44723 (N_44723,N_42203,N_43154);
nand U44724 (N_44724,N_43870,N_42282);
nor U44725 (N_44725,N_42686,N_43489);
xnor U44726 (N_44726,N_43268,N_42445);
nand U44727 (N_44727,N_42930,N_43465);
or U44728 (N_44728,N_42130,N_43959);
nor U44729 (N_44729,N_43086,N_42894);
and U44730 (N_44730,N_43296,N_43881);
nand U44731 (N_44731,N_42972,N_42976);
nor U44732 (N_44732,N_43979,N_42389);
or U44733 (N_44733,N_42363,N_42344);
or U44734 (N_44734,N_42910,N_43579);
xnor U44735 (N_44735,N_43823,N_42646);
nor U44736 (N_44736,N_43559,N_42783);
nand U44737 (N_44737,N_42312,N_43089);
and U44738 (N_44738,N_43834,N_43241);
xor U44739 (N_44739,N_42951,N_43070);
or U44740 (N_44740,N_42193,N_43122);
nand U44741 (N_44741,N_43693,N_43459);
xnor U44742 (N_44742,N_43682,N_42752);
xnor U44743 (N_44743,N_43946,N_43139);
nand U44744 (N_44744,N_42798,N_43499);
and U44745 (N_44745,N_43369,N_43368);
or U44746 (N_44746,N_43050,N_42104);
and U44747 (N_44747,N_43116,N_42252);
and U44748 (N_44748,N_43159,N_42965);
xor U44749 (N_44749,N_43606,N_42688);
nand U44750 (N_44750,N_42174,N_43273);
nor U44751 (N_44751,N_43111,N_42936);
nor U44752 (N_44752,N_42012,N_42701);
nand U44753 (N_44753,N_43263,N_43069);
xor U44754 (N_44754,N_42842,N_42892);
nor U44755 (N_44755,N_42846,N_43841);
and U44756 (N_44756,N_42647,N_42321);
or U44757 (N_44757,N_42045,N_43030);
nor U44758 (N_44758,N_42720,N_42632);
nand U44759 (N_44759,N_43323,N_43896);
xnor U44760 (N_44760,N_43243,N_42348);
or U44761 (N_44761,N_43552,N_42274);
xor U44762 (N_44762,N_43980,N_42357);
xor U44763 (N_44763,N_42141,N_43872);
nand U44764 (N_44764,N_43186,N_42430);
nand U44765 (N_44765,N_43634,N_43386);
xor U44766 (N_44766,N_42238,N_43346);
or U44767 (N_44767,N_42114,N_42583);
xnor U44768 (N_44768,N_43633,N_43835);
nand U44769 (N_44769,N_43752,N_43614);
xor U44770 (N_44770,N_42808,N_42328);
xnor U44771 (N_44771,N_42737,N_42645);
xnor U44772 (N_44772,N_43464,N_43091);
xor U44773 (N_44773,N_43561,N_42347);
and U44774 (N_44774,N_43566,N_42422);
or U44775 (N_44775,N_43940,N_42190);
xnor U44776 (N_44776,N_42495,N_42409);
nand U44777 (N_44777,N_42959,N_42260);
or U44778 (N_44778,N_42345,N_43783);
or U44779 (N_44779,N_43866,N_43653);
and U44780 (N_44780,N_43972,N_42366);
nand U44781 (N_44781,N_43529,N_43819);
xnor U44782 (N_44782,N_43004,N_43045);
nor U44783 (N_44783,N_43792,N_43143);
nor U44784 (N_44784,N_43885,N_43888);
xnor U44785 (N_44785,N_43611,N_42198);
xnor U44786 (N_44786,N_42743,N_43351);
or U44787 (N_44787,N_43907,N_42578);
nand U44788 (N_44788,N_42523,N_43668);
xor U44789 (N_44789,N_43121,N_42349);
and U44790 (N_44790,N_42309,N_43036);
xnor U44791 (N_44791,N_43574,N_43417);
and U44792 (N_44792,N_42534,N_42202);
nand U44793 (N_44793,N_43502,N_43175);
xor U44794 (N_44794,N_43746,N_42729);
xor U44795 (N_44795,N_42971,N_43684);
xnor U44796 (N_44796,N_43672,N_43476);
xor U44797 (N_44797,N_42228,N_42217);
nand U44798 (N_44798,N_43731,N_42579);
nor U44799 (N_44799,N_43620,N_43915);
and U44800 (N_44800,N_42844,N_42254);
nor U44801 (N_44801,N_43740,N_42184);
nor U44802 (N_44802,N_42324,N_43738);
and U44803 (N_44803,N_43954,N_42197);
or U44804 (N_44804,N_43324,N_42481);
nand U44805 (N_44805,N_43478,N_42760);
or U44806 (N_44806,N_43925,N_43131);
nand U44807 (N_44807,N_42673,N_42858);
nor U44808 (N_44808,N_42248,N_42683);
or U44809 (N_44809,N_42755,N_42832);
nand U44810 (N_44810,N_42159,N_42542);
and U44811 (N_44811,N_43133,N_43544);
xnor U44812 (N_44812,N_42315,N_42697);
and U44813 (N_44813,N_43641,N_43103);
nor U44814 (N_44814,N_43098,N_43012);
xnor U44815 (N_44815,N_43922,N_42459);
nand U44816 (N_44816,N_43421,N_43443);
xor U44817 (N_44817,N_43193,N_43661);
and U44818 (N_44818,N_42757,N_43914);
or U44819 (N_44819,N_43375,N_42016);
xor U44820 (N_44820,N_43399,N_42962);
and U44821 (N_44821,N_42167,N_43916);
and U44822 (N_44822,N_42470,N_42682);
nor U44823 (N_44823,N_43261,N_42786);
xor U44824 (N_44824,N_42668,N_43924);
nor U44825 (N_44825,N_42504,N_42218);
or U44826 (N_44826,N_43591,N_42934);
nor U44827 (N_44827,N_42255,N_43806);
nor U44828 (N_44828,N_42873,N_42948);
xor U44829 (N_44829,N_43700,N_42070);
and U44830 (N_44830,N_43242,N_43998);
or U44831 (N_44831,N_43755,N_43549);
nor U44832 (N_44832,N_43162,N_42277);
and U44833 (N_44833,N_43240,N_43556);
nand U44834 (N_44834,N_43635,N_42847);
nor U44835 (N_44835,N_43303,N_42146);
and U44836 (N_44836,N_42360,N_42186);
nand U44837 (N_44837,N_42497,N_43543);
or U44838 (N_44838,N_43372,N_42598);
xor U44839 (N_44839,N_42787,N_43172);
and U44840 (N_44840,N_43984,N_42945);
or U44841 (N_44841,N_42229,N_42902);
and U44842 (N_44842,N_42151,N_42819);
or U44843 (N_44843,N_42600,N_43316);
nor U44844 (N_44844,N_43398,N_43442);
xnor U44845 (N_44845,N_42516,N_42876);
and U44846 (N_44846,N_43938,N_42201);
or U44847 (N_44847,N_42660,N_42296);
and U44848 (N_44848,N_42226,N_42297);
nand U44849 (N_44849,N_43209,N_43308);
and U44850 (N_44850,N_43335,N_43260);
and U44851 (N_44851,N_43864,N_42984);
nor U44852 (N_44852,N_42998,N_42144);
nor U44853 (N_44853,N_43704,N_42980);
nand U44854 (N_44854,N_43166,N_43720);
nand U44855 (N_44855,N_42915,N_43840);
and U44856 (N_44856,N_42127,N_42338);
nor U44857 (N_44857,N_43601,N_42341);
or U44858 (N_44858,N_42364,N_42825);
xor U44859 (N_44859,N_43928,N_43894);
or U44860 (N_44860,N_43768,N_42630);
xnor U44861 (N_44861,N_43145,N_43440);
or U44862 (N_44862,N_42828,N_43290);
and U44863 (N_44863,N_43516,N_42283);
or U44864 (N_44864,N_43483,N_42812);
or U44865 (N_44865,N_43627,N_42675);
xor U44866 (N_44866,N_42099,N_43033);
nor U44867 (N_44867,N_43759,N_42591);
and U44868 (N_44868,N_43191,N_42702);
and U44869 (N_44869,N_42468,N_42785);
xor U44870 (N_44870,N_43203,N_43078);
xor U44871 (N_44871,N_42149,N_42036);
xor U44872 (N_44872,N_43825,N_43939);
or U44873 (N_44873,N_43956,N_43434);
nor U44874 (N_44874,N_42463,N_42942);
or U44875 (N_44875,N_43723,N_42653);
nor U44876 (N_44876,N_42552,N_42462);
xor U44877 (N_44877,N_42708,N_43788);
nor U44878 (N_44878,N_43097,N_42019);
xor U44879 (N_44879,N_43420,N_42285);
or U44880 (N_44880,N_43965,N_43473);
nand U44881 (N_44881,N_42055,N_42590);
nand U44882 (N_44882,N_42822,N_43493);
xor U44883 (N_44883,N_42920,N_42090);
xnor U44884 (N_44884,N_42622,N_43953);
or U44885 (N_44885,N_42080,N_42805);
xnor U44886 (N_44886,N_42369,N_42950);
nand U44887 (N_44887,N_43148,N_43748);
xnor U44888 (N_44888,N_43079,N_42631);
nor U44889 (N_44889,N_43047,N_43730);
nor U44890 (N_44890,N_42063,N_42071);
nor U44891 (N_44891,N_43747,N_43115);
or U44892 (N_44892,N_42770,N_42212);
xnor U44893 (N_44893,N_42476,N_42771);
nor U44894 (N_44894,N_42572,N_43167);
xor U44895 (N_44895,N_43540,N_42208);
nor U44896 (N_44896,N_43000,N_43105);
nand U44897 (N_44897,N_42650,N_43225);
nand U44898 (N_44898,N_42327,N_43090);
xor U44899 (N_44899,N_42302,N_43814);
or U44900 (N_44900,N_42000,N_43461);
nand U44901 (N_44901,N_42427,N_42923);
nor U44902 (N_44902,N_43997,N_43003);
xnor U44903 (N_44903,N_43163,N_43524);
xor U44904 (N_44904,N_43265,N_43477);
xor U44905 (N_44905,N_43803,N_43640);
xor U44906 (N_44906,N_42576,N_43655);
and U44907 (N_44907,N_43742,N_42612);
xor U44908 (N_44908,N_43118,N_42009);
nor U44909 (N_44909,N_42175,N_42903);
or U44910 (N_44910,N_43660,N_42442);
or U44911 (N_44911,N_42739,N_43766);
or U44912 (N_44912,N_42707,N_42512);
or U44913 (N_44913,N_43936,N_43318);
xnor U44914 (N_44914,N_42116,N_43820);
and U44915 (N_44915,N_42077,N_42478);
or U44916 (N_44916,N_42749,N_42257);
or U44917 (N_44917,N_43218,N_43769);
or U44918 (N_44918,N_43177,N_43890);
or U44919 (N_44919,N_42838,N_42305);
nor U44920 (N_44920,N_42935,N_42083);
nand U44921 (N_44921,N_42618,N_43480);
xnor U44922 (N_44922,N_42741,N_43173);
or U44923 (N_44923,N_43645,N_42711);
xor U44924 (N_44924,N_42335,N_43234);
nand U44925 (N_44925,N_42763,N_43832);
nand U44926 (N_44926,N_43858,N_43647);
nand U44927 (N_44927,N_42659,N_42467);
xor U44928 (N_44928,N_42397,N_42913);
xor U44929 (N_44929,N_42249,N_43501);
and U44930 (N_44930,N_42863,N_43557);
xor U44931 (N_44931,N_43319,N_42056);
nor U44932 (N_44932,N_42566,N_42251);
nor U44933 (N_44933,N_42947,N_42011);
or U44934 (N_44934,N_43822,N_43013);
nand U44935 (N_44935,N_42636,N_42018);
nand U44936 (N_44936,N_43874,N_43631);
nand U44937 (N_44937,N_43582,N_43594);
xnor U44938 (N_44938,N_42661,N_43472);
nand U44939 (N_44939,N_43232,N_43854);
or U44940 (N_44940,N_43276,N_42223);
xnor U44941 (N_44941,N_42466,N_43040);
nor U44942 (N_44942,N_43598,N_42582);
or U44943 (N_44943,N_43534,N_43057);
nor U44944 (N_44944,N_42925,N_42580);
nor U44945 (N_44945,N_43542,N_42235);
and U44946 (N_44946,N_43414,N_43941);
nand U44947 (N_44947,N_42874,N_42428);
xor U44948 (N_44948,N_42888,N_43199);
nand U44949 (N_44949,N_43223,N_42809);
and U44950 (N_44950,N_42109,N_43157);
and U44951 (N_44951,N_42840,N_43010);
and U44952 (N_44952,N_42050,N_42157);
nand U44953 (N_44953,N_42441,N_43326);
nor U44954 (N_44954,N_42408,N_42607);
nor U44955 (N_44955,N_43884,N_43082);
and U44956 (N_44956,N_43666,N_42006);
and U44957 (N_44957,N_43359,N_43246);
nor U44958 (N_44958,N_43016,N_42259);
nand U44959 (N_44959,N_43289,N_43130);
or U44960 (N_44960,N_43333,N_43879);
xnor U44961 (N_44961,N_42521,N_42875);
or U44962 (N_44962,N_43923,N_43739);
or U44963 (N_44963,N_42539,N_42040);
or U44964 (N_44964,N_42101,N_42048);
or U44965 (N_44965,N_42717,N_43338);
nor U44966 (N_44966,N_43798,N_42028);
or U44967 (N_44967,N_42536,N_42371);
nand U44968 (N_44968,N_43575,N_42596);
xnor U44969 (N_44969,N_43906,N_42147);
and U44970 (N_44970,N_42039,N_43675);
nor U44971 (N_44971,N_43773,N_42059);
or U44972 (N_44972,N_43535,N_43717);
nand U44973 (N_44973,N_43952,N_43548);
nand U44974 (N_44974,N_43431,N_43339);
nand U44975 (N_44975,N_42999,N_43061);
or U44976 (N_44976,N_42826,N_43531);
or U44977 (N_44977,N_42931,N_43947);
nor U44978 (N_44978,N_43897,N_43150);
xnor U44979 (N_44979,N_43836,N_42041);
and U44980 (N_44980,N_43538,N_42715);
and U44981 (N_44981,N_43212,N_42933);
and U44982 (N_44982,N_42423,N_42800);
and U44983 (N_44983,N_42185,N_43934);
and U44984 (N_44984,N_42824,N_43991);
and U44985 (N_44985,N_42359,N_42938);
xnor U44986 (N_44986,N_43573,N_42691);
xnor U44987 (N_44987,N_42634,N_43795);
and U44988 (N_44988,N_42391,N_42390);
xor U44989 (N_44989,N_43758,N_42485);
nand U44990 (N_44990,N_43153,N_43712);
nor U44991 (N_44991,N_43988,N_43474);
and U44992 (N_44992,N_42261,N_43721);
nand U44993 (N_44993,N_43365,N_42690);
or U44994 (N_44994,N_42075,N_43176);
or U44995 (N_44995,N_42897,N_42727);
or U44996 (N_44996,N_42275,N_42814);
or U44997 (N_44997,N_42135,N_42899);
xnor U44998 (N_44998,N_43920,N_43642);
nor U44999 (N_44999,N_43735,N_43075);
xnor U45000 (N_45000,N_43411,N_43975);
nor U45001 (N_45001,N_43601,N_42618);
xor U45002 (N_45002,N_43331,N_42050);
nand U45003 (N_45003,N_42774,N_42011);
xnor U45004 (N_45004,N_43457,N_42947);
and U45005 (N_45005,N_43730,N_43139);
and U45006 (N_45006,N_42350,N_42681);
or U45007 (N_45007,N_42940,N_42574);
or U45008 (N_45008,N_43659,N_43733);
xnor U45009 (N_45009,N_43854,N_42897);
or U45010 (N_45010,N_43485,N_42424);
and U45011 (N_45011,N_43283,N_43733);
or U45012 (N_45012,N_43882,N_42380);
xor U45013 (N_45013,N_43848,N_43937);
or U45014 (N_45014,N_43184,N_43796);
nand U45015 (N_45015,N_42263,N_43789);
and U45016 (N_45016,N_43334,N_43608);
and U45017 (N_45017,N_42515,N_43219);
xnor U45018 (N_45018,N_43193,N_42717);
xor U45019 (N_45019,N_42999,N_42022);
and U45020 (N_45020,N_42342,N_42391);
nand U45021 (N_45021,N_43832,N_42100);
xor U45022 (N_45022,N_43431,N_42710);
or U45023 (N_45023,N_43246,N_42875);
nand U45024 (N_45024,N_42002,N_43236);
and U45025 (N_45025,N_42970,N_43284);
xnor U45026 (N_45026,N_43009,N_42968);
xnor U45027 (N_45027,N_42631,N_42681);
nand U45028 (N_45028,N_43689,N_43678);
xnor U45029 (N_45029,N_42740,N_42937);
nor U45030 (N_45030,N_42687,N_42107);
nand U45031 (N_45031,N_43550,N_42193);
nor U45032 (N_45032,N_43408,N_42486);
and U45033 (N_45033,N_43852,N_42124);
and U45034 (N_45034,N_43998,N_43912);
nor U45035 (N_45035,N_43186,N_43005);
and U45036 (N_45036,N_42940,N_43360);
nand U45037 (N_45037,N_42458,N_42653);
nand U45038 (N_45038,N_42603,N_43196);
nor U45039 (N_45039,N_42617,N_43169);
nand U45040 (N_45040,N_42628,N_43434);
xnor U45041 (N_45041,N_43804,N_43576);
nor U45042 (N_45042,N_43239,N_43497);
nor U45043 (N_45043,N_42696,N_43779);
nand U45044 (N_45044,N_42389,N_42520);
or U45045 (N_45045,N_43631,N_42493);
nand U45046 (N_45046,N_43412,N_42709);
and U45047 (N_45047,N_42446,N_43035);
xnor U45048 (N_45048,N_43068,N_43975);
nand U45049 (N_45049,N_42249,N_42796);
xnor U45050 (N_45050,N_42702,N_43242);
or U45051 (N_45051,N_43900,N_42565);
nor U45052 (N_45052,N_42722,N_43071);
and U45053 (N_45053,N_43122,N_42797);
nor U45054 (N_45054,N_42855,N_43005);
or U45055 (N_45055,N_43970,N_42427);
and U45056 (N_45056,N_43352,N_43996);
or U45057 (N_45057,N_43160,N_42552);
or U45058 (N_45058,N_42527,N_43696);
or U45059 (N_45059,N_43095,N_43827);
or U45060 (N_45060,N_43052,N_42607);
or U45061 (N_45061,N_43108,N_42875);
or U45062 (N_45062,N_43636,N_42411);
nor U45063 (N_45063,N_42204,N_43809);
and U45064 (N_45064,N_42372,N_43069);
nor U45065 (N_45065,N_43012,N_43918);
nand U45066 (N_45066,N_42158,N_42421);
nand U45067 (N_45067,N_43557,N_43187);
and U45068 (N_45068,N_43898,N_43357);
and U45069 (N_45069,N_43474,N_43745);
nand U45070 (N_45070,N_42463,N_42761);
xnor U45071 (N_45071,N_43813,N_43071);
nor U45072 (N_45072,N_42365,N_43460);
nor U45073 (N_45073,N_42815,N_42603);
xor U45074 (N_45074,N_42654,N_42511);
nor U45075 (N_45075,N_43682,N_43212);
or U45076 (N_45076,N_42316,N_42759);
and U45077 (N_45077,N_42948,N_42237);
xor U45078 (N_45078,N_42883,N_43719);
nand U45079 (N_45079,N_42196,N_42987);
nor U45080 (N_45080,N_43057,N_43390);
or U45081 (N_45081,N_42997,N_43084);
nand U45082 (N_45082,N_43620,N_43867);
and U45083 (N_45083,N_43357,N_43477);
nor U45084 (N_45084,N_43437,N_42110);
nand U45085 (N_45085,N_42977,N_43754);
or U45086 (N_45086,N_43597,N_43712);
or U45087 (N_45087,N_42663,N_42542);
or U45088 (N_45088,N_43824,N_42149);
or U45089 (N_45089,N_42057,N_42718);
xnor U45090 (N_45090,N_43214,N_42894);
and U45091 (N_45091,N_43599,N_43293);
nor U45092 (N_45092,N_43831,N_42634);
or U45093 (N_45093,N_42847,N_43791);
xnor U45094 (N_45094,N_43645,N_43078);
nor U45095 (N_45095,N_43931,N_43863);
xnor U45096 (N_45096,N_43690,N_42312);
xor U45097 (N_45097,N_42190,N_43451);
xor U45098 (N_45098,N_43875,N_42000);
nor U45099 (N_45099,N_42558,N_42360);
nor U45100 (N_45100,N_42809,N_43940);
nand U45101 (N_45101,N_43279,N_43911);
or U45102 (N_45102,N_42944,N_42029);
and U45103 (N_45103,N_42189,N_42905);
or U45104 (N_45104,N_43077,N_42531);
xor U45105 (N_45105,N_43686,N_43145);
nand U45106 (N_45106,N_43691,N_43352);
nand U45107 (N_45107,N_42831,N_43743);
and U45108 (N_45108,N_42634,N_42197);
nor U45109 (N_45109,N_43614,N_43205);
or U45110 (N_45110,N_43407,N_42262);
and U45111 (N_45111,N_43657,N_42075);
and U45112 (N_45112,N_43875,N_42490);
and U45113 (N_45113,N_43282,N_43039);
or U45114 (N_45114,N_42395,N_43593);
nor U45115 (N_45115,N_42228,N_42702);
or U45116 (N_45116,N_42824,N_43473);
or U45117 (N_45117,N_42506,N_43771);
nand U45118 (N_45118,N_43584,N_42725);
nand U45119 (N_45119,N_43486,N_43891);
xnor U45120 (N_45120,N_42302,N_43124);
nor U45121 (N_45121,N_42454,N_43348);
nor U45122 (N_45122,N_42492,N_42173);
and U45123 (N_45123,N_42069,N_43611);
or U45124 (N_45124,N_42085,N_43476);
xnor U45125 (N_45125,N_43137,N_43487);
nor U45126 (N_45126,N_42027,N_42758);
nand U45127 (N_45127,N_42766,N_42173);
nand U45128 (N_45128,N_42011,N_43795);
or U45129 (N_45129,N_42911,N_43763);
and U45130 (N_45130,N_42062,N_42302);
nor U45131 (N_45131,N_43043,N_42492);
nor U45132 (N_45132,N_42023,N_43620);
xor U45133 (N_45133,N_42940,N_43814);
nand U45134 (N_45134,N_43865,N_43771);
xor U45135 (N_45135,N_43411,N_42419);
and U45136 (N_45136,N_43480,N_42919);
nand U45137 (N_45137,N_42189,N_43065);
or U45138 (N_45138,N_43488,N_43030);
xor U45139 (N_45139,N_43359,N_42843);
nor U45140 (N_45140,N_43280,N_43527);
xnor U45141 (N_45141,N_43253,N_42870);
and U45142 (N_45142,N_42950,N_42802);
xor U45143 (N_45143,N_42464,N_42848);
or U45144 (N_45144,N_43256,N_42976);
nor U45145 (N_45145,N_43304,N_43839);
or U45146 (N_45146,N_42653,N_43474);
and U45147 (N_45147,N_43691,N_43356);
xor U45148 (N_45148,N_43262,N_43369);
xor U45149 (N_45149,N_42776,N_43630);
xnor U45150 (N_45150,N_42117,N_43600);
or U45151 (N_45151,N_43852,N_42299);
and U45152 (N_45152,N_43945,N_43217);
nand U45153 (N_45153,N_42211,N_43777);
and U45154 (N_45154,N_43906,N_42956);
xnor U45155 (N_45155,N_42369,N_42210);
or U45156 (N_45156,N_43328,N_42634);
xor U45157 (N_45157,N_42275,N_42079);
nor U45158 (N_45158,N_42340,N_43074);
or U45159 (N_45159,N_43680,N_43465);
nor U45160 (N_45160,N_42839,N_43606);
and U45161 (N_45161,N_43338,N_42459);
xnor U45162 (N_45162,N_42980,N_42586);
xnor U45163 (N_45163,N_42874,N_43226);
xor U45164 (N_45164,N_43038,N_42286);
xor U45165 (N_45165,N_42150,N_42007);
and U45166 (N_45166,N_43912,N_42019);
xnor U45167 (N_45167,N_43492,N_42702);
or U45168 (N_45168,N_43829,N_42311);
xnor U45169 (N_45169,N_42005,N_43524);
nor U45170 (N_45170,N_42679,N_43922);
xnor U45171 (N_45171,N_42270,N_43590);
nand U45172 (N_45172,N_43632,N_42192);
and U45173 (N_45173,N_43906,N_43472);
and U45174 (N_45174,N_42508,N_43283);
nor U45175 (N_45175,N_42803,N_42548);
xnor U45176 (N_45176,N_42554,N_42399);
or U45177 (N_45177,N_42368,N_42889);
nor U45178 (N_45178,N_42608,N_43830);
nand U45179 (N_45179,N_43936,N_43788);
or U45180 (N_45180,N_43626,N_43686);
nor U45181 (N_45181,N_43089,N_43406);
nand U45182 (N_45182,N_42052,N_42779);
or U45183 (N_45183,N_43566,N_42909);
xnor U45184 (N_45184,N_42938,N_42807);
or U45185 (N_45185,N_42999,N_42857);
nand U45186 (N_45186,N_43138,N_42835);
or U45187 (N_45187,N_43190,N_42112);
xor U45188 (N_45188,N_43805,N_43211);
nor U45189 (N_45189,N_43879,N_42511);
xnor U45190 (N_45190,N_43376,N_42926);
nand U45191 (N_45191,N_43268,N_43036);
nor U45192 (N_45192,N_42900,N_42634);
and U45193 (N_45193,N_42764,N_42661);
nor U45194 (N_45194,N_42319,N_42221);
nand U45195 (N_45195,N_42291,N_42721);
xnor U45196 (N_45196,N_42055,N_42990);
or U45197 (N_45197,N_42226,N_43871);
nand U45198 (N_45198,N_42748,N_42786);
or U45199 (N_45199,N_42009,N_42856);
or U45200 (N_45200,N_42150,N_42248);
nor U45201 (N_45201,N_43059,N_43661);
nand U45202 (N_45202,N_43699,N_43107);
xnor U45203 (N_45203,N_42540,N_42340);
or U45204 (N_45204,N_43860,N_42274);
nand U45205 (N_45205,N_42585,N_42895);
nand U45206 (N_45206,N_42996,N_42373);
nand U45207 (N_45207,N_42666,N_42908);
xor U45208 (N_45208,N_42692,N_43952);
or U45209 (N_45209,N_42872,N_42729);
or U45210 (N_45210,N_42705,N_42491);
xor U45211 (N_45211,N_43023,N_43621);
nand U45212 (N_45212,N_43223,N_42127);
xor U45213 (N_45213,N_42389,N_43224);
and U45214 (N_45214,N_43263,N_42884);
nor U45215 (N_45215,N_42566,N_43145);
xnor U45216 (N_45216,N_43581,N_43425);
xnor U45217 (N_45217,N_42632,N_43655);
nor U45218 (N_45218,N_42067,N_43410);
or U45219 (N_45219,N_43892,N_42565);
and U45220 (N_45220,N_43442,N_42099);
nand U45221 (N_45221,N_42597,N_42145);
nand U45222 (N_45222,N_43243,N_42190);
and U45223 (N_45223,N_42279,N_42090);
nor U45224 (N_45224,N_42081,N_43584);
and U45225 (N_45225,N_43298,N_43743);
nor U45226 (N_45226,N_42887,N_43818);
nand U45227 (N_45227,N_43276,N_42511);
xnor U45228 (N_45228,N_43863,N_42454);
xor U45229 (N_45229,N_42213,N_42787);
and U45230 (N_45230,N_43644,N_43941);
and U45231 (N_45231,N_42228,N_42170);
and U45232 (N_45232,N_43047,N_42842);
nand U45233 (N_45233,N_43463,N_43913);
xnor U45234 (N_45234,N_43250,N_42430);
nor U45235 (N_45235,N_42669,N_42583);
nor U45236 (N_45236,N_42129,N_43312);
or U45237 (N_45237,N_43830,N_43144);
or U45238 (N_45238,N_43118,N_42070);
and U45239 (N_45239,N_42582,N_42523);
and U45240 (N_45240,N_43410,N_43408);
xor U45241 (N_45241,N_43012,N_43306);
nor U45242 (N_45242,N_43772,N_43649);
or U45243 (N_45243,N_42078,N_43173);
or U45244 (N_45244,N_42092,N_43246);
or U45245 (N_45245,N_42486,N_42605);
nand U45246 (N_45246,N_42288,N_43340);
and U45247 (N_45247,N_43493,N_43149);
nand U45248 (N_45248,N_42462,N_42061);
or U45249 (N_45249,N_42747,N_42929);
or U45250 (N_45250,N_43886,N_43021);
xor U45251 (N_45251,N_43153,N_43576);
and U45252 (N_45252,N_42880,N_42112);
nor U45253 (N_45253,N_42148,N_43863);
nor U45254 (N_45254,N_43532,N_42168);
or U45255 (N_45255,N_43210,N_42313);
and U45256 (N_45256,N_43766,N_43425);
and U45257 (N_45257,N_43603,N_42118);
and U45258 (N_45258,N_42022,N_42004);
or U45259 (N_45259,N_43068,N_42763);
nand U45260 (N_45260,N_43472,N_42183);
and U45261 (N_45261,N_42792,N_42411);
xnor U45262 (N_45262,N_43474,N_43312);
or U45263 (N_45263,N_43147,N_43960);
nor U45264 (N_45264,N_43875,N_43416);
xnor U45265 (N_45265,N_43533,N_43916);
nor U45266 (N_45266,N_43868,N_43965);
nor U45267 (N_45267,N_43117,N_42131);
xor U45268 (N_45268,N_43593,N_42208);
nor U45269 (N_45269,N_43795,N_42642);
or U45270 (N_45270,N_43974,N_43997);
or U45271 (N_45271,N_43875,N_42925);
nand U45272 (N_45272,N_42752,N_43347);
xnor U45273 (N_45273,N_43640,N_42328);
nor U45274 (N_45274,N_43954,N_43159);
and U45275 (N_45275,N_42637,N_43634);
or U45276 (N_45276,N_43457,N_42687);
nand U45277 (N_45277,N_43757,N_42019);
nand U45278 (N_45278,N_43223,N_42738);
nor U45279 (N_45279,N_42264,N_43200);
and U45280 (N_45280,N_42350,N_42904);
nand U45281 (N_45281,N_43073,N_43691);
nand U45282 (N_45282,N_43451,N_43942);
nand U45283 (N_45283,N_42202,N_43429);
xnor U45284 (N_45284,N_43121,N_42653);
and U45285 (N_45285,N_43456,N_43793);
or U45286 (N_45286,N_43137,N_42214);
or U45287 (N_45287,N_42849,N_43538);
or U45288 (N_45288,N_43834,N_43178);
or U45289 (N_45289,N_43968,N_43085);
nand U45290 (N_45290,N_43703,N_43872);
xnor U45291 (N_45291,N_43221,N_43547);
and U45292 (N_45292,N_43981,N_42708);
and U45293 (N_45293,N_42293,N_43476);
or U45294 (N_45294,N_43540,N_43858);
xor U45295 (N_45295,N_43803,N_42239);
and U45296 (N_45296,N_43750,N_43085);
xor U45297 (N_45297,N_43808,N_42435);
nor U45298 (N_45298,N_42849,N_43235);
nor U45299 (N_45299,N_43662,N_42233);
or U45300 (N_45300,N_42128,N_42761);
or U45301 (N_45301,N_43562,N_43479);
xor U45302 (N_45302,N_43552,N_42852);
or U45303 (N_45303,N_42797,N_42097);
nand U45304 (N_45304,N_43692,N_43235);
xor U45305 (N_45305,N_42715,N_42341);
nor U45306 (N_45306,N_43804,N_43233);
or U45307 (N_45307,N_42642,N_42651);
xor U45308 (N_45308,N_43347,N_43216);
nand U45309 (N_45309,N_43184,N_43678);
and U45310 (N_45310,N_42295,N_42022);
and U45311 (N_45311,N_42142,N_42872);
nor U45312 (N_45312,N_42790,N_42406);
nor U45313 (N_45313,N_42954,N_43005);
and U45314 (N_45314,N_43407,N_42048);
nand U45315 (N_45315,N_42057,N_42563);
nand U45316 (N_45316,N_42296,N_42781);
or U45317 (N_45317,N_42337,N_43613);
xor U45318 (N_45318,N_42210,N_43229);
or U45319 (N_45319,N_43243,N_43683);
or U45320 (N_45320,N_42408,N_43980);
nor U45321 (N_45321,N_42238,N_42062);
xor U45322 (N_45322,N_42820,N_43384);
or U45323 (N_45323,N_42355,N_43604);
or U45324 (N_45324,N_42270,N_42458);
nor U45325 (N_45325,N_43094,N_43794);
nor U45326 (N_45326,N_43824,N_42009);
nor U45327 (N_45327,N_43626,N_42568);
xor U45328 (N_45328,N_42890,N_42718);
or U45329 (N_45329,N_43577,N_43250);
and U45330 (N_45330,N_43644,N_43585);
nor U45331 (N_45331,N_42279,N_43706);
xnor U45332 (N_45332,N_42598,N_43256);
and U45333 (N_45333,N_42438,N_43384);
nand U45334 (N_45334,N_42310,N_43204);
nor U45335 (N_45335,N_42479,N_43556);
or U45336 (N_45336,N_43131,N_42556);
xnor U45337 (N_45337,N_43506,N_42248);
nand U45338 (N_45338,N_42366,N_42467);
xnor U45339 (N_45339,N_42302,N_43448);
nor U45340 (N_45340,N_43155,N_42585);
nand U45341 (N_45341,N_42163,N_43226);
and U45342 (N_45342,N_42590,N_42506);
and U45343 (N_45343,N_43578,N_43911);
nor U45344 (N_45344,N_43925,N_43236);
nor U45345 (N_45345,N_43145,N_43350);
nor U45346 (N_45346,N_42369,N_43364);
and U45347 (N_45347,N_43669,N_42581);
or U45348 (N_45348,N_42291,N_42915);
or U45349 (N_45349,N_42763,N_42701);
nor U45350 (N_45350,N_42281,N_43786);
or U45351 (N_45351,N_42790,N_42070);
nand U45352 (N_45352,N_43118,N_42030);
xnor U45353 (N_45353,N_42274,N_43160);
xor U45354 (N_45354,N_42637,N_42667);
nand U45355 (N_45355,N_43158,N_43305);
nor U45356 (N_45356,N_43672,N_43905);
and U45357 (N_45357,N_43190,N_42403);
xnor U45358 (N_45358,N_43228,N_42845);
nor U45359 (N_45359,N_43939,N_42041);
xnor U45360 (N_45360,N_43595,N_42873);
nand U45361 (N_45361,N_43668,N_43800);
nor U45362 (N_45362,N_42956,N_43553);
xor U45363 (N_45363,N_42079,N_43837);
nor U45364 (N_45364,N_43074,N_42581);
nand U45365 (N_45365,N_43078,N_42608);
or U45366 (N_45366,N_42108,N_43432);
nor U45367 (N_45367,N_42274,N_42126);
and U45368 (N_45368,N_42679,N_42200);
nand U45369 (N_45369,N_42902,N_43062);
nand U45370 (N_45370,N_42332,N_42796);
and U45371 (N_45371,N_42118,N_42958);
nand U45372 (N_45372,N_42419,N_42581);
nand U45373 (N_45373,N_43491,N_42142);
xor U45374 (N_45374,N_42755,N_42115);
xnor U45375 (N_45375,N_42263,N_43549);
or U45376 (N_45376,N_42746,N_43154);
nor U45377 (N_45377,N_42628,N_43706);
nor U45378 (N_45378,N_42175,N_42239);
nand U45379 (N_45379,N_42283,N_42787);
nand U45380 (N_45380,N_43766,N_42209);
and U45381 (N_45381,N_42823,N_43715);
or U45382 (N_45382,N_42315,N_42175);
or U45383 (N_45383,N_43344,N_43392);
and U45384 (N_45384,N_43748,N_43077);
nor U45385 (N_45385,N_43771,N_43677);
and U45386 (N_45386,N_42426,N_42707);
nor U45387 (N_45387,N_43354,N_42844);
xnor U45388 (N_45388,N_42687,N_43575);
xnor U45389 (N_45389,N_42078,N_42510);
nor U45390 (N_45390,N_42240,N_43567);
and U45391 (N_45391,N_43005,N_42225);
or U45392 (N_45392,N_42674,N_42503);
nor U45393 (N_45393,N_43387,N_43763);
or U45394 (N_45394,N_43168,N_43238);
or U45395 (N_45395,N_43020,N_43703);
and U45396 (N_45396,N_43641,N_43650);
nand U45397 (N_45397,N_42570,N_42366);
or U45398 (N_45398,N_42267,N_42937);
nor U45399 (N_45399,N_42228,N_42405);
nor U45400 (N_45400,N_42465,N_42130);
nor U45401 (N_45401,N_43311,N_42497);
xor U45402 (N_45402,N_42162,N_42371);
or U45403 (N_45403,N_43244,N_42372);
or U45404 (N_45404,N_42831,N_42461);
nor U45405 (N_45405,N_43594,N_42478);
and U45406 (N_45406,N_42431,N_42116);
nor U45407 (N_45407,N_42956,N_43097);
nand U45408 (N_45408,N_42592,N_43084);
nor U45409 (N_45409,N_43727,N_43005);
and U45410 (N_45410,N_43162,N_43524);
nand U45411 (N_45411,N_42009,N_43773);
nor U45412 (N_45412,N_43161,N_43208);
xnor U45413 (N_45413,N_42435,N_43115);
xnor U45414 (N_45414,N_42553,N_42173);
and U45415 (N_45415,N_42704,N_43526);
xnor U45416 (N_45416,N_42506,N_43033);
nor U45417 (N_45417,N_43240,N_42236);
or U45418 (N_45418,N_42455,N_43537);
and U45419 (N_45419,N_43057,N_43820);
nand U45420 (N_45420,N_43887,N_42433);
and U45421 (N_45421,N_42205,N_43339);
or U45422 (N_45422,N_43035,N_42302);
and U45423 (N_45423,N_43829,N_43884);
nand U45424 (N_45424,N_42260,N_43773);
nand U45425 (N_45425,N_43236,N_43062);
xnor U45426 (N_45426,N_43983,N_42927);
nor U45427 (N_45427,N_43876,N_42447);
nand U45428 (N_45428,N_42288,N_42001);
nand U45429 (N_45429,N_43659,N_42517);
nor U45430 (N_45430,N_43788,N_43125);
nand U45431 (N_45431,N_43611,N_42346);
or U45432 (N_45432,N_42597,N_42441);
and U45433 (N_45433,N_42747,N_42097);
and U45434 (N_45434,N_42509,N_42982);
xnor U45435 (N_45435,N_42493,N_42895);
nand U45436 (N_45436,N_43300,N_43057);
nand U45437 (N_45437,N_43064,N_43923);
nand U45438 (N_45438,N_42883,N_43692);
or U45439 (N_45439,N_43342,N_42804);
nand U45440 (N_45440,N_42348,N_42954);
xnor U45441 (N_45441,N_43030,N_42396);
or U45442 (N_45442,N_43291,N_43843);
and U45443 (N_45443,N_43453,N_42464);
and U45444 (N_45444,N_42308,N_42927);
or U45445 (N_45445,N_42464,N_43938);
nand U45446 (N_45446,N_43737,N_43871);
and U45447 (N_45447,N_42688,N_43999);
and U45448 (N_45448,N_43255,N_42308);
xor U45449 (N_45449,N_43481,N_43010);
nor U45450 (N_45450,N_42313,N_42599);
and U45451 (N_45451,N_43128,N_42194);
and U45452 (N_45452,N_43522,N_42793);
or U45453 (N_45453,N_43860,N_43837);
nand U45454 (N_45454,N_42410,N_43584);
nand U45455 (N_45455,N_43320,N_43594);
and U45456 (N_45456,N_43608,N_42750);
or U45457 (N_45457,N_42712,N_43959);
or U45458 (N_45458,N_42076,N_42607);
xnor U45459 (N_45459,N_43171,N_42484);
and U45460 (N_45460,N_43037,N_42810);
nand U45461 (N_45461,N_42154,N_42537);
nor U45462 (N_45462,N_43919,N_43378);
or U45463 (N_45463,N_43364,N_42425);
nand U45464 (N_45464,N_42999,N_43424);
and U45465 (N_45465,N_43949,N_43127);
xnor U45466 (N_45466,N_43257,N_43344);
and U45467 (N_45467,N_42256,N_42556);
nand U45468 (N_45468,N_42727,N_43378);
xnor U45469 (N_45469,N_43741,N_43117);
or U45470 (N_45470,N_43262,N_42556);
nand U45471 (N_45471,N_42315,N_42089);
and U45472 (N_45472,N_43073,N_42163);
or U45473 (N_45473,N_43962,N_43515);
nand U45474 (N_45474,N_42433,N_43229);
or U45475 (N_45475,N_42769,N_43384);
and U45476 (N_45476,N_43750,N_42234);
and U45477 (N_45477,N_42095,N_42979);
and U45478 (N_45478,N_42967,N_43797);
xnor U45479 (N_45479,N_43873,N_42816);
nor U45480 (N_45480,N_43684,N_42767);
or U45481 (N_45481,N_43049,N_42085);
nor U45482 (N_45482,N_42569,N_43987);
nor U45483 (N_45483,N_43595,N_43313);
nand U45484 (N_45484,N_42416,N_42527);
or U45485 (N_45485,N_42060,N_43981);
or U45486 (N_45486,N_42825,N_43173);
and U45487 (N_45487,N_42441,N_42176);
and U45488 (N_45488,N_43837,N_42746);
nand U45489 (N_45489,N_42936,N_43589);
nor U45490 (N_45490,N_42108,N_43709);
and U45491 (N_45491,N_43213,N_42442);
nor U45492 (N_45492,N_42613,N_43966);
nand U45493 (N_45493,N_43476,N_43848);
nor U45494 (N_45494,N_42218,N_43888);
nor U45495 (N_45495,N_42724,N_42415);
or U45496 (N_45496,N_43324,N_42469);
nand U45497 (N_45497,N_42051,N_42990);
xnor U45498 (N_45498,N_42333,N_42759);
nor U45499 (N_45499,N_43980,N_43248);
xor U45500 (N_45500,N_42908,N_42445);
nand U45501 (N_45501,N_42995,N_42403);
and U45502 (N_45502,N_42116,N_42421);
nand U45503 (N_45503,N_42714,N_42234);
and U45504 (N_45504,N_43300,N_43315);
or U45505 (N_45505,N_42635,N_43472);
nand U45506 (N_45506,N_43823,N_43085);
nor U45507 (N_45507,N_43469,N_43709);
nor U45508 (N_45508,N_42563,N_43868);
nand U45509 (N_45509,N_43897,N_43353);
xnor U45510 (N_45510,N_42278,N_43071);
nand U45511 (N_45511,N_42334,N_42987);
nor U45512 (N_45512,N_43529,N_43235);
nand U45513 (N_45513,N_42506,N_42717);
and U45514 (N_45514,N_42872,N_43679);
xnor U45515 (N_45515,N_42158,N_43260);
nor U45516 (N_45516,N_42222,N_43536);
nand U45517 (N_45517,N_42372,N_42221);
or U45518 (N_45518,N_43452,N_42131);
and U45519 (N_45519,N_43042,N_43160);
and U45520 (N_45520,N_42442,N_43971);
xnor U45521 (N_45521,N_42153,N_42421);
nor U45522 (N_45522,N_43204,N_43035);
nand U45523 (N_45523,N_43027,N_42595);
or U45524 (N_45524,N_42289,N_43190);
nor U45525 (N_45525,N_43432,N_43251);
nor U45526 (N_45526,N_42020,N_42243);
and U45527 (N_45527,N_42481,N_42234);
nand U45528 (N_45528,N_43245,N_42164);
or U45529 (N_45529,N_43286,N_42719);
or U45530 (N_45530,N_42075,N_42445);
or U45531 (N_45531,N_42813,N_43431);
nand U45532 (N_45532,N_43314,N_42681);
nand U45533 (N_45533,N_42581,N_43412);
or U45534 (N_45534,N_43039,N_43313);
nor U45535 (N_45535,N_43068,N_43056);
and U45536 (N_45536,N_42936,N_43569);
and U45537 (N_45537,N_43615,N_42758);
nor U45538 (N_45538,N_43540,N_42535);
and U45539 (N_45539,N_42082,N_43065);
and U45540 (N_45540,N_43271,N_43109);
xnor U45541 (N_45541,N_42701,N_43977);
xor U45542 (N_45542,N_42141,N_43940);
nor U45543 (N_45543,N_42792,N_43433);
xor U45544 (N_45544,N_43582,N_42547);
or U45545 (N_45545,N_42631,N_42936);
nor U45546 (N_45546,N_42062,N_42612);
or U45547 (N_45547,N_42692,N_42257);
nand U45548 (N_45548,N_43001,N_42613);
and U45549 (N_45549,N_43382,N_43789);
nor U45550 (N_45550,N_43773,N_42179);
or U45551 (N_45551,N_43301,N_43663);
and U45552 (N_45552,N_42345,N_42995);
nand U45553 (N_45553,N_42518,N_43300);
xnor U45554 (N_45554,N_42246,N_43221);
nor U45555 (N_45555,N_43730,N_43925);
and U45556 (N_45556,N_42950,N_42349);
xnor U45557 (N_45557,N_43707,N_42381);
or U45558 (N_45558,N_42953,N_42132);
nand U45559 (N_45559,N_43503,N_43659);
nor U45560 (N_45560,N_42488,N_42674);
or U45561 (N_45561,N_42200,N_43115);
and U45562 (N_45562,N_42504,N_42354);
nor U45563 (N_45563,N_43620,N_43425);
nor U45564 (N_45564,N_42183,N_43308);
nor U45565 (N_45565,N_43372,N_43378);
nand U45566 (N_45566,N_43516,N_43157);
nor U45567 (N_45567,N_42001,N_43080);
or U45568 (N_45568,N_42481,N_42389);
xor U45569 (N_45569,N_43906,N_43824);
nor U45570 (N_45570,N_42433,N_42396);
nor U45571 (N_45571,N_43741,N_42416);
and U45572 (N_45572,N_42763,N_43555);
xor U45573 (N_45573,N_42622,N_43886);
nand U45574 (N_45574,N_43364,N_42671);
and U45575 (N_45575,N_42811,N_42006);
nand U45576 (N_45576,N_42650,N_43460);
nor U45577 (N_45577,N_43863,N_42111);
or U45578 (N_45578,N_43619,N_42189);
and U45579 (N_45579,N_42334,N_43164);
xnor U45580 (N_45580,N_42857,N_42292);
nand U45581 (N_45581,N_43250,N_43552);
nand U45582 (N_45582,N_43256,N_42236);
nor U45583 (N_45583,N_43970,N_42824);
xnor U45584 (N_45584,N_43323,N_43153);
xnor U45585 (N_45585,N_43797,N_43236);
nor U45586 (N_45586,N_42970,N_42371);
and U45587 (N_45587,N_43503,N_42891);
nor U45588 (N_45588,N_43031,N_43211);
xnor U45589 (N_45589,N_42227,N_43791);
and U45590 (N_45590,N_43162,N_43656);
and U45591 (N_45591,N_43351,N_42688);
and U45592 (N_45592,N_42604,N_43467);
nor U45593 (N_45593,N_42527,N_42583);
nor U45594 (N_45594,N_42702,N_42737);
xnor U45595 (N_45595,N_42652,N_43179);
xor U45596 (N_45596,N_43247,N_43709);
nor U45597 (N_45597,N_42935,N_43984);
nand U45598 (N_45598,N_42869,N_42199);
or U45599 (N_45599,N_42404,N_43539);
and U45600 (N_45600,N_42589,N_42945);
nand U45601 (N_45601,N_42908,N_42491);
nand U45602 (N_45602,N_42765,N_42672);
xor U45603 (N_45603,N_43616,N_43896);
nor U45604 (N_45604,N_42508,N_43013);
nor U45605 (N_45605,N_43349,N_43934);
or U45606 (N_45606,N_42550,N_43672);
nor U45607 (N_45607,N_42598,N_42169);
nand U45608 (N_45608,N_43518,N_43719);
and U45609 (N_45609,N_43853,N_43413);
nor U45610 (N_45610,N_43159,N_42570);
or U45611 (N_45611,N_42823,N_42114);
nor U45612 (N_45612,N_43480,N_43951);
and U45613 (N_45613,N_43299,N_43051);
and U45614 (N_45614,N_42144,N_42961);
nor U45615 (N_45615,N_42695,N_43938);
nor U45616 (N_45616,N_42274,N_42456);
and U45617 (N_45617,N_42841,N_42056);
and U45618 (N_45618,N_43563,N_42172);
and U45619 (N_45619,N_43885,N_43937);
or U45620 (N_45620,N_42976,N_43139);
nand U45621 (N_45621,N_42240,N_43808);
xor U45622 (N_45622,N_43338,N_42501);
xor U45623 (N_45623,N_42853,N_42558);
and U45624 (N_45624,N_43316,N_43180);
and U45625 (N_45625,N_43800,N_42822);
and U45626 (N_45626,N_43707,N_43586);
nor U45627 (N_45627,N_43061,N_43956);
and U45628 (N_45628,N_43808,N_43686);
and U45629 (N_45629,N_42608,N_42078);
and U45630 (N_45630,N_43232,N_43104);
nor U45631 (N_45631,N_42230,N_43512);
xnor U45632 (N_45632,N_43922,N_42149);
nor U45633 (N_45633,N_42679,N_42238);
and U45634 (N_45634,N_43271,N_43325);
nor U45635 (N_45635,N_42623,N_42047);
nand U45636 (N_45636,N_43709,N_43968);
nand U45637 (N_45637,N_42001,N_43573);
and U45638 (N_45638,N_43007,N_42313);
nand U45639 (N_45639,N_42049,N_43774);
or U45640 (N_45640,N_43783,N_42320);
nor U45641 (N_45641,N_42031,N_42991);
and U45642 (N_45642,N_43333,N_43491);
xnor U45643 (N_45643,N_43943,N_43881);
or U45644 (N_45644,N_43542,N_43056);
xor U45645 (N_45645,N_42761,N_42621);
or U45646 (N_45646,N_43113,N_42232);
xor U45647 (N_45647,N_43205,N_43073);
or U45648 (N_45648,N_42605,N_42655);
nand U45649 (N_45649,N_43101,N_43233);
or U45650 (N_45650,N_42917,N_42394);
nand U45651 (N_45651,N_43018,N_42814);
or U45652 (N_45652,N_43975,N_42522);
xnor U45653 (N_45653,N_43223,N_43315);
xnor U45654 (N_45654,N_42610,N_42607);
nand U45655 (N_45655,N_43899,N_43801);
and U45656 (N_45656,N_43232,N_42618);
nand U45657 (N_45657,N_42955,N_42501);
nand U45658 (N_45658,N_42988,N_42056);
xor U45659 (N_45659,N_42883,N_42469);
nand U45660 (N_45660,N_43450,N_43666);
or U45661 (N_45661,N_43151,N_42653);
and U45662 (N_45662,N_42545,N_43289);
nor U45663 (N_45663,N_42145,N_42547);
nand U45664 (N_45664,N_42897,N_42297);
nand U45665 (N_45665,N_42661,N_42698);
nand U45666 (N_45666,N_42253,N_43293);
or U45667 (N_45667,N_43476,N_43091);
and U45668 (N_45668,N_42825,N_43126);
nand U45669 (N_45669,N_42157,N_42108);
xnor U45670 (N_45670,N_43073,N_43146);
and U45671 (N_45671,N_43755,N_42591);
or U45672 (N_45672,N_43904,N_42931);
or U45673 (N_45673,N_43231,N_42953);
nand U45674 (N_45674,N_43506,N_43372);
xnor U45675 (N_45675,N_43159,N_43204);
xnor U45676 (N_45676,N_43626,N_42258);
and U45677 (N_45677,N_43823,N_42487);
nor U45678 (N_45678,N_42042,N_42776);
or U45679 (N_45679,N_42212,N_42833);
and U45680 (N_45680,N_43344,N_42500);
nand U45681 (N_45681,N_42042,N_42546);
nand U45682 (N_45682,N_42116,N_43451);
nor U45683 (N_45683,N_43032,N_42291);
nand U45684 (N_45684,N_43737,N_43307);
nor U45685 (N_45685,N_43967,N_42712);
or U45686 (N_45686,N_43335,N_43432);
nand U45687 (N_45687,N_43701,N_42894);
nand U45688 (N_45688,N_43905,N_42025);
nand U45689 (N_45689,N_43463,N_42574);
and U45690 (N_45690,N_42051,N_43108);
or U45691 (N_45691,N_43231,N_42252);
or U45692 (N_45692,N_42559,N_43072);
or U45693 (N_45693,N_42808,N_42401);
nand U45694 (N_45694,N_43200,N_42310);
nand U45695 (N_45695,N_42522,N_42037);
nor U45696 (N_45696,N_43957,N_42322);
and U45697 (N_45697,N_42432,N_43210);
xnor U45698 (N_45698,N_42633,N_42743);
nor U45699 (N_45699,N_43979,N_43350);
or U45700 (N_45700,N_43911,N_42073);
or U45701 (N_45701,N_42726,N_43155);
or U45702 (N_45702,N_43905,N_42751);
nand U45703 (N_45703,N_43738,N_42766);
and U45704 (N_45704,N_42881,N_42649);
or U45705 (N_45705,N_42665,N_42926);
and U45706 (N_45706,N_42346,N_43964);
nor U45707 (N_45707,N_42772,N_42296);
xnor U45708 (N_45708,N_42978,N_42927);
nor U45709 (N_45709,N_42908,N_42375);
and U45710 (N_45710,N_43693,N_42501);
xor U45711 (N_45711,N_43233,N_43493);
xor U45712 (N_45712,N_42386,N_43964);
nand U45713 (N_45713,N_43223,N_43642);
xor U45714 (N_45714,N_43926,N_43464);
nor U45715 (N_45715,N_42984,N_43332);
nor U45716 (N_45716,N_43199,N_43428);
nor U45717 (N_45717,N_42820,N_43767);
or U45718 (N_45718,N_43696,N_43971);
or U45719 (N_45719,N_43271,N_43119);
and U45720 (N_45720,N_42097,N_43435);
nor U45721 (N_45721,N_43592,N_43654);
nor U45722 (N_45722,N_43608,N_43643);
nor U45723 (N_45723,N_42844,N_43638);
xor U45724 (N_45724,N_43902,N_42132);
or U45725 (N_45725,N_43383,N_42127);
or U45726 (N_45726,N_43619,N_43896);
xnor U45727 (N_45727,N_42688,N_43334);
xor U45728 (N_45728,N_43316,N_43916);
and U45729 (N_45729,N_43384,N_42211);
nor U45730 (N_45730,N_42653,N_43482);
nor U45731 (N_45731,N_42694,N_42680);
and U45732 (N_45732,N_42074,N_42574);
or U45733 (N_45733,N_43333,N_42595);
xnor U45734 (N_45734,N_43108,N_42250);
and U45735 (N_45735,N_43988,N_42877);
and U45736 (N_45736,N_43036,N_43460);
or U45737 (N_45737,N_42106,N_43048);
xnor U45738 (N_45738,N_42045,N_42665);
nor U45739 (N_45739,N_43480,N_43943);
or U45740 (N_45740,N_43925,N_43410);
nand U45741 (N_45741,N_42870,N_42828);
and U45742 (N_45742,N_43353,N_43676);
or U45743 (N_45743,N_42252,N_42040);
nor U45744 (N_45744,N_43319,N_43280);
nor U45745 (N_45745,N_43942,N_43292);
and U45746 (N_45746,N_42967,N_42612);
and U45747 (N_45747,N_43483,N_42128);
nor U45748 (N_45748,N_42269,N_42005);
nor U45749 (N_45749,N_42396,N_43275);
or U45750 (N_45750,N_42321,N_42689);
nor U45751 (N_45751,N_42752,N_42178);
or U45752 (N_45752,N_42250,N_42192);
nand U45753 (N_45753,N_43360,N_42413);
or U45754 (N_45754,N_43863,N_42939);
or U45755 (N_45755,N_43906,N_43303);
xnor U45756 (N_45756,N_43638,N_42251);
or U45757 (N_45757,N_43078,N_42341);
nor U45758 (N_45758,N_43464,N_42874);
xnor U45759 (N_45759,N_43236,N_43667);
or U45760 (N_45760,N_42185,N_42909);
xnor U45761 (N_45761,N_42984,N_43698);
and U45762 (N_45762,N_43402,N_43976);
or U45763 (N_45763,N_43731,N_43494);
xor U45764 (N_45764,N_42140,N_42869);
xor U45765 (N_45765,N_43157,N_42888);
or U45766 (N_45766,N_43699,N_42349);
nand U45767 (N_45767,N_43416,N_42112);
nor U45768 (N_45768,N_43715,N_43438);
and U45769 (N_45769,N_42918,N_43228);
nor U45770 (N_45770,N_43330,N_42859);
nand U45771 (N_45771,N_42251,N_43778);
or U45772 (N_45772,N_42386,N_43603);
nand U45773 (N_45773,N_43617,N_42116);
nand U45774 (N_45774,N_43803,N_43025);
xor U45775 (N_45775,N_43496,N_43968);
nor U45776 (N_45776,N_42824,N_43352);
nand U45777 (N_45777,N_42951,N_42079);
nor U45778 (N_45778,N_42086,N_43609);
and U45779 (N_45779,N_42319,N_42789);
or U45780 (N_45780,N_42115,N_42979);
or U45781 (N_45781,N_43420,N_43225);
nor U45782 (N_45782,N_42143,N_42946);
or U45783 (N_45783,N_42618,N_42347);
xnor U45784 (N_45784,N_43213,N_42362);
or U45785 (N_45785,N_42112,N_43630);
or U45786 (N_45786,N_43979,N_42237);
nor U45787 (N_45787,N_43479,N_42730);
or U45788 (N_45788,N_42446,N_42519);
or U45789 (N_45789,N_43734,N_42142);
and U45790 (N_45790,N_43971,N_43847);
nor U45791 (N_45791,N_42952,N_42694);
or U45792 (N_45792,N_42012,N_43486);
xor U45793 (N_45793,N_43206,N_42676);
or U45794 (N_45794,N_42386,N_43572);
xnor U45795 (N_45795,N_43866,N_43878);
and U45796 (N_45796,N_43336,N_42285);
nor U45797 (N_45797,N_43716,N_43264);
and U45798 (N_45798,N_43259,N_42737);
xor U45799 (N_45799,N_43430,N_42044);
nor U45800 (N_45800,N_43749,N_43174);
and U45801 (N_45801,N_42083,N_42150);
or U45802 (N_45802,N_42483,N_42847);
nand U45803 (N_45803,N_43265,N_43116);
xnor U45804 (N_45804,N_43158,N_43295);
xnor U45805 (N_45805,N_43610,N_43922);
nor U45806 (N_45806,N_43149,N_43484);
nor U45807 (N_45807,N_43603,N_42339);
or U45808 (N_45808,N_42645,N_42945);
xor U45809 (N_45809,N_42029,N_42668);
and U45810 (N_45810,N_43883,N_42595);
xor U45811 (N_45811,N_43302,N_43326);
xor U45812 (N_45812,N_43063,N_42749);
xor U45813 (N_45813,N_43369,N_43734);
nand U45814 (N_45814,N_43643,N_42588);
xor U45815 (N_45815,N_43742,N_42746);
nor U45816 (N_45816,N_42569,N_43287);
xor U45817 (N_45817,N_42587,N_42502);
xnor U45818 (N_45818,N_42314,N_42833);
nand U45819 (N_45819,N_43740,N_43729);
nor U45820 (N_45820,N_43653,N_43294);
nor U45821 (N_45821,N_43133,N_42130);
xor U45822 (N_45822,N_42476,N_42972);
nor U45823 (N_45823,N_42840,N_43660);
nand U45824 (N_45824,N_42305,N_43729);
xnor U45825 (N_45825,N_42585,N_43682);
or U45826 (N_45826,N_43171,N_43243);
or U45827 (N_45827,N_42973,N_43461);
and U45828 (N_45828,N_42786,N_43256);
or U45829 (N_45829,N_43792,N_43019);
and U45830 (N_45830,N_43323,N_42813);
and U45831 (N_45831,N_43418,N_42862);
nor U45832 (N_45832,N_43293,N_43991);
nor U45833 (N_45833,N_43052,N_42699);
xor U45834 (N_45834,N_42832,N_42768);
or U45835 (N_45835,N_43599,N_42647);
and U45836 (N_45836,N_42283,N_43742);
nand U45837 (N_45837,N_43442,N_42395);
or U45838 (N_45838,N_42179,N_42127);
or U45839 (N_45839,N_43366,N_43800);
xnor U45840 (N_45840,N_43189,N_42727);
nand U45841 (N_45841,N_42187,N_42788);
xnor U45842 (N_45842,N_42696,N_43214);
xor U45843 (N_45843,N_42284,N_43901);
nand U45844 (N_45844,N_43722,N_42036);
xnor U45845 (N_45845,N_42360,N_43702);
and U45846 (N_45846,N_43103,N_42800);
xnor U45847 (N_45847,N_42321,N_43866);
xor U45848 (N_45848,N_42783,N_42917);
and U45849 (N_45849,N_43575,N_42529);
nand U45850 (N_45850,N_43280,N_43166);
or U45851 (N_45851,N_42216,N_43641);
nor U45852 (N_45852,N_43600,N_43603);
nor U45853 (N_45853,N_42096,N_42045);
nand U45854 (N_45854,N_42013,N_42193);
nand U45855 (N_45855,N_43433,N_42541);
or U45856 (N_45856,N_42254,N_42043);
or U45857 (N_45857,N_43837,N_43763);
or U45858 (N_45858,N_43242,N_42561);
or U45859 (N_45859,N_42032,N_43642);
nor U45860 (N_45860,N_42401,N_42205);
nor U45861 (N_45861,N_42747,N_42384);
or U45862 (N_45862,N_43506,N_42549);
and U45863 (N_45863,N_43305,N_43119);
xnor U45864 (N_45864,N_43578,N_42441);
nor U45865 (N_45865,N_43128,N_43467);
nor U45866 (N_45866,N_42583,N_43600);
nand U45867 (N_45867,N_43318,N_42881);
xor U45868 (N_45868,N_43382,N_42449);
and U45869 (N_45869,N_43729,N_42048);
nor U45870 (N_45870,N_43866,N_43507);
and U45871 (N_45871,N_43143,N_43168);
or U45872 (N_45872,N_42716,N_43731);
or U45873 (N_45873,N_43642,N_43491);
or U45874 (N_45874,N_43889,N_42634);
nor U45875 (N_45875,N_43297,N_42852);
nor U45876 (N_45876,N_42550,N_43581);
nor U45877 (N_45877,N_42312,N_42961);
and U45878 (N_45878,N_42227,N_43793);
nand U45879 (N_45879,N_43964,N_43441);
and U45880 (N_45880,N_43686,N_42328);
or U45881 (N_45881,N_42780,N_42012);
or U45882 (N_45882,N_42127,N_43564);
xor U45883 (N_45883,N_42146,N_42715);
or U45884 (N_45884,N_42615,N_43227);
xnor U45885 (N_45885,N_43294,N_43782);
and U45886 (N_45886,N_42110,N_42802);
xor U45887 (N_45887,N_43198,N_43782);
nor U45888 (N_45888,N_42112,N_42035);
and U45889 (N_45889,N_42475,N_43913);
or U45890 (N_45890,N_42801,N_42551);
nor U45891 (N_45891,N_42100,N_42530);
or U45892 (N_45892,N_43189,N_43762);
nor U45893 (N_45893,N_42435,N_43326);
xnor U45894 (N_45894,N_43819,N_42453);
nor U45895 (N_45895,N_42739,N_43039);
xnor U45896 (N_45896,N_42903,N_43395);
nor U45897 (N_45897,N_42526,N_42589);
and U45898 (N_45898,N_42006,N_43502);
and U45899 (N_45899,N_42789,N_43508);
or U45900 (N_45900,N_43676,N_42521);
nor U45901 (N_45901,N_42030,N_43035);
and U45902 (N_45902,N_43184,N_42135);
or U45903 (N_45903,N_42445,N_43208);
or U45904 (N_45904,N_42626,N_43947);
nor U45905 (N_45905,N_42345,N_42543);
nor U45906 (N_45906,N_42883,N_42530);
xor U45907 (N_45907,N_42360,N_42794);
or U45908 (N_45908,N_43308,N_43420);
and U45909 (N_45909,N_42947,N_42427);
nand U45910 (N_45910,N_42923,N_42831);
xor U45911 (N_45911,N_42665,N_42166);
or U45912 (N_45912,N_43740,N_42554);
xor U45913 (N_45913,N_42660,N_42559);
nor U45914 (N_45914,N_43577,N_42933);
nand U45915 (N_45915,N_43136,N_42102);
nand U45916 (N_45916,N_43730,N_43351);
and U45917 (N_45917,N_43689,N_42640);
and U45918 (N_45918,N_42697,N_43550);
or U45919 (N_45919,N_42103,N_43002);
or U45920 (N_45920,N_43555,N_43091);
nand U45921 (N_45921,N_42451,N_43711);
or U45922 (N_45922,N_42952,N_42321);
nor U45923 (N_45923,N_43887,N_42638);
or U45924 (N_45924,N_43833,N_43974);
or U45925 (N_45925,N_42587,N_42695);
and U45926 (N_45926,N_42401,N_43287);
and U45927 (N_45927,N_42417,N_42573);
and U45928 (N_45928,N_42718,N_43974);
and U45929 (N_45929,N_42082,N_42979);
nor U45930 (N_45930,N_43201,N_43937);
nor U45931 (N_45931,N_42759,N_43794);
and U45932 (N_45932,N_43402,N_42981);
xor U45933 (N_45933,N_43113,N_42929);
or U45934 (N_45934,N_43806,N_42781);
and U45935 (N_45935,N_42316,N_43753);
xnor U45936 (N_45936,N_42979,N_43354);
xor U45937 (N_45937,N_42863,N_43397);
nand U45938 (N_45938,N_42954,N_43412);
xnor U45939 (N_45939,N_42467,N_42255);
nand U45940 (N_45940,N_42086,N_42376);
nor U45941 (N_45941,N_43642,N_43379);
nand U45942 (N_45942,N_42007,N_43829);
or U45943 (N_45943,N_42405,N_43317);
nor U45944 (N_45944,N_42894,N_43457);
nand U45945 (N_45945,N_42393,N_43419);
and U45946 (N_45946,N_42891,N_42157);
xnor U45947 (N_45947,N_42870,N_42703);
nor U45948 (N_45948,N_43544,N_42376);
nor U45949 (N_45949,N_43541,N_43391);
nor U45950 (N_45950,N_43127,N_43139);
nand U45951 (N_45951,N_42314,N_42074);
nand U45952 (N_45952,N_42168,N_42709);
and U45953 (N_45953,N_42183,N_42160);
or U45954 (N_45954,N_43060,N_42263);
and U45955 (N_45955,N_43259,N_43207);
xor U45956 (N_45956,N_43679,N_43646);
or U45957 (N_45957,N_42300,N_43361);
and U45958 (N_45958,N_43472,N_43483);
nand U45959 (N_45959,N_43113,N_42768);
nor U45960 (N_45960,N_43724,N_43555);
xnor U45961 (N_45961,N_43243,N_42446);
and U45962 (N_45962,N_43720,N_42309);
and U45963 (N_45963,N_42619,N_42421);
nand U45964 (N_45964,N_42076,N_42235);
nand U45965 (N_45965,N_43916,N_43717);
or U45966 (N_45966,N_42337,N_42462);
xor U45967 (N_45967,N_43179,N_42624);
or U45968 (N_45968,N_42831,N_42393);
and U45969 (N_45969,N_43434,N_42984);
and U45970 (N_45970,N_43730,N_43930);
or U45971 (N_45971,N_42867,N_43163);
or U45972 (N_45972,N_43709,N_42818);
and U45973 (N_45973,N_43521,N_42018);
or U45974 (N_45974,N_42957,N_42288);
nand U45975 (N_45975,N_43144,N_43770);
xor U45976 (N_45976,N_42600,N_43984);
xor U45977 (N_45977,N_42568,N_42477);
xor U45978 (N_45978,N_43361,N_43654);
and U45979 (N_45979,N_42737,N_43127);
nand U45980 (N_45980,N_43879,N_43078);
and U45981 (N_45981,N_42128,N_43466);
xnor U45982 (N_45982,N_42518,N_43522);
nand U45983 (N_45983,N_43411,N_42650);
nand U45984 (N_45984,N_42684,N_42756);
or U45985 (N_45985,N_42570,N_43580);
and U45986 (N_45986,N_42759,N_42613);
or U45987 (N_45987,N_43708,N_42908);
or U45988 (N_45988,N_43581,N_43015);
xnor U45989 (N_45989,N_42455,N_43283);
or U45990 (N_45990,N_42676,N_43287);
nand U45991 (N_45991,N_42236,N_43215);
or U45992 (N_45992,N_42513,N_43311);
and U45993 (N_45993,N_42866,N_43192);
or U45994 (N_45994,N_42139,N_42703);
nor U45995 (N_45995,N_43134,N_43948);
or U45996 (N_45996,N_43199,N_42222);
nand U45997 (N_45997,N_42308,N_43905);
xnor U45998 (N_45998,N_43735,N_43268);
and U45999 (N_45999,N_42426,N_43043);
or U46000 (N_46000,N_44229,N_45402);
and U46001 (N_46001,N_44130,N_44627);
nor U46002 (N_46002,N_45542,N_45761);
nand U46003 (N_46003,N_44828,N_45458);
nand U46004 (N_46004,N_44315,N_44392);
nor U46005 (N_46005,N_45438,N_44393);
nand U46006 (N_46006,N_44641,N_44072);
nor U46007 (N_46007,N_45798,N_45487);
or U46008 (N_46008,N_44712,N_45215);
nand U46009 (N_46009,N_45660,N_44269);
nand U46010 (N_46010,N_45342,N_45519);
nand U46011 (N_46011,N_44900,N_45777);
and U46012 (N_46012,N_44964,N_44423);
nor U46013 (N_46013,N_44736,N_44203);
nand U46014 (N_46014,N_44924,N_44613);
nor U46015 (N_46015,N_45966,N_44446);
and U46016 (N_46016,N_45277,N_44618);
nor U46017 (N_46017,N_44375,N_44011);
nand U46018 (N_46018,N_44010,N_44471);
or U46019 (N_46019,N_44501,N_44510);
and U46020 (N_46020,N_45117,N_45228);
or U46021 (N_46021,N_44268,N_45085);
xor U46022 (N_46022,N_45591,N_44147);
xnor U46023 (N_46023,N_44711,N_45401);
and U46024 (N_46024,N_44397,N_44673);
xnor U46025 (N_46025,N_45294,N_45807);
xnor U46026 (N_46026,N_44063,N_45831);
or U46027 (N_46027,N_44132,N_45996);
xnor U46028 (N_46028,N_45185,N_44639);
xnor U46029 (N_46029,N_45230,N_44430);
xnor U46030 (N_46030,N_45167,N_44133);
nand U46031 (N_46031,N_45558,N_45281);
or U46032 (N_46032,N_45297,N_45544);
nand U46033 (N_46033,N_45221,N_45472);
and U46034 (N_46034,N_45408,N_45992);
nor U46035 (N_46035,N_44722,N_44880);
nand U46036 (N_46036,N_44438,N_45262);
and U46037 (N_46037,N_45148,N_44633);
nand U46038 (N_46038,N_45843,N_44756);
xnor U46039 (N_46039,N_45583,N_44976);
nor U46040 (N_46040,N_45555,N_45766);
or U46041 (N_46041,N_45114,N_44889);
or U46042 (N_46042,N_44272,N_45033);
and U46043 (N_46043,N_45416,N_44293);
xor U46044 (N_46044,N_45720,N_44239);
nand U46045 (N_46045,N_45822,N_44770);
and U46046 (N_46046,N_45028,N_44359);
and U46047 (N_46047,N_45653,N_45156);
nor U46048 (N_46048,N_44300,N_45675);
nor U46049 (N_46049,N_45980,N_44585);
nand U46050 (N_46050,N_45677,N_45504);
or U46051 (N_46051,N_44674,N_45526);
nor U46052 (N_46052,N_44812,N_45573);
xor U46053 (N_46053,N_45227,N_45122);
xor U46054 (N_46054,N_44034,N_44526);
xor U46055 (N_46055,N_45743,N_44102);
nand U46056 (N_46056,N_45674,N_45726);
and U46057 (N_46057,N_44313,N_44329);
nand U46058 (N_46058,N_45550,N_44140);
and U46059 (N_46059,N_44979,N_44197);
nand U46060 (N_46060,N_44436,N_44823);
and U46061 (N_46061,N_45810,N_44824);
nand U46062 (N_46062,N_45833,N_45999);
or U46063 (N_46063,N_44541,N_44009);
nor U46064 (N_46064,N_45234,N_45264);
and U46065 (N_46065,N_44449,N_44251);
and U46066 (N_46066,N_45902,N_45232);
nand U46067 (N_46067,N_44017,N_45723);
nor U46068 (N_46068,N_44018,N_44084);
or U46069 (N_46069,N_44958,N_44307);
or U46070 (N_46070,N_45708,N_45521);
or U46071 (N_46071,N_44914,N_45590);
nand U46072 (N_46072,N_44169,N_45935);
xor U46073 (N_46073,N_44917,N_44925);
and U46074 (N_46074,N_45929,N_44400);
xnor U46075 (N_46075,N_45460,N_45933);
xor U46076 (N_46076,N_44894,N_45658);
nor U46077 (N_46077,N_45256,N_45151);
nor U46078 (N_46078,N_44886,N_44418);
xnor U46079 (N_46079,N_45701,N_44544);
nand U46080 (N_46080,N_45961,N_45862);
nor U46081 (N_46081,N_44245,N_45662);
xor U46082 (N_46082,N_44749,N_44699);
and U46083 (N_46083,N_45199,N_45671);
and U46084 (N_46084,N_45391,N_45161);
or U46085 (N_46085,N_44746,N_44226);
and U46086 (N_46086,N_45224,N_45038);
nor U46087 (N_46087,N_45271,N_45687);
or U46088 (N_46088,N_45017,N_45955);
and U46089 (N_46089,N_44915,N_45174);
or U46090 (N_46090,N_44762,N_44153);
nand U46091 (N_46091,N_44214,N_45871);
nand U46092 (N_46092,N_45008,N_45093);
nor U46093 (N_46093,N_44387,N_44345);
and U46094 (N_46094,N_44983,N_44957);
nand U46095 (N_46095,N_45339,N_45285);
nand U46096 (N_46096,N_45859,N_44683);
xnor U46097 (N_46097,N_44281,N_45059);
nand U46098 (N_46098,N_44076,N_44177);
nand U46099 (N_46099,N_45042,N_45388);
or U46100 (N_46100,N_44342,N_44079);
and U46101 (N_46101,N_45823,N_45900);
nor U46102 (N_46102,N_45879,N_44919);
xor U46103 (N_46103,N_44086,N_45066);
nor U46104 (N_46104,N_44678,N_44932);
and U46105 (N_46105,N_44789,N_45787);
nor U46106 (N_46106,N_44440,N_45268);
and U46107 (N_46107,N_44649,N_45856);
xor U46108 (N_46108,N_44877,N_44971);
and U46109 (N_46109,N_45877,N_44224);
or U46110 (N_46110,N_45169,N_45347);
nor U46111 (N_46111,N_44625,N_45063);
and U46112 (N_46112,N_44007,N_44171);
and U46113 (N_46113,N_45914,N_44991);
and U46114 (N_46114,N_44481,N_44259);
and U46115 (N_46115,N_45097,N_44710);
nor U46116 (N_46116,N_44173,N_44998);
or U46117 (N_46117,N_44391,N_45025);
nand U46118 (N_46118,N_45554,N_45340);
and U46119 (N_46119,N_44858,N_44614);
and U46120 (N_46120,N_45686,N_45067);
and U46121 (N_46121,N_45390,N_44439);
and U46122 (N_46122,N_45361,N_44583);
nor U46123 (N_46123,N_44396,N_45456);
or U46124 (N_46124,N_45868,N_44031);
and U46125 (N_46125,N_44250,N_44491);
nand U46126 (N_46126,N_45894,N_45680);
nor U46127 (N_46127,N_45690,N_45733);
and U46128 (N_46128,N_44708,N_45382);
xnor U46129 (N_46129,N_44427,N_45683);
and U46130 (N_46130,N_45596,N_44518);
nor U46131 (N_46131,N_44747,N_44111);
and U46132 (N_46132,N_45629,N_44097);
nor U46133 (N_46133,N_45747,N_44955);
nor U46134 (N_46134,N_44498,N_45560);
and U46135 (N_46135,N_45474,N_45600);
xnor U46136 (N_46136,N_44208,N_44800);
nor U46137 (N_46137,N_45570,N_45483);
xnor U46138 (N_46138,N_45247,N_45096);
nor U46139 (N_46139,N_45193,N_44271);
xor U46140 (N_46140,N_44118,N_44782);
or U46141 (N_46141,N_45730,N_45092);
or U46142 (N_46142,N_45449,N_44941);
or U46143 (N_46143,N_44107,N_44228);
nand U46144 (N_46144,N_44929,N_45517);
and U46145 (N_46145,N_44455,N_44277);
nand U46146 (N_46146,N_45429,N_44287);
xor U46147 (N_46147,N_45749,N_45322);
nand U46148 (N_46148,N_44165,N_45495);
nor U46149 (N_46149,N_45901,N_44787);
nand U46150 (N_46150,N_45255,N_45086);
nor U46151 (N_46151,N_44089,N_45163);
nand U46152 (N_46152,N_44116,N_45126);
or U46153 (N_46153,N_44167,N_45592);
xnor U46154 (N_46154,N_45303,N_45398);
nand U46155 (N_46155,N_44316,N_45707);
xor U46156 (N_46156,N_45187,N_45734);
xnor U46157 (N_46157,N_44205,N_45279);
and U46158 (N_46158,N_45562,N_44586);
xnor U46159 (N_46159,N_45800,N_44443);
nor U46160 (N_46160,N_44795,N_44818);
xor U46161 (N_46161,N_44637,N_45503);
xnor U46162 (N_46162,N_44942,N_44821);
or U46163 (N_46163,N_45643,N_44552);
or U46164 (N_46164,N_45657,N_45007);
or U46165 (N_46165,N_45353,N_44069);
nor U46166 (N_46166,N_45949,N_44847);
and U46167 (N_46167,N_45226,N_44211);
or U46168 (N_46168,N_45292,N_45509);
and U46169 (N_46169,N_45317,N_45426);
or U46170 (N_46170,N_44696,N_45754);
and U46171 (N_46171,N_44144,N_44270);
nand U46172 (N_46172,N_44934,N_45113);
and U46173 (N_46173,N_44148,N_44970);
nor U46174 (N_46174,N_45359,N_45225);
and U46175 (N_46175,N_44508,N_45385);
and U46176 (N_46176,N_44032,N_45891);
and U46177 (N_46177,N_45697,N_45885);
xor U46178 (N_46178,N_45988,N_44549);
or U46179 (N_46179,N_44528,N_45500);
nor U46180 (N_46180,N_45586,N_45621);
nor U46181 (N_46181,N_44283,N_45420);
nor U46182 (N_46182,N_45842,N_44968);
nor U46183 (N_46183,N_44462,N_45642);
nand U46184 (N_46184,N_45441,N_45880);
nand U46185 (N_46185,N_45186,N_45357);
xnor U46186 (N_46186,N_44406,N_45159);
xnor U46187 (N_46187,N_44965,N_45065);
nor U46188 (N_46188,N_45107,N_45947);
nand U46189 (N_46189,N_44309,N_45080);
xor U46190 (N_46190,N_45537,N_44050);
and U46191 (N_46191,N_45418,N_45133);
or U46192 (N_46192,N_44382,N_45507);
nand U46193 (N_46193,N_45329,N_45424);
nand U46194 (N_46194,N_45684,N_44906);
and U46195 (N_46195,N_45918,N_45534);
nand U46196 (N_46196,N_44398,N_45379);
nor U46197 (N_46197,N_44442,N_45470);
xnor U46198 (N_46198,N_44274,N_45541);
or U46199 (N_46199,N_45516,N_44394);
and U46200 (N_46200,N_44853,N_45981);
xor U46201 (N_46201,N_45756,N_44936);
nand U46202 (N_46202,N_45714,N_44928);
and U46203 (N_46203,N_44368,N_44253);
or U46204 (N_46204,N_44456,N_45864);
xnor U46205 (N_46205,N_44682,N_44164);
and U46206 (N_46206,N_45805,N_44183);
or U46207 (N_46207,N_44220,N_45445);
or U46208 (N_46208,N_44356,N_45791);
nor U46209 (N_46209,N_45259,N_45157);
and U46210 (N_46210,N_44833,N_44679);
nand U46211 (N_46211,N_44230,N_45404);
nand U46212 (N_46212,N_45464,N_45443);
nor U46213 (N_46213,N_44232,N_45165);
and U46214 (N_46214,N_44690,N_44026);
and U46215 (N_46215,N_44347,N_44059);
and U46216 (N_46216,N_45923,N_44502);
xor U46217 (N_46217,N_44995,N_45220);
and U46218 (N_46218,N_44516,N_44348);
or U46219 (N_46219,N_45752,N_44545);
nand U46220 (N_46220,N_44567,N_45813);
or U46221 (N_46221,N_45857,N_44176);
nand U46222 (N_46222,N_44306,N_44045);
nand U46223 (N_46223,N_45615,N_44014);
nor U46224 (N_46224,N_45288,N_44562);
xor U46225 (N_46225,N_45531,N_44967);
xor U46226 (N_46226,N_45207,N_45164);
nand U46227 (N_46227,N_44969,N_44351);
xor U46228 (N_46228,N_44154,N_45200);
xnor U46229 (N_46229,N_45741,N_44681);
nor U46230 (N_46230,N_44033,N_44486);
nand U46231 (N_46231,N_45839,N_45814);
or U46232 (N_46232,N_44987,N_44006);
nand U46233 (N_46233,N_44522,N_45269);
nor U46234 (N_46234,N_45291,N_44371);
xnor U46235 (N_46235,N_44772,N_44067);
nor U46236 (N_46236,N_44403,N_44814);
xor U46237 (N_46237,N_45552,N_44338);
xor U46238 (N_46238,N_45599,N_45780);
xor U46239 (N_46239,N_45532,N_44466);
xnor U46240 (N_46240,N_45146,N_45032);
xor U46241 (N_46241,N_45711,N_45089);
xor U46242 (N_46242,N_44706,N_44628);
and U46243 (N_46243,N_44038,N_45760);
xnor U46244 (N_46244,N_45926,N_44723);
xor U46245 (N_46245,N_45804,N_45852);
and U46246 (N_46246,N_44694,N_45276);
or U46247 (N_46247,N_45070,N_44576);
or U46248 (N_46248,N_44948,N_45533);
or U46249 (N_46249,N_44499,N_45904);
and U46250 (N_46250,N_45568,N_44667);
and U46251 (N_46251,N_45216,N_45850);
nor U46252 (N_46252,N_45841,N_45640);
and U46253 (N_46253,N_45771,N_44360);
nor U46254 (N_46254,N_45727,N_45044);
nor U46255 (N_46255,N_45309,N_45109);
xor U46256 (N_46256,N_45770,N_45689);
xor U46257 (N_46257,N_45972,N_44222);
or U46258 (N_46258,N_44512,N_45742);
nor U46259 (N_46259,N_45616,N_45134);
or U46260 (N_46260,N_44785,N_44389);
nand U46261 (N_46261,N_45628,N_44720);
and U46262 (N_46262,N_44135,N_45283);
xnor U46263 (N_46263,N_45459,N_45272);
and U46264 (N_46264,N_45239,N_45890);
nor U46265 (N_46265,N_45931,N_44700);
nor U46266 (N_46266,N_44920,N_45647);
xnor U46267 (N_46267,N_44632,N_45040);
nor U46268 (N_46268,N_44421,N_44902);
xnor U46269 (N_46269,N_44468,N_44659);
xor U46270 (N_46270,N_44944,N_45061);
xnor U46271 (N_46271,N_44424,N_44207);
and U46272 (N_46272,N_45762,N_44266);
and U46273 (N_46273,N_45054,N_44642);
and U46274 (N_46274,N_44843,N_45506);
nand U46275 (N_46275,N_44101,N_44620);
nand U46276 (N_46276,N_44740,N_44907);
xnor U46277 (N_46277,N_45411,N_45062);
and U46278 (N_46278,N_45368,N_44536);
nand U46279 (N_46279,N_45130,N_45545);
and U46280 (N_46280,N_45384,N_45029);
nor U46281 (N_46281,N_44538,N_44454);
nor U46282 (N_46282,N_44553,N_45406);
nand U46283 (N_46283,N_45826,N_45518);
nand U46284 (N_46284,N_45101,N_45913);
nand U46285 (N_46285,N_45998,N_45293);
xnor U46286 (N_46286,N_44664,N_45115);
nor U46287 (N_46287,N_44136,N_45289);
nand U46288 (N_46288,N_45392,N_45188);
and U46289 (N_46289,N_45034,N_44325);
or U46290 (N_46290,N_45419,N_44482);
nand U46291 (N_46291,N_45275,N_45736);
or U46292 (N_46292,N_45442,N_44310);
nor U46293 (N_46293,N_45719,N_45481);
xor U46294 (N_46294,N_45373,N_44529);
and U46295 (N_46295,N_45860,N_45344);
nand U46296 (N_46296,N_45953,N_45799);
and U46297 (N_46297,N_45336,N_44114);
or U46298 (N_46298,N_45983,N_44851);
or U46299 (N_46299,N_44046,N_44697);
or U46300 (N_46300,N_45605,N_44592);
nor U46301 (N_46301,N_44012,N_45312);
nand U46302 (N_46302,N_44384,N_44015);
or U46303 (N_46303,N_45630,N_45367);
xor U46304 (N_46304,N_45299,N_44370);
or U46305 (N_46305,N_45104,N_45676);
xor U46306 (N_46306,N_45985,N_45698);
and U46307 (N_46307,N_44363,N_44863);
xnor U46308 (N_46308,N_45479,N_45784);
and U46309 (N_46309,N_44796,N_45377);
nor U46310 (N_46310,N_44206,N_44662);
xor U46311 (N_46311,N_45502,N_45136);
and U46312 (N_46312,N_45827,N_44766);
or U46313 (N_46313,N_45606,N_44194);
or U46314 (N_46314,N_45975,N_44419);
or U46315 (N_46315,N_44013,N_45649);
xnor U46316 (N_46316,N_45997,N_44333);
and U46317 (N_46317,N_44314,N_44523);
and U46318 (N_46318,N_44138,N_45057);
nor U46319 (N_46319,N_44754,N_44755);
nand U46320 (N_46320,N_44750,N_44112);
nor U46321 (N_46321,N_45043,N_45713);
or U46322 (N_46322,N_45772,N_45564);
or U46323 (N_46323,N_45233,N_44852);
or U46324 (N_46324,N_45439,N_45444);
or U46325 (N_46325,N_45348,N_44304);
nand U46326 (N_46326,N_45549,N_44096);
and U46327 (N_46327,N_44686,N_44267);
nand U46328 (N_46328,N_44509,N_45855);
and U46329 (N_46329,N_45971,N_44024);
nand U46330 (N_46330,N_45872,N_45103);
and U46331 (N_46331,N_45538,N_44609);
nor U46332 (N_46332,N_44185,N_44569);
nor U46333 (N_46333,N_45990,N_45131);
nand U46334 (N_46334,N_44844,N_44385);
nand U46335 (N_46335,N_44874,N_45962);
nor U46336 (N_46336,N_45540,N_45100);
or U46337 (N_46337,N_44103,N_44956);
and U46338 (N_46338,N_44744,N_44822);
and U46339 (N_46339,N_45248,N_45327);
and U46340 (N_46340,N_44278,N_44182);
nor U46341 (N_46341,N_45844,N_45982);
nor U46342 (N_46342,N_45433,N_44379);
nand U46343 (N_46343,N_45738,N_45037);
nor U46344 (N_46344,N_45882,N_45052);
xor U46345 (N_46345,N_45422,N_45819);
nor U46346 (N_46346,N_44826,N_44275);
or U46347 (N_46347,N_44435,N_45462);
xnor U46348 (N_46348,N_45323,N_45056);
nor U46349 (N_46349,N_44433,N_44078);
xor U46350 (N_46350,N_45582,N_44407);
or U46351 (N_46351,N_44236,N_45637);
or U46352 (N_46352,N_44660,N_45112);
and U46353 (N_46353,N_44931,N_45091);
and U46354 (N_46354,N_45204,N_45405);
nand U46355 (N_46355,N_45641,N_45529);
nand U46356 (N_46356,N_44878,N_45319);
or U46357 (N_46357,N_44946,N_44105);
and U46358 (N_46358,N_44425,N_45380);
and U46359 (N_46359,N_44781,N_45491);
nand U46360 (N_46360,N_44817,N_45712);
or U46361 (N_46361,N_45768,N_44186);
nand U46362 (N_46362,N_45946,N_44238);
or U46363 (N_46363,N_45895,N_44157);
nand U46364 (N_46364,N_45598,N_44428);
nor U46365 (N_46365,N_44606,N_44568);
xor U46366 (N_46366,N_44743,N_44252);
nor U46367 (N_46367,N_44655,N_44029);
nor U46368 (N_46368,N_45524,N_45030);
xnor U46369 (N_46369,N_45527,N_44035);
xor U46370 (N_46370,N_45654,N_44286);
nor U46371 (N_46371,N_44566,N_45927);
xnor U46372 (N_46372,N_44860,N_44301);
or U46373 (N_46373,N_44985,N_45270);
or U46374 (N_46374,N_44193,N_44816);
and U46375 (N_46375,N_44048,N_45617);
xor U46376 (N_46376,N_45450,N_44765);
and U46377 (N_46377,N_45203,N_45494);
nand U46378 (N_46378,N_45682,N_44589);
nand U46379 (N_46379,N_45574,N_45967);
xnor U46380 (N_46380,N_44792,N_44413);
or U46381 (N_46381,N_45601,N_44607);
or U46382 (N_46382,N_45166,N_44790);
and U46383 (N_46383,N_45979,N_44794);
nand U46384 (N_46384,N_45498,N_44982);
or U46385 (N_46385,N_45121,N_45832);
and U46386 (N_46386,N_45964,N_44064);
or U46387 (N_46387,N_45775,N_44893);
nand U46388 (N_46388,N_45932,N_45162);
and U46389 (N_46389,N_44237,N_44085);
nand U46390 (N_46390,N_45119,N_44916);
nor U46391 (N_46391,N_44040,N_45808);
and U46392 (N_46392,N_45535,N_44353);
nand U46393 (N_46393,N_44705,N_44142);
and U46394 (N_46394,N_44836,N_44088);
or U46395 (N_46395,N_44718,N_44016);
or U46396 (N_46396,N_44732,N_45525);
and U46397 (N_46397,N_44675,N_45608);
nand U46398 (N_46398,N_45035,N_44093);
or U46399 (N_46399,N_44357,N_44962);
and U46400 (N_46400,N_44261,N_44870);
nor U46401 (N_46401,N_44719,N_44108);
xor U46402 (N_46402,N_44051,N_44656);
xor U46403 (N_46403,N_44819,N_45878);
nand U46404 (N_46404,N_44726,N_45195);
xnor U46405 (N_46405,N_45974,N_44596);
and U46406 (N_46406,N_44517,N_45243);
and U46407 (N_46407,N_44626,N_44158);
nor U46408 (N_46408,N_44244,N_45453);
and U46409 (N_46409,N_44563,N_45265);
and U46410 (N_46410,N_45023,N_44291);
nand U46411 (N_46411,N_44350,N_45510);
xnor U46412 (N_46412,N_44511,N_45757);
xnor U46413 (N_46413,N_45031,N_44935);
nor U46414 (N_46414,N_44825,N_45646);
or U46415 (N_46415,N_44809,N_44741);
and U46416 (N_46416,N_45168,N_45047);
nor U46417 (N_46417,N_44940,N_44328);
and U46418 (N_46418,N_45489,N_45728);
or U46419 (N_46419,N_44850,N_45142);
and U46420 (N_46420,N_45310,N_44094);
or U46421 (N_46421,N_44557,N_44448);
or U46422 (N_46422,N_45447,N_44610);
or U46423 (N_46423,N_44161,N_44087);
or U46424 (N_46424,N_44615,N_44636);
or U46425 (N_46425,N_45170,N_44349);
or U46426 (N_46426,N_45847,N_45938);
or U46427 (N_46427,N_45386,N_44764);
or U46428 (N_46428,N_45302,N_44525);
and U46429 (N_46429,N_45022,N_44721);
and U46430 (N_46430,N_44514,N_45095);
or U46431 (N_46431,N_44531,N_44835);
or U46432 (N_46432,N_44725,N_44980);
nor U46433 (N_46433,N_44830,N_44621);
xnor U46434 (N_46434,N_44404,N_45795);
nor U46435 (N_46435,N_44540,N_45238);
and U46436 (N_46436,N_44692,N_44515);
and U46437 (N_46437,N_44128,N_44556);
nand U46438 (N_46438,N_45970,N_45407);
xnor U46439 (N_46439,N_44184,N_44125);
or U46440 (N_46440,N_45015,N_44487);
nand U46441 (N_46441,N_44963,N_45625);
xnor U46442 (N_46442,N_45128,N_45421);
xnor U46443 (N_46443,N_44883,N_45330);
nor U46444 (N_46444,N_44380,N_44885);
nor U46445 (N_46445,N_45428,N_45298);
nor U46446 (N_46446,N_44441,N_45235);
or U46447 (N_46447,N_45295,N_44288);
or U46448 (N_46448,N_45594,N_45349);
or U46449 (N_46449,N_44871,N_45334);
xor U46450 (N_46450,N_44730,N_44868);
nand U46451 (N_46451,N_45475,N_44729);
nor U46452 (N_46452,N_44174,N_45722);
nand U46453 (N_46453,N_45071,N_45505);
or U46454 (N_46454,N_44783,N_45661);
nand U46455 (N_46455,N_45378,N_44802);
or U46456 (N_46456,N_45249,N_44469);
xor U46457 (N_46457,N_45806,N_45484);
nand U46458 (N_46458,N_44324,N_45024);
or U46459 (N_46459,N_44168,N_44254);
nand U46460 (N_46460,N_44319,N_44534);
nor U46461 (N_46461,N_45365,N_45468);
xor U46462 (N_46462,N_44865,N_44779);
nand U46463 (N_46463,N_45731,N_45547);
or U46464 (N_46464,N_45324,N_45026);
nor U46465 (N_46465,N_45496,N_44864);
nor U46466 (N_46466,N_45769,N_44395);
xor U46467 (N_46467,N_44539,N_45371);
xor U46468 (N_46468,N_44002,N_44475);
xor U46469 (N_46469,N_44260,N_45567);
nor U46470 (N_46470,N_45362,N_44905);
nand U46471 (N_46471,N_44601,N_45889);
or U46472 (N_46472,N_44580,N_45655);
xnor U46473 (N_46473,N_45412,N_45884);
xor U46474 (N_46474,N_44318,N_45252);
and U46475 (N_46475,N_44670,N_44106);
nand U46476 (N_46476,N_44284,N_44200);
nand U46477 (N_46477,N_44680,N_45118);
nand U46478 (N_46478,N_44776,N_45011);
or U46479 (N_46479,N_44005,N_45211);
or U46480 (N_46480,N_45845,N_44055);
xnor U46481 (N_46481,N_45634,N_44612);
nor U46482 (N_46482,N_45282,N_45465);
and U46483 (N_46483,N_44074,N_45820);
and U46484 (N_46484,N_44849,N_45693);
xnor U46485 (N_46485,N_45198,N_45448);
nand U46486 (N_46486,N_44383,N_44992);
xor U46487 (N_46487,N_45651,N_45160);
and U46488 (N_46488,N_44110,N_45790);
xor U46489 (N_46489,N_44388,N_45815);
xnor U46490 (N_46490,N_44156,N_44547);
and U46491 (N_46491,N_44506,N_44631);
xor U46492 (N_46492,N_45811,N_44500);
xnor U46493 (N_46493,N_45286,N_44340);
and U46494 (N_46494,N_44654,N_45969);
or U46495 (N_46495,N_44882,N_45987);
or U46496 (N_46496,N_45925,N_44204);
and U46497 (N_46497,N_44952,N_45956);
nor U46498 (N_46498,N_44248,N_45120);
nor U46499 (N_46499,N_45139,N_44330);
nor U46500 (N_46500,N_44143,N_44221);
nor U46501 (N_46501,N_45685,N_45589);
or U46502 (N_46502,N_44362,N_44996);
nand U46503 (N_46503,N_44426,N_44903);
and U46504 (N_46504,N_44652,N_45587);
xnor U46505 (N_46505,N_44657,N_44604);
nor U46506 (N_46506,N_44966,N_45332);
and U46507 (N_46507,N_45488,N_44339);
nand U46508 (N_46508,N_45704,N_44414);
nor U46509 (N_46509,N_44530,N_44797);
nand U46510 (N_46510,N_45906,N_44263);
and U46511 (N_46511,N_44786,N_45993);
or U46512 (N_46512,N_45764,N_44634);
and U46513 (N_46513,N_45179,N_45939);
and U46514 (N_46514,N_45776,N_44036);
and U46515 (N_46515,N_44008,N_45633);
nor U46516 (N_46516,N_45326,N_44827);
or U46517 (N_46517,N_45018,N_44457);
xor U46518 (N_46518,N_45194,N_44974);
and U46519 (N_46519,N_45223,N_44241);
and U46520 (N_46520,N_45765,N_44650);
nor U46521 (N_46521,N_44412,N_45180);
or U46522 (N_46522,N_45273,N_45206);
or U46523 (N_46523,N_45865,N_44030);
xor U46524 (N_46524,N_45783,N_45858);
xor U46525 (N_46525,N_45076,N_44311);
nand U46526 (N_46526,N_44289,N_45695);
and U46527 (N_46527,N_44806,N_44070);
and U46528 (N_46528,N_44513,N_45088);
nand U46529 (N_46529,N_45921,N_44565);
nor U46530 (N_46530,N_44975,N_45381);
nor U46531 (N_46531,N_44671,N_44904);
and U46532 (N_46532,N_44181,N_44131);
or U46533 (N_46533,N_44047,N_44505);
and U46534 (N_46534,N_44734,N_45585);
nor U46535 (N_46535,N_44364,N_44450);
and U46536 (N_46536,N_44577,N_45048);
xnor U46537 (N_46537,N_44139,N_45250);
xor U46538 (N_46538,N_44122,N_44605);
xor U46539 (N_46539,N_44417,N_45732);
and U46540 (N_46540,N_45579,N_44264);
or U46541 (N_46541,N_44003,N_45036);
nor U46542 (N_46542,N_45907,N_45644);
and U46543 (N_46543,N_45218,N_45619);
and U46544 (N_46544,N_44923,N_45520);
and U46545 (N_46545,N_44867,N_44240);
nand U46546 (N_46546,N_44570,N_45014);
nor U46547 (N_46547,N_45267,N_44742);
nand U46548 (N_46548,N_45803,N_44305);
xor U46549 (N_46549,N_45548,N_44839);
and U46550 (N_46550,N_44179,N_45455);
or U46551 (N_46551,N_44082,N_44753);
nor U46552 (N_46552,N_45905,N_44622);
nor U46553 (N_46553,N_44542,N_44752);
or U46554 (N_46554,N_44716,N_44960);
or U46555 (N_46555,N_45132,N_44668);
and U46556 (N_46556,N_45748,N_44496);
and U46557 (N_46557,N_45229,N_44160);
nand U46558 (N_46558,N_45836,N_45755);
nor U46559 (N_46559,N_44120,N_44098);
and U46560 (N_46560,N_45577,N_44255);
or U46561 (N_46561,N_44876,N_45110);
nor U46562 (N_46562,N_44262,N_44335);
nand U46563 (N_46563,N_44296,N_45473);
xnor U46564 (N_46564,N_44945,N_44912);
nor U46565 (N_46565,N_44151,N_45678);
and U46566 (N_46566,N_45158,N_45861);
or U46567 (N_46567,N_45241,N_45613);
and U46568 (N_46568,N_45778,N_45111);
or U46569 (N_46569,N_45141,N_45837);
xnor U46570 (N_46570,N_44875,N_45937);
and U46571 (N_46571,N_45436,N_44218);
nor U46572 (N_46572,N_44129,N_45372);
nand U46573 (N_46573,N_44608,N_44294);
or U46574 (N_46574,N_45400,N_45236);
xnor U46575 (N_46575,N_45137,N_44408);
xor U46576 (N_46576,N_45515,N_44124);
nor U46577 (N_46577,N_44180,N_45739);
nand U46578 (N_46578,N_44422,N_44559);
and U46579 (N_46579,N_44676,N_45514);
or U46580 (N_46580,N_45300,N_44258);
xnor U46581 (N_46581,N_45352,N_45074);
nor U46582 (N_46582,N_45078,N_45692);
xor U46583 (N_46583,N_44405,N_45930);
or U46584 (N_46584,N_45102,N_44233);
xor U46585 (N_46585,N_44953,N_44981);
and U46586 (N_46586,N_44493,N_44479);
or U46587 (N_46587,N_45740,N_45716);
or U46588 (N_46588,N_45888,N_44921);
and U46589 (N_46589,N_44355,N_45659);
nand U46590 (N_46590,N_45213,N_45476);
or U46591 (N_46591,N_45457,N_44480);
nor U46592 (N_46592,N_44838,N_44595);
and U46593 (N_46593,N_45437,N_44444);
or U46594 (N_46594,N_44593,N_45563);
and U46595 (N_46595,N_45278,N_44178);
nand U46596 (N_46596,N_44581,N_45467);
and U46597 (N_46597,N_45050,N_45667);
nor U46598 (N_46598,N_44763,N_45333);
xor U46599 (N_46599,N_44862,N_44774);
and U46600 (N_46600,N_44658,N_44665);
or U46601 (N_46601,N_44972,N_45584);
and U46602 (N_46602,N_45106,N_45363);
and U46603 (N_46603,N_44100,N_45825);
nand U46604 (N_46604,N_45366,N_45125);
and U46605 (N_46605,N_45454,N_45557);
nand U46606 (N_46606,N_44242,N_45345);
nand U46607 (N_46607,N_45003,N_44748);
or U46608 (N_46608,N_45639,N_45994);
nor U46609 (N_46609,N_45108,N_45417);
or U46610 (N_46610,N_44434,N_44464);
and U46611 (N_46611,N_45002,N_45758);
and U46612 (N_46612,N_44840,N_44551);
nand U46613 (N_46613,N_45854,N_44054);
nor U46614 (N_46614,N_45672,N_44698);
and U46615 (N_46615,N_45870,N_44366);
or U46616 (N_46616,N_45263,N_44869);
or U46617 (N_46617,N_45152,N_44898);
or U46618 (N_46618,N_45597,N_44856);
or U46619 (N_46619,N_44246,N_45954);
nand U46620 (N_46620,N_45090,N_45237);
xnor U46621 (N_46621,N_45853,N_45261);
nand U46622 (N_46622,N_45338,N_45656);
or U46623 (N_46623,N_45724,N_44080);
xor U46624 (N_46624,N_44810,N_45337);
nor U46625 (N_46625,N_45869,N_44999);
nor U46626 (N_46626,N_45191,N_44155);
nand U46627 (N_46627,N_44846,N_44192);
and U46628 (N_46628,N_45941,N_44702);
xnor U46629 (N_46629,N_45315,N_44401);
xnor U46630 (N_46630,N_45423,N_45668);
xor U46631 (N_46631,N_44761,N_44599);
or U46632 (N_46632,N_44854,N_45543);
nand U46633 (N_46633,N_44687,N_44494);
xor U46634 (N_46634,N_44411,N_45387);
xnor U46635 (N_46635,N_44990,N_44757);
xor U46636 (N_46636,N_44630,N_44065);
nor U46637 (N_46637,N_45307,N_45005);
and U46638 (N_46638,N_45721,N_45508);
nor U46639 (N_46639,N_45960,N_45916);
or U46640 (N_46640,N_45620,N_44092);
nor U46641 (N_46641,N_45965,N_45446);
or U46642 (N_46642,N_44778,N_45976);
nor U46643 (N_46643,N_44490,N_44378);
xor U46644 (N_46644,N_44461,N_45266);
xnor U46645 (N_46645,N_45881,N_44791);
nand U46646 (N_46646,N_45945,N_44768);
or U46647 (N_46647,N_45360,N_44459);
nand U46648 (N_46648,N_45624,N_45952);
and U46649 (N_46649,N_45546,N_44954);
nand U46650 (N_46650,N_45306,N_45325);
and U46651 (N_46651,N_45849,N_45094);
nor U46652 (N_46652,N_45049,N_44191);
xor U46653 (N_46653,N_44477,N_45892);
nor U46654 (N_46654,N_45669,N_44043);
nand U46655 (N_46655,N_44558,N_44057);
nand U46656 (N_46656,N_45511,N_44042);
and U46657 (N_46657,N_44811,N_45631);
nor U46658 (N_46658,N_44777,N_45251);
xnor U46659 (N_46659,N_45991,N_44451);
xor U46660 (N_46660,N_45873,N_45331);
nor U46661 (N_46661,N_45082,N_44947);
nor U46662 (N_46662,N_44021,N_45897);
nor U46663 (N_46663,N_45963,N_45027);
nand U46664 (N_46664,N_45463,N_45480);
nand U46665 (N_46665,N_44337,N_44703);
or U46666 (N_46666,N_45350,N_44150);
xor U46667 (N_46667,N_45581,N_44372);
nand U46668 (N_46668,N_45150,N_44879);
or U46669 (N_46669,N_45816,N_45149);
and U46670 (N_46670,N_44978,N_45155);
or U46671 (N_46671,N_45469,N_44465);
xor U46672 (N_46672,N_45875,N_44861);
and U46673 (N_46673,N_44892,N_45673);
nand U46674 (N_46674,N_45355,N_44453);
nor U46675 (N_46675,N_44472,N_45138);
and U46676 (N_46676,N_45729,N_44829);
xnor U46677 (N_46677,N_45039,N_44602);
nor U46678 (N_46678,N_45700,N_44066);
xnor U46679 (N_46679,N_45393,N_44273);
nand U46680 (N_46680,N_44369,N_45290);
xnor U46681 (N_46681,N_44918,N_45835);
nand U46682 (N_46682,N_44520,N_44257);
and U46683 (N_46683,N_45356,N_44053);
nand U46684 (N_46684,N_44573,N_45214);
and U46685 (N_46685,N_45745,N_44028);
nor U46686 (N_46686,N_45060,N_45181);
and U46687 (N_46687,N_44056,N_45580);
xor U46688 (N_46688,N_44993,N_45072);
nor U46689 (N_46689,N_44109,N_44488);
and U46690 (N_46690,N_44492,N_45124);
xnor U46691 (N_46691,N_45626,N_44452);
xnor U46692 (N_46692,N_44004,N_44470);
nor U46693 (N_46693,N_45486,N_45793);
or U46694 (N_46694,N_45512,N_45717);
nor U46695 (N_46695,N_44099,N_45280);
nor U46696 (N_46696,N_45192,N_44647);
xor U46697 (N_46697,N_45409,N_45670);
or U46698 (N_46698,N_45973,N_44141);
nor U46699 (N_46699,N_44187,N_45208);
and U46700 (N_46700,N_45909,N_45922);
or U46701 (N_46701,N_45848,N_45984);
and U46702 (N_46702,N_45950,N_45559);
xor U46703 (N_46703,N_44888,N_44227);
or U46704 (N_46704,N_45830,N_44346);
or U46705 (N_46705,N_44611,N_45209);
nor U46706 (N_46706,N_45490,N_45190);
or U46707 (N_46707,N_45354,N_45706);
or U46708 (N_46708,N_45565,N_45320);
xor U46709 (N_46709,N_44859,N_45274);
xnor U46710 (N_46710,N_44429,N_44077);
nand U46711 (N_46711,N_45522,N_44503);
and U46712 (N_46712,N_45172,N_45665);
xor U46713 (N_46713,N_45477,N_45715);
and U46714 (N_46714,N_44624,N_44210);
nand U46715 (N_46715,N_44832,N_44073);
or U46716 (N_46716,N_44695,N_44709);
nand U46717 (N_46717,N_44090,N_44590);
and U46718 (N_46718,N_44467,N_45725);
and U46719 (N_46719,N_45750,N_45603);
or U46720 (N_46720,N_44881,N_45802);
nand U46721 (N_46721,N_44619,N_45959);
or U46722 (N_46722,N_45886,N_44805);
and U46723 (N_46723,N_44661,N_44841);
nand U46724 (N_46724,N_45773,N_45478);
and U46725 (N_46725,N_45681,N_44137);
and U46726 (N_46726,N_44617,N_44485);
and U46727 (N_46727,N_44039,N_45140);
or U46728 (N_46728,N_45197,N_44463);
nor U46729 (N_46729,N_44693,N_45341);
and U46730 (N_46730,N_45081,N_44738);
nor U46731 (N_46731,N_45222,N_45205);
and U46732 (N_46732,N_45308,N_44815);
nand U46733 (N_46733,N_45055,N_44437);
xor U46734 (N_46734,N_44000,N_45663);
or U46735 (N_46735,N_45838,N_45328);
xor U46736 (N_46736,N_45851,N_44943);
or U46737 (N_46737,N_44701,N_44684);
and U46738 (N_46738,N_44504,N_45789);
xnor U46739 (N_46739,N_45084,N_44988);
nand U46740 (N_46740,N_44873,N_44276);
nor U46741 (N_46741,N_44416,N_45435);
nand U46742 (N_46742,N_44344,N_45296);
xor U46743 (N_46743,N_44292,N_44219);
nor U46744 (N_46744,N_45652,N_44707);
xnor U46745 (N_46745,N_45231,N_45779);
xor U46746 (N_46746,N_44025,N_44095);
and U46747 (N_46747,N_44579,N_45370);
nor U46748 (N_46748,N_45899,N_45184);
and U46749 (N_46749,N_44648,N_44555);
nand U46750 (N_46750,N_45751,N_44022);
xor U46751 (N_46751,N_44638,N_45876);
and U46752 (N_46752,N_45915,N_44195);
xor U46753 (N_46753,N_45201,N_45928);
nor U46754 (N_46754,N_44001,N_45812);
and U46755 (N_46755,N_44149,N_44119);
and U46756 (N_46756,N_45182,N_44672);
xnor U46757 (N_46757,N_44784,N_45173);
nand U46758 (N_46758,N_44280,N_45105);
or U46759 (N_46759,N_45389,N_45415);
nand U46760 (N_46760,N_45523,N_44949);
xor U46761 (N_46761,N_45702,N_44265);
and U46762 (N_46762,N_45863,N_45912);
or U46763 (N_46763,N_44973,N_45240);
and U46764 (N_46764,N_44431,N_44432);
nand U46765 (N_46765,N_44788,N_45153);
nand U46766 (N_46766,N_44733,N_45253);
xnor U46767 (N_46767,N_45501,N_44104);
or U46768 (N_46768,N_44212,N_44666);
nand U46769 (N_46769,N_44188,N_44535);
nand U46770 (N_46770,N_44049,N_44365);
nand U46771 (N_46771,N_44415,N_45189);
or U46772 (N_46772,N_45217,N_45145);
nand U46773 (N_46773,N_45499,N_45575);
nor U46774 (N_46774,N_45821,N_45553);
xnor U46775 (N_46775,N_44121,N_44170);
nand U46776 (N_46776,N_44813,N_45431);
and U46777 (N_46777,N_44603,N_44977);
or U46778 (N_46778,N_44175,N_45245);
or U46779 (N_46779,N_44199,N_45650);
nor U46780 (N_46780,N_45020,N_45788);
xor U46781 (N_46781,N_45364,N_45316);
xor U46782 (N_46782,N_44062,N_44361);
nand U46783 (N_46783,N_45202,N_45254);
nor U46784 (N_46784,N_44341,N_45828);
and U46785 (N_46785,N_45143,N_44691);
nor U46786 (N_46786,N_45759,N_45942);
nand U46787 (N_46787,N_44484,N_45593);
or U46788 (N_46788,N_44727,N_45019);
or U46789 (N_46789,N_45343,N_44279);
nor U46790 (N_46790,N_44521,N_45817);
and U46791 (N_46791,N_45782,N_45099);
xor U46792 (N_46792,N_45632,N_44927);
xor U46793 (N_46793,N_44489,N_45566);
nor U46794 (N_46794,N_44922,N_44247);
or U46795 (N_46795,N_45430,N_45177);
nor U46796 (N_46796,N_44798,N_45399);
or U46797 (N_46797,N_44234,N_45171);
or U46798 (N_46798,N_45718,N_44651);
xor U46799 (N_46799,N_44172,N_45414);
nand U46800 (N_46800,N_44402,N_44961);
or U46801 (N_46801,N_45595,N_45774);
or U46802 (N_46802,N_45485,N_44582);
nand U46803 (N_46803,N_44646,N_45703);
and U46804 (N_46804,N_44939,N_45934);
xor U46805 (N_46805,N_45571,N_45311);
or U46806 (N_46806,N_45986,N_44071);
nand U46807 (N_46807,N_45083,N_44235);
or U46808 (N_46808,N_44578,N_44290);
nand U46809 (N_46809,N_45679,N_45792);
nor U46810 (N_46810,N_44409,N_44587);
nand U46811 (N_46811,N_44037,N_44994);
or U46812 (N_46812,N_45077,N_45539);
nor U46813 (N_46813,N_45318,N_44377);
or U46814 (N_46814,N_45609,N_44780);
xor U46815 (N_46815,N_45614,N_44745);
and U46816 (N_46816,N_44913,N_45051);
nand U46817 (N_46817,N_44495,N_45840);
nand U46818 (N_46818,N_45069,N_44323);
and U46819 (N_46819,N_44554,N_44213);
and U46820 (N_46820,N_45427,N_45210);
xor U46821 (N_46821,N_45978,N_44845);
nand U46822 (N_46822,N_44527,N_45796);
xnor U46823 (N_46823,N_44986,N_45452);
and U46824 (N_46824,N_45753,N_45786);
and U46825 (N_46825,N_44951,N_45867);
or U46826 (N_46826,N_44731,N_44243);
nor U46827 (N_46827,N_44460,N_45403);
and U46828 (N_46828,N_45305,N_44507);
nor U46829 (N_46829,N_45995,N_44201);
or U46830 (N_46830,N_44689,N_44930);
xnor U46831 (N_46831,N_45940,N_45175);
or U46832 (N_46832,N_44548,N_44163);
or U46833 (N_46833,N_45968,N_44837);
or U46834 (N_46834,N_45242,N_45129);
or U46835 (N_46835,N_45920,N_45735);
and U46836 (N_46836,N_45611,N_44367);
or U46837 (N_46837,N_45461,N_44196);
or U46838 (N_46838,N_44704,N_44134);
and U46839 (N_46839,N_45287,N_45910);
or U46840 (N_46840,N_45781,N_45369);
nor U46841 (N_46841,N_45824,N_45513);
xor U46842 (N_46842,N_44285,N_45917);
nand U46843 (N_46843,N_44123,N_44793);
nor U46844 (N_46844,N_44591,N_44336);
xor U46845 (N_46845,N_45135,N_44584);
nand U46846 (N_46846,N_45394,N_45434);
nor U46847 (N_46847,N_44560,N_45046);
and U46848 (N_46848,N_45785,N_44476);
nor U46849 (N_46849,N_44997,N_44831);
and U46850 (N_46850,N_44399,N_45413);
xor U46851 (N_46851,N_44834,N_44358);
or U46852 (N_46852,N_44231,N_44801);
or U46853 (N_46853,N_44332,N_45321);
xor U46854 (N_46854,N_44052,N_45045);
nand U46855 (N_46855,N_45466,N_44724);
xor U46856 (N_46856,N_44644,N_45012);
or U46857 (N_46857,N_44751,N_44373);
or U46858 (N_46858,N_45536,N_44458);
nor U46859 (N_46859,N_45551,N_45410);
and U46860 (N_46860,N_44911,N_44908);
nor U46861 (N_46861,N_45176,N_45395);
nor U46862 (N_46862,N_44896,N_44594);
nor U46863 (N_46863,N_44225,N_45396);
nand U46864 (N_46864,N_44113,N_45809);
nand U46865 (N_46865,N_44343,N_45260);
and U46866 (N_46866,N_44117,N_44984);
xor U46867 (N_46867,N_44717,N_44302);
and U46868 (N_46868,N_44759,N_45258);
nand U46869 (N_46869,N_45376,N_44543);
and U46870 (N_46870,N_44713,N_44623);
nand U46871 (N_46871,N_44075,N_45818);
nor U46872 (N_46872,N_44663,N_45696);
and U46873 (N_46873,N_44223,N_44887);
nor U46874 (N_46874,N_45154,N_44669);
xor U46875 (N_46875,N_44321,N_44381);
xnor U46876 (N_46876,N_45144,N_45602);
nand U46877 (N_46877,N_45746,N_45578);
nor U46878 (N_46878,N_44572,N_44532);
nand U46879 (N_46879,N_45896,N_44322);
or U46880 (N_46880,N_44162,N_44909);
nand U46881 (N_46881,N_44474,N_44897);
and U46882 (N_46882,N_44890,N_45178);
nand U46883 (N_46883,N_44326,N_45604);
or U46884 (N_46884,N_44571,N_44857);
and U46885 (N_46885,N_45041,N_44803);
xnor U46886 (N_46886,N_45898,N_45924);
or U46887 (N_46887,N_45893,N_45147);
xor U46888 (N_46888,N_45627,N_44297);
nand U46889 (N_46889,N_44023,N_44937);
nor U46890 (N_46890,N_45666,N_44166);
nand U46891 (N_46891,N_45709,N_45951);
and U46892 (N_46892,N_44497,N_45053);
nor U46893 (N_46893,N_45425,N_45001);
and U46894 (N_46894,N_44848,N_44390);
nand U46895 (N_46895,N_45688,N_44933);
nand U46896 (N_46896,N_44629,N_44282);
and U46897 (N_46897,N_45911,N_44410);
or U46898 (N_46898,N_44027,N_45073);
xnor U46899 (N_46899,N_44420,N_44447);
xor U46900 (N_46900,N_44209,N_44217);
and U46901 (N_46901,N_44295,N_45087);
nor U46902 (N_46902,N_45244,N_44899);
xor U46903 (N_46903,N_45763,N_44256);
nand U46904 (N_46904,N_45335,N_44068);
or U46905 (N_46905,N_45010,N_44308);
nor U46906 (N_46906,N_44061,N_44202);
and U46907 (N_46907,N_44189,N_44127);
or U46908 (N_46908,N_44653,N_44564);
xor U46909 (N_46909,N_44760,N_44019);
xor U46910 (N_46910,N_44483,N_45797);
and U46911 (N_46911,N_45021,N_45116);
xor U46912 (N_46912,N_44775,N_44334);
nand U46913 (N_46913,N_45358,N_44640);
nand U46914 (N_46914,N_44866,N_45530);
nand U46915 (N_46915,N_45482,N_45556);
nand U46916 (N_46916,N_44715,N_45846);
xnor U46917 (N_46917,N_44737,N_45313);
and U46918 (N_46918,N_45383,N_45013);
nand U46919 (N_46919,N_45622,N_45301);
nor U46920 (N_46920,N_45958,N_45000);
nand U46921 (N_46921,N_45636,N_45576);
nor U46922 (N_46922,N_45623,N_45919);
or U46923 (N_46923,N_44190,N_44910);
nand U46924 (N_46924,N_45064,N_44215);
nor U46925 (N_46925,N_45068,N_44317);
nor U46926 (N_46926,N_44739,N_44842);
or U46927 (N_46927,N_44635,N_44597);
nand U46928 (N_46928,N_44685,N_45493);
or U46929 (N_46929,N_44895,N_45737);
and U46930 (N_46930,N_45079,N_45183);
nor U46931 (N_46931,N_44299,N_44950);
and U46932 (N_46932,N_45016,N_44959);
xnor U46933 (N_46933,N_45284,N_44799);
nand U46934 (N_46934,N_44804,N_45767);
xor U46935 (N_46935,N_44938,N_45705);
and U46936 (N_46936,N_44891,N_44598);
xnor U46937 (N_46937,N_44767,N_45492);
or U46938 (N_46938,N_45075,N_45451);
and U46939 (N_46939,N_45944,N_45618);
xnor U46940 (N_46940,N_44820,N_44884);
and U46941 (N_46941,N_45572,N_45866);
nand U46942 (N_46942,N_44808,N_44041);
or U46943 (N_46943,N_45635,N_44376);
xor U46944 (N_46944,N_45834,N_45694);
nand U46945 (N_46945,N_45346,N_45351);
nor U46946 (N_46946,N_45691,N_44574);
or U46947 (N_46947,N_44327,N_45374);
xor U46948 (N_46948,N_44807,N_44091);
xnor U46949 (N_46949,N_44386,N_45710);
and U46950 (N_46950,N_44645,N_44044);
and U46951 (N_46951,N_44758,N_44600);
or U46952 (N_46952,N_44728,N_45908);
nand U46953 (N_46953,N_44575,N_44546);
xor U46954 (N_46954,N_44115,N_44126);
nor U46955 (N_46955,N_45098,N_44374);
and U46956 (N_46956,N_45645,N_44901);
xor U46957 (N_46957,N_45903,N_44354);
or U46958 (N_46958,N_45440,N_44688);
nor U46959 (N_46959,N_44855,N_45314);
or U46960 (N_46960,N_44989,N_44677);
xnor U46961 (N_46961,N_45607,N_45196);
and U46962 (N_46962,N_45123,N_45648);
xnor U46963 (N_46963,N_44537,N_45009);
or U46964 (N_46964,N_45610,N_44216);
nand U46965 (N_46965,N_44872,N_45375);
nor U46966 (N_46966,N_44473,N_45127);
nor U46967 (N_46967,N_45989,N_45612);
xnor U46968 (N_46968,N_45471,N_45699);
nor U46969 (N_46969,N_44561,N_45528);
nand U46970 (N_46970,N_44352,N_44519);
nor U46971 (N_46971,N_44159,N_44020);
and U46972 (N_46972,N_44303,N_44524);
and U46973 (N_46973,N_44588,N_44083);
nand U46974 (N_46974,N_45212,N_44478);
and U46975 (N_46975,N_44298,N_45004);
nand U46976 (N_46976,N_44249,N_45887);
nand U46977 (N_46977,N_45664,N_45246);
and U46978 (N_46978,N_45432,N_44152);
and U46979 (N_46979,N_44769,N_45638);
nand U46980 (N_46980,N_44533,N_45569);
and U46981 (N_46981,N_44058,N_45058);
nor U46982 (N_46982,N_45497,N_44445);
nor U46983 (N_46983,N_44331,N_44550);
nand U46984 (N_46984,N_44145,N_44060);
and U46985 (N_46985,N_45977,N_45006);
and U46986 (N_46986,N_45801,N_45948);
and U46987 (N_46987,N_45397,N_44081);
nand U46988 (N_46988,N_44616,N_45304);
or U46989 (N_46989,N_44771,N_45588);
or U46990 (N_46990,N_45257,N_45943);
xor U46991 (N_46991,N_44312,N_45936);
xnor U46992 (N_46992,N_44926,N_44643);
or U46993 (N_46993,N_45874,N_45883);
nand U46994 (N_46994,N_45829,N_44320);
nand U46995 (N_46995,N_44146,N_44198);
xor U46996 (N_46996,N_45744,N_45794);
and U46997 (N_46997,N_45561,N_45219);
or U46998 (N_46998,N_44773,N_44714);
or U46999 (N_46999,N_44735,N_45957);
or U47000 (N_47000,N_44985,N_44125);
nor U47001 (N_47001,N_44593,N_44731);
nor U47002 (N_47002,N_45299,N_45569);
nor U47003 (N_47003,N_45447,N_45274);
nor U47004 (N_47004,N_44951,N_44160);
nand U47005 (N_47005,N_44028,N_44644);
and U47006 (N_47006,N_45798,N_44496);
xnor U47007 (N_47007,N_45958,N_45567);
and U47008 (N_47008,N_45235,N_45968);
and U47009 (N_47009,N_44550,N_44629);
nand U47010 (N_47010,N_44082,N_45616);
or U47011 (N_47011,N_44781,N_44744);
nor U47012 (N_47012,N_44255,N_44108);
nand U47013 (N_47013,N_45124,N_45306);
or U47014 (N_47014,N_44709,N_45448);
or U47015 (N_47015,N_45414,N_45603);
nand U47016 (N_47016,N_45840,N_44408);
nand U47017 (N_47017,N_44890,N_45335);
and U47018 (N_47018,N_44215,N_44473);
or U47019 (N_47019,N_44702,N_45551);
nand U47020 (N_47020,N_45456,N_45554);
and U47021 (N_47021,N_45750,N_44594);
nand U47022 (N_47022,N_44047,N_45702);
and U47023 (N_47023,N_44595,N_44506);
and U47024 (N_47024,N_44792,N_45355);
xor U47025 (N_47025,N_44815,N_45989);
xnor U47026 (N_47026,N_45518,N_44395);
or U47027 (N_47027,N_44541,N_45347);
xor U47028 (N_47028,N_45924,N_45403);
nand U47029 (N_47029,N_44623,N_44632);
and U47030 (N_47030,N_45401,N_45468);
nand U47031 (N_47031,N_45621,N_45183);
and U47032 (N_47032,N_44382,N_44989);
nor U47033 (N_47033,N_45035,N_45513);
xor U47034 (N_47034,N_45469,N_44964);
nor U47035 (N_47035,N_45594,N_44322);
and U47036 (N_47036,N_44964,N_45136);
or U47037 (N_47037,N_44359,N_44099);
and U47038 (N_47038,N_44069,N_45527);
nor U47039 (N_47039,N_44311,N_44742);
or U47040 (N_47040,N_44889,N_44687);
nand U47041 (N_47041,N_44955,N_44891);
or U47042 (N_47042,N_44593,N_45667);
nor U47043 (N_47043,N_44985,N_45116);
xnor U47044 (N_47044,N_44533,N_44563);
or U47045 (N_47045,N_45244,N_44366);
nand U47046 (N_47046,N_45995,N_45063);
nor U47047 (N_47047,N_44182,N_44390);
and U47048 (N_47048,N_45165,N_45208);
and U47049 (N_47049,N_45459,N_44121);
and U47050 (N_47050,N_45767,N_45812);
or U47051 (N_47051,N_45366,N_45026);
xnor U47052 (N_47052,N_44871,N_45100);
nor U47053 (N_47053,N_45993,N_44307);
nand U47054 (N_47054,N_45890,N_45143);
nor U47055 (N_47055,N_44592,N_45739);
and U47056 (N_47056,N_45456,N_44981);
and U47057 (N_47057,N_44882,N_45637);
and U47058 (N_47058,N_44252,N_44124);
and U47059 (N_47059,N_45464,N_45010);
xnor U47060 (N_47060,N_45946,N_44767);
nand U47061 (N_47061,N_44391,N_45899);
and U47062 (N_47062,N_45998,N_44271);
nor U47063 (N_47063,N_45371,N_44136);
or U47064 (N_47064,N_44019,N_44577);
or U47065 (N_47065,N_44445,N_44612);
nor U47066 (N_47066,N_45426,N_45522);
and U47067 (N_47067,N_45599,N_45211);
or U47068 (N_47068,N_44912,N_45371);
nor U47069 (N_47069,N_45741,N_45110);
and U47070 (N_47070,N_44584,N_45853);
or U47071 (N_47071,N_45386,N_44650);
nand U47072 (N_47072,N_44639,N_44178);
or U47073 (N_47073,N_45234,N_45598);
nand U47074 (N_47074,N_45332,N_44854);
nor U47075 (N_47075,N_45991,N_45552);
or U47076 (N_47076,N_45609,N_45223);
and U47077 (N_47077,N_44633,N_45647);
nand U47078 (N_47078,N_44304,N_44862);
nand U47079 (N_47079,N_44762,N_44623);
and U47080 (N_47080,N_45828,N_44463);
xor U47081 (N_47081,N_44574,N_44977);
or U47082 (N_47082,N_44717,N_44747);
or U47083 (N_47083,N_44926,N_45264);
nand U47084 (N_47084,N_44604,N_44711);
nand U47085 (N_47085,N_44630,N_45971);
nand U47086 (N_47086,N_45297,N_44371);
and U47087 (N_47087,N_44910,N_44462);
nand U47088 (N_47088,N_45883,N_44512);
or U47089 (N_47089,N_45876,N_45411);
nand U47090 (N_47090,N_44700,N_45632);
nor U47091 (N_47091,N_44335,N_44975);
xor U47092 (N_47092,N_44995,N_44119);
nand U47093 (N_47093,N_44352,N_45867);
nand U47094 (N_47094,N_44062,N_44916);
and U47095 (N_47095,N_44620,N_44662);
xor U47096 (N_47096,N_45966,N_45400);
nand U47097 (N_47097,N_44355,N_45442);
xnor U47098 (N_47098,N_44502,N_44440);
nor U47099 (N_47099,N_45285,N_45547);
nand U47100 (N_47100,N_45675,N_45771);
and U47101 (N_47101,N_45683,N_45839);
xor U47102 (N_47102,N_45913,N_45596);
and U47103 (N_47103,N_44097,N_44666);
xnor U47104 (N_47104,N_45950,N_45382);
or U47105 (N_47105,N_44851,N_45610);
nor U47106 (N_47106,N_44554,N_45555);
and U47107 (N_47107,N_45856,N_44067);
nand U47108 (N_47108,N_44823,N_44835);
nand U47109 (N_47109,N_45027,N_45553);
nor U47110 (N_47110,N_44607,N_45310);
nand U47111 (N_47111,N_44962,N_45444);
nor U47112 (N_47112,N_45159,N_45982);
nor U47113 (N_47113,N_44456,N_44980);
xor U47114 (N_47114,N_45164,N_44220);
nand U47115 (N_47115,N_45919,N_45651);
xnor U47116 (N_47116,N_44704,N_45771);
nand U47117 (N_47117,N_45684,N_44030);
and U47118 (N_47118,N_45142,N_44873);
or U47119 (N_47119,N_45815,N_44767);
or U47120 (N_47120,N_45178,N_45834);
or U47121 (N_47121,N_44222,N_44273);
nor U47122 (N_47122,N_45041,N_45824);
or U47123 (N_47123,N_45718,N_44923);
and U47124 (N_47124,N_44605,N_45434);
xnor U47125 (N_47125,N_45825,N_44083);
xor U47126 (N_47126,N_45529,N_45764);
or U47127 (N_47127,N_45402,N_44991);
and U47128 (N_47128,N_45415,N_45566);
or U47129 (N_47129,N_45458,N_44298);
nor U47130 (N_47130,N_45650,N_44137);
xor U47131 (N_47131,N_45555,N_44490);
xor U47132 (N_47132,N_44180,N_44832);
nor U47133 (N_47133,N_44159,N_44263);
or U47134 (N_47134,N_44017,N_44949);
and U47135 (N_47135,N_45235,N_44927);
nand U47136 (N_47136,N_44859,N_45137);
xor U47137 (N_47137,N_45551,N_45557);
xnor U47138 (N_47138,N_45166,N_45280);
xor U47139 (N_47139,N_44404,N_45863);
nand U47140 (N_47140,N_45650,N_45266);
nor U47141 (N_47141,N_44094,N_44785);
nand U47142 (N_47142,N_45430,N_45419);
and U47143 (N_47143,N_45162,N_45998);
nor U47144 (N_47144,N_44292,N_44217);
nand U47145 (N_47145,N_44219,N_45125);
xnor U47146 (N_47146,N_44099,N_45737);
or U47147 (N_47147,N_44933,N_44872);
xor U47148 (N_47148,N_44851,N_45653);
nand U47149 (N_47149,N_44200,N_44593);
or U47150 (N_47150,N_44181,N_44035);
nand U47151 (N_47151,N_44423,N_44458);
nand U47152 (N_47152,N_45878,N_45128);
and U47153 (N_47153,N_45586,N_45406);
and U47154 (N_47154,N_45396,N_45839);
and U47155 (N_47155,N_44496,N_44168);
and U47156 (N_47156,N_44336,N_45618);
xnor U47157 (N_47157,N_45348,N_45422);
nand U47158 (N_47158,N_45201,N_45988);
nor U47159 (N_47159,N_44004,N_45580);
xnor U47160 (N_47160,N_45384,N_45581);
or U47161 (N_47161,N_45659,N_45096);
nor U47162 (N_47162,N_44030,N_45336);
nor U47163 (N_47163,N_45666,N_45745);
xnor U47164 (N_47164,N_44715,N_44460);
xor U47165 (N_47165,N_45723,N_44071);
nor U47166 (N_47166,N_45560,N_44354);
or U47167 (N_47167,N_44626,N_45599);
and U47168 (N_47168,N_44317,N_45089);
nand U47169 (N_47169,N_45250,N_44619);
or U47170 (N_47170,N_45853,N_45752);
nor U47171 (N_47171,N_44617,N_44755);
or U47172 (N_47172,N_44772,N_45818);
xor U47173 (N_47173,N_45746,N_45626);
nand U47174 (N_47174,N_44340,N_45829);
nor U47175 (N_47175,N_44192,N_44502);
or U47176 (N_47176,N_44187,N_45926);
nand U47177 (N_47177,N_45901,N_45023);
nor U47178 (N_47178,N_44922,N_45440);
or U47179 (N_47179,N_45722,N_45889);
xor U47180 (N_47180,N_44080,N_44065);
and U47181 (N_47181,N_45742,N_44211);
xor U47182 (N_47182,N_44508,N_45492);
nor U47183 (N_47183,N_45585,N_44992);
nor U47184 (N_47184,N_45622,N_44952);
nand U47185 (N_47185,N_45652,N_44715);
nand U47186 (N_47186,N_44762,N_44840);
nor U47187 (N_47187,N_44126,N_45314);
nand U47188 (N_47188,N_44197,N_45197);
or U47189 (N_47189,N_44739,N_45026);
nand U47190 (N_47190,N_44830,N_44328);
or U47191 (N_47191,N_45728,N_45425);
nor U47192 (N_47192,N_45028,N_45026);
and U47193 (N_47193,N_45928,N_45142);
nand U47194 (N_47194,N_44924,N_44507);
nand U47195 (N_47195,N_44648,N_45105);
or U47196 (N_47196,N_44170,N_44042);
and U47197 (N_47197,N_44240,N_44990);
or U47198 (N_47198,N_45177,N_44477);
xor U47199 (N_47199,N_45338,N_45530);
xnor U47200 (N_47200,N_44172,N_45052);
nand U47201 (N_47201,N_44805,N_44266);
nor U47202 (N_47202,N_44337,N_44080);
or U47203 (N_47203,N_44217,N_45491);
and U47204 (N_47204,N_44636,N_45882);
and U47205 (N_47205,N_45633,N_44701);
nor U47206 (N_47206,N_44000,N_45201);
and U47207 (N_47207,N_45835,N_44332);
xnor U47208 (N_47208,N_44107,N_44432);
nand U47209 (N_47209,N_45717,N_45848);
or U47210 (N_47210,N_45782,N_44370);
nor U47211 (N_47211,N_45036,N_44327);
nand U47212 (N_47212,N_44282,N_44912);
xnor U47213 (N_47213,N_45554,N_45010);
or U47214 (N_47214,N_44521,N_44904);
nor U47215 (N_47215,N_45213,N_45723);
or U47216 (N_47216,N_44528,N_45111);
nor U47217 (N_47217,N_44718,N_45088);
and U47218 (N_47218,N_45048,N_45621);
or U47219 (N_47219,N_45358,N_45751);
and U47220 (N_47220,N_44388,N_45624);
nand U47221 (N_47221,N_45219,N_45525);
or U47222 (N_47222,N_45893,N_45659);
and U47223 (N_47223,N_44345,N_45959);
and U47224 (N_47224,N_44556,N_45282);
xor U47225 (N_47225,N_44957,N_45725);
xor U47226 (N_47226,N_44461,N_44551);
nor U47227 (N_47227,N_45972,N_45660);
nor U47228 (N_47228,N_45846,N_45247);
nand U47229 (N_47229,N_45294,N_44508);
nand U47230 (N_47230,N_45585,N_44469);
xnor U47231 (N_47231,N_45444,N_44330);
nand U47232 (N_47232,N_45326,N_45140);
and U47233 (N_47233,N_44045,N_45522);
or U47234 (N_47234,N_45142,N_45350);
and U47235 (N_47235,N_44878,N_44698);
nand U47236 (N_47236,N_45437,N_45478);
xnor U47237 (N_47237,N_45855,N_44167);
nand U47238 (N_47238,N_45284,N_45649);
nand U47239 (N_47239,N_44808,N_44002);
nand U47240 (N_47240,N_45559,N_45760);
and U47241 (N_47241,N_44919,N_44908);
nand U47242 (N_47242,N_44863,N_45094);
nand U47243 (N_47243,N_45861,N_45385);
or U47244 (N_47244,N_44231,N_45240);
or U47245 (N_47245,N_44609,N_45247);
or U47246 (N_47246,N_44903,N_45308);
nor U47247 (N_47247,N_44246,N_44280);
nor U47248 (N_47248,N_45596,N_44418);
xor U47249 (N_47249,N_44204,N_45824);
xor U47250 (N_47250,N_44657,N_45502);
and U47251 (N_47251,N_45555,N_45387);
or U47252 (N_47252,N_44459,N_44105);
xnor U47253 (N_47253,N_44100,N_44816);
nor U47254 (N_47254,N_45456,N_45896);
or U47255 (N_47255,N_44534,N_44812);
nor U47256 (N_47256,N_45201,N_44303);
or U47257 (N_47257,N_44447,N_44314);
nor U47258 (N_47258,N_45247,N_45181);
nor U47259 (N_47259,N_44677,N_44253);
xnor U47260 (N_47260,N_45989,N_45583);
nor U47261 (N_47261,N_45565,N_45576);
xnor U47262 (N_47262,N_44546,N_44788);
or U47263 (N_47263,N_44968,N_44505);
or U47264 (N_47264,N_44656,N_45353);
and U47265 (N_47265,N_44810,N_44406);
nor U47266 (N_47266,N_44281,N_44008);
nor U47267 (N_47267,N_44549,N_44226);
and U47268 (N_47268,N_45201,N_45821);
or U47269 (N_47269,N_44511,N_45252);
nor U47270 (N_47270,N_44147,N_44597);
xnor U47271 (N_47271,N_45287,N_44339);
nand U47272 (N_47272,N_45919,N_45766);
nor U47273 (N_47273,N_45536,N_44976);
and U47274 (N_47274,N_45160,N_44099);
or U47275 (N_47275,N_45463,N_44381);
or U47276 (N_47276,N_44736,N_45371);
and U47277 (N_47277,N_45761,N_44252);
or U47278 (N_47278,N_45781,N_44605);
or U47279 (N_47279,N_45937,N_45982);
nand U47280 (N_47280,N_44826,N_45656);
nand U47281 (N_47281,N_45202,N_44087);
and U47282 (N_47282,N_44659,N_45570);
or U47283 (N_47283,N_44697,N_44631);
or U47284 (N_47284,N_44314,N_45472);
nand U47285 (N_47285,N_44441,N_44181);
and U47286 (N_47286,N_45545,N_45264);
or U47287 (N_47287,N_44722,N_44417);
or U47288 (N_47288,N_44981,N_44043);
nand U47289 (N_47289,N_45941,N_45876);
or U47290 (N_47290,N_44717,N_45826);
nor U47291 (N_47291,N_45812,N_44737);
and U47292 (N_47292,N_45317,N_44635);
nor U47293 (N_47293,N_44825,N_45121);
nor U47294 (N_47294,N_44705,N_44636);
or U47295 (N_47295,N_44129,N_44381);
or U47296 (N_47296,N_44680,N_45267);
or U47297 (N_47297,N_44329,N_45478);
and U47298 (N_47298,N_44784,N_44802);
nand U47299 (N_47299,N_44225,N_44497);
xnor U47300 (N_47300,N_44223,N_44910);
and U47301 (N_47301,N_44220,N_45891);
xnor U47302 (N_47302,N_44007,N_44902);
nor U47303 (N_47303,N_45859,N_45480);
or U47304 (N_47304,N_45772,N_45897);
xor U47305 (N_47305,N_45819,N_44457);
nand U47306 (N_47306,N_45582,N_44072);
nor U47307 (N_47307,N_45496,N_44349);
nand U47308 (N_47308,N_45220,N_45810);
nor U47309 (N_47309,N_44213,N_44966);
and U47310 (N_47310,N_45250,N_44768);
xor U47311 (N_47311,N_44278,N_44579);
nand U47312 (N_47312,N_44067,N_45659);
and U47313 (N_47313,N_45578,N_44160);
and U47314 (N_47314,N_45313,N_44816);
and U47315 (N_47315,N_44516,N_45886);
and U47316 (N_47316,N_45711,N_44607);
nand U47317 (N_47317,N_45861,N_44862);
or U47318 (N_47318,N_45006,N_45212);
nor U47319 (N_47319,N_45223,N_44542);
nor U47320 (N_47320,N_44552,N_44609);
nand U47321 (N_47321,N_45661,N_45790);
nor U47322 (N_47322,N_45808,N_45702);
nand U47323 (N_47323,N_44598,N_44670);
nand U47324 (N_47324,N_45169,N_44692);
nand U47325 (N_47325,N_44367,N_45313);
or U47326 (N_47326,N_45965,N_44364);
nand U47327 (N_47327,N_45720,N_45784);
nor U47328 (N_47328,N_44446,N_45877);
xnor U47329 (N_47329,N_45151,N_44782);
nand U47330 (N_47330,N_44275,N_44501);
xor U47331 (N_47331,N_44173,N_45340);
or U47332 (N_47332,N_45869,N_45845);
xor U47333 (N_47333,N_44425,N_44635);
xor U47334 (N_47334,N_44966,N_44969);
and U47335 (N_47335,N_44559,N_45078);
and U47336 (N_47336,N_44183,N_45480);
and U47337 (N_47337,N_44939,N_45483);
xnor U47338 (N_47338,N_44392,N_44556);
nand U47339 (N_47339,N_45339,N_45694);
nand U47340 (N_47340,N_44394,N_44211);
and U47341 (N_47341,N_45188,N_45058);
or U47342 (N_47342,N_45113,N_45954);
nand U47343 (N_47343,N_45119,N_45227);
and U47344 (N_47344,N_45609,N_44944);
or U47345 (N_47345,N_44078,N_45805);
or U47346 (N_47346,N_45021,N_45220);
nor U47347 (N_47347,N_45271,N_45822);
nor U47348 (N_47348,N_44533,N_44640);
nor U47349 (N_47349,N_45710,N_45246);
xor U47350 (N_47350,N_45123,N_44651);
and U47351 (N_47351,N_45023,N_45441);
or U47352 (N_47352,N_45476,N_44719);
or U47353 (N_47353,N_45233,N_44489);
xnor U47354 (N_47354,N_44596,N_45678);
nand U47355 (N_47355,N_45232,N_44110);
nand U47356 (N_47356,N_44344,N_44894);
xor U47357 (N_47357,N_44893,N_45104);
or U47358 (N_47358,N_45617,N_45443);
nor U47359 (N_47359,N_44038,N_45740);
and U47360 (N_47360,N_44312,N_45209);
or U47361 (N_47361,N_44715,N_44542);
and U47362 (N_47362,N_44785,N_44632);
nand U47363 (N_47363,N_45529,N_45008);
nand U47364 (N_47364,N_44251,N_45686);
or U47365 (N_47365,N_45974,N_44567);
xnor U47366 (N_47366,N_45010,N_45911);
xnor U47367 (N_47367,N_44470,N_45836);
or U47368 (N_47368,N_44102,N_44671);
xor U47369 (N_47369,N_44861,N_45465);
nand U47370 (N_47370,N_44072,N_45901);
nand U47371 (N_47371,N_45620,N_45384);
and U47372 (N_47372,N_44833,N_45162);
nand U47373 (N_47373,N_45499,N_45011);
xnor U47374 (N_47374,N_45950,N_44475);
nand U47375 (N_47375,N_44953,N_45997);
nor U47376 (N_47376,N_45660,N_44444);
nand U47377 (N_47377,N_44894,N_45369);
nand U47378 (N_47378,N_45276,N_45105);
nand U47379 (N_47379,N_45319,N_44207);
or U47380 (N_47380,N_44982,N_44727);
xor U47381 (N_47381,N_44335,N_44892);
xnor U47382 (N_47382,N_45273,N_44535);
nand U47383 (N_47383,N_45644,N_44212);
nand U47384 (N_47384,N_44373,N_45518);
or U47385 (N_47385,N_44505,N_44830);
or U47386 (N_47386,N_45766,N_44018);
or U47387 (N_47387,N_45730,N_45832);
or U47388 (N_47388,N_45620,N_45396);
xnor U47389 (N_47389,N_45226,N_45380);
nor U47390 (N_47390,N_44544,N_45171);
nand U47391 (N_47391,N_45645,N_44461);
or U47392 (N_47392,N_44928,N_45636);
nor U47393 (N_47393,N_44584,N_44840);
and U47394 (N_47394,N_45841,N_44514);
or U47395 (N_47395,N_44890,N_44689);
and U47396 (N_47396,N_45298,N_44228);
nand U47397 (N_47397,N_44364,N_44702);
or U47398 (N_47398,N_44165,N_45223);
nor U47399 (N_47399,N_45035,N_45776);
xnor U47400 (N_47400,N_45635,N_44551);
nor U47401 (N_47401,N_44522,N_44921);
nor U47402 (N_47402,N_45452,N_45775);
and U47403 (N_47403,N_44170,N_44468);
nor U47404 (N_47404,N_44772,N_45211);
or U47405 (N_47405,N_44131,N_44366);
nor U47406 (N_47406,N_44428,N_45979);
nand U47407 (N_47407,N_45637,N_44965);
and U47408 (N_47408,N_45278,N_44093);
nor U47409 (N_47409,N_44098,N_44460);
nand U47410 (N_47410,N_44102,N_45749);
nand U47411 (N_47411,N_44967,N_44662);
nand U47412 (N_47412,N_44934,N_44640);
nor U47413 (N_47413,N_45071,N_45683);
nand U47414 (N_47414,N_45915,N_45246);
and U47415 (N_47415,N_45959,N_44550);
nand U47416 (N_47416,N_45149,N_44824);
and U47417 (N_47417,N_44327,N_45846);
or U47418 (N_47418,N_44199,N_44620);
nand U47419 (N_47419,N_44932,N_45313);
nor U47420 (N_47420,N_44839,N_45179);
xor U47421 (N_47421,N_45772,N_45052);
or U47422 (N_47422,N_45250,N_44903);
nand U47423 (N_47423,N_44206,N_44634);
and U47424 (N_47424,N_44799,N_44899);
nor U47425 (N_47425,N_45990,N_45600);
and U47426 (N_47426,N_45735,N_44211);
and U47427 (N_47427,N_44449,N_44677);
nand U47428 (N_47428,N_44169,N_45872);
or U47429 (N_47429,N_44698,N_44279);
nand U47430 (N_47430,N_44052,N_45740);
nand U47431 (N_47431,N_45484,N_44029);
and U47432 (N_47432,N_45521,N_45991);
xnor U47433 (N_47433,N_44671,N_45885);
and U47434 (N_47434,N_45318,N_44197);
nor U47435 (N_47435,N_45706,N_45877);
nand U47436 (N_47436,N_44615,N_44435);
nand U47437 (N_47437,N_45586,N_44236);
and U47438 (N_47438,N_45013,N_45019);
nand U47439 (N_47439,N_44241,N_45833);
nor U47440 (N_47440,N_44927,N_45868);
nor U47441 (N_47441,N_45552,N_45915);
nor U47442 (N_47442,N_44539,N_44572);
nand U47443 (N_47443,N_44647,N_45689);
and U47444 (N_47444,N_45305,N_45371);
nand U47445 (N_47445,N_45357,N_45931);
xor U47446 (N_47446,N_44862,N_44132);
xor U47447 (N_47447,N_44748,N_45968);
xor U47448 (N_47448,N_45070,N_44148);
or U47449 (N_47449,N_44514,N_44115);
xnor U47450 (N_47450,N_44933,N_44765);
nor U47451 (N_47451,N_45534,N_44132);
nand U47452 (N_47452,N_45376,N_45087);
and U47453 (N_47453,N_44207,N_45705);
or U47454 (N_47454,N_44185,N_44622);
and U47455 (N_47455,N_45717,N_45836);
and U47456 (N_47456,N_44505,N_44840);
xnor U47457 (N_47457,N_45867,N_44750);
xnor U47458 (N_47458,N_44533,N_45072);
xor U47459 (N_47459,N_45439,N_44381);
nand U47460 (N_47460,N_45197,N_45064);
nor U47461 (N_47461,N_45727,N_45462);
and U47462 (N_47462,N_44143,N_44552);
nor U47463 (N_47463,N_45598,N_45421);
and U47464 (N_47464,N_44385,N_44470);
or U47465 (N_47465,N_44126,N_45218);
nor U47466 (N_47466,N_44458,N_44633);
xnor U47467 (N_47467,N_44334,N_45807);
nor U47468 (N_47468,N_45857,N_44787);
or U47469 (N_47469,N_45437,N_45762);
nand U47470 (N_47470,N_45389,N_44457);
nor U47471 (N_47471,N_44815,N_44990);
nand U47472 (N_47472,N_44736,N_45127);
or U47473 (N_47473,N_45494,N_44711);
and U47474 (N_47474,N_45140,N_44239);
or U47475 (N_47475,N_44952,N_44363);
nor U47476 (N_47476,N_44345,N_44352);
nand U47477 (N_47477,N_45768,N_45866);
and U47478 (N_47478,N_45248,N_45875);
xnor U47479 (N_47479,N_44347,N_44288);
nand U47480 (N_47480,N_45065,N_45894);
nand U47481 (N_47481,N_44734,N_45138);
nand U47482 (N_47482,N_44467,N_44361);
or U47483 (N_47483,N_44768,N_44763);
nor U47484 (N_47484,N_44613,N_44618);
or U47485 (N_47485,N_44304,N_45727);
nand U47486 (N_47486,N_44791,N_44952);
and U47487 (N_47487,N_45221,N_45063);
and U47488 (N_47488,N_45409,N_44856);
and U47489 (N_47489,N_44135,N_45712);
or U47490 (N_47490,N_44535,N_44300);
nor U47491 (N_47491,N_45778,N_45811);
nor U47492 (N_47492,N_44890,N_45525);
and U47493 (N_47493,N_45865,N_44744);
or U47494 (N_47494,N_45538,N_45450);
or U47495 (N_47495,N_45628,N_45792);
xor U47496 (N_47496,N_44124,N_45328);
nor U47497 (N_47497,N_45980,N_45868);
xnor U47498 (N_47498,N_45660,N_45393);
nand U47499 (N_47499,N_44486,N_45411);
and U47500 (N_47500,N_45372,N_44133);
nand U47501 (N_47501,N_44689,N_44058);
nand U47502 (N_47502,N_44354,N_45294);
xor U47503 (N_47503,N_45731,N_45143);
nor U47504 (N_47504,N_44143,N_44301);
and U47505 (N_47505,N_45884,N_44935);
nor U47506 (N_47506,N_44612,N_45046);
and U47507 (N_47507,N_44045,N_45376);
and U47508 (N_47508,N_44059,N_45196);
and U47509 (N_47509,N_45835,N_45049);
xor U47510 (N_47510,N_44830,N_45054);
and U47511 (N_47511,N_45254,N_45480);
nand U47512 (N_47512,N_45873,N_45707);
nand U47513 (N_47513,N_44935,N_45194);
or U47514 (N_47514,N_45166,N_44641);
nand U47515 (N_47515,N_44077,N_44245);
and U47516 (N_47516,N_44360,N_44876);
nand U47517 (N_47517,N_45894,N_44456);
xor U47518 (N_47518,N_45146,N_44486);
xor U47519 (N_47519,N_45301,N_45321);
nand U47520 (N_47520,N_45967,N_44286);
xnor U47521 (N_47521,N_44937,N_44999);
nor U47522 (N_47522,N_45552,N_44266);
nand U47523 (N_47523,N_45362,N_45768);
nand U47524 (N_47524,N_45492,N_44672);
or U47525 (N_47525,N_45936,N_44439);
or U47526 (N_47526,N_44372,N_45110);
nand U47527 (N_47527,N_44225,N_45668);
or U47528 (N_47528,N_44000,N_45158);
or U47529 (N_47529,N_44634,N_44808);
xnor U47530 (N_47530,N_44548,N_45809);
nor U47531 (N_47531,N_45864,N_45225);
nand U47532 (N_47532,N_45694,N_44654);
nand U47533 (N_47533,N_44275,N_45848);
nor U47534 (N_47534,N_44479,N_44199);
and U47535 (N_47535,N_44641,N_45192);
and U47536 (N_47536,N_45660,N_45533);
and U47537 (N_47537,N_45201,N_45188);
nor U47538 (N_47538,N_45900,N_45327);
and U47539 (N_47539,N_45877,N_45615);
or U47540 (N_47540,N_44103,N_44436);
xor U47541 (N_47541,N_45926,N_44254);
nor U47542 (N_47542,N_44735,N_44995);
xor U47543 (N_47543,N_44903,N_44736);
or U47544 (N_47544,N_44954,N_44448);
nor U47545 (N_47545,N_45506,N_44168);
xnor U47546 (N_47546,N_45457,N_45181);
xor U47547 (N_47547,N_45118,N_45923);
and U47548 (N_47548,N_44143,N_44665);
nand U47549 (N_47549,N_45413,N_44045);
nand U47550 (N_47550,N_45409,N_44539);
and U47551 (N_47551,N_44063,N_44540);
nand U47552 (N_47552,N_45959,N_44605);
or U47553 (N_47553,N_44154,N_45669);
xnor U47554 (N_47554,N_44011,N_44117);
or U47555 (N_47555,N_45935,N_45988);
nand U47556 (N_47556,N_45319,N_44944);
nand U47557 (N_47557,N_45177,N_44535);
xor U47558 (N_47558,N_45900,N_44511);
nor U47559 (N_47559,N_45042,N_45292);
and U47560 (N_47560,N_44514,N_44051);
and U47561 (N_47561,N_45713,N_45560);
nand U47562 (N_47562,N_44495,N_45571);
nand U47563 (N_47563,N_44112,N_44692);
or U47564 (N_47564,N_45677,N_44276);
nand U47565 (N_47565,N_44248,N_44969);
xnor U47566 (N_47566,N_44826,N_45635);
and U47567 (N_47567,N_44110,N_44184);
nor U47568 (N_47568,N_45540,N_45875);
nand U47569 (N_47569,N_44391,N_45819);
nand U47570 (N_47570,N_44897,N_45399);
and U47571 (N_47571,N_45442,N_44760);
nand U47572 (N_47572,N_44934,N_44262);
and U47573 (N_47573,N_44052,N_44010);
nand U47574 (N_47574,N_45363,N_45767);
or U47575 (N_47575,N_45222,N_44245);
and U47576 (N_47576,N_45095,N_44284);
nand U47577 (N_47577,N_44511,N_44704);
nand U47578 (N_47578,N_44140,N_45979);
nor U47579 (N_47579,N_44226,N_45485);
and U47580 (N_47580,N_45336,N_44794);
nand U47581 (N_47581,N_44479,N_45402);
and U47582 (N_47582,N_45945,N_45201);
and U47583 (N_47583,N_44951,N_45690);
nor U47584 (N_47584,N_44266,N_44593);
xor U47585 (N_47585,N_45260,N_45646);
nand U47586 (N_47586,N_44325,N_44899);
nor U47587 (N_47587,N_45293,N_45835);
or U47588 (N_47588,N_45818,N_45738);
xnor U47589 (N_47589,N_44635,N_45992);
or U47590 (N_47590,N_45554,N_44562);
and U47591 (N_47591,N_44690,N_45935);
xnor U47592 (N_47592,N_45120,N_44132);
nand U47593 (N_47593,N_45595,N_44010);
or U47594 (N_47594,N_45142,N_44581);
nand U47595 (N_47595,N_45328,N_44822);
xnor U47596 (N_47596,N_45686,N_45282);
nand U47597 (N_47597,N_45649,N_44012);
or U47598 (N_47598,N_44053,N_45588);
or U47599 (N_47599,N_44800,N_45377);
xor U47600 (N_47600,N_45682,N_45871);
nand U47601 (N_47601,N_45025,N_45636);
or U47602 (N_47602,N_44699,N_45702);
or U47603 (N_47603,N_45899,N_44512);
xor U47604 (N_47604,N_45847,N_44759);
and U47605 (N_47605,N_44961,N_44279);
nand U47606 (N_47606,N_45568,N_45919);
xnor U47607 (N_47607,N_45850,N_44561);
nor U47608 (N_47608,N_44908,N_45910);
or U47609 (N_47609,N_44631,N_45149);
or U47610 (N_47610,N_45063,N_44649);
and U47611 (N_47611,N_44268,N_45678);
xnor U47612 (N_47612,N_44793,N_45364);
nor U47613 (N_47613,N_44684,N_44481);
nand U47614 (N_47614,N_44831,N_44151);
and U47615 (N_47615,N_45041,N_44215);
or U47616 (N_47616,N_44771,N_44839);
nand U47617 (N_47617,N_44029,N_45278);
nor U47618 (N_47618,N_44584,N_45154);
and U47619 (N_47619,N_45329,N_45938);
nand U47620 (N_47620,N_44574,N_45505);
or U47621 (N_47621,N_45626,N_44697);
or U47622 (N_47622,N_44227,N_45254);
nor U47623 (N_47623,N_45814,N_45940);
or U47624 (N_47624,N_44789,N_44546);
nand U47625 (N_47625,N_45255,N_45368);
and U47626 (N_47626,N_45113,N_45984);
nor U47627 (N_47627,N_45944,N_45853);
and U47628 (N_47628,N_44326,N_45553);
and U47629 (N_47629,N_44736,N_45066);
and U47630 (N_47630,N_45554,N_44487);
nand U47631 (N_47631,N_45127,N_45409);
and U47632 (N_47632,N_44277,N_44096);
xor U47633 (N_47633,N_44879,N_45028);
xor U47634 (N_47634,N_45816,N_45833);
and U47635 (N_47635,N_45513,N_45533);
and U47636 (N_47636,N_45165,N_44511);
xor U47637 (N_47637,N_45391,N_44537);
nor U47638 (N_47638,N_44061,N_44320);
nor U47639 (N_47639,N_45180,N_44669);
nand U47640 (N_47640,N_44952,N_45281);
xor U47641 (N_47641,N_45103,N_44829);
or U47642 (N_47642,N_44647,N_45911);
nor U47643 (N_47643,N_45107,N_44182);
xor U47644 (N_47644,N_44720,N_44724);
nor U47645 (N_47645,N_45224,N_45242);
nand U47646 (N_47646,N_44705,N_44288);
or U47647 (N_47647,N_44147,N_45174);
xor U47648 (N_47648,N_44402,N_44498);
nor U47649 (N_47649,N_44102,N_44940);
nor U47650 (N_47650,N_45623,N_45251);
nand U47651 (N_47651,N_44500,N_44356);
xnor U47652 (N_47652,N_45113,N_45841);
or U47653 (N_47653,N_45197,N_44189);
and U47654 (N_47654,N_45326,N_45885);
xnor U47655 (N_47655,N_44047,N_44583);
and U47656 (N_47656,N_44747,N_45183);
and U47657 (N_47657,N_45234,N_44153);
and U47658 (N_47658,N_45427,N_44580);
xnor U47659 (N_47659,N_44741,N_44456);
nand U47660 (N_47660,N_44808,N_44035);
nand U47661 (N_47661,N_45150,N_45042);
and U47662 (N_47662,N_44418,N_45653);
or U47663 (N_47663,N_45030,N_45228);
or U47664 (N_47664,N_44190,N_44751);
and U47665 (N_47665,N_44797,N_45971);
and U47666 (N_47666,N_44635,N_44212);
nor U47667 (N_47667,N_44568,N_44502);
nand U47668 (N_47668,N_45565,N_44242);
or U47669 (N_47669,N_44489,N_44920);
xnor U47670 (N_47670,N_45238,N_44137);
nor U47671 (N_47671,N_44384,N_45039);
nand U47672 (N_47672,N_45831,N_44134);
or U47673 (N_47673,N_45759,N_45777);
nand U47674 (N_47674,N_45316,N_45643);
and U47675 (N_47675,N_45776,N_44756);
xor U47676 (N_47676,N_45038,N_44320);
and U47677 (N_47677,N_44625,N_44236);
and U47678 (N_47678,N_44323,N_45551);
nand U47679 (N_47679,N_45310,N_44211);
nand U47680 (N_47680,N_44540,N_45397);
xor U47681 (N_47681,N_44615,N_44077);
and U47682 (N_47682,N_45778,N_45976);
and U47683 (N_47683,N_45311,N_44338);
or U47684 (N_47684,N_45608,N_44318);
xnor U47685 (N_47685,N_45934,N_45367);
and U47686 (N_47686,N_44967,N_44113);
nor U47687 (N_47687,N_45898,N_45214);
or U47688 (N_47688,N_45855,N_45075);
nor U47689 (N_47689,N_44218,N_44744);
or U47690 (N_47690,N_44009,N_44184);
or U47691 (N_47691,N_45904,N_44668);
nor U47692 (N_47692,N_44378,N_45717);
xnor U47693 (N_47693,N_44840,N_44837);
nand U47694 (N_47694,N_45906,N_45422);
nor U47695 (N_47695,N_45297,N_44612);
nor U47696 (N_47696,N_44341,N_45063);
and U47697 (N_47697,N_44149,N_44798);
or U47698 (N_47698,N_44198,N_45866);
or U47699 (N_47699,N_45437,N_45232);
nand U47700 (N_47700,N_44821,N_44902);
xor U47701 (N_47701,N_44418,N_44123);
xnor U47702 (N_47702,N_44423,N_44002);
or U47703 (N_47703,N_45343,N_45441);
or U47704 (N_47704,N_44269,N_44867);
nor U47705 (N_47705,N_44599,N_44552);
and U47706 (N_47706,N_44120,N_45591);
and U47707 (N_47707,N_45216,N_44369);
or U47708 (N_47708,N_45478,N_45837);
and U47709 (N_47709,N_45945,N_45121);
nor U47710 (N_47710,N_44460,N_44100);
or U47711 (N_47711,N_45368,N_45985);
nand U47712 (N_47712,N_45517,N_45819);
or U47713 (N_47713,N_45258,N_44439);
nor U47714 (N_47714,N_44975,N_45018);
nor U47715 (N_47715,N_44233,N_44311);
xnor U47716 (N_47716,N_45665,N_44728);
or U47717 (N_47717,N_44446,N_44126);
xnor U47718 (N_47718,N_45326,N_44284);
nand U47719 (N_47719,N_44317,N_44734);
and U47720 (N_47720,N_44402,N_44755);
nor U47721 (N_47721,N_45547,N_45620);
xnor U47722 (N_47722,N_45390,N_45776);
nor U47723 (N_47723,N_44542,N_45832);
and U47724 (N_47724,N_45065,N_45603);
or U47725 (N_47725,N_44966,N_44788);
and U47726 (N_47726,N_45746,N_45940);
nor U47727 (N_47727,N_45627,N_45623);
nand U47728 (N_47728,N_45391,N_44839);
nand U47729 (N_47729,N_45064,N_45791);
nor U47730 (N_47730,N_44159,N_44313);
nor U47731 (N_47731,N_44405,N_44887);
xnor U47732 (N_47732,N_44195,N_44776);
nand U47733 (N_47733,N_44110,N_44585);
nor U47734 (N_47734,N_44399,N_44378);
xor U47735 (N_47735,N_44338,N_44172);
nor U47736 (N_47736,N_45350,N_44634);
nor U47737 (N_47737,N_44201,N_45627);
xor U47738 (N_47738,N_45017,N_44888);
and U47739 (N_47739,N_45249,N_45466);
xor U47740 (N_47740,N_45231,N_45500);
nor U47741 (N_47741,N_45408,N_45526);
nand U47742 (N_47742,N_45873,N_45000);
xor U47743 (N_47743,N_44429,N_45780);
and U47744 (N_47744,N_44829,N_44452);
nand U47745 (N_47745,N_45270,N_44522);
nor U47746 (N_47746,N_45971,N_44265);
nand U47747 (N_47747,N_45932,N_44610);
or U47748 (N_47748,N_44697,N_45612);
xnor U47749 (N_47749,N_44514,N_44227);
nand U47750 (N_47750,N_45757,N_45406);
xnor U47751 (N_47751,N_45097,N_44561);
xnor U47752 (N_47752,N_45438,N_44344);
or U47753 (N_47753,N_45326,N_45739);
and U47754 (N_47754,N_45790,N_44563);
and U47755 (N_47755,N_45531,N_44042);
nand U47756 (N_47756,N_44629,N_45794);
nor U47757 (N_47757,N_45991,N_45427);
nand U47758 (N_47758,N_45995,N_45344);
xor U47759 (N_47759,N_44618,N_44413);
and U47760 (N_47760,N_45518,N_45191);
nand U47761 (N_47761,N_44676,N_44164);
nor U47762 (N_47762,N_45482,N_45144);
nand U47763 (N_47763,N_44993,N_44454);
or U47764 (N_47764,N_45387,N_45524);
xnor U47765 (N_47765,N_44519,N_45769);
nor U47766 (N_47766,N_44997,N_44529);
and U47767 (N_47767,N_45663,N_45275);
xnor U47768 (N_47768,N_45087,N_45451);
or U47769 (N_47769,N_44965,N_44095);
xnor U47770 (N_47770,N_45117,N_44079);
nor U47771 (N_47771,N_44816,N_44410);
and U47772 (N_47772,N_45316,N_44225);
or U47773 (N_47773,N_45962,N_45097);
nand U47774 (N_47774,N_45751,N_44041);
or U47775 (N_47775,N_45544,N_45844);
or U47776 (N_47776,N_44089,N_44364);
nor U47777 (N_47777,N_44203,N_44813);
and U47778 (N_47778,N_45449,N_44353);
or U47779 (N_47779,N_44794,N_44759);
xor U47780 (N_47780,N_45489,N_44043);
and U47781 (N_47781,N_45071,N_44862);
nor U47782 (N_47782,N_44577,N_44612);
or U47783 (N_47783,N_45081,N_44487);
or U47784 (N_47784,N_45609,N_44642);
nand U47785 (N_47785,N_44914,N_45443);
nand U47786 (N_47786,N_44194,N_44917);
nor U47787 (N_47787,N_45588,N_45142);
xor U47788 (N_47788,N_45216,N_45041);
nand U47789 (N_47789,N_44475,N_44713);
and U47790 (N_47790,N_44400,N_45279);
or U47791 (N_47791,N_44634,N_44285);
and U47792 (N_47792,N_45137,N_44902);
nor U47793 (N_47793,N_44213,N_45350);
xnor U47794 (N_47794,N_44829,N_45058);
nor U47795 (N_47795,N_45884,N_45837);
and U47796 (N_47796,N_44865,N_45502);
nor U47797 (N_47797,N_44923,N_44499);
or U47798 (N_47798,N_45711,N_45266);
nand U47799 (N_47799,N_44201,N_45229);
or U47800 (N_47800,N_45384,N_44129);
nor U47801 (N_47801,N_44637,N_45922);
or U47802 (N_47802,N_45465,N_45661);
and U47803 (N_47803,N_44860,N_44912);
nor U47804 (N_47804,N_44438,N_45575);
nor U47805 (N_47805,N_45984,N_45730);
nand U47806 (N_47806,N_44346,N_45319);
and U47807 (N_47807,N_44332,N_45248);
xor U47808 (N_47808,N_44887,N_45280);
or U47809 (N_47809,N_45756,N_45774);
or U47810 (N_47810,N_44260,N_44120);
and U47811 (N_47811,N_45847,N_45939);
nand U47812 (N_47812,N_45956,N_44669);
nor U47813 (N_47813,N_45219,N_45514);
nand U47814 (N_47814,N_45785,N_45788);
and U47815 (N_47815,N_44453,N_44324);
xor U47816 (N_47816,N_44219,N_44407);
or U47817 (N_47817,N_45317,N_45560);
or U47818 (N_47818,N_44203,N_45470);
nand U47819 (N_47819,N_44274,N_45956);
xor U47820 (N_47820,N_44721,N_44681);
nand U47821 (N_47821,N_45632,N_44666);
nor U47822 (N_47822,N_44181,N_45138);
nor U47823 (N_47823,N_44029,N_45343);
or U47824 (N_47824,N_45026,N_45726);
nor U47825 (N_47825,N_44687,N_45462);
or U47826 (N_47826,N_44701,N_45057);
nand U47827 (N_47827,N_45376,N_45586);
and U47828 (N_47828,N_45505,N_44171);
xnor U47829 (N_47829,N_45035,N_44549);
and U47830 (N_47830,N_44871,N_45223);
and U47831 (N_47831,N_44025,N_44872);
and U47832 (N_47832,N_44207,N_44843);
nor U47833 (N_47833,N_45963,N_45732);
nor U47834 (N_47834,N_45316,N_44026);
or U47835 (N_47835,N_44336,N_44315);
and U47836 (N_47836,N_44918,N_45501);
nand U47837 (N_47837,N_45255,N_45743);
and U47838 (N_47838,N_44652,N_45796);
nor U47839 (N_47839,N_45164,N_44668);
xor U47840 (N_47840,N_44518,N_44614);
nand U47841 (N_47841,N_44790,N_45611);
and U47842 (N_47842,N_44531,N_45090);
nor U47843 (N_47843,N_44495,N_44665);
or U47844 (N_47844,N_44930,N_45127);
nor U47845 (N_47845,N_44476,N_45623);
or U47846 (N_47846,N_45136,N_44536);
nor U47847 (N_47847,N_45723,N_44940);
nor U47848 (N_47848,N_45267,N_44521);
xor U47849 (N_47849,N_44419,N_44224);
nor U47850 (N_47850,N_45051,N_44789);
and U47851 (N_47851,N_45932,N_45846);
nand U47852 (N_47852,N_45091,N_44489);
nor U47853 (N_47853,N_45732,N_44279);
xnor U47854 (N_47854,N_44748,N_45742);
nor U47855 (N_47855,N_44801,N_44513);
and U47856 (N_47856,N_45827,N_44296);
nand U47857 (N_47857,N_44884,N_44759);
xnor U47858 (N_47858,N_45985,N_45475);
and U47859 (N_47859,N_45929,N_44024);
nor U47860 (N_47860,N_44363,N_44589);
nor U47861 (N_47861,N_44171,N_44746);
nand U47862 (N_47862,N_45635,N_44907);
and U47863 (N_47863,N_45342,N_45138);
and U47864 (N_47864,N_45089,N_44985);
or U47865 (N_47865,N_44528,N_44759);
and U47866 (N_47866,N_45457,N_44852);
nor U47867 (N_47867,N_45949,N_45364);
nand U47868 (N_47868,N_44656,N_44710);
or U47869 (N_47869,N_45240,N_45170);
xor U47870 (N_47870,N_44842,N_44571);
or U47871 (N_47871,N_45003,N_44139);
xor U47872 (N_47872,N_44514,N_45650);
or U47873 (N_47873,N_44846,N_44686);
or U47874 (N_47874,N_44530,N_45203);
nor U47875 (N_47875,N_44858,N_44733);
xnor U47876 (N_47876,N_45612,N_45107);
or U47877 (N_47877,N_44786,N_45197);
nor U47878 (N_47878,N_45554,N_45938);
nand U47879 (N_47879,N_44370,N_45623);
and U47880 (N_47880,N_44780,N_45063);
and U47881 (N_47881,N_45873,N_44239);
and U47882 (N_47882,N_45421,N_44948);
xnor U47883 (N_47883,N_45310,N_45771);
nand U47884 (N_47884,N_44077,N_45663);
nor U47885 (N_47885,N_44965,N_45647);
nor U47886 (N_47886,N_45265,N_44168);
or U47887 (N_47887,N_44788,N_44125);
or U47888 (N_47888,N_44784,N_44670);
and U47889 (N_47889,N_44003,N_44229);
and U47890 (N_47890,N_45718,N_44684);
xor U47891 (N_47891,N_44636,N_44318);
and U47892 (N_47892,N_44883,N_44228);
nand U47893 (N_47893,N_44968,N_44021);
nor U47894 (N_47894,N_44028,N_45697);
xor U47895 (N_47895,N_44549,N_44572);
or U47896 (N_47896,N_44982,N_45377);
nor U47897 (N_47897,N_44821,N_45424);
nor U47898 (N_47898,N_45296,N_45237);
or U47899 (N_47899,N_45715,N_45847);
xnor U47900 (N_47900,N_44094,N_45127);
xnor U47901 (N_47901,N_45799,N_44489);
nand U47902 (N_47902,N_44362,N_44771);
xnor U47903 (N_47903,N_45844,N_45809);
or U47904 (N_47904,N_45937,N_44853);
and U47905 (N_47905,N_45284,N_44094);
xor U47906 (N_47906,N_44266,N_44493);
nand U47907 (N_47907,N_45045,N_45248);
nand U47908 (N_47908,N_44193,N_45521);
or U47909 (N_47909,N_44087,N_45843);
and U47910 (N_47910,N_45675,N_45781);
and U47911 (N_47911,N_45024,N_44669);
or U47912 (N_47912,N_44830,N_45657);
and U47913 (N_47913,N_45679,N_45300);
nand U47914 (N_47914,N_45117,N_44148);
xnor U47915 (N_47915,N_44385,N_44959);
nor U47916 (N_47916,N_44580,N_45970);
nand U47917 (N_47917,N_44800,N_44563);
or U47918 (N_47918,N_44369,N_44624);
or U47919 (N_47919,N_45212,N_44343);
nor U47920 (N_47920,N_44790,N_45892);
and U47921 (N_47921,N_44019,N_44118);
and U47922 (N_47922,N_44309,N_44063);
xor U47923 (N_47923,N_44443,N_45596);
xor U47924 (N_47924,N_44127,N_44985);
xor U47925 (N_47925,N_44292,N_44606);
or U47926 (N_47926,N_45819,N_44091);
or U47927 (N_47927,N_44237,N_45837);
nand U47928 (N_47928,N_45444,N_45003);
nor U47929 (N_47929,N_45172,N_44461);
and U47930 (N_47930,N_44781,N_45354);
nand U47931 (N_47931,N_44320,N_44183);
nand U47932 (N_47932,N_44349,N_45242);
and U47933 (N_47933,N_45027,N_45342);
nor U47934 (N_47934,N_45149,N_44470);
xor U47935 (N_47935,N_45653,N_45264);
nand U47936 (N_47936,N_44460,N_44010);
or U47937 (N_47937,N_44525,N_44033);
xor U47938 (N_47938,N_45555,N_45452);
nand U47939 (N_47939,N_45866,N_45009);
and U47940 (N_47940,N_44180,N_44994);
and U47941 (N_47941,N_44633,N_45109);
nor U47942 (N_47942,N_45097,N_44290);
or U47943 (N_47943,N_44704,N_45089);
nor U47944 (N_47944,N_45569,N_45816);
or U47945 (N_47945,N_44301,N_45914);
xnor U47946 (N_47946,N_45797,N_45264);
and U47947 (N_47947,N_44664,N_45433);
and U47948 (N_47948,N_44284,N_45130);
or U47949 (N_47949,N_44174,N_44293);
or U47950 (N_47950,N_44344,N_45628);
nand U47951 (N_47951,N_44513,N_45002);
or U47952 (N_47952,N_45020,N_45410);
nand U47953 (N_47953,N_44030,N_44422);
and U47954 (N_47954,N_45001,N_44394);
and U47955 (N_47955,N_45510,N_45040);
or U47956 (N_47956,N_44323,N_44738);
and U47957 (N_47957,N_45478,N_44603);
xnor U47958 (N_47958,N_44011,N_44366);
or U47959 (N_47959,N_45402,N_45061);
nor U47960 (N_47960,N_44949,N_45973);
nor U47961 (N_47961,N_44153,N_45902);
nor U47962 (N_47962,N_45793,N_45380);
nor U47963 (N_47963,N_45587,N_45720);
xnor U47964 (N_47964,N_45945,N_44859);
nor U47965 (N_47965,N_44843,N_45979);
and U47966 (N_47966,N_44954,N_45366);
nor U47967 (N_47967,N_44367,N_44812);
nand U47968 (N_47968,N_44682,N_44947);
and U47969 (N_47969,N_45225,N_45459);
or U47970 (N_47970,N_45326,N_45978);
nand U47971 (N_47971,N_45686,N_44346);
or U47972 (N_47972,N_44143,N_44881);
and U47973 (N_47973,N_45930,N_45854);
xnor U47974 (N_47974,N_45931,N_44634);
nand U47975 (N_47975,N_44219,N_45849);
and U47976 (N_47976,N_44884,N_45997);
and U47977 (N_47977,N_44622,N_45728);
and U47978 (N_47978,N_44955,N_45404);
xor U47979 (N_47979,N_45768,N_45360);
or U47980 (N_47980,N_45696,N_45553);
and U47981 (N_47981,N_44733,N_44985);
xor U47982 (N_47982,N_44599,N_45936);
nand U47983 (N_47983,N_45805,N_44870);
or U47984 (N_47984,N_45107,N_44189);
xor U47985 (N_47985,N_45457,N_44084);
nand U47986 (N_47986,N_44963,N_45189);
and U47987 (N_47987,N_44712,N_44215);
nand U47988 (N_47988,N_45570,N_45945);
xor U47989 (N_47989,N_45475,N_45598);
xnor U47990 (N_47990,N_45618,N_44766);
and U47991 (N_47991,N_45122,N_44040);
or U47992 (N_47992,N_44075,N_45685);
nor U47993 (N_47993,N_45268,N_45607);
xnor U47994 (N_47994,N_45202,N_44661);
nand U47995 (N_47995,N_45115,N_45941);
and U47996 (N_47996,N_45455,N_44565);
xor U47997 (N_47997,N_44794,N_44626);
or U47998 (N_47998,N_45797,N_44927);
xnor U47999 (N_47999,N_44338,N_44904);
xnor U48000 (N_48000,N_47919,N_46135);
or U48001 (N_48001,N_47833,N_47343);
nand U48002 (N_48002,N_46531,N_46198);
nor U48003 (N_48003,N_47757,N_46015);
xor U48004 (N_48004,N_46069,N_47299);
nor U48005 (N_48005,N_46151,N_46967);
nand U48006 (N_48006,N_46991,N_47674);
nor U48007 (N_48007,N_47787,N_46109);
nor U48008 (N_48008,N_47776,N_46825);
nor U48009 (N_48009,N_47871,N_47835);
nor U48010 (N_48010,N_46017,N_47305);
nor U48011 (N_48011,N_47275,N_46316);
xor U48012 (N_48012,N_47592,N_46053);
nand U48013 (N_48013,N_46243,N_46369);
xnor U48014 (N_48014,N_46468,N_47785);
or U48015 (N_48015,N_46735,N_47556);
nor U48016 (N_48016,N_46363,N_47762);
or U48017 (N_48017,N_46122,N_47620);
nor U48018 (N_48018,N_46663,N_46617);
nand U48019 (N_48019,N_47035,N_47547);
nand U48020 (N_48020,N_47790,N_47499);
nand U48021 (N_48021,N_47064,N_46219);
xnor U48022 (N_48022,N_46434,N_46562);
or U48023 (N_48023,N_47791,N_46733);
nor U48024 (N_48024,N_47622,N_47680);
xnor U48025 (N_48025,N_46577,N_46235);
nor U48026 (N_48026,N_47151,N_46538);
or U48027 (N_48027,N_47312,N_46454);
and U48028 (N_48028,N_47117,N_47624);
nand U48029 (N_48029,N_46585,N_47551);
and U48030 (N_48030,N_46910,N_47068);
or U48031 (N_48031,N_46848,N_47682);
nor U48032 (N_48032,N_46838,N_46817);
and U48033 (N_48033,N_47948,N_47500);
nand U48034 (N_48034,N_46082,N_47361);
xor U48035 (N_48035,N_47257,N_47975);
xnor U48036 (N_48036,N_47079,N_46270);
nor U48037 (N_48037,N_47375,N_46321);
nand U48038 (N_48038,N_47213,N_47742);
or U48039 (N_48039,N_46982,N_46252);
and U48040 (N_48040,N_47492,N_46775);
xor U48041 (N_48041,N_46561,N_47171);
nor U48042 (N_48042,N_46798,N_47600);
xnor U48043 (N_48043,N_46615,N_46089);
or U48044 (N_48044,N_47471,N_46856);
or U48045 (N_48045,N_47777,N_46756);
and U48046 (N_48046,N_47850,N_46556);
and U48047 (N_48047,N_46546,N_46867);
nand U48048 (N_48048,N_46949,N_46224);
xor U48049 (N_48049,N_47251,N_47432);
xor U48050 (N_48050,N_47408,N_47739);
or U48051 (N_48051,N_47502,N_46380);
xnor U48052 (N_48052,N_47057,N_46984);
and U48053 (N_48053,N_47889,N_46841);
or U48054 (N_48054,N_47255,N_47411);
xnor U48055 (N_48055,N_46569,N_47761);
xor U48056 (N_48056,N_46085,N_46463);
xnor U48057 (N_48057,N_46778,N_47144);
or U48058 (N_48058,N_46277,N_46532);
xor U48059 (N_48059,N_47961,N_47883);
nand U48060 (N_48060,N_47763,N_47067);
or U48061 (N_48061,N_46586,N_46939);
nor U48062 (N_48062,N_46943,N_47435);
and U48063 (N_48063,N_46707,N_47759);
xnor U48064 (N_48064,N_46891,N_46671);
nand U48065 (N_48065,N_46533,N_47808);
nand U48066 (N_48066,N_47594,N_46888);
nand U48067 (N_48067,N_47350,N_47369);
nand U48068 (N_48068,N_46377,N_47216);
or U48069 (N_48069,N_47112,N_47076);
or U48070 (N_48070,N_47641,N_46427);
nand U48071 (N_48071,N_46651,N_47491);
or U48072 (N_48072,N_47095,N_46900);
and U48073 (N_48073,N_47297,N_46200);
or U48074 (N_48074,N_47482,N_47967);
and U48075 (N_48075,N_46297,N_46242);
and U48076 (N_48076,N_46452,N_46782);
and U48077 (N_48077,N_46348,N_47501);
xor U48078 (N_48078,N_47453,N_46280);
nor U48079 (N_48079,N_47041,N_46604);
nand U48080 (N_48080,N_46361,N_47404);
or U48081 (N_48081,N_47496,N_47925);
and U48082 (N_48082,N_47320,N_47798);
or U48083 (N_48083,N_47395,N_47632);
nor U48084 (N_48084,N_46088,N_46314);
and U48085 (N_48085,N_47339,N_46853);
or U48086 (N_48086,N_47828,N_46788);
or U48087 (N_48087,N_46974,N_46642);
and U48088 (N_48088,N_46123,N_46655);
nor U48089 (N_48089,N_47352,N_47944);
xor U48090 (N_48090,N_46295,N_47839);
nor U48091 (N_48091,N_46041,N_46000);
nand U48092 (N_48092,N_47414,N_46773);
or U48093 (N_48093,N_47456,N_47376);
xor U48094 (N_48094,N_47630,N_47027);
or U48095 (N_48095,N_47329,N_46784);
xor U48096 (N_48096,N_46961,N_46886);
nor U48097 (N_48097,N_46657,N_47053);
or U48098 (N_48098,N_47434,N_46550);
nor U48099 (N_48099,N_46215,N_47654);
or U48100 (N_48100,N_47999,N_46946);
xnor U48101 (N_48101,N_47303,N_46703);
and U48102 (N_48102,N_46667,N_46096);
xnor U48103 (N_48103,N_47950,N_47034);
and U48104 (N_48104,N_47832,N_46399);
or U48105 (N_48105,N_46739,N_46881);
nor U48106 (N_48106,N_46937,N_47497);
xnor U48107 (N_48107,N_46554,N_46723);
nor U48108 (N_48108,N_47439,N_47483);
nand U48109 (N_48109,N_46814,N_47646);
or U48110 (N_48110,N_47236,N_47892);
nand U48111 (N_48111,N_47764,N_47406);
nor U48112 (N_48112,N_47970,N_47959);
or U48113 (N_48113,N_47609,N_47979);
and U48114 (N_48114,N_46402,N_47280);
and U48115 (N_48115,N_47325,N_46444);
nor U48116 (N_48116,N_46666,N_47346);
nand U48117 (N_48117,N_47030,N_46034);
nand U48118 (N_48118,N_47814,N_47410);
nor U48119 (N_48119,N_47170,N_47331);
nand U48120 (N_48120,N_47254,N_46973);
nor U48121 (N_48121,N_47570,N_47664);
nand U48122 (N_48122,N_46345,N_46734);
nand U48123 (N_48123,N_46653,N_47514);
nand U48124 (N_48124,N_47844,N_47773);
xnor U48125 (N_48125,N_47327,N_47550);
or U48126 (N_48126,N_46749,N_47473);
nor U48127 (N_48127,N_47983,N_46490);
nand U48128 (N_48128,N_46207,N_46058);
and U48129 (N_48129,N_47381,N_46512);
xor U48130 (N_48130,N_46266,N_47077);
xnor U48131 (N_48131,N_47815,N_47207);
xor U48132 (N_48132,N_46634,N_46603);
nand U48133 (N_48133,N_46160,N_46744);
xor U48134 (N_48134,N_46992,N_46352);
nor U48135 (N_48135,N_46376,N_47477);
nand U48136 (N_48136,N_47282,N_47908);
or U48137 (N_48137,N_46736,N_47032);
xnor U48138 (N_48138,N_47962,N_46826);
or U48139 (N_48139,N_47868,N_47723);
and U48140 (N_48140,N_46405,N_47878);
nand U48141 (N_48141,N_46322,N_46180);
nor U48142 (N_48142,N_47652,N_46385);
or U48143 (N_48143,N_46037,N_47090);
and U48144 (N_48144,N_46648,N_46933);
or U48145 (N_48145,N_46870,N_47227);
or U48146 (N_48146,N_46003,N_46232);
and U48147 (N_48147,N_47972,N_47548);
and U48148 (N_48148,N_46776,N_47138);
or U48149 (N_48149,N_47240,N_47210);
or U48150 (N_48150,N_46124,N_46181);
xnor U48151 (N_48151,N_46247,N_47534);
and U48152 (N_48152,N_47267,N_47677);
nor U48153 (N_48153,N_46493,N_46112);
xor U48154 (N_48154,N_46504,N_47960);
or U48155 (N_48155,N_47356,N_47572);
nand U48156 (N_48156,N_47903,N_46865);
xnor U48157 (N_48157,N_47136,N_46308);
or U48158 (N_48158,N_47180,N_47279);
xor U48159 (N_48159,N_47049,N_47513);
and U48160 (N_48160,N_46465,N_46284);
xor U48161 (N_48161,N_47001,N_47011);
xnor U48162 (N_48162,N_46372,N_47161);
and U48163 (N_48163,N_46597,N_47607);
nand U48164 (N_48164,N_47708,N_46726);
and U48165 (N_48165,N_47805,N_47143);
or U48166 (N_48166,N_47158,N_47403);
nor U48167 (N_48167,N_46065,N_47374);
and U48168 (N_48168,N_46489,N_46662);
nand U48169 (N_48169,N_46898,N_46647);
nor U48170 (N_48170,N_46311,N_47223);
or U48171 (N_48171,N_47372,N_46713);
nor U48172 (N_48172,N_47448,N_46134);
nand U48173 (N_48173,N_46186,N_46095);
nor U48174 (N_48174,N_47703,N_46794);
xnor U48175 (N_48175,N_46936,N_46954);
xnor U48176 (N_48176,N_47073,N_46429);
and U48177 (N_48177,N_46695,N_46478);
xnor U48178 (N_48178,N_46128,N_47233);
nor U48179 (N_48179,N_46012,N_47334);
nor U48180 (N_48180,N_46686,N_46384);
nor U48181 (N_48181,N_46170,N_46175);
and U48182 (N_48182,N_46981,N_46285);
or U48183 (N_48183,N_47281,N_47155);
nand U48184 (N_48184,N_46633,N_47431);
nor U48185 (N_48185,N_47553,N_47596);
nor U48186 (N_48186,N_47123,N_47531);
nand U48187 (N_48187,N_47159,N_46854);
or U48188 (N_48188,N_46801,N_47089);
and U48189 (N_48189,N_47188,N_47066);
and U48190 (N_48190,N_47509,N_46500);
xnor U48191 (N_48191,N_47028,N_47666);
xor U48192 (N_48192,N_46809,N_46459);
nor U48193 (N_48193,N_46457,N_47394);
or U48194 (N_48194,N_47181,N_46863);
or U48195 (N_48195,N_47611,N_46211);
xnor U48196 (N_48196,N_47792,N_46110);
nand U48197 (N_48197,N_47603,N_47310);
and U48198 (N_48198,N_46618,N_47587);
nand U48199 (N_48199,N_47347,N_47451);
nor U48200 (N_48200,N_47809,N_46791);
xnor U48201 (N_48201,N_46872,N_47019);
and U48202 (N_48202,N_47508,N_46583);
or U48203 (N_48203,N_47396,N_47535);
nand U48204 (N_48204,N_46480,N_46233);
nand U48205 (N_48205,N_46456,N_47737);
nand U48206 (N_48206,N_47175,N_47389);
or U48207 (N_48207,N_47845,N_47400);
xor U48208 (N_48208,N_46205,N_47194);
and U48209 (N_48209,N_47463,N_46333);
nand U48210 (N_48210,N_47261,N_46165);
nor U48211 (N_48211,N_47031,N_46673);
or U48212 (N_48212,N_46932,N_47494);
nor U48213 (N_48213,N_47588,N_47520);
nor U48214 (N_48214,N_46283,N_47314);
nor U48215 (N_48215,N_46753,N_47012);
or U48216 (N_48216,N_46400,N_47493);
and U48217 (N_48217,N_46137,N_47409);
and U48218 (N_48218,N_47419,N_47552);
xnor U48219 (N_48219,N_46077,N_46516);
and U48220 (N_48220,N_46092,N_46737);
nand U48221 (N_48221,N_46862,N_47229);
or U48222 (N_48222,N_47848,N_46606);
xnor U48223 (N_48223,N_46397,N_46097);
nor U48224 (N_48224,N_46694,N_47930);
xnor U48225 (N_48225,N_46482,N_46039);
nand U48226 (N_48226,N_46157,N_47638);
or U48227 (N_48227,N_46393,N_47797);
nor U48228 (N_48228,N_47820,N_47527);
or U48229 (N_48229,N_47445,N_47881);
or U48230 (N_48230,N_47420,N_46447);
and U48231 (N_48231,N_47528,N_47103);
and U48232 (N_48232,N_46078,N_46995);
nand U48233 (N_48233,N_46559,N_46325);
nand U48234 (N_48234,N_47266,N_46743);
xnor U48235 (N_48235,N_47072,N_46381);
nand U48236 (N_48236,N_47885,N_46938);
and U48237 (N_48237,N_47046,N_46392);
or U48238 (N_48238,N_47847,N_47078);
and U48239 (N_48239,N_46271,N_47734);
or U48240 (N_48240,N_47813,N_46644);
and U48241 (N_48241,N_46747,N_47231);
nor U48242 (N_48242,N_47965,N_47009);
and U48243 (N_48243,N_46787,N_47595);
xor U48244 (N_48244,N_47020,N_46373);
or U48245 (N_48245,N_46008,N_46786);
nor U48246 (N_48246,N_46805,N_46724);
or U48247 (N_48247,N_47021,N_47767);
xor U48248 (N_48248,N_46684,N_47099);
and U48249 (N_48249,N_46761,N_46989);
and U48250 (N_48250,N_46721,N_47849);
nand U48251 (N_48251,N_46050,N_46529);
xnor U48252 (N_48252,N_47729,N_46859);
nor U48253 (N_48253,N_46437,N_47023);
or U48254 (N_48254,N_47830,N_47914);
xor U48255 (N_48255,N_47058,N_46631);
and U48256 (N_48256,N_46844,N_47142);
and U48257 (N_48257,N_47354,N_46571);
and U48258 (N_48258,N_46331,N_46965);
nor U48259 (N_48259,N_46835,N_46244);
nand U48260 (N_48260,N_46741,N_47397);
nand U48261 (N_48261,N_46602,N_47841);
nand U48262 (N_48262,N_46896,N_47932);
and U48263 (N_48263,N_47943,N_47920);
nor U48264 (N_48264,N_46698,N_46922);
nand U48265 (N_48265,N_47048,N_47523);
and U48266 (N_48266,N_47751,N_47189);
and U48267 (N_48267,N_46423,N_46199);
nand U48268 (N_48268,N_46803,N_46351);
or U48269 (N_48269,N_47793,N_47307);
or U48270 (N_48270,N_47662,N_46057);
nor U48271 (N_48271,N_46189,N_47537);
and U48272 (N_48272,N_46362,N_47198);
or U48273 (N_48273,N_46484,N_46979);
xnor U48274 (N_48274,N_47877,N_46868);
xor U48275 (N_48275,N_46464,N_47899);
and U48276 (N_48276,N_46171,N_46153);
nor U48277 (N_48277,N_46138,N_46884);
and U48278 (N_48278,N_46245,N_47366);
and U48279 (N_48279,N_46745,N_47316);
nor U48280 (N_48280,N_46009,N_46415);
nor U48281 (N_48281,N_47447,N_46612);
and U48282 (N_48282,N_47427,N_47516);
and U48283 (N_48283,N_46952,N_46760);
nor U48284 (N_48284,N_47752,N_46730);
and U48285 (N_48285,N_46026,N_47711);
xnor U48286 (N_48286,N_47713,N_46904);
xnor U48287 (N_48287,N_47160,N_46195);
or U48288 (N_48288,N_46090,N_46279);
xnor U48289 (N_48289,N_47760,N_47699);
and U48290 (N_48290,N_46978,N_46668);
nand U48291 (N_48291,N_46469,N_46909);
or U48292 (N_48292,N_47628,N_47165);
nor U48293 (N_48293,N_47554,N_46491);
xor U48294 (N_48294,N_46169,N_46338);
nor U48295 (N_48295,N_46441,N_46526);
xor U48296 (N_48296,N_47164,N_46980);
nor U48297 (N_48297,N_46116,N_46320);
xor U48298 (N_48298,N_47119,N_46764);
nor U48299 (N_48299,N_46840,N_46300);
nor U48300 (N_48300,N_46074,N_46687);
or U48301 (N_48301,N_47024,N_46313);
nor U48302 (N_48302,N_46388,N_46403);
nor U48303 (N_48303,N_46565,N_46833);
and U48304 (N_48304,N_46985,N_47659);
or U48305 (N_48305,N_46353,N_47230);
nor U48306 (N_48306,N_47051,N_47033);
nand U48307 (N_48307,N_46401,N_47913);
or U48308 (N_48308,N_47132,N_47192);
and U48309 (N_48309,N_46416,N_47799);
xor U48310 (N_48310,N_47821,N_46107);
nor U48311 (N_48311,N_47610,N_47226);
nor U48312 (N_48312,N_47720,N_47363);
nand U48313 (N_48313,N_46310,N_46640);
nor U48314 (N_48314,N_46332,N_46425);
or U48315 (N_48315,N_46335,N_47789);
and U48316 (N_48316,N_47156,N_46410);
and U48317 (N_48317,N_47616,N_46810);
xor U48318 (N_48318,N_46860,N_46146);
xnor U48319 (N_48319,N_47179,N_46010);
nor U48320 (N_48320,N_46681,N_47982);
xnor U48321 (N_48321,N_47529,N_47005);
and U48322 (N_48322,N_46850,N_47007);
xnor U48323 (N_48323,N_46911,N_46458);
nand U48324 (N_48324,N_47228,N_46975);
nor U48325 (N_48325,N_46424,N_47166);
nand U48326 (N_48326,N_47481,N_46638);
or U48327 (N_48327,N_46168,N_46129);
nand U48328 (N_48328,N_46173,N_47963);
and U48329 (N_48329,N_46696,N_46610);
and U48330 (N_48330,N_47843,N_47585);
xor U48331 (N_48331,N_46689,N_46774);
nand U48332 (N_48332,N_47893,N_46682);
and U48333 (N_48333,N_47582,N_46710);
xor U48334 (N_48334,N_46395,N_47459);
nand U48335 (N_48335,N_47232,N_47876);
or U48336 (N_48336,N_47846,N_46573);
nand U48337 (N_48337,N_47125,N_47429);
and U48338 (N_48338,N_47526,N_46238);
or U48339 (N_48339,N_46930,N_46976);
and U48340 (N_48340,N_46792,N_46349);
nor U48341 (N_48341,N_46318,N_46517);
nand U48342 (N_48342,N_46849,N_46264);
xor U48343 (N_48343,N_46236,N_46438);
xnor U48344 (N_48344,N_46094,N_46507);
nor U48345 (N_48345,N_47239,N_47359);
nor U48346 (N_48346,N_47904,N_47649);
nand U48347 (N_48347,N_47416,N_47627);
nand U48348 (N_48348,N_46148,N_46346);
or U48349 (N_48349,N_46025,N_46204);
xnor U48350 (N_48350,N_46832,N_46344);
xnor U48351 (N_48351,N_47308,N_47446);
or U48352 (N_48352,N_47525,N_47656);
nor U48353 (N_48353,N_47924,N_46357);
xnor U48354 (N_48354,N_46303,N_47698);
or U48355 (N_48355,N_46780,N_47321);
xnor U48356 (N_48356,N_47045,N_46894);
or U48357 (N_48357,N_46190,N_47387);
nand U48358 (N_48358,N_46476,N_47643);
and U48359 (N_48359,N_47601,N_47399);
or U48360 (N_48360,N_47612,N_47278);
nand U48361 (N_48361,N_46834,N_46923);
nor U48362 (N_48362,N_46907,N_46688);
nor U48363 (N_48363,N_46222,N_46903);
or U48364 (N_48364,N_46382,N_47786);
nor U48365 (N_48365,N_46893,N_46758);
or U48366 (N_48366,N_46433,N_47348);
nor U48367 (N_48367,N_47141,N_46679);
xor U48368 (N_48368,N_46364,N_47626);
and U48369 (N_48369,N_47104,N_46899);
and U48370 (N_48370,N_46558,N_47289);
nor U48371 (N_48371,N_47378,N_47301);
nor U48372 (N_48372,N_46449,N_46166);
xnor U48373 (N_48373,N_46968,N_47544);
nand U48374 (N_48374,N_47695,N_46312);
and U48375 (N_48375,N_46154,N_46004);
xnor U48376 (N_48376,N_47842,N_46054);
nor U48377 (N_48377,N_46185,N_46599);
nor U48378 (N_48378,N_47436,N_47006);
or U48379 (N_48379,N_47536,N_47215);
xnor U48380 (N_48380,N_46473,N_46187);
and U48381 (N_48381,N_46676,N_47515);
or U48382 (N_48382,N_47238,N_46093);
or U48383 (N_48383,N_46969,N_47867);
xor U48384 (N_48384,N_46113,N_46496);
and U48385 (N_48385,N_47300,N_46406);
and U48386 (N_48386,N_47110,N_46267);
and U48387 (N_48387,N_47807,N_46821);
nor U48388 (N_48388,N_47222,N_46196);
and U48389 (N_48389,N_47597,N_46986);
xnor U48390 (N_48390,N_47184,N_47201);
nand U48391 (N_48391,N_47302,N_46519);
xnor U48392 (N_48392,N_47811,N_47940);
xor U48393 (N_48393,N_46646,N_47096);
xnor U48394 (N_48394,N_47978,N_46567);
xor U48395 (N_48395,N_47689,N_46389);
or U48396 (N_48396,N_47579,N_47665);
and U48397 (N_48397,N_47748,N_46763);
or U48398 (N_48398,N_46118,N_46685);
or U48399 (N_48399,N_47398,N_46824);
xnor U48400 (N_48400,N_47413,N_46049);
or U48401 (N_48401,N_46518,N_46495);
nand U48402 (N_48402,N_46060,N_47246);
xor U48403 (N_48403,N_47108,N_46874);
nand U48404 (N_48404,N_47524,N_47083);
xor U48405 (N_48405,N_47178,N_47706);
nand U48406 (N_48406,N_46309,N_47360);
nand U48407 (N_48407,N_46715,N_47693);
nor U48408 (N_48408,N_46839,N_47357);
and U48409 (N_48409,N_47485,N_46430);
xor U48410 (N_48410,N_47185,N_47621);
and U48411 (N_48411,N_47478,N_47898);
and U48412 (N_48412,N_46751,N_47146);
or U48413 (N_48413,N_47644,N_46523);
nor U48414 (N_48414,N_47801,N_46011);
or U48415 (N_48415,N_46260,N_47517);
nor U48416 (N_48416,N_47495,N_46230);
and U48417 (N_48417,N_47162,N_46105);
xor U48418 (N_48418,N_46150,N_47237);
xnor U48419 (N_48419,N_46117,N_47969);
or U48420 (N_48420,N_47512,N_47576);
xnor U48421 (N_48421,N_47056,N_46347);
and U48422 (N_48422,N_46925,N_47137);
nor U48423 (N_48423,N_47992,N_46391);
and U48424 (N_48424,N_46184,N_46435);
nor U48425 (N_48425,N_47705,N_46258);
nor U48426 (N_48426,N_47560,N_46001);
or U48427 (N_48427,N_47598,N_47687);
nand U48428 (N_48428,N_46278,N_47062);
or U48429 (N_48429,N_46906,N_47377);
nor U48430 (N_48430,N_47326,N_47522);
or U48431 (N_48431,N_47870,N_47315);
xor U48432 (N_48432,N_47530,N_46203);
nor U48433 (N_48433,N_46557,N_47974);
nand U48434 (N_48434,N_46358,N_46595);
nor U48435 (N_48435,N_46298,N_46993);
xor U48436 (N_48436,N_47407,N_47667);
and U48437 (N_48437,N_47284,N_47724);
nand U48438 (N_48438,N_47422,N_47163);
and U48439 (N_48439,N_46367,N_47174);
nand U48440 (N_48440,N_46609,N_47268);
nor U48441 (N_48441,N_46649,N_46404);
and U48442 (N_48442,N_47016,N_47367);
xnor U48443 (N_48443,N_46935,N_46605);
nor U48444 (N_48444,N_46047,N_47273);
or U48445 (N_48445,N_46071,N_46115);
and U48446 (N_48446,N_46997,N_46063);
and U48447 (N_48447,N_47697,N_47298);
or U48448 (N_48448,N_46183,N_47264);
or U48449 (N_48449,N_47853,N_47953);
xnor U48450 (N_48450,N_47084,N_47126);
or U48451 (N_48451,N_47637,N_47717);
and U48452 (N_48452,N_47911,N_46365);
nand U48453 (N_48453,N_47441,N_46193);
and U48454 (N_48454,N_46164,N_46873);
and U48455 (N_48455,N_47725,N_47683);
or U48456 (N_48456,N_46255,N_47470);
xnor U48457 (N_48457,N_46951,N_47984);
nand U48458 (N_48458,N_47614,N_46188);
xnor U48459 (N_48459,N_46142,N_46218);
xor U48460 (N_48460,N_46072,N_47958);
nor U48461 (N_48461,N_47274,N_47017);
xnor U48462 (N_48462,N_46555,N_47475);
nor U48463 (N_48463,N_47202,N_46498);
or U48464 (N_48464,N_47539,N_46908);
or U48465 (N_48465,N_46522,N_46330);
nor U48466 (N_48466,N_46040,N_46846);
xor U48467 (N_48467,N_46262,N_46729);
nor U48468 (N_48468,N_46917,N_47765);
or U48469 (N_48469,N_46971,N_46947);
or U48470 (N_48470,N_47599,N_46656);
or U48471 (N_48471,N_46802,N_47145);
xnor U48472 (N_48472,N_46757,N_47946);
nor U48473 (N_48473,N_47922,N_46806);
nor U48474 (N_48474,N_46716,N_47129);
or U48475 (N_48475,N_47749,N_46336);
nand U48476 (N_48476,N_46560,N_46772);
and U48477 (N_48477,N_46918,N_47474);
or U48478 (N_48478,N_47935,N_46643);
or U48479 (N_48479,N_46926,N_47902);
xor U48480 (N_48480,N_47069,N_47113);
nand U48481 (N_48481,N_47541,N_47247);
nand U48482 (N_48482,N_47504,N_47740);
or U48483 (N_48483,N_47388,N_46940);
xor U48484 (N_48484,N_47670,N_47910);
xor U48485 (N_48485,N_47121,N_46665);
nor U48486 (N_48486,N_46289,N_46342);
or U48487 (N_48487,N_46174,N_46419);
nand U48488 (N_48488,N_47252,N_46875);
nor U48489 (N_48489,N_46087,N_46386);
nand U48490 (N_48490,N_46119,N_46256);
nand U48491 (N_48491,N_46483,N_47219);
and U48492 (N_48492,N_47443,N_47873);
nand U48493 (N_48493,N_47382,N_47709);
xnor U48494 (N_48494,N_46485,N_46201);
nor U48495 (N_48495,N_47657,N_46102);
and U48496 (N_48496,N_46996,N_47002);
nor U48497 (N_48497,N_47296,N_47968);
nor U48498 (N_48498,N_47371,N_47070);
or U48499 (N_48499,N_46368,N_47018);
nand U48500 (N_48500,N_46547,N_47263);
or U48501 (N_48501,N_47584,N_46611);
xnor U48502 (N_48502,N_47593,N_47696);
nor U48503 (N_48503,N_46864,N_47022);
and U48504 (N_48504,N_46378,N_46159);
or U48505 (N_48505,N_46650,N_47014);
xnor U48506 (N_48506,N_47039,N_47342);
xnor U48507 (N_48507,N_47109,N_47629);
or U48508 (N_48508,N_47258,N_47778);
xnor U48509 (N_48509,N_46125,N_47886);
nand U48510 (N_48510,N_47127,N_47613);
and U48511 (N_48511,N_47276,N_47825);
nor U48512 (N_48512,N_46924,N_47936);
or U48513 (N_48513,N_46439,N_46674);
nand U48514 (N_48514,N_47433,N_47952);
xor U48515 (N_48515,N_47988,N_47140);
nand U48516 (N_48516,N_47879,N_47183);
xnor U48517 (N_48517,N_46334,N_47362);
or U48518 (N_48518,N_46221,N_46286);
and U48519 (N_48519,N_47452,N_47506);
and U48520 (N_48520,N_47424,N_46499);
nand U48521 (N_48521,N_47618,N_47097);
and U48522 (N_48522,N_46781,N_47800);
nand U48523 (N_48523,N_47461,N_47428);
or U48524 (N_48524,N_46813,N_46534);
or U48525 (N_48525,N_46005,N_46294);
or U48526 (N_48526,N_47209,N_47575);
or U48527 (N_48527,N_46167,N_46214);
nor U48528 (N_48528,N_46127,N_47154);
nor U48529 (N_48529,N_46052,N_46528);
or U48530 (N_48530,N_47635,N_47311);
or U48531 (N_48531,N_46067,N_47107);
nand U48532 (N_48532,N_47956,N_46738);
xnor U48533 (N_48533,N_47087,N_47197);
and U48534 (N_48534,N_47928,N_46350);
xor U48535 (N_48535,N_47176,N_47650);
and U48536 (N_48536,N_46191,N_46426);
and U48537 (N_48537,N_47918,N_46847);
or U48538 (N_48538,N_47673,N_46535);
xnor U48539 (N_48539,N_46234,N_46861);
nand U48540 (N_48540,N_47379,N_46766);
or U48541 (N_48541,N_46680,N_47338);
and U48542 (N_48542,N_46988,N_46770);
nor U48543 (N_48543,N_47469,N_46587);
xnor U48544 (N_48544,N_47557,N_47417);
nand U48545 (N_48545,N_47283,N_46596);
xor U48546 (N_48546,N_47681,N_46845);
or U48547 (N_48547,N_46987,N_47771);
nand U48548 (N_48548,N_46409,N_47462);
nand U48549 (N_48549,N_46672,N_46746);
or U48550 (N_48550,N_46945,N_46527);
and U48551 (N_48551,N_46210,N_46579);
and U48552 (N_48552,N_46136,N_47647);
xor U48553 (N_48553,N_46530,N_47212);
nor U48554 (N_48554,N_47479,N_46869);
xor U48555 (N_48555,N_46970,N_46056);
xor U48556 (N_48556,N_47906,N_46273);
xnor U48557 (N_48557,N_47243,N_46871);
and U48558 (N_48558,N_46179,N_46006);
nand U48559 (N_48559,N_47555,N_47775);
and U48560 (N_48560,N_46488,N_47341);
or U48561 (N_48561,N_47966,N_46251);
nand U48562 (N_48562,N_47405,N_46711);
or U48563 (N_48563,N_47054,N_47128);
xor U48564 (N_48564,N_46675,N_47648);
nor U48565 (N_48565,N_46706,N_47571);
nand U48566 (N_48566,N_46014,N_47819);
nand U48567 (N_48567,N_47880,N_46261);
nor U48568 (N_48568,N_47081,N_46066);
or U48569 (N_48569,N_46287,N_46795);
or U48570 (N_48570,N_46645,N_47816);
or U48571 (N_48571,N_46209,N_47476);
or U48572 (N_48572,N_46035,N_46818);
or U48573 (N_48573,N_46654,N_46598);
nor U48574 (N_48574,N_46799,N_47604);
xnor U48575 (N_48575,N_47082,N_47025);
xor U48576 (N_48576,N_47900,N_46614);
nand U48577 (N_48577,N_47488,N_47887);
nor U48578 (N_48578,N_46820,N_47384);
nor U48579 (N_48579,N_46866,N_47364);
and U48580 (N_48580,N_47457,N_46525);
or U48581 (N_48581,N_47727,N_47738);
nor U48582 (N_48582,N_46690,N_46239);
nand U48583 (N_48583,N_47772,N_47716);
nor U48584 (N_48584,N_47086,N_46228);
xor U48585 (N_48585,N_47542,N_46227);
or U48586 (N_48586,N_47147,N_47454);
nand U48587 (N_48587,N_47874,N_46337);
xnor U48588 (N_48588,N_47393,N_46461);
xor U48589 (N_48589,N_47323,N_47574);
nand U48590 (N_48590,N_46472,N_46360);
nor U48591 (N_48591,N_46549,N_47294);
and U48592 (N_48592,N_46632,N_47199);
and U48593 (N_48593,N_46324,N_47259);
or U48594 (N_48594,N_46291,N_47423);
nor U48595 (N_48595,N_47938,N_47116);
nand U48596 (N_48596,N_47768,N_46269);
xor U48597 (N_48597,N_46966,N_46206);
xnor U48598 (N_48598,N_46293,N_47964);
nor U48599 (N_48599,N_46027,N_47206);
nand U48600 (N_48600,N_47971,N_47661);
xnor U48601 (N_48601,N_47245,N_46624);
nand U48602 (N_48602,N_46492,N_46217);
and U48603 (N_48603,N_47309,N_47466);
xor U48604 (N_48604,N_47645,N_47583);
or U48605 (N_48605,N_46619,N_46213);
xor U48606 (N_48606,N_46414,N_46804);
or U48607 (N_48607,N_47234,N_47047);
nor U48608 (N_48608,N_46543,N_46371);
or U48609 (N_48609,N_47859,N_46921);
nand U48610 (N_48610,N_47015,N_46075);
and U48611 (N_48611,N_47059,N_46202);
or U48612 (N_48612,N_46145,N_47577);
or U48613 (N_48613,N_46323,N_47931);
or U48614 (N_48614,N_47344,N_46783);
nor U48615 (N_48615,N_46390,N_46510);
nand U48616 (N_48616,N_46912,N_46719);
nand U48617 (N_48617,N_46100,N_47074);
or U48618 (N_48618,N_46038,N_47134);
and U48619 (N_48619,N_47769,N_47205);
and U48620 (N_48620,N_47602,N_46212);
nor U48621 (N_48621,N_46591,N_46158);
nor U48622 (N_48622,N_46216,N_47581);
xor U48623 (N_48623,N_46443,N_47707);
nand U48624 (N_48624,N_46445,N_47003);
nand U48625 (N_48625,N_46103,N_46086);
nand U48626 (N_48626,N_46446,N_47455);
and U48627 (N_48627,N_47980,N_47712);
nor U48628 (N_48628,N_46268,N_47855);
xor U48629 (N_48629,N_47854,N_46249);
or U48630 (N_48630,N_46641,N_47937);
and U48631 (N_48631,N_47736,N_46431);
or U48632 (N_48632,N_46520,N_46942);
and U48633 (N_48633,N_46466,N_47655);
nor U48634 (N_48634,N_46501,N_46545);
and U48635 (N_48635,N_46566,N_47779);
xnor U48636 (N_48636,N_46048,N_46702);
and U48637 (N_48637,N_47755,N_47242);
xor U48638 (N_48638,N_47942,N_46326);
or U48639 (N_48639,N_47065,N_46927);
and U48640 (N_48640,N_47169,N_46575);
nand U48641 (N_48641,N_46132,N_47244);
nand U48642 (N_48642,N_47660,N_47402);
and U48643 (N_48643,N_46099,N_46417);
nor U48644 (N_48644,N_47195,N_46720);
nand U48645 (N_48645,N_47167,N_47562);
and U48646 (N_48646,N_46220,N_47182);
or U48647 (N_48647,N_47345,N_46637);
xor U48648 (N_48648,N_47133,N_46607);
nor U48649 (N_48649,N_47824,N_46223);
nor U48650 (N_48650,N_46728,N_46301);
or U48651 (N_48651,N_47383,N_46241);
or U48652 (N_48652,N_47000,N_46664);
and U48653 (N_48653,N_46622,N_47976);
xnor U48654 (N_48654,N_47826,N_47901);
nor U48655 (N_48655,N_46477,N_47285);
or U48656 (N_48656,N_46570,N_47545);
xnor U48657 (N_48657,N_46315,N_47861);
and U48658 (N_48658,N_46576,N_46023);
or U48659 (N_48659,N_47688,N_46765);
xor U48660 (N_48660,N_46076,N_47700);
nor U48661 (N_48661,N_47869,N_47784);
xor U48662 (N_48662,N_47758,N_46704);
or U48663 (N_48663,N_47440,N_47224);
nand U48664 (N_48664,N_47998,N_46511);
xnor U48665 (N_48665,N_47671,N_46513);
and U48666 (N_48666,N_47973,N_47766);
nand U48667 (N_48667,N_46141,N_47391);
or U48668 (N_48668,N_46827,N_47955);
and U48669 (N_48669,N_47947,N_46621);
nor U48670 (N_48670,N_46019,N_46383);
or U48671 (N_48671,N_46740,N_46539);
nand U48672 (N_48672,N_46084,N_47860);
or U48673 (N_48673,N_46420,N_46509);
nand U48674 (N_48674,N_46502,N_47430);
nor U48675 (N_48675,N_46275,N_47685);
nand U48676 (N_48676,N_47991,N_47115);
or U48677 (N_48677,N_47995,N_46958);
and U48678 (N_48678,N_47957,N_47153);
xnor U48679 (N_48679,N_47114,N_47250);
nor U48680 (N_48680,N_46083,N_47313);
and U48681 (N_48681,N_46521,N_47679);
xor U48682 (N_48682,N_47586,N_47449);
or U48683 (N_48683,N_46340,N_47105);
nor U48684 (N_48684,N_47425,N_47701);
nand U48685 (N_48685,N_47684,N_46475);
nand U48686 (N_48686,N_47663,N_47894);
and U48687 (N_48687,N_47538,N_46536);
nand U48688 (N_48688,N_47905,N_46830);
or U48689 (N_48689,N_47804,N_46901);
nand U48690 (N_48690,N_47573,N_47642);
nand U48691 (N_48691,N_47186,N_47858);
nand U48692 (N_48692,N_46752,N_46304);
or U48693 (N_48693,N_46379,N_47631);
or U48694 (N_48694,N_47013,N_46588);
and U48695 (N_48695,N_46616,N_47390);
nand U48696 (N_48696,N_47218,N_46876);
or U48697 (N_48697,N_47149,N_46343);
and U48698 (N_48698,N_47633,N_47337);
or U48699 (N_48699,N_47330,N_46064);
or U48700 (N_48700,N_47890,N_46016);
nor U48701 (N_48701,N_46111,N_46036);
nand U48702 (N_48702,N_46592,N_47822);
nor U48703 (N_48703,N_46029,N_47636);
xnor U48704 (N_48704,N_47124,N_47929);
or U48705 (N_48705,N_47521,N_47566);
or U48706 (N_48706,N_47211,N_46257);
and U48707 (N_48707,N_47823,N_47235);
nand U48708 (N_48708,N_47640,N_46341);
xnor U48709 (N_48709,N_47884,N_47608);
or U48710 (N_48710,N_47863,N_47370);
nand U48711 (N_48711,N_47442,N_46018);
and U48712 (N_48712,N_47157,N_47385);
and U48713 (N_48713,N_47029,N_47203);
xor U48714 (N_48714,N_47829,N_46754);
xnor U48715 (N_48715,N_47718,N_46553);
nand U48716 (N_48716,N_47060,N_47071);
nor U48717 (N_48717,N_47401,N_47996);
or U48718 (N_48718,N_46474,N_46759);
or U48719 (N_48719,N_47270,N_47728);
nand U48720 (N_48720,N_47038,N_47945);
or U48721 (N_48721,N_47565,N_47004);
or U48722 (N_48722,N_47484,N_47675);
or U48723 (N_48723,N_47559,N_47426);
nand U48724 (N_48724,N_47026,N_46366);
nor U48725 (N_48725,N_47190,N_46237);
nand U48726 (N_48726,N_46878,N_46963);
nor U48727 (N_48727,N_46882,N_47840);
or U48728 (N_48728,N_46091,N_47812);
xnor U48729 (N_48729,N_47464,N_46727);
or U48730 (N_48730,N_46374,N_47120);
xor U48731 (N_48731,N_46081,N_47796);
nor U48732 (N_48732,N_47304,N_46994);
or U48733 (N_48733,N_47563,N_46288);
xor U48734 (N_48734,N_47668,N_46306);
nand U48735 (N_48735,N_46660,N_46462);
and U48736 (N_48736,N_47546,N_47856);
or U48737 (N_48737,N_47365,N_46370);
xnor U48738 (N_48738,N_47907,N_46934);
xor U48739 (N_48739,N_47533,N_46544);
nor U48740 (N_48740,N_46411,N_47851);
nor U48741 (N_48741,N_47241,N_46879);
or U48742 (N_48742,N_46807,N_47438);
or U48743 (N_48743,N_46692,N_46842);
and U48744 (N_48744,N_47510,N_46486);
and U48745 (N_48745,N_46505,N_46948);
nor U48746 (N_48746,N_46584,N_47111);
xor U48747 (N_48747,N_46131,N_47897);
and U48748 (N_48748,N_46777,N_47692);
and U48749 (N_48749,N_46162,N_47010);
and U48750 (N_48750,N_47704,N_47322);
or U48751 (N_48751,N_46897,N_46328);
nand U48752 (N_48752,N_47997,N_46471);
nor U48753 (N_48753,N_47567,N_47590);
and U48754 (N_48754,N_46953,N_46231);
and U48755 (N_48755,N_47355,N_46652);
nand U48756 (N_48756,N_46104,N_46636);
and U48757 (N_48757,N_47008,N_46121);
xor U48758 (N_48758,N_47265,N_46307);
or U48759 (N_48759,N_46412,N_46156);
or U48760 (N_48760,N_46319,N_47750);
nand U48761 (N_48761,N_46828,N_47615);
xnor U48762 (N_48762,N_47487,N_46902);
nor U48763 (N_48763,N_46451,N_47933);
xor U48764 (N_48764,N_47332,N_47694);
and U48765 (N_48765,N_46831,N_47498);
nor U48766 (N_48766,N_47754,N_46079);
nor U48767 (N_48767,N_46068,N_47063);
and U48768 (N_48768,N_46032,N_46497);
nand U48769 (N_48769,N_46418,N_46149);
or U48770 (N_48770,N_46140,N_46829);
or U48771 (N_48771,N_46811,N_47392);
xnor U48772 (N_48772,N_46329,N_46790);
and U48773 (N_48773,N_47949,N_46812);
xor U48774 (N_48774,N_47150,N_46002);
nor U48775 (N_48775,N_46240,N_47040);
or U48776 (N_48776,N_46450,N_47286);
or U48777 (N_48777,N_47731,N_46182);
and U48778 (N_48778,N_46693,N_46022);
nor U48779 (N_48779,N_47921,N_46552);
nor U48780 (N_48780,N_47131,N_46327);
xnor U48781 (N_48781,N_47044,N_47561);
and U48782 (N_48782,N_47486,N_46700);
xor U48783 (N_48783,N_46608,N_47916);
nand U48784 (N_48784,N_47292,N_46046);
xor U48785 (N_48785,N_47719,N_47187);
or U48786 (N_48786,N_47744,N_47172);
xor U48787 (N_48787,N_47135,N_47106);
nor U48788 (N_48788,N_47954,N_47368);
or U48789 (N_48789,N_46880,N_47091);
nor U48790 (N_48790,N_46428,N_46479);
and U48791 (N_48791,N_47817,N_47721);
or U48792 (N_48792,N_47248,N_47421);
and U48793 (N_48793,N_46944,N_46133);
xor U48794 (N_48794,N_47122,N_47335);
and U48795 (N_48795,N_47118,N_47990);
nor U48796 (N_48796,N_47743,N_47676);
and U48797 (N_48797,N_47380,N_47770);
and U48798 (N_48798,N_47619,N_47730);
xnor U48799 (N_48799,N_47795,N_47503);
xor U48800 (N_48800,N_47200,N_47746);
nand U48801 (N_48801,N_46931,N_47225);
or U48802 (N_48802,N_46836,N_46051);
nor U48803 (N_48803,N_46013,N_46895);
nand U48804 (N_48804,N_46061,N_46421);
and U48805 (N_48805,N_46796,N_46494);
and U48806 (N_48806,N_46797,N_46413);
nand U48807 (N_48807,N_47037,N_47061);
and U48808 (N_48808,N_47625,N_46769);
or U48809 (N_48809,N_46356,N_46722);
nand U48810 (N_48810,N_47865,N_47340);
nand U48811 (N_48811,N_46062,N_47460);
xor U48812 (N_48812,N_46959,N_47152);
and U48813 (N_48813,N_46106,N_46714);
xnor U48814 (N_48814,N_47653,N_46957);
and U48815 (N_48815,N_47468,N_46152);
nor U48816 (N_48816,N_47986,N_47669);
and U48817 (N_48817,N_47353,N_47173);
nand U48818 (N_48818,N_47702,N_47912);
xor U48819 (N_48819,N_46837,N_46767);
or U48820 (N_48820,N_47917,N_47891);
and U48821 (N_48821,N_47480,N_47458);
xor U48822 (N_48822,N_47295,N_46916);
xnor U48823 (N_48823,N_46467,N_46120);
nor U48824 (N_48824,N_47862,N_47852);
or U48825 (N_48825,N_47714,N_47569);
or U48826 (N_48826,N_47732,N_47269);
nand U48827 (N_48827,N_47781,N_46021);
xor U48828 (N_48828,N_46941,N_46354);
nor U48829 (N_48829,N_47196,N_46627);
nor U48830 (N_48830,N_47710,N_46055);
nor U48831 (N_48831,N_47139,N_46246);
nor U48832 (N_48832,N_46920,N_46225);
and U48833 (N_48833,N_46659,N_47489);
nand U48834 (N_48834,N_47806,N_47490);
and U48835 (N_48835,N_46590,N_46274);
and U48836 (N_48836,N_47088,N_47549);
or U48837 (N_48837,N_46043,N_46551);
nand U48838 (N_48838,N_46742,N_46254);
xor U48839 (N_48839,N_47634,N_47864);
xor U48840 (N_48840,N_46114,N_47092);
or U48841 (N_48841,N_47558,N_47589);
and U48842 (N_48842,N_46683,N_46030);
nand U48843 (N_48843,N_46705,N_47836);
nor U48844 (N_48844,N_47951,N_46276);
and U48845 (N_48845,N_47827,N_47467);
and U48846 (N_48846,N_46582,N_47994);
nand U48847 (N_48847,N_46669,N_46851);
and U48848 (N_48848,N_47277,N_46139);
xor U48849 (N_48849,N_47741,N_46155);
nor U48850 (N_48850,N_47939,N_47036);
or U48851 (N_48851,N_46563,N_46470);
and U48852 (N_48852,N_47818,N_47102);
xor U48853 (N_48853,N_46625,N_46915);
and U48854 (N_48854,N_46709,N_46126);
or U48855 (N_48855,N_47606,N_46282);
nor U48856 (N_48856,N_47290,N_47328);
and U48857 (N_48857,N_46108,N_46919);
or U48858 (N_48858,N_46192,N_47412);
xor U48859 (N_48859,N_46670,N_46677);
xnor U48860 (N_48860,N_46178,N_46375);
xor U48861 (N_48861,N_46020,N_46635);
and U48862 (N_48862,N_47260,N_47872);
or U48863 (N_48863,N_46541,N_47055);
and U48864 (N_48864,N_47272,N_46460);
nor U48865 (N_48865,N_46793,N_47505);
or U48866 (N_48866,N_47735,N_47715);
and U48867 (N_48867,N_46355,N_46725);
nor U48868 (N_48868,N_47774,N_47658);
nor U48869 (N_48869,N_47101,N_47220);
and U48870 (N_48870,N_46515,N_46691);
nor U48871 (N_48871,N_46855,N_46613);
nand U48872 (N_48872,N_47511,N_47191);
nand U48873 (N_48873,N_47989,N_46785);
and U48874 (N_48874,N_46524,N_46593);
and U48875 (N_48875,N_47386,N_47287);
xor U48876 (N_48876,N_47802,N_47540);
xnor U48877 (N_48877,N_46455,N_46568);
and U48878 (N_48878,N_47794,N_46073);
and U48879 (N_48879,N_47780,N_47333);
nor U48880 (N_48880,N_46852,N_47834);
nand U48881 (N_48881,N_46177,N_46998);
xor U48882 (N_48882,N_46024,N_46630);
or U48883 (N_48883,N_47788,N_46387);
xor U48884 (N_48884,N_46701,N_46819);
nor U48885 (N_48885,N_46250,N_47617);
nor U48886 (N_48886,N_47518,N_47672);
and U48887 (N_48887,N_47100,N_47993);
nand U48888 (N_48888,N_46144,N_47753);
nor U48889 (N_48889,N_46589,N_46503);
or U48890 (N_48890,N_47987,N_46080);
and U48891 (N_48891,N_47177,N_46732);
xnor U48892 (N_48892,N_46453,N_46983);
and U48893 (N_48893,N_46889,N_46626);
xor U48894 (N_48894,N_47927,N_46628);
nor U48895 (N_48895,N_47075,N_46808);
or U48896 (N_48896,N_46977,N_47985);
xor U48897 (N_48897,N_47543,N_46537);
and U48898 (N_48898,N_46317,N_47094);
or U48899 (N_48899,N_46928,N_47217);
and U48900 (N_48900,N_46028,N_47733);
xor U48901 (N_48901,N_46574,N_47318);
nor U48902 (N_48902,N_47288,N_46768);
nand U48903 (N_48903,N_46359,N_46163);
nand U48904 (N_48904,N_46197,N_47042);
nand U48905 (N_48905,N_47747,N_46890);
nor U48906 (N_48906,N_46962,N_46731);
xnor U48907 (N_48907,N_46396,N_47256);
nand U48908 (N_48908,N_46581,N_47722);
nor U48909 (N_48909,N_47888,N_47745);
nand U48910 (N_48910,N_47349,N_47909);
xnor U48911 (N_48911,N_46964,N_46398);
or U48912 (N_48912,N_46779,N_46408);
or U48913 (N_48913,N_46639,N_47934);
or U48914 (N_48914,N_46623,N_46914);
xnor U48915 (N_48915,N_46999,N_46678);
or U48916 (N_48916,N_47926,N_46718);
nand U48917 (N_48917,N_46843,N_47043);
nand U48918 (N_48918,N_46564,N_47437);
or U48919 (N_48919,N_47373,N_47691);
or U48920 (N_48920,N_46007,N_47351);
nand U48921 (N_48921,N_47317,N_47981);
nor U48922 (N_48922,N_46292,N_47130);
nor U48923 (N_48923,N_46101,N_47803);
xnor U48924 (N_48924,N_46905,N_46658);
xor U48925 (N_48925,N_46990,N_47756);
xor U48926 (N_48926,N_46542,N_46290);
nand U48927 (N_48927,N_47221,N_47450);
and U48928 (N_48928,N_46800,N_47726);
nor U48929 (N_48929,N_46031,N_46600);
xnor U48930 (N_48930,N_46762,N_47882);
and U48931 (N_48931,N_46580,N_46816);
and U48932 (N_48932,N_46750,N_47262);
xnor U48933 (N_48933,N_46789,N_46771);
xnor U48934 (N_48934,N_46620,N_47336);
and U48935 (N_48935,N_47052,N_46877);
and U48936 (N_48936,N_46272,N_47915);
and U48937 (N_48937,N_46044,N_46712);
nand U48938 (N_48938,N_46253,N_47050);
or U48939 (N_48939,N_47578,N_47564);
nor U48940 (N_48940,N_46481,N_46857);
and U48941 (N_48941,N_47465,N_46305);
and U48942 (N_48942,N_47651,N_46059);
xor U48943 (N_48943,N_46302,N_46822);
nor U48944 (N_48944,N_46161,N_46572);
xnor U48945 (N_48945,N_47568,N_47977);
nand U48946 (N_48946,N_47148,N_46259);
or U48947 (N_48947,N_46176,N_47271);
or U48948 (N_48948,N_46263,N_46130);
nor U48949 (N_48949,N_47214,N_46033);
or U48950 (N_48950,N_46815,N_47923);
xnor U48951 (N_48951,N_46717,N_46226);
xor U48952 (N_48952,N_46487,N_47472);
nand U48953 (N_48953,N_46432,N_46748);
xnor U48954 (N_48954,N_47580,N_46913);
nand U48955 (N_48955,N_47507,N_46422);
nand U48956 (N_48956,N_46950,N_46299);
nor U48957 (N_48957,N_47098,N_47080);
and U48958 (N_48958,N_47418,N_47415);
nor U48959 (N_48959,N_46708,N_47857);
nor U48960 (N_48960,N_46755,N_46960);
nand U48961 (N_48961,N_46883,N_47866);
xor U48962 (N_48962,N_46892,N_47519);
or U48963 (N_48963,N_47639,N_47319);
nor U48964 (N_48964,N_47623,N_46661);
or U48965 (N_48965,N_46506,N_47293);
nor U48966 (N_48966,N_46956,N_47204);
and U48967 (N_48967,N_46955,N_46407);
nor U48968 (N_48968,N_46578,N_46098);
or U48969 (N_48969,N_46442,N_47810);
nor U48970 (N_48970,N_47896,N_46972);
and U48971 (N_48971,N_46508,N_47782);
nand U48972 (N_48972,N_46440,N_47249);
or U48973 (N_48973,N_47291,N_46147);
xnor U48974 (N_48974,N_47168,N_47532);
and U48975 (N_48975,N_46887,N_47444);
nand U48976 (N_48976,N_46143,N_46281);
xor U48977 (N_48977,N_47831,N_46042);
and U48978 (N_48978,N_47895,N_47253);
nor U48979 (N_48979,N_46885,N_47358);
nor U48980 (N_48980,N_47306,N_46172);
and U48981 (N_48981,N_47591,N_46448);
and U48982 (N_48982,N_46697,N_46601);
or U48983 (N_48983,N_46045,N_46699);
or U48984 (N_48984,N_46436,N_46858);
nor U48985 (N_48985,N_47678,N_47093);
nor U48986 (N_48986,N_47690,N_47783);
and U48987 (N_48987,N_47085,N_47875);
xor U48988 (N_48988,N_47941,N_47324);
nor U48989 (N_48989,N_46265,N_46296);
nand U48990 (N_48990,N_47208,N_46514);
nor U48991 (N_48991,N_46339,N_46548);
or U48992 (N_48992,N_46394,N_46248);
xnor U48993 (N_48993,N_46540,N_46194);
and U48994 (N_48994,N_47837,N_46594);
and U48995 (N_48995,N_46229,N_46070);
nand U48996 (N_48996,N_47193,N_46208);
nand U48997 (N_48997,N_46629,N_47686);
xnor U48998 (N_48998,N_47605,N_47838);
nand U48999 (N_48999,N_46823,N_46929);
nor U49000 (N_49000,N_47909,N_46007);
xnor U49001 (N_49001,N_46807,N_47230);
nor U49002 (N_49002,N_47277,N_46601);
xnor U49003 (N_49003,N_47918,N_47821);
or U49004 (N_49004,N_47156,N_47382);
nor U49005 (N_49005,N_47163,N_47520);
nor U49006 (N_49006,N_46037,N_46346);
xnor U49007 (N_49007,N_46032,N_46565);
nor U49008 (N_49008,N_46337,N_47086);
or U49009 (N_49009,N_46806,N_47625);
or U49010 (N_49010,N_46254,N_47673);
xor U49011 (N_49011,N_46019,N_47940);
nand U49012 (N_49012,N_47794,N_47138);
xnor U49013 (N_49013,N_47336,N_47338);
xor U49014 (N_49014,N_47942,N_47030);
xnor U49015 (N_49015,N_46551,N_47806);
xnor U49016 (N_49016,N_47860,N_46807);
xor U49017 (N_49017,N_46565,N_47882);
or U49018 (N_49018,N_47188,N_47187);
and U49019 (N_49019,N_47280,N_47302);
and U49020 (N_49020,N_47861,N_46361);
xor U49021 (N_49021,N_47862,N_46001);
or U49022 (N_49022,N_47400,N_47662);
and U49023 (N_49023,N_47255,N_46509);
and U49024 (N_49024,N_47273,N_46304);
nor U49025 (N_49025,N_46016,N_47945);
or U49026 (N_49026,N_47007,N_47130);
nand U49027 (N_49027,N_47614,N_47989);
xor U49028 (N_49028,N_47577,N_47430);
or U49029 (N_49029,N_46468,N_47659);
xnor U49030 (N_49030,N_46375,N_47348);
and U49031 (N_49031,N_47026,N_47444);
nor U49032 (N_49032,N_46362,N_46497);
xor U49033 (N_49033,N_47341,N_47086);
or U49034 (N_49034,N_47055,N_46513);
or U49035 (N_49035,N_47145,N_46780);
and U49036 (N_49036,N_46437,N_46405);
and U49037 (N_49037,N_46256,N_47928);
nand U49038 (N_49038,N_47259,N_46841);
and U49039 (N_49039,N_47680,N_46865);
nor U49040 (N_49040,N_47693,N_47042);
and U49041 (N_49041,N_46099,N_47766);
and U49042 (N_49042,N_46425,N_47245);
nor U49043 (N_49043,N_46742,N_46294);
or U49044 (N_49044,N_46251,N_46016);
or U49045 (N_49045,N_46738,N_47702);
or U49046 (N_49046,N_47779,N_47169);
nand U49047 (N_49047,N_46831,N_47575);
and U49048 (N_49048,N_47030,N_47749);
nand U49049 (N_49049,N_47752,N_46907);
nand U49050 (N_49050,N_47587,N_47465);
xnor U49051 (N_49051,N_46784,N_47470);
nand U49052 (N_49052,N_46787,N_47203);
xor U49053 (N_49053,N_46374,N_47500);
nand U49054 (N_49054,N_47297,N_47906);
nor U49055 (N_49055,N_47155,N_46969);
nor U49056 (N_49056,N_46679,N_46960);
nand U49057 (N_49057,N_47724,N_47975);
or U49058 (N_49058,N_47909,N_46341);
or U49059 (N_49059,N_46842,N_47111);
nor U49060 (N_49060,N_47811,N_46214);
or U49061 (N_49061,N_46537,N_47711);
and U49062 (N_49062,N_46735,N_46919);
and U49063 (N_49063,N_46276,N_46835);
nor U49064 (N_49064,N_46283,N_46761);
or U49065 (N_49065,N_47833,N_46141);
or U49066 (N_49066,N_47904,N_46142);
nand U49067 (N_49067,N_46187,N_47258);
or U49068 (N_49068,N_47679,N_46646);
nand U49069 (N_49069,N_46032,N_47911);
or U49070 (N_49070,N_47222,N_47437);
and U49071 (N_49071,N_47704,N_47843);
and U49072 (N_49072,N_46740,N_47711);
or U49073 (N_49073,N_46597,N_47652);
and U49074 (N_49074,N_47396,N_46220);
xor U49075 (N_49075,N_47270,N_46673);
nor U49076 (N_49076,N_47593,N_47852);
and U49077 (N_49077,N_47288,N_47579);
or U49078 (N_49078,N_46898,N_47579);
or U49079 (N_49079,N_46485,N_47290);
nand U49080 (N_49080,N_46461,N_46837);
or U49081 (N_49081,N_46170,N_46469);
xor U49082 (N_49082,N_47937,N_46242);
or U49083 (N_49083,N_46601,N_47561);
or U49084 (N_49084,N_47225,N_46178);
nand U49085 (N_49085,N_47530,N_46187);
nor U49086 (N_49086,N_47995,N_47503);
xnor U49087 (N_49087,N_46953,N_46537);
nor U49088 (N_49088,N_47850,N_47160);
or U49089 (N_49089,N_47082,N_46708);
nor U49090 (N_49090,N_47962,N_47103);
xor U49091 (N_49091,N_46787,N_46428);
nor U49092 (N_49092,N_46412,N_46439);
nor U49093 (N_49093,N_46644,N_47480);
and U49094 (N_49094,N_46661,N_47782);
xor U49095 (N_49095,N_47109,N_47285);
nand U49096 (N_49096,N_47325,N_46812);
xor U49097 (N_49097,N_47554,N_46052);
nand U49098 (N_49098,N_47244,N_46143);
and U49099 (N_49099,N_47159,N_47659);
xnor U49100 (N_49100,N_46606,N_47423);
xnor U49101 (N_49101,N_47428,N_47687);
xor U49102 (N_49102,N_47007,N_46815);
or U49103 (N_49103,N_47344,N_46870);
nand U49104 (N_49104,N_46952,N_46471);
and U49105 (N_49105,N_47394,N_47033);
nand U49106 (N_49106,N_47716,N_47021);
or U49107 (N_49107,N_46053,N_46670);
and U49108 (N_49108,N_46734,N_46992);
and U49109 (N_49109,N_46755,N_47484);
nand U49110 (N_49110,N_47215,N_46286);
nand U49111 (N_49111,N_46569,N_46038);
or U49112 (N_49112,N_46431,N_47807);
nand U49113 (N_49113,N_46661,N_46468);
xor U49114 (N_49114,N_46227,N_47486);
xor U49115 (N_49115,N_46421,N_46661);
xnor U49116 (N_49116,N_47172,N_46739);
nand U49117 (N_49117,N_47851,N_46217);
or U49118 (N_49118,N_46270,N_47051);
xor U49119 (N_49119,N_47584,N_47640);
nand U49120 (N_49120,N_46355,N_47823);
nor U49121 (N_49121,N_47995,N_46003);
nor U49122 (N_49122,N_46661,N_47188);
nor U49123 (N_49123,N_46106,N_47816);
and U49124 (N_49124,N_47998,N_46621);
nor U49125 (N_49125,N_46649,N_46327);
nand U49126 (N_49126,N_47607,N_46300);
nand U49127 (N_49127,N_46245,N_46085);
and U49128 (N_49128,N_47998,N_47586);
or U49129 (N_49129,N_46988,N_46981);
xnor U49130 (N_49130,N_46090,N_46251);
xor U49131 (N_49131,N_46825,N_46875);
nand U49132 (N_49132,N_47631,N_47260);
nand U49133 (N_49133,N_46068,N_46803);
and U49134 (N_49134,N_46660,N_47258);
xnor U49135 (N_49135,N_46706,N_46559);
and U49136 (N_49136,N_46125,N_46392);
xor U49137 (N_49137,N_47840,N_46224);
nand U49138 (N_49138,N_47524,N_46910);
nand U49139 (N_49139,N_47890,N_46400);
xor U49140 (N_49140,N_47558,N_47432);
xnor U49141 (N_49141,N_46934,N_46068);
nand U49142 (N_49142,N_47812,N_46642);
xor U49143 (N_49143,N_47555,N_47748);
and U49144 (N_49144,N_47139,N_47658);
or U49145 (N_49145,N_46133,N_46658);
or U49146 (N_49146,N_47127,N_46594);
nor U49147 (N_49147,N_47550,N_46754);
xor U49148 (N_49148,N_46159,N_47753);
or U49149 (N_49149,N_46158,N_46692);
nand U49150 (N_49150,N_47656,N_47487);
nor U49151 (N_49151,N_46955,N_47845);
nand U49152 (N_49152,N_46172,N_47947);
xnor U49153 (N_49153,N_46995,N_47098);
nor U49154 (N_49154,N_47657,N_46565);
nand U49155 (N_49155,N_46960,N_46567);
nand U49156 (N_49156,N_47044,N_46520);
and U49157 (N_49157,N_47641,N_47366);
xor U49158 (N_49158,N_46097,N_46098);
nor U49159 (N_49159,N_46320,N_46582);
nor U49160 (N_49160,N_47192,N_46415);
and U49161 (N_49161,N_46048,N_47664);
or U49162 (N_49162,N_46489,N_46876);
and U49163 (N_49163,N_46441,N_46523);
and U49164 (N_49164,N_46600,N_47713);
and U49165 (N_49165,N_47920,N_46071);
xor U49166 (N_49166,N_47610,N_47707);
nor U49167 (N_49167,N_47029,N_47961);
or U49168 (N_49168,N_46950,N_46864);
xor U49169 (N_49169,N_46274,N_47185);
nand U49170 (N_49170,N_47417,N_46116);
and U49171 (N_49171,N_46772,N_46806);
nand U49172 (N_49172,N_47302,N_47379);
nand U49173 (N_49173,N_46649,N_46315);
nor U49174 (N_49174,N_46745,N_47381);
xor U49175 (N_49175,N_47974,N_47567);
nand U49176 (N_49176,N_46628,N_47556);
nor U49177 (N_49177,N_46839,N_47362);
nand U49178 (N_49178,N_47993,N_47908);
xnor U49179 (N_49179,N_46223,N_46697);
nor U49180 (N_49180,N_46897,N_46936);
nor U49181 (N_49181,N_47616,N_46782);
or U49182 (N_49182,N_46158,N_47315);
nand U49183 (N_49183,N_46789,N_47399);
nand U49184 (N_49184,N_47538,N_46135);
nor U49185 (N_49185,N_47107,N_47057);
xnor U49186 (N_49186,N_47460,N_46834);
and U49187 (N_49187,N_46203,N_46944);
and U49188 (N_49188,N_47797,N_47431);
or U49189 (N_49189,N_47514,N_46826);
nand U49190 (N_49190,N_47949,N_46220);
xnor U49191 (N_49191,N_47524,N_46294);
or U49192 (N_49192,N_46311,N_46775);
or U49193 (N_49193,N_46236,N_47288);
and U49194 (N_49194,N_46378,N_47883);
xnor U49195 (N_49195,N_46569,N_47298);
or U49196 (N_49196,N_46183,N_46622);
nor U49197 (N_49197,N_47485,N_46272);
nor U49198 (N_49198,N_46761,N_46865);
xor U49199 (N_49199,N_47408,N_47788);
and U49200 (N_49200,N_46365,N_47320);
xnor U49201 (N_49201,N_47794,N_46317);
nand U49202 (N_49202,N_46792,N_47171);
and U49203 (N_49203,N_47768,N_46851);
nor U49204 (N_49204,N_47891,N_46423);
or U49205 (N_49205,N_47941,N_46208);
nor U49206 (N_49206,N_46065,N_46542);
and U49207 (N_49207,N_46961,N_46072);
nand U49208 (N_49208,N_46293,N_47550);
or U49209 (N_49209,N_47914,N_47254);
and U49210 (N_49210,N_46881,N_46468);
nor U49211 (N_49211,N_46093,N_47660);
or U49212 (N_49212,N_47010,N_46324);
nor U49213 (N_49213,N_46439,N_46451);
or U49214 (N_49214,N_47193,N_46305);
and U49215 (N_49215,N_47945,N_46878);
and U49216 (N_49216,N_47945,N_47665);
xnor U49217 (N_49217,N_47510,N_46739);
nor U49218 (N_49218,N_46198,N_46004);
and U49219 (N_49219,N_47794,N_46585);
nor U49220 (N_49220,N_46291,N_47146);
nand U49221 (N_49221,N_47720,N_47499);
or U49222 (N_49222,N_47242,N_46079);
or U49223 (N_49223,N_46477,N_47965);
and U49224 (N_49224,N_46779,N_47304);
and U49225 (N_49225,N_46440,N_47119);
nor U49226 (N_49226,N_46894,N_47992);
and U49227 (N_49227,N_46428,N_47822);
xor U49228 (N_49228,N_47544,N_46098);
and U49229 (N_49229,N_47196,N_47078);
nor U49230 (N_49230,N_47003,N_47258);
or U49231 (N_49231,N_46415,N_46405);
or U49232 (N_49232,N_46358,N_46135);
and U49233 (N_49233,N_46945,N_47325);
nand U49234 (N_49234,N_47375,N_46777);
and U49235 (N_49235,N_46687,N_46789);
nor U49236 (N_49236,N_47503,N_46124);
nor U49237 (N_49237,N_46074,N_47963);
and U49238 (N_49238,N_47339,N_47727);
nor U49239 (N_49239,N_47060,N_47706);
xnor U49240 (N_49240,N_46645,N_47441);
xor U49241 (N_49241,N_47904,N_47751);
nor U49242 (N_49242,N_46073,N_47898);
nand U49243 (N_49243,N_46576,N_47490);
nand U49244 (N_49244,N_47589,N_46681);
nor U49245 (N_49245,N_47218,N_47668);
and U49246 (N_49246,N_46098,N_46961);
nor U49247 (N_49247,N_46816,N_46683);
or U49248 (N_49248,N_47529,N_47057);
or U49249 (N_49249,N_47905,N_47233);
xor U49250 (N_49250,N_46040,N_46243);
nor U49251 (N_49251,N_47185,N_47733);
nand U49252 (N_49252,N_46780,N_46858);
or U49253 (N_49253,N_46036,N_47985);
or U49254 (N_49254,N_47823,N_47464);
or U49255 (N_49255,N_47409,N_46722);
or U49256 (N_49256,N_47870,N_46064);
and U49257 (N_49257,N_46110,N_46615);
nand U49258 (N_49258,N_46432,N_46586);
or U49259 (N_49259,N_46597,N_47667);
nor U49260 (N_49260,N_47933,N_47744);
nor U49261 (N_49261,N_46935,N_46824);
and U49262 (N_49262,N_46624,N_47313);
or U49263 (N_49263,N_47309,N_46335);
and U49264 (N_49264,N_46841,N_46931);
xor U49265 (N_49265,N_46446,N_47989);
or U49266 (N_49266,N_47301,N_46717);
nor U49267 (N_49267,N_47158,N_47366);
nand U49268 (N_49268,N_47514,N_47516);
or U49269 (N_49269,N_46412,N_47568);
nand U49270 (N_49270,N_46175,N_46389);
nor U49271 (N_49271,N_47731,N_46726);
nor U49272 (N_49272,N_46434,N_47599);
nand U49273 (N_49273,N_47311,N_47386);
nand U49274 (N_49274,N_47191,N_46377);
or U49275 (N_49275,N_47017,N_46940);
or U49276 (N_49276,N_46422,N_46500);
xor U49277 (N_49277,N_47957,N_47074);
and U49278 (N_49278,N_47704,N_46444);
and U49279 (N_49279,N_47048,N_46353);
nand U49280 (N_49280,N_46630,N_47029);
nor U49281 (N_49281,N_46523,N_46432);
or U49282 (N_49282,N_47882,N_47287);
nand U49283 (N_49283,N_46603,N_47274);
xnor U49284 (N_49284,N_46544,N_47421);
xnor U49285 (N_49285,N_47577,N_47260);
or U49286 (N_49286,N_46340,N_47269);
nor U49287 (N_49287,N_46411,N_46658);
or U49288 (N_49288,N_46615,N_46417);
or U49289 (N_49289,N_46674,N_46684);
and U49290 (N_49290,N_46629,N_47217);
nand U49291 (N_49291,N_47679,N_47156);
or U49292 (N_49292,N_47841,N_46047);
nor U49293 (N_49293,N_47915,N_47445);
and U49294 (N_49294,N_46157,N_46626);
nor U49295 (N_49295,N_47704,N_47577);
nor U49296 (N_49296,N_46492,N_47300);
nor U49297 (N_49297,N_47739,N_47105);
nor U49298 (N_49298,N_47310,N_46600);
nor U49299 (N_49299,N_47748,N_46417);
or U49300 (N_49300,N_46351,N_46377);
nor U49301 (N_49301,N_47806,N_47614);
or U49302 (N_49302,N_46174,N_47617);
or U49303 (N_49303,N_46191,N_46689);
nor U49304 (N_49304,N_47179,N_46036);
and U49305 (N_49305,N_47294,N_46565);
nor U49306 (N_49306,N_47423,N_46859);
nand U49307 (N_49307,N_46606,N_46908);
nand U49308 (N_49308,N_47261,N_46243);
nor U49309 (N_49309,N_46202,N_46519);
nand U49310 (N_49310,N_46202,N_47145);
and U49311 (N_49311,N_46955,N_47894);
and U49312 (N_49312,N_46191,N_47947);
or U49313 (N_49313,N_46285,N_46910);
and U49314 (N_49314,N_47100,N_47411);
or U49315 (N_49315,N_46487,N_46952);
xnor U49316 (N_49316,N_46672,N_46960);
nor U49317 (N_49317,N_46261,N_47760);
nand U49318 (N_49318,N_47243,N_46485);
nand U49319 (N_49319,N_47571,N_46538);
nand U49320 (N_49320,N_46926,N_46941);
nand U49321 (N_49321,N_46754,N_46847);
xnor U49322 (N_49322,N_47385,N_46772);
nand U49323 (N_49323,N_47353,N_46419);
and U49324 (N_49324,N_46670,N_46485);
and U49325 (N_49325,N_47650,N_46223);
nor U49326 (N_49326,N_46801,N_47384);
xnor U49327 (N_49327,N_46576,N_47148);
xor U49328 (N_49328,N_47022,N_47883);
nor U49329 (N_49329,N_46027,N_46433);
or U49330 (N_49330,N_46531,N_46581);
nor U49331 (N_49331,N_46073,N_46576);
nor U49332 (N_49332,N_47467,N_47521);
nor U49333 (N_49333,N_46011,N_46213);
and U49334 (N_49334,N_46378,N_47039);
and U49335 (N_49335,N_47677,N_47363);
nor U49336 (N_49336,N_46577,N_47625);
and U49337 (N_49337,N_46999,N_47917);
nor U49338 (N_49338,N_46737,N_47959);
or U49339 (N_49339,N_46603,N_47765);
or U49340 (N_49340,N_46654,N_47652);
xnor U49341 (N_49341,N_46187,N_46207);
xnor U49342 (N_49342,N_47110,N_47034);
nor U49343 (N_49343,N_47506,N_47547);
or U49344 (N_49344,N_47352,N_47960);
and U49345 (N_49345,N_47163,N_46196);
and U49346 (N_49346,N_47580,N_46784);
xnor U49347 (N_49347,N_46609,N_47195);
xor U49348 (N_49348,N_47177,N_47392);
nor U49349 (N_49349,N_46388,N_47234);
or U49350 (N_49350,N_46200,N_47853);
nor U49351 (N_49351,N_46664,N_46393);
and U49352 (N_49352,N_47506,N_47251);
nor U49353 (N_49353,N_47781,N_46190);
nor U49354 (N_49354,N_47901,N_46356);
or U49355 (N_49355,N_47901,N_47256);
nand U49356 (N_49356,N_47586,N_46531);
nor U49357 (N_49357,N_47382,N_47113);
nor U49358 (N_49358,N_46736,N_46949);
or U49359 (N_49359,N_46604,N_47505);
and U49360 (N_49360,N_46757,N_47527);
xnor U49361 (N_49361,N_46528,N_47128);
or U49362 (N_49362,N_46096,N_46861);
or U49363 (N_49363,N_46435,N_46375);
nor U49364 (N_49364,N_47405,N_46029);
and U49365 (N_49365,N_47241,N_46655);
and U49366 (N_49366,N_47597,N_47944);
xnor U49367 (N_49367,N_46331,N_46211);
nor U49368 (N_49368,N_47384,N_46781);
xnor U49369 (N_49369,N_46708,N_47121);
nor U49370 (N_49370,N_47465,N_47093);
nand U49371 (N_49371,N_47443,N_47258);
or U49372 (N_49372,N_47078,N_47515);
nand U49373 (N_49373,N_46879,N_46591);
or U49374 (N_49374,N_47278,N_47817);
nand U49375 (N_49375,N_47141,N_46407);
and U49376 (N_49376,N_47594,N_47401);
nor U49377 (N_49377,N_46991,N_47771);
or U49378 (N_49378,N_47739,N_47365);
nand U49379 (N_49379,N_47037,N_46971);
nand U49380 (N_49380,N_47569,N_46338);
xnor U49381 (N_49381,N_46160,N_47704);
or U49382 (N_49382,N_46441,N_47834);
xnor U49383 (N_49383,N_46927,N_46136);
nor U49384 (N_49384,N_47932,N_47383);
or U49385 (N_49385,N_47167,N_47192);
nor U49386 (N_49386,N_47114,N_47988);
or U49387 (N_49387,N_46118,N_46671);
or U49388 (N_49388,N_47147,N_46790);
or U49389 (N_49389,N_47441,N_46055);
nand U49390 (N_49390,N_47129,N_46755);
and U49391 (N_49391,N_46723,N_46801);
or U49392 (N_49392,N_46847,N_47483);
xnor U49393 (N_49393,N_47782,N_46181);
nand U49394 (N_49394,N_46039,N_47909);
or U49395 (N_49395,N_46357,N_46257);
nor U49396 (N_49396,N_46529,N_46239);
nor U49397 (N_49397,N_46286,N_47477);
xor U49398 (N_49398,N_46138,N_47269);
xor U49399 (N_49399,N_47648,N_46435);
and U49400 (N_49400,N_46623,N_47913);
or U49401 (N_49401,N_47494,N_46562);
nor U49402 (N_49402,N_47690,N_46787);
xor U49403 (N_49403,N_46326,N_46026);
or U49404 (N_49404,N_46761,N_47067);
nand U49405 (N_49405,N_47552,N_47116);
and U49406 (N_49406,N_47338,N_47849);
xnor U49407 (N_49407,N_46245,N_47877);
xor U49408 (N_49408,N_46131,N_46055);
nor U49409 (N_49409,N_47544,N_47093);
or U49410 (N_49410,N_47643,N_46435);
nor U49411 (N_49411,N_47487,N_46158);
nor U49412 (N_49412,N_47097,N_46646);
and U49413 (N_49413,N_46945,N_46968);
and U49414 (N_49414,N_47680,N_47090);
or U49415 (N_49415,N_46075,N_46434);
nor U49416 (N_49416,N_46177,N_47569);
and U49417 (N_49417,N_47057,N_47708);
xnor U49418 (N_49418,N_47377,N_47178);
nand U49419 (N_49419,N_47766,N_46154);
nand U49420 (N_49420,N_47798,N_46133);
or U49421 (N_49421,N_47714,N_46149);
nor U49422 (N_49422,N_46140,N_47818);
or U49423 (N_49423,N_47997,N_47501);
nor U49424 (N_49424,N_47632,N_47450);
nor U49425 (N_49425,N_46318,N_47518);
nor U49426 (N_49426,N_46902,N_47861);
xnor U49427 (N_49427,N_47724,N_47955);
nand U49428 (N_49428,N_47607,N_46400);
or U49429 (N_49429,N_47746,N_47521);
and U49430 (N_49430,N_46747,N_46292);
xor U49431 (N_49431,N_46441,N_46905);
nand U49432 (N_49432,N_47872,N_46380);
nor U49433 (N_49433,N_47184,N_46769);
or U49434 (N_49434,N_47958,N_47014);
xor U49435 (N_49435,N_47298,N_46764);
or U49436 (N_49436,N_47153,N_46019);
nor U49437 (N_49437,N_47660,N_46772);
or U49438 (N_49438,N_47453,N_46815);
nor U49439 (N_49439,N_46016,N_46229);
nand U49440 (N_49440,N_47532,N_47592);
or U49441 (N_49441,N_47418,N_46354);
nor U49442 (N_49442,N_46423,N_46002);
and U49443 (N_49443,N_46803,N_46571);
and U49444 (N_49444,N_46904,N_46705);
xor U49445 (N_49445,N_46458,N_46422);
nor U49446 (N_49446,N_46499,N_46410);
and U49447 (N_49447,N_46187,N_46949);
xor U49448 (N_49448,N_47576,N_47991);
nand U49449 (N_49449,N_47683,N_46142);
xor U49450 (N_49450,N_46530,N_47485);
and U49451 (N_49451,N_47495,N_47869);
or U49452 (N_49452,N_47330,N_47509);
or U49453 (N_49453,N_46037,N_47300);
xor U49454 (N_49454,N_47527,N_47141);
or U49455 (N_49455,N_46176,N_46458);
nand U49456 (N_49456,N_46107,N_46374);
nand U49457 (N_49457,N_46956,N_47968);
and U49458 (N_49458,N_46693,N_46827);
xor U49459 (N_49459,N_46155,N_46303);
and U49460 (N_49460,N_47453,N_47208);
nor U49461 (N_49461,N_47136,N_46664);
nand U49462 (N_49462,N_47092,N_47386);
xor U49463 (N_49463,N_46612,N_46281);
nor U49464 (N_49464,N_46532,N_46460);
and U49465 (N_49465,N_46639,N_47738);
and U49466 (N_49466,N_47908,N_47332);
or U49467 (N_49467,N_46958,N_46955);
or U49468 (N_49468,N_46151,N_46605);
nand U49469 (N_49469,N_46706,N_47772);
and U49470 (N_49470,N_47504,N_47877);
nand U49471 (N_49471,N_47140,N_47150);
xnor U49472 (N_49472,N_47566,N_47499);
xor U49473 (N_49473,N_47560,N_46426);
nand U49474 (N_49474,N_46204,N_47921);
and U49475 (N_49475,N_47759,N_46571);
nor U49476 (N_49476,N_46973,N_47422);
xor U49477 (N_49477,N_46681,N_46137);
and U49478 (N_49478,N_47121,N_47674);
nor U49479 (N_49479,N_47319,N_46551);
nand U49480 (N_49480,N_47026,N_47318);
nor U49481 (N_49481,N_47031,N_47355);
or U49482 (N_49482,N_47947,N_47692);
nand U49483 (N_49483,N_47378,N_46485);
nor U49484 (N_49484,N_47777,N_47193);
and U49485 (N_49485,N_46702,N_47774);
or U49486 (N_49486,N_46989,N_46806);
nor U49487 (N_49487,N_46503,N_46258);
or U49488 (N_49488,N_47090,N_46428);
xnor U49489 (N_49489,N_47934,N_46393);
xor U49490 (N_49490,N_46128,N_46586);
nor U49491 (N_49491,N_47864,N_47379);
nor U49492 (N_49492,N_46445,N_47895);
or U49493 (N_49493,N_47361,N_47832);
or U49494 (N_49494,N_46235,N_47179);
xnor U49495 (N_49495,N_46352,N_47819);
or U49496 (N_49496,N_47811,N_47030);
or U49497 (N_49497,N_47953,N_46671);
nand U49498 (N_49498,N_46280,N_46609);
or U49499 (N_49499,N_47873,N_47368);
nand U49500 (N_49500,N_46855,N_46592);
nor U49501 (N_49501,N_47658,N_47065);
xnor U49502 (N_49502,N_46006,N_47695);
nor U49503 (N_49503,N_46232,N_46430);
xor U49504 (N_49504,N_46358,N_46025);
nand U49505 (N_49505,N_46981,N_46257);
nand U49506 (N_49506,N_47803,N_47111);
xor U49507 (N_49507,N_47418,N_46200);
and U49508 (N_49508,N_47224,N_46224);
nor U49509 (N_49509,N_46238,N_47343);
and U49510 (N_49510,N_46705,N_47323);
nor U49511 (N_49511,N_47538,N_46807);
xor U49512 (N_49512,N_46438,N_46220);
and U49513 (N_49513,N_46709,N_47135);
and U49514 (N_49514,N_47160,N_46332);
nor U49515 (N_49515,N_47911,N_46619);
or U49516 (N_49516,N_46539,N_47254);
nand U49517 (N_49517,N_46624,N_47742);
and U49518 (N_49518,N_47813,N_46532);
nor U49519 (N_49519,N_46328,N_47149);
and U49520 (N_49520,N_47578,N_46284);
or U49521 (N_49521,N_46081,N_47873);
xnor U49522 (N_49522,N_46419,N_47123);
xor U49523 (N_49523,N_47259,N_46120);
xnor U49524 (N_49524,N_46076,N_46090);
xor U49525 (N_49525,N_47129,N_47206);
xor U49526 (N_49526,N_47416,N_47688);
nor U49527 (N_49527,N_47435,N_47528);
and U49528 (N_49528,N_47473,N_46721);
xor U49529 (N_49529,N_47113,N_46075);
nor U49530 (N_49530,N_46734,N_46311);
xor U49531 (N_49531,N_47334,N_47692);
xnor U49532 (N_49532,N_46647,N_46512);
and U49533 (N_49533,N_47454,N_46886);
or U49534 (N_49534,N_47057,N_46831);
xnor U49535 (N_49535,N_47228,N_47919);
and U49536 (N_49536,N_47619,N_46765);
xor U49537 (N_49537,N_47170,N_46796);
or U49538 (N_49538,N_46496,N_47701);
and U49539 (N_49539,N_47112,N_47926);
nand U49540 (N_49540,N_47349,N_46535);
or U49541 (N_49541,N_47091,N_46730);
nor U49542 (N_49542,N_47490,N_47553);
or U49543 (N_49543,N_47894,N_47506);
and U49544 (N_49544,N_46537,N_46055);
nor U49545 (N_49545,N_47477,N_47905);
and U49546 (N_49546,N_46606,N_46104);
nor U49547 (N_49547,N_47142,N_47404);
nor U49548 (N_49548,N_47321,N_47656);
or U49549 (N_49549,N_47836,N_47848);
and U49550 (N_49550,N_46439,N_47190);
or U49551 (N_49551,N_46495,N_46546);
nor U49552 (N_49552,N_46704,N_47035);
xnor U49553 (N_49553,N_47941,N_47264);
and U49554 (N_49554,N_47779,N_47386);
and U49555 (N_49555,N_47026,N_47878);
or U49556 (N_49556,N_47339,N_47683);
nand U49557 (N_49557,N_47273,N_46965);
xor U49558 (N_49558,N_46927,N_46919);
xor U49559 (N_49559,N_47729,N_47632);
xor U49560 (N_49560,N_47067,N_46042);
nand U49561 (N_49561,N_47138,N_46511);
xor U49562 (N_49562,N_46767,N_47004);
and U49563 (N_49563,N_47710,N_46377);
and U49564 (N_49564,N_47410,N_46797);
nand U49565 (N_49565,N_46588,N_46875);
and U49566 (N_49566,N_47129,N_47727);
nand U49567 (N_49567,N_46159,N_46255);
nand U49568 (N_49568,N_46072,N_47956);
and U49569 (N_49569,N_47795,N_47076);
xnor U49570 (N_49570,N_46517,N_47631);
and U49571 (N_49571,N_47027,N_46391);
nor U49572 (N_49572,N_47374,N_47835);
or U49573 (N_49573,N_47459,N_47543);
xor U49574 (N_49574,N_46274,N_46490);
and U49575 (N_49575,N_47044,N_47582);
or U49576 (N_49576,N_47291,N_47930);
and U49577 (N_49577,N_47131,N_46970);
nor U49578 (N_49578,N_47546,N_47273);
nand U49579 (N_49579,N_46647,N_47083);
xor U49580 (N_49580,N_47622,N_47837);
or U49581 (N_49581,N_46796,N_46532);
or U49582 (N_49582,N_47018,N_47089);
nand U49583 (N_49583,N_46763,N_47358);
nand U49584 (N_49584,N_47126,N_47752);
and U49585 (N_49585,N_47766,N_46334);
nand U49586 (N_49586,N_47947,N_46210);
nand U49587 (N_49587,N_47531,N_46980);
or U49588 (N_49588,N_46231,N_46178);
nor U49589 (N_49589,N_46427,N_47530);
nand U49590 (N_49590,N_46478,N_47664);
nand U49591 (N_49591,N_47322,N_47862);
nor U49592 (N_49592,N_46405,N_47420);
nor U49593 (N_49593,N_47148,N_47256);
xor U49594 (N_49594,N_46545,N_46048);
nor U49595 (N_49595,N_46549,N_47311);
or U49596 (N_49596,N_46121,N_47097);
xnor U49597 (N_49597,N_46923,N_47098);
xnor U49598 (N_49598,N_46377,N_47776);
nor U49599 (N_49599,N_46560,N_47623);
or U49600 (N_49600,N_46980,N_46209);
or U49601 (N_49601,N_47939,N_47229);
nor U49602 (N_49602,N_46541,N_46318);
or U49603 (N_49603,N_47791,N_47334);
xor U49604 (N_49604,N_46554,N_46011);
nand U49605 (N_49605,N_46296,N_47897);
nand U49606 (N_49606,N_47822,N_46152);
or U49607 (N_49607,N_47286,N_46202);
or U49608 (N_49608,N_46408,N_46567);
and U49609 (N_49609,N_47238,N_46398);
nand U49610 (N_49610,N_47062,N_47631);
nor U49611 (N_49611,N_46314,N_46659);
nand U49612 (N_49612,N_46675,N_47148);
nand U49613 (N_49613,N_47120,N_46262);
nor U49614 (N_49614,N_47878,N_47656);
xnor U49615 (N_49615,N_46239,N_47897);
or U49616 (N_49616,N_47378,N_47068);
nor U49617 (N_49617,N_47937,N_47361);
nor U49618 (N_49618,N_47838,N_46508);
or U49619 (N_49619,N_46644,N_46684);
or U49620 (N_49620,N_46981,N_46944);
or U49621 (N_49621,N_46893,N_47972);
or U49622 (N_49622,N_47870,N_46806);
nand U49623 (N_49623,N_47513,N_46066);
and U49624 (N_49624,N_47939,N_46444);
nor U49625 (N_49625,N_47189,N_47977);
or U49626 (N_49626,N_46072,N_47819);
xnor U49627 (N_49627,N_46489,N_46922);
nand U49628 (N_49628,N_46195,N_47423);
nor U49629 (N_49629,N_47949,N_46649);
nand U49630 (N_49630,N_46074,N_46350);
xnor U49631 (N_49631,N_46932,N_47065);
or U49632 (N_49632,N_47598,N_46779);
and U49633 (N_49633,N_46143,N_46750);
nor U49634 (N_49634,N_46400,N_46286);
nor U49635 (N_49635,N_46283,N_46070);
or U49636 (N_49636,N_47572,N_46635);
and U49637 (N_49637,N_47724,N_47530);
or U49638 (N_49638,N_46347,N_46678);
nor U49639 (N_49639,N_46865,N_46498);
and U49640 (N_49640,N_46068,N_47250);
xnor U49641 (N_49641,N_46908,N_46667);
and U49642 (N_49642,N_47543,N_46424);
or U49643 (N_49643,N_46848,N_46132);
nand U49644 (N_49644,N_46526,N_47645);
or U49645 (N_49645,N_47916,N_47718);
nor U49646 (N_49646,N_46320,N_47162);
nand U49647 (N_49647,N_46031,N_46099);
and U49648 (N_49648,N_46209,N_47566);
nor U49649 (N_49649,N_46493,N_47784);
xor U49650 (N_49650,N_47351,N_46019);
nor U49651 (N_49651,N_47162,N_46268);
nand U49652 (N_49652,N_46092,N_47569);
nor U49653 (N_49653,N_47100,N_46000);
nor U49654 (N_49654,N_46169,N_46749);
and U49655 (N_49655,N_47798,N_47789);
nand U49656 (N_49656,N_47095,N_47892);
or U49657 (N_49657,N_46812,N_47512);
nor U49658 (N_49658,N_47962,N_47077);
and U49659 (N_49659,N_46866,N_46056);
nand U49660 (N_49660,N_46276,N_47548);
and U49661 (N_49661,N_46569,N_46587);
and U49662 (N_49662,N_47039,N_46043);
or U49663 (N_49663,N_46888,N_46357);
and U49664 (N_49664,N_46727,N_47362);
nand U49665 (N_49665,N_46016,N_47377);
nor U49666 (N_49666,N_47117,N_46552);
nand U49667 (N_49667,N_47440,N_47218);
and U49668 (N_49668,N_47570,N_46654);
nor U49669 (N_49669,N_47647,N_46199);
nor U49670 (N_49670,N_47575,N_46197);
xor U49671 (N_49671,N_46056,N_47399);
nor U49672 (N_49672,N_47640,N_47172);
and U49673 (N_49673,N_47107,N_46442);
and U49674 (N_49674,N_47175,N_47405);
and U49675 (N_49675,N_46757,N_47548);
or U49676 (N_49676,N_47598,N_47160);
xor U49677 (N_49677,N_46221,N_46055);
nor U49678 (N_49678,N_46580,N_47177);
xor U49679 (N_49679,N_46592,N_46702);
or U49680 (N_49680,N_46872,N_46294);
and U49681 (N_49681,N_46536,N_46443);
and U49682 (N_49682,N_47819,N_47731);
and U49683 (N_49683,N_46664,N_47264);
nand U49684 (N_49684,N_47869,N_47302);
or U49685 (N_49685,N_47945,N_46204);
nor U49686 (N_49686,N_46507,N_47158);
nand U49687 (N_49687,N_47156,N_47840);
nor U49688 (N_49688,N_46560,N_47895);
or U49689 (N_49689,N_46725,N_46926);
nand U49690 (N_49690,N_46356,N_47540);
or U49691 (N_49691,N_46559,N_46662);
xnor U49692 (N_49692,N_46641,N_47271);
and U49693 (N_49693,N_46096,N_46412);
nand U49694 (N_49694,N_46228,N_46167);
or U49695 (N_49695,N_46671,N_47490);
and U49696 (N_49696,N_47679,N_46754);
and U49697 (N_49697,N_46420,N_47963);
xnor U49698 (N_49698,N_47711,N_46856);
nand U49699 (N_49699,N_47753,N_46063);
nor U49700 (N_49700,N_47078,N_47493);
nor U49701 (N_49701,N_47156,N_47761);
or U49702 (N_49702,N_46900,N_46154);
xor U49703 (N_49703,N_47967,N_47564);
or U49704 (N_49704,N_46312,N_47702);
nor U49705 (N_49705,N_47208,N_47093);
or U49706 (N_49706,N_47894,N_47626);
xnor U49707 (N_49707,N_46932,N_46387);
xnor U49708 (N_49708,N_46557,N_46780);
nor U49709 (N_49709,N_46537,N_46358);
and U49710 (N_49710,N_46318,N_47006);
nor U49711 (N_49711,N_47724,N_46115);
nand U49712 (N_49712,N_47768,N_46587);
nand U49713 (N_49713,N_47330,N_46626);
and U49714 (N_49714,N_46274,N_46638);
xor U49715 (N_49715,N_46776,N_46015);
or U49716 (N_49716,N_47067,N_46052);
xor U49717 (N_49717,N_46676,N_47513);
nand U49718 (N_49718,N_47785,N_47752);
nor U49719 (N_49719,N_46518,N_46383);
and U49720 (N_49720,N_47867,N_47916);
and U49721 (N_49721,N_47993,N_46603);
nor U49722 (N_49722,N_46367,N_46377);
xnor U49723 (N_49723,N_46475,N_46588);
or U49724 (N_49724,N_46896,N_47745);
and U49725 (N_49725,N_46352,N_46833);
and U49726 (N_49726,N_47169,N_47125);
nand U49727 (N_49727,N_46969,N_47878);
nand U49728 (N_49728,N_47952,N_46382);
nor U49729 (N_49729,N_46909,N_47411);
nand U49730 (N_49730,N_47769,N_47384);
and U49731 (N_49731,N_47508,N_46048);
nand U49732 (N_49732,N_46077,N_47996);
or U49733 (N_49733,N_47574,N_47903);
xnor U49734 (N_49734,N_47195,N_46088);
nand U49735 (N_49735,N_47931,N_47032);
nand U49736 (N_49736,N_47697,N_46338);
xor U49737 (N_49737,N_46243,N_46752);
xor U49738 (N_49738,N_46338,N_47627);
and U49739 (N_49739,N_46048,N_47600);
and U49740 (N_49740,N_47007,N_46465);
or U49741 (N_49741,N_46269,N_47194);
nand U49742 (N_49742,N_47326,N_47432);
nand U49743 (N_49743,N_46890,N_46780);
xor U49744 (N_49744,N_46467,N_46634);
nand U49745 (N_49745,N_46682,N_47854);
nor U49746 (N_49746,N_47756,N_47287);
nor U49747 (N_49747,N_47163,N_46896);
and U49748 (N_49748,N_47721,N_46606);
nor U49749 (N_49749,N_47353,N_46822);
nor U49750 (N_49750,N_46062,N_46345);
and U49751 (N_49751,N_46398,N_46672);
nand U49752 (N_49752,N_46609,N_47990);
and U49753 (N_49753,N_46136,N_46882);
nand U49754 (N_49754,N_47847,N_47419);
and U49755 (N_49755,N_46410,N_47863);
or U49756 (N_49756,N_47454,N_47636);
nand U49757 (N_49757,N_46156,N_46643);
nand U49758 (N_49758,N_47129,N_46534);
nor U49759 (N_49759,N_47117,N_46613);
nor U49760 (N_49760,N_46083,N_46682);
nor U49761 (N_49761,N_47088,N_46053);
nor U49762 (N_49762,N_46843,N_46754);
xor U49763 (N_49763,N_47176,N_46027);
or U49764 (N_49764,N_47673,N_46531);
or U49765 (N_49765,N_47340,N_46557);
or U49766 (N_49766,N_47227,N_47352);
and U49767 (N_49767,N_47827,N_46998);
and U49768 (N_49768,N_47296,N_46473);
xnor U49769 (N_49769,N_47504,N_46665);
nand U49770 (N_49770,N_46866,N_47175);
or U49771 (N_49771,N_47000,N_46742);
and U49772 (N_49772,N_46740,N_46945);
nor U49773 (N_49773,N_47932,N_47192);
nand U49774 (N_49774,N_46669,N_47693);
or U49775 (N_49775,N_47159,N_46120);
nand U49776 (N_49776,N_47012,N_46247);
xor U49777 (N_49777,N_46339,N_46081);
nand U49778 (N_49778,N_46822,N_47877);
xor U49779 (N_49779,N_47240,N_47152);
xor U49780 (N_49780,N_47221,N_47588);
xnor U49781 (N_49781,N_46956,N_47305);
nand U49782 (N_49782,N_47209,N_47861);
and U49783 (N_49783,N_46581,N_46681);
nor U49784 (N_49784,N_47413,N_47724);
nor U49785 (N_49785,N_47261,N_47502);
nor U49786 (N_49786,N_46371,N_46265);
and U49787 (N_49787,N_46188,N_46012);
xnor U49788 (N_49788,N_46673,N_47032);
nand U49789 (N_49789,N_47476,N_47741);
or U49790 (N_49790,N_46353,N_47496);
xor U49791 (N_49791,N_47701,N_47521);
xnor U49792 (N_49792,N_47394,N_46352);
xor U49793 (N_49793,N_47033,N_46866);
or U49794 (N_49794,N_46553,N_47315);
nor U49795 (N_49795,N_47555,N_46809);
nor U49796 (N_49796,N_46401,N_47904);
and U49797 (N_49797,N_46861,N_47719);
nand U49798 (N_49798,N_47169,N_46671);
and U49799 (N_49799,N_47227,N_47057);
or U49800 (N_49800,N_47311,N_46989);
and U49801 (N_49801,N_46568,N_46426);
xnor U49802 (N_49802,N_47242,N_46597);
nand U49803 (N_49803,N_47693,N_46789);
nor U49804 (N_49804,N_46910,N_46128);
or U49805 (N_49805,N_46543,N_47914);
or U49806 (N_49806,N_46334,N_47945);
xor U49807 (N_49807,N_46268,N_47415);
xor U49808 (N_49808,N_46797,N_47468);
and U49809 (N_49809,N_46307,N_46913);
xor U49810 (N_49810,N_46142,N_47894);
nand U49811 (N_49811,N_46842,N_47491);
and U49812 (N_49812,N_46054,N_47633);
xor U49813 (N_49813,N_46101,N_46485);
xnor U49814 (N_49814,N_46676,N_47695);
nand U49815 (N_49815,N_47182,N_47691);
or U49816 (N_49816,N_46016,N_46442);
xor U49817 (N_49817,N_47160,N_47781);
xnor U49818 (N_49818,N_46109,N_47747);
and U49819 (N_49819,N_47249,N_47227);
xnor U49820 (N_49820,N_46925,N_46684);
and U49821 (N_49821,N_46236,N_46327);
or U49822 (N_49822,N_46637,N_46670);
nor U49823 (N_49823,N_47398,N_46818);
and U49824 (N_49824,N_46283,N_46791);
xor U49825 (N_49825,N_47916,N_46284);
or U49826 (N_49826,N_47035,N_47280);
and U49827 (N_49827,N_47996,N_46692);
and U49828 (N_49828,N_47514,N_46952);
xnor U49829 (N_49829,N_46499,N_46189);
or U49830 (N_49830,N_46354,N_46285);
xnor U49831 (N_49831,N_47915,N_47417);
and U49832 (N_49832,N_47473,N_46246);
xor U49833 (N_49833,N_46596,N_46406);
xor U49834 (N_49834,N_47923,N_47243);
xor U49835 (N_49835,N_47725,N_46811);
or U49836 (N_49836,N_47255,N_46808);
nor U49837 (N_49837,N_47582,N_46894);
and U49838 (N_49838,N_46302,N_46571);
nor U49839 (N_49839,N_46797,N_46776);
or U49840 (N_49840,N_46352,N_47380);
and U49841 (N_49841,N_47408,N_46782);
nor U49842 (N_49842,N_46870,N_46930);
or U49843 (N_49843,N_47774,N_47162);
nand U49844 (N_49844,N_46520,N_47155);
xor U49845 (N_49845,N_46663,N_47499);
nand U49846 (N_49846,N_47157,N_47989);
or U49847 (N_49847,N_47097,N_47591);
xor U49848 (N_49848,N_46218,N_47050);
and U49849 (N_49849,N_47557,N_46403);
nand U49850 (N_49850,N_46689,N_46150);
xnor U49851 (N_49851,N_46119,N_47785);
nand U49852 (N_49852,N_47757,N_47314);
nand U49853 (N_49853,N_46308,N_46918);
or U49854 (N_49854,N_47008,N_47569);
or U49855 (N_49855,N_46276,N_46448);
nand U49856 (N_49856,N_47851,N_46932);
or U49857 (N_49857,N_46893,N_46321);
or U49858 (N_49858,N_47293,N_47284);
nor U49859 (N_49859,N_47464,N_47214);
nor U49860 (N_49860,N_46946,N_47075);
and U49861 (N_49861,N_47737,N_47368);
nand U49862 (N_49862,N_47720,N_47505);
xnor U49863 (N_49863,N_47564,N_47713);
nand U49864 (N_49864,N_46043,N_46554);
or U49865 (N_49865,N_47383,N_46106);
nor U49866 (N_49866,N_46257,N_47377);
or U49867 (N_49867,N_47684,N_47973);
or U49868 (N_49868,N_47045,N_47252);
or U49869 (N_49869,N_47333,N_47554);
and U49870 (N_49870,N_47837,N_47117);
or U49871 (N_49871,N_47618,N_46899);
nand U49872 (N_49872,N_46284,N_47759);
and U49873 (N_49873,N_46483,N_47746);
or U49874 (N_49874,N_47528,N_47465);
nor U49875 (N_49875,N_47352,N_47699);
nand U49876 (N_49876,N_47898,N_46037);
or U49877 (N_49877,N_46540,N_46793);
and U49878 (N_49878,N_46842,N_47392);
nand U49879 (N_49879,N_47654,N_47566);
xnor U49880 (N_49880,N_47555,N_46213);
and U49881 (N_49881,N_46571,N_47911);
and U49882 (N_49882,N_46883,N_47428);
nand U49883 (N_49883,N_47205,N_46452);
xnor U49884 (N_49884,N_47676,N_46183);
xnor U49885 (N_49885,N_47285,N_46549);
nor U49886 (N_49886,N_46933,N_46847);
or U49887 (N_49887,N_47642,N_47628);
nor U49888 (N_49888,N_46309,N_46103);
or U49889 (N_49889,N_47594,N_46949);
or U49890 (N_49890,N_46860,N_47848);
and U49891 (N_49891,N_46482,N_46368);
nand U49892 (N_49892,N_46616,N_47569);
nor U49893 (N_49893,N_47639,N_46068);
or U49894 (N_49894,N_47559,N_47384);
nand U49895 (N_49895,N_46229,N_46448);
and U49896 (N_49896,N_47612,N_47368);
nand U49897 (N_49897,N_46291,N_47029);
nor U49898 (N_49898,N_46419,N_47094);
xnor U49899 (N_49899,N_47169,N_46851);
and U49900 (N_49900,N_46753,N_46983);
or U49901 (N_49901,N_46325,N_47354);
xor U49902 (N_49902,N_46481,N_47364);
and U49903 (N_49903,N_47108,N_47081);
or U49904 (N_49904,N_46137,N_47792);
nor U49905 (N_49905,N_46531,N_46384);
and U49906 (N_49906,N_47436,N_47539);
and U49907 (N_49907,N_46380,N_47751);
nand U49908 (N_49908,N_47199,N_47553);
xnor U49909 (N_49909,N_47846,N_46841);
nand U49910 (N_49910,N_46585,N_47892);
xnor U49911 (N_49911,N_46309,N_47381);
or U49912 (N_49912,N_46254,N_46991);
or U49913 (N_49913,N_47950,N_47733);
nand U49914 (N_49914,N_47062,N_47298);
xor U49915 (N_49915,N_46917,N_46641);
nor U49916 (N_49916,N_47091,N_46759);
nor U49917 (N_49917,N_47607,N_47421);
or U49918 (N_49918,N_46519,N_47994);
nor U49919 (N_49919,N_46726,N_47092);
and U49920 (N_49920,N_47119,N_46781);
nor U49921 (N_49921,N_46815,N_47131);
nor U49922 (N_49922,N_47184,N_47258);
nor U49923 (N_49923,N_47393,N_47486);
or U49924 (N_49924,N_46048,N_46109);
and U49925 (N_49925,N_47163,N_46484);
or U49926 (N_49926,N_46831,N_46845);
nand U49927 (N_49927,N_47346,N_47415);
and U49928 (N_49928,N_47517,N_47792);
and U49929 (N_49929,N_46866,N_46040);
nor U49930 (N_49930,N_46634,N_46977);
xnor U49931 (N_49931,N_47891,N_47746);
or U49932 (N_49932,N_46293,N_47496);
nor U49933 (N_49933,N_47513,N_46329);
and U49934 (N_49934,N_47815,N_46604);
xnor U49935 (N_49935,N_47252,N_46611);
nand U49936 (N_49936,N_47597,N_46157);
xnor U49937 (N_49937,N_47621,N_46236);
or U49938 (N_49938,N_46016,N_47146);
or U49939 (N_49939,N_46522,N_46069);
and U49940 (N_49940,N_47266,N_47510);
and U49941 (N_49941,N_47139,N_46612);
or U49942 (N_49942,N_47606,N_47850);
and U49943 (N_49943,N_47117,N_46786);
and U49944 (N_49944,N_46764,N_46173);
nand U49945 (N_49945,N_46579,N_46343);
and U49946 (N_49946,N_47018,N_46103);
and U49947 (N_49947,N_46419,N_46629);
or U49948 (N_49948,N_46578,N_46257);
and U49949 (N_49949,N_46702,N_46764);
nand U49950 (N_49950,N_47238,N_46220);
nor U49951 (N_49951,N_47093,N_47484);
nor U49952 (N_49952,N_47388,N_47881);
xor U49953 (N_49953,N_46740,N_46503);
or U49954 (N_49954,N_47143,N_46996);
or U49955 (N_49955,N_47158,N_46307);
and U49956 (N_49956,N_47901,N_46996);
nor U49957 (N_49957,N_47838,N_46253);
xor U49958 (N_49958,N_46810,N_47596);
and U49959 (N_49959,N_46402,N_46642);
and U49960 (N_49960,N_47195,N_47595);
or U49961 (N_49961,N_47103,N_47918);
nor U49962 (N_49962,N_46952,N_46071);
xnor U49963 (N_49963,N_47056,N_47897);
nand U49964 (N_49964,N_47664,N_47504);
nand U49965 (N_49965,N_47151,N_47660);
and U49966 (N_49966,N_46805,N_47459);
or U49967 (N_49967,N_47533,N_46837);
xnor U49968 (N_49968,N_46657,N_46014);
xnor U49969 (N_49969,N_46174,N_47014);
and U49970 (N_49970,N_47324,N_46326);
nor U49971 (N_49971,N_46509,N_46874);
or U49972 (N_49972,N_47612,N_47031);
or U49973 (N_49973,N_47458,N_46450);
or U49974 (N_49974,N_46359,N_46356);
nor U49975 (N_49975,N_46176,N_47825);
xnor U49976 (N_49976,N_46758,N_46667);
xnor U49977 (N_49977,N_46382,N_46504);
nand U49978 (N_49978,N_46452,N_47411);
or U49979 (N_49979,N_46178,N_46373);
nand U49980 (N_49980,N_46666,N_46468);
and U49981 (N_49981,N_46504,N_47721);
xnor U49982 (N_49982,N_47746,N_46850);
nand U49983 (N_49983,N_47585,N_46802);
and U49984 (N_49984,N_47207,N_47775);
nor U49985 (N_49985,N_47963,N_47985);
nor U49986 (N_49986,N_47803,N_46628);
xnor U49987 (N_49987,N_47736,N_47546);
nand U49988 (N_49988,N_47134,N_46289);
nor U49989 (N_49989,N_47995,N_47762);
and U49990 (N_49990,N_46752,N_46728);
nor U49991 (N_49991,N_47667,N_47733);
nor U49992 (N_49992,N_47566,N_46736);
nor U49993 (N_49993,N_47415,N_47229);
or U49994 (N_49994,N_47947,N_47324);
xor U49995 (N_49995,N_46580,N_46235);
or U49996 (N_49996,N_46154,N_47219);
nor U49997 (N_49997,N_47556,N_46564);
and U49998 (N_49998,N_47062,N_47376);
and U49999 (N_49999,N_46236,N_46533);
nor UO_0 (O_0,N_48636,N_49787);
and UO_1 (O_1,N_49749,N_49444);
and UO_2 (O_2,N_49562,N_49069);
or UO_3 (O_3,N_49360,N_49619);
or UO_4 (O_4,N_49384,N_49366);
nor UO_5 (O_5,N_48971,N_49648);
or UO_6 (O_6,N_49371,N_49029);
xnor UO_7 (O_7,N_48118,N_48615);
nor UO_8 (O_8,N_48890,N_48722);
nand UO_9 (O_9,N_49299,N_49599);
and UO_10 (O_10,N_49842,N_49095);
and UO_11 (O_11,N_49850,N_48016);
nand UO_12 (O_12,N_48338,N_49829);
and UO_13 (O_13,N_48641,N_49542);
xor UO_14 (O_14,N_49779,N_49194);
or UO_15 (O_15,N_48965,N_49965);
and UO_16 (O_16,N_48117,N_48024);
or UO_17 (O_17,N_48047,N_48483);
nand UO_18 (O_18,N_48484,N_49598);
xor UO_19 (O_19,N_49810,N_49730);
or UO_20 (O_20,N_49313,N_49783);
nand UO_21 (O_21,N_49034,N_49953);
and UO_22 (O_22,N_49644,N_48838);
nor UO_23 (O_23,N_48967,N_49685);
and UO_24 (O_24,N_49691,N_48089);
and UO_25 (O_25,N_49778,N_49800);
nand UO_26 (O_26,N_48699,N_48240);
and UO_27 (O_27,N_49132,N_49245);
or UO_28 (O_28,N_48646,N_48752);
and UO_29 (O_29,N_49884,N_48873);
or UO_30 (O_30,N_49792,N_49474);
xnor UO_31 (O_31,N_49471,N_49250);
or UO_32 (O_32,N_49001,N_48523);
xor UO_33 (O_33,N_49498,N_48499);
and UO_34 (O_34,N_49586,N_48195);
nor UO_35 (O_35,N_49834,N_49646);
nor UO_36 (O_36,N_48329,N_48356);
nand UO_37 (O_37,N_48554,N_48177);
and UO_38 (O_38,N_49900,N_49895);
nand UO_39 (O_39,N_48757,N_48001);
and UO_40 (O_40,N_48015,N_48389);
nand UO_41 (O_41,N_49093,N_49486);
xnor UO_42 (O_42,N_48468,N_49566);
and UO_43 (O_43,N_48900,N_48938);
nand UO_44 (O_44,N_49941,N_49460);
nor UO_45 (O_45,N_48798,N_48827);
or UO_46 (O_46,N_49237,N_48303);
nand UO_47 (O_47,N_49359,N_48841);
nand UO_48 (O_48,N_49382,N_49883);
nor UO_49 (O_49,N_48559,N_49665);
or UO_50 (O_50,N_49153,N_49113);
and UO_51 (O_51,N_48272,N_49048);
nor UO_52 (O_52,N_48660,N_49228);
or UO_53 (O_53,N_48341,N_48916);
nor UO_54 (O_54,N_49833,N_49706);
nor UO_55 (O_55,N_48004,N_49750);
nor UO_56 (O_56,N_49671,N_49137);
nor UO_57 (O_57,N_49441,N_48300);
nor UO_58 (O_58,N_48951,N_48179);
xnor UO_59 (O_59,N_48534,N_48365);
xnor UO_60 (O_60,N_49826,N_48745);
and UO_61 (O_61,N_49183,N_49812);
nand UO_62 (O_62,N_49236,N_48350);
and UO_63 (O_63,N_49933,N_48762);
xor UO_64 (O_64,N_48183,N_48302);
nand UO_65 (O_65,N_48562,N_48498);
nand UO_66 (O_66,N_49035,N_48934);
xnor UO_67 (O_67,N_49744,N_49535);
nor UO_68 (O_68,N_49006,N_49369);
xnor UO_69 (O_69,N_49929,N_49672);
nor UO_70 (O_70,N_49641,N_49627);
nand UO_71 (O_71,N_49769,N_49289);
nand UO_72 (O_72,N_49851,N_49476);
nand UO_73 (O_73,N_49815,N_48882);
or UO_74 (O_74,N_48829,N_48895);
xor UO_75 (O_75,N_48424,N_48783);
xor UO_76 (O_76,N_48011,N_49904);
nor UO_77 (O_77,N_48230,N_49793);
xor UO_78 (O_78,N_49024,N_48789);
nand UO_79 (O_79,N_48621,N_48128);
nand UO_80 (O_80,N_49721,N_48961);
and UO_81 (O_81,N_49465,N_49439);
xnor UO_82 (O_82,N_48754,N_48505);
and UO_83 (O_83,N_48792,N_49688);
xnor UO_84 (O_84,N_48864,N_48355);
xnor UO_85 (O_85,N_48919,N_48325);
or UO_86 (O_86,N_49058,N_48824);
xor UO_87 (O_87,N_48512,N_48605);
nor UO_88 (O_88,N_49604,N_49072);
nand UO_89 (O_89,N_49856,N_48431);
xnor UO_90 (O_90,N_49433,N_48393);
and UO_91 (O_91,N_49008,N_48171);
and UO_92 (O_92,N_48821,N_49189);
nor UO_93 (O_93,N_49896,N_49378);
nand UO_94 (O_94,N_49526,N_49507);
xnor UO_95 (O_95,N_48593,N_49985);
or UO_96 (O_96,N_49108,N_48173);
nand UO_97 (O_97,N_49572,N_48475);
or UO_98 (O_98,N_48655,N_49797);
and UO_99 (O_99,N_48202,N_49949);
and UO_100 (O_100,N_48102,N_48763);
nor UO_101 (O_101,N_48734,N_48027);
nor UO_102 (O_102,N_48150,N_48620);
nand UO_103 (O_103,N_48228,N_48345);
xnor UO_104 (O_104,N_48408,N_48247);
and UO_105 (O_105,N_49261,N_48962);
or UO_106 (O_106,N_48954,N_48776);
nor UO_107 (O_107,N_49412,N_49063);
and UO_108 (O_108,N_48755,N_49068);
nand UO_109 (O_109,N_48887,N_48489);
and UO_110 (O_110,N_48811,N_49794);
nor UO_111 (O_111,N_48284,N_49753);
or UO_112 (O_112,N_49925,N_49716);
and UO_113 (O_113,N_48306,N_48623);
xnor UO_114 (O_114,N_48957,N_48617);
and UO_115 (O_115,N_49807,N_49528);
nand UO_116 (O_116,N_48320,N_48067);
nor UO_117 (O_117,N_48270,N_48736);
nand UO_118 (O_118,N_49402,N_48438);
xnor UO_119 (O_119,N_49473,N_48628);
nand UO_120 (O_120,N_48361,N_48137);
nor UO_121 (O_121,N_49011,N_49032);
xnor UO_122 (O_122,N_48869,N_48216);
or UO_123 (O_123,N_48423,N_49695);
nor UO_124 (O_124,N_48791,N_49987);
or UO_125 (O_125,N_48400,N_49544);
and UO_126 (O_126,N_49491,N_49130);
xnor UO_127 (O_127,N_48407,N_49106);
nand UO_128 (O_128,N_48766,N_49855);
and UO_129 (O_129,N_49760,N_49004);
xnor UO_130 (O_130,N_48127,N_48552);
xnor UO_131 (O_131,N_48019,N_49578);
xor UO_132 (O_132,N_49150,N_49867);
and UO_133 (O_133,N_49204,N_48040);
or UO_134 (O_134,N_49222,N_48348);
nand UO_135 (O_135,N_49386,N_48850);
and UO_136 (O_136,N_49496,N_48086);
nand UO_137 (O_137,N_48382,N_49983);
or UO_138 (O_138,N_49423,N_48099);
nand UO_139 (O_139,N_48835,N_48362);
and UO_140 (O_140,N_49935,N_48104);
nand UO_141 (O_141,N_49472,N_49061);
nand UO_142 (O_142,N_48070,N_49873);
xnor UO_143 (O_143,N_49969,N_49639);
nor UO_144 (O_144,N_49347,N_48669);
xor UO_145 (O_145,N_49515,N_48075);
or UO_146 (O_146,N_48364,N_48910);
nor UO_147 (O_147,N_48684,N_49543);
xor UO_148 (O_148,N_48115,N_48807);
xor UO_149 (O_149,N_48458,N_48426);
or UO_150 (O_150,N_48588,N_49495);
xor UO_151 (O_151,N_48170,N_49406);
and UO_152 (O_152,N_48637,N_48278);
nor UO_153 (O_153,N_49519,N_48773);
nand UO_154 (O_154,N_49101,N_48994);
xnor UO_155 (O_155,N_48721,N_49588);
nand UO_156 (O_156,N_49692,N_49861);
nand UO_157 (O_157,N_49321,N_49538);
xor UO_158 (O_158,N_49616,N_48031);
xnor UO_159 (O_159,N_49979,N_48956);
nor UO_160 (O_160,N_49265,N_48907);
and UO_161 (O_161,N_48132,N_49612);
nor UO_162 (O_162,N_48580,N_49383);
nor UO_163 (O_163,N_49550,N_48276);
or UO_164 (O_164,N_49144,N_48052);
nand UO_165 (O_165,N_49147,N_49451);
nor UO_166 (O_166,N_49757,N_49482);
and UO_167 (O_167,N_48218,N_49954);
nand UO_168 (O_168,N_48330,N_48264);
xor UO_169 (O_169,N_48913,N_49539);
nor UO_170 (O_170,N_49821,N_48622);
nand UO_171 (O_171,N_48050,N_48583);
nand UO_172 (O_172,N_48336,N_49279);
or UO_173 (O_173,N_48940,N_49152);
nand UO_174 (O_174,N_48538,N_49919);
or UO_175 (O_175,N_49116,N_49494);
nand UO_176 (O_176,N_49389,N_49000);
or UO_177 (O_177,N_48160,N_48058);
nor UO_178 (O_178,N_49015,N_49039);
xnor UO_179 (O_179,N_48813,N_48323);
and UO_180 (O_180,N_49732,N_49914);
nor UO_181 (O_181,N_49668,N_48561);
and UO_182 (O_182,N_48235,N_49866);
or UO_183 (O_183,N_48417,N_49697);
or UO_184 (O_184,N_48949,N_49045);
xnor UO_185 (O_185,N_49959,N_48905);
and UO_186 (O_186,N_49809,N_48647);
and UO_187 (O_187,N_48248,N_49891);
nand UO_188 (O_188,N_48074,N_49994);
nand UO_189 (O_189,N_48800,N_49838);
and UO_190 (O_190,N_49666,N_48888);
and UO_191 (O_191,N_48809,N_49163);
and UO_192 (O_192,N_48756,N_48060);
nand UO_193 (O_193,N_49468,N_49067);
or UO_194 (O_194,N_49435,N_48377);
nand UO_195 (O_195,N_48402,N_49234);
and UO_196 (O_196,N_48713,N_49117);
nor UO_197 (O_197,N_48644,N_48654);
or UO_198 (O_198,N_49844,N_48814);
and UO_199 (O_199,N_48045,N_49316);
nand UO_200 (O_200,N_48319,N_48502);
and UO_201 (O_201,N_48532,N_49715);
nor UO_202 (O_202,N_49514,N_49537);
nand UO_203 (O_203,N_49429,N_49643);
and UO_204 (O_204,N_48563,N_49018);
or UO_205 (O_205,N_49022,N_48056);
or UO_206 (O_206,N_48448,N_49879);
and UO_207 (O_207,N_48275,N_49013);
and UO_208 (O_208,N_49180,N_48161);
or UO_209 (O_209,N_48979,N_49466);
xnor UO_210 (O_210,N_49215,N_49874);
and UO_211 (O_211,N_48988,N_49893);
xor UO_212 (O_212,N_48480,N_49346);
nand UO_213 (O_213,N_48942,N_48078);
xnor UO_214 (O_214,N_48051,N_49531);
or UO_215 (O_215,N_49372,N_49023);
nor UO_216 (O_216,N_49567,N_49853);
nor UO_217 (O_217,N_48030,N_49859);
and UO_218 (O_218,N_49611,N_48172);
xnor UO_219 (O_219,N_49541,N_49452);
xor UO_220 (O_220,N_48120,N_49823);
nand UO_221 (O_221,N_49256,N_49774);
nand UO_222 (O_222,N_49816,N_49796);
and UO_223 (O_223,N_49506,N_49808);
and UO_224 (O_224,N_49027,N_49285);
and UO_225 (O_225,N_49705,N_48168);
nand UO_226 (O_226,N_48514,N_48582);
nand UO_227 (O_227,N_48085,N_48221);
nor UO_228 (O_228,N_48372,N_49380);
or UO_229 (O_229,N_48640,N_49766);
nand UO_230 (O_230,N_49247,N_48993);
or UO_231 (O_231,N_48317,N_48590);
and UO_232 (O_232,N_48193,N_49684);
xnor UO_233 (O_233,N_49126,N_49966);
and UO_234 (O_234,N_49928,N_48639);
or UO_235 (O_235,N_49263,N_48233);
or UO_236 (O_236,N_49290,N_48494);
xor UO_237 (O_237,N_49573,N_49618);
nand UO_238 (O_238,N_48281,N_48642);
nand UO_239 (O_239,N_49418,N_48017);
and UO_240 (O_240,N_49581,N_48737);
nor UO_241 (O_241,N_48781,N_48964);
xnor UO_242 (O_242,N_48860,N_49663);
xor UO_243 (O_243,N_48148,N_49040);
nor UO_244 (O_244,N_48316,N_48528);
xnor UO_245 (O_245,N_48619,N_49902);
nand UO_246 (O_246,N_48698,N_48986);
or UO_247 (O_247,N_49890,N_48541);
or UO_248 (O_248,N_48923,N_48381);
xnor UO_249 (O_249,N_48491,N_49308);
and UO_250 (O_250,N_48189,N_49786);
nand UO_251 (O_251,N_48404,N_49119);
nand UO_252 (O_252,N_48421,N_48805);
nor UO_253 (O_253,N_48263,N_49081);
nor UO_254 (O_254,N_48474,N_48718);
or UO_255 (O_255,N_49259,N_48097);
xor UO_256 (O_256,N_49761,N_48894);
or UO_257 (O_257,N_49177,N_48454);
nor UO_258 (O_258,N_48455,N_48871);
xor UO_259 (O_259,N_48662,N_48996);
nand UO_260 (O_260,N_48818,N_49508);
nand UO_261 (O_261,N_49273,N_49249);
and UO_262 (O_262,N_49052,N_49440);
nand UO_263 (O_263,N_48510,N_48927);
xor UO_264 (O_264,N_48761,N_49437);
or UO_265 (O_265,N_48094,N_48481);
xnor UO_266 (O_266,N_48587,N_48003);
nand UO_267 (O_267,N_48113,N_48542);
or UO_268 (O_268,N_49336,N_49521);
nand UO_269 (O_269,N_48520,N_49790);
nand UO_270 (O_270,N_49074,N_48719);
and UO_271 (O_271,N_49583,N_49140);
nor UO_272 (O_272,N_48395,N_49518);
nor UO_273 (O_273,N_49590,N_49062);
and UO_274 (O_274,N_48439,N_49300);
and UO_275 (O_275,N_48100,N_49197);
nor UO_276 (O_276,N_49777,N_48570);
or UO_277 (O_277,N_48391,N_48997);
or UO_278 (O_278,N_48777,N_49202);
xor UO_279 (O_279,N_48169,N_48139);
or UO_280 (O_280,N_48708,N_48206);
and UO_281 (O_281,N_48311,N_49620);
and UO_282 (O_282,N_48236,N_48522);
and UO_283 (O_283,N_49320,N_49199);
or UO_284 (O_284,N_48544,N_48631);
nand UO_285 (O_285,N_48154,N_49513);
nand UO_286 (O_286,N_48354,N_49175);
and UO_287 (O_287,N_49765,N_49626);
or UO_288 (O_288,N_48668,N_48799);
xor UO_289 (O_289,N_48209,N_49960);
nand UO_290 (O_290,N_48591,N_48376);
xor UO_291 (O_291,N_49558,N_49835);
nand UO_292 (O_292,N_48511,N_49781);
nand UO_293 (O_293,N_49819,N_48344);
and UO_294 (O_294,N_49575,N_48877);
nand UO_295 (O_295,N_49394,N_48255);
and UO_296 (O_296,N_48497,N_48597);
nor UO_297 (O_297,N_48269,N_48863);
and UO_298 (O_298,N_48486,N_48677);
or UO_299 (O_299,N_49178,N_49333);
or UO_300 (O_300,N_48346,N_48479);
nor UO_301 (O_301,N_49814,N_48865);
or UO_302 (O_302,N_48191,N_49037);
nand UO_303 (O_303,N_48749,N_48730);
and UO_304 (O_304,N_48147,N_48398);
and UO_305 (O_305,N_49090,N_48608);
and UO_306 (O_306,N_48337,N_48280);
and UO_307 (O_307,N_49179,N_48711);
nor UO_308 (O_308,N_49773,N_49978);
nor UO_309 (O_309,N_48769,N_49111);
or UO_310 (O_310,N_48679,N_49990);
or UO_311 (O_311,N_48326,N_49683);
nor UO_312 (O_312,N_48268,N_48924);
nand UO_313 (O_313,N_49257,N_48690);
or UO_314 (O_314,N_49190,N_49141);
or UO_315 (O_315,N_48731,N_48293);
and UO_316 (O_316,N_48930,N_48902);
or UO_317 (O_317,N_48116,N_49951);
and UO_318 (O_318,N_48692,N_49266);
nand UO_319 (O_319,N_49446,N_49789);
and UO_320 (O_320,N_48140,N_49899);
nand UO_321 (O_321,N_48485,N_48257);
or UO_322 (O_322,N_49365,N_48014);
nor UO_323 (O_323,N_48613,N_49129);
nand UO_324 (O_324,N_49432,N_49229);
xnor UO_325 (O_325,N_48166,N_49373);
or UO_326 (O_326,N_48005,N_49758);
or UO_327 (O_327,N_49736,N_49702);
or UO_328 (O_328,N_49780,N_49510);
xor UO_329 (O_329,N_48163,N_49288);
xor UO_330 (O_330,N_49121,N_49863);
nand UO_331 (O_331,N_49699,N_48854);
nor UO_332 (O_332,N_49381,N_49995);
and UO_333 (O_333,N_48695,N_49326);
nand UO_334 (O_334,N_49332,N_48999);
nor UO_335 (O_335,N_48224,N_49788);
nor UO_336 (O_336,N_48771,N_48419);
or UO_337 (O_337,N_49589,N_48142);
or UO_338 (O_338,N_49828,N_48611);
nor UO_339 (O_339,N_48678,N_48420);
or UO_340 (O_340,N_49157,N_49426);
nor UO_341 (O_341,N_48700,N_48703);
nor UO_342 (O_342,N_48564,N_48328);
and UO_343 (O_343,N_48090,N_49030);
nor UO_344 (O_344,N_49967,N_48530);
or UO_345 (O_345,N_48616,N_49049);
nor UO_346 (O_346,N_49145,N_49877);
xor UO_347 (O_347,N_48691,N_48025);
and UO_348 (O_348,N_49210,N_49595);
nor UO_349 (O_349,N_48515,N_48855);
and UO_350 (O_350,N_49950,N_48405);
xnor UO_351 (O_351,N_48950,N_49139);
or UO_352 (O_352,N_48518,N_49657);
nand UO_353 (O_353,N_48650,N_49020);
nand UO_354 (O_354,N_49637,N_49443);
nor UO_355 (O_355,N_48250,N_49176);
nand UO_356 (O_356,N_48251,N_49294);
nand UO_357 (O_357,N_49354,N_49645);
or UO_358 (O_358,N_49881,N_49517);
and UO_359 (O_359,N_48111,N_48077);
xnor UO_360 (O_360,N_49161,N_49858);
nand UO_361 (O_361,N_48982,N_48671);
or UO_362 (O_362,N_48312,N_49393);
or UO_363 (O_363,N_49667,N_49630);
nand UO_364 (O_364,N_48686,N_48852);
and UO_365 (O_365,N_49596,N_49219);
nor UO_366 (O_366,N_49310,N_48868);
nor UO_367 (O_367,N_48299,N_48308);
xor UO_368 (O_368,N_48277,N_48282);
nor UO_369 (O_369,N_49785,N_49591);
or UO_370 (O_370,N_48618,N_49122);
nor UO_371 (O_371,N_49170,N_49876);
xor UO_372 (O_372,N_48291,N_48036);
nand UO_373 (O_373,N_48213,N_49377);
and UO_374 (O_374,N_48609,N_49169);
nor UO_375 (O_375,N_48985,N_48215);
and UO_376 (O_376,N_48467,N_49056);
nand UO_377 (O_377,N_49010,N_49298);
xnor UO_378 (O_378,N_49271,N_48288);
nor UO_379 (O_379,N_49862,N_49128);
nor UO_380 (O_380,N_48449,N_49231);
nand UO_381 (O_381,N_49097,N_48219);
and UO_382 (O_382,N_48343,N_49917);
and UO_383 (O_383,N_48658,N_49258);
nor UO_384 (O_384,N_48008,N_49014);
nand UO_385 (O_385,N_49831,N_48849);
or UO_386 (O_386,N_49564,N_49687);
nand UO_387 (O_387,N_48307,N_49171);
xor UO_388 (O_388,N_48672,N_49167);
nand UO_389 (O_389,N_48796,N_49220);
nor UO_390 (O_390,N_49434,N_49376);
and UO_391 (O_391,N_48959,N_49500);
and UO_392 (O_392,N_48470,N_48939);
nor UO_393 (O_393,N_48130,N_48101);
or UO_394 (O_394,N_49295,N_48028);
nand UO_395 (O_395,N_49860,N_48782);
and UO_396 (O_396,N_48596,N_48886);
nand UO_397 (O_397,N_48106,N_49091);
and UO_398 (O_398,N_49520,N_48152);
nor UO_399 (O_399,N_48918,N_48851);
nand UO_400 (O_400,N_48088,N_48462);
and UO_401 (O_401,N_49363,N_49213);
xor UO_402 (O_402,N_49908,N_49038);
nor UO_403 (O_403,N_48182,N_49704);
or UO_404 (O_404,N_49092,N_48764);
xnor UO_405 (O_405,N_48197,N_49784);
xor UO_406 (O_406,N_48790,N_49487);
xor UO_407 (O_407,N_49502,N_49934);
and UO_408 (O_408,N_49043,N_49416);
nand UO_409 (O_409,N_48237,N_49751);
and UO_410 (O_410,N_49525,N_49962);
nor UO_411 (O_411,N_49854,N_48984);
nand UO_412 (O_412,N_49557,N_48975);
nor UO_413 (O_413,N_49455,N_48178);
nand UO_414 (O_414,N_49885,N_49421);
nand UO_415 (O_415,N_49799,N_48225);
or UO_416 (O_416,N_48048,N_48492);
and UO_417 (O_417,N_49009,N_48774);
and UO_418 (O_418,N_49690,N_48847);
nand UO_419 (O_419,N_48205,N_48856);
nor UO_420 (O_420,N_48187,N_49405);
and UO_421 (O_421,N_49723,N_49331);
or UO_422 (O_422,N_48578,N_49811);
and UO_423 (O_423,N_49105,N_48663);
xor UO_424 (O_424,N_49553,N_49267);
nor UO_425 (O_425,N_49770,N_49469);
and UO_426 (O_426,N_49529,N_48870);
nand UO_427 (O_427,N_49230,N_49592);
and UO_428 (O_428,N_49255,N_49127);
or UO_429 (O_429,N_48819,N_48445);
or UO_430 (O_430,N_49442,N_48380);
xnor UO_431 (O_431,N_49103,N_49973);
nand UO_432 (O_432,N_48352,N_49738);
xor UO_433 (O_433,N_48249,N_49387);
and UO_434 (O_434,N_48947,N_49481);
nor UO_435 (O_435,N_48753,N_48203);
nor UO_436 (O_436,N_48815,N_48124);
or UO_437 (O_437,N_49042,N_48453);
nand UO_438 (O_438,N_48371,N_48735);
xor UO_439 (O_439,N_48061,N_48638);
nor UO_440 (O_440,N_49560,N_49070);
nand UO_441 (O_441,N_49549,N_48676);
and UO_442 (O_442,N_48759,N_48020);
nor UO_443 (O_443,N_48707,N_49635);
or UO_444 (O_444,N_48357,N_48080);
and UO_445 (O_445,N_49677,N_48645);
or UO_446 (O_446,N_49303,N_49742);
nor UO_447 (O_447,N_49209,N_48509);
nand UO_448 (O_448,N_49124,N_49135);
xor UO_449 (O_449,N_49390,N_49275);
nor UO_450 (O_450,N_49109,N_48351);
or UO_451 (O_451,N_49680,N_48848);
nor UO_452 (O_452,N_49901,N_49223);
and UO_453 (O_453,N_48643,N_49806);
or UO_454 (O_454,N_48861,N_48876);
or UO_455 (O_455,N_48274,N_48441);
nand UO_456 (O_456,N_48112,N_49729);
nand UO_457 (O_457,N_49395,N_48283);
nand UO_458 (O_458,N_49345,N_49207);
and UO_459 (O_459,N_49798,N_49041);
and UO_460 (O_460,N_49459,N_49277);
nor UO_461 (O_461,N_49849,N_49497);
xor UO_462 (O_462,N_48180,N_49311);
nor UO_463 (O_463,N_49110,N_48023);
nand UO_464 (O_464,N_49102,N_48612);
and UO_465 (O_465,N_48729,N_49449);
nand UO_466 (O_466,N_49570,N_49536);
and UO_467 (O_467,N_49887,N_48944);
xnor UO_468 (O_468,N_48149,N_49601);
nand UO_469 (O_469,N_49046,N_49755);
and UO_470 (O_470,N_48546,N_48242);
or UO_471 (O_471,N_48903,N_48788);
or UO_472 (O_472,N_48301,N_49089);
nor UO_473 (O_473,N_49464,N_49036);
nor UO_474 (O_474,N_49927,N_49114);
nand UO_475 (O_475,N_48747,N_48429);
or UO_476 (O_476,N_49328,N_48210);
or UO_477 (O_477,N_49533,N_48627);
or UO_478 (O_478,N_49980,N_48141);
or UO_479 (O_479,N_49989,N_48911);
or UO_480 (O_480,N_49756,N_49852);
xnor UO_481 (O_481,N_49512,N_48929);
xnor UO_482 (O_482,N_48524,N_49244);
and UO_483 (O_483,N_48842,N_49670);
or UO_484 (O_484,N_49339,N_48192);
xor UO_485 (O_485,N_49605,N_48367);
nor UO_486 (O_486,N_48839,N_48804);
nand UO_487 (O_487,N_48874,N_48295);
and UO_488 (O_488,N_48872,N_48673);
and UO_489 (O_489,N_48867,N_49571);
nand UO_490 (O_490,N_48937,N_48488);
and UO_491 (O_491,N_49278,N_49477);
nor UO_492 (O_492,N_49782,N_49349);
or UO_493 (O_493,N_49868,N_49628);
or UO_494 (O_494,N_49206,N_49865);
nor UO_495 (O_495,N_49694,N_49357);
and UO_496 (O_496,N_48935,N_48879);
or UO_497 (O_497,N_48568,N_49080);
or UO_498 (O_498,N_49286,N_48266);
and UO_499 (O_499,N_48185,N_49136);
nor UO_500 (O_500,N_48156,N_48566);
and UO_501 (O_501,N_49897,N_49073);
or UO_502 (O_502,N_48581,N_49651);
nor UO_503 (O_503,N_49915,N_49554);
xor UO_504 (O_504,N_49375,N_49463);
and UO_505 (O_505,N_48450,N_49972);
nand UO_506 (O_506,N_49568,N_48253);
nor UO_507 (O_507,N_48878,N_49945);
and UO_508 (O_508,N_49939,N_48359);
nand UO_509 (O_509,N_48009,N_49740);
nor UO_510 (O_510,N_49314,N_48884);
and UO_511 (O_511,N_48010,N_49752);
xor UO_512 (O_512,N_48055,N_48661);
nand UO_513 (O_513,N_48109,N_48531);
or UO_514 (O_514,N_49087,N_49869);
nor UO_515 (O_515,N_49975,N_49686);
and UO_516 (O_516,N_48503,N_48914);
and UO_517 (O_517,N_49615,N_49159);
and UO_518 (O_518,N_49597,N_48599);
or UO_519 (O_519,N_49580,N_49226);
and UO_520 (O_520,N_48535,N_48478);
nor UO_521 (O_521,N_48368,N_48793);
nand UO_522 (O_522,N_49243,N_48899);
nor UO_523 (O_523,N_49624,N_49238);
or UO_524 (O_524,N_48748,N_49242);
and UO_525 (O_525,N_48705,N_48548);
and UO_526 (O_526,N_49470,N_49415);
xnor UO_527 (O_527,N_49276,N_48960);
and UO_528 (O_528,N_49511,N_49552);
xnor UO_529 (O_529,N_49696,N_49188);
nor UO_530 (O_530,N_49174,N_49485);
xor UO_531 (O_531,N_49974,N_48259);
nor UO_532 (O_532,N_49425,N_49625);
and UO_533 (O_533,N_49239,N_49727);
nor UO_534 (O_534,N_49312,N_49191);
nor UO_535 (O_535,N_48286,N_49417);
and UO_536 (O_536,N_49196,N_49392);
xnor UO_537 (O_537,N_48875,N_49710);
nor UO_538 (O_538,N_48844,N_48057);
xnor UO_539 (O_539,N_48134,N_48318);
or UO_540 (O_540,N_48410,N_48649);
nand UO_541 (O_541,N_49493,N_48968);
nor UO_542 (O_542,N_49916,N_48092);
nand UO_543 (O_543,N_48657,N_48490);
nand UO_544 (O_544,N_49924,N_49240);
and UO_545 (O_545,N_49028,N_49475);
and UO_546 (O_546,N_49031,N_49282);
and UO_547 (O_547,N_48349,N_49154);
and UO_548 (O_548,N_48504,N_49050);
and UO_549 (O_549,N_49227,N_48446);
and UO_550 (O_550,N_49864,N_49361);
xor UO_551 (O_551,N_48334,N_49920);
or UO_552 (O_552,N_49524,N_49120);
and UO_553 (O_553,N_48208,N_48465);
nand UO_554 (O_554,N_48477,N_48652);
xnor UO_555 (O_555,N_48243,N_48435);
or UO_556 (O_556,N_48026,N_48443);
nand UO_557 (O_557,N_49938,N_49608);
or UO_558 (O_558,N_48241,N_49713);
xnor UO_559 (O_559,N_48958,N_48825);
and UO_560 (O_560,N_48659,N_48029);
and UO_561 (O_561,N_49430,N_49981);
nand UO_562 (O_562,N_48724,N_48388);
or UO_563 (O_563,N_48709,N_49958);
nand UO_564 (O_564,N_49205,N_48332);
nor UO_565 (O_565,N_49996,N_49556);
nor UO_566 (O_566,N_49836,N_49055);
and UO_567 (O_567,N_49772,N_49991);
or UO_568 (O_568,N_48806,N_48767);
xnor UO_569 (O_569,N_49579,N_49398);
and UO_570 (O_570,N_49225,N_48415);
nand UO_571 (O_571,N_49131,N_49252);
or UO_572 (O_572,N_49293,N_49530);
nor UO_573 (O_573,N_48292,N_48482);
xor UO_574 (O_574,N_48751,N_48574);
nand UO_575 (O_575,N_49658,N_48537);
nor UO_576 (O_576,N_49334,N_49351);
nor UO_577 (O_577,N_48770,N_49676);
nand UO_578 (O_578,N_48459,N_48741);
nand UO_579 (O_579,N_49355,N_48602);
or UO_580 (O_580,N_48720,N_48188);
nand UO_581 (O_581,N_48493,N_49012);
and UO_582 (O_582,N_48897,N_48063);
and UO_583 (O_583,N_48557,N_49587);
or UO_584 (O_584,N_49060,N_48012);
and UO_585 (O_585,N_49805,N_49832);
or UO_586 (O_586,N_48091,N_48595);
and UO_587 (O_587,N_49675,N_48227);
nor UO_588 (O_588,N_49795,N_49044);
or UO_589 (O_589,N_48199,N_48945);
xor UO_590 (O_590,N_48428,N_49309);
and UO_591 (O_591,N_49457,N_48190);
nor UO_592 (O_592,N_48181,N_49649);
nand UO_593 (O_593,N_49364,N_49467);
nor UO_594 (O_594,N_49385,N_49638);
nand UO_595 (O_595,N_49593,N_49728);
and UO_596 (O_596,N_48107,N_49703);
and UO_597 (O_597,N_48555,N_49846);
and UO_598 (O_598,N_48928,N_49906);
xnor UO_599 (O_599,N_48340,N_49143);
nor UO_600 (O_600,N_48853,N_49146);
xor UO_601 (O_601,N_48339,N_49976);
xnor UO_602 (O_602,N_49817,N_49843);
xnor UO_603 (O_603,N_49764,N_49970);
nor UO_604 (O_604,N_49066,N_48466);
xnor UO_605 (O_605,N_48506,N_48068);
or UO_606 (O_606,N_48904,N_48810);
xnor UO_607 (O_607,N_49913,N_48779);
nand UO_608 (O_608,N_49633,N_48196);
or UO_609 (O_609,N_49957,N_49427);
or UO_610 (O_610,N_48526,N_48000);
xor UO_611 (O_611,N_48217,N_48717);
nand UO_612 (O_612,N_48129,N_49984);
and UO_613 (O_613,N_49669,N_49614);
or UO_614 (O_614,N_48464,N_48296);
xnor UO_615 (O_615,N_48159,N_48823);
and UO_616 (O_616,N_48694,N_48119);
nor UO_617 (O_617,N_48401,N_49971);
nand UO_618 (O_618,N_48701,N_49963);
or UO_619 (O_619,N_48081,N_48803);
or UO_620 (O_620,N_48083,N_48353);
xnor UO_621 (O_621,N_49413,N_49775);
nand UO_622 (O_622,N_48324,N_49490);
nand UO_623 (O_623,N_48594,N_48164);
nor UO_624 (O_624,N_48843,N_49480);
xnor UO_625 (O_625,N_48932,N_48035);
or UO_626 (O_626,N_49399,N_49253);
nor UO_627 (O_627,N_48840,N_48989);
nand UO_628 (O_628,N_48122,N_48966);
or UO_629 (O_629,N_49791,N_49322);
nand UO_630 (O_630,N_49431,N_49414);
nor UO_631 (O_631,N_48501,N_49149);
xor UO_632 (O_632,N_48606,N_48540);
xnor UO_633 (O_633,N_49342,N_49166);
nand UO_634 (O_634,N_49193,N_49892);
or UO_635 (O_635,N_48271,N_49329);
nor UO_636 (O_636,N_49005,N_49759);
nor UO_637 (O_637,N_49982,N_49138);
or UO_638 (O_638,N_49725,N_48496);
xor UO_639 (O_639,N_48648,N_48262);
xor UO_640 (O_640,N_48403,N_49148);
or UO_641 (O_641,N_48093,N_49268);
xnor UO_642 (O_642,N_49115,N_49660);
nand UO_643 (O_643,N_48411,N_49623);
or UO_644 (O_644,N_49501,N_49195);
xor UO_645 (O_645,N_48434,N_48577);
or UO_646 (O_646,N_48032,N_49164);
or UO_647 (O_647,N_48157,N_48575);
nor UO_648 (O_648,N_48135,N_49898);
or UO_649 (O_649,N_48567,N_48980);
xor UO_650 (O_650,N_48413,N_48948);
nor UO_651 (O_651,N_48858,N_49813);
xor UO_652 (O_652,N_49450,N_48385);
and UO_653 (O_653,N_49947,N_49396);
nand UO_654 (O_654,N_48399,N_48558);
xor UO_655 (O_655,N_49021,N_49634);
or UO_656 (O_656,N_49754,N_48079);
xor UO_657 (O_657,N_49582,N_48909);
or UO_658 (O_658,N_49337,N_48396);
xnor UO_659 (O_659,N_48795,N_48397);
or UO_660 (O_660,N_48333,N_48238);
xnor UO_661 (O_661,N_49574,N_48366);
xnor UO_662 (O_662,N_48740,N_48831);
xnor UO_663 (O_663,N_48576,N_48013);
nand UO_664 (O_664,N_49033,N_48778);
nor UO_665 (O_665,N_49653,N_48315);
nor UO_666 (O_666,N_49104,N_49118);
and UO_667 (O_667,N_49492,N_49158);
and UO_668 (O_668,N_48044,N_49878);
or UO_669 (O_669,N_48955,N_49162);
xor UO_670 (O_670,N_49632,N_48002);
xnor UO_671 (O_671,N_48926,N_48452);
or UO_672 (O_672,N_49585,N_48816);
xnor UO_673 (O_673,N_48565,N_48906);
and UO_674 (O_674,N_48513,N_49997);
and UO_675 (O_675,N_49462,N_48901);
nor UO_676 (O_676,N_49112,N_48922);
xnor UO_677 (O_677,N_49400,N_49584);
or UO_678 (O_678,N_49254,N_48933);
and UO_679 (O_679,N_49882,N_48881);
nand UO_680 (O_680,N_49540,N_48744);
or UO_681 (O_681,N_48880,N_49260);
and UO_682 (O_682,N_48681,N_48634);
nor UO_683 (O_683,N_48812,N_48977);
xor UO_684 (O_684,N_49160,N_49085);
nand UO_685 (O_685,N_49301,N_49561);
or UO_686 (O_686,N_48006,N_49304);
nand UO_687 (O_687,N_49340,N_49609);
nor UO_688 (O_688,N_48891,N_48136);
xor UO_689 (O_689,N_48290,N_49292);
and UO_690 (O_690,N_49461,N_48232);
or UO_691 (O_691,N_49323,N_48670);
and UO_692 (O_692,N_49344,N_48912);
or UO_693 (O_693,N_49679,N_49746);
nor UO_694 (O_694,N_48049,N_49262);
and UO_695 (O_695,N_48817,N_49932);
and UO_696 (O_696,N_49857,N_49374);
or UO_697 (O_697,N_49930,N_49248);
xor UO_698 (O_698,N_48885,N_49217);
and UO_699 (O_699,N_48444,N_48667);
nor UO_700 (O_700,N_48666,N_49698);
xor UO_701 (O_701,N_48298,N_49889);
nand UO_702 (O_702,N_48064,N_48289);
xnor UO_703 (O_703,N_49306,N_49025);
xnor UO_704 (O_704,N_48043,N_48545);
and UO_705 (O_705,N_48801,N_48110);
and UO_706 (O_706,N_48500,N_48460);
nand UO_707 (O_707,N_48126,N_49317);
or UO_708 (O_708,N_49356,N_48373);
xnor UO_709 (O_709,N_48551,N_49007);
xnor UO_710 (O_710,N_48437,N_49840);
xnor UO_711 (O_711,N_49762,N_48042);
xnor UO_712 (O_712,N_48607,N_48723);
or UO_713 (O_713,N_49888,N_49409);
and UO_714 (O_714,N_49367,N_49717);
nor UO_715 (O_715,N_48374,N_48516);
or UO_716 (O_716,N_49955,N_48832);
xnor UO_717 (O_717,N_48394,N_48990);
nand UO_718 (O_718,N_49722,N_48584);
or UO_719 (O_719,N_49918,N_48772);
or UO_720 (O_720,N_49636,N_48733);
xor UO_721 (O_721,N_48715,N_48787);
or UO_722 (O_722,N_49909,N_48369);
nor UO_723 (O_723,N_49894,N_49078);
or UO_724 (O_724,N_49338,N_49458);
nand UO_725 (O_725,N_48234,N_49133);
nand UO_726 (O_726,N_48550,N_48201);
nand UO_727 (O_727,N_48245,N_48963);
nand UO_728 (O_728,N_49305,N_49335);
nor UO_729 (O_729,N_48693,N_49187);
nand UO_730 (O_730,N_48279,N_48738);
nand UO_731 (O_731,N_48917,N_49516);
xnor UO_732 (O_732,N_49505,N_48614);
or UO_733 (O_733,N_49082,N_49407);
xnor UO_734 (O_734,N_48716,N_49921);
nor UO_735 (O_735,N_48571,N_49871);
nor UO_736 (O_736,N_49281,N_49576);
nand UO_737 (O_737,N_48664,N_49931);
and UO_738 (O_738,N_48680,N_48833);
nor UO_739 (O_739,N_48155,N_49848);
and UO_740 (O_740,N_48222,N_49820);
xnor UO_741 (O_741,N_49019,N_48144);
or UO_742 (O_742,N_49522,N_49839);
and UO_743 (O_743,N_48946,N_49348);
xnor UO_744 (O_744,N_48521,N_49532);
nand UO_745 (O_745,N_49741,N_49173);
xnor UO_746 (O_746,N_49600,N_49968);
nor UO_747 (O_747,N_48331,N_48335);
or UO_748 (O_748,N_49047,N_48527);
nor UO_749 (O_749,N_49940,N_49681);
and UO_750 (O_750,N_49603,N_48018);
nor UO_751 (O_751,N_49483,N_48952);
nor UO_752 (O_752,N_48347,N_49743);
and UO_753 (O_753,N_48732,N_49404);
nand UO_754 (O_754,N_49640,N_49546);
and UO_755 (O_755,N_49693,N_48073);
xnor UO_756 (O_756,N_49192,N_49912);
xnor UO_757 (O_757,N_48370,N_49993);
xor UO_758 (O_758,N_48712,N_48223);
nor UO_759 (O_759,N_48378,N_48007);
xor UO_760 (O_760,N_49961,N_48176);
or UO_761 (O_761,N_49084,N_48688);
or UO_762 (O_762,N_49656,N_49324);
and UO_763 (O_763,N_49438,N_48414);
and UO_764 (O_764,N_49100,N_49952);
nand UO_765 (O_765,N_48038,N_48921);
and UO_766 (O_766,N_48992,N_48601);
nor UO_767 (O_767,N_49422,N_48087);
nand UO_768 (O_768,N_48974,N_48529);
xor UO_769 (O_769,N_49379,N_49718);
or UO_770 (O_770,N_48727,N_49563);
and UO_771 (O_771,N_49269,N_49720);
or UO_772 (O_772,N_49534,N_49977);
nand UO_773 (O_773,N_48714,N_49569);
xor UO_774 (O_774,N_48383,N_48589);
and UO_775 (O_775,N_49327,N_49391);
nor UO_776 (O_776,N_48743,N_49224);
and UO_777 (O_777,N_49186,N_48473);
nand UO_778 (O_778,N_48165,N_49936);
xnor UO_779 (O_779,N_49088,N_48784);
nor UO_780 (O_780,N_49707,N_49673);
or UO_781 (O_781,N_49296,N_48592);
xnor UO_782 (O_782,N_49478,N_48543);
xor UO_783 (O_783,N_48547,N_48041);
or UO_784 (O_784,N_48651,N_49845);
nand UO_785 (O_785,N_49922,N_49079);
nor UO_786 (O_786,N_48387,N_48069);
and UO_787 (O_787,N_49448,N_49401);
xnor UO_788 (O_788,N_49594,N_49251);
and UO_789 (O_789,N_48153,N_49076);
nand UO_790 (O_790,N_49992,N_49847);
xor UO_791 (O_791,N_49218,N_49923);
xnor UO_792 (O_792,N_48697,N_49674);
nor UO_793 (O_793,N_49235,N_49098);
or UO_794 (O_794,N_49201,N_48146);
and UO_795 (O_795,N_48167,N_48517);
or UO_796 (O_796,N_49964,N_49094);
or UO_797 (O_797,N_48936,N_48071);
xor UO_798 (O_798,N_48386,N_48162);
and UO_799 (O_799,N_49999,N_48310);
or UO_800 (O_800,N_48972,N_49003);
and UO_801 (O_801,N_48342,N_49436);
xor UO_802 (O_802,N_49910,N_48495);
nand UO_803 (O_803,N_49731,N_48685);
nand UO_804 (O_804,N_48204,N_48258);
nor UO_805 (O_805,N_49509,N_49325);
xnor UO_806 (O_806,N_49075,N_48200);
xor UO_807 (O_807,N_48476,N_49610);
or UO_808 (O_808,N_48054,N_49942);
nor UO_809 (O_809,N_48533,N_49353);
and UO_810 (O_810,N_49343,N_48991);
nor UO_811 (O_811,N_49701,N_49662);
nor UO_812 (O_812,N_48033,N_48442);
nor UO_813 (O_813,N_49221,N_49801);
or UO_814 (O_814,N_48261,N_48941);
or UO_815 (O_815,N_48797,N_49488);
nor UO_816 (O_816,N_48212,N_48226);
nor UO_817 (O_817,N_49559,N_48987);
xor UO_818 (O_818,N_49272,N_48943);
or UO_819 (O_819,N_49659,N_48586);
xor UO_820 (O_820,N_49988,N_48683);
nand UO_821 (O_821,N_49944,N_49071);
and UO_822 (O_822,N_49903,N_48925);
and UO_823 (O_823,N_49125,N_48696);
or UO_824 (O_824,N_48560,N_49291);
and UO_825 (O_825,N_49719,N_49142);
nand UO_826 (O_826,N_49802,N_49886);
nand UO_827 (O_827,N_49948,N_49748);
nor UO_828 (O_828,N_49661,N_49712);
or UO_829 (O_829,N_49054,N_48746);
xnor UO_830 (O_830,N_48256,N_49527);
xnor UO_831 (O_831,N_49211,N_49607);
and UO_832 (O_832,N_48610,N_48463);
nor UO_833 (O_833,N_49123,N_49002);
and UO_834 (O_834,N_48846,N_49682);
xnor UO_835 (O_835,N_48314,N_49315);
nand UO_836 (O_836,N_49504,N_49956);
and UO_837 (O_837,N_49484,N_49737);
nand UO_838 (O_838,N_48630,N_49420);
and UO_839 (O_839,N_48254,N_48653);
nor UO_840 (O_840,N_48556,N_48211);
nor UO_841 (O_841,N_49771,N_48632);
or UO_842 (O_842,N_49181,N_48121);
nand UO_843 (O_843,N_48265,N_48931);
nor UO_844 (O_844,N_48704,N_48304);
and UO_845 (O_845,N_48037,N_48138);
xnor UO_846 (O_846,N_48392,N_48579);
xnor UO_847 (O_847,N_48440,N_49368);
or UO_848 (O_848,N_48186,N_48866);
nor UO_849 (O_849,N_48836,N_48604);
nand UO_850 (O_850,N_48953,N_48084);
xnor UO_851 (O_851,N_48313,N_49330);
xor UO_852 (O_852,N_48425,N_48739);
xnor UO_853 (O_853,N_48065,N_48553);
or UO_854 (O_854,N_49241,N_48427);
nor UO_855 (O_855,N_48406,N_48573);
or UO_856 (O_856,N_48287,N_48758);
nand UO_857 (O_857,N_48656,N_49410);
xor UO_858 (O_858,N_48469,N_48059);
or UO_859 (O_859,N_48859,N_49822);
or UO_860 (O_860,N_49547,N_49358);
and UO_861 (O_861,N_49051,N_48760);
xor UO_862 (O_862,N_48585,N_48828);
nor UO_863 (O_863,N_49911,N_49053);
and UO_864 (O_864,N_49827,N_49350);
nor UO_865 (O_865,N_48321,N_48072);
or UO_866 (O_866,N_49246,N_48322);
nor UO_867 (O_867,N_49841,N_48363);
nor UO_868 (O_868,N_49388,N_49872);
and UO_869 (O_869,N_49065,N_48451);
nor UO_870 (O_870,N_48379,N_48820);
nor UO_871 (O_871,N_48883,N_48808);
xor UO_872 (O_872,N_48845,N_48066);
nand UO_873 (O_873,N_49096,N_48327);
nor UO_874 (O_874,N_48039,N_49830);
and UO_875 (O_875,N_48834,N_48471);
xor UO_876 (O_876,N_48096,N_48175);
nand UO_877 (O_877,N_48105,N_49307);
xor UO_878 (O_878,N_49926,N_48624);
nand UO_879 (O_879,N_48447,N_48239);
nor UO_880 (O_880,N_48267,N_49203);
or UO_881 (O_881,N_49503,N_49151);
xnor UO_882 (O_882,N_49155,N_49185);
and UO_883 (O_883,N_49613,N_49318);
and UO_884 (O_884,N_49763,N_48198);
or UO_885 (O_885,N_48915,N_49523);
xnor UO_886 (O_886,N_48983,N_49776);
or UO_887 (O_887,N_48430,N_48572);
xnor UO_888 (O_888,N_48889,N_49479);
or UO_889 (O_889,N_48433,N_48687);
nor UO_890 (O_890,N_49734,N_49652);
or UO_891 (O_891,N_49489,N_48231);
xor UO_892 (O_892,N_49804,N_49629);
nor UO_893 (O_893,N_48133,N_49986);
xnor UO_894 (O_894,N_49768,N_49565);
nor UO_895 (O_895,N_49907,N_48768);
nand UO_896 (O_896,N_49208,N_48525);
nor UO_897 (O_897,N_49655,N_49214);
nand UO_898 (O_898,N_48022,N_49447);
xor UO_899 (O_899,N_48123,N_49216);
nand UO_900 (O_900,N_48461,N_48131);
and UO_901 (O_901,N_49184,N_49424);
and UO_902 (O_902,N_48973,N_49408);
and UO_903 (O_903,N_49134,N_48726);
and UO_904 (O_904,N_49733,N_48285);
nor UO_905 (O_905,N_48549,N_49602);
or UO_906 (O_906,N_48893,N_48390);
or UO_907 (O_907,N_48976,N_48765);
or UO_908 (O_908,N_49264,N_48830);
and UO_909 (O_909,N_49319,N_49714);
nand UO_910 (O_910,N_48742,N_49107);
or UO_911 (O_911,N_49689,N_48603);
and UO_912 (O_912,N_48360,N_49650);
or UO_913 (O_913,N_48422,N_49064);
and UO_914 (O_914,N_48970,N_48775);
or UO_915 (O_915,N_48725,N_49709);
xnor UO_916 (O_916,N_48519,N_48674);
or UO_917 (O_917,N_49621,N_49642);
xnor UO_918 (O_918,N_49370,N_48384);
and UO_919 (O_919,N_48981,N_48920);
nand UO_920 (O_920,N_48472,N_49545);
xnor UO_921 (O_921,N_48625,N_48125);
and UO_922 (O_922,N_49937,N_48794);
and UO_923 (O_923,N_49026,N_48689);
nand UO_924 (O_924,N_48098,N_49654);
nand UO_925 (O_925,N_49099,N_48082);
nand UO_926 (O_926,N_48053,N_49551);
and UO_927 (O_927,N_49678,N_49077);
or UO_928 (O_928,N_48436,N_48539);
nor UO_929 (O_929,N_49453,N_48244);
xor UO_930 (O_930,N_49456,N_49200);
xor UO_931 (O_931,N_48207,N_49297);
nand UO_932 (O_932,N_49499,N_48108);
or UO_933 (O_933,N_49724,N_49274);
or UO_934 (O_934,N_49837,N_48309);
nand UO_935 (O_935,N_49083,N_48536);
or UO_936 (O_936,N_49445,N_48892);
and UO_937 (O_937,N_48432,N_48802);
or UO_938 (O_938,N_48076,N_48418);
or UO_939 (O_939,N_49747,N_49172);
xor UO_940 (O_940,N_49825,N_48569);
or UO_941 (O_941,N_48409,N_48706);
nor UO_942 (O_942,N_49352,N_49341);
or UO_943 (O_943,N_48184,N_49880);
nand UO_944 (O_944,N_48969,N_48785);
nand UO_945 (O_945,N_49735,N_48862);
nor UO_946 (O_946,N_48273,N_48626);
and UO_947 (O_947,N_49411,N_49165);
and UO_948 (O_948,N_48633,N_49212);
xor UO_949 (O_949,N_49287,N_49086);
nand UO_950 (O_950,N_49946,N_49577);
xor UO_951 (O_951,N_48143,N_48898);
xnor UO_952 (O_952,N_49270,N_48978);
nor UO_953 (O_953,N_48246,N_49555);
or UO_954 (O_954,N_49198,N_48103);
and UO_955 (O_955,N_49232,N_48822);
xnor UO_956 (O_956,N_49156,N_49875);
nor UO_957 (O_957,N_48682,N_48151);
xnor UO_958 (O_958,N_49419,N_49943);
xor UO_959 (O_959,N_49745,N_48508);
nand UO_960 (O_960,N_48750,N_49803);
or UO_961 (O_961,N_48114,N_49059);
nand UO_962 (O_962,N_48786,N_48158);
and UO_963 (O_963,N_49606,N_48896);
nor UO_964 (O_964,N_49905,N_49767);
and UO_965 (O_965,N_48908,N_48780);
or UO_966 (O_966,N_49302,N_49818);
and UO_967 (O_967,N_49726,N_49280);
nor UO_968 (O_968,N_49739,N_48034);
nor UO_969 (O_969,N_49617,N_48174);
nand UO_970 (O_970,N_48629,N_48252);
nor UO_971 (O_971,N_49057,N_49631);
nand UO_972 (O_972,N_48837,N_49824);
xnor UO_973 (O_973,N_48095,N_48305);
nor UO_974 (O_974,N_48260,N_49397);
or UO_975 (O_975,N_48507,N_48062);
xor UO_976 (O_976,N_49362,N_48635);
nand UO_977 (O_977,N_49647,N_48995);
xor UO_978 (O_978,N_48145,N_49664);
or UO_979 (O_979,N_48220,N_49870);
or UO_980 (O_980,N_49233,N_49454);
or UO_981 (O_981,N_48702,N_48665);
nor UO_982 (O_982,N_49700,N_49017);
nand UO_983 (O_983,N_48728,N_48487);
nand UO_984 (O_984,N_48194,N_48416);
nand UO_985 (O_985,N_49708,N_48857);
nor UO_986 (O_986,N_49283,N_48358);
or UO_987 (O_987,N_49016,N_48456);
xor UO_988 (O_988,N_48998,N_49622);
and UO_989 (O_989,N_49428,N_48297);
nand UO_990 (O_990,N_49284,N_48412);
nand UO_991 (O_991,N_49403,N_48710);
or UO_992 (O_992,N_48600,N_49168);
nor UO_993 (O_993,N_48021,N_49711);
and UO_994 (O_994,N_48675,N_48294);
nand UO_995 (O_995,N_48375,N_48598);
nand UO_996 (O_996,N_48457,N_49182);
nand UO_997 (O_997,N_48214,N_49548);
nor UO_998 (O_998,N_48046,N_48229);
nand UO_999 (O_999,N_49998,N_48826);
xnor UO_1000 (O_1000,N_48230,N_49238);
nor UO_1001 (O_1001,N_48697,N_49083);
and UO_1002 (O_1002,N_48686,N_49512);
nor UO_1003 (O_1003,N_49437,N_49978);
nor UO_1004 (O_1004,N_49068,N_48817);
nand UO_1005 (O_1005,N_48806,N_48999);
xor UO_1006 (O_1006,N_49865,N_48137);
nor UO_1007 (O_1007,N_48179,N_48694);
nand UO_1008 (O_1008,N_48232,N_48247);
nor UO_1009 (O_1009,N_49824,N_48605);
and UO_1010 (O_1010,N_49415,N_48152);
nor UO_1011 (O_1011,N_49506,N_49902);
xnor UO_1012 (O_1012,N_48779,N_48358);
nor UO_1013 (O_1013,N_49110,N_49989);
or UO_1014 (O_1014,N_48918,N_49371);
and UO_1015 (O_1015,N_48479,N_48883);
and UO_1016 (O_1016,N_49194,N_48234);
xnor UO_1017 (O_1017,N_49439,N_48721);
or UO_1018 (O_1018,N_49858,N_48926);
nor UO_1019 (O_1019,N_49816,N_48243);
and UO_1020 (O_1020,N_49125,N_49704);
xnor UO_1021 (O_1021,N_49634,N_49186);
and UO_1022 (O_1022,N_48490,N_49085);
and UO_1023 (O_1023,N_49218,N_49452);
nor UO_1024 (O_1024,N_49481,N_49333);
xnor UO_1025 (O_1025,N_49201,N_48898);
nor UO_1026 (O_1026,N_48035,N_49108);
or UO_1027 (O_1027,N_49666,N_48249);
nor UO_1028 (O_1028,N_49406,N_48661);
xor UO_1029 (O_1029,N_49525,N_49424);
xor UO_1030 (O_1030,N_49824,N_48095);
nand UO_1031 (O_1031,N_48467,N_48278);
and UO_1032 (O_1032,N_49060,N_48154);
and UO_1033 (O_1033,N_48113,N_48391);
and UO_1034 (O_1034,N_48847,N_49841);
nor UO_1035 (O_1035,N_48278,N_49682);
or UO_1036 (O_1036,N_49124,N_49663);
xor UO_1037 (O_1037,N_48668,N_48792);
nor UO_1038 (O_1038,N_48728,N_49656);
and UO_1039 (O_1039,N_48672,N_48743);
nand UO_1040 (O_1040,N_48823,N_49777);
nand UO_1041 (O_1041,N_49107,N_48441);
and UO_1042 (O_1042,N_49008,N_48512);
nand UO_1043 (O_1043,N_48127,N_49465);
nor UO_1044 (O_1044,N_49024,N_49462);
xor UO_1045 (O_1045,N_49055,N_49228);
nand UO_1046 (O_1046,N_48804,N_49334);
xor UO_1047 (O_1047,N_49190,N_48378);
or UO_1048 (O_1048,N_49991,N_48269);
and UO_1049 (O_1049,N_49690,N_49599);
nand UO_1050 (O_1050,N_49071,N_48399);
nor UO_1051 (O_1051,N_48237,N_48112);
xor UO_1052 (O_1052,N_49241,N_48853);
xor UO_1053 (O_1053,N_48995,N_48686);
or UO_1054 (O_1054,N_49660,N_49274);
or UO_1055 (O_1055,N_49782,N_49929);
or UO_1056 (O_1056,N_48463,N_48885);
or UO_1057 (O_1057,N_48425,N_49568);
and UO_1058 (O_1058,N_48571,N_49298);
xor UO_1059 (O_1059,N_48393,N_49317);
xnor UO_1060 (O_1060,N_49901,N_48176);
nor UO_1061 (O_1061,N_49985,N_48460);
or UO_1062 (O_1062,N_48079,N_49027);
xor UO_1063 (O_1063,N_49198,N_49776);
and UO_1064 (O_1064,N_48748,N_48152);
nor UO_1065 (O_1065,N_48973,N_48802);
nor UO_1066 (O_1066,N_49345,N_49348);
nor UO_1067 (O_1067,N_48273,N_49057);
and UO_1068 (O_1068,N_49576,N_48649);
or UO_1069 (O_1069,N_48644,N_49834);
xnor UO_1070 (O_1070,N_48367,N_49013);
nor UO_1071 (O_1071,N_49977,N_48033);
nand UO_1072 (O_1072,N_48321,N_48948);
nor UO_1073 (O_1073,N_49166,N_48523);
nor UO_1074 (O_1074,N_49081,N_48641);
nor UO_1075 (O_1075,N_49771,N_48464);
xnor UO_1076 (O_1076,N_48989,N_49669);
or UO_1077 (O_1077,N_49692,N_48776);
nor UO_1078 (O_1078,N_49615,N_49766);
nor UO_1079 (O_1079,N_48273,N_48962);
or UO_1080 (O_1080,N_49161,N_48231);
or UO_1081 (O_1081,N_48812,N_48052);
and UO_1082 (O_1082,N_48236,N_49249);
nor UO_1083 (O_1083,N_49601,N_48090);
and UO_1084 (O_1084,N_48279,N_49731);
xnor UO_1085 (O_1085,N_48277,N_48679);
xor UO_1086 (O_1086,N_49650,N_48914);
and UO_1087 (O_1087,N_49160,N_49320);
and UO_1088 (O_1088,N_48262,N_48998);
or UO_1089 (O_1089,N_48232,N_49859);
or UO_1090 (O_1090,N_49974,N_48072);
nand UO_1091 (O_1091,N_49908,N_49631);
nor UO_1092 (O_1092,N_48626,N_48865);
or UO_1093 (O_1093,N_49878,N_49347);
and UO_1094 (O_1094,N_49503,N_48182);
xnor UO_1095 (O_1095,N_49586,N_49650);
nor UO_1096 (O_1096,N_49473,N_48031);
and UO_1097 (O_1097,N_48054,N_49175);
and UO_1098 (O_1098,N_48464,N_49187);
xnor UO_1099 (O_1099,N_48551,N_48338);
xor UO_1100 (O_1100,N_48524,N_48375);
nand UO_1101 (O_1101,N_48270,N_49536);
or UO_1102 (O_1102,N_49452,N_48781);
or UO_1103 (O_1103,N_49904,N_49446);
nand UO_1104 (O_1104,N_49191,N_48001);
nand UO_1105 (O_1105,N_48028,N_48953);
nand UO_1106 (O_1106,N_49190,N_49243);
and UO_1107 (O_1107,N_49904,N_49116);
nand UO_1108 (O_1108,N_48500,N_49841);
or UO_1109 (O_1109,N_49750,N_49055);
and UO_1110 (O_1110,N_49056,N_48923);
and UO_1111 (O_1111,N_48655,N_48648);
xnor UO_1112 (O_1112,N_48580,N_48323);
nand UO_1113 (O_1113,N_48489,N_49607);
nor UO_1114 (O_1114,N_48353,N_48824);
nor UO_1115 (O_1115,N_49212,N_48351);
nor UO_1116 (O_1116,N_49448,N_49030);
nor UO_1117 (O_1117,N_49547,N_49439);
or UO_1118 (O_1118,N_48710,N_48792);
or UO_1119 (O_1119,N_49320,N_48389);
and UO_1120 (O_1120,N_48299,N_49839);
nand UO_1121 (O_1121,N_49084,N_49285);
or UO_1122 (O_1122,N_48054,N_48597);
nor UO_1123 (O_1123,N_48733,N_48426);
xor UO_1124 (O_1124,N_49048,N_49965);
xnor UO_1125 (O_1125,N_48191,N_48236);
nand UO_1126 (O_1126,N_49302,N_49536);
xor UO_1127 (O_1127,N_48891,N_48110);
nor UO_1128 (O_1128,N_49273,N_48754);
nand UO_1129 (O_1129,N_49671,N_49769);
or UO_1130 (O_1130,N_49310,N_49454);
or UO_1131 (O_1131,N_48953,N_49439);
and UO_1132 (O_1132,N_48859,N_49120);
nand UO_1133 (O_1133,N_48558,N_48046);
nor UO_1134 (O_1134,N_48687,N_49282);
xor UO_1135 (O_1135,N_48096,N_49677);
nand UO_1136 (O_1136,N_48404,N_48782);
or UO_1137 (O_1137,N_49737,N_49036);
and UO_1138 (O_1138,N_49824,N_48246);
nor UO_1139 (O_1139,N_48321,N_49182);
xnor UO_1140 (O_1140,N_48663,N_48261);
xnor UO_1141 (O_1141,N_49814,N_49697);
or UO_1142 (O_1142,N_48365,N_48267);
and UO_1143 (O_1143,N_48252,N_49126);
nand UO_1144 (O_1144,N_48737,N_49937);
or UO_1145 (O_1145,N_49955,N_49182);
or UO_1146 (O_1146,N_49662,N_49661);
or UO_1147 (O_1147,N_49512,N_49936);
xor UO_1148 (O_1148,N_49698,N_49510);
nor UO_1149 (O_1149,N_49702,N_49831);
and UO_1150 (O_1150,N_49009,N_48043);
and UO_1151 (O_1151,N_48092,N_49908);
and UO_1152 (O_1152,N_49257,N_48956);
nor UO_1153 (O_1153,N_48744,N_48381);
nand UO_1154 (O_1154,N_48091,N_48621);
nor UO_1155 (O_1155,N_48619,N_49572);
or UO_1156 (O_1156,N_48546,N_49949);
nor UO_1157 (O_1157,N_49618,N_48418);
xnor UO_1158 (O_1158,N_49963,N_48336);
nor UO_1159 (O_1159,N_49208,N_48458);
and UO_1160 (O_1160,N_49367,N_48765);
nor UO_1161 (O_1161,N_48596,N_48176);
or UO_1162 (O_1162,N_48761,N_49057);
nor UO_1163 (O_1163,N_49446,N_48749);
nand UO_1164 (O_1164,N_49422,N_49206);
nand UO_1165 (O_1165,N_48187,N_49168);
xnor UO_1166 (O_1166,N_49132,N_49509);
xor UO_1167 (O_1167,N_49382,N_49550);
xor UO_1168 (O_1168,N_48568,N_49135);
nand UO_1169 (O_1169,N_48021,N_48037);
nor UO_1170 (O_1170,N_48888,N_49857);
or UO_1171 (O_1171,N_49446,N_49130);
nand UO_1172 (O_1172,N_49008,N_49964);
or UO_1173 (O_1173,N_48928,N_48473);
xnor UO_1174 (O_1174,N_48798,N_48159);
xnor UO_1175 (O_1175,N_48043,N_48618);
and UO_1176 (O_1176,N_49224,N_49788);
xor UO_1177 (O_1177,N_49879,N_49343);
or UO_1178 (O_1178,N_48742,N_48555);
xnor UO_1179 (O_1179,N_48883,N_49171);
and UO_1180 (O_1180,N_49304,N_49575);
xor UO_1181 (O_1181,N_48854,N_49525);
nand UO_1182 (O_1182,N_49288,N_49946);
nor UO_1183 (O_1183,N_48877,N_48564);
and UO_1184 (O_1184,N_49133,N_49030);
nor UO_1185 (O_1185,N_49326,N_48082);
or UO_1186 (O_1186,N_49336,N_49782);
nor UO_1187 (O_1187,N_48667,N_49835);
nor UO_1188 (O_1188,N_49944,N_48404);
xnor UO_1189 (O_1189,N_48893,N_48830);
xor UO_1190 (O_1190,N_48816,N_49524);
nand UO_1191 (O_1191,N_48623,N_48983);
and UO_1192 (O_1192,N_49446,N_48549);
and UO_1193 (O_1193,N_49465,N_49669);
xor UO_1194 (O_1194,N_49535,N_48768);
nand UO_1195 (O_1195,N_49111,N_48106);
xnor UO_1196 (O_1196,N_49141,N_49932);
nand UO_1197 (O_1197,N_49206,N_48657);
nor UO_1198 (O_1198,N_49716,N_48845);
and UO_1199 (O_1199,N_49906,N_49257);
xor UO_1200 (O_1200,N_49476,N_49478);
nand UO_1201 (O_1201,N_49110,N_49147);
or UO_1202 (O_1202,N_49316,N_48562);
nand UO_1203 (O_1203,N_49270,N_49614);
nand UO_1204 (O_1204,N_49661,N_48973);
and UO_1205 (O_1205,N_49539,N_48674);
nand UO_1206 (O_1206,N_48441,N_49918);
and UO_1207 (O_1207,N_48324,N_49444);
nor UO_1208 (O_1208,N_49705,N_48131);
xor UO_1209 (O_1209,N_49511,N_48903);
and UO_1210 (O_1210,N_49584,N_48138);
nand UO_1211 (O_1211,N_48506,N_48714);
nand UO_1212 (O_1212,N_48701,N_49721);
nand UO_1213 (O_1213,N_48052,N_49956);
nor UO_1214 (O_1214,N_49770,N_49492);
nor UO_1215 (O_1215,N_48805,N_49666);
nor UO_1216 (O_1216,N_49838,N_49235);
or UO_1217 (O_1217,N_49683,N_48772);
and UO_1218 (O_1218,N_49494,N_48508);
xnor UO_1219 (O_1219,N_49499,N_49554);
nand UO_1220 (O_1220,N_49716,N_49157);
nand UO_1221 (O_1221,N_48323,N_48587);
xor UO_1222 (O_1222,N_48435,N_48935);
or UO_1223 (O_1223,N_48697,N_49686);
nand UO_1224 (O_1224,N_48724,N_48698);
and UO_1225 (O_1225,N_49036,N_49211);
xnor UO_1226 (O_1226,N_49494,N_49493);
xnor UO_1227 (O_1227,N_48181,N_48622);
nor UO_1228 (O_1228,N_49879,N_48217);
or UO_1229 (O_1229,N_49070,N_49942);
and UO_1230 (O_1230,N_48278,N_48829);
or UO_1231 (O_1231,N_48808,N_48581);
xor UO_1232 (O_1232,N_49516,N_48511);
nor UO_1233 (O_1233,N_49575,N_49468);
nor UO_1234 (O_1234,N_49809,N_49890);
xor UO_1235 (O_1235,N_48529,N_49003);
nor UO_1236 (O_1236,N_48963,N_48017);
and UO_1237 (O_1237,N_48711,N_48992);
or UO_1238 (O_1238,N_48033,N_49548);
nand UO_1239 (O_1239,N_49638,N_48598);
nand UO_1240 (O_1240,N_48380,N_48658);
or UO_1241 (O_1241,N_48030,N_48283);
nor UO_1242 (O_1242,N_48698,N_48718);
xor UO_1243 (O_1243,N_49834,N_49338);
or UO_1244 (O_1244,N_49995,N_49963);
and UO_1245 (O_1245,N_49743,N_49394);
and UO_1246 (O_1246,N_48009,N_48169);
nand UO_1247 (O_1247,N_48739,N_49969);
or UO_1248 (O_1248,N_49233,N_48525);
and UO_1249 (O_1249,N_48367,N_48462);
nor UO_1250 (O_1250,N_49051,N_48535);
or UO_1251 (O_1251,N_48253,N_48952);
and UO_1252 (O_1252,N_48395,N_49914);
nand UO_1253 (O_1253,N_48896,N_48500);
nand UO_1254 (O_1254,N_49137,N_48251);
xor UO_1255 (O_1255,N_48709,N_49719);
xor UO_1256 (O_1256,N_48559,N_48520);
xnor UO_1257 (O_1257,N_49732,N_49105);
nor UO_1258 (O_1258,N_48127,N_49842);
xor UO_1259 (O_1259,N_49623,N_49545);
or UO_1260 (O_1260,N_49896,N_49959);
nand UO_1261 (O_1261,N_49011,N_48524);
xnor UO_1262 (O_1262,N_49336,N_48349);
or UO_1263 (O_1263,N_49360,N_49527);
and UO_1264 (O_1264,N_48637,N_49858);
nor UO_1265 (O_1265,N_48879,N_48733);
or UO_1266 (O_1266,N_48871,N_49774);
xor UO_1267 (O_1267,N_49161,N_49577);
and UO_1268 (O_1268,N_48216,N_48926);
nor UO_1269 (O_1269,N_48953,N_49060);
and UO_1270 (O_1270,N_48064,N_49632);
nand UO_1271 (O_1271,N_48303,N_48328);
nand UO_1272 (O_1272,N_48729,N_49382);
or UO_1273 (O_1273,N_49070,N_49091);
nor UO_1274 (O_1274,N_48953,N_48335);
xnor UO_1275 (O_1275,N_49385,N_49178);
nor UO_1276 (O_1276,N_48850,N_49722);
nor UO_1277 (O_1277,N_49754,N_48460);
xnor UO_1278 (O_1278,N_48508,N_48918);
xnor UO_1279 (O_1279,N_49765,N_48364);
or UO_1280 (O_1280,N_48387,N_49376);
and UO_1281 (O_1281,N_48005,N_48123);
or UO_1282 (O_1282,N_48395,N_49368);
xnor UO_1283 (O_1283,N_48027,N_49673);
nand UO_1284 (O_1284,N_48664,N_48088);
nand UO_1285 (O_1285,N_49663,N_48914);
xor UO_1286 (O_1286,N_48919,N_48435);
nand UO_1287 (O_1287,N_49847,N_48465);
nand UO_1288 (O_1288,N_48932,N_49496);
and UO_1289 (O_1289,N_49007,N_48562);
nand UO_1290 (O_1290,N_49509,N_48296);
nand UO_1291 (O_1291,N_49853,N_49958);
and UO_1292 (O_1292,N_48115,N_49179);
and UO_1293 (O_1293,N_48627,N_48681);
nand UO_1294 (O_1294,N_49972,N_49213);
nor UO_1295 (O_1295,N_49194,N_48455);
nand UO_1296 (O_1296,N_49368,N_49565);
xnor UO_1297 (O_1297,N_48364,N_48137);
nand UO_1298 (O_1298,N_48564,N_49696);
or UO_1299 (O_1299,N_48060,N_49145);
nand UO_1300 (O_1300,N_49374,N_49843);
or UO_1301 (O_1301,N_49916,N_48216);
or UO_1302 (O_1302,N_49138,N_49018);
or UO_1303 (O_1303,N_49632,N_48125);
or UO_1304 (O_1304,N_49926,N_48951);
nand UO_1305 (O_1305,N_49491,N_49419);
and UO_1306 (O_1306,N_49735,N_48898);
or UO_1307 (O_1307,N_48016,N_49824);
nand UO_1308 (O_1308,N_48485,N_48577);
xor UO_1309 (O_1309,N_48232,N_48313);
nor UO_1310 (O_1310,N_48684,N_49846);
nand UO_1311 (O_1311,N_49009,N_48126);
or UO_1312 (O_1312,N_48564,N_49805);
or UO_1313 (O_1313,N_49926,N_48736);
or UO_1314 (O_1314,N_48001,N_48060);
nor UO_1315 (O_1315,N_48821,N_48325);
or UO_1316 (O_1316,N_49429,N_49012);
xor UO_1317 (O_1317,N_48347,N_48915);
or UO_1318 (O_1318,N_48251,N_49641);
nor UO_1319 (O_1319,N_49606,N_49851);
and UO_1320 (O_1320,N_49023,N_48775);
xor UO_1321 (O_1321,N_49020,N_48847);
nand UO_1322 (O_1322,N_49248,N_49149);
nand UO_1323 (O_1323,N_49372,N_48320);
nand UO_1324 (O_1324,N_48778,N_48125);
and UO_1325 (O_1325,N_48995,N_48475);
and UO_1326 (O_1326,N_49666,N_48476);
and UO_1327 (O_1327,N_49934,N_49268);
nor UO_1328 (O_1328,N_48450,N_48108);
xnor UO_1329 (O_1329,N_48058,N_49042);
nor UO_1330 (O_1330,N_49318,N_49003);
xnor UO_1331 (O_1331,N_48259,N_48939);
nand UO_1332 (O_1332,N_48161,N_48260);
nor UO_1333 (O_1333,N_49335,N_49817);
xnor UO_1334 (O_1334,N_49585,N_48040);
or UO_1335 (O_1335,N_48797,N_48250);
xor UO_1336 (O_1336,N_48369,N_48259);
and UO_1337 (O_1337,N_48860,N_48329);
or UO_1338 (O_1338,N_48475,N_48480);
nor UO_1339 (O_1339,N_49342,N_49467);
and UO_1340 (O_1340,N_49107,N_49434);
or UO_1341 (O_1341,N_49341,N_49855);
nand UO_1342 (O_1342,N_49462,N_49584);
xnor UO_1343 (O_1343,N_49629,N_48356);
or UO_1344 (O_1344,N_48100,N_49863);
nor UO_1345 (O_1345,N_48748,N_48010);
nand UO_1346 (O_1346,N_49175,N_48088);
and UO_1347 (O_1347,N_49292,N_48108);
nor UO_1348 (O_1348,N_49934,N_49293);
or UO_1349 (O_1349,N_49594,N_48050);
xor UO_1350 (O_1350,N_49111,N_49105);
nand UO_1351 (O_1351,N_49017,N_48400);
nand UO_1352 (O_1352,N_49444,N_48257);
or UO_1353 (O_1353,N_49971,N_48094);
nor UO_1354 (O_1354,N_49851,N_49808);
nor UO_1355 (O_1355,N_48893,N_49851);
nor UO_1356 (O_1356,N_49499,N_48401);
nor UO_1357 (O_1357,N_48797,N_48171);
and UO_1358 (O_1358,N_49746,N_49784);
or UO_1359 (O_1359,N_48507,N_48056);
or UO_1360 (O_1360,N_48203,N_48297);
xor UO_1361 (O_1361,N_49850,N_48970);
nand UO_1362 (O_1362,N_49636,N_48827);
xor UO_1363 (O_1363,N_48097,N_49338);
and UO_1364 (O_1364,N_49002,N_48836);
and UO_1365 (O_1365,N_49209,N_49325);
xnor UO_1366 (O_1366,N_49730,N_48218);
xor UO_1367 (O_1367,N_49987,N_49992);
nand UO_1368 (O_1368,N_49287,N_48905);
xnor UO_1369 (O_1369,N_49990,N_49313);
nand UO_1370 (O_1370,N_49176,N_49136);
and UO_1371 (O_1371,N_49865,N_48426);
nand UO_1372 (O_1372,N_48229,N_48919);
nor UO_1373 (O_1373,N_49679,N_48518);
or UO_1374 (O_1374,N_48278,N_49781);
nand UO_1375 (O_1375,N_49185,N_49903);
nand UO_1376 (O_1376,N_48817,N_49494);
xor UO_1377 (O_1377,N_48236,N_48250);
nand UO_1378 (O_1378,N_49245,N_49572);
and UO_1379 (O_1379,N_49212,N_48469);
xor UO_1380 (O_1380,N_48770,N_49412);
nand UO_1381 (O_1381,N_48877,N_49465);
xnor UO_1382 (O_1382,N_48488,N_49538);
nand UO_1383 (O_1383,N_48027,N_48390);
or UO_1384 (O_1384,N_48145,N_49604);
xor UO_1385 (O_1385,N_49348,N_49178);
nor UO_1386 (O_1386,N_49732,N_49540);
xnor UO_1387 (O_1387,N_49680,N_49609);
xor UO_1388 (O_1388,N_49294,N_48330);
nand UO_1389 (O_1389,N_48232,N_48755);
xor UO_1390 (O_1390,N_49919,N_48188);
or UO_1391 (O_1391,N_49267,N_48338);
nor UO_1392 (O_1392,N_49217,N_48532);
and UO_1393 (O_1393,N_49453,N_49407);
and UO_1394 (O_1394,N_48149,N_48805);
or UO_1395 (O_1395,N_49799,N_48676);
nand UO_1396 (O_1396,N_49518,N_49901);
and UO_1397 (O_1397,N_48556,N_49066);
xor UO_1398 (O_1398,N_48374,N_49014);
or UO_1399 (O_1399,N_48836,N_48244);
xnor UO_1400 (O_1400,N_49049,N_49446);
or UO_1401 (O_1401,N_49203,N_49577);
nand UO_1402 (O_1402,N_49465,N_49281);
and UO_1403 (O_1403,N_48314,N_49789);
and UO_1404 (O_1404,N_48090,N_49569);
nor UO_1405 (O_1405,N_49912,N_49449);
nor UO_1406 (O_1406,N_49685,N_49698);
xor UO_1407 (O_1407,N_49974,N_48006);
and UO_1408 (O_1408,N_48757,N_49133);
or UO_1409 (O_1409,N_49365,N_48707);
nor UO_1410 (O_1410,N_49697,N_48343);
or UO_1411 (O_1411,N_49734,N_49233);
xnor UO_1412 (O_1412,N_48087,N_48842);
and UO_1413 (O_1413,N_48304,N_49461);
nor UO_1414 (O_1414,N_48437,N_48277);
and UO_1415 (O_1415,N_49493,N_49825);
xor UO_1416 (O_1416,N_48441,N_48850);
nand UO_1417 (O_1417,N_49691,N_48431);
or UO_1418 (O_1418,N_48971,N_49038);
nand UO_1419 (O_1419,N_48144,N_49998);
or UO_1420 (O_1420,N_48037,N_49102);
xor UO_1421 (O_1421,N_48021,N_49050);
nor UO_1422 (O_1422,N_48596,N_49555);
nand UO_1423 (O_1423,N_48737,N_49293);
or UO_1424 (O_1424,N_49281,N_49181);
and UO_1425 (O_1425,N_48776,N_48900);
or UO_1426 (O_1426,N_49153,N_49018);
nor UO_1427 (O_1427,N_48690,N_49200);
nor UO_1428 (O_1428,N_49621,N_49705);
or UO_1429 (O_1429,N_49704,N_49910);
nor UO_1430 (O_1430,N_49185,N_48297);
nand UO_1431 (O_1431,N_48717,N_48678);
xnor UO_1432 (O_1432,N_48104,N_48560);
xnor UO_1433 (O_1433,N_48627,N_48673);
or UO_1434 (O_1434,N_48889,N_48646);
nand UO_1435 (O_1435,N_49372,N_48994);
xor UO_1436 (O_1436,N_48347,N_49886);
nor UO_1437 (O_1437,N_49363,N_49488);
xnor UO_1438 (O_1438,N_49589,N_49092);
nor UO_1439 (O_1439,N_49613,N_48864);
or UO_1440 (O_1440,N_48327,N_48065);
or UO_1441 (O_1441,N_48714,N_49109);
or UO_1442 (O_1442,N_48642,N_49309);
nor UO_1443 (O_1443,N_48693,N_48143);
nand UO_1444 (O_1444,N_48634,N_48552);
nor UO_1445 (O_1445,N_48188,N_49281);
or UO_1446 (O_1446,N_49675,N_49353);
or UO_1447 (O_1447,N_48703,N_49018);
nand UO_1448 (O_1448,N_49522,N_49220);
nand UO_1449 (O_1449,N_48611,N_49091);
and UO_1450 (O_1450,N_48731,N_49770);
nand UO_1451 (O_1451,N_48399,N_48460);
xor UO_1452 (O_1452,N_49590,N_49066);
nand UO_1453 (O_1453,N_49750,N_48333);
or UO_1454 (O_1454,N_49115,N_49434);
nor UO_1455 (O_1455,N_49082,N_48771);
nor UO_1456 (O_1456,N_48253,N_48979);
xor UO_1457 (O_1457,N_49385,N_49564);
nand UO_1458 (O_1458,N_48294,N_49621);
nand UO_1459 (O_1459,N_48085,N_49019);
xor UO_1460 (O_1460,N_49553,N_48291);
nor UO_1461 (O_1461,N_48947,N_48772);
nor UO_1462 (O_1462,N_49134,N_48328);
and UO_1463 (O_1463,N_48532,N_48860);
and UO_1464 (O_1464,N_48196,N_49905);
nand UO_1465 (O_1465,N_48897,N_49658);
nor UO_1466 (O_1466,N_48143,N_48593);
and UO_1467 (O_1467,N_48437,N_49948);
and UO_1468 (O_1468,N_48771,N_48023);
or UO_1469 (O_1469,N_48010,N_49066);
nor UO_1470 (O_1470,N_48355,N_49937);
nand UO_1471 (O_1471,N_48029,N_49258);
and UO_1472 (O_1472,N_48944,N_48990);
nand UO_1473 (O_1473,N_49532,N_49698);
nor UO_1474 (O_1474,N_48289,N_48384);
xor UO_1475 (O_1475,N_48169,N_49682);
and UO_1476 (O_1476,N_49346,N_48642);
and UO_1477 (O_1477,N_49046,N_49153);
and UO_1478 (O_1478,N_49081,N_49228);
nor UO_1479 (O_1479,N_49708,N_49021);
xnor UO_1480 (O_1480,N_49717,N_48638);
nand UO_1481 (O_1481,N_49097,N_49383);
nand UO_1482 (O_1482,N_48031,N_49564);
or UO_1483 (O_1483,N_49100,N_49646);
xor UO_1484 (O_1484,N_49355,N_48725);
and UO_1485 (O_1485,N_48517,N_49462);
xor UO_1486 (O_1486,N_48812,N_48924);
nor UO_1487 (O_1487,N_49247,N_48279);
or UO_1488 (O_1488,N_49834,N_49395);
nor UO_1489 (O_1489,N_48332,N_49114);
nand UO_1490 (O_1490,N_49733,N_49647);
or UO_1491 (O_1491,N_48269,N_49423);
and UO_1492 (O_1492,N_48714,N_49880);
nor UO_1493 (O_1493,N_49811,N_48114);
nor UO_1494 (O_1494,N_49179,N_49267);
nor UO_1495 (O_1495,N_49209,N_48959);
and UO_1496 (O_1496,N_49574,N_49844);
xnor UO_1497 (O_1497,N_49771,N_48770);
nand UO_1498 (O_1498,N_49745,N_48645);
and UO_1499 (O_1499,N_49509,N_49488);
nor UO_1500 (O_1500,N_49617,N_48708);
and UO_1501 (O_1501,N_49804,N_48443);
nor UO_1502 (O_1502,N_48276,N_49022);
or UO_1503 (O_1503,N_49802,N_48272);
nand UO_1504 (O_1504,N_49437,N_48465);
xor UO_1505 (O_1505,N_48705,N_48107);
nand UO_1506 (O_1506,N_49133,N_49843);
and UO_1507 (O_1507,N_48516,N_49361);
or UO_1508 (O_1508,N_48582,N_48736);
xor UO_1509 (O_1509,N_48188,N_48250);
xor UO_1510 (O_1510,N_49231,N_49089);
xnor UO_1511 (O_1511,N_49997,N_48583);
nand UO_1512 (O_1512,N_49417,N_49879);
xor UO_1513 (O_1513,N_48354,N_48993);
nor UO_1514 (O_1514,N_49316,N_48964);
and UO_1515 (O_1515,N_48078,N_49869);
nor UO_1516 (O_1516,N_48702,N_49939);
nor UO_1517 (O_1517,N_48832,N_49478);
nand UO_1518 (O_1518,N_48532,N_48009);
nor UO_1519 (O_1519,N_48801,N_48394);
and UO_1520 (O_1520,N_48142,N_49723);
and UO_1521 (O_1521,N_49103,N_49866);
xor UO_1522 (O_1522,N_49132,N_49581);
xor UO_1523 (O_1523,N_48126,N_49999);
or UO_1524 (O_1524,N_48219,N_49705);
or UO_1525 (O_1525,N_49370,N_49515);
xnor UO_1526 (O_1526,N_49934,N_48855);
xnor UO_1527 (O_1527,N_48121,N_49565);
nand UO_1528 (O_1528,N_48451,N_49494);
or UO_1529 (O_1529,N_49303,N_48874);
or UO_1530 (O_1530,N_48553,N_48709);
and UO_1531 (O_1531,N_49205,N_48660);
xor UO_1532 (O_1532,N_49691,N_48906);
or UO_1533 (O_1533,N_49102,N_48082);
and UO_1534 (O_1534,N_49980,N_48481);
and UO_1535 (O_1535,N_48911,N_49206);
nor UO_1536 (O_1536,N_49918,N_48501);
nand UO_1537 (O_1537,N_48804,N_49303);
and UO_1538 (O_1538,N_48260,N_48661);
or UO_1539 (O_1539,N_48330,N_49988);
or UO_1540 (O_1540,N_49360,N_49637);
xor UO_1541 (O_1541,N_49647,N_49570);
nor UO_1542 (O_1542,N_48124,N_49035);
nand UO_1543 (O_1543,N_48808,N_48782);
xnor UO_1544 (O_1544,N_49737,N_49562);
or UO_1545 (O_1545,N_48768,N_48705);
xor UO_1546 (O_1546,N_49393,N_48748);
nand UO_1547 (O_1547,N_49281,N_48183);
xor UO_1548 (O_1548,N_49407,N_49187);
and UO_1549 (O_1549,N_49970,N_49139);
nand UO_1550 (O_1550,N_49664,N_49782);
xor UO_1551 (O_1551,N_48247,N_48532);
xnor UO_1552 (O_1552,N_48524,N_48803);
xor UO_1553 (O_1553,N_49432,N_48029);
nand UO_1554 (O_1554,N_49113,N_48362);
nand UO_1555 (O_1555,N_49185,N_48079);
nand UO_1556 (O_1556,N_48691,N_48798);
or UO_1557 (O_1557,N_48194,N_49013);
nand UO_1558 (O_1558,N_49104,N_49718);
nor UO_1559 (O_1559,N_48546,N_48392);
nor UO_1560 (O_1560,N_49634,N_49430);
nand UO_1561 (O_1561,N_48986,N_48554);
nor UO_1562 (O_1562,N_49851,N_49119);
nor UO_1563 (O_1563,N_49066,N_49803);
xnor UO_1564 (O_1564,N_48057,N_49910);
nand UO_1565 (O_1565,N_48817,N_49771);
or UO_1566 (O_1566,N_49009,N_49226);
and UO_1567 (O_1567,N_49819,N_48769);
or UO_1568 (O_1568,N_48954,N_48628);
nor UO_1569 (O_1569,N_48130,N_49493);
xnor UO_1570 (O_1570,N_48079,N_48906);
and UO_1571 (O_1571,N_49772,N_48534);
and UO_1572 (O_1572,N_49843,N_48037);
and UO_1573 (O_1573,N_48267,N_48579);
and UO_1574 (O_1574,N_48636,N_48641);
nor UO_1575 (O_1575,N_49003,N_48863);
xor UO_1576 (O_1576,N_48695,N_49436);
nor UO_1577 (O_1577,N_48536,N_48983);
nand UO_1578 (O_1578,N_48302,N_49432);
or UO_1579 (O_1579,N_49661,N_48085);
nor UO_1580 (O_1580,N_49862,N_49170);
and UO_1581 (O_1581,N_48980,N_49728);
xor UO_1582 (O_1582,N_48958,N_49878);
and UO_1583 (O_1583,N_48199,N_49222);
or UO_1584 (O_1584,N_49125,N_49697);
xor UO_1585 (O_1585,N_49144,N_49495);
and UO_1586 (O_1586,N_49734,N_48296);
nand UO_1587 (O_1587,N_48998,N_48870);
xor UO_1588 (O_1588,N_48303,N_49778);
xnor UO_1589 (O_1589,N_49862,N_48798);
and UO_1590 (O_1590,N_48546,N_48781);
nand UO_1591 (O_1591,N_49821,N_48764);
and UO_1592 (O_1592,N_49770,N_49587);
or UO_1593 (O_1593,N_48964,N_48638);
xor UO_1594 (O_1594,N_49537,N_48365);
and UO_1595 (O_1595,N_48451,N_48864);
nor UO_1596 (O_1596,N_49132,N_48440);
nand UO_1597 (O_1597,N_49888,N_48426);
xnor UO_1598 (O_1598,N_49195,N_48941);
and UO_1599 (O_1599,N_49578,N_49316);
xor UO_1600 (O_1600,N_49328,N_48643);
nand UO_1601 (O_1601,N_49754,N_49484);
and UO_1602 (O_1602,N_49918,N_49993);
nand UO_1603 (O_1603,N_49820,N_48832);
nor UO_1604 (O_1604,N_48866,N_49643);
or UO_1605 (O_1605,N_48868,N_49532);
nand UO_1606 (O_1606,N_48455,N_49004);
xor UO_1607 (O_1607,N_48186,N_49556);
or UO_1608 (O_1608,N_49670,N_48150);
xnor UO_1609 (O_1609,N_49181,N_49666);
xnor UO_1610 (O_1610,N_48803,N_48450);
xor UO_1611 (O_1611,N_48094,N_48864);
or UO_1612 (O_1612,N_49591,N_49130);
xor UO_1613 (O_1613,N_48240,N_48902);
nand UO_1614 (O_1614,N_49853,N_48942);
or UO_1615 (O_1615,N_49676,N_48053);
xnor UO_1616 (O_1616,N_48547,N_48671);
and UO_1617 (O_1617,N_48170,N_49427);
or UO_1618 (O_1618,N_49273,N_48681);
xnor UO_1619 (O_1619,N_48004,N_49667);
nor UO_1620 (O_1620,N_48832,N_49201);
xnor UO_1621 (O_1621,N_48842,N_48048);
nand UO_1622 (O_1622,N_49208,N_48584);
nand UO_1623 (O_1623,N_48202,N_49673);
nand UO_1624 (O_1624,N_48384,N_49132);
and UO_1625 (O_1625,N_48645,N_48895);
nand UO_1626 (O_1626,N_48483,N_49015);
nor UO_1627 (O_1627,N_48040,N_49148);
nor UO_1628 (O_1628,N_49009,N_49202);
nor UO_1629 (O_1629,N_48829,N_48279);
xor UO_1630 (O_1630,N_48176,N_48535);
nor UO_1631 (O_1631,N_49466,N_49628);
nand UO_1632 (O_1632,N_48628,N_48766);
and UO_1633 (O_1633,N_48199,N_49133);
nand UO_1634 (O_1634,N_48244,N_49630);
or UO_1635 (O_1635,N_48745,N_49345);
or UO_1636 (O_1636,N_48785,N_49554);
and UO_1637 (O_1637,N_48756,N_48497);
or UO_1638 (O_1638,N_49803,N_48644);
and UO_1639 (O_1639,N_48094,N_48242);
nor UO_1640 (O_1640,N_49063,N_48988);
nand UO_1641 (O_1641,N_49361,N_48803);
and UO_1642 (O_1642,N_48965,N_48659);
xnor UO_1643 (O_1643,N_49948,N_48897);
nor UO_1644 (O_1644,N_48243,N_49824);
and UO_1645 (O_1645,N_49108,N_49840);
nand UO_1646 (O_1646,N_49721,N_48455);
xor UO_1647 (O_1647,N_48918,N_49640);
nand UO_1648 (O_1648,N_48884,N_48659);
or UO_1649 (O_1649,N_49585,N_48153);
and UO_1650 (O_1650,N_49736,N_49740);
or UO_1651 (O_1651,N_49526,N_49400);
and UO_1652 (O_1652,N_49514,N_48298);
and UO_1653 (O_1653,N_49975,N_49932);
nor UO_1654 (O_1654,N_48063,N_49422);
and UO_1655 (O_1655,N_49589,N_48207);
nor UO_1656 (O_1656,N_49725,N_48120);
and UO_1657 (O_1657,N_49558,N_48448);
nor UO_1658 (O_1658,N_48397,N_49083);
or UO_1659 (O_1659,N_48807,N_48995);
xnor UO_1660 (O_1660,N_49633,N_48563);
or UO_1661 (O_1661,N_48653,N_49791);
nand UO_1662 (O_1662,N_49303,N_48822);
nand UO_1663 (O_1663,N_48336,N_49801);
xor UO_1664 (O_1664,N_48744,N_49218);
nor UO_1665 (O_1665,N_48216,N_48229);
or UO_1666 (O_1666,N_48963,N_49709);
nor UO_1667 (O_1667,N_49636,N_49363);
xnor UO_1668 (O_1668,N_48901,N_49777);
nor UO_1669 (O_1669,N_48210,N_49360);
xnor UO_1670 (O_1670,N_49112,N_48474);
nor UO_1671 (O_1671,N_48236,N_48036);
and UO_1672 (O_1672,N_49684,N_48056);
nand UO_1673 (O_1673,N_48300,N_49109);
nand UO_1674 (O_1674,N_48098,N_48619);
and UO_1675 (O_1675,N_49286,N_48966);
xor UO_1676 (O_1676,N_49219,N_49968);
xnor UO_1677 (O_1677,N_49230,N_49657);
nor UO_1678 (O_1678,N_48269,N_48403);
nand UO_1679 (O_1679,N_48256,N_49600);
xor UO_1680 (O_1680,N_48116,N_49551);
nand UO_1681 (O_1681,N_48437,N_48840);
or UO_1682 (O_1682,N_48210,N_49076);
nand UO_1683 (O_1683,N_48847,N_49879);
nand UO_1684 (O_1684,N_48097,N_48765);
nor UO_1685 (O_1685,N_49091,N_49238);
xor UO_1686 (O_1686,N_48699,N_48579);
nand UO_1687 (O_1687,N_49200,N_48691);
nor UO_1688 (O_1688,N_49575,N_48825);
and UO_1689 (O_1689,N_49907,N_48939);
and UO_1690 (O_1690,N_49126,N_48771);
nand UO_1691 (O_1691,N_48804,N_49373);
nor UO_1692 (O_1692,N_49096,N_48865);
or UO_1693 (O_1693,N_48324,N_48583);
nor UO_1694 (O_1694,N_49748,N_48321);
nand UO_1695 (O_1695,N_48737,N_48230);
xnor UO_1696 (O_1696,N_48270,N_48771);
nor UO_1697 (O_1697,N_48260,N_48083);
or UO_1698 (O_1698,N_49274,N_48308);
nand UO_1699 (O_1699,N_48886,N_48217);
and UO_1700 (O_1700,N_48168,N_48285);
xor UO_1701 (O_1701,N_49075,N_49563);
and UO_1702 (O_1702,N_48983,N_48120);
xnor UO_1703 (O_1703,N_48911,N_48760);
nand UO_1704 (O_1704,N_48039,N_48775);
nor UO_1705 (O_1705,N_49109,N_49870);
xnor UO_1706 (O_1706,N_49305,N_48186);
nand UO_1707 (O_1707,N_48043,N_49299);
or UO_1708 (O_1708,N_49113,N_48878);
nand UO_1709 (O_1709,N_49744,N_48037);
and UO_1710 (O_1710,N_49614,N_49742);
xnor UO_1711 (O_1711,N_48669,N_49068);
or UO_1712 (O_1712,N_48471,N_48463);
or UO_1713 (O_1713,N_48687,N_48265);
and UO_1714 (O_1714,N_48422,N_48849);
or UO_1715 (O_1715,N_48109,N_49249);
nor UO_1716 (O_1716,N_48449,N_49626);
nor UO_1717 (O_1717,N_49385,N_48004);
nand UO_1718 (O_1718,N_48797,N_48491);
or UO_1719 (O_1719,N_48636,N_48582);
and UO_1720 (O_1720,N_49789,N_48498);
nand UO_1721 (O_1721,N_49773,N_48138);
nor UO_1722 (O_1722,N_48548,N_49910);
and UO_1723 (O_1723,N_48269,N_48074);
nand UO_1724 (O_1724,N_48975,N_49877);
nor UO_1725 (O_1725,N_49440,N_49187);
or UO_1726 (O_1726,N_49363,N_49476);
nand UO_1727 (O_1727,N_49189,N_49176);
xor UO_1728 (O_1728,N_49952,N_49868);
and UO_1729 (O_1729,N_48444,N_49437);
xnor UO_1730 (O_1730,N_49242,N_49675);
nand UO_1731 (O_1731,N_49231,N_48245);
or UO_1732 (O_1732,N_48653,N_48738);
and UO_1733 (O_1733,N_48537,N_48032);
and UO_1734 (O_1734,N_48376,N_48280);
nand UO_1735 (O_1735,N_48129,N_49740);
xor UO_1736 (O_1736,N_49359,N_48767);
xor UO_1737 (O_1737,N_49552,N_49858);
or UO_1738 (O_1738,N_49069,N_49480);
and UO_1739 (O_1739,N_48846,N_48894);
xnor UO_1740 (O_1740,N_48901,N_48474);
nor UO_1741 (O_1741,N_48371,N_49881);
and UO_1742 (O_1742,N_48709,N_49350);
nor UO_1743 (O_1743,N_49319,N_49408);
nand UO_1744 (O_1744,N_49274,N_48654);
or UO_1745 (O_1745,N_48385,N_49576);
xor UO_1746 (O_1746,N_49378,N_48327);
and UO_1747 (O_1747,N_48469,N_48681);
and UO_1748 (O_1748,N_48698,N_48827);
nand UO_1749 (O_1749,N_49270,N_48314);
xor UO_1750 (O_1750,N_48335,N_49536);
and UO_1751 (O_1751,N_48264,N_49572);
xor UO_1752 (O_1752,N_49159,N_49881);
nand UO_1753 (O_1753,N_49887,N_49255);
and UO_1754 (O_1754,N_48357,N_48614);
or UO_1755 (O_1755,N_49836,N_48251);
nand UO_1756 (O_1756,N_49813,N_48733);
and UO_1757 (O_1757,N_48022,N_49340);
or UO_1758 (O_1758,N_49303,N_48062);
and UO_1759 (O_1759,N_48791,N_48647);
and UO_1760 (O_1760,N_49164,N_49214);
or UO_1761 (O_1761,N_49794,N_49108);
and UO_1762 (O_1762,N_48664,N_49270);
and UO_1763 (O_1763,N_48037,N_49733);
nor UO_1764 (O_1764,N_49835,N_49421);
and UO_1765 (O_1765,N_49698,N_49560);
xnor UO_1766 (O_1766,N_49888,N_48368);
or UO_1767 (O_1767,N_49980,N_49585);
xnor UO_1768 (O_1768,N_49093,N_48977);
or UO_1769 (O_1769,N_48157,N_48365);
and UO_1770 (O_1770,N_49241,N_49278);
or UO_1771 (O_1771,N_49535,N_49870);
nand UO_1772 (O_1772,N_49730,N_48702);
nor UO_1773 (O_1773,N_48062,N_48940);
nor UO_1774 (O_1774,N_48481,N_49857);
or UO_1775 (O_1775,N_48024,N_48601);
nor UO_1776 (O_1776,N_48088,N_48182);
nor UO_1777 (O_1777,N_49574,N_48692);
nor UO_1778 (O_1778,N_49465,N_48068);
or UO_1779 (O_1779,N_48050,N_49756);
or UO_1780 (O_1780,N_49869,N_49518);
xor UO_1781 (O_1781,N_48942,N_48961);
nand UO_1782 (O_1782,N_48828,N_48659);
and UO_1783 (O_1783,N_49323,N_49688);
nor UO_1784 (O_1784,N_49897,N_49166);
and UO_1785 (O_1785,N_48138,N_48077);
and UO_1786 (O_1786,N_48175,N_49971);
or UO_1787 (O_1787,N_48935,N_48395);
nand UO_1788 (O_1788,N_49354,N_49051);
nand UO_1789 (O_1789,N_48149,N_48547);
nor UO_1790 (O_1790,N_49430,N_49284);
nand UO_1791 (O_1791,N_49740,N_49262);
nand UO_1792 (O_1792,N_48789,N_49656);
and UO_1793 (O_1793,N_49901,N_49808);
or UO_1794 (O_1794,N_49513,N_49945);
nand UO_1795 (O_1795,N_49636,N_48964);
or UO_1796 (O_1796,N_49907,N_48195);
nand UO_1797 (O_1797,N_48887,N_48864);
xor UO_1798 (O_1798,N_49038,N_49622);
or UO_1799 (O_1799,N_48385,N_48628);
and UO_1800 (O_1800,N_48452,N_48374);
or UO_1801 (O_1801,N_49945,N_48199);
and UO_1802 (O_1802,N_49866,N_49602);
nor UO_1803 (O_1803,N_49607,N_48069);
xnor UO_1804 (O_1804,N_48520,N_49420);
or UO_1805 (O_1805,N_48817,N_49618);
nand UO_1806 (O_1806,N_48740,N_49724);
or UO_1807 (O_1807,N_48656,N_49160);
and UO_1808 (O_1808,N_48300,N_48089);
xor UO_1809 (O_1809,N_48354,N_48157);
or UO_1810 (O_1810,N_49571,N_48786);
nor UO_1811 (O_1811,N_49465,N_49728);
or UO_1812 (O_1812,N_48988,N_49644);
nor UO_1813 (O_1813,N_48164,N_49943);
xnor UO_1814 (O_1814,N_49935,N_48401);
nand UO_1815 (O_1815,N_49358,N_49847);
or UO_1816 (O_1816,N_49579,N_48942);
or UO_1817 (O_1817,N_49752,N_49965);
and UO_1818 (O_1818,N_49256,N_48146);
xnor UO_1819 (O_1819,N_49430,N_48476);
and UO_1820 (O_1820,N_49295,N_49104);
or UO_1821 (O_1821,N_48183,N_48466);
nand UO_1822 (O_1822,N_48065,N_49591);
nand UO_1823 (O_1823,N_49488,N_49452);
nor UO_1824 (O_1824,N_49222,N_49338);
nand UO_1825 (O_1825,N_48824,N_48956);
and UO_1826 (O_1826,N_48033,N_49901);
nor UO_1827 (O_1827,N_48647,N_48696);
nand UO_1828 (O_1828,N_48875,N_49840);
nor UO_1829 (O_1829,N_48808,N_48500);
and UO_1830 (O_1830,N_48051,N_49505);
or UO_1831 (O_1831,N_48322,N_48151);
or UO_1832 (O_1832,N_48460,N_49860);
or UO_1833 (O_1833,N_49843,N_48685);
nor UO_1834 (O_1834,N_48673,N_49346);
nor UO_1835 (O_1835,N_49856,N_48288);
xnor UO_1836 (O_1836,N_49061,N_48302);
xnor UO_1837 (O_1837,N_48584,N_48871);
or UO_1838 (O_1838,N_48683,N_49208);
xnor UO_1839 (O_1839,N_48352,N_48306);
and UO_1840 (O_1840,N_49594,N_49180);
and UO_1841 (O_1841,N_49226,N_48673);
or UO_1842 (O_1842,N_49518,N_48666);
nand UO_1843 (O_1843,N_49122,N_48300);
nor UO_1844 (O_1844,N_48494,N_48268);
and UO_1845 (O_1845,N_48809,N_49239);
nor UO_1846 (O_1846,N_49989,N_48713);
nand UO_1847 (O_1847,N_48975,N_48597);
xnor UO_1848 (O_1848,N_48525,N_48231);
nand UO_1849 (O_1849,N_49212,N_48588);
nor UO_1850 (O_1850,N_49103,N_49778);
and UO_1851 (O_1851,N_48636,N_49141);
nor UO_1852 (O_1852,N_49661,N_49385);
xnor UO_1853 (O_1853,N_49880,N_48201);
or UO_1854 (O_1854,N_49581,N_48974);
and UO_1855 (O_1855,N_48882,N_49441);
nand UO_1856 (O_1856,N_49458,N_49405);
and UO_1857 (O_1857,N_48573,N_49549);
nor UO_1858 (O_1858,N_48317,N_49503);
nor UO_1859 (O_1859,N_49038,N_48678);
xnor UO_1860 (O_1860,N_49917,N_49066);
and UO_1861 (O_1861,N_49291,N_49469);
nand UO_1862 (O_1862,N_48626,N_49407);
and UO_1863 (O_1863,N_49373,N_48405);
nor UO_1864 (O_1864,N_49237,N_49236);
nand UO_1865 (O_1865,N_48041,N_49666);
xnor UO_1866 (O_1866,N_48416,N_49609);
nand UO_1867 (O_1867,N_49544,N_49785);
xnor UO_1868 (O_1868,N_48670,N_49180);
or UO_1869 (O_1869,N_48405,N_49732);
and UO_1870 (O_1870,N_49779,N_49996);
and UO_1871 (O_1871,N_48704,N_48515);
xnor UO_1872 (O_1872,N_48668,N_48160);
or UO_1873 (O_1873,N_49234,N_48901);
xor UO_1874 (O_1874,N_49680,N_48166);
or UO_1875 (O_1875,N_48055,N_48999);
or UO_1876 (O_1876,N_49775,N_49791);
or UO_1877 (O_1877,N_48198,N_49487);
nand UO_1878 (O_1878,N_49384,N_49856);
and UO_1879 (O_1879,N_49276,N_49864);
or UO_1880 (O_1880,N_49209,N_49094);
or UO_1881 (O_1881,N_48794,N_48576);
nor UO_1882 (O_1882,N_49868,N_48658);
or UO_1883 (O_1883,N_49889,N_49324);
nand UO_1884 (O_1884,N_49380,N_48034);
and UO_1885 (O_1885,N_49662,N_49594);
or UO_1886 (O_1886,N_48446,N_48355);
nand UO_1887 (O_1887,N_49704,N_49788);
nor UO_1888 (O_1888,N_49919,N_49927);
xor UO_1889 (O_1889,N_48675,N_49380);
and UO_1890 (O_1890,N_49227,N_48462);
or UO_1891 (O_1891,N_49573,N_49514);
nor UO_1892 (O_1892,N_49331,N_48124);
or UO_1893 (O_1893,N_49547,N_49858);
or UO_1894 (O_1894,N_49355,N_48790);
nor UO_1895 (O_1895,N_49092,N_49471);
nor UO_1896 (O_1896,N_48501,N_48181);
and UO_1897 (O_1897,N_49286,N_48610);
or UO_1898 (O_1898,N_48910,N_48888);
and UO_1899 (O_1899,N_48127,N_48228);
or UO_1900 (O_1900,N_49865,N_49472);
and UO_1901 (O_1901,N_49971,N_48455);
and UO_1902 (O_1902,N_48619,N_48718);
nor UO_1903 (O_1903,N_48194,N_49040);
nand UO_1904 (O_1904,N_49352,N_48802);
and UO_1905 (O_1905,N_49065,N_48200);
nor UO_1906 (O_1906,N_48733,N_49941);
or UO_1907 (O_1907,N_48782,N_48090);
or UO_1908 (O_1908,N_49621,N_48492);
and UO_1909 (O_1909,N_49218,N_49940);
nor UO_1910 (O_1910,N_49021,N_49321);
or UO_1911 (O_1911,N_48876,N_49934);
xnor UO_1912 (O_1912,N_49758,N_49315);
nor UO_1913 (O_1913,N_49633,N_49525);
nor UO_1914 (O_1914,N_49054,N_49646);
xor UO_1915 (O_1915,N_48683,N_48173);
or UO_1916 (O_1916,N_48533,N_48989);
and UO_1917 (O_1917,N_48492,N_49137);
and UO_1918 (O_1918,N_49210,N_48898);
nor UO_1919 (O_1919,N_49797,N_49000);
and UO_1920 (O_1920,N_48159,N_48181);
and UO_1921 (O_1921,N_49603,N_49122);
and UO_1922 (O_1922,N_48509,N_48881);
or UO_1923 (O_1923,N_48311,N_49106);
and UO_1924 (O_1924,N_48334,N_48229);
or UO_1925 (O_1925,N_48610,N_49429);
or UO_1926 (O_1926,N_48487,N_49941);
or UO_1927 (O_1927,N_49292,N_48234);
nand UO_1928 (O_1928,N_48901,N_49996);
nand UO_1929 (O_1929,N_49109,N_48916);
and UO_1930 (O_1930,N_49260,N_49329);
nand UO_1931 (O_1931,N_49977,N_48543);
and UO_1932 (O_1932,N_49977,N_49588);
nand UO_1933 (O_1933,N_49456,N_48908);
nor UO_1934 (O_1934,N_49058,N_48883);
nand UO_1935 (O_1935,N_49673,N_49010);
nand UO_1936 (O_1936,N_49525,N_49551);
and UO_1937 (O_1937,N_49642,N_48162);
nor UO_1938 (O_1938,N_49816,N_48390);
or UO_1939 (O_1939,N_49797,N_49705);
and UO_1940 (O_1940,N_48385,N_49242);
nor UO_1941 (O_1941,N_49571,N_48386);
nor UO_1942 (O_1942,N_48977,N_49106);
xor UO_1943 (O_1943,N_49789,N_48709);
nor UO_1944 (O_1944,N_48947,N_49580);
and UO_1945 (O_1945,N_49241,N_49668);
and UO_1946 (O_1946,N_49590,N_48481);
nor UO_1947 (O_1947,N_48513,N_48966);
nand UO_1948 (O_1948,N_49448,N_48210);
xor UO_1949 (O_1949,N_49690,N_49110);
nand UO_1950 (O_1950,N_48189,N_48111);
and UO_1951 (O_1951,N_48529,N_48192);
nand UO_1952 (O_1952,N_49220,N_48901);
and UO_1953 (O_1953,N_49802,N_48718);
nor UO_1954 (O_1954,N_48150,N_49091);
nand UO_1955 (O_1955,N_49770,N_49881);
or UO_1956 (O_1956,N_49838,N_49497);
or UO_1957 (O_1957,N_49053,N_49572);
and UO_1958 (O_1958,N_48669,N_48356);
or UO_1959 (O_1959,N_48726,N_48296);
and UO_1960 (O_1960,N_49641,N_48504);
nor UO_1961 (O_1961,N_48007,N_48196);
and UO_1962 (O_1962,N_48134,N_49902);
and UO_1963 (O_1963,N_48153,N_49081);
nor UO_1964 (O_1964,N_49761,N_48247);
nand UO_1965 (O_1965,N_49396,N_49516);
xnor UO_1966 (O_1966,N_48656,N_48971);
nor UO_1967 (O_1967,N_48673,N_48193);
nor UO_1968 (O_1968,N_49683,N_49987);
nor UO_1969 (O_1969,N_49006,N_48193);
and UO_1970 (O_1970,N_49069,N_48415);
xnor UO_1971 (O_1971,N_49471,N_49821);
nor UO_1972 (O_1972,N_49373,N_48272);
and UO_1973 (O_1973,N_48287,N_49342);
or UO_1974 (O_1974,N_48111,N_49982);
and UO_1975 (O_1975,N_48866,N_49249);
and UO_1976 (O_1976,N_49340,N_48620);
nand UO_1977 (O_1977,N_48359,N_48791);
or UO_1978 (O_1978,N_49064,N_49715);
nand UO_1979 (O_1979,N_48430,N_49825);
and UO_1980 (O_1980,N_49739,N_49300);
or UO_1981 (O_1981,N_49145,N_49258);
nor UO_1982 (O_1982,N_49730,N_48945);
xnor UO_1983 (O_1983,N_49654,N_49067);
xor UO_1984 (O_1984,N_48010,N_48176);
nor UO_1985 (O_1985,N_49946,N_48011);
xor UO_1986 (O_1986,N_49259,N_49750);
or UO_1987 (O_1987,N_49484,N_48731);
and UO_1988 (O_1988,N_49272,N_49688);
nand UO_1989 (O_1989,N_48193,N_49558);
or UO_1990 (O_1990,N_49673,N_49163);
and UO_1991 (O_1991,N_49577,N_49988);
or UO_1992 (O_1992,N_48560,N_49073);
xnor UO_1993 (O_1993,N_48946,N_48827);
nand UO_1994 (O_1994,N_49894,N_48278);
and UO_1995 (O_1995,N_49159,N_48124);
xor UO_1996 (O_1996,N_48714,N_49380);
or UO_1997 (O_1997,N_48889,N_49808);
or UO_1998 (O_1998,N_49866,N_48868);
nor UO_1999 (O_1999,N_49193,N_48272);
xnor UO_2000 (O_2000,N_48776,N_48675);
and UO_2001 (O_2001,N_48704,N_49376);
nor UO_2002 (O_2002,N_48225,N_49570);
and UO_2003 (O_2003,N_49018,N_49911);
nor UO_2004 (O_2004,N_48628,N_49887);
xor UO_2005 (O_2005,N_48755,N_48531);
nand UO_2006 (O_2006,N_49629,N_48897);
and UO_2007 (O_2007,N_49892,N_49741);
xor UO_2008 (O_2008,N_49767,N_49728);
or UO_2009 (O_2009,N_48851,N_48370);
and UO_2010 (O_2010,N_49465,N_48133);
or UO_2011 (O_2011,N_48442,N_49551);
nor UO_2012 (O_2012,N_48235,N_49992);
xnor UO_2013 (O_2013,N_48240,N_48646);
nor UO_2014 (O_2014,N_48377,N_49234);
and UO_2015 (O_2015,N_49928,N_49171);
nand UO_2016 (O_2016,N_49998,N_48234);
nor UO_2017 (O_2017,N_48253,N_49812);
nand UO_2018 (O_2018,N_49038,N_48871);
nand UO_2019 (O_2019,N_49765,N_49359);
and UO_2020 (O_2020,N_48579,N_48708);
nor UO_2021 (O_2021,N_48511,N_49986);
xor UO_2022 (O_2022,N_49426,N_48528);
nand UO_2023 (O_2023,N_48270,N_49058);
and UO_2024 (O_2024,N_48917,N_48969);
nand UO_2025 (O_2025,N_48320,N_49527);
nor UO_2026 (O_2026,N_49714,N_48860);
xor UO_2027 (O_2027,N_49060,N_48107);
or UO_2028 (O_2028,N_48219,N_49287);
nand UO_2029 (O_2029,N_49365,N_48592);
nand UO_2030 (O_2030,N_48441,N_49467);
or UO_2031 (O_2031,N_48346,N_49750);
or UO_2032 (O_2032,N_49550,N_49788);
or UO_2033 (O_2033,N_48042,N_49030);
and UO_2034 (O_2034,N_49088,N_49691);
nand UO_2035 (O_2035,N_49045,N_49971);
and UO_2036 (O_2036,N_49907,N_48158);
nor UO_2037 (O_2037,N_48200,N_48571);
xor UO_2038 (O_2038,N_48411,N_49367);
and UO_2039 (O_2039,N_48438,N_49227);
and UO_2040 (O_2040,N_49594,N_48487);
xor UO_2041 (O_2041,N_49393,N_48049);
xnor UO_2042 (O_2042,N_48375,N_48311);
xnor UO_2043 (O_2043,N_48045,N_48514);
xnor UO_2044 (O_2044,N_49046,N_48624);
and UO_2045 (O_2045,N_49390,N_48405);
or UO_2046 (O_2046,N_48483,N_48854);
or UO_2047 (O_2047,N_49713,N_49165);
or UO_2048 (O_2048,N_49273,N_49543);
xnor UO_2049 (O_2049,N_48861,N_48737);
nor UO_2050 (O_2050,N_49423,N_48772);
nand UO_2051 (O_2051,N_48627,N_49879);
xnor UO_2052 (O_2052,N_49244,N_48083);
xor UO_2053 (O_2053,N_49563,N_49006);
or UO_2054 (O_2054,N_48476,N_49083);
nand UO_2055 (O_2055,N_48700,N_48551);
and UO_2056 (O_2056,N_49052,N_49275);
xnor UO_2057 (O_2057,N_49233,N_49085);
and UO_2058 (O_2058,N_49625,N_48383);
nor UO_2059 (O_2059,N_48230,N_48741);
and UO_2060 (O_2060,N_48353,N_49298);
xor UO_2061 (O_2061,N_48841,N_49826);
and UO_2062 (O_2062,N_48412,N_48832);
xor UO_2063 (O_2063,N_49005,N_49782);
or UO_2064 (O_2064,N_49764,N_49769);
or UO_2065 (O_2065,N_49074,N_48428);
nor UO_2066 (O_2066,N_49910,N_48016);
and UO_2067 (O_2067,N_48774,N_48698);
nand UO_2068 (O_2068,N_48040,N_49902);
xor UO_2069 (O_2069,N_48395,N_49600);
xnor UO_2070 (O_2070,N_49602,N_49673);
and UO_2071 (O_2071,N_48025,N_49410);
or UO_2072 (O_2072,N_48288,N_49742);
and UO_2073 (O_2073,N_49537,N_49976);
xor UO_2074 (O_2074,N_48438,N_49943);
nand UO_2075 (O_2075,N_49621,N_49429);
or UO_2076 (O_2076,N_49591,N_48162);
or UO_2077 (O_2077,N_49506,N_49557);
nand UO_2078 (O_2078,N_49878,N_48295);
xnor UO_2079 (O_2079,N_49321,N_48578);
nand UO_2080 (O_2080,N_48925,N_49558);
xnor UO_2081 (O_2081,N_49093,N_49345);
nor UO_2082 (O_2082,N_48249,N_48166);
nor UO_2083 (O_2083,N_48331,N_48615);
nor UO_2084 (O_2084,N_48372,N_49813);
xnor UO_2085 (O_2085,N_48520,N_48259);
nor UO_2086 (O_2086,N_49187,N_48580);
and UO_2087 (O_2087,N_48190,N_49391);
or UO_2088 (O_2088,N_49178,N_49286);
nand UO_2089 (O_2089,N_48196,N_48908);
xnor UO_2090 (O_2090,N_48065,N_49863);
and UO_2091 (O_2091,N_49736,N_48349);
xor UO_2092 (O_2092,N_48529,N_49819);
xor UO_2093 (O_2093,N_48795,N_48587);
nor UO_2094 (O_2094,N_49816,N_49926);
and UO_2095 (O_2095,N_49528,N_49945);
or UO_2096 (O_2096,N_49214,N_48048);
and UO_2097 (O_2097,N_49738,N_49765);
and UO_2098 (O_2098,N_49973,N_49609);
xnor UO_2099 (O_2099,N_49147,N_49075);
nor UO_2100 (O_2100,N_48539,N_48649);
nor UO_2101 (O_2101,N_49103,N_49007);
nand UO_2102 (O_2102,N_48802,N_49221);
or UO_2103 (O_2103,N_48092,N_48434);
nand UO_2104 (O_2104,N_48647,N_49191);
or UO_2105 (O_2105,N_49936,N_48210);
nand UO_2106 (O_2106,N_49584,N_49062);
nand UO_2107 (O_2107,N_48475,N_49990);
and UO_2108 (O_2108,N_49225,N_48232);
xnor UO_2109 (O_2109,N_49764,N_48917);
xnor UO_2110 (O_2110,N_48555,N_48576);
nor UO_2111 (O_2111,N_48108,N_49705);
or UO_2112 (O_2112,N_49669,N_48767);
nor UO_2113 (O_2113,N_49877,N_49890);
nand UO_2114 (O_2114,N_49244,N_48252);
and UO_2115 (O_2115,N_49543,N_48928);
nand UO_2116 (O_2116,N_48417,N_49749);
nor UO_2117 (O_2117,N_49675,N_49786);
or UO_2118 (O_2118,N_49400,N_49742);
and UO_2119 (O_2119,N_48367,N_48219);
and UO_2120 (O_2120,N_48398,N_48635);
and UO_2121 (O_2121,N_49045,N_49576);
nand UO_2122 (O_2122,N_48098,N_49769);
and UO_2123 (O_2123,N_49473,N_49625);
xor UO_2124 (O_2124,N_48761,N_49060);
nand UO_2125 (O_2125,N_48255,N_48308);
and UO_2126 (O_2126,N_49435,N_48621);
xnor UO_2127 (O_2127,N_48760,N_49960);
nand UO_2128 (O_2128,N_48088,N_49385);
nor UO_2129 (O_2129,N_49773,N_48707);
nand UO_2130 (O_2130,N_48480,N_48384);
and UO_2131 (O_2131,N_49472,N_49633);
or UO_2132 (O_2132,N_48734,N_48791);
nand UO_2133 (O_2133,N_48770,N_49053);
nand UO_2134 (O_2134,N_48961,N_49840);
xor UO_2135 (O_2135,N_48175,N_49574);
or UO_2136 (O_2136,N_49256,N_48705);
or UO_2137 (O_2137,N_48490,N_49152);
and UO_2138 (O_2138,N_49224,N_49248);
and UO_2139 (O_2139,N_48009,N_49656);
xor UO_2140 (O_2140,N_48789,N_48893);
nand UO_2141 (O_2141,N_49258,N_48816);
or UO_2142 (O_2142,N_48479,N_49560);
or UO_2143 (O_2143,N_48001,N_49186);
xor UO_2144 (O_2144,N_49224,N_48945);
nand UO_2145 (O_2145,N_49034,N_48671);
nand UO_2146 (O_2146,N_49501,N_48913);
nor UO_2147 (O_2147,N_48423,N_48344);
nor UO_2148 (O_2148,N_48760,N_48823);
and UO_2149 (O_2149,N_49329,N_48242);
and UO_2150 (O_2150,N_49892,N_49549);
and UO_2151 (O_2151,N_48681,N_49494);
and UO_2152 (O_2152,N_49158,N_49219);
xor UO_2153 (O_2153,N_49873,N_49423);
nand UO_2154 (O_2154,N_48226,N_48568);
xnor UO_2155 (O_2155,N_48065,N_48676);
nand UO_2156 (O_2156,N_48287,N_48663);
nand UO_2157 (O_2157,N_49529,N_49801);
nand UO_2158 (O_2158,N_48574,N_49728);
or UO_2159 (O_2159,N_48204,N_49360);
and UO_2160 (O_2160,N_48823,N_48026);
nor UO_2161 (O_2161,N_49817,N_48886);
and UO_2162 (O_2162,N_49552,N_48366);
nor UO_2163 (O_2163,N_49461,N_49162);
nand UO_2164 (O_2164,N_48400,N_49729);
nor UO_2165 (O_2165,N_48676,N_48729);
nor UO_2166 (O_2166,N_48913,N_49719);
nor UO_2167 (O_2167,N_49999,N_48249);
nor UO_2168 (O_2168,N_48124,N_48209);
xor UO_2169 (O_2169,N_48627,N_48111);
nor UO_2170 (O_2170,N_48122,N_48080);
nor UO_2171 (O_2171,N_49785,N_49071);
xor UO_2172 (O_2172,N_48726,N_49207);
nor UO_2173 (O_2173,N_48365,N_49338);
nor UO_2174 (O_2174,N_49720,N_48024);
nor UO_2175 (O_2175,N_49868,N_49270);
and UO_2176 (O_2176,N_49905,N_48038);
nand UO_2177 (O_2177,N_48322,N_48851);
or UO_2178 (O_2178,N_48741,N_49721);
nor UO_2179 (O_2179,N_48347,N_48763);
xnor UO_2180 (O_2180,N_48871,N_48362);
xnor UO_2181 (O_2181,N_48087,N_49629);
nand UO_2182 (O_2182,N_48540,N_48539);
nand UO_2183 (O_2183,N_48020,N_49080);
or UO_2184 (O_2184,N_49140,N_49235);
and UO_2185 (O_2185,N_49727,N_48346);
xnor UO_2186 (O_2186,N_49699,N_48411);
xnor UO_2187 (O_2187,N_49619,N_48407);
and UO_2188 (O_2188,N_48527,N_48517);
nand UO_2189 (O_2189,N_49594,N_48950);
xor UO_2190 (O_2190,N_48756,N_49416);
nand UO_2191 (O_2191,N_48679,N_49201);
xor UO_2192 (O_2192,N_49189,N_48856);
nand UO_2193 (O_2193,N_48364,N_49419);
or UO_2194 (O_2194,N_48870,N_49444);
and UO_2195 (O_2195,N_49477,N_48999);
nand UO_2196 (O_2196,N_49283,N_48279);
or UO_2197 (O_2197,N_48209,N_48621);
nand UO_2198 (O_2198,N_49417,N_49654);
nand UO_2199 (O_2199,N_49257,N_48588);
nor UO_2200 (O_2200,N_49957,N_49361);
and UO_2201 (O_2201,N_49173,N_48881);
nor UO_2202 (O_2202,N_48179,N_48668);
and UO_2203 (O_2203,N_48466,N_48609);
nor UO_2204 (O_2204,N_49606,N_49844);
xnor UO_2205 (O_2205,N_48761,N_49396);
or UO_2206 (O_2206,N_48142,N_48404);
xor UO_2207 (O_2207,N_49442,N_49684);
nor UO_2208 (O_2208,N_49703,N_49164);
nand UO_2209 (O_2209,N_49313,N_48672);
and UO_2210 (O_2210,N_49413,N_49679);
nand UO_2211 (O_2211,N_48174,N_49923);
or UO_2212 (O_2212,N_48772,N_48558);
and UO_2213 (O_2213,N_49412,N_49657);
nor UO_2214 (O_2214,N_48750,N_49459);
and UO_2215 (O_2215,N_48546,N_48165);
xor UO_2216 (O_2216,N_48574,N_49846);
nor UO_2217 (O_2217,N_49968,N_48988);
xor UO_2218 (O_2218,N_49899,N_48454);
nor UO_2219 (O_2219,N_48521,N_49597);
nand UO_2220 (O_2220,N_48646,N_49513);
or UO_2221 (O_2221,N_49712,N_48649);
nor UO_2222 (O_2222,N_49163,N_48360);
xnor UO_2223 (O_2223,N_48926,N_49722);
xnor UO_2224 (O_2224,N_48208,N_49140);
and UO_2225 (O_2225,N_49643,N_48161);
nand UO_2226 (O_2226,N_48029,N_48597);
nand UO_2227 (O_2227,N_49990,N_48695);
nor UO_2228 (O_2228,N_48470,N_49643);
nand UO_2229 (O_2229,N_48862,N_49633);
xor UO_2230 (O_2230,N_48882,N_49539);
nor UO_2231 (O_2231,N_48579,N_49971);
or UO_2232 (O_2232,N_48987,N_48624);
xnor UO_2233 (O_2233,N_48803,N_49122);
nand UO_2234 (O_2234,N_49420,N_48819);
xnor UO_2235 (O_2235,N_48666,N_49449);
nor UO_2236 (O_2236,N_48037,N_48262);
nand UO_2237 (O_2237,N_49687,N_48676);
nand UO_2238 (O_2238,N_49587,N_49418);
or UO_2239 (O_2239,N_49497,N_48736);
xor UO_2240 (O_2240,N_49263,N_49069);
xor UO_2241 (O_2241,N_49046,N_49079);
and UO_2242 (O_2242,N_48058,N_48407);
xor UO_2243 (O_2243,N_48437,N_48246);
or UO_2244 (O_2244,N_48776,N_49946);
xnor UO_2245 (O_2245,N_48094,N_48875);
xnor UO_2246 (O_2246,N_48318,N_48379);
and UO_2247 (O_2247,N_48342,N_48999);
and UO_2248 (O_2248,N_48834,N_49172);
xor UO_2249 (O_2249,N_48006,N_49541);
nand UO_2250 (O_2250,N_48393,N_49004);
and UO_2251 (O_2251,N_49812,N_48508);
or UO_2252 (O_2252,N_48895,N_49112);
nand UO_2253 (O_2253,N_49400,N_48464);
nor UO_2254 (O_2254,N_48899,N_48883);
nand UO_2255 (O_2255,N_48709,N_48311);
xor UO_2256 (O_2256,N_49042,N_48507);
xor UO_2257 (O_2257,N_48189,N_48691);
or UO_2258 (O_2258,N_49353,N_49207);
nor UO_2259 (O_2259,N_48039,N_49154);
or UO_2260 (O_2260,N_49549,N_49641);
and UO_2261 (O_2261,N_48833,N_48305);
nand UO_2262 (O_2262,N_49470,N_49887);
and UO_2263 (O_2263,N_48913,N_48508);
nand UO_2264 (O_2264,N_48603,N_49433);
and UO_2265 (O_2265,N_49823,N_48744);
and UO_2266 (O_2266,N_49512,N_48107);
xor UO_2267 (O_2267,N_49581,N_49670);
nand UO_2268 (O_2268,N_49803,N_49881);
xnor UO_2269 (O_2269,N_48309,N_48769);
nor UO_2270 (O_2270,N_49532,N_48516);
xnor UO_2271 (O_2271,N_49346,N_48166);
xnor UO_2272 (O_2272,N_49190,N_48785);
nor UO_2273 (O_2273,N_48467,N_48220);
or UO_2274 (O_2274,N_48472,N_49740);
or UO_2275 (O_2275,N_49545,N_48430);
xor UO_2276 (O_2276,N_49769,N_49150);
nor UO_2277 (O_2277,N_48977,N_48756);
nand UO_2278 (O_2278,N_48203,N_48680);
nand UO_2279 (O_2279,N_48122,N_49485);
nor UO_2280 (O_2280,N_48752,N_48556);
nand UO_2281 (O_2281,N_49831,N_48109);
nor UO_2282 (O_2282,N_48350,N_49635);
and UO_2283 (O_2283,N_48805,N_49011);
or UO_2284 (O_2284,N_48870,N_49731);
xnor UO_2285 (O_2285,N_49636,N_48109);
and UO_2286 (O_2286,N_49864,N_49968);
and UO_2287 (O_2287,N_49276,N_48346);
nand UO_2288 (O_2288,N_49963,N_48988);
nand UO_2289 (O_2289,N_48183,N_48566);
nor UO_2290 (O_2290,N_49432,N_48221);
and UO_2291 (O_2291,N_49227,N_48321);
nand UO_2292 (O_2292,N_48851,N_48661);
or UO_2293 (O_2293,N_48927,N_49617);
xnor UO_2294 (O_2294,N_49964,N_48097);
and UO_2295 (O_2295,N_48884,N_48508);
nor UO_2296 (O_2296,N_48327,N_48217);
or UO_2297 (O_2297,N_48577,N_48764);
xnor UO_2298 (O_2298,N_49666,N_49962);
or UO_2299 (O_2299,N_48977,N_49651);
nand UO_2300 (O_2300,N_49331,N_48969);
xor UO_2301 (O_2301,N_49966,N_49887);
or UO_2302 (O_2302,N_49718,N_48196);
or UO_2303 (O_2303,N_48428,N_49042);
or UO_2304 (O_2304,N_49215,N_49019);
or UO_2305 (O_2305,N_49496,N_48246);
or UO_2306 (O_2306,N_49470,N_49721);
nor UO_2307 (O_2307,N_48454,N_48230);
nor UO_2308 (O_2308,N_48812,N_49098);
xor UO_2309 (O_2309,N_49758,N_48098);
nand UO_2310 (O_2310,N_49796,N_48968);
nor UO_2311 (O_2311,N_48783,N_49166);
nand UO_2312 (O_2312,N_48483,N_49848);
and UO_2313 (O_2313,N_49261,N_49326);
and UO_2314 (O_2314,N_48145,N_49647);
xnor UO_2315 (O_2315,N_48213,N_49313);
nor UO_2316 (O_2316,N_49361,N_48200);
nand UO_2317 (O_2317,N_48771,N_48571);
or UO_2318 (O_2318,N_49797,N_48292);
or UO_2319 (O_2319,N_49138,N_48739);
xnor UO_2320 (O_2320,N_49774,N_48518);
nand UO_2321 (O_2321,N_49055,N_48300);
or UO_2322 (O_2322,N_48826,N_49389);
or UO_2323 (O_2323,N_48456,N_48965);
or UO_2324 (O_2324,N_49717,N_48912);
nand UO_2325 (O_2325,N_48183,N_48122);
nor UO_2326 (O_2326,N_49765,N_49497);
or UO_2327 (O_2327,N_48212,N_49468);
and UO_2328 (O_2328,N_48867,N_48290);
nand UO_2329 (O_2329,N_48956,N_49155);
nor UO_2330 (O_2330,N_49057,N_48873);
or UO_2331 (O_2331,N_48155,N_48594);
or UO_2332 (O_2332,N_48382,N_48064);
xnor UO_2333 (O_2333,N_48755,N_48587);
xor UO_2334 (O_2334,N_49715,N_48152);
or UO_2335 (O_2335,N_48690,N_48225);
xor UO_2336 (O_2336,N_49284,N_48202);
nor UO_2337 (O_2337,N_48762,N_48320);
xnor UO_2338 (O_2338,N_48513,N_49927);
xnor UO_2339 (O_2339,N_49940,N_48632);
nand UO_2340 (O_2340,N_48121,N_49030);
nand UO_2341 (O_2341,N_49029,N_49805);
nand UO_2342 (O_2342,N_49902,N_48341);
or UO_2343 (O_2343,N_49280,N_49889);
nor UO_2344 (O_2344,N_48783,N_48924);
nand UO_2345 (O_2345,N_48233,N_49561);
nand UO_2346 (O_2346,N_48063,N_48890);
and UO_2347 (O_2347,N_49198,N_48211);
and UO_2348 (O_2348,N_49045,N_49596);
and UO_2349 (O_2349,N_49179,N_49221);
and UO_2350 (O_2350,N_48222,N_48951);
nor UO_2351 (O_2351,N_48070,N_48902);
xnor UO_2352 (O_2352,N_48430,N_48370);
nand UO_2353 (O_2353,N_48319,N_49218);
and UO_2354 (O_2354,N_49656,N_49758);
nor UO_2355 (O_2355,N_48876,N_49764);
xnor UO_2356 (O_2356,N_49568,N_48863);
nor UO_2357 (O_2357,N_49021,N_48734);
and UO_2358 (O_2358,N_49964,N_49662);
or UO_2359 (O_2359,N_49983,N_49205);
nor UO_2360 (O_2360,N_49526,N_48119);
nor UO_2361 (O_2361,N_49543,N_49089);
and UO_2362 (O_2362,N_49604,N_49938);
or UO_2363 (O_2363,N_48647,N_49273);
nand UO_2364 (O_2364,N_49570,N_48743);
nor UO_2365 (O_2365,N_49797,N_49146);
or UO_2366 (O_2366,N_48127,N_48018);
xor UO_2367 (O_2367,N_48579,N_49589);
xnor UO_2368 (O_2368,N_48714,N_49387);
nor UO_2369 (O_2369,N_49781,N_48165);
xnor UO_2370 (O_2370,N_49303,N_49462);
nand UO_2371 (O_2371,N_48720,N_49797);
nor UO_2372 (O_2372,N_49518,N_49520);
nor UO_2373 (O_2373,N_48741,N_48990);
nand UO_2374 (O_2374,N_48484,N_48615);
nor UO_2375 (O_2375,N_48139,N_49686);
or UO_2376 (O_2376,N_48450,N_49602);
nor UO_2377 (O_2377,N_48810,N_48283);
nand UO_2378 (O_2378,N_48826,N_48804);
or UO_2379 (O_2379,N_49690,N_49338);
or UO_2380 (O_2380,N_48364,N_49763);
nor UO_2381 (O_2381,N_49883,N_49606);
nor UO_2382 (O_2382,N_49378,N_49439);
nor UO_2383 (O_2383,N_49970,N_48587);
and UO_2384 (O_2384,N_49331,N_48878);
and UO_2385 (O_2385,N_48838,N_49741);
nor UO_2386 (O_2386,N_49111,N_48452);
nand UO_2387 (O_2387,N_49965,N_48042);
nand UO_2388 (O_2388,N_48972,N_48782);
nand UO_2389 (O_2389,N_49631,N_49950);
or UO_2390 (O_2390,N_49790,N_48613);
nand UO_2391 (O_2391,N_48914,N_48813);
or UO_2392 (O_2392,N_49610,N_48403);
nand UO_2393 (O_2393,N_49835,N_49431);
and UO_2394 (O_2394,N_49830,N_49153);
and UO_2395 (O_2395,N_49092,N_48644);
or UO_2396 (O_2396,N_49540,N_48778);
xor UO_2397 (O_2397,N_48441,N_49116);
nand UO_2398 (O_2398,N_49514,N_48856);
xnor UO_2399 (O_2399,N_48264,N_49116);
or UO_2400 (O_2400,N_49506,N_49776);
xnor UO_2401 (O_2401,N_48014,N_48021);
xor UO_2402 (O_2402,N_48350,N_49356);
xor UO_2403 (O_2403,N_48344,N_49132);
nand UO_2404 (O_2404,N_48627,N_48730);
nand UO_2405 (O_2405,N_49685,N_48091);
xnor UO_2406 (O_2406,N_49835,N_49573);
and UO_2407 (O_2407,N_48303,N_48728);
and UO_2408 (O_2408,N_48372,N_49952);
nand UO_2409 (O_2409,N_49811,N_49410);
and UO_2410 (O_2410,N_48799,N_48150);
or UO_2411 (O_2411,N_49682,N_48313);
nand UO_2412 (O_2412,N_49639,N_48580);
xor UO_2413 (O_2413,N_48778,N_49869);
and UO_2414 (O_2414,N_49647,N_48319);
xor UO_2415 (O_2415,N_48763,N_48198);
nor UO_2416 (O_2416,N_48645,N_48079);
and UO_2417 (O_2417,N_48005,N_48627);
xnor UO_2418 (O_2418,N_48929,N_48218);
or UO_2419 (O_2419,N_49745,N_48689);
xnor UO_2420 (O_2420,N_49566,N_49180);
or UO_2421 (O_2421,N_49325,N_48645);
nand UO_2422 (O_2422,N_49562,N_48814);
or UO_2423 (O_2423,N_49489,N_48725);
and UO_2424 (O_2424,N_48595,N_48178);
nand UO_2425 (O_2425,N_49993,N_48774);
or UO_2426 (O_2426,N_49667,N_49991);
nand UO_2427 (O_2427,N_48346,N_49134);
nor UO_2428 (O_2428,N_49579,N_48696);
xnor UO_2429 (O_2429,N_49330,N_49150);
and UO_2430 (O_2430,N_49111,N_48977);
or UO_2431 (O_2431,N_49539,N_49797);
xnor UO_2432 (O_2432,N_48945,N_48112);
or UO_2433 (O_2433,N_49104,N_49778);
and UO_2434 (O_2434,N_48094,N_49887);
xor UO_2435 (O_2435,N_49999,N_49949);
nor UO_2436 (O_2436,N_49461,N_49013);
nor UO_2437 (O_2437,N_48273,N_48264);
nand UO_2438 (O_2438,N_48469,N_49342);
nor UO_2439 (O_2439,N_49816,N_49958);
or UO_2440 (O_2440,N_48325,N_48335);
nand UO_2441 (O_2441,N_49525,N_48105);
xor UO_2442 (O_2442,N_49233,N_48568);
xnor UO_2443 (O_2443,N_49101,N_49622);
xnor UO_2444 (O_2444,N_48818,N_49397);
xnor UO_2445 (O_2445,N_49206,N_49840);
and UO_2446 (O_2446,N_48147,N_49858);
nand UO_2447 (O_2447,N_48025,N_49181);
and UO_2448 (O_2448,N_49304,N_48176);
and UO_2449 (O_2449,N_48661,N_48924);
nor UO_2450 (O_2450,N_49734,N_49053);
nand UO_2451 (O_2451,N_48325,N_48813);
or UO_2452 (O_2452,N_49905,N_49439);
and UO_2453 (O_2453,N_48552,N_49888);
and UO_2454 (O_2454,N_49314,N_48307);
xor UO_2455 (O_2455,N_48742,N_49512);
and UO_2456 (O_2456,N_48353,N_48847);
or UO_2457 (O_2457,N_49642,N_49604);
nor UO_2458 (O_2458,N_48967,N_48474);
or UO_2459 (O_2459,N_48256,N_49011);
nand UO_2460 (O_2460,N_49558,N_49307);
nor UO_2461 (O_2461,N_48133,N_49602);
nand UO_2462 (O_2462,N_49836,N_49186);
or UO_2463 (O_2463,N_49932,N_49103);
nand UO_2464 (O_2464,N_48526,N_48140);
or UO_2465 (O_2465,N_49834,N_48962);
nor UO_2466 (O_2466,N_49660,N_48537);
and UO_2467 (O_2467,N_49876,N_49862);
xnor UO_2468 (O_2468,N_49697,N_48076);
and UO_2469 (O_2469,N_48001,N_48787);
nand UO_2470 (O_2470,N_48671,N_48041);
or UO_2471 (O_2471,N_48340,N_48173);
nand UO_2472 (O_2472,N_48794,N_49978);
or UO_2473 (O_2473,N_48818,N_48664);
nand UO_2474 (O_2474,N_49784,N_48035);
and UO_2475 (O_2475,N_48076,N_49417);
nor UO_2476 (O_2476,N_49290,N_49612);
xor UO_2477 (O_2477,N_49889,N_49184);
or UO_2478 (O_2478,N_49341,N_48539);
xor UO_2479 (O_2479,N_48683,N_48704);
nor UO_2480 (O_2480,N_49223,N_48169);
or UO_2481 (O_2481,N_48848,N_48978);
nor UO_2482 (O_2482,N_49647,N_48693);
xor UO_2483 (O_2483,N_48970,N_48210);
or UO_2484 (O_2484,N_48774,N_48457);
nand UO_2485 (O_2485,N_48855,N_49741);
or UO_2486 (O_2486,N_48088,N_49446);
nor UO_2487 (O_2487,N_49268,N_48255);
and UO_2488 (O_2488,N_48930,N_49793);
and UO_2489 (O_2489,N_49541,N_49770);
or UO_2490 (O_2490,N_48661,N_49037);
xor UO_2491 (O_2491,N_48473,N_48474);
or UO_2492 (O_2492,N_48782,N_48422);
xor UO_2493 (O_2493,N_48477,N_49744);
and UO_2494 (O_2494,N_48084,N_49845);
and UO_2495 (O_2495,N_48760,N_48261);
or UO_2496 (O_2496,N_49033,N_48111);
nand UO_2497 (O_2497,N_48747,N_49313);
nand UO_2498 (O_2498,N_49934,N_48641);
nor UO_2499 (O_2499,N_48718,N_49662);
and UO_2500 (O_2500,N_49145,N_48474);
nor UO_2501 (O_2501,N_49343,N_49259);
nor UO_2502 (O_2502,N_48417,N_48749);
and UO_2503 (O_2503,N_48791,N_48067);
nand UO_2504 (O_2504,N_49400,N_49765);
nand UO_2505 (O_2505,N_49920,N_48194);
and UO_2506 (O_2506,N_48247,N_49419);
and UO_2507 (O_2507,N_48634,N_48278);
or UO_2508 (O_2508,N_48124,N_48199);
xor UO_2509 (O_2509,N_49548,N_49058);
nand UO_2510 (O_2510,N_49938,N_49137);
nand UO_2511 (O_2511,N_49737,N_48584);
nand UO_2512 (O_2512,N_48824,N_48707);
nor UO_2513 (O_2513,N_49638,N_48129);
nand UO_2514 (O_2514,N_49574,N_49259);
xnor UO_2515 (O_2515,N_49343,N_48116);
and UO_2516 (O_2516,N_48964,N_49062);
nand UO_2517 (O_2517,N_48598,N_48642);
and UO_2518 (O_2518,N_49019,N_49010);
nand UO_2519 (O_2519,N_48278,N_48783);
xor UO_2520 (O_2520,N_49706,N_49249);
nor UO_2521 (O_2521,N_48861,N_48078);
xnor UO_2522 (O_2522,N_49345,N_49339);
or UO_2523 (O_2523,N_48977,N_49311);
xnor UO_2524 (O_2524,N_49486,N_48437);
nand UO_2525 (O_2525,N_49809,N_48500);
nor UO_2526 (O_2526,N_49835,N_49994);
and UO_2527 (O_2527,N_49618,N_49243);
and UO_2528 (O_2528,N_49864,N_49088);
nand UO_2529 (O_2529,N_49439,N_49194);
or UO_2530 (O_2530,N_48032,N_49448);
xor UO_2531 (O_2531,N_48723,N_48397);
nand UO_2532 (O_2532,N_48778,N_49747);
and UO_2533 (O_2533,N_48225,N_49252);
or UO_2534 (O_2534,N_48273,N_49990);
xor UO_2535 (O_2535,N_49667,N_49678);
and UO_2536 (O_2536,N_49859,N_48656);
or UO_2537 (O_2537,N_49625,N_48540);
and UO_2538 (O_2538,N_49284,N_49167);
nand UO_2539 (O_2539,N_49502,N_48573);
xnor UO_2540 (O_2540,N_49166,N_49290);
nand UO_2541 (O_2541,N_49792,N_49352);
nand UO_2542 (O_2542,N_48996,N_49287);
and UO_2543 (O_2543,N_49523,N_49426);
nand UO_2544 (O_2544,N_49570,N_48408);
nand UO_2545 (O_2545,N_49359,N_49445);
and UO_2546 (O_2546,N_48477,N_48313);
nor UO_2547 (O_2547,N_49658,N_48212);
and UO_2548 (O_2548,N_48156,N_48328);
nand UO_2549 (O_2549,N_48284,N_49471);
nand UO_2550 (O_2550,N_48588,N_49543);
and UO_2551 (O_2551,N_48954,N_49367);
xnor UO_2552 (O_2552,N_48315,N_49629);
and UO_2553 (O_2553,N_48910,N_49192);
or UO_2554 (O_2554,N_49209,N_48674);
nand UO_2555 (O_2555,N_48645,N_49591);
or UO_2556 (O_2556,N_49361,N_49099);
nand UO_2557 (O_2557,N_49182,N_48808);
xor UO_2558 (O_2558,N_48818,N_49791);
nor UO_2559 (O_2559,N_48767,N_48473);
and UO_2560 (O_2560,N_48659,N_48027);
xnor UO_2561 (O_2561,N_49852,N_49400);
nand UO_2562 (O_2562,N_49493,N_48713);
or UO_2563 (O_2563,N_48111,N_48320);
or UO_2564 (O_2564,N_49292,N_48141);
and UO_2565 (O_2565,N_48987,N_49244);
xor UO_2566 (O_2566,N_48399,N_48093);
nand UO_2567 (O_2567,N_49522,N_48999);
and UO_2568 (O_2568,N_48143,N_49630);
nand UO_2569 (O_2569,N_49262,N_49907);
or UO_2570 (O_2570,N_49373,N_48551);
nand UO_2571 (O_2571,N_49121,N_49599);
or UO_2572 (O_2572,N_49122,N_49072);
nand UO_2573 (O_2573,N_48174,N_48717);
or UO_2574 (O_2574,N_49491,N_48785);
xor UO_2575 (O_2575,N_49096,N_49650);
or UO_2576 (O_2576,N_48222,N_49129);
or UO_2577 (O_2577,N_48712,N_49894);
xor UO_2578 (O_2578,N_49248,N_49630);
and UO_2579 (O_2579,N_48474,N_49945);
nor UO_2580 (O_2580,N_49759,N_48748);
nand UO_2581 (O_2581,N_48979,N_48754);
nand UO_2582 (O_2582,N_49671,N_49929);
nor UO_2583 (O_2583,N_49103,N_49389);
and UO_2584 (O_2584,N_48164,N_49848);
and UO_2585 (O_2585,N_48484,N_48752);
and UO_2586 (O_2586,N_49147,N_48030);
or UO_2587 (O_2587,N_48221,N_49375);
nor UO_2588 (O_2588,N_49869,N_48361);
and UO_2589 (O_2589,N_48287,N_49216);
xnor UO_2590 (O_2590,N_49618,N_48571);
nand UO_2591 (O_2591,N_49042,N_49352);
or UO_2592 (O_2592,N_49333,N_48551);
nor UO_2593 (O_2593,N_48361,N_49973);
nor UO_2594 (O_2594,N_48884,N_49567);
nand UO_2595 (O_2595,N_49240,N_48630);
and UO_2596 (O_2596,N_49226,N_49144);
or UO_2597 (O_2597,N_48823,N_48592);
and UO_2598 (O_2598,N_49738,N_49295);
and UO_2599 (O_2599,N_49121,N_49630);
xnor UO_2600 (O_2600,N_49052,N_48929);
xor UO_2601 (O_2601,N_48032,N_49519);
xor UO_2602 (O_2602,N_49494,N_49773);
and UO_2603 (O_2603,N_49858,N_49896);
nor UO_2604 (O_2604,N_49715,N_48586);
nand UO_2605 (O_2605,N_49134,N_49694);
xor UO_2606 (O_2606,N_48041,N_48317);
xor UO_2607 (O_2607,N_48171,N_48841);
nand UO_2608 (O_2608,N_48123,N_48805);
nand UO_2609 (O_2609,N_49530,N_48207);
xor UO_2610 (O_2610,N_49748,N_49632);
and UO_2611 (O_2611,N_49961,N_49088);
nand UO_2612 (O_2612,N_49872,N_49364);
nor UO_2613 (O_2613,N_49252,N_49469);
xnor UO_2614 (O_2614,N_48396,N_48763);
nand UO_2615 (O_2615,N_49979,N_48056);
or UO_2616 (O_2616,N_49432,N_48538);
nand UO_2617 (O_2617,N_49069,N_48221);
nor UO_2618 (O_2618,N_49716,N_49840);
and UO_2619 (O_2619,N_48265,N_48866);
and UO_2620 (O_2620,N_48574,N_49412);
nor UO_2621 (O_2621,N_49838,N_48682);
or UO_2622 (O_2622,N_49862,N_49010);
xor UO_2623 (O_2623,N_48213,N_48086);
and UO_2624 (O_2624,N_48171,N_48384);
nand UO_2625 (O_2625,N_49427,N_48386);
and UO_2626 (O_2626,N_48591,N_48309);
nand UO_2627 (O_2627,N_49442,N_49765);
and UO_2628 (O_2628,N_48606,N_49793);
nand UO_2629 (O_2629,N_49830,N_49301);
and UO_2630 (O_2630,N_49546,N_48831);
xnor UO_2631 (O_2631,N_48669,N_49274);
xor UO_2632 (O_2632,N_48408,N_48664);
nor UO_2633 (O_2633,N_48237,N_49749);
xnor UO_2634 (O_2634,N_48730,N_48227);
nand UO_2635 (O_2635,N_49612,N_48102);
xnor UO_2636 (O_2636,N_49980,N_48289);
and UO_2637 (O_2637,N_48864,N_48550);
or UO_2638 (O_2638,N_48528,N_48726);
nand UO_2639 (O_2639,N_49554,N_48398);
and UO_2640 (O_2640,N_48678,N_48519);
xor UO_2641 (O_2641,N_48717,N_49413);
and UO_2642 (O_2642,N_49932,N_49274);
nor UO_2643 (O_2643,N_49253,N_49374);
and UO_2644 (O_2644,N_49849,N_49890);
xor UO_2645 (O_2645,N_48757,N_48716);
nand UO_2646 (O_2646,N_49641,N_49582);
nor UO_2647 (O_2647,N_48909,N_49370);
nand UO_2648 (O_2648,N_48814,N_48029);
or UO_2649 (O_2649,N_49515,N_49498);
nand UO_2650 (O_2650,N_49902,N_48123);
or UO_2651 (O_2651,N_48519,N_48211);
or UO_2652 (O_2652,N_48655,N_48842);
or UO_2653 (O_2653,N_48507,N_49432);
nand UO_2654 (O_2654,N_48596,N_48846);
and UO_2655 (O_2655,N_49393,N_49812);
and UO_2656 (O_2656,N_48991,N_48838);
nand UO_2657 (O_2657,N_48892,N_48307);
nor UO_2658 (O_2658,N_48132,N_49990);
nand UO_2659 (O_2659,N_48881,N_48902);
nor UO_2660 (O_2660,N_49130,N_49597);
nor UO_2661 (O_2661,N_48546,N_49205);
nor UO_2662 (O_2662,N_48590,N_49928);
and UO_2663 (O_2663,N_48701,N_48905);
nand UO_2664 (O_2664,N_49289,N_49152);
and UO_2665 (O_2665,N_48263,N_49334);
xnor UO_2666 (O_2666,N_48925,N_48812);
nand UO_2667 (O_2667,N_48457,N_48814);
and UO_2668 (O_2668,N_49459,N_48495);
xnor UO_2669 (O_2669,N_48544,N_48304);
or UO_2670 (O_2670,N_48359,N_49575);
nor UO_2671 (O_2671,N_48359,N_48684);
or UO_2672 (O_2672,N_49163,N_48860);
xnor UO_2673 (O_2673,N_49489,N_48353);
nand UO_2674 (O_2674,N_48407,N_49256);
and UO_2675 (O_2675,N_49308,N_49729);
xor UO_2676 (O_2676,N_48463,N_48786);
nor UO_2677 (O_2677,N_49158,N_48995);
nor UO_2678 (O_2678,N_48737,N_49161);
xnor UO_2679 (O_2679,N_48744,N_49141);
or UO_2680 (O_2680,N_49651,N_49414);
or UO_2681 (O_2681,N_49312,N_49863);
xnor UO_2682 (O_2682,N_49426,N_48907);
xnor UO_2683 (O_2683,N_49243,N_49778);
and UO_2684 (O_2684,N_49792,N_48811);
xnor UO_2685 (O_2685,N_49646,N_48113);
and UO_2686 (O_2686,N_49513,N_49283);
xor UO_2687 (O_2687,N_49260,N_49958);
nand UO_2688 (O_2688,N_49272,N_48868);
xnor UO_2689 (O_2689,N_48815,N_48791);
xor UO_2690 (O_2690,N_48558,N_49445);
nand UO_2691 (O_2691,N_48072,N_49824);
nand UO_2692 (O_2692,N_49619,N_49566);
xnor UO_2693 (O_2693,N_49397,N_49087);
and UO_2694 (O_2694,N_49636,N_49215);
xor UO_2695 (O_2695,N_48654,N_49312);
nand UO_2696 (O_2696,N_48375,N_49848);
nor UO_2697 (O_2697,N_48348,N_49365);
or UO_2698 (O_2698,N_49680,N_49948);
or UO_2699 (O_2699,N_48502,N_49726);
or UO_2700 (O_2700,N_48217,N_48126);
nand UO_2701 (O_2701,N_49323,N_49309);
nor UO_2702 (O_2702,N_49292,N_49589);
and UO_2703 (O_2703,N_49956,N_48729);
and UO_2704 (O_2704,N_48924,N_49434);
xnor UO_2705 (O_2705,N_49938,N_48093);
or UO_2706 (O_2706,N_49038,N_48951);
nor UO_2707 (O_2707,N_49255,N_48497);
nor UO_2708 (O_2708,N_49869,N_49322);
or UO_2709 (O_2709,N_49683,N_48821);
and UO_2710 (O_2710,N_49711,N_49255);
and UO_2711 (O_2711,N_48967,N_48510);
nor UO_2712 (O_2712,N_48018,N_48757);
nor UO_2713 (O_2713,N_49835,N_49771);
and UO_2714 (O_2714,N_49962,N_48357);
or UO_2715 (O_2715,N_48944,N_49536);
nand UO_2716 (O_2716,N_48934,N_48580);
nand UO_2717 (O_2717,N_48018,N_48382);
nor UO_2718 (O_2718,N_49221,N_48765);
nor UO_2719 (O_2719,N_49573,N_49671);
or UO_2720 (O_2720,N_49979,N_49474);
xnor UO_2721 (O_2721,N_49918,N_48119);
and UO_2722 (O_2722,N_48310,N_48316);
and UO_2723 (O_2723,N_49500,N_49252);
nor UO_2724 (O_2724,N_48952,N_48223);
or UO_2725 (O_2725,N_48773,N_49670);
nor UO_2726 (O_2726,N_49193,N_49371);
xnor UO_2727 (O_2727,N_48892,N_49763);
nor UO_2728 (O_2728,N_49853,N_49348);
nand UO_2729 (O_2729,N_48705,N_49760);
xor UO_2730 (O_2730,N_49601,N_48639);
and UO_2731 (O_2731,N_49262,N_49675);
nor UO_2732 (O_2732,N_48013,N_48698);
and UO_2733 (O_2733,N_48685,N_48047);
nor UO_2734 (O_2734,N_48895,N_48880);
xnor UO_2735 (O_2735,N_48929,N_48499);
and UO_2736 (O_2736,N_49982,N_48286);
xnor UO_2737 (O_2737,N_49987,N_48513);
nand UO_2738 (O_2738,N_48872,N_49953);
or UO_2739 (O_2739,N_49819,N_49375);
and UO_2740 (O_2740,N_48929,N_49550);
nor UO_2741 (O_2741,N_49306,N_48967);
and UO_2742 (O_2742,N_49592,N_49731);
and UO_2743 (O_2743,N_49715,N_49982);
nor UO_2744 (O_2744,N_49282,N_49616);
nand UO_2745 (O_2745,N_48189,N_49157);
nor UO_2746 (O_2746,N_48263,N_48631);
and UO_2747 (O_2747,N_48137,N_49174);
nand UO_2748 (O_2748,N_48491,N_48948);
or UO_2749 (O_2749,N_49290,N_49362);
nor UO_2750 (O_2750,N_48712,N_49264);
nand UO_2751 (O_2751,N_48254,N_48092);
xor UO_2752 (O_2752,N_48288,N_49563);
xnor UO_2753 (O_2753,N_49716,N_48634);
and UO_2754 (O_2754,N_49793,N_49523);
nand UO_2755 (O_2755,N_48977,N_48475);
nor UO_2756 (O_2756,N_49163,N_48961);
or UO_2757 (O_2757,N_49192,N_48402);
and UO_2758 (O_2758,N_48402,N_48027);
xnor UO_2759 (O_2759,N_48832,N_49096);
and UO_2760 (O_2760,N_49981,N_48064);
and UO_2761 (O_2761,N_48527,N_49754);
and UO_2762 (O_2762,N_49316,N_49264);
or UO_2763 (O_2763,N_48619,N_48067);
nand UO_2764 (O_2764,N_49668,N_49537);
xnor UO_2765 (O_2765,N_49680,N_48608);
nand UO_2766 (O_2766,N_49142,N_49218);
xnor UO_2767 (O_2767,N_49989,N_49707);
or UO_2768 (O_2768,N_49669,N_48442);
nand UO_2769 (O_2769,N_48226,N_49226);
xor UO_2770 (O_2770,N_49209,N_49940);
xor UO_2771 (O_2771,N_49943,N_48923);
or UO_2772 (O_2772,N_49631,N_48332);
xor UO_2773 (O_2773,N_48833,N_49168);
nand UO_2774 (O_2774,N_49992,N_49403);
or UO_2775 (O_2775,N_48709,N_48584);
or UO_2776 (O_2776,N_48293,N_48470);
nor UO_2777 (O_2777,N_48744,N_49545);
nor UO_2778 (O_2778,N_49533,N_49397);
xnor UO_2779 (O_2779,N_49366,N_49804);
and UO_2780 (O_2780,N_49711,N_48351);
nor UO_2781 (O_2781,N_49850,N_49058);
xor UO_2782 (O_2782,N_48524,N_48807);
and UO_2783 (O_2783,N_49197,N_49068);
or UO_2784 (O_2784,N_49469,N_49761);
or UO_2785 (O_2785,N_49490,N_48994);
xor UO_2786 (O_2786,N_49474,N_49341);
nor UO_2787 (O_2787,N_49401,N_48230);
or UO_2788 (O_2788,N_48235,N_48795);
nor UO_2789 (O_2789,N_48571,N_49591);
or UO_2790 (O_2790,N_49459,N_48413);
and UO_2791 (O_2791,N_48964,N_49103);
nand UO_2792 (O_2792,N_49053,N_49857);
and UO_2793 (O_2793,N_48288,N_49335);
or UO_2794 (O_2794,N_48897,N_48366);
or UO_2795 (O_2795,N_49204,N_49349);
nand UO_2796 (O_2796,N_49279,N_49253);
and UO_2797 (O_2797,N_49079,N_49350);
nand UO_2798 (O_2798,N_48613,N_48881);
nand UO_2799 (O_2799,N_49491,N_48323);
nor UO_2800 (O_2800,N_48710,N_49901);
nor UO_2801 (O_2801,N_49519,N_48550);
nand UO_2802 (O_2802,N_49095,N_48248);
or UO_2803 (O_2803,N_48627,N_48929);
nor UO_2804 (O_2804,N_49764,N_49876);
nand UO_2805 (O_2805,N_49973,N_49721);
or UO_2806 (O_2806,N_48267,N_49170);
nand UO_2807 (O_2807,N_48817,N_48949);
nor UO_2808 (O_2808,N_49332,N_48885);
and UO_2809 (O_2809,N_49945,N_48658);
xnor UO_2810 (O_2810,N_48412,N_48752);
nand UO_2811 (O_2811,N_49957,N_48951);
or UO_2812 (O_2812,N_49689,N_48613);
and UO_2813 (O_2813,N_49836,N_48115);
nor UO_2814 (O_2814,N_48001,N_49333);
or UO_2815 (O_2815,N_48106,N_49706);
and UO_2816 (O_2816,N_48423,N_49051);
nor UO_2817 (O_2817,N_49471,N_48137);
or UO_2818 (O_2818,N_49261,N_48950);
or UO_2819 (O_2819,N_48100,N_48544);
and UO_2820 (O_2820,N_48296,N_49628);
and UO_2821 (O_2821,N_48113,N_48797);
xnor UO_2822 (O_2822,N_48099,N_49002);
or UO_2823 (O_2823,N_49501,N_48994);
xnor UO_2824 (O_2824,N_49507,N_48930);
or UO_2825 (O_2825,N_49338,N_48779);
nand UO_2826 (O_2826,N_49733,N_48749);
xnor UO_2827 (O_2827,N_48460,N_49089);
or UO_2828 (O_2828,N_48408,N_49930);
or UO_2829 (O_2829,N_48328,N_48251);
and UO_2830 (O_2830,N_49675,N_49915);
nand UO_2831 (O_2831,N_48571,N_49127);
xor UO_2832 (O_2832,N_48273,N_48968);
or UO_2833 (O_2833,N_48147,N_48939);
nor UO_2834 (O_2834,N_48409,N_48187);
or UO_2835 (O_2835,N_48793,N_48380);
nor UO_2836 (O_2836,N_48613,N_49570);
xnor UO_2837 (O_2837,N_49964,N_49795);
and UO_2838 (O_2838,N_48702,N_48050);
xnor UO_2839 (O_2839,N_49935,N_48869);
xnor UO_2840 (O_2840,N_48485,N_48709);
or UO_2841 (O_2841,N_48895,N_49964);
and UO_2842 (O_2842,N_48527,N_48207);
or UO_2843 (O_2843,N_49064,N_48101);
or UO_2844 (O_2844,N_48565,N_48202);
and UO_2845 (O_2845,N_48227,N_48797);
nor UO_2846 (O_2846,N_49248,N_48287);
and UO_2847 (O_2847,N_48832,N_48491);
nand UO_2848 (O_2848,N_48417,N_49666);
and UO_2849 (O_2849,N_48059,N_48125);
nand UO_2850 (O_2850,N_48724,N_49440);
nand UO_2851 (O_2851,N_48763,N_48929);
and UO_2852 (O_2852,N_49481,N_49843);
xor UO_2853 (O_2853,N_48515,N_48138);
or UO_2854 (O_2854,N_49576,N_49524);
nor UO_2855 (O_2855,N_49791,N_49661);
and UO_2856 (O_2856,N_49285,N_48777);
xor UO_2857 (O_2857,N_48428,N_48934);
or UO_2858 (O_2858,N_48410,N_49300);
xor UO_2859 (O_2859,N_49711,N_48926);
nand UO_2860 (O_2860,N_48638,N_48813);
nand UO_2861 (O_2861,N_48721,N_48730);
xor UO_2862 (O_2862,N_48507,N_48289);
and UO_2863 (O_2863,N_49994,N_49580);
nand UO_2864 (O_2864,N_48515,N_48727);
or UO_2865 (O_2865,N_49497,N_49714);
nand UO_2866 (O_2866,N_48499,N_48655);
nand UO_2867 (O_2867,N_49835,N_48032);
xnor UO_2868 (O_2868,N_49930,N_49326);
xnor UO_2869 (O_2869,N_48534,N_49900);
nor UO_2870 (O_2870,N_48942,N_49208);
and UO_2871 (O_2871,N_48840,N_48720);
and UO_2872 (O_2872,N_49852,N_48684);
nand UO_2873 (O_2873,N_49319,N_49017);
nand UO_2874 (O_2874,N_48287,N_49141);
and UO_2875 (O_2875,N_49642,N_49211);
nor UO_2876 (O_2876,N_48599,N_49943);
nand UO_2877 (O_2877,N_49950,N_48073);
or UO_2878 (O_2878,N_48063,N_48638);
and UO_2879 (O_2879,N_48602,N_48423);
nor UO_2880 (O_2880,N_49415,N_48430);
nand UO_2881 (O_2881,N_48982,N_49488);
and UO_2882 (O_2882,N_48912,N_48824);
nor UO_2883 (O_2883,N_49589,N_49529);
nand UO_2884 (O_2884,N_49195,N_48889);
nand UO_2885 (O_2885,N_49530,N_48717);
or UO_2886 (O_2886,N_49029,N_49906);
nand UO_2887 (O_2887,N_49062,N_49246);
nor UO_2888 (O_2888,N_48452,N_48623);
and UO_2889 (O_2889,N_49688,N_49367);
nor UO_2890 (O_2890,N_48900,N_49911);
nand UO_2891 (O_2891,N_49623,N_48475);
or UO_2892 (O_2892,N_49688,N_48303);
nand UO_2893 (O_2893,N_48937,N_48025);
or UO_2894 (O_2894,N_48757,N_49332);
or UO_2895 (O_2895,N_48902,N_49893);
or UO_2896 (O_2896,N_48489,N_49386);
or UO_2897 (O_2897,N_48430,N_49630);
or UO_2898 (O_2898,N_49904,N_49250);
nand UO_2899 (O_2899,N_48632,N_49157);
and UO_2900 (O_2900,N_49060,N_48735);
nor UO_2901 (O_2901,N_49624,N_49447);
nor UO_2902 (O_2902,N_48433,N_49964);
or UO_2903 (O_2903,N_48669,N_49067);
and UO_2904 (O_2904,N_48555,N_48802);
and UO_2905 (O_2905,N_48357,N_48555);
xor UO_2906 (O_2906,N_49960,N_49395);
nand UO_2907 (O_2907,N_48890,N_48381);
nand UO_2908 (O_2908,N_48977,N_48825);
or UO_2909 (O_2909,N_48155,N_48238);
and UO_2910 (O_2910,N_49327,N_48049);
nor UO_2911 (O_2911,N_49475,N_48795);
xnor UO_2912 (O_2912,N_48811,N_48261);
or UO_2913 (O_2913,N_48400,N_49718);
nand UO_2914 (O_2914,N_48204,N_49004);
xor UO_2915 (O_2915,N_49471,N_49322);
or UO_2916 (O_2916,N_49688,N_49053);
nand UO_2917 (O_2917,N_48167,N_48159);
or UO_2918 (O_2918,N_48159,N_49971);
xor UO_2919 (O_2919,N_49195,N_49812);
nor UO_2920 (O_2920,N_49233,N_49053);
or UO_2921 (O_2921,N_48138,N_48687);
or UO_2922 (O_2922,N_49321,N_49501);
and UO_2923 (O_2923,N_48330,N_49287);
nor UO_2924 (O_2924,N_49235,N_49042);
xnor UO_2925 (O_2925,N_49181,N_48547);
or UO_2926 (O_2926,N_48763,N_49939);
nand UO_2927 (O_2927,N_48160,N_49238);
and UO_2928 (O_2928,N_49944,N_48973);
or UO_2929 (O_2929,N_48903,N_48710);
xor UO_2930 (O_2930,N_49508,N_49094);
nor UO_2931 (O_2931,N_49217,N_48930);
nor UO_2932 (O_2932,N_48090,N_49732);
nor UO_2933 (O_2933,N_49320,N_48585);
nand UO_2934 (O_2934,N_49518,N_48904);
and UO_2935 (O_2935,N_49560,N_48377);
or UO_2936 (O_2936,N_48812,N_49382);
and UO_2937 (O_2937,N_49981,N_48726);
and UO_2938 (O_2938,N_48268,N_49098);
or UO_2939 (O_2939,N_49874,N_49157);
and UO_2940 (O_2940,N_49925,N_48199);
nor UO_2941 (O_2941,N_49079,N_48440);
nand UO_2942 (O_2942,N_48595,N_49915);
or UO_2943 (O_2943,N_49237,N_48797);
and UO_2944 (O_2944,N_49309,N_48157);
and UO_2945 (O_2945,N_48624,N_48709);
nor UO_2946 (O_2946,N_49331,N_49629);
and UO_2947 (O_2947,N_49376,N_48880);
or UO_2948 (O_2948,N_48569,N_49945);
or UO_2949 (O_2949,N_49172,N_49188);
xor UO_2950 (O_2950,N_49312,N_48757);
xor UO_2951 (O_2951,N_48474,N_49328);
and UO_2952 (O_2952,N_49573,N_49518);
nand UO_2953 (O_2953,N_49168,N_49081);
or UO_2954 (O_2954,N_48864,N_48478);
or UO_2955 (O_2955,N_48761,N_48363);
xnor UO_2956 (O_2956,N_48376,N_49360);
nor UO_2957 (O_2957,N_48421,N_48700);
nand UO_2958 (O_2958,N_49860,N_48090);
nor UO_2959 (O_2959,N_49878,N_48252);
and UO_2960 (O_2960,N_48463,N_49536);
and UO_2961 (O_2961,N_48015,N_48656);
xnor UO_2962 (O_2962,N_49030,N_48511);
and UO_2963 (O_2963,N_48759,N_49071);
nor UO_2964 (O_2964,N_48455,N_48505);
nor UO_2965 (O_2965,N_49918,N_48893);
or UO_2966 (O_2966,N_49856,N_49550);
nand UO_2967 (O_2967,N_48307,N_48925);
xor UO_2968 (O_2968,N_49899,N_48950);
xor UO_2969 (O_2969,N_48930,N_49988);
or UO_2970 (O_2970,N_49753,N_49205);
nor UO_2971 (O_2971,N_49907,N_48851);
and UO_2972 (O_2972,N_49674,N_49101);
nor UO_2973 (O_2973,N_48401,N_49373);
xor UO_2974 (O_2974,N_49317,N_49030);
or UO_2975 (O_2975,N_48664,N_49126);
xnor UO_2976 (O_2976,N_49404,N_48470);
and UO_2977 (O_2977,N_49536,N_49304);
nand UO_2978 (O_2978,N_49520,N_49731);
or UO_2979 (O_2979,N_48670,N_48566);
nand UO_2980 (O_2980,N_49532,N_48750);
xnor UO_2981 (O_2981,N_49830,N_49471);
and UO_2982 (O_2982,N_49943,N_49836);
nor UO_2983 (O_2983,N_49273,N_49593);
xor UO_2984 (O_2984,N_48972,N_48074);
or UO_2985 (O_2985,N_48921,N_48507);
nor UO_2986 (O_2986,N_49875,N_49830);
nand UO_2987 (O_2987,N_49456,N_49797);
nor UO_2988 (O_2988,N_49876,N_49602);
nor UO_2989 (O_2989,N_48525,N_49305);
or UO_2990 (O_2990,N_49651,N_49582);
or UO_2991 (O_2991,N_48884,N_49586);
or UO_2992 (O_2992,N_48931,N_48738);
nand UO_2993 (O_2993,N_48293,N_48003);
or UO_2994 (O_2994,N_48873,N_49647);
nand UO_2995 (O_2995,N_48002,N_48059);
xor UO_2996 (O_2996,N_49066,N_48328);
nand UO_2997 (O_2997,N_49473,N_48797);
xnor UO_2998 (O_2998,N_48383,N_48892);
nand UO_2999 (O_2999,N_48094,N_49986);
and UO_3000 (O_3000,N_48028,N_48255);
nor UO_3001 (O_3001,N_49761,N_48434);
xnor UO_3002 (O_3002,N_48436,N_48880);
nand UO_3003 (O_3003,N_49125,N_48175);
nor UO_3004 (O_3004,N_48355,N_48502);
xor UO_3005 (O_3005,N_48593,N_48814);
nand UO_3006 (O_3006,N_48600,N_48317);
xor UO_3007 (O_3007,N_48443,N_48884);
or UO_3008 (O_3008,N_48553,N_49772);
nand UO_3009 (O_3009,N_49196,N_49248);
xor UO_3010 (O_3010,N_49562,N_48200);
xor UO_3011 (O_3011,N_48595,N_49811);
and UO_3012 (O_3012,N_48765,N_48067);
xnor UO_3013 (O_3013,N_49843,N_49498);
xor UO_3014 (O_3014,N_49419,N_49800);
and UO_3015 (O_3015,N_49774,N_48080);
nor UO_3016 (O_3016,N_48148,N_48581);
xor UO_3017 (O_3017,N_49696,N_48448);
xnor UO_3018 (O_3018,N_48486,N_48944);
or UO_3019 (O_3019,N_48395,N_49704);
and UO_3020 (O_3020,N_48955,N_49975);
nor UO_3021 (O_3021,N_49361,N_48827);
xor UO_3022 (O_3022,N_48610,N_49806);
nand UO_3023 (O_3023,N_49625,N_49272);
and UO_3024 (O_3024,N_48416,N_48069);
or UO_3025 (O_3025,N_48128,N_49727);
nor UO_3026 (O_3026,N_48632,N_49898);
nor UO_3027 (O_3027,N_48942,N_49739);
or UO_3028 (O_3028,N_48693,N_48548);
nor UO_3029 (O_3029,N_48666,N_49893);
nor UO_3030 (O_3030,N_48313,N_49928);
nor UO_3031 (O_3031,N_49199,N_48148);
and UO_3032 (O_3032,N_49422,N_49221);
or UO_3033 (O_3033,N_48815,N_48170);
nand UO_3034 (O_3034,N_48715,N_48160);
xor UO_3035 (O_3035,N_49932,N_48343);
and UO_3036 (O_3036,N_48391,N_49388);
or UO_3037 (O_3037,N_48432,N_49816);
and UO_3038 (O_3038,N_48253,N_48986);
or UO_3039 (O_3039,N_49407,N_48949);
nor UO_3040 (O_3040,N_49195,N_48984);
nor UO_3041 (O_3041,N_48186,N_48248);
nor UO_3042 (O_3042,N_48755,N_48065);
or UO_3043 (O_3043,N_49192,N_48108);
xor UO_3044 (O_3044,N_49438,N_49467);
xor UO_3045 (O_3045,N_48669,N_49941);
nor UO_3046 (O_3046,N_49851,N_49397);
and UO_3047 (O_3047,N_49284,N_49164);
nor UO_3048 (O_3048,N_48217,N_48022);
and UO_3049 (O_3049,N_48723,N_48832);
xor UO_3050 (O_3050,N_49317,N_48601);
xor UO_3051 (O_3051,N_48170,N_49665);
nand UO_3052 (O_3052,N_48094,N_49587);
and UO_3053 (O_3053,N_48474,N_48880);
or UO_3054 (O_3054,N_48100,N_49883);
or UO_3055 (O_3055,N_48944,N_49409);
nor UO_3056 (O_3056,N_48435,N_49218);
nor UO_3057 (O_3057,N_48477,N_49606);
nand UO_3058 (O_3058,N_49424,N_49818);
nor UO_3059 (O_3059,N_49966,N_49843);
nand UO_3060 (O_3060,N_49961,N_48074);
or UO_3061 (O_3061,N_49534,N_48530);
or UO_3062 (O_3062,N_48145,N_48319);
and UO_3063 (O_3063,N_49359,N_49571);
or UO_3064 (O_3064,N_48131,N_48086);
nand UO_3065 (O_3065,N_49016,N_49878);
nand UO_3066 (O_3066,N_49238,N_48625);
nor UO_3067 (O_3067,N_48597,N_48275);
xor UO_3068 (O_3068,N_49475,N_48114);
and UO_3069 (O_3069,N_49013,N_48999);
nor UO_3070 (O_3070,N_48447,N_48785);
xnor UO_3071 (O_3071,N_49093,N_49638);
nor UO_3072 (O_3072,N_48010,N_49344);
and UO_3073 (O_3073,N_49438,N_49612);
or UO_3074 (O_3074,N_49712,N_48068);
or UO_3075 (O_3075,N_48802,N_49290);
and UO_3076 (O_3076,N_48771,N_48724);
nor UO_3077 (O_3077,N_48289,N_48202);
nor UO_3078 (O_3078,N_49894,N_48179);
nor UO_3079 (O_3079,N_48482,N_49688);
and UO_3080 (O_3080,N_49874,N_48278);
and UO_3081 (O_3081,N_48239,N_48284);
and UO_3082 (O_3082,N_48035,N_48461);
or UO_3083 (O_3083,N_49559,N_48747);
nand UO_3084 (O_3084,N_48246,N_49643);
nor UO_3085 (O_3085,N_49545,N_48933);
or UO_3086 (O_3086,N_49681,N_48319);
xnor UO_3087 (O_3087,N_48227,N_49858);
nand UO_3088 (O_3088,N_48298,N_48416);
nor UO_3089 (O_3089,N_48411,N_48623);
nand UO_3090 (O_3090,N_49892,N_49500);
and UO_3091 (O_3091,N_49134,N_49211);
nand UO_3092 (O_3092,N_49175,N_49214);
and UO_3093 (O_3093,N_49544,N_48738);
xor UO_3094 (O_3094,N_49777,N_48574);
and UO_3095 (O_3095,N_48982,N_48024);
and UO_3096 (O_3096,N_49377,N_49446);
and UO_3097 (O_3097,N_49299,N_49498);
nand UO_3098 (O_3098,N_48844,N_48423);
nand UO_3099 (O_3099,N_48344,N_49928);
or UO_3100 (O_3100,N_49372,N_49324);
and UO_3101 (O_3101,N_48295,N_49159);
nor UO_3102 (O_3102,N_49118,N_49454);
xor UO_3103 (O_3103,N_48686,N_49250);
nor UO_3104 (O_3104,N_48931,N_49766);
nor UO_3105 (O_3105,N_48865,N_48534);
nand UO_3106 (O_3106,N_48275,N_49961);
nor UO_3107 (O_3107,N_49675,N_48939);
or UO_3108 (O_3108,N_49648,N_48861);
or UO_3109 (O_3109,N_48566,N_48464);
and UO_3110 (O_3110,N_49685,N_48844);
nand UO_3111 (O_3111,N_49200,N_49579);
or UO_3112 (O_3112,N_48838,N_49139);
nand UO_3113 (O_3113,N_48477,N_48896);
nor UO_3114 (O_3114,N_49175,N_48190);
nor UO_3115 (O_3115,N_49275,N_49017);
and UO_3116 (O_3116,N_49859,N_48440);
nand UO_3117 (O_3117,N_49446,N_49385);
xnor UO_3118 (O_3118,N_48996,N_48400);
nor UO_3119 (O_3119,N_49251,N_49513);
or UO_3120 (O_3120,N_49536,N_48301);
and UO_3121 (O_3121,N_49078,N_48025);
nor UO_3122 (O_3122,N_48720,N_49830);
nand UO_3123 (O_3123,N_49090,N_48197);
nor UO_3124 (O_3124,N_48251,N_49275);
nand UO_3125 (O_3125,N_48663,N_49562);
and UO_3126 (O_3126,N_49938,N_48628);
nor UO_3127 (O_3127,N_48441,N_49597);
nor UO_3128 (O_3128,N_49165,N_49171);
or UO_3129 (O_3129,N_49168,N_49558);
xor UO_3130 (O_3130,N_48371,N_49961);
nand UO_3131 (O_3131,N_49587,N_48355);
xnor UO_3132 (O_3132,N_49931,N_48879);
xor UO_3133 (O_3133,N_49071,N_48420);
xor UO_3134 (O_3134,N_48062,N_49292);
and UO_3135 (O_3135,N_49566,N_49074);
nand UO_3136 (O_3136,N_48129,N_49870);
and UO_3137 (O_3137,N_49570,N_49529);
and UO_3138 (O_3138,N_48057,N_48063);
or UO_3139 (O_3139,N_49493,N_49469);
and UO_3140 (O_3140,N_48908,N_48009);
nor UO_3141 (O_3141,N_48334,N_49810);
and UO_3142 (O_3142,N_49646,N_48700);
and UO_3143 (O_3143,N_48894,N_49255);
xor UO_3144 (O_3144,N_49114,N_49827);
and UO_3145 (O_3145,N_48876,N_48820);
xnor UO_3146 (O_3146,N_48353,N_49979);
or UO_3147 (O_3147,N_48824,N_49647);
nor UO_3148 (O_3148,N_48367,N_48284);
nand UO_3149 (O_3149,N_49300,N_48012);
nand UO_3150 (O_3150,N_48258,N_48904);
or UO_3151 (O_3151,N_48820,N_48841);
and UO_3152 (O_3152,N_48562,N_48698);
nand UO_3153 (O_3153,N_48015,N_48223);
nor UO_3154 (O_3154,N_48220,N_49492);
and UO_3155 (O_3155,N_49784,N_48241);
or UO_3156 (O_3156,N_48279,N_48281);
xnor UO_3157 (O_3157,N_48550,N_48020);
nor UO_3158 (O_3158,N_48433,N_49523);
nor UO_3159 (O_3159,N_48286,N_49101);
nor UO_3160 (O_3160,N_48181,N_48665);
nand UO_3161 (O_3161,N_49189,N_48796);
xnor UO_3162 (O_3162,N_49482,N_49025);
and UO_3163 (O_3163,N_48693,N_48219);
xor UO_3164 (O_3164,N_49321,N_49970);
and UO_3165 (O_3165,N_48875,N_48982);
nor UO_3166 (O_3166,N_49925,N_49783);
nand UO_3167 (O_3167,N_48197,N_48840);
or UO_3168 (O_3168,N_49733,N_49766);
and UO_3169 (O_3169,N_49383,N_48637);
nor UO_3170 (O_3170,N_49139,N_49651);
nor UO_3171 (O_3171,N_49788,N_49847);
and UO_3172 (O_3172,N_48834,N_49263);
or UO_3173 (O_3173,N_48507,N_48680);
and UO_3174 (O_3174,N_49149,N_49039);
and UO_3175 (O_3175,N_49486,N_48737);
nor UO_3176 (O_3176,N_48087,N_49540);
nand UO_3177 (O_3177,N_49422,N_49801);
or UO_3178 (O_3178,N_48585,N_49792);
and UO_3179 (O_3179,N_48124,N_48778);
nand UO_3180 (O_3180,N_49446,N_49015);
and UO_3181 (O_3181,N_49840,N_49208);
nor UO_3182 (O_3182,N_49190,N_48179);
nor UO_3183 (O_3183,N_49355,N_48157);
nand UO_3184 (O_3184,N_49014,N_48969);
xor UO_3185 (O_3185,N_48879,N_48675);
and UO_3186 (O_3186,N_49391,N_48743);
xnor UO_3187 (O_3187,N_48496,N_49764);
and UO_3188 (O_3188,N_49965,N_48060);
xnor UO_3189 (O_3189,N_49828,N_48623);
nor UO_3190 (O_3190,N_48709,N_48222);
nand UO_3191 (O_3191,N_49878,N_48840);
and UO_3192 (O_3192,N_48912,N_49830);
nand UO_3193 (O_3193,N_49505,N_48837);
and UO_3194 (O_3194,N_49069,N_48787);
and UO_3195 (O_3195,N_48979,N_49817);
xnor UO_3196 (O_3196,N_49473,N_49570);
and UO_3197 (O_3197,N_49884,N_48210);
xor UO_3198 (O_3198,N_49723,N_48747);
nand UO_3199 (O_3199,N_48630,N_48665);
nor UO_3200 (O_3200,N_48595,N_48327);
nor UO_3201 (O_3201,N_48580,N_49105);
nor UO_3202 (O_3202,N_49598,N_48451);
xnor UO_3203 (O_3203,N_48208,N_49335);
or UO_3204 (O_3204,N_48439,N_49798);
nor UO_3205 (O_3205,N_48001,N_49701);
and UO_3206 (O_3206,N_49917,N_49725);
or UO_3207 (O_3207,N_49761,N_49301);
or UO_3208 (O_3208,N_48609,N_48430);
nand UO_3209 (O_3209,N_49263,N_48592);
or UO_3210 (O_3210,N_49402,N_49017);
xor UO_3211 (O_3211,N_49073,N_48996);
xor UO_3212 (O_3212,N_48775,N_49178);
and UO_3213 (O_3213,N_49442,N_49099);
nor UO_3214 (O_3214,N_49403,N_49336);
nor UO_3215 (O_3215,N_48922,N_49100);
or UO_3216 (O_3216,N_48126,N_49428);
nand UO_3217 (O_3217,N_48605,N_49933);
and UO_3218 (O_3218,N_49073,N_48161);
or UO_3219 (O_3219,N_48345,N_48879);
and UO_3220 (O_3220,N_49186,N_48372);
xnor UO_3221 (O_3221,N_48268,N_48334);
nor UO_3222 (O_3222,N_49768,N_49715);
and UO_3223 (O_3223,N_49151,N_49197);
or UO_3224 (O_3224,N_48484,N_48189);
or UO_3225 (O_3225,N_48571,N_49038);
nor UO_3226 (O_3226,N_48694,N_49052);
nor UO_3227 (O_3227,N_48608,N_48828);
xnor UO_3228 (O_3228,N_49701,N_49194);
nor UO_3229 (O_3229,N_48260,N_49698);
nand UO_3230 (O_3230,N_48406,N_48619);
nand UO_3231 (O_3231,N_49435,N_49220);
or UO_3232 (O_3232,N_48984,N_48661);
nand UO_3233 (O_3233,N_49925,N_48060);
or UO_3234 (O_3234,N_48979,N_49093);
nand UO_3235 (O_3235,N_49007,N_48359);
and UO_3236 (O_3236,N_49263,N_49406);
and UO_3237 (O_3237,N_49352,N_48601);
or UO_3238 (O_3238,N_48150,N_49209);
and UO_3239 (O_3239,N_48226,N_48021);
nor UO_3240 (O_3240,N_48740,N_48106);
xnor UO_3241 (O_3241,N_48708,N_48375);
xnor UO_3242 (O_3242,N_48620,N_49606);
xor UO_3243 (O_3243,N_49045,N_48546);
and UO_3244 (O_3244,N_49001,N_48771);
and UO_3245 (O_3245,N_49362,N_49658);
nand UO_3246 (O_3246,N_49694,N_49822);
xnor UO_3247 (O_3247,N_48760,N_49211);
and UO_3248 (O_3248,N_48205,N_49212);
or UO_3249 (O_3249,N_49452,N_48471);
xor UO_3250 (O_3250,N_49526,N_48014);
and UO_3251 (O_3251,N_49411,N_49531);
xnor UO_3252 (O_3252,N_49621,N_48609);
or UO_3253 (O_3253,N_49742,N_48856);
xnor UO_3254 (O_3254,N_48374,N_48953);
xnor UO_3255 (O_3255,N_49678,N_49103);
xnor UO_3256 (O_3256,N_48048,N_49793);
or UO_3257 (O_3257,N_49448,N_49195);
xnor UO_3258 (O_3258,N_48962,N_49908);
nand UO_3259 (O_3259,N_48390,N_48098);
or UO_3260 (O_3260,N_48424,N_48456);
and UO_3261 (O_3261,N_48273,N_48848);
or UO_3262 (O_3262,N_49305,N_49370);
or UO_3263 (O_3263,N_48499,N_49520);
nor UO_3264 (O_3264,N_49264,N_49442);
xor UO_3265 (O_3265,N_48646,N_49931);
nor UO_3266 (O_3266,N_49910,N_49273);
and UO_3267 (O_3267,N_48476,N_48650);
nor UO_3268 (O_3268,N_48563,N_49901);
nor UO_3269 (O_3269,N_49811,N_49116);
nor UO_3270 (O_3270,N_48257,N_48891);
or UO_3271 (O_3271,N_49199,N_49671);
xor UO_3272 (O_3272,N_49669,N_49684);
nand UO_3273 (O_3273,N_49371,N_49284);
nand UO_3274 (O_3274,N_48493,N_49195);
xnor UO_3275 (O_3275,N_49981,N_49291);
and UO_3276 (O_3276,N_48223,N_48259);
nor UO_3277 (O_3277,N_49373,N_48482);
nor UO_3278 (O_3278,N_49540,N_48737);
nand UO_3279 (O_3279,N_48376,N_49133);
xor UO_3280 (O_3280,N_49470,N_49676);
nand UO_3281 (O_3281,N_48047,N_48681);
xnor UO_3282 (O_3282,N_48458,N_49140);
nand UO_3283 (O_3283,N_49825,N_49538);
nor UO_3284 (O_3284,N_49242,N_48108);
xor UO_3285 (O_3285,N_49208,N_49858);
and UO_3286 (O_3286,N_48225,N_48870);
xor UO_3287 (O_3287,N_48922,N_48862);
nand UO_3288 (O_3288,N_48837,N_49478);
nand UO_3289 (O_3289,N_49339,N_48830);
xor UO_3290 (O_3290,N_48201,N_48683);
or UO_3291 (O_3291,N_48842,N_49249);
nand UO_3292 (O_3292,N_48311,N_48655);
nand UO_3293 (O_3293,N_48891,N_48340);
nand UO_3294 (O_3294,N_49014,N_48050);
or UO_3295 (O_3295,N_48387,N_49289);
or UO_3296 (O_3296,N_48272,N_48903);
nand UO_3297 (O_3297,N_48605,N_48414);
xnor UO_3298 (O_3298,N_49571,N_48573);
nand UO_3299 (O_3299,N_48074,N_48836);
xor UO_3300 (O_3300,N_49642,N_48849);
or UO_3301 (O_3301,N_49569,N_48056);
nor UO_3302 (O_3302,N_49670,N_48061);
or UO_3303 (O_3303,N_49161,N_48735);
nor UO_3304 (O_3304,N_48866,N_48720);
nor UO_3305 (O_3305,N_49287,N_48702);
or UO_3306 (O_3306,N_49028,N_49951);
nand UO_3307 (O_3307,N_49102,N_48290);
or UO_3308 (O_3308,N_49745,N_48303);
nor UO_3309 (O_3309,N_49636,N_48115);
and UO_3310 (O_3310,N_49921,N_48778);
nor UO_3311 (O_3311,N_48899,N_49697);
xnor UO_3312 (O_3312,N_49685,N_49845);
and UO_3313 (O_3313,N_49549,N_49932);
or UO_3314 (O_3314,N_49627,N_48704);
xor UO_3315 (O_3315,N_49369,N_49133);
xnor UO_3316 (O_3316,N_48655,N_48156);
nand UO_3317 (O_3317,N_48009,N_48997);
nand UO_3318 (O_3318,N_49000,N_49989);
and UO_3319 (O_3319,N_48382,N_48788);
xnor UO_3320 (O_3320,N_49548,N_48258);
nor UO_3321 (O_3321,N_48931,N_49644);
or UO_3322 (O_3322,N_49782,N_49442);
nand UO_3323 (O_3323,N_49220,N_49606);
or UO_3324 (O_3324,N_48902,N_49665);
or UO_3325 (O_3325,N_49224,N_49077);
xnor UO_3326 (O_3326,N_48929,N_48335);
xnor UO_3327 (O_3327,N_49675,N_49896);
nand UO_3328 (O_3328,N_49970,N_48021);
nor UO_3329 (O_3329,N_49598,N_49301);
xor UO_3330 (O_3330,N_48077,N_49157);
xnor UO_3331 (O_3331,N_48764,N_49672);
or UO_3332 (O_3332,N_49805,N_49768);
or UO_3333 (O_3333,N_49229,N_49005);
or UO_3334 (O_3334,N_48989,N_48052);
and UO_3335 (O_3335,N_48512,N_49228);
or UO_3336 (O_3336,N_48151,N_49018);
nand UO_3337 (O_3337,N_49152,N_48050);
nor UO_3338 (O_3338,N_49682,N_48256);
xnor UO_3339 (O_3339,N_49115,N_49436);
or UO_3340 (O_3340,N_49736,N_48308);
nand UO_3341 (O_3341,N_48655,N_48509);
or UO_3342 (O_3342,N_48693,N_48516);
xor UO_3343 (O_3343,N_49364,N_49335);
nor UO_3344 (O_3344,N_48595,N_48504);
and UO_3345 (O_3345,N_49566,N_49101);
xnor UO_3346 (O_3346,N_48923,N_49263);
nand UO_3347 (O_3347,N_48642,N_49796);
or UO_3348 (O_3348,N_48437,N_48386);
nand UO_3349 (O_3349,N_48405,N_49649);
nand UO_3350 (O_3350,N_48323,N_49374);
or UO_3351 (O_3351,N_49741,N_48739);
or UO_3352 (O_3352,N_48603,N_49168);
and UO_3353 (O_3353,N_48612,N_49608);
and UO_3354 (O_3354,N_48473,N_48000);
and UO_3355 (O_3355,N_49719,N_49776);
xnor UO_3356 (O_3356,N_48248,N_48278);
and UO_3357 (O_3357,N_48337,N_49730);
nor UO_3358 (O_3358,N_48974,N_48822);
or UO_3359 (O_3359,N_48632,N_48214);
nor UO_3360 (O_3360,N_48733,N_49114);
nand UO_3361 (O_3361,N_48919,N_49396);
nor UO_3362 (O_3362,N_49707,N_49850);
nor UO_3363 (O_3363,N_49989,N_48320);
and UO_3364 (O_3364,N_49792,N_49359);
nor UO_3365 (O_3365,N_48360,N_48534);
and UO_3366 (O_3366,N_49938,N_48896);
or UO_3367 (O_3367,N_49469,N_49851);
nand UO_3368 (O_3368,N_48453,N_49271);
and UO_3369 (O_3369,N_49920,N_48474);
or UO_3370 (O_3370,N_48340,N_49107);
nand UO_3371 (O_3371,N_48931,N_48319);
and UO_3372 (O_3372,N_49810,N_48190);
and UO_3373 (O_3373,N_48518,N_49537);
xor UO_3374 (O_3374,N_48981,N_49442);
nor UO_3375 (O_3375,N_49188,N_48011);
or UO_3376 (O_3376,N_48105,N_49054);
and UO_3377 (O_3377,N_49595,N_49435);
nand UO_3378 (O_3378,N_48726,N_48479);
or UO_3379 (O_3379,N_49509,N_49724);
nand UO_3380 (O_3380,N_48291,N_49467);
nand UO_3381 (O_3381,N_48270,N_48114);
nand UO_3382 (O_3382,N_48705,N_49920);
xor UO_3383 (O_3383,N_49416,N_48863);
and UO_3384 (O_3384,N_48329,N_49973);
nor UO_3385 (O_3385,N_48808,N_49691);
xnor UO_3386 (O_3386,N_49416,N_48658);
nor UO_3387 (O_3387,N_48517,N_49227);
xnor UO_3388 (O_3388,N_49270,N_48042);
nand UO_3389 (O_3389,N_48777,N_49638);
nand UO_3390 (O_3390,N_49658,N_48615);
and UO_3391 (O_3391,N_48746,N_48537);
and UO_3392 (O_3392,N_49092,N_49525);
or UO_3393 (O_3393,N_48994,N_49482);
and UO_3394 (O_3394,N_48011,N_48042);
nor UO_3395 (O_3395,N_48753,N_49416);
nand UO_3396 (O_3396,N_49785,N_49417);
nand UO_3397 (O_3397,N_49061,N_48547);
nor UO_3398 (O_3398,N_48221,N_49060);
or UO_3399 (O_3399,N_49564,N_49055);
xor UO_3400 (O_3400,N_49392,N_49020);
nor UO_3401 (O_3401,N_49451,N_48585);
and UO_3402 (O_3402,N_48404,N_48666);
or UO_3403 (O_3403,N_49061,N_49069);
nand UO_3404 (O_3404,N_49441,N_49746);
or UO_3405 (O_3405,N_49653,N_48904);
and UO_3406 (O_3406,N_49885,N_48845);
and UO_3407 (O_3407,N_49671,N_49672);
and UO_3408 (O_3408,N_49796,N_49230);
nor UO_3409 (O_3409,N_48054,N_49155);
nor UO_3410 (O_3410,N_49341,N_48288);
or UO_3411 (O_3411,N_49771,N_49768);
nor UO_3412 (O_3412,N_49226,N_48310);
xnor UO_3413 (O_3413,N_49687,N_49912);
nand UO_3414 (O_3414,N_49123,N_49202);
nor UO_3415 (O_3415,N_49070,N_48052);
and UO_3416 (O_3416,N_49033,N_49825);
and UO_3417 (O_3417,N_48326,N_49725);
xor UO_3418 (O_3418,N_49547,N_49026);
nand UO_3419 (O_3419,N_48408,N_48901);
and UO_3420 (O_3420,N_49507,N_49483);
xnor UO_3421 (O_3421,N_49149,N_49935);
and UO_3422 (O_3422,N_48336,N_48276);
nor UO_3423 (O_3423,N_48644,N_49387);
nand UO_3424 (O_3424,N_48126,N_48760);
or UO_3425 (O_3425,N_48797,N_49920);
or UO_3426 (O_3426,N_49017,N_48981);
and UO_3427 (O_3427,N_48435,N_49885);
nand UO_3428 (O_3428,N_49036,N_48122);
nand UO_3429 (O_3429,N_49266,N_48575);
nand UO_3430 (O_3430,N_49811,N_49196);
or UO_3431 (O_3431,N_48970,N_48344);
xnor UO_3432 (O_3432,N_49444,N_48181);
xor UO_3433 (O_3433,N_48959,N_48694);
and UO_3434 (O_3434,N_49179,N_49584);
and UO_3435 (O_3435,N_49875,N_48290);
nand UO_3436 (O_3436,N_49754,N_49287);
nor UO_3437 (O_3437,N_49907,N_49062);
nand UO_3438 (O_3438,N_49151,N_49638);
nor UO_3439 (O_3439,N_48213,N_48877);
nand UO_3440 (O_3440,N_49662,N_48543);
and UO_3441 (O_3441,N_48670,N_49322);
and UO_3442 (O_3442,N_49115,N_49817);
nand UO_3443 (O_3443,N_49476,N_49348);
xor UO_3444 (O_3444,N_49014,N_48660);
or UO_3445 (O_3445,N_48603,N_48554);
and UO_3446 (O_3446,N_49706,N_49758);
nor UO_3447 (O_3447,N_48343,N_48825);
and UO_3448 (O_3448,N_48777,N_49933);
xor UO_3449 (O_3449,N_49781,N_49752);
nand UO_3450 (O_3450,N_49660,N_49766);
xor UO_3451 (O_3451,N_49709,N_48132);
and UO_3452 (O_3452,N_48302,N_49619);
or UO_3453 (O_3453,N_48910,N_49424);
nand UO_3454 (O_3454,N_49649,N_49136);
xor UO_3455 (O_3455,N_48352,N_48608);
nor UO_3456 (O_3456,N_48690,N_49155);
xnor UO_3457 (O_3457,N_48535,N_49587);
or UO_3458 (O_3458,N_49385,N_48819);
and UO_3459 (O_3459,N_49765,N_49902);
nand UO_3460 (O_3460,N_49375,N_48081);
and UO_3461 (O_3461,N_49826,N_48213);
or UO_3462 (O_3462,N_48368,N_49121);
or UO_3463 (O_3463,N_48808,N_49104);
nor UO_3464 (O_3464,N_49351,N_49601);
nand UO_3465 (O_3465,N_49586,N_49901);
or UO_3466 (O_3466,N_48506,N_49161);
or UO_3467 (O_3467,N_48816,N_48924);
nand UO_3468 (O_3468,N_49093,N_48279);
or UO_3469 (O_3469,N_49425,N_48519);
or UO_3470 (O_3470,N_48541,N_48003);
nand UO_3471 (O_3471,N_48064,N_48092);
and UO_3472 (O_3472,N_48797,N_49838);
or UO_3473 (O_3473,N_49522,N_49792);
nor UO_3474 (O_3474,N_49893,N_49166);
xor UO_3475 (O_3475,N_48188,N_48471);
or UO_3476 (O_3476,N_49112,N_48451);
xnor UO_3477 (O_3477,N_49390,N_48919);
nand UO_3478 (O_3478,N_49970,N_48822);
nor UO_3479 (O_3479,N_49885,N_48086);
or UO_3480 (O_3480,N_48390,N_49053);
xnor UO_3481 (O_3481,N_49902,N_49776);
xor UO_3482 (O_3482,N_48411,N_49324);
nand UO_3483 (O_3483,N_49734,N_49402);
xor UO_3484 (O_3484,N_48350,N_49632);
xnor UO_3485 (O_3485,N_48292,N_49534);
or UO_3486 (O_3486,N_48430,N_48812);
and UO_3487 (O_3487,N_48365,N_48900);
or UO_3488 (O_3488,N_48659,N_48597);
or UO_3489 (O_3489,N_48844,N_48704);
nand UO_3490 (O_3490,N_49215,N_48903);
or UO_3491 (O_3491,N_48195,N_49746);
xor UO_3492 (O_3492,N_49196,N_49354);
or UO_3493 (O_3493,N_48413,N_49307);
and UO_3494 (O_3494,N_48541,N_48710);
or UO_3495 (O_3495,N_48660,N_49375);
nand UO_3496 (O_3496,N_49776,N_48626);
nand UO_3497 (O_3497,N_49244,N_48574);
nor UO_3498 (O_3498,N_48351,N_49392);
or UO_3499 (O_3499,N_49239,N_48019);
or UO_3500 (O_3500,N_49660,N_49680);
nor UO_3501 (O_3501,N_48335,N_48567);
xor UO_3502 (O_3502,N_48161,N_48089);
and UO_3503 (O_3503,N_48032,N_49588);
nand UO_3504 (O_3504,N_48778,N_48946);
nand UO_3505 (O_3505,N_48570,N_48386);
nand UO_3506 (O_3506,N_48148,N_49609);
nand UO_3507 (O_3507,N_49984,N_49619);
xor UO_3508 (O_3508,N_48821,N_49933);
or UO_3509 (O_3509,N_49774,N_49007);
nand UO_3510 (O_3510,N_49786,N_49461);
or UO_3511 (O_3511,N_48388,N_49098);
or UO_3512 (O_3512,N_48060,N_48936);
and UO_3513 (O_3513,N_48952,N_49814);
nor UO_3514 (O_3514,N_49638,N_48986);
nand UO_3515 (O_3515,N_48429,N_49188);
xnor UO_3516 (O_3516,N_48810,N_49507);
nand UO_3517 (O_3517,N_48978,N_48857);
and UO_3518 (O_3518,N_48840,N_48686);
or UO_3519 (O_3519,N_48449,N_48096);
xnor UO_3520 (O_3520,N_48508,N_49376);
or UO_3521 (O_3521,N_48361,N_48999);
nand UO_3522 (O_3522,N_48926,N_48860);
nand UO_3523 (O_3523,N_48593,N_48217);
or UO_3524 (O_3524,N_49632,N_49604);
and UO_3525 (O_3525,N_49299,N_49303);
or UO_3526 (O_3526,N_49156,N_49070);
and UO_3527 (O_3527,N_48574,N_49702);
nor UO_3528 (O_3528,N_48163,N_49560);
or UO_3529 (O_3529,N_49512,N_49009);
nor UO_3530 (O_3530,N_49183,N_49606);
xor UO_3531 (O_3531,N_49531,N_48211);
and UO_3532 (O_3532,N_49449,N_48794);
or UO_3533 (O_3533,N_48727,N_49312);
xor UO_3534 (O_3534,N_48827,N_49586);
xnor UO_3535 (O_3535,N_48287,N_49688);
nor UO_3536 (O_3536,N_49637,N_48017);
and UO_3537 (O_3537,N_48856,N_48867);
nor UO_3538 (O_3538,N_48617,N_49363);
xor UO_3539 (O_3539,N_49109,N_48070);
nor UO_3540 (O_3540,N_49420,N_49035);
and UO_3541 (O_3541,N_48050,N_49158);
nand UO_3542 (O_3542,N_49890,N_48124);
xnor UO_3543 (O_3543,N_49430,N_48961);
and UO_3544 (O_3544,N_49595,N_48492);
and UO_3545 (O_3545,N_48338,N_48119);
nor UO_3546 (O_3546,N_49119,N_48230);
xnor UO_3547 (O_3547,N_48732,N_49706);
and UO_3548 (O_3548,N_48747,N_48202);
nand UO_3549 (O_3549,N_49079,N_49528);
and UO_3550 (O_3550,N_49795,N_49438);
nor UO_3551 (O_3551,N_48811,N_48916);
or UO_3552 (O_3552,N_48326,N_49640);
or UO_3553 (O_3553,N_49492,N_48082);
and UO_3554 (O_3554,N_48643,N_49768);
nor UO_3555 (O_3555,N_48022,N_49466);
nor UO_3556 (O_3556,N_48932,N_49326);
or UO_3557 (O_3557,N_48035,N_49417);
nand UO_3558 (O_3558,N_48372,N_48434);
xnor UO_3559 (O_3559,N_48417,N_49445);
xor UO_3560 (O_3560,N_48220,N_48023);
and UO_3561 (O_3561,N_49435,N_49479);
nor UO_3562 (O_3562,N_49527,N_49681);
or UO_3563 (O_3563,N_49359,N_49863);
and UO_3564 (O_3564,N_48742,N_49249);
or UO_3565 (O_3565,N_49909,N_48033);
xor UO_3566 (O_3566,N_48101,N_48933);
xnor UO_3567 (O_3567,N_49273,N_49790);
nand UO_3568 (O_3568,N_49042,N_48245);
xnor UO_3569 (O_3569,N_49196,N_48653);
xor UO_3570 (O_3570,N_49401,N_49788);
and UO_3571 (O_3571,N_48515,N_49802);
nand UO_3572 (O_3572,N_48439,N_49799);
and UO_3573 (O_3573,N_48864,N_49893);
nor UO_3574 (O_3574,N_48544,N_49850);
or UO_3575 (O_3575,N_49500,N_49701);
nor UO_3576 (O_3576,N_48539,N_49828);
or UO_3577 (O_3577,N_49946,N_49023);
nand UO_3578 (O_3578,N_48014,N_48485);
or UO_3579 (O_3579,N_48209,N_49339);
or UO_3580 (O_3580,N_49627,N_48619);
nand UO_3581 (O_3581,N_49494,N_49629);
xnor UO_3582 (O_3582,N_48956,N_48852);
or UO_3583 (O_3583,N_48386,N_49806);
or UO_3584 (O_3584,N_49858,N_48481);
or UO_3585 (O_3585,N_48343,N_49583);
xnor UO_3586 (O_3586,N_49187,N_48315);
nor UO_3587 (O_3587,N_48162,N_48284);
or UO_3588 (O_3588,N_49829,N_48271);
nand UO_3589 (O_3589,N_49087,N_49674);
and UO_3590 (O_3590,N_48995,N_48523);
or UO_3591 (O_3591,N_48149,N_48027);
or UO_3592 (O_3592,N_49579,N_48571);
or UO_3593 (O_3593,N_49485,N_48633);
or UO_3594 (O_3594,N_48094,N_49338);
or UO_3595 (O_3595,N_48615,N_49625);
or UO_3596 (O_3596,N_48764,N_49393);
and UO_3597 (O_3597,N_49379,N_48066);
nor UO_3598 (O_3598,N_48049,N_48457);
or UO_3599 (O_3599,N_48478,N_48093);
nand UO_3600 (O_3600,N_48234,N_48281);
and UO_3601 (O_3601,N_48237,N_49042);
or UO_3602 (O_3602,N_49145,N_49931);
xnor UO_3603 (O_3603,N_49003,N_49015);
and UO_3604 (O_3604,N_49867,N_49425);
nor UO_3605 (O_3605,N_48725,N_49980);
nor UO_3606 (O_3606,N_48955,N_49274);
nor UO_3607 (O_3607,N_49233,N_49103);
and UO_3608 (O_3608,N_48977,N_48080);
or UO_3609 (O_3609,N_49639,N_48466);
nor UO_3610 (O_3610,N_48656,N_49752);
nand UO_3611 (O_3611,N_48162,N_48211);
and UO_3612 (O_3612,N_49734,N_48817);
xnor UO_3613 (O_3613,N_48242,N_49644);
or UO_3614 (O_3614,N_49927,N_49235);
xor UO_3615 (O_3615,N_49744,N_49609);
nand UO_3616 (O_3616,N_49109,N_48540);
and UO_3617 (O_3617,N_48812,N_49628);
or UO_3618 (O_3618,N_48175,N_49852);
and UO_3619 (O_3619,N_48345,N_49218);
nand UO_3620 (O_3620,N_48861,N_48096);
or UO_3621 (O_3621,N_49234,N_49810);
nand UO_3622 (O_3622,N_48103,N_48497);
nor UO_3623 (O_3623,N_49601,N_48989);
xor UO_3624 (O_3624,N_48239,N_48687);
nor UO_3625 (O_3625,N_48963,N_49480);
and UO_3626 (O_3626,N_49954,N_48637);
nor UO_3627 (O_3627,N_49854,N_48335);
and UO_3628 (O_3628,N_49168,N_49677);
and UO_3629 (O_3629,N_49098,N_49460);
xor UO_3630 (O_3630,N_48881,N_49071);
or UO_3631 (O_3631,N_48818,N_49153);
nand UO_3632 (O_3632,N_49165,N_48426);
or UO_3633 (O_3633,N_49059,N_49708);
or UO_3634 (O_3634,N_48920,N_49433);
xnor UO_3635 (O_3635,N_49192,N_48344);
or UO_3636 (O_3636,N_49930,N_48933);
or UO_3637 (O_3637,N_49484,N_49044);
or UO_3638 (O_3638,N_48966,N_48925);
nand UO_3639 (O_3639,N_48540,N_49108);
nand UO_3640 (O_3640,N_49912,N_48036);
nand UO_3641 (O_3641,N_49536,N_48636);
or UO_3642 (O_3642,N_48027,N_49112);
and UO_3643 (O_3643,N_49265,N_49211);
or UO_3644 (O_3644,N_48694,N_49161);
or UO_3645 (O_3645,N_48424,N_49874);
xor UO_3646 (O_3646,N_48161,N_49084);
nand UO_3647 (O_3647,N_49622,N_49464);
or UO_3648 (O_3648,N_48258,N_49593);
or UO_3649 (O_3649,N_48671,N_48447);
xor UO_3650 (O_3650,N_48187,N_49918);
nor UO_3651 (O_3651,N_48473,N_48938);
and UO_3652 (O_3652,N_48382,N_49672);
and UO_3653 (O_3653,N_49707,N_48002);
or UO_3654 (O_3654,N_48564,N_49593);
nor UO_3655 (O_3655,N_48825,N_48098);
nor UO_3656 (O_3656,N_48304,N_49476);
nand UO_3657 (O_3657,N_48656,N_48493);
or UO_3658 (O_3658,N_48843,N_48992);
and UO_3659 (O_3659,N_49166,N_49541);
nand UO_3660 (O_3660,N_48127,N_48355);
and UO_3661 (O_3661,N_49986,N_49736);
and UO_3662 (O_3662,N_48922,N_48568);
and UO_3663 (O_3663,N_49367,N_49706);
and UO_3664 (O_3664,N_48392,N_48378);
and UO_3665 (O_3665,N_49989,N_48638);
and UO_3666 (O_3666,N_49835,N_48654);
nand UO_3667 (O_3667,N_49257,N_49639);
and UO_3668 (O_3668,N_49827,N_48854);
xnor UO_3669 (O_3669,N_48782,N_49350);
nand UO_3670 (O_3670,N_49545,N_49002);
nor UO_3671 (O_3671,N_48382,N_48600);
nor UO_3672 (O_3672,N_49278,N_49537);
or UO_3673 (O_3673,N_49198,N_49150);
xor UO_3674 (O_3674,N_49997,N_48029);
nand UO_3675 (O_3675,N_48681,N_49258);
nand UO_3676 (O_3676,N_48968,N_48734);
or UO_3677 (O_3677,N_48605,N_48697);
nor UO_3678 (O_3678,N_49949,N_48835);
and UO_3679 (O_3679,N_48166,N_48211);
and UO_3680 (O_3680,N_48912,N_49733);
xor UO_3681 (O_3681,N_49629,N_48516);
xnor UO_3682 (O_3682,N_49427,N_49426);
nor UO_3683 (O_3683,N_49825,N_49066);
xor UO_3684 (O_3684,N_48492,N_49730);
and UO_3685 (O_3685,N_48413,N_48230);
nand UO_3686 (O_3686,N_49155,N_48815);
and UO_3687 (O_3687,N_48695,N_49803);
and UO_3688 (O_3688,N_49794,N_49613);
or UO_3689 (O_3689,N_48628,N_49361);
nor UO_3690 (O_3690,N_49469,N_48875);
and UO_3691 (O_3691,N_48882,N_48446);
or UO_3692 (O_3692,N_48533,N_48890);
xor UO_3693 (O_3693,N_48566,N_49811);
xor UO_3694 (O_3694,N_49913,N_48434);
xor UO_3695 (O_3695,N_49071,N_49956);
and UO_3696 (O_3696,N_48370,N_49309);
nand UO_3697 (O_3697,N_49274,N_48247);
xor UO_3698 (O_3698,N_49218,N_49440);
xor UO_3699 (O_3699,N_49207,N_49972);
nor UO_3700 (O_3700,N_48221,N_49809);
or UO_3701 (O_3701,N_48090,N_49292);
xnor UO_3702 (O_3702,N_48719,N_49998);
nand UO_3703 (O_3703,N_48896,N_48336);
and UO_3704 (O_3704,N_49786,N_48925);
or UO_3705 (O_3705,N_48778,N_49947);
and UO_3706 (O_3706,N_48347,N_48076);
xnor UO_3707 (O_3707,N_49351,N_49855);
nand UO_3708 (O_3708,N_49612,N_49905);
xnor UO_3709 (O_3709,N_48888,N_48146);
nand UO_3710 (O_3710,N_48219,N_49822);
or UO_3711 (O_3711,N_48399,N_48712);
nand UO_3712 (O_3712,N_48528,N_49918);
nor UO_3713 (O_3713,N_49141,N_49614);
nand UO_3714 (O_3714,N_48894,N_48028);
xor UO_3715 (O_3715,N_49507,N_49009);
xnor UO_3716 (O_3716,N_48855,N_49794);
nor UO_3717 (O_3717,N_48400,N_49130);
nand UO_3718 (O_3718,N_48831,N_48819);
nand UO_3719 (O_3719,N_49744,N_48885);
and UO_3720 (O_3720,N_48028,N_48471);
nand UO_3721 (O_3721,N_49220,N_48840);
or UO_3722 (O_3722,N_49607,N_48483);
and UO_3723 (O_3723,N_48166,N_49608);
and UO_3724 (O_3724,N_49880,N_48805);
nand UO_3725 (O_3725,N_48197,N_48470);
xnor UO_3726 (O_3726,N_49857,N_48108);
nand UO_3727 (O_3727,N_49203,N_48379);
xnor UO_3728 (O_3728,N_48696,N_48638);
nand UO_3729 (O_3729,N_49843,N_48580);
xor UO_3730 (O_3730,N_49169,N_49259);
and UO_3731 (O_3731,N_48667,N_48791);
xnor UO_3732 (O_3732,N_48665,N_49968);
xor UO_3733 (O_3733,N_49457,N_49461);
and UO_3734 (O_3734,N_49321,N_48292);
nor UO_3735 (O_3735,N_49013,N_49667);
xnor UO_3736 (O_3736,N_49823,N_48312);
nand UO_3737 (O_3737,N_49026,N_49642);
xnor UO_3738 (O_3738,N_48509,N_48440);
nor UO_3739 (O_3739,N_48257,N_49142);
nor UO_3740 (O_3740,N_49153,N_49130);
xor UO_3741 (O_3741,N_48411,N_48441);
or UO_3742 (O_3742,N_49864,N_49058);
xor UO_3743 (O_3743,N_49409,N_49285);
and UO_3744 (O_3744,N_48381,N_49437);
or UO_3745 (O_3745,N_49579,N_49839);
or UO_3746 (O_3746,N_49745,N_48409);
xnor UO_3747 (O_3747,N_49465,N_49908);
nor UO_3748 (O_3748,N_48398,N_48909);
xnor UO_3749 (O_3749,N_48499,N_49044);
and UO_3750 (O_3750,N_49530,N_49083);
nand UO_3751 (O_3751,N_48188,N_49679);
and UO_3752 (O_3752,N_49474,N_48775);
or UO_3753 (O_3753,N_49708,N_49287);
or UO_3754 (O_3754,N_48602,N_49779);
or UO_3755 (O_3755,N_48963,N_49661);
xor UO_3756 (O_3756,N_48456,N_48352);
and UO_3757 (O_3757,N_48118,N_49043);
xnor UO_3758 (O_3758,N_49223,N_48816);
nor UO_3759 (O_3759,N_49556,N_49243);
nand UO_3760 (O_3760,N_49697,N_48023);
nand UO_3761 (O_3761,N_49786,N_48072);
or UO_3762 (O_3762,N_48177,N_48963);
or UO_3763 (O_3763,N_48923,N_48102);
or UO_3764 (O_3764,N_48435,N_49567);
or UO_3765 (O_3765,N_48773,N_49826);
xor UO_3766 (O_3766,N_48265,N_48429);
or UO_3767 (O_3767,N_49768,N_48477);
xor UO_3768 (O_3768,N_49070,N_48186);
xor UO_3769 (O_3769,N_49628,N_48492);
xnor UO_3770 (O_3770,N_49516,N_49199);
nor UO_3771 (O_3771,N_49207,N_48797);
nor UO_3772 (O_3772,N_48353,N_49638);
or UO_3773 (O_3773,N_48100,N_48977);
nor UO_3774 (O_3774,N_49179,N_49482);
xor UO_3775 (O_3775,N_48378,N_48918);
xnor UO_3776 (O_3776,N_49448,N_49368);
xnor UO_3777 (O_3777,N_49651,N_48915);
xor UO_3778 (O_3778,N_48327,N_48791);
and UO_3779 (O_3779,N_48321,N_49522);
xnor UO_3780 (O_3780,N_48800,N_48872);
or UO_3781 (O_3781,N_49754,N_48732);
xor UO_3782 (O_3782,N_49836,N_49513);
nor UO_3783 (O_3783,N_49586,N_48704);
xnor UO_3784 (O_3784,N_48126,N_49441);
nor UO_3785 (O_3785,N_48793,N_48782);
and UO_3786 (O_3786,N_49038,N_49246);
or UO_3787 (O_3787,N_49231,N_48093);
and UO_3788 (O_3788,N_48830,N_48471);
nand UO_3789 (O_3789,N_48510,N_48238);
nor UO_3790 (O_3790,N_48315,N_48517);
and UO_3791 (O_3791,N_48086,N_49520);
nor UO_3792 (O_3792,N_48740,N_48985);
nor UO_3793 (O_3793,N_48112,N_48269);
nor UO_3794 (O_3794,N_48068,N_49999);
and UO_3795 (O_3795,N_49311,N_49986);
nand UO_3796 (O_3796,N_48580,N_48887);
nor UO_3797 (O_3797,N_49226,N_48014);
and UO_3798 (O_3798,N_49060,N_48460);
or UO_3799 (O_3799,N_48784,N_49333);
or UO_3800 (O_3800,N_48981,N_48408);
or UO_3801 (O_3801,N_49639,N_49499);
and UO_3802 (O_3802,N_49138,N_48272);
or UO_3803 (O_3803,N_48534,N_48883);
nand UO_3804 (O_3804,N_49950,N_49002);
or UO_3805 (O_3805,N_49661,N_48282);
or UO_3806 (O_3806,N_48365,N_49004);
xor UO_3807 (O_3807,N_49341,N_49918);
or UO_3808 (O_3808,N_48417,N_49505);
xnor UO_3809 (O_3809,N_48245,N_48006);
nand UO_3810 (O_3810,N_49063,N_49911);
or UO_3811 (O_3811,N_49771,N_48057);
nor UO_3812 (O_3812,N_48636,N_48480);
nand UO_3813 (O_3813,N_48935,N_49036);
and UO_3814 (O_3814,N_48403,N_49149);
nor UO_3815 (O_3815,N_49616,N_48710);
xnor UO_3816 (O_3816,N_49229,N_48210);
nor UO_3817 (O_3817,N_48829,N_49441);
nor UO_3818 (O_3818,N_49245,N_48809);
nand UO_3819 (O_3819,N_48076,N_49027);
or UO_3820 (O_3820,N_49801,N_49296);
or UO_3821 (O_3821,N_49245,N_48730);
nand UO_3822 (O_3822,N_49937,N_48387);
or UO_3823 (O_3823,N_48150,N_48925);
nor UO_3824 (O_3824,N_49648,N_48019);
nor UO_3825 (O_3825,N_48938,N_48970);
nand UO_3826 (O_3826,N_48594,N_49415);
or UO_3827 (O_3827,N_49030,N_49306);
nor UO_3828 (O_3828,N_48043,N_48155);
and UO_3829 (O_3829,N_49284,N_49225);
or UO_3830 (O_3830,N_49215,N_48792);
xnor UO_3831 (O_3831,N_49654,N_48561);
or UO_3832 (O_3832,N_49177,N_49482);
nand UO_3833 (O_3833,N_49329,N_49357);
or UO_3834 (O_3834,N_49041,N_49275);
nand UO_3835 (O_3835,N_49262,N_49040);
and UO_3836 (O_3836,N_49222,N_48549);
xnor UO_3837 (O_3837,N_49897,N_48402);
nor UO_3838 (O_3838,N_49454,N_48027);
xor UO_3839 (O_3839,N_48879,N_49405);
xnor UO_3840 (O_3840,N_48837,N_49041);
or UO_3841 (O_3841,N_48338,N_48885);
xor UO_3842 (O_3842,N_48622,N_49116);
and UO_3843 (O_3843,N_49965,N_48254);
xor UO_3844 (O_3844,N_48528,N_48640);
xnor UO_3845 (O_3845,N_49869,N_48993);
and UO_3846 (O_3846,N_49761,N_49900);
and UO_3847 (O_3847,N_49348,N_48287);
nand UO_3848 (O_3848,N_48601,N_48740);
nand UO_3849 (O_3849,N_49700,N_49620);
nor UO_3850 (O_3850,N_48971,N_49136);
nor UO_3851 (O_3851,N_49364,N_48659);
and UO_3852 (O_3852,N_49215,N_48629);
and UO_3853 (O_3853,N_48478,N_48842);
nand UO_3854 (O_3854,N_48580,N_48292);
and UO_3855 (O_3855,N_49475,N_48717);
or UO_3856 (O_3856,N_49514,N_49540);
nand UO_3857 (O_3857,N_49436,N_48174);
xnor UO_3858 (O_3858,N_48844,N_48714);
or UO_3859 (O_3859,N_48720,N_49208);
nand UO_3860 (O_3860,N_49441,N_49116);
nand UO_3861 (O_3861,N_49166,N_48214);
xor UO_3862 (O_3862,N_48349,N_49142);
nor UO_3863 (O_3863,N_49885,N_49599);
xor UO_3864 (O_3864,N_49205,N_48743);
nand UO_3865 (O_3865,N_48443,N_48763);
and UO_3866 (O_3866,N_48077,N_48644);
or UO_3867 (O_3867,N_48557,N_49099);
and UO_3868 (O_3868,N_48373,N_49609);
xnor UO_3869 (O_3869,N_49481,N_48437);
or UO_3870 (O_3870,N_49972,N_48358);
and UO_3871 (O_3871,N_48816,N_48709);
nor UO_3872 (O_3872,N_49589,N_48625);
nand UO_3873 (O_3873,N_49546,N_48721);
xor UO_3874 (O_3874,N_49007,N_48684);
nand UO_3875 (O_3875,N_49701,N_49071);
nor UO_3876 (O_3876,N_48941,N_49391);
and UO_3877 (O_3877,N_48327,N_49714);
and UO_3878 (O_3878,N_49471,N_48614);
or UO_3879 (O_3879,N_49128,N_48796);
xor UO_3880 (O_3880,N_48500,N_48170);
nand UO_3881 (O_3881,N_49890,N_48720);
nor UO_3882 (O_3882,N_48526,N_49829);
or UO_3883 (O_3883,N_48540,N_49980);
nor UO_3884 (O_3884,N_48976,N_48567);
nor UO_3885 (O_3885,N_49294,N_49279);
nor UO_3886 (O_3886,N_48102,N_48862);
and UO_3887 (O_3887,N_48372,N_49859);
nand UO_3888 (O_3888,N_49907,N_48760);
and UO_3889 (O_3889,N_48789,N_48624);
and UO_3890 (O_3890,N_48379,N_49063);
xnor UO_3891 (O_3891,N_49108,N_48482);
and UO_3892 (O_3892,N_48264,N_48093);
and UO_3893 (O_3893,N_49905,N_49079);
or UO_3894 (O_3894,N_49302,N_48991);
xor UO_3895 (O_3895,N_48493,N_48596);
nand UO_3896 (O_3896,N_49413,N_48835);
xor UO_3897 (O_3897,N_48113,N_49106);
nand UO_3898 (O_3898,N_48037,N_48820);
and UO_3899 (O_3899,N_48095,N_49778);
nor UO_3900 (O_3900,N_49941,N_49573);
or UO_3901 (O_3901,N_49535,N_48567);
nand UO_3902 (O_3902,N_48623,N_49078);
nor UO_3903 (O_3903,N_48030,N_48099);
xor UO_3904 (O_3904,N_48297,N_49237);
nand UO_3905 (O_3905,N_48407,N_49078);
xor UO_3906 (O_3906,N_48115,N_48649);
nand UO_3907 (O_3907,N_48037,N_48986);
nand UO_3908 (O_3908,N_48589,N_48643);
nor UO_3909 (O_3909,N_49320,N_48895);
or UO_3910 (O_3910,N_49884,N_48057);
nor UO_3911 (O_3911,N_48673,N_49295);
xnor UO_3912 (O_3912,N_49722,N_49791);
nor UO_3913 (O_3913,N_48666,N_49735);
nand UO_3914 (O_3914,N_48593,N_48695);
xnor UO_3915 (O_3915,N_49626,N_48680);
nor UO_3916 (O_3916,N_48674,N_48511);
and UO_3917 (O_3917,N_48390,N_48391);
or UO_3918 (O_3918,N_49908,N_48742);
and UO_3919 (O_3919,N_48965,N_48415);
or UO_3920 (O_3920,N_49962,N_48042);
and UO_3921 (O_3921,N_49021,N_48007);
xor UO_3922 (O_3922,N_48289,N_48737);
nor UO_3923 (O_3923,N_48336,N_48505);
or UO_3924 (O_3924,N_48558,N_48391);
xor UO_3925 (O_3925,N_48079,N_49947);
or UO_3926 (O_3926,N_48038,N_49151);
nor UO_3927 (O_3927,N_48868,N_48900);
nand UO_3928 (O_3928,N_48649,N_49245);
nor UO_3929 (O_3929,N_48820,N_49341);
xnor UO_3930 (O_3930,N_48722,N_49202);
nor UO_3931 (O_3931,N_49387,N_48689);
nand UO_3932 (O_3932,N_48821,N_49537);
and UO_3933 (O_3933,N_49292,N_49975);
nand UO_3934 (O_3934,N_48867,N_49700);
nor UO_3935 (O_3935,N_48428,N_49107);
xnor UO_3936 (O_3936,N_49700,N_49831);
nor UO_3937 (O_3937,N_48694,N_49392);
nand UO_3938 (O_3938,N_49481,N_48028);
nor UO_3939 (O_3939,N_49575,N_48961);
nor UO_3940 (O_3940,N_48723,N_48468);
nand UO_3941 (O_3941,N_49752,N_49785);
nor UO_3942 (O_3942,N_48009,N_49870);
nand UO_3943 (O_3943,N_49195,N_49670);
nor UO_3944 (O_3944,N_48259,N_49860);
nand UO_3945 (O_3945,N_49523,N_48019);
and UO_3946 (O_3946,N_48568,N_49782);
xor UO_3947 (O_3947,N_48127,N_49899);
nor UO_3948 (O_3948,N_49568,N_49368);
xnor UO_3949 (O_3949,N_48382,N_48894);
or UO_3950 (O_3950,N_48840,N_49982);
nor UO_3951 (O_3951,N_49935,N_48383);
xnor UO_3952 (O_3952,N_48857,N_49203);
xnor UO_3953 (O_3953,N_48627,N_49428);
xor UO_3954 (O_3954,N_49825,N_48532);
xnor UO_3955 (O_3955,N_48701,N_49222);
xnor UO_3956 (O_3956,N_48316,N_49553);
nand UO_3957 (O_3957,N_49438,N_48312);
xor UO_3958 (O_3958,N_48023,N_49407);
xor UO_3959 (O_3959,N_48770,N_49195);
nand UO_3960 (O_3960,N_48964,N_48798);
nor UO_3961 (O_3961,N_48149,N_48028);
nor UO_3962 (O_3962,N_48240,N_49551);
nor UO_3963 (O_3963,N_49298,N_49119);
or UO_3964 (O_3964,N_48848,N_49098);
nand UO_3965 (O_3965,N_48017,N_49168);
and UO_3966 (O_3966,N_48928,N_48446);
nand UO_3967 (O_3967,N_49482,N_49736);
nand UO_3968 (O_3968,N_48463,N_48017);
nor UO_3969 (O_3969,N_49841,N_48539);
or UO_3970 (O_3970,N_48950,N_48298);
and UO_3971 (O_3971,N_49862,N_49473);
xnor UO_3972 (O_3972,N_49402,N_49427);
and UO_3973 (O_3973,N_48832,N_48737);
nand UO_3974 (O_3974,N_48469,N_48617);
xor UO_3975 (O_3975,N_49844,N_49151);
or UO_3976 (O_3976,N_49170,N_48493);
xor UO_3977 (O_3977,N_49858,N_48754);
nor UO_3978 (O_3978,N_49256,N_49088);
xnor UO_3979 (O_3979,N_48755,N_48144);
or UO_3980 (O_3980,N_49502,N_48770);
and UO_3981 (O_3981,N_48351,N_48387);
nand UO_3982 (O_3982,N_48084,N_49802);
or UO_3983 (O_3983,N_48382,N_49971);
nor UO_3984 (O_3984,N_48309,N_49873);
or UO_3985 (O_3985,N_49692,N_48044);
nand UO_3986 (O_3986,N_49453,N_48283);
nand UO_3987 (O_3987,N_49007,N_49414);
nand UO_3988 (O_3988,N_48150,N_49487);
xor UO_3989 (O_3989,N_48170,N_49325);
xnor UO_3990 (O_3990,N_48386,N_48975);
or UO_3991 (O_3991,N_49481,N_48076);
nor UO_3992 (O_3992,N_49473,N_49790);
nor UO_3993 (O_3993,N_48540,N_49761);
or UO_3994 (O_3994,N_48509,N_49338);
nor UO_3995 (O_3995,N_49726,N_48348);
and UO_3996 (O_3996,N_48242,N_48817);
nor UO_3997 (O_3997,N_48530,N_48362);
or UO_3998 (O_3998,N_49033,N_49178);
nand UO_3999 (O_3999,N_48592,N_49600);
or UO_4000 (O_4000,N_48143,N_49414);
xnor UO_4001 (O_4001,N_48747,N_49196);
or UO_4002 (O_4002,N_48960,N_49445);
nand UO_4003 (O_4003,N_49151,N_49467);
nor UO_4004 (O_4004,N_48970,N_48678);
nor UO_4005 (O_4005,N_48776,N_48887);
or UO_4006 (O_4006,N_48268,N_49754);
xor UO_4007 (O_4007,N_48915,N_49075);
nand UO_4008 (O_4008,N_48435,N_48260);
or UO_4009 (O_4009,N_49938,N_48847);
or UO_4010 (O_4010,N_49350,N_48098);
nor UO_4011 (O_4011,N_49528,N_48752);
nand UO_4012 (O_4012,N_49013,N_48015);
and UO_4013 (O_4013,N_49025,N_49382);
or UO_4014 (O_4014,N_49807,N_48394);
or UO_4015 (O_4015,N_48665,N_49674);
xnor UO_4016 (O_4016,N_49437,N_48336);
and UO_4017 (O_4017,N_48364,N_49702);
nand UO_4018 (O_4018,N_49525,N_49453);
xnor UO_4019 (O_4019,N_48010,N_48051);
nand UO_4020 (O_4020,N_48299,N_49895);
or UO_4021 (O_4021,N_48313,N_48767);
xnor UO_4022 (O_4022,N_49298,N_48703);
nor UO_4023 (O_4023,N_48090,N_49008);
and UO_4024 (O_4024,N_49838,N_48764);
nand UO_4025 (O_4025,N_49441,N_48915);
or UO_4026 (O_4026,N_48160,N_49656);
or UO_4027 (O_4027,N_49126,N_48202);
nor UO_4028 (O_4028,N_48292,N_49709);
nor UO_4029 (O_4029,N_49533,N_49068);
nand UO_4030 (O_4030,N_48089,N_49242);
nor UO_4031 (O_4031,N_48410,N_48541);
xor UO_4032 (O_4032,N_48637,N_48964);
and UO_4033 (O_4033,N_48699,N_48048);
nand UO_4034 (O_4034,N_49562,N_48793);
xor UO_4035 (O_4035,N_49879,N_49144);
xnor UO_4036 (O_4036,N_48664,N_49976);
or UO_4037 (O_4037,N_49781,N_48679);
and UO_4038 (O_4038,N_49997,N_49345);
nor UO_4039 (O_4039,N_48430,N_49115);
xor UO_4040 (O_4040,N_48995,N_48826);
xor UO_4041 (O_4041,N_49523,N_49126);
and UO_4042 (O_4042,N_48498,N_48893);
or UO_4043 (O_4043,N_48469,N_49669);
xor UO_4044 (O_4044,N_49709,N_49863);
nand UO_4045 (O_4045,N_49335,N_49908);
xnor UO_4046 (O_4046,N_48510,N_49410);
or UO_4047 (O_4047,N_49985,N_48311);
nor UO_4048 (O_4048,N_49580,N_48481);
or UO_4049 (O_4049,N_49626,N_49952);
and UO_4050 (O_4050,N_48439,N_49708);
and UO_4051 (O_4051,N_48465,N_49429);
or UO_4052 (O_4052,N_49339,N_48715);
and UO_4053 (O_4053,N_48785,N_48552);
nor UO_4054 (O_4054,N_48252,N_49330);
and UO_4055 (O_4055,N_49860,N_49706);
or UO_4056 (O_4056,N_49673,N_48032);
and UO_4057 (O_4057,N_49440,N_49918);
or UO_4058 (O_4058,N_49279,N_49385);
or UO_4059 (O_4059,N_49233,N_49922);
nand UO_4060 (O_4060,N_48104,N_48591);
or UO_4061 (O_4061,N_49630,N_48218);
and UO_4062 (O_4062,N_49279,N_48320);
nor UO_4063 (O_4063,N_48629,N_48376);
nand UO_4064 (O_4064,N_49219,N_48809);
nor UO_4065 (O_4065,N_49457,N_49292);
and UO_4066 (O_4066,N_48824,N_48723);
xor UO_4067 (O_4067,N_48827,N_49352);
xnor UO_4068 (O_4068,N_49377,N_49384);
nand UO_4069 (O_4069,N_48343,N_48969);
and UO_4070 (O_4070,N_48596,N_49770);
xor UO_4071 (O_4071,N_48723,N_49914);
xnor UO_4072 (O_4072,N_48350,N_48550);
xor UO_4073 (O_4073,N_48764,N_48907);
or UO_4074 (O_4074,N_49880,N_48746);
or UO_4075 (O_4075,N_49210,N_49649);
nor UO_4076 (O_4076,N_48345,N_49551);
xnor UO_4077 (O_4077,N_48761,N_49913);
or UO_4078 (O_4078,N_48720,N_48230);
and UO_4079 (O_4079,N_48304,N_48454);
xor UO_4080 (O_4080,N_49049,N_48279);
or UO_4081 (O_4081,N_48180,N_48361);
or UO_4082 (O_4082,N_48657,N_49775);
nor UO_4083 (O_4083,N_49452,N_49160);
or UO_4084 (O_4084,N_49119,N_49745);
and UO_4085 (O_4085,N_49043,N_48935);
xor UO_4086 (O_4086,N_48533,N_49234);
or UO_4087 (O_4087,N_48309,N_49180);
and UO_4088 (O_4088,N_48395,N_49190);
nor UO_4089 (O_4089,N_48645,N_49111);
and UO_4090 (O_4090,N_48007,N_49614);
or UO_4091 (O_4091,N_48153,N_49637);
nor UO_4092 (O_4092,N_48861,N_48918);
nand UO_4093 (O_4093,N_48494,N_49488);
nand UO_4094 (O_4094,N_48323,N_48531);
and UO_4095 (O_4095,N_49099,N_48381);
nor UO_4096 (O_4096,N_49538,N_48209);
or UO_4097 (O_4097,N_48186,N_49641);
and UO_4098 (O_4098,N_48039,N_48460);
nand UO_4099 (O_4099,N_49535,N_49854);
xor UO_4100 (O_4100,N_48010,N_48133);
nor UO_4101 (O_4101,N_48210,N_48287);
or UO_4102 (O_4102,N_48871,N_49104);
xnor UO_4103 (O_4103,N_48014,N_48858);
nand UO_4104 (O_4104,N_48908,N_48106);
nand UO_4105 (O_4105,N_48023,N_49054);
and UO_4106 (O_4106,N_49200,N_49464);
nand UO_4107 (O_4107,N_49013,N_49211);
and UO_4108 (O_4108,N_48756,N_48428);
xnor UO_4109 (O_4109,N_48236,N_48424);
xnor UO_4110 (O_4110,N_49435,N_49657);
or UO_4111 (O_4111,N_49359,N_49335);
and UO_4112 (O_4112,N_48143,N_48509);
xor UO_4113 (O_4113,N_49940,N_49509);
and UO_4114 (O_4114,N_49177,N_48180);
xor UO_4115 (O_4115,N_48165,N_48941);
or UO_4116 (O_4116,N_48855,N_49173);
or UO_4117 (O_4117,N_49140,N_48354);
nand UO_4118 (O_4118,N_48286,N_49147);
nor UO_4119 (O_4119,N_48827,N_49372);
xor UO_4120 (O_4120,N_48204,N_49561);
nand UO_4121 (O_4121,N_48482,N_48716);
or UO_4122 (O_4122,N_49982,N_49500);
nand UO_4123 (O_4123,N_48450,N_49984);
and UO_4124 (O_4124,N_48782,N_49336);
xor UO_4125 (O_4125,N_49098,N_49855);
nand UO_4126 (O_4126,N_49970,N_48739);
or UO_4127 (O_4127,N_48140,N_49858);
nor UO_4128 (O_4128,N_48586,N_49632);
nor UO_4129 (O_4129,N_48466,N_49775);
and UO_4130 (O_4130,N_49221,N_49300);
nor UO_4131 (O_4131,N_49924,N_49802);
nor UO_4132 (O_4132,N_48298,N_49996);
xnor UO_4133 (O_4133,N_48920,N_49783);
or UO_4134 (O_4134,N_48754,N_49076);
nand UO_4135 (O_4135,N_49037,N_49867);
xor UO_4136 (O_4136,N_48453,N_49507);
nand UO_4137 (O_4137,N_49967,N_48346);
nand UO_4138 (O_4138,N_49112,N_48931);
xor UO_4139 (O_4139,N_48148,N_49281);
xor UO_4140 (O_4140,N_49293,N_48155);
and UO_4141 (O_4141,N_48989,N_49938);
or UO_4142 (O_4142,N_48019,N_49900);
nand UO_4143 (O_4143,N_49416,N_48907);
and UO_4144 (O_4144,N_48737,N_49675);
nor UO_4145 (O_4145,N_49796,N_48163);
nand UO_4146 (O_4146,N_48769,N_49883);
and UO_4147 (O_4147,N_49221,N_49983);
nand UO_4148 (O_4148,N_49137,N_49491);
nand UO_4149 (O_4149,N_49219,N_48151);
or UO_4150 (O_4150,N_48887,N_48655);
and UO_4151 (O_4151,N_48647,N_49997);
nand UO_4152 (O_4152,N_48849,N_49829);
nor UO_4153 (O_4153,N_48874,N_48528);
xor UO_4154 (O_4154,N_48889,N_48075);
xor UO_4155 (O_4155,N_48213,N_48786);
nor UO_4156 (O_4156,N_48069,N_49002);
xnor UO_4157 (O_4157,N_48669,N_48146);
nand UO_4158 (O_4158,N_48103,N_49557);
and UO_4159 (O_4159,N_48991,N_48931);
xnor UO_4160 (O_4160,N_48060,N_48003);
and UO_4161 (O_4161,N_48394,N_48764);
xor UO_4162 (O_4162,N_48351,N_48235);
nor UO_4163 (O_4163,N_49844,N_49373);
nand UO_4164 (O_4164,N_48212,N_48625);
xnor UO_4165 (O_4165,N_49756,N_49380);
and UO_4166 (O_4166,N_48392,N_48796);
nor UO_4167 (O_4167,N_49268,N_49270);
or UO_4168 (O_4168,N_48647,N_48707);
xnor UO_4169 (O_4169,N_48519,N_48824);
nand UO_4170 (O_4170,N_48771,N_48110);
nor UO_4171 (O_4171,N_49727,N_49564);
or UO_4172 (O_4172,N_48150,N_48923);
nand UO_4173 (O_4173,N_48769,N_49079);
or UO_4174 (O_4174,N_48672,N_48021);
nand UO_4175 (O_4175,N_48810,N_49714);
or UO_4176 (O_4176,N_48979,N_49215);
nor UO_4177 (O_4177,N_49840,N_48331);
nor UO_4178 (O_4178,N_48023,N_49408);
or UO_4179 (O_4179,N_48475,N_48159);
nand UO_4180 (O_4180,N_49414,N_48526);
xnor UO_4181 (O_4181,N_48381,N_49487);
nor UO_4182 (O_4182,N_49585,N_48310);
nand UO_4183 (O_4183,N_48214,N_49077);
or UO_4184 (O_4184,N_49874,N_48024);
xnor UO_4185 (O_4185,N_48111,N_48760);
or UO_4186 (O_4186,N_48885,N_49802);
and UO_4187 (O_4187,N_48334,N_48500);
or UO_4188 (O_4188,N_49136,N_49617);
nor UO_4189 (O_4189,N_48687,N_49447);
nor UO_4190 (O_4190,N_48962,N_49565);
and UO_4191 (O_4191,N_48961,N_48126);
and UO_4192 (O_4192,N_48326,N_49730);
xnor UO_4193 (O_4193,N_48455,N_49426);
nand UO_4194 (O_4194,N_48498,N_48396);
nor UO_4195 (O_4195,N_49117,N_49061);
or UO_4196 (O_4196,N_49299,N_48282);
nand UO_4197 (O_4197,N_48520,N_48334);
or UO_4198 (O_4198,N_49107,N_48710);
nor UO_4199 (O_4199,N_49443,N_49685);
or UO_4200 (O_4200,N_48472,N_49796);
nor UO_4201 (O_4201,N_49890,N_49587);
xor UO_4202 (O_4202,N_48791,N_48129);
and UO_4203 (O_4203,N_48379,N_49839);
and UO_4204 (O_4204,N_48108,N_48065);
xnor UO_4205 (O_4205,N_49162,N_48360);
and UO_4206 (O_4206,N_49248,N_49461);
xnor UO_4207 (O_4207,N_48340,N_49618);
nor UO_4208 (O_4208,N_48435,N_49601);
xor UO_4209 (O_4209,N_48057,N_48180);
and UO_4210 (O_4210,N_48318,N_49212);
nor UO_4211 (O_4211,N_48769,N_49757);
and UO_4212 (O_4212,N_48645,N_48354);
or UO_4213 (O_4213,N_49701,N_48046);
xor UO_4214 (O_4214,N_49052,N_49966);
xor UO_4215 (O_4215,N_49949,N_48163);
nor UO_4216 (O_4216,N_48646,N_48007);
or UO_4217 (O_4217,N_48119,N_48632);
xor UO_4218 (O_4218,N_49746,N_48456);
and UO_4219 (O_4219,N_49361,N_48450);
or UO_4220 (O_4220,N_49289,N_48403);
nand UO_4221 (O_4221,N_48060,N_49267);
or UO_4222 (O_4222,N_48629,N_48691);
and UO_4223 (O_4223,N_48383,N_49668);
xnor UO_4224 (O_4224,N_49132,N_49678);
or UO_4225 (O_4225,N_48243,N_49438);
or UO_4226 (O_4226,N_49915,N_48361);
nor UO_4227 (O_4227,N_49403,N_49845);
nor UO_4228 (O_4228,N_49652,N_48354);
and UO_4229 (O_4229,N_49762,N_48391);
nand UO_4230 (O_4230,N_48803,N_49455);
or UO_4231 (O_4231,N_49428,N_48682);
nor UO_4232 (O_4232,N_48850,N_49692);
and UO_4233 (O_4233,N_48131,N_49452);
nand UO_4234 (O_4234,N_48325,N_48326);
nor UO_4235 (O_4235,N_49986,N_49075);
nor UO_4236 (O_4236,N_49906,N_49993);
and UO_4237 (O_4237,N_49900,N_49602);
or UO_4238 (O_4238,N_48388,N_49534);
xnor UO_4239 (O_4239,N_48075,N_48029);
nand UO_4240 (O_4240,N_48421,N_48653);
or UO_4241 (O_4241,N_48029,N_49696);
xnor UO_4242 (O_4242,N_48037,N_48018);
xor UO_4243 (O_4243,N_48851,N_48031);
and UO_4244 (O_4244,N_48039,N_49604);
nor UO_4245 (O_4245,N_49331,N_48418);
nor UO_4246 (O_4246,N_49432,N_49403);
or UO_4247 (O_4247,N_49311,N_49401);
xnor UO_4248 (O_4248,N_49863,N_48202);
nor UO_4249 (O_4249,N_48671,N_49537);
nand UO_4250 (O_4250,N_49697,N_48897);
and UO_4251 (O_4251,N_48311,N_48044);
nand UO_4252 (O_4252,N_49872,N_49308);
and UO_4253 (O_4253,N_48987,N_49381);
xnor UO_4254 (O_4254,N_48280,N_49618);
nand UO_4255 (O_4255,N_49474,N_49863);
and UO_4256 (O_4256,N_49611,N_48507);
nor UO_4257 (O_4257,N_49912,N_49984);
or UO_4258 (O_4258,N_49020,N_48891);
nor UO_4259 (O_4259,N_48532,N_49981);
and UO_4260 (O_4260,N_49808,N_48796);
nor UO_4261 (O_4261,N_49966,N_48796);
nor UO_4262 (O_4262,N_49469,N_48514);
or UO_4263 (O_4263,N_49244,N_48662);
nor UO_4264 (O_4264,N_49455,N_48007);
and UO_4265 (O_4265,N_49192,N_48710);
nor UO_4266 (O_4266,N_48470,N_48376);
nor UO_4267 (O_4267,N_49576,N_48862);
and UO_4268 (O_4268,N_49471,N_49895);
xor UO_4269 (O_4269,N_49573,N_48848);
nand UO_4270 (O_4270,N_49992,N_48964);
nand UO_4271 (O_4271,N_48488,N_49796);
nor UO_4272 (O_4272,N_48215,N_49143);
nor UO_4273 (O_4273,N_49497,N_49298);
or UO_4274 (O_4274,N_48078,N_48349);
or UO_4275 (O_4275,N_48455,N_49367);
or UO_4276 (O_4276,N_48286,N_49966);
or UO_4277 (O_4277,N_49113,N_49205);
nor UO_4278 (O_4278,N_49890,N_48968);
nand UO_4279 (O_4279,N_49522,N_48414);
xor UO_4280 (O_4280,N_49210,N_48688);
and UO_4281 (O_4281,N_48201,N_48932);
nand UO_4282 (O_4282,N_49343,N_49022);
nand UO_4283 (O_4283,N_48319,N_49284);
nor UO_4284 (O_4284,N_48542,N_49081);
xor UO_4285 (O_4285,N_48181,N_49807);
nand UO_4286 (O_4286,N_48227,N_49552);
or UO_4287 (O_4287,N_48675,N_48884);
nand UO_4288 (O_4288,N_49274,N_49968);
and UO_4289 (O_4289,N_49147,N_49721);
and UO_4290 (O_4290,N_48315,N_48885);
or UO_4291 (O_4291,N_49379,N_49524);
nand UO_4292 (O_4292,N_48807,N_49814);
and UO_4293 (O_4293,N_48628,N_48994);
nor UO_4294 (O_4294,N_48092,N_49412);
and UO_4295 (O_4295,N_49683,N_49784);
and UO_4296 (O_4296,N_48089,N_49511);
or UO_4297 (O_4297,N_49605,N_48221);
or UO_4298 (O_4298,N_48302,N_49394);
nand UO_4299 (O_4299,N_48304,N_49603);
or UO_4300 (O_4300,N_48447,N_49462);
nor UO_4301 (O_4301,N_49942,N_49950);
and UO_4302 (O_4302,N_49948,N_49145);
or UO_4303 (O_4303,N_49019,N_49615);
xor UO_4304 (O_4304,N_48163,N_49520);
nor UO_4305 (O_4305,N_48211,N_48993);
or UO_4306 (O_4306,N_49764,N_49790);
and UO_4307 (O_4307,N_49717,N_49585);
nor UO_4308 (O_4308,N_49941,N_49727);
xnor UO_4309 (O_4309,N_48095,N_49091);
and UO_4310 (O_4310,N_48053,N_48957);
nand UO_4311 (O_4311,N_48848,N_49195);
or UO_4312 (O_4312,N_49232,N_49262);
nand UO_4313 (O_4313,N_48859,N_49260);
xnor UO_4314 (O_4314,N_49918,N_49172);
xor UO_4315 (O_4315,N_48654,N_48248);
xor UO_4316 (O_4316,N_48099,N_49323);
nor UO_4317 (O_4317,N_49871,N_49401);
or UO_4318 (O_4318,N_48718,N_48123);
nor UO_4319 (O_4319,N_49391,N_48510);
nand UO_4320 (O_4320,N_49345,N_48182);
and UO_4321 (O_4321,N_48014,N_49415);
or UO_4322 (O_4322,N_49297,N_48080);
nor UO_4323 (O_4323,N_49884,N_48004);
nor UO_4324 (O_4324,N_49619,N_49391);
or UO_4325 (O_4325,N_49274,N_49066);
or UO_4326 (O_4326,N_49564,N_48217);
xnor UO_4327 (O_4327,N_49984,N_48841);
and UO_4328 (O_4328,N_48222,N_48151);
and UO_4329 (O_4329,N_48662,N_48978);
and UO_4330 (O_4330,N_48799,N_49631);
or UO_4331 (O_4331,N_49449,N_49533);
nand UO_4332 (O_4332,N_48740,N_48145);
nor UO_4333 (O_4333,N_49227,N_49403);
nand UO_4334 (O_4334,N_49295,N_48804);
xor UO_4335 (O_4335,N_49846,N_49614);
and UO_4336 (O_4336,N_48758,N_49643);
nor UO_4337 (O_4337,N_48997,N_48574);
or UO_4338 (O_4338,N_49745,N_49985);
nand UO_4339 (O_4339,N_48675,N_48927);
nand UO_4340 (O_4340,N_48908,N_49711);
or UO_4341 (O_4341,N_49027,N_49449);
nand UO_4342 (O_4342,N_49648,N_48209);
and UO_4343 (O_4343,N_49951,N_49834);
xnor UO_4344 (O_4344,N_48879,N_48296);
xnor UO_4345 (O_4345,N_49802,N_49678);
nand UO_4346 (O_4346,N_48138,N_49319);
and UO_4347 (O_4347,N_49688,N_49444);
and UO_4348 (O_4348,N_49702,N_48579);
nand UO_4349 (O_4349,N_48931,N_49459);
or UO_4350 (O_4350,N_49804,N_48086);
nor UO_4351 (O_4351,N_49572,N_49840);
nor UO_4352 (O_4352,N_48984,N_49174);
xor UO_4353 (O_4353,N_49207,N_49107);
or UO_4354 (O_4354,N_49435,N_48575);
nor UO_4355 (O_4355,N_48539,N_49147);
and UO_4356 (O_4356,N_49502,N_48542);
nand UO_4357 (O_4357,N_48037,N_49568);
nor UO_4358 (O_4358,N_49541,N_48318);
nand UO_4359 (O_4359,N_48970,N_48504);
or UO_4360 (O_4360,N_48860,N_48291);
nand UO_4361 (O_4361,N_48655,N_48298);
xor UO_4362 (O_4362,N_49814,N_48671);
nor UO_4363 (O_4363,N_49399,N_48816);
nor UO_4364 (O_4364,N_49469,N_48081);
nand UO_4365 (O_4365,N_48232,N_49249);
nor UO_4366 (O_4366,N_48634,N_48503);
nand UO_4367 (O_4367,N_49241,N_48170);
and UO_4368 (O_4368,N_49888,N_49650);
nor UO_4369 (O_4369,N_48310,N_48552);
and UO_4370 (O_4370,N_49200,N_49563);
and UO_4371 (O_4371,N_49453,N_48389);
and UO_4372 (O_4372,N_49069,N_49425);
or UO_4373 (O_4373,N_49055,N_48497);
nand UO_4374 (O_4374,N_49539,N_48522);
xor UO_4375 (O_4375,N_48109,N_48714);
xnor UO_4376 (O_4376,N_48380,N_48274);
xnor UO_4377 (O_4377,N_49783,N_48242);
or UO_4378 (O_4378,N_49133,N_48064);
xor UO_4379 (O_4379,N_48601,N_48609);
or UO_4380 (O_4380,N_48672,N_49732);
nor UO_4381 (O_4381,N_48248,N_48880);
nand UO_4382 (O_4382,N_48575,N_48718);
or UO_4383 (O_4383,N_48094,N_49523);
nand UO_4384 (O_4384,N_48140,N_49754);
and UO_4385 (O_4385,N_49237,N_49808);
xor UO_4386 (O_4386,N_48844,N_48875);
xor UO_4387 (O_4387,N_48580,N_49320);
or UO_4388 (O_4388,N_49367,N_49492);
nand UO_4389 (O_4389,N_49755,N_48033);
and UO_4390 (O_4390,N_48101,N_49816);
and UO_4391 (O_4391,N_49595,N_49020);
or UO_4392 (O_4392,N_48314,N_49887);
or UO_4393 (O_4393,N_48298,N_49866);
or UO_4394 (O_4394,N_48489,N_48403);
xnor UO_4395 (O_4395,N_48213,N_49954);
nor UO_4396 (O_4396,N_48735,N_49372);
and UO_4397 (O_4397,N_49460,N_48208);
and UO_4398 (O_4398,N_49404,N_48969);
and UO_4399 (O_4399,N_48175,N_48432);
nor UO_4400 (O_4400,N_48203,N_49429);
nand UO_4401 (O_4401,N_48412,N_48915);
nor UO_4402 (O_4402,N_48351,N_49694);
and UO_4403 (O_4403,N_48215,N_49706);
and UO_4404 (O_4404,N_48296,N_49344);
or UO_4405 (O_4405,N_49600,N_48258);
nand UO_4406 (O_4406,N_48184,N_49394);
and UO_4407 (O_4407,N_48607,N_49908);
nand UO_4408 (O_4408,N_49145,N_49058);
xor UO_4409 (O_4409,N_48847,N_49555);
nand UO_4410 (O_4410,N_48221,N_49530);
xnor UO_4411 (O_4411,N_48029,N_48716);
and UO_4412 (O_4412,N_49679,N_48137);
nor UO_4413 (O_4413,N_48844,N_48113);
or UO_4414 (O_4414,N_48543,N_49421);
xor UO_4415 (O_4415,N_49435,N_48039);
or UO_4416 (O_4416,N_48503,N_48103);
nand UO_4417 (O_4417,N_49079,N_48331);
and UO_4418 (O_4418,N_49424,N_48524);
xnor UO_4419 (O_4419,N_49250,N_49070);
or UO_4420 (O_4420,N_48697,N_49210);
and UO_4421 (O_4421,N_48722,N_49499);
nand UO_4422 (O_4422,N_49225,N_48034);
nor UO_4423 (O_4423,N_49217,N_48049);
and UO_4424 (O_4424,N_49365,N_48949);
nand UO_4425 (O_4425,N_48765,N_49263);
xnor UO_4426 (O_4426,N_49827,N_49952);
xnor UO_4427 (O_4427,N_48845,N_48856);
and UO_4428 (O_4428,N_49483,N_48697);
nand UO_4429 (O_4429,N_49147,N_49890);
nor UO_4430 (O_4430,N_49579,N_49343);
or UO_4431 (O_4431,N_49642,N_49001);
xnor UO_4432 (O_4432,N_49545,N_48785);
xnor UO_4433 (O_4433,N_48035,N_48991);
xnor UO_4434 (O_4434,N_48285,N_48673);
xor UO_4435 (O_4435,N_48452,N_48546);
nand UO_4436 (O_4436,N_49275,N_49669);
xnor UO_4437 (O_4437,N_49824,N_49979);
nor UO_4438 (O_4438,N_48968,N_49755);
and UO_4439 (O_4439,N_49348,N_49017);
nor UO_4440 (O_4440,N_49030,N_49964);
xor UO_4441 (O_4441,N_49927,N_49849);
xnor UO_4442 (O_4442,N_49697,N_49296);
xnor UO_4443 (O_4443,N_49569,N_48878);
and UO_4444 (O_4444,N_48521,N_49390);
nand UO_4445 (O_4445,N_49056,N_49071);
nor UO_4446 (O_4446,N_48300,N_49130);
nand UO_4447 (O_4447,N_48853,N_48588);
nand UO_4448 (O_4448,N_48175,N_48627);
nand UO_4449 (O_4449,N_49552,N_49040);
xor UO_4450 (O_4450,N_48675,N_48465);
xor UO_4451 (O_4451,N_48023,N_49213);
or UO_4452 (O_4452,N_48707,N_49019);
and UO_4453 (O_4453,N_48343,N_49447);
nor UO_4454 (O_4454,N_48421,N_48685);
nand UO_4455 (O_4455,N_48206,N_49362);
or UO_4456 (O_4456,N_48094,N_48798);
or UO_4457 (O_4457,N_49870,N_48576);
nand UO_4458 (O_4458,N_49986,N_49431);
xor UO_4459 (O_4459,N_49390,N_49750);
or UO_4460 (O_4460,N_48835,N_48003);
nor UO_4461 (O_4461,N_49089,N_49913);
nand UO_4462 (O_4462,N_48444,N_49993);
and UO_4463 (O_4463,N_49190,N_49450);
or UO_4464 (O_4464,N_49101,N_48294);
xor UO_4465 (O_4465,N_48426,N_48591);
or UO_4466 (O_4466,N_49923,N_48303);
and UO_4467 (O_4467,N_48450,N_48483);
or UO_4468 (O_4468,N_48924,N_48762);
nand UO_4469 (O_4469,N_49811,N_48557);
or UO_4470 (O_4470,N_49899,N_48275);
xnor UO_4471 (O_4471,N_48598,N_48771);
xor UO_4472 (O_4472,N_48638,N_48911);
xor UO_4473 (O_4473,N_48517,N_49088);
nor UO_4474 (O_4474,N_49530,N_48434);
xor UO_4475 (O_4475,N_49073,N_49999);
nor UO_4476 (O_4476,N_48835,N_49638);
and UO_4477 (O_4477,N_48289,N_48319);
xor UO_4478 (O_4478,N_49863,N_48424);
and UO_4479 (O_4479,N_48560,N_49569);
or UO_4480 (O_4480,N_49364,N_49092);
nand UO_4481 (O_4481,N_49174,N_49323);
nor UO_4482 (O_4482,N_48303,N_49085);
nand UO_4483 (O_4483,N_48690,N_49450);
and UO_4484 (O_4484,N_49581,N_48666);
nand UO_4485 (O_4485,N_49707,N_48828);
nor UO_4486 (O_4486,N_48499,N_48858);
xnor UO_4487 (O_4487,N_49567,N_48180);
or UO_4488 (O_4488,N_49008,N_49707);
or UO_4489 (O_4489,N_49366,N_49951);
nor UO_4490 (O_4490,N_48375,N_49062);
nor UO_4491 (O_4491,N_49401,N_48729);
and UO_4492 (O_4492,N_49476,N_48299);
nor UO_4493 (O_4493,N_48657,N_48231);
or UO_4494 (O_4494,N_49386,N_48233);
nor UO_4495 (O_4495,N_48759,N_49215);
nand UO_4496 (O_4496,N_49358,N_48853);
and UO_4497 (O_4497,N_48394,N_48513);
nand UO_4498 (O_4498,N_48059,N_48761);
or UO_4499 (O_4499,N_49695,N_48184);
or UO_4500 (O_4500,N_48462,N_49307);
nor UO_4501 (O_4501,N_49915,N_49234);
nor UO_4502 (O_4502,N_49851,N_48597);
and UO_4503 (O_4503,N_49384,N_49311);
xor UO_4504 (O_4504,N_49375,N_48055);
and UO_4505 (O_4505,N_49157,N_49769);
and UO_4506 (O_4506,N_49289,N_48043);
or UO_4507 (O_4507,N_49282,N_49742);
nand UO_4508 (O_4508,N_48590,N_49005);
nand UO_4509 (O_4509,N_48345,N_49711);
nor UO_4510 (O_4510,N_48072,N_48710);
and UO_4511 (O_4511,N_49047,N_48576);
xor UO_4512 (O_4512,N_49553,N_49296);
nor UO_4513 (O_4513,N_49263,N_49199);
nand UO_4514 (O_4514,N_49153,N_49105);
nand UO_4515 (O_4515,N_48483,N_49816);
nor UO_4516 (O_4516,N_48345,N_48456);
and UO_4517 (O_4517,N_49965,N_48290);
and UO_4518 (O_4518,N_49830,N_48779);
or UO_4519 (O_4519,N_48514,N_49970);
nand UO_4520 (O_4520,N_49335,N_49240);
nand UO_4521 (O_4521,N_48496,N_49590);
or UO_4522 (O_4522,N_49476,N_48775);
xor UO_4523 (O_4523,N_49453,N_48860);
or UO_4524 (O_4524,N_49482,N_48606);
and UO_4525 (O_4525,N_49101,N_48923);
xnor UO_4526 (O_4526,N_48605,N_48574);
and UO_4527 (O_4527,N_49278,N_49429);
nor UO_4528 (O_4528,N_48057,N_49569);
nand UO_4529 (O_4529,N_49938,N_48421);
nand UO_4530 (O_4530,N_49362,N_48787);
or UO_4531 (O_4531,N_48142,N_48481);
nand UO_4532 (O_4532,N_48302,N_48083);
nand UO_4533 (O_4533,N_49422,N_48884);
xnor UO_4534 (O_4534,N_49399,N_48377);
and UO_4535 (O_4535,N_49098,N_49353);
nand UO_4536 (O_4536,N_48478,N_48962);
nor UO_4537 (O_4537,N_48789,N_49717);
and UO_4538 (O_4538,N_49722,N_48399);
and UO_4539 (O_4539,N_49147,N_49801);
nor UO_4540 (O_4540,N_49154,N_49683);
nor UO_4541 (O_4541,N_48391,N_49688);
nor UO_4542 (O_4542,N_48073,N_49037);
nand UO_4543 (O_4543,N_48405,N_49303);
xnor UO_4544 (O_4544,N_49995,N_49594);
nor UO_4545 (O_4545,N_49057,N_48242);
xor UO_4546 (O_4546,N_49748,N_49808);
or UO_4547 (O_4547,N_49017,N_49809);
and UO_4548 (O_4548,N_49285,N_49979);
and UO_4549 (O_4549,N_49627,N_49188);
nand UO_4550 (O_4550,N_48430,N_48111);
and UO_4551 (O_4551,N_49310,N_49541);
or UO_4552 (O_4552,N_48728,N_49310);
nand UO_4553 (O_4553,N_48002,N_48009);
nor UO_4554 (O_4554,N_48456,N_48524);
nor UO_4555 (O_4555,N_49337,N_48337);
and UO_4556 (O_4556,N_49504,N_48590);
and UO_4557 (O_4557,N_48270,N_48116);
or UO_4558 (O_4558,N_48359,N_49345);
and UO_4559 (O_4559,N_48579,N_48599);
or UO_4560 (O_4560,N_48413,N_49515);
and UO_4561 (O_4561,N_49885,N_48880);
nand UO_4562 (O_4562,N_49488,N_49941);
nor UO_4563 (O_4563,N_48777,N_49999);
or UO_4564 (O_4564,N_48083,N_49206);
nand UO_4565 (O_4565,N_49386,N_48654);
nand UO_4566 (O_4566,N_49915,N_48366);
xnor UO_4567 (O_4567,N_48665,N_48138);
nor UO_4568 (O_4568,N_49315,N_48430);
and UO_4569 (O_4569,N_48635,N_48035);
or UO_4570 (O_4570,N_49628,N_49658);
xor UO_4571 (O_4571,N_49451,N_48595);
and UO_4572 (O_4572,N_49686,N_49747);
and UO_4573 (O_4573,N_49172,N_49550);
or UO_4574 (O_4574,N_48950,N_49114);
xor UO_4575 (O_4575,N_49804,N_49036);
xnor UO_4576 (O_4576,N_48359,N_49075);
or UO_4577 (O_4577,N_48657,N_49939);
nor UO_4578 (O_4578,N_48960,N_49835);
or UO_4579 (O_4579,N_48567,N_49442);
or UO_4580 (O_4580,N_48519,N_48077);
nand UO_4581 (O_4581,N_49816,N_48779);
nand UO_4582 (O_4582,N_48246,N_48358);
nor UO_4583 (O_4583,N_48503,N_48337);
or UO_4584 (O_4584,N_48089,N_48633);
nand UO_4585 (O_4585,N_49924,N_49801);
nor UO_4586 (O_4586,N_49558,N_48818);
and UO_4587 (O_4587,N_48305,N_49076);
nand UO_4588 (O_4588,N_49496,N_49517);
xor UO_4589 (O_4589,N_49699,N_48109);
nor UO_4590 (O_4590,N_48901,N_49122);
xor UO_4591 (O_4591,N_48391,N_49527);
or UO_4592 (O_4592,N_49545,N_49440);
or UO_4593 (O_4593,N_48345,N_48683);
xnor UO_4594 (O_4594,N_49957,N_48388);
xor UO_4595 (O_4595,N_49298,N_48150);
or UO_4596 (O_4596,N_49244,N_49167);
nor UO_4597 (O_4597,N_49023,N_49189);
and UO_4598 (O_4598,N_48432,N_49511);
nand UO_4599 (O_4599,N_49540,N_49914);
nor UO_4600 (O_4600,N_48595,N_48669);
and UO_4601 (O_4601,N_48724,N_48258);
and UO_4602 (O_4602,N_49022,N_48734);
and UO_4603 (O_4603,N_49529,N_48096);
or UO_4604 (O_4604,N_48517,N_49520);
and UO_4605 (O_4605,N_48551,N_48975);
nand UO_4606 (O_4606,N_49050,N_48685);
nor UO_4607 (O_4607,N_48106,N_49715);
nand UO_4608 (O_4608,N_48155,N_49430);
and UO_4609 (O_4609,N_49321,N_49628);
nor UO_4610 (O_4610,N_49629,N_49945);
xor UO_4611 (O_4611,N_49219,N_49690);
xor UO_4612 (O_4612,N_49678,N_48217);
nand UO_4613 (O_4613,N_48285,N_48031);
nand UO_4614 (O_4614,N_49149,N_49033);
nor UO_4615 (O_4615,N_49553,N_49473);
nand UO_4616 (O_4616,N_48116,N_49647);
xnor UO_4617 (O_4617,N_49396,N_48912);
nand UO_4618 (O_4618,N_48907,N_49328);
nand UO_4619 (O_4619,N_48406,N_48679);
and UO_4620 (O_4620,N_48880,N_49308);
and UO_4621 (O_4621,N_48308,N_49791);
and UO_4622 (O_4622,N_48538,N_49364);
and UO_4623 (O_4623,N_49832,N_48729);
nand UO_4624 (O_4624,N_49639,N_48784);
nor UO_4625 (O_4625,N_48703,N_48138);
or UO_4626 (O_4626,N_49526,N_49123);
and UO_4627 (O_4627,N_48030,N_48785);
and UO_4628 (O_4628,N_48046,N_49256);
nor UO_4629 (O_4629,N_49381,N_49973);
nor UO_4630 (O_4630,N_49787,N_48505);
nor UO_4631 (O_4631,N_48179,N_48615);
xnor UO_4632 (O_4632,N_49705,N_48994);
nand UO_4633 (O_4633,N_48623,N_49629);
nand UO_4634 (O_4634,N_48491,N_49293);
or UO_4635 (O_4635,N_48851,N_49856);
nand UO_4636 (O_4636,N_49567,N_49850);
or UO_4637 (O_4637,N_48363,N_48714);
and UO_4638 (O_4638,N_48785,N_49993);
nand UO_4639 (O_4639,N_48748,N_48357);
or UO_4640 (O_4640,N_48262,N_48071);
xnor UO_4641 (O_4641,N_49151,N_49367);
nor UO_4642 (O_4642,N_48941,N_49927);
nand UO_4643 (O_4643,N_48280,N_49102);
nor UO_4644 (O_4644,N_49230,N_49794);
and UO_4645 (O_4645,N_48091,N_49683);
xnor UO_4646 (O_4646,N_48332,N_48126);
nor UO_4647 (O_4647,N_49649,N_49677);
xnor UO_4648 (O_4648,N_48369,N_49954);
nor UO_4649 (O_4649,N_49000,N_49543);
xnor UO_4650 (O_4650,N_49782,N_48527);
nand UO_4651 (O_4651,N_49856,N_49104);
xor UO_4652 (O_4652,N_48991,N_48144);
or UO_4653 (O_4653,N_48658,N_49261);
nor UO_4654 (O_4654,N_49911,N_49722);
and UO_4655 (O_4655,N_49686,N_49991);
or UO_4656 (O_4656,N_49291,N_49951);
and UO_4657 (O_4657,N_48986,N_48346);
nor UO_4658 (O_4658,N_49489,N_49134);
nor UO_4659 (O_4659,N_49214,N_49027);
xor UO_4660 (O_4660,N_49380,N_49178);
nor UO_4661 (O_4661,N_48179,N_48351);
xor UO_4662 (O_4662,N_48914,N_48095);
xor UO_4663 (O_4663,N_49669,N_49981);
and UO_4664 (O_4664,N_49544,N_49771);
and UO_4665 (O_4665,N_48456,N_48131);
and UO_4666 (O_4666,N_49626,N_48327);
or UO_4667 (O_4667,N_48024,N_48337);
xnor UO_4668 (O_4668,N_49895,N_48654);
xnor UO_4669 (O_4669,N_48427,N_48654);
xor UO_4670 (O_4670,N_48273,N_48378);
nor UO_4671 (O_4671,N_48283,N_49939);
nor UO_4672 (O_4672,N_49182,N_49699);
xor UO_4673 (O_4673,N_48250,N_49422);
or UO_4674 (O_4674,N_49731,N_49423);
nand UO_4675 (O_4675,N_49148,N_49851);
and UO_4676 (O_4676,N_48791,N_49573);
and UO_4677 (O_4677,N_49405,N_49453);
or UO_4678 (O_4678,N_48478,N_48469);
nand UO_4679 (O_4679,N_48327,N_49824);
xnor UO_4680 (O_4680,N_49830,N_48611);
nand UO_4681 (O_4681,N_48101,N_49988);
and UO_4682 (O_4682,N_49636,N_49386);
nor UO_4683 (O_4683,N_49931,N_48920);
nor UO_4684 (O_4684,N_48204,N_48286);
nand UO_4685 (O_4685,N_49199,N_48399);
and UO_4686 (O_4686,N_49843,N_48226);
xnor UO_4687 (O_4687,N_48919,N_49502);
xor UO_4688 (O_4688,N_48039,N_49409);
xnor UO_4689 (O_4689,N_49877,N_49021);
nand UO_4690 (O_4690,N_49180,N_49187);
nand UO_4691 (O_4691,N_49445,N_48987);
nor UO_4692 (O_4692,N_49885,N_49221);
xor UO_4693 (O_4693,N_49329,N_49914);
or UO_4694 (O_4694,N_49990,N_49012);
or UO_4695 (O_4695,N_49020,N_48093);
nand UO_4696 (O_4696,N_49368,N_48864);
and UO_4697 (O_4697,N_49693,N_48655);
xnor UO_4698 (O_4698,N_49647,N_48728);
xor UO_4699 (O_4699,N_48767,N_49895);
xnor UO_4700 (O_4700,N_48239,N_49840);
nand UO_4701 (O_4701,N_48541,N_48353);
and UO_4702 (O_4702,N_49584,N_49172);
xnor UO_4703 (O_4703,N_48438,N_48716);
or UO_4704 (O_4704,N_49951,N_49187);
or UO_4705 (O_4705,N_49653,N_48075);
and UO_4706 (O_4706,N_48507,N_49213);
xor UO_4707 (O_4707,N_49136,N_48461);
nor UO_4708 (O_4708,N_49713,N_48975);
nor UO_4709 (O_4709,N_48784,N_48175);
nand UO_4710 (O_4710,N_49174,N_49875);
xor UO_4711 (O_4711,N_49066,N_48654);
and UO_4712 (O_4712,N_49406,N_48584);
or UO_4713 (O_4713,N_48339,N_48844);
nor UO_4714 (O_4714,N_48364,N_49505);
nor UO_4715 (O_4715,N_48701,N_49736);
or UO_4716 (O_4716,N_48234,N_48833);
xor UO_4717 (O_4717,N_48264,N_49545);
nor UO_4718 (O_4718,N_48279,N_49236);
nor UO_4719 (O_4719,N_49659,N_48285);
nor UO_4720 (O_4720,N_49885,N_48257);
xor UO_4721 (O_4721,N_48701,N_49720);
and UO_4722 (O_4722,N_49369,N_48350);
and UO_4723 (O_4723,N_49904,N_49345);
or UO_4724 (O_4724,N_48195,N_49971);
xor UO_4725 (O_4725,N_49652,N_48892);
or UO_4726 (O_4726,N_48545,N_48649);
nand UO_4727 (O_4727,N_48158,N_49873);
or UO_4728 (O_4728,N_48290,N_48066);
and UO_4729 (O_4729,N_49610,N_49592);
and UO_4730 (O_4730,N_49101,N_49362);
nand UO_4731 (O_4731,N_49624,N_49571);
nand UO_4732 (O_4732,N_49963,N_48503);
nand UO_4733 (O_4733,N_49887,N_49967);
nor UO_4734 (O_4734,N_49732,N_49705);
nor UO_4735 (O_4735,N_48617,N_48475);
and UO_4736 (O_4736,N_48078,N_49554);
nor UO_4737 (O_4737,N_49311,N_49014);
nor UO_4738 (O_4738,N_48914,N_49836);
and UO_4739 (O_4739,N_49227,N_48679);
or UO_4740 (O_4740,N_49388,N_49822);
or UO_4741 (O_4741,N_48102,N_49613);
or UO_4742 (O_4742,N_48336,N_49364);
xor UO_4743 (O_4743,N_48211,N_48229);
and UO_4744 (O_4744,N_48956,N_48545);
and UO_4745 (O_4745,N_49389,N_49481);
xor UO_4746 (O_4746,N_49754,N_48154);
or UO_4747 (O_4747,N_49533,N_48521);
and UO_4748 (O_4748,N_48166,N_49442);
nor UO_4749 (O_4749,N_48216,N_48473);
and UO_4750 (O_4750,N_49039,N_49227);
xor UO_4751 (O_4751,N_48807,N_49949);
nand UO_4752 (O_4752,N_49757,N_49199);
nand UO_4753 (O_4753,N_48770,N_48799);
nor UO_4754 (O_4754,N_49363,N_49769);
nand UO_4755 (O_4755,N_49721,N_48506);
nor UO_4756 (O_4756,N_48852,N_48364);
nand UO_4757 (O_4757,N_49044,N_48303);
nor UO_4758 (O_4758,N_48779,N_49724);
nand UO_4759 (O_4759,N_48448,N_48337);
and UO_4760 (O_4760,N_48597,N_48214);
nor UO_4761 (O_4761,N_49127,N_48502);
or UO_4762 (O_4762,N_49564,N_48110);
or UO_4763 (O_4763,N_48274,N_49038);
nor UO_4764 (O_4764,N_49034,N_48502);
nor UO_4765 (O_4765,N_49954,N_49753);
nand UO_4766 (O_4766,N_48426,N_49986);
or UO_4767 (O_4767,N_48135,N_49083);
and UO_4768 (O_4768,N_49486,N_48528);
nor UO_4769 (O_4769,N_49123,N_49090);
nand UO_4770 (O_4770,N_48408,N_48564);
or UO_4771 (O_4771,N_48394,N_49405);
xnor UO_4772 (O_4772,N_48898,N_49167);
or UO_4773 (O_4773,N_49431,N_49812);
and UO_4774 (O_4774,N_49537,N_49948);
xor UO_4775 (O_4775,N_49656,N_48562);
nand UO_4776 (O_4776,N_48627,N_48225);
nor UO_4777 (O_4777,N_49176,N_49512);
nor UO_4778 (O_4778,N_48449,N_49957);
nand UO_4779 (O_4779,N_48424,N_49016);
nand UO_4780 (O_4780,N_48186,N_48093);
xor UO_4781 (O_4781,N_49932,N_48537);
nand UO_4782 (O_4782,N_48467,N_49504);
or UO_4783 (O_4783,N_49725,N_49852);
and UO_4784 (O_4784,N_48326,N_48467);
nor UO_4785 (O_4785,N_48999,N_49262);
and UO_4786 (O_4786,N_49742,N_48109);
nand UO_4787 (O_4787,N_49548,N_48470);
nor UO_4788 (O_4788,N_49164,N_48974);
nor UO_4789 (O_4789,N_49146,N_49068);
or UO_4790 (O_4790,N_49762,N_48908);
nor UO_4791 (O_4791,N_48870,N_48005);
and UO_4792 (O_4792,N_48962,N_49795);
or UO_4793 (O_4793,N_48657,N_48124);
nand UO_4794 (O_4794,N_49640,N_48203);
nand UO_4795 (O_4795,N_49408,N_49449);
nor UO_4796 (O_4796,N_49981,N_48575);
and UO_4797 (O_4797,N_49427,N_49304);
and UO_4798 (O_4798,N_48872,N_48809);
nor UO_4799 (O_4799,N_49269,N_49842);
nand UO_4800 (O_4800,N_48714,N_49912);
nor UO_4801 (O_4801,N_48284,N_48994);
or UO_4802 (O_4802,N_49549,N_48461);
nor UO_4803 (O_4803,N_49718,N_48079);
and UO_4804 (O_4804,N_48384,N_48528);
and UO_4805 (O_4805,N_49356,N_48169);
and UO_4806 (O_4806,N_49999,N_49907);
or UO_4807 (O_4807,N_48830,N_49293);
and UO_4808 (O_4808,N_49676,N_48212);
xnor UO_4809 (O_4809,N_48196,N_49639);
nor UO_4810 (O_4810,N_48100,N_49283);
nand UO_4811 (O_4811,N_49339,N_48064);
xnor UO_4812 (O_4812,N_49317,N_48682);
nand UO_4813 (O_4813,N_48817,N_49775);
xnor UO_4814 (O_4814,N_49414,N_48030);
or UO_4815 (O_4815,N_48381,N_48327);
or UO_4816 (O_4816,N_49291,N_49712);
nand UO_4817 (O_4817,N_48111,N_48619);
nor UO_4818 (O_4818,N_49010,N_48748);
xnor UO_4819 (O_4819,N_49909,N_49694);
xnor UO_4820 (O_4820,N_48437,N_48742);
nand UO_4821 (O_4821,N_48780,N_48914);
or UO_4822 (O_4822,N_48185,N_49336);
or UO_4823 (O_4823,N_49932,N_49114);
nand UO_4824 (O_4824,N_48107,N_49307);
or UO_4825 (O_4825,N_49528,N_48816);
and UO_4826 (O_4826,N_49132,N_48588);
nand UO_4827 (O_4827,N_49211,N_48684);
nor UO_4828 (O_4828,N_48358,N_48990);
nor UO_4829 (O_4829,N_49871,N_48258);
or UO_4830 (O_4830,N_48151,N_49313);
or UO_4831 (O_4831,N_49151,N_49551);
and UO_4832 (O_4832,N_49639,N_49006);
and UO_4833 (O_4833,N_48288,N_48347);
or UO_4834 (O_4834,N_48774,N_48983);
and UO_4835 (O_4835,N_49090,N_49240);
or UO_4836 (O_4836,N_48063,N_49308);
and UO_4837 (O_4837,N_49588,N_49580);
nor UO_4838 (O_4838,N_48861,N_49689);
nand UO_4839 (O_4839,N_48670,N_49425);
xnor UO_4840 (O_4840,N_49985,N_49316);
xor UO_4841 (O_4841,N_48087,N_48849);
nor UO_4842 (O_4842,N_49782,N_49149);
and UO_4843 (O_4843,N_49209,N_48168);
nor UO_4844 (O_4844,N_49838,N_49022);
nand UO_4845 (O_4845,N_49201,N_49801);
and UO_4846 (O_4846,N_48371,N_48146);
xor UO_4847 (O_4847,N_49570,N_48806);
nand UO_4848 (O_4848,N_48839,N_49303);
nand UO_4849 (O_4849,N_48964,N_48136);
or UO_4850 (O_4850,N_48916,N_49009);
or UO_4851 (O_4851,N_48490,N_49857);
or UO_4852 (O_4852,N_48030,N_49728);
xnor UO_4853 (O_4853,N_49426,N_48562);
nand UO_4854 (O_4854,N_48860,N_49901);
nor UO_4855 (O_4855,N_49697,N_49765);
or UO_4856 (O_4856,N_49293,N_48159);
and UO_4857 (O_4857,N_48159,N_49028);
or UO_4858 (O_4858,N_49621,N_48430);
nand UO_4859 (O_4859,N_48637,N_48124);
or UO_4860 (O_4860,N_48656,N_48835);
or UO_4861 (O_4861,N_48979,N_48717);
and UO_4862 (O_4862,N_49574,N_49492);
nand UO_4863 (O_4863,N_49707,N_49011);
or UO_4864 (O_4864,N_49652,N_49387);
or UO_4865 (O_4865,N_49803,N_48055);
and UO_4866 (O_4866,N_48493,N_49908);
and UO_4867 (O_4867,N_49916,N_48267);
nand UO_4868 (O_4868,N_48099,N_48536);
or UO_4869 (O_4869,N_48211,N_48863);
xor UO_4870 (O_4870,N_49077,N_48006);
xnor UO_4871 (O_4871,N_49661,N_48612);
nor UO_4872 (O_4872,N_48334,N_48242);
nand UO_4873 (O_4873,N_49158,N_48700);
xor UO_4874 (O_4874,N_49953,N_49005);
nor UO_4875 (O_4875,N_48871,N_49421);
nor UO_4876 (O_4876,N_48619,N_48016);
or UO_4877 (O_4877,N_48192,N_48195);
nor UO_4878 (O_4878,N_48716,N_49621);
and UO_4879 (O_4879,N_48927,N_49665);
nor UO_4880 (O_4880,N_48695,N_48277);
nand UO_4881 (O_4881,N_49948,N_49855);
nor UO_4882 (O_4882,N_48294,N_48007);
nor UO_4883 (O_4883,N_48800,N_49332);
nor UO_4884 (O_4884,N_49853,N_48260);
xor UO_4885 (O_4885,N_49558,N_48184);
or UO_4886 (O_4886,N_48099,N_48479);
and UO_4887 (O_4887,N_49385,N_48124);
nor UO_4888 (O_4888,N_49845,N_48229);
xor UO_4889 (O_4889,N_49098,N_49386);
nand UO_4890 (O_4890,N_48843,N_48046);
or UO_4891 (O_4891,N_48382,N_49460);
nor UO_4892 (O_4892,N_48821,N_48328);
or UO_4893 (O_4893,N_49378,N_48674);
nor UO_4894 (O_4894,N_49747,N_48047);
nor UO_4895 (O_4895,N_49967,N_49252);
or UO_4896 (O_4896,N_49841,N_49822);
xnor UO_4897 (O_4897,N_49230,N_49374);
nor UO_4898 (O_4898,N_49214,N_49043);
nor UO_4899 (O_4899,N_49230,N_49455);
or UO_4900 (O_4900,N_49536,N_49503);
nand UO_4901 (O_4901,N_49543,N_48666);
nor UO_4902 (O_4902,N_48743,N_49428);
nor UO_4903 (O_4903,N_48516,N_49501);
xor UO_4904 (O_4904,N_49609,N_48026);
nor UO_4905 (O_4905,N_48099,N_48132);
xor UO_4906 (O_4906,N_48739,N_49100);
xnor UO_4907 (O_4907,N_49775,N_48699);
or UO_4908 (O_4908,N_48773,N_48260);
xor UO_4909 (O_4909,N_49114,N_49665);
nand UO_4910 (O_4910,N_49262,N_49522);
and UO_4911 (O_4911,N_49663,N_48201);
xor UO_4912 (O_4912,N_49769,N_49732);
xnor UO_4913 (O_4913,N_48474,N_48795);
or UO_4914 (O_4914,N_49343,N_49726);
and UO_4915 (O_4915,N_48178,N_48869);
xor UO_4916 (O_4916,N_49045,N_48583);
or UO_4917 (O_4917,N_48487,N_48479);
xor UO_4918 (O_4918,N_48846,N_48544);
xor UO_4919 (O_4919,N_49283,N_49566);
xor UO_4920 (O_4920,N_49695,N_48726);
and UO_4921 (O_4921,N_49211,N_49018);
xor UO_4922 (O_4922,N_48001,N_49776);
nor UO_4923 (O_4923,N_49025,N_49174);
and UO_4924 (O_4924,N_48945,N_48340);
xor UO_4925 (O_4925,N_48857,N_49425);
xor UO_4926 (O_4926,N_48703,N_48344);
and UO_4927 (O_4927,N_48463,N_48745);
nand UO_4928 (O_4928,N_49926,N_48635);
or UO_4929 (O_4929,N_48677,N_48007);
nand UO_4930 (O_4930,N_49613,N_48934);
and UO_4931 (O_4931,N_49298,N_49290);
xor UO_4932 (O_4932,N_49606,N_49927);
or UO_4933 (O_4933,N_49217,N_49340);
nor UO_4934 (O_4934,N_48685,N_48872);
and UO_4935 (O_4935,N_49664,N_49212);
xnor UO_4936 (O_4936,N_49330,N_49975);
nor UO_4937 (O_4937,N_48518,N_48666);
and UO_4938 (O_4938,N_49288,N_49701);
and UO_4939 (O_4939,N_48710,N_48449);
or UO_4940 (O_4940,N_48672,N_48939);
nand UO_4941 (O_4941,N_49395,N_49778);
nand UO_4942 (O_4942,N_49226,N_49415);
nand UO_4943 (O_4943,N_48665,N_49580);
nand UO_4944 (O_4944,N_49739,N_49118);
and UO_4945 (O_4945,N_49033,N_49525);
and UO_4946 (O_4946,N_48407,N_48394);
or UO_4947 (O_4947,N_49438,N_48191);
nor UO_4948 (O_4948,N_49753,N_48831);
nand UO_4949 (O_4949,N_48551,N_48715);
or UO_4950 (O_4950,N_49354,N_49318);
or UO_4951 (O_4951,N_48472,N_48603);
nor UO_4952 (O_4952,N_48741,N_49482);
nand UO_4953 (O_4953,N_49253,N_49413);
nand UO_4954 (O_4954,N_49840,N_48924);
or UO_4955 (O_4955,N_48519,N_49288);
and UO_4956 (O_4956,N_48175,N_48303);
xor UO_4957 (O_4957,N_49983,N_49402);
nor UO_4958 (O_4958,N_49840,N_48332);
nand UO_4959 (O_4959,N_49286,N_48139);
nor UO_4960 (O_4960,N_49649,N_49514);
xnor UO_4961 (O_4961,N_49947,N_48121);
and UO_4962 (O_4962,N_48166,N_49898);
xor UO_4963 (O_4963,N_48633,N_48375);
nor UO_4964 (O_4964,N_49638,N_49629);
xor UO_4965 (O_4965,N_49726,N_49503);
and UO_4966 (O_4966,N_48900,N_48522);
or UO_4967 (O_4967,N_48778,N_49198);
and UO_4968 (O_4968,N_49820,N_48814);
and UO_4969 (O_4969,N_49704,N_48157);
or UO_4970 (O_4970,N_48641,N_49855);
nand UO_4971 (O_4971,N_49088,N_49248);
and UO_4972 (O_4972,N_49469,N_49841);
xor UO_4973 (O_4973,N_49332,N_49947);
nand UO_4974 (O_4974,N_48625,N_49718);
nor UO_4975 (O_4975,N_48790,N_48327);
nor UO_4976 (O_4976,N_49625,N_48690);
nor UO_4977 (O_4977,N_48474,N_49148);
xor UO_4978 (O_4978,N_48210,N_49344);
and UO_4979 (O_4979,N_49868,N_48726);
or UO_4980 (O_4980,N_49821,N_49539);
xnor UO_4981 (O_4981,N_49521,N_48169);
or UO_4982 (O_4982,N_48479,N_48928);
or UO_4983 (O_4983,N_49095,N_48566);
nand UO_4984 (O_4984,N_48425,N_49955);
and UO_4985 (O_4985,N_49213,N_48265);
nor UO_4986 (O_4986,N_49100,N_49343);
xnor UO_4987 (O_4987,N_48184,N_49647);
and UO_4988 (O_4988,N_49139,N_49502);
or UO_4989 (O_4989,N_49894,N_48076);
or UO_4990 (O_4990,N_48837,N_48698);
nor UO_4991 (O_4991,N_48961,N_48888);
nand UO_4992 (O_4992,N_49382,N_49352);
and UO_4993 (O_4993,N_49335,N_48464);
nor UO_4994 (O_4994,N_49360,N_48521);
nand UO_4995 (O_4995,N_48457,N_48962);
nand UO_4996 (O_4996,N_49481,N_48444);
xor UO_4997 (O_4997,N_48132,N_48563);
xor UO_4998 (O_4998,N_48919,N_48683);
and UO_4999 (O_4999,N_49534,N_49609);
endmodule