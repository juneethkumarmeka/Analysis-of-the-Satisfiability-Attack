module basic_2000_20000_2500_5_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1504,In_580);
or U1 (N_1,In_1676,In_184);
and U2 (N_2,In_1476,In_1085);
and U3 (N_3,In_1649,In_1180);
nand U4 (N_4,In_1708,In_966);
or U5 (N_5,In_222,In_1909);
nor U6 (N_6,In_1287,In_1789);
and U7 (N_7,In_1162,In_1128);
nand U8 (N_8,In_1556,In_1099);
or U9 (N_9,In_479,In_169);
and U10 (N_10,In_1996,In_216);
or U11 (N_11,In_288,In_1665);
nor U12 (N_12,In_827,In_1381);
or U13 (N_13,In_395,In_1118);
or U14 (N_14,In_563,In_562);
nor U15 (N_15,In_694,In_1343);
and U16 (N_16,In_1150,In_1368);
nand U17 (N_17,In_592,In_1011);
and U18 (N_18,In_1643,In_1289);
nor U19 (N_19,In_30,In_205);
or U20 (N_20,In_1443,In_241);
or U21 (N_21,In_27,In_1861);
nor U22 (N_22,In_412,In_746);
and U23 (N_23,In_1897,In_75);
or U24 (N_24,In_1550,In_1396);
or U25 (N_25,In_564,In_1592);
nor U26 (N_26,In_541,In_76);
nor U27 (N_27,In_835,In_788);
and U28 (N_28,In_194,In_1639);
and U29 (N_29,In_1572,In_1647);
nand U30 (N_30,In_140,In_1108);
and U31 (N_31,In_1153,In_1740);
nor U32 (N_32,In_1765,In_1246);
and U33 (N_33,In_1406,In_1815);
and U34 (N_34,In_547,In_203);
nor U35 (N_35,In_1673,In_1116);
and U36 (N_36,In_1501,In_1972);
nor U37 (N_37,In_17,In_1553);
nand U38 (N_38,In_709,In_1030);
nor U39 (N_39,In_811,In_891);
and U40 (N_40,In_881,In_814);
and U41 (N_41,In_62,In_807);
and U42 (N_42,In_1320,In_929);
or U43 (N_43,In_857,In_1859);
nand U44 (N_44,In_1088,In_1399);
or U45 (N_45,In_317,In_283);
and U46 (N_46,In_1461,In_634);
nor U47 (N_47,In_1973,In_383);
and U48 (N_48,In_110,In_1791);
and U49 (N_49,In_1210,In_561);
and U50 (N_50,In_644,In_752);
or U51 (N_51,In_389,In_526);
and U52 (N_52,In_687,In_1355);
or U53 (N_53,In_1640,In_1818);
nor U54 (N_54,In_147,In_1117);
and U55 (N_55,In_825,In_408);
and U56 (N_56,In_287,In_204);
and U57 (N_57,In_809,In_94);
nand U58 (N_58,In_1232,In_1826);
or U59 (N_59,In_1025,In_1426);
and U60 (N_60,In_760,In_1956);
and U61 (N_61,In_294,In_1042);
nor U62 (N_62,In_1615,In_625);
xnor U63 (N_63,In_1159,In_1823);
or U64 (N_64,In_1415,In_742);
xor U65 (N_65,In_1876,In_1067);
or U66 (N_66,In_1429,In_103);
nand U67 (N_67,In_1090,In_1397);
xor U68 (N_68,In_804,In_696);
or U69 (N_69,In_961,In_1837);
and U70 (N_70,In_165,In_445);
nor U71 (N_71,In_1511,In_671);
nor U72 (N_72,In_2,In_869);
nor U73 (N_73,In_47,In_1980);
and U74 (N_74,In_1022,In_1908);
or U75 (N_75,In_1546,In_496);
or U76 (N_76,In_1277,In_1294);
and U77 (N_77,In_1903,In_985);
and U78 (N_78,In_873,In_1228);
nor U79 (N_79,In_552,In_1189);
nand U80 (N_80,In_720,In_1080);
and U81 (N_81,In_1267,In_144);
or U82 (N_82,In_1796,In_289);
nand U83 (N_83,In_594,In_844);
nand U84 (N_84,In_1503,In_1238);
and U85 (N_85,In_500,In_662);
or U86 (N_86,In_315,In_1590);
and U87 (N_87,In_1328,In_485);
nand U88 (N_88,In_1004,In_64);
xor U89 (N_89,In_793,In_557);
and U90 (N_90,In_196,In_1253);
or U91 (N_91,In_1687,In_1341);
xnor U92 (N_92,In_1037,In_1220);
or U93 (N_93,In_1339,In_1691);
xnor U94 (N_94,In_36,In_134);
nor U95 (N_95,In_1035,In_1172);
and U96 (N_96,In_708,In_753);
nor U97 (N_97,In_1878,In_382);
or U98 (N_98,In_319,In_763);
and U99 (N_99,In_1616,In_642);
or U100 (N_100,In_1833,In_1979);
or U101 (N_101,In_729,In_798);
nand U102 (N_102,In_695,In_422);
and U103 (N_103,In_1281,In_356);
nor U104 (N_104,In_750,In_1974);
and U105 (N_105,In_385,In_164);
xnor U106 (N_106,In_322,In_1070);
nand U107 (N_107,In_89,In_1419);
nand U108 (N_108,In_0,In_840);
or U109 (N_109,In_1138,In_107);
xnor U110 (N_110,In_578,In_1911);
xnor U111 (N_111,In_431,In_972);
nor U112 (N_112,In_1050,In_1717);
or U113 (N_113,In_1814,In_468);
nand U114 (N_114,In_55,In_1068);
and U115 (N_115,In_1268,In_1186);
nand U116 (N_116,In_1191,In_900);
nor U117 (N_117,In_1678,In_157);
xnor U118 (N_118,In_499,In_1155);
nor U119 (N_119,In_1487,In_1283);
nand U120 (N_120,In_1872,In_178);
nor U121 (N_121,In_1599,In_968);
nand U122 (N_122,In_1907,In_704);
nor U123 (N_123,In_1927,In_1243);
or U124 (N_124,In_1889,In_1266);
nand U125 (N_125,In_1654,In_1557);
and U126 (N_126,In_964,In_1611);
and U127 (N_127,In_1223,In_778);
and U128 (N_128,In_576,In_1888);
nor U129 (N_129,In_1910,In_718);
nor U130 (N_130,In_569,In_609);
or U131 (N_131,In_1177,In_1646);
or U132 (N_132,In_1916,In_1655);
nand U133 (N_133,In_273,In_138);
nor U134 (N_134,In_951,In_214);
or U135 (N_135,In_618,In_751);
and U136 (N_136,In_975,In_652);
and U137 (N_137,In_1602,In_1432);
nor U138 (N_138,In_713,In_610);
and U139 (N_139,In_691,In_769);
and U140 (N_140,In_643,In_1403);
nand U141 (N_141,In_1781,In_1902);
or U142 (N_142,In_785,In_675);
nand U143 (N_143,In_1650,In_724);
or U144 (N_144,In_1523,In_1212);
xor U145 (N_145,In_321,In_1808);
and U146 (N_146,In_1024,In_682);
nor U147 (N_147,In_1695,In_854);
nand U148 (N_148,In_1554,In_1405);
and U149 (N_149,In_297,In_882);
or U150 (N_150,In_145,In_721);
nor U151 (N_151,In_3,In_84);
and U152 (N_152,In_1510,In_1113);
nor U153 (N_153,In_52,In_1997);
or U154 (N_154,In_1658,In_166);
and U155 (N_155,In_1385,In_684);
nand U156 (N_156,In_626,In_417);
nand U157 (N_157,In_822,In_60);
nand U158 (N_158,In_660,In_98);
xor U159 (N_159,In_1652,In_1474);
nor U160 (N_160,In_1747,In_1761);
and U161 (N_161,In_1087,In_1959);
nor U162 (N_162,In_1059,In_1240);
nand U163 (N_163,In_1352,In_109);
or U164 (N_164,In_1924,In_767);
or U165 (N_165,In_1757,In_1058);
nor U166 (N_166,In_1401,In_935);
nor U167 (N_167,In_722,In_1104);
nor U168 (N_168,In_1567,In_1288);
and U169 (N_169,In_1192,In_108);
and U170 (N_170,In_1096,In_88);
xor U171 (N_171,In_1386,In_1136);
nand U172 (N_172,In_1930,In_1482);
and U173 (N_173,In_359,In_1026);
nor U174 (N_174,In_510,In_1142);
nand U175 (N_175,In_544,In_1200);
nand U176 (N_176,In_673,In_39);
and U177 (N_177,In_43,In_1871);
and U178 (N_178,In_1347,In_1437);
nor U179 (N_179,In_1251,In_1873);
nand U180 (N_180,In_1485,In_787);
and U181 (N_181,In_930,In_1923);
and U182 (N_182,In_831,In_1097);
nand U183 (N_183,In_1756,In_387);
xor U184 (N_184,In_1742,In_1867);
xor U185 (N_185,In_796,In_608);
nor U186 (N_186,In_1530,In_71);
or U187 (N_187,In_1129,In_1904);
or U188 (N_188,In_363,In_1741);
nand U189 (N_189,In_953,In_845);
xnor U190 (N_190,In_493,In_365);
nand U191 (N_191,In_420,In_1311);
nor U192 (N_192,In_350,In_1976);
xnor U193 (N_193,In_1651,In_923);
or U194 (N_194,In_364,In_1953);
or U195 (N_195,In_1774,In_1008);
and U196 (N_196,In_1166,In_316);
and U197 (N_197,In_1679,In_534);
and U198 (N_198,In_484,In_1753);
nor U199 (N_199,In_902,In_864);
and U200 (N_200,In_791,In_1086);
nand U201 (N_201,In_4,In_946);
or U202 (N_202,In_1064,In_952);
nand U203 (N_203,In_1562,In_1805);
and U204 (N_204,In_162,In_1028);
and U205 (N_205,In_1460,In_16);
and U206 (N_206,In_1854,In_325);
nor U207 (N_207,In_1327,In_593);
nor U208 (N_208,In_310,In_498);
or U209 (N_209,In_1293,In_1879);
or U210 (N_210,In_253,In_1962);
nor U211 (N_211,In_72,In_1614);
nand U212 (N_212,In_358,In_768);
and U213 (N_213,In_1817,In_1473);
nor U214 (N_214,In_1792,In_56);
or U215 (N_215,In_1754,In_1298);
nand U216 (N_216,In_225,In_1937);
and U217 (N_217,In_1414,In_1346);
nand U218 (N_218,In_1221,In_320);
nand U219 (N_219,In_40,In_471);
nor U220 (N_220,In_1842,In_220);
nand U221 (N_221,In_1998,In_1899);
and U222 (N_222,In_601,In_1621);
or U223 (N_223,In_828,In_209);
and U224 (N_224,In_1834,In_1604);
and U225 (N_225,In_855,In_597);
or U226 (N_226,In_1526,In_432);
nand U227 (N_227,In_217,In_105);
or U228 (N_228,In_1069,In_1380);
and U229 (N_229,In_53,In_697);
or U230 (N_230,In_558,In_1536);
and U231 (N_231,In_243,In_415);
or U232 (N_232,In_1093,In_1292);
or U233 (N_233,In_645,In_237);
and U234 (N_234,In_372,In_1726);
nand U235 (N_235,In_714,In_1723);
xnor U236 (N_236,In_546,In_911);
or U237 (N_237,In_780,In_48);
nand U238 (N_238,In_648,In_1768);
nand U239 (N_239,In_1775,In_565);
nor U240 (N_240,In_837,In_1565);
or U241 (N_241,In_206,In_1217);
or U242 (N_242,In_13,In_1417);
or U243 (N_243,In_1811,In_1544);
and U244 (N_244,In_1140,In_374);
xor U245 (N_245,In_477,In_616);
nor U246 (N_246,In_438,In_161);
and U247 (N_247,In_117,In_605);
nor U248 (N_248,In_1705,In_611);
nor U249 (N_249,In_1364,In_1706);
nand U250 (N_250,In_1115,In_1812);
nand U251 (N_251,In_1609,In_1079);
nor U252 (N_252,In_454,In_330);
xnor U253 (N_253,In_1048,In_517);
or U254 (N_254,In_235,In_37);
or U255 (N_255,In_81,In_1569);
and U256 (N_256,In_153,In_1944);
nand U257 (N_257,In_1170,In_581);
xnor U258 (N_258,In_1558,In_1940);
nand U259 (N_259,In_497,In_888);
nor U260 (N_260,In_529,In_451);
or U261 (N_261,In_921,In_1074);
or U262 (N_262,In_1901,In_1126);
or U263 (N_263,In_1769,In_537);
xor U264 (N_264,In_749,In_1946);
xnor U265 (N_265,In_180,In_1636);
and U266 (N_266,In_360,In_1955);
and U267 (N_267,In_327,In_1310);
xor U268 (N_268,In_743,In_1506);
and U269 (N_269,In_667,In_647);
nor U270 (N_270,In_489,In_1541);
and U271 (N_271,In_514,In_460);
nand U272 (N_272,In_1454,In_1653);
nand U273 (N_273,In_851,In_223);
nand U274 (N_274,In_755,In_914);
nand U275 (N_275,In_137,In_861);
nand U276 (N_276,In_308,In_1110);
or U277 (N_277,In_349,In_817);
or U278 (N_278,In_1819,In_1794);
and U279 (N_279,In_1407,In_920);
or U280 (N_280,In_1813,In_839);
or U281 (N_281,In_1578,In_1438);
or U282 (N_282,In_1807,In_1488);
nand U283 (N_283,In_1296,In_1049);
and U284 (N_284,In_764,In_1896);
or U285 (N_285,In_118,In_516);
nand U286 (N_286,In_324,In_1617);
nand U287 (N_287,In_434,In_450);
and U288 (N_288,In_1598,In_1696);
and U289 (N_289,In_1333,In_448);
nor U290 (N_290,In_182,In_1480);
nor U291 (N_291,In_958,In_249);
and U292 (N_292,In_1949,In_407);
or U293 (N_293,In_741,In_1683);
nand U294 (N_294,In_543,In_300);
nor U295 (N_295,In_136,In_1728);
nor U296 (N_296,In_1408,In_1999);
nor U297 (N_297,In_115,In_266);
nand U298 (N_298,In_379,In_1763);
nor U299 (N_299,In_1375,In_1202);
nand U300 (N_300,In_329,In_1785);
nand U301 (N_301,In_1083,In_1795);
nand U302 (N_302,In_1362,In_1669);
xor U303 (N_303,In_766,In_783);
and U304 (N_304,In_1969,In_1325);
nor U305 (N_305,In_442,In_1513);
nor U306 (N_306,In_863,In_1174);
or U307 (N_307,In_258,In_919);
and U308 (N_308,In_1077,In_171);
and U309 (N_309,In_1727,In_1701);
xnor U310 (N_310,In_802,In_1539);
or U311 (N_311,In_1305,In_1533);
or U312 (N_312,In_228,In_1231);
nand U313 (N_313,In_259,In_1951);
and U314 (N_314,In_439,In_824);
nor U315 (N_315,In_1936,In_1431);
and U316 (N_316,In_706,In_1627);
nor U317 (N_317,In_402,In_733);
nand U318 (N_318,In_712,In_621);
and U319 (N_319,In_245,In_511);
nor U320 (N_320,In_1586,In_1448);
xor U321 (N_321,In_1743,In_613);
nand U322 (N_322,In_1986,In_730);
and U323 (N_323,In_1787,In_1499);
nand U324 (N_324,In_624,In_686);
and U325 (N_325,In_1848,In_932);
nor U326 (N_326,In_1278,In_1199);
nand U327 (N_327,In_956,In_1442);
nor U328 (N_328,In_1032,In_1606);
or U329 (N_329,In_1856,In_1449);
nand U330 (N_330,In_1847,In_688);
nand U331 (N_331,In_163,In_111);
nor U332 (N_332,In_812,In_530);
or U333 (N_333,In_343,In_907);
xor U334 (N_334,In_1423,In_1486);
nor U335 (N_335,In_1481,In_1470);
or U336 (N_336,In_1056,In_1608);
xnor U337 (N_337,In_549,In_1379);
and U338 (N_338,In_872,In_1149);
or U339 (N_339,In_101,In_1773);
xor U340 (N_340,In_1273,In_1832);
nand U341 (N_341,In_1326,In_1033);
nor U342 (N_342,In_1181,In_1524);
xnor U343 (N_343,In_1988,In_925);
nor U344 (N_344,In_233,In_280);
and U345 (N_345,In_1182,In_1560);
or U346 (N_346,In_944,In_1404);
or U347 (N_347,In_650,In_191);
nand U348 (N_348,In_1134,In_1619);
nor U349 (N_349,In_1271,In_33);
nor U350 (N_350,In_1752,In_1600);
nand U351 (N_351,In_1017,In_1866);
nor U352 (N_352,In_1103,In_738);
and U353 (N_353,In_1451,In_843);
and U354 (N_354,In_285,In_1205);
and U355 (N_355,In_125,In_1816);
or U356 (N_356,In_1635,In_775);
nor U357 (N_357,In_674,In_370);
nand U358 (N_358,In_393,In_29);
nor U359 (N_359,In_988,In_571);
and U360 (N_360,In_1187,In_998);
nand U361 (N_361,In_232,In_403);
nor U362 (N_362,In_470,In_1314);
and U363 (N_363,In_1075,In_346);
xnor U364 (N_364,In_1633,In_1793);
and U365 (N_365,In_423,In_116);
nor U366 (N_366,In_1540,In_92);
nor U367 (N_367,In_969,In_1555);
nand U368 (N_368,In_1829,In_1915);
xnor U369 (N_369,In_1124,In_278);
nand U370 (N_370,In_995,In_1644);
nor U371 (N_371,In_661,In_70);
or U372 (N_372,In_416,In_1759);
nor U373 (N_373,In_1254,In_1632);
and U374 (N_374,In_1900,In_1534);
and U375 (N_375,In_1670,In_1421);
or U376 (N_376,In_1014,In_1393);
nor U377 (N_377,In_747,In_45);
and U378 (N_378,In_380,In_1006);
and U379 (N_379,In_937,In_1256);
nand U380 (N_380,In_539,In_362);
nor U381 (N_381,In_336,In_505);
and U382 (N_382,In_124,In_922);
and U383 (N_383,In_692,In_700);
and U384 (N_384,In_264,In_1309);
and U385 (N_385,In_1772,In_267);
and U386 (N_386,In_716,In_596);
or U387 (N_387,In_1089,In_281);
xnor U388 (N_388,In_1169,In_936);
nor U389 (N_389,In_392,In_1360);
and U390 (N_390,In_1013,In_523);
and U391 (N_391,In_1857,In_10);
xor U392 (N_392,In_1710,In_868);
nand U393 (N_393,In_462,In_666);
and U394 (N_394,In_390,In_51);
or U395 (N_395,In_1151,In_573);
nand U396 (N_396,In_1156,In_156);
or U397 (N_397,In_1890,In_1594);
or U398 (N_398,In_1722,In_1991);
nor U399 (N_399,In_1331,In_1363);
and U400 (N_400,In_351,In_229);
and U401 (N_401,In_1537,In_1342);
nand U402 (N_402,In_1402,In_1139);
or U403 (N_403,In_1265,In_1585);
xnor U404 (N_404,In_446,In_699);
nand U405 (N_405,In_1383,In_943);
and U406 (N_406,In_1841,In_1685);
nor U407 (N_407,In_876,In_779);
nor U408 (N_408,In_1167,In_1441);
and U409 (N_409,In_1471,In_856);
nand U410 (N_410,In_794,In_1580);
and U411 (N_411,In_848,In_1948);
nor U412 (N_412,In_348,In_503);
nand U413 (N_413,In_1332,In_1628);
nand U414 (N_414,In_834,In_1300);
nand U415 (N_415,In_1957,In_896);
nand U416 (N_416,In_1378,In_494);
nand U417 (N_417,In_104,In_1248);
nor U418 (N_418,In_120,In_352);
nor U419 (N_419,In_354,In_1637);
and U420 (N_420,In_332,In_1514);
and U421 (N_421,In_1307,In_1349);
xnor U422 (N_422,In_893,In_1564);
nand U423 (N_423,In_1881,In_355);
and U424 (N_424,In_1922,In_1786);
or U425 (N_425,In_252,In_1102);
nor U426 (N_426,In_464,In_1178);
nand U427 (N_427,In_967,In_149);
nor U428 (N_428,In_810,In_1713);
nand U429 (N_429,In_1960,In_274);
and U430 (N_430,In_765,In_1978);
nor U431 (N_431,In_121,In_654);
and U432 (N_432,In_1428,In_1027);
xor U433 (N_433,In_1329,In_521);
or U434 (N_434,In_1052,In_1122);
and U435 (N_435,In_282,In_665);
and U436 (N_436,In_759,In_212);
or U437 (N_437,In_299,In_97);
xor U438 (N_438,In_1509,In_744);
or U439 (N_439,In_1316,In_1472);
nor U440 (N_440,In_1954,In_1684);
or U441 (N_441,In_1571,In_1450);
and U442 (N_442,In_246,In_106);
or U443 (N_443,In_155,In_640);
xor U444 (N_444,In_532,In_1838);
and U445 (N_445,In_268,In_545);
and U446 (N_446,In_813,In_1098);
nor U447 (N_447,In_711,In_1719);
nor U448 (N_448,In_483,In_1931);
and U449 (N_449,In_1222,In_559);
nor U450 (N_450,In_427,In_1276);
and U451 (N_451,In_1970,In_1797);
and U452 (N_452,In_1395,In_1051);
nand U453 (N_453,In_1622,In_1733);
nand U454 (N_454,In_242,In_1041);
nor U455 (N_455,In_880,In_632);
and U456 (N_456,In_947,In_172);
and U457 (N_457,In_1508,In_1100);
nand U458 (N_458,In_916,In_1777);
and U459 (N_459,In_179,In_1947);
xnor U460 (N_460,In_502,In_435);
nor U461 (N_461,In_1681,In_1799);
nor U462 (N_462,In_1433,In_177);
and U463 (N_463,In_1965,In_1732);
xor U464 (N_464,In_1301,In_112);
or U465 (N_465,In_1870,In_1840);
and U466 (N_466,In_962,In_1993);
xnor U467 (N_467,In_871,In_955);
nand U468 (N_468,In_1709,In_821);
and U469 (N_469,In_91,In_82);
or U470 (N_470,In_1642,In_1591);
nor U471 (N_471,In_527,In_95);
or U472 (N_472,In_404,In_41);
nand U473 (N_473,In_192,In_1843);
or U474 (N_474,In_1892,In_135);
xor U475 (N_475,In_1945,In_1929);
xnor U476 (N_476,In_859,In_79);
nand U477 (N_477,In_984,In_368);
and U478 (N_478,In_226,In_548);
and U479 (N_479,In_1519,In_1858);
or U480 (N_480,In_619,In_1559);
or U481 (N_481,In_1545,In_1928);
and U482 (N_482,In_1682,In_44);
or U483 (N_483,In_1127,In_478);
and U484 (N_484,In_1498,In_829);
or U485 (N_485,In_334,In_982);
and U486 (N_486,In_614,In_940);
or U487 (N_487,In_1109,In_292);
nand U488 (N_488,In_606,In_1912);
or U489 (N_489,In_838,In_1365);
nand U490 (N_490,In_1680,In_1737);
and U491 (N_491,In_1641,In_690);
nor U492 (N_492,In_1358,In_1666);
nor U493 (N_493,In_1895,In_1446);
and U494 (N_494,In_1515,In_656);
and U495 (N_495,In_1891,In_1764);
and U496 (N_496,In_141,In_50);
and U497 (N_497,In_1313,In_18);
xor U498 (N_498,In_190,In_286);
and U499 (N_499,In_90,In_1547);
xor U500 (N_500,In_586,In_1259);
nor U501 (N_501,In_202,In_1361);
nor U502 (N_502,In_1040,In_1146);
and U503 (N_503,In_1111,In_14);
or U504 (N_504,In_490,In_131);
nand U505 (N_505,In_1046,In_87);
xnor U506 (N_506,In_506,In_8);
nand U507 (N_507,In_1703,In_792);
and U508 (N_508,In_1625,In_1168);
nor U509 (N_509,In_790,In_465);
nand U510 (N_510,In_1001,In_1880);
nand U511 (N_511,In_1274,In_1661);
and U512 (N_512,In_1983,In_1822);
and U513 (N_513,In_1464,In_992);
and U514 (N_514,In_1458,In_928);
and U515 (N_515,In_627,In_1018);
and U516 (N_516,In_1073,In_1282);
xnor U517 (N_517,In_649,In_361);
xor U518 (N_518,In_1055,In_1101);
nor U519 (N_519,In_58,In_1179);
nor U520 (N_520,In_1106,In_1260);
nor U521 (N_521,In_1543,In_870);
nand U522 (N_522,In_425,In_776);
and U523 (N_523,In_1914,In_1053);
nor U524 (N_524,In_452,In_1502);
or U525 (N_525,In_1987,In_1345);
nand U526 (N_526,In_414,In_187);
nor U527 (N_527,In_1425,In_257);
and U528 (N_528,In_378,In_710);
or U529 (N_529,In_1739,In_398);
and U530 (N_530,In_1551,In_23);
nand U531 (N_531,In_189,In_1734);
xor U532 (N_532,In_68,In_622);
or U533 (N_533,In_1092,In_1123);
and U534 (N_534,In_528,In_1330);
nor U535 (N_535,In_1452,In_1218);
or U536 (N_536,In_175,In_657);
and U537 (N_537,In_1771,In_284);
nor U538 (N_538,In_1459,In_1766);
or U539 (N_539,In_1917,In_188);
nand U540 (N_540,In_717,In_1337);
or U541 (N_541,In_251,In_1427);
nand U542 (N_542,In_1020,In_472);
or U543 (N_543,In_1664,In_1424);
nor U544 (N_544,In_1029,In_1262);
nand U545 (N_545,In_467,In_1357);
or U546 (N_546,In_1236,In_1318);
nor U547 (N_547,In_1207,In_719);
nand U548 (N_548,In_5,In_331);
or U549 (N_549,In_1645,In_1820);
or U550 (N_550,In_949,In_799);
and U551 (N_551,In_1835,In_400);
or U552 (N_552,In_860,In_1084);
or U553 (N_553,In_1469,In_1152);
nor U554 (N_554,In_974,In_1216);
or U555 (N_555,In_1894,In_739);
and U556 (N_556,In_602,In_761);
nand U557 (N_557,In_1990,In_455);
xor U558 (N_558,In_231,In_173);
nor U559 (N_559,In_1694,In_453);
nor U560 (N_560,In_1392,In_1164);
and U561 (N_561,In_195,In_1264);
nand U562 (N_562,In_852,In_1938);
or U563 (N_563,In_1648,In_123);
nor U564 (N_564,In_979,In_1755);
and U565 (N_565,In_1776,In_1354);
nor U566 (N_566,In_1490,In_1507);
nor U567 (N_567,In_1574,In_818);
or U568 (N_568,In_910,In_890);
and U569 (N_569,In_1675,In_976);
nor U570 (N_570,In_883,In_617);
and U571 (N_571,In_1570,In_129);
and U572 (N_572,In_1725,In_1994);
or U573 (N_573,In_826,In_1114);
and U574 (N_574,In_1010,In_1319);
or U575 (N_575,In_815,In_1925);
nand U576 (N_576,In_1731,In_1984);
nand U577 (N_577,In_1370,In_1334);
nor U578 (N_578,In_1071,In_1121);
nand U579 (N_579,In_1107,In_784);
and U580 (N_580,In_723,In_1561);
nor U581 (N_581,In_1105,In_1824);
or U582 (N_582,In_1809,In_1291);
xor U583 (N_583,In_1657,In_1788);
nor U584 (N_584,In_1783,In_1157);
nor U585 (N_585,In_1275,In_369);
nor U586 (N_586,In_1453,In_1389);
or U587 (N_587,In_554,In_1981);
or U588 (N_588,In_1827,In_905);
xor U589 (N_589,In_1631,In_126);
nand U590 (N_590,In_208,In_1801);
nor U591 (N_591,In_227,In_1230);
and U592 (N_592,In_1692,In_938);
or U593 (N_593,In_1885,In_522);
and U594 (N_594,In_1005,In_913);
xor U595 (N_595,In_1237,In_19);
and U596 (N_596,In_629,In_1009);
and U597 (N_597,In_1875,In_1435);
or U598 (N_598,In_1197,In_430);
xnor U599 (N_599,In_707,In_850);
nor U600 (N_600,In_591,In_1031);
nand U601 (N_601,In_1884,In_1462);
or U602 (N_602,In_428,In_1712);
nand U603 (N_603,In_1702,In_1057);
or U604 (N_604,In_1868,In_770);
and U605 (N_605,In_12,In_312);
xor U606 (N_606,In_1803,In_1295);
nor U607 (N_607,In_1760,In_1985);
and U608 (N_608,In_1527,In_970);
and U609 (N_609,In_26,In_550);
nand U610 (N_610,In_933,In_449);
nor U611 (N_611,In_376,In_1410);
and U612 (N_612,In_1376,In_1601);
nor U613 (N_613,In_1855,In_1623);
and U614 (N_614,In_1227,In_122);
nor U615 (N_615,In_858,In_474);
xor U616 (N_616,In_1893,In_210);
or U617 (N_617,In_1290,In_1700);
nand U618 (N_618,In_1196,In_85);
nor U619 (N_619,In_65,In_386);
or U620 (N_620,In_291,In_909);
and U621 (N_621,In_808,In_1491);
and U622 (N_622,In_168,In_1467);
or U623 (N_623,In_1577,In_1047);
xor U624 (N_624,In_328,In_1500);
and U625 (N_625,In_820,In_6);
nand U626 (N_626,In_67,In_1918);
nor U627 (N_627,In_139,In_555);
and U628 (N_628,In_978,In_679);
nand U629 (N_629,In_1939,In_680);
nand U630 (N_630,In_1758,In_823);
nor U631 (N_631,In_574,In_1384);
and U632 (N_632,In_1255,In_260);
and U633 (N_633,In_1249,In_832);
nand U634 (N_634,In_1887,In_797);
nand U635 (N_635,In_32,In_1724);
nor U636 (N_636,In_996,In_639);
nor U637 (N_637,In_469,In_1548);
nor U638 (N_638,In_303,In_424);
xnor U639 (N_639,In_481,In_941);
and U640 (N_640,In_1188,In_774);
nor U641 (N_641,In_333,In_276);
or U642 (N_642,In_1081,In_904);
nand U643 (N_643,In_250,In_583);
nand U644 (N_644,In_142,In_884);
xor U645 (N_645,In_167,In_781);
and U646 (N_646,In_339,In_119);
nand U647 (N_647,In_311,In_1831);
or U648 (N_648,In_304,In_296);
and U649 (N_649,In_1942,In_1697);
or U650 (N_650,In_1340,In_1324);
or U651 (N_651,In_256,In_1613);
or U652 (N_652,In_1012,In_501);
xor U653 (N_653,In_1517,In_293);
nor U654 (N_654,In_1494,In_239);
xnor U655 (N_655,In_1373,In_1213);
or U656 (N_656,In_748,In_672);
xor U657 (N_657,In_1371,In_1804);
and U658 (N_658,In_277,In_1475);
nand U659 (N_659,In_1308,In_185);
xor U660 (N_660,In_1416,In_1610);
xor U661 (N_661,In_556,In_1286);
and U662 (N_662,In_519,In_159);
or U663 (N_663,In_491,In_344);
or U664 (N_664,In_1806,In_35);
nand U665 (N_665,In_1798,In_418);
and U666 (N_666,In_732,In_531);
nor U667 (N_667,In_301,In_1226);
nand U668 (N_668,In_1618,In_197);
and U669 (N_669,In_960,In_1964);
xnor U670 (N_670,In_198,In_49);
nand U671 (N_671,In_1312,In_1961);
and U672 (N_672,In_240,In_86);
xor U673 (N_673,In_411,In_758);
nor U674 (N_674,In_509,In_1748);
nor U675 (N_675,In_410,In_1483);
nand U676 (N_676,In_560,In_1626);
and U677 (N_677,In_512,In_736);
xor U678 (N_678,In_1579,In_1778);
nand U679 (N_679,In_575,In_939);
xor U680 (N_680,In_1575,In_1261);
or U681 (N_681,In_927,In_1496);
nor U682 (N_682,In_1629,In_771);
nor U683 (N_683,In_623,In_803);
or U684 (N_684,In_683,In_590);
nor U685 (N_685,In_515,In_384);
and U686 (N_686,In_1689,In_875);
and U687 (N_687,In_314,In_444);
nand U688 (N_688,In_495,In_1821);
and U689 (N_689,In_1699,In_57);
and U690 (N_690,In_7,In_698);
nand U691 (N_691,In_1662,In_199);
nand U692 (N_692,In_1780,In_1412);
nand U693 (N_693,In_347,In_1456);
nand U694 (N_694,In_337,In_419);
or U695 (N_695,In_399,In_375);
or U696 (N_696,In_263,In_1002);
or U697 (N_697,In_646,In_518);
xnor U698 (N_698,In_1315,In_1409);
nor U699 (N_699,In_305,In_1247);
or U700 (N_700,In_957,In_388);
xor U701 (N_701,In_440,In_806);
xor U702 (N_702,In_740,In_486);
nand U703 (N_703,In_1219,In_551);
nor U704 (N_704,In_487,In_1913);
or U705 (N_705,In_841,In_213);
nand U706 (N_706,In_1698,In_1239);
nor U707 (N_707,In_577,In_373);
or U708 (N_708,In_986,In_433);
nor U709 (N_709,In_1779,In_1860);
or U710 (N_710,In_833,In_878);
nand U711 (N_711,In_1883,In_394);
nand U712 (N_712,In_441,In_366);
nor U713 (N_713,In_603,In_261);
nand U714 (N_714,In_1145,In_1588);
and U715 (N_715,In_1137,In_102);
nor U716 (N_716,In_1244,In_1413);
and U717 (N_717,In_1306,In_1297);
nor U718 (N_718,In_520,In_186);
xnor U719 (N_719,In_525,In_93);
or U720 (N_720,In_201,In_991);
xor U721 (N_721,In_466,In_595);
nor U722 (N_722,In_1388,In_685);
and U723 (N_723,In_1076,In_1082);
xnor U724 (N_724,In_306,In_973);
nand U725 (N_725,In_1518,In_1154);
xor U726 (N_726,In_401,In_1720);
and U727 (N_727,In_492,In_1563);
nand U728 (N_728,In_777,In_1529);
and U729 (N_729,In_1367,In_1120);
or U730 (N_730,In_152,In_945);
and U731 (N_731,In_816,In_1716);
xnor U732 (N_732,In_1420,In_926);
xnor U733 (N_733,In_1836,In_1135);
or U734 (N_734,In_1532,In_1285);
nor U735 (N_735,In_1484,In_745);
nor U736 (N_736,In_899,In_669);
or U737 (N_737,In_323,In_100);
or U738 (N_738,In_54,In_1686);
or U739 (N_739,In_38,In_918);
nand U740 (N_740,In_200,In_20);
and U741 (N_741,In_1214,In_397);
nor U742 (N_742,In_735,In_1603);
nand U743 (N_743,In_1250,In_971);
and U744 (N_744,In_703,In_867);
nand U745 (N_745,In_1,In_338);
xnor U746 (N_746,In_1800,In_1463);
and U747 (N_747,In_1468,In_154);
or U748 (N_748,In_579,In_1853);
or U749 (N_749,In_728,In_248);
nand U750 (N_750,In_615,In_307);
nand U751 (N_751,In_994,In_773);
or U752 (N_752,In_1322,In_1235);
nand U753 (N_753,In_1148,In_1593);
nor U754 (N_754,In_1224,In_950);
and U755 (N_755,In_128,In_1422);
nor U756 (N_756,In_598,In_342);
nor U757 (N_757,In_901,In_1338);
or U758 (N_758,In_1336,In_1971);
nand U759 (N_759,In_1882,In_113);
nor U760 (N_760,In_889,In_981);
xor U761 (N_761,In_1258,In_151);
nand U762 (N_762,In_1839,In_1440);
nor U763 (N_763,In_607,In_585);
nand U764 (N_764,In_737,In_114);
nor U765 (N_765,In_1455,In_1095);
nor U766 (N_766,In_1926,In_894);
xor U767 (N_767,In_1016,In_1762);
xor U768 (N_768,In_1744,In_1846);
or U769 (N_769,In_849,In_1280);
nand U770 (N_770,In_636,In_819);
and U771 (N_771,In_570,In_1321);
and U772 (N_772,In_1538,In_1038);
or U773 (N_773,In_1369,In_866);
nor U774 (N_774,In_658,In_1206);
or U775 (N_775,In_1525,In_1941);
nor U776 (N_776,In_69,In_1252);
or U777 (N_777,In_726,In_224);
nand U778 (N_778,In_1119,In_25);
and U779 (N_779,In_236,In_447);
and U780 (N_780,In_638,In_1898);
and U781 (N_781,In_1382,In_99);
nor U782 (N_782,In_1877,In_1356);
or U783 (N_783,In_1810,In_805);
nand U784 (N_784,In_1173,In_1886);
nor U785 (N_785,In_997,In_1920);
and U786 (N_786,In_897,In_59);
and U787 (N_787,In_1387,In_1372);
or U788 (N_788,In_1094,In_1400);
nor U789 (N_789,In_1967,In_1852);
nor U790 (N_790,In_1176,In_1489);
xnor U791 (N_791,In_589,In_272);
nor U792 (N_792,In_1039,In_318);
xnor U793 (N_793,In_1531,In_1241);
xnor U794 (N_794,In_1062,In_1663);
nor U795 (N_795,In_275,In_1958);
nor U796 (N_796,In_143,In_1693);
and U797 (N_797,In_1596,In_11);
and U798 (N_798,In_1668,In_279);
nor U799 (N_799,In_959,In_218);
nor U800 (N_800,In_80,In_887);
nand U801 (N_801,In_786,In_584);
or U802 (N_802,In_475,In_1263);
and U803 (N_803,In_1576,In_668);
nand U804 (N_804,In_653,In_270);
nor U805 (N_805,In_1198,In_676);
or U806 (N_806,In_1943,In_795);
or U807 (N_807,In_158,In_1659);
and U808 (N_808,In_1209,In_437);
xor U809 (N_809,In_1715,In_588);
nand U810 (N_810,In_1495,In_1072);
nor U811 (N_811,In_193,In_160);
or U812 (N_812,In_1790,In_989);
nand U813 (N_813,In_1521,In_892);
nor U814 (N_814,In_762,In_1394);
nor U815 (N_815,In_567,In_1522);
and U816 (N_816,In_1161,In_572);
nand U817 (N_817,In_1582,In_1634);
or U818 (N_818,In_1444,In_1034);
nand U819 (N_819,In_915,In_1845);
or U820 (N_820,In_265,In_1802);
and U821 (N_821,In_1036,In_309);
and U822 (N_822,In_1587,In_1411);
nand U823 (N_823,In_1982,In_1989);
nor U824 (N_824,In_895,In_1171);
xnor U825 (N_825,In_1745,In_504);
nand U826 (N_826,In_757,In_1185);
nand U827 (N_827,In_1390,In_247);
xor U828 (N_828,In_488,In_181);
and U829 (N_829,In_409,In_132);
nand U830 (N_830,In_1434,In_46);
or U831 (N_831,In_604,In_1078);
nand U832 (N_832,In_715,In_1000);
nor U833 (N_833,In_651,In_847);
nand U834 (N_834,In_1043,In_1581);
or U835 (N_835,In_9,In_1735);
and U836 (N_836,In_1516,In_1479);
or U837 (N_837,In_1736,In_800);
and U838 (N_838,In_965,In_1597);
nor U839 (N_839,In_234,In_221);
or U840 (N_840,In_862,In_948);
nor U841 (N_841,In_353,In_1112);
and U842 (N_842,In_1711,In_566);
nor U843 (N_843,In_1595,In_553);
or U844 (N_844,In_963,In_1542);
nor U845 (N_845,In_290,In_1934);
or U846 (N_846,In_295,In_533);
or U847 (N_847,In_1874,In_1465);
nor U848 (N_848,In_1688,In_1607);
and U849 (N_849,In_1624,In_148);
and U850 (N_850,In_853,In_789);
or U851 (N_851,In_130,In_877);
nand U852 (N_852,In_255,In_1125);
nor U853 (N_853,In_1667,In_1977);
nand U854 (N_854,In_886,In_1935);
or U855 (N_855,In_1007,In_513);
nor U856 (N_856,In_670,In_734);
or U857 (N_857,In_1505,In_230);
nand U858 (N_858,In_1184,In_1374);
nor U859 (N_859,In_406,In_371);
nand U860 (N_860,In_1677,In_269);
and U861 (N_861,In_1377,In_628);
and U862 (N_862,In_1272,In_1660);
xor U863 (N_863,In_1535,In_1270);
nor U864 (N_864,In_396,In_980);
nand U865 (N_865,In_456,In_987);
xnor U866 (N_866,In_1919,In_254);
and U867 (N_867,In_262,In_663);
nand U868 (N_868,In_725,In_1144);
or U869 (N_869,In_1750,In_1143);
and U870 (N_870,In_176,In_74);
nor U871 (N_871,In_681,In_1477);
nand U872 (N_872,In_906,In_507);
or U873 (N_873,In_1021,In_1584);
nand U874 (N_874,In_413,In_1767);
and U875 (N_875,In_1350,In_1851);
nor U876 (N_876,In_898,In_620);
nor U877 (N_877,In_1850,In_1302);
and U878 (N_878,In_1165,In_540);
and U879 (N_879,In_1671,In_782);
xnor U880 (N_880,In_457,In_83);
nor U881 (N_881,In_1418,In_1436);
xnor U882 (N_882,In_405,In_1044);
and U883 (N_883,In_1299,In_637);
nand U884 (N_884,In_1828,In_1921);
and U885 (N_885,In_1770,In_1520);
nand U886 (N_886,In_1497,In_508);
nand U887 (N_887,In_133,In_1160);
nand U888 (N_888,In_459,In_846);
or U889 (N_889,In_1975,In_1620);
nor U890 (N_890,In_1353,In_993);
nor U891 (N_891,In_1233,In_538);
xor U892 (N_892,In_463,In_756);
and U893 (N_893,In_1612,In_345);
nor U894 (N_894,In_1638,In_1583);
and U895 (N_895,In_830,In_1864);
nor U896 (N_896,In_1317,In_1746);
nand U897 (N_897,In_524,In_1549);
nor U898 (N_898,In_1674,In_1445);
nor U899 (N_899,In_1215,In_1323);
or U900 (N_900,In_24,In_731);
or U901 (N_901,In_21,In_1348);
nand U902 (N_902,In_1242,In_1690);
and U903 (N_903,In_357,In_536);
or U904 (N_904,In_1995,In_1147);
or U905 (N_905,In_482,In_931);
nor U906 (N_906,In_77,In_1568);
and U907 (N_907,In_1091,In_1065);
and U908 (N_908,In_1204,In_78);
nor U909 (N_909,In_1208,In_630);
or U910 (N_910,In_801,In_1749);
xnor U911 (N_911,In_1466,In_1869);
or U912 (N_912,In_426,In_1284);
nand U913 (N_913,In_1492,In_535);
nand U914 (N_914,In_473,In_1493);
nand U915 (N_915,In_1751,In_63);
or U916 (N_916,In_1721,In_28);
nand U917 (N_917,In_1992,In_865);
nand U918 (N_918,In_1211,In_183);
or U919 (N_919,In_903,In_391);
or U920 (N_920,In_1175,In_461);
or U921 (N_921,In_879,In_1865);
and U922 (N_922,In_1707,In_1862);
nand U923 (N_923,In_335,In_271);
xnor U924 (N_924,In_977,In_1201);
nor U925 (N_925,In_1672,In_659);
and U926 (N_926,In_1738,In_1359);
xnor U927 (N_927,In_1963,In_1257);
or U928 (N_928,In_1573,In_1131);
and U929 (N_929,In_443,In_1528);
nand U930 (N_930,In_1730,In_326);
and U931 (N_931,In_1183,In_631);
nand U932 (N_932,In_1552,In_702);
nor U933 (N_933,In_664,In_211);
or U934 (N_934,In_174,In_1060);
nand U935 (N_935,In_1830,In_1966);
or U936 (N_936,In_689,In_244);
nor U937 (N_937,In_298,In_1447);
xnor U938 (N_938,In_1457,In_61);
nand U939 (N_939,In_772,In_1225);
nor U940 (N_940,In_421,In_635);
and U941 (N_941,In_1439,In_1229);
nand U942 (N_942,In_1163,In_924);
or U943 (N_943,In_476,In_1304);
nand U944 (N_944,In_908,In_1344);
nand U945 (N_945,In_73,In_1279);
nand U946 (N_946,In_1269,In_1430);
nand U947 (N_947,In_568,In_31);
and U948 (N_948,In_22,In_1932);
xnor U949 (N_949,In_66,In_1194);
nor U950 (N_950,In_542,In_341);
nor U951 (N_951,In_1023,In_146);
or U952 (N_952,In_1630,In_480);
and U953 (N_953,In_1952,In_340);
nor U954 (N_954,In_1968,In_1061);
and U955 (N_955,In_96,In_612);
nand U956 (N_956,In_1714,In_912);
nor U957 (N_957,In_1335,In_633);
nand U958 (N_958,In_1605,In_641);
xnor U959 (N_959,In_1933,In_42);
xor U960 (N_960,In_942,In_1782);
and U961 (N_961,In_934,In_1003);
nor U962 (N_962,In_582,In_1303);
nor U963 (N_963,In_954,In_1015);
or U964 (N_964,In_1844,In_127);
nor U965 (N_965,In_1729,In_1849);
nand U966 (N_966,In_207,In_677);
and U967 (N_967,In_1478,In_1589);
nand U968 (N_968,In_1950,In_600);
nand U969 (N_969,In_1141,In_150);
nand U970 (N_970,In_1190,In_313);
nor U971 (N_971,In_1825,In_34);
nor U972 (N_972,In_1863,In_999);
and U973 (N_973,In_219,In_1234);
and U974 (N_974,In_1398,In_381);
nand U975 (N_975,In_215,In_705);
or U976 (N_976,In_1566,In_1718);
nor U977 (N_977,In_983,In_1133);
nor U978 (N_978,In_727,In_1906);
nor U979 (N_979,In_1158,In_302);
xor U980 (N_980,In_655,In_754);
or U981 (N_981,In_587,In_1019);
or U982 (N_982,In_1905,In_429);
nand U983 (N_983,In_1391,In_693);
xnor U984 (N_984,In_1351,In_1063);
nand U985 (N_985,In_377,In_1132);
nor U986 (N_986,In_1245,In_238);
and U987 (N_987,In_1193,In_170);
xnor U988 (N_988,In_1054,In_701);
nand U989 (N_989,In_1784,In_990);
nor U990 (N_990,In_367,In_1195);
nand U991 (N_991,In_874,In_1130);
nor U992 (N_992,In_678,In_836);
nand U993 (N_993,In_1512,In_1366);
or U994 (N_994,In_1203,In_1704);
or U995 (N_995,In_842,In_917);
and U996 (N_996,In_1045,In_15);
xnor U997 (N_997,In_436,In_1066);
nor U998 (N_998,In_458,In_599);
nand U999 (N_999,In_885,In_1656);
nand U1000 (N_1000,In_633,In_1753);
and U1001 (N_1001,In_445,In_393);
and U1002 (N_1002,In_1782,In_1492);
nor U1003 (N_1003,In_149,In_1152);
nor U1004 (N_1004,In_150,In_674);
nor U1005 (N_1005,In_1945,In_1723);
and U1006 (N_1006,In_1748,In_986);
and U1007 (N_1007,In_1388,In_790);
nor U1008 (N_1008,In_1808,In_44);
nor U1009 (N_1009,In_1213,In_619);
and U1010 (N_1010,In_184,In_820);
and U1011 (N_1011,In_1802,In_1507);
and U1012 (N_1012,In_1216,In_185);
nand U1013 (N_1013,In_1380,In_1264);
nor U1014 (N_1014,In_53,In_1626);
nand U1015 (N_1015,In_1999,In_590);
and U1016 (N_1016,In_617,In_1536);
or U1017 (N_1017,In_1410,In_100);
and U1018 (N_1018,In_1904,In_1849);
nand U1019 (N_1019,In_1166,In_49);
nor U1020 (N_1020,In_1612,In_1080);
nor U1021 (N_1021,In_1563,In_1786);
or U1022 (N_1022,In_204,In_1802);
and U1023 (N_1023,In_1146,In_898);
nand U1024 (N_1024,In_854,In_797);
nand U1025 (N_1025,In_1440,In_856);
and U1026 (N_1026,In_1984,In_447);
nand U1027 (N_1027,In_718,In_271);
or U1028 (N_1028,In_1426,In_423);
nor U1029 (N_1029,In_1817,In_1228);
nand U1030 (N_1030,In_802,In_403);
xnor U1031 (N_1031,In_1124,In_1856);
and U1032 (N_1032,In_1965,In_1017);
nor U1033 (N_1033,In_1663,In_1715);
and U1034 (N_1034,In_1870,In_1191);
and U1035 (N_1035,In_1597,In_306);
or U1036 (N_1036,In_1446,In_1722);
or U1037 (N_1037,In_509,In_68);
nor U1038 (N_1038,In_1951,In_656);
nand U1039 (N_1039,In_1418,In_328);
nor U1040 (N_1040,In_1948,In_1366);
and U1041 (N_1041,In_571,In_777);
nor U1042 (N_1042,In_1315,In_333);
nor U1043 (N_1043,In_742,In_1426);
nor U1044 (N_1044,In_865,In_620);
nand U1045 (N_1045,In_14,In_718);
nand U1046 (N_1046,In_1448,In_1038);
or U1047 (N_1047,In_1122,In_636);
or U1048 (N_1048,In_315,In_1845);
nor U1049 (N_1049,In_1256,In_599);
nor U1050 (N_1050,In_831,In_91);
or U1051 (N_1051,In_700,In_1403);
nor U1052 (N_1052,In_490,In_1865);
nand U1053 (N_1053,In_274,In_516);
or U1054 (N_1054,In_750,In_776);
or U1055 (N_1055,In_62,In_718);
and U1056 (N_1056,In_1538,In_1848);
xor U1057 (N_1057,In_888,In_808);
nand U1058 (N_1058,In_905,In_625);
nor U1059 (N_1059,In_431,In_1842);
nor U1060 (N_1060,In_1381,In_1635);
nor U1061 (N_1061,In_1866,In_613);
or U1062 (N_1062,In_907,In_1327);
nand U1063 (N_1063,In_204,In_141);
and U1064 (N_1064,In_348,In_1434);
nand U1065 (N_1065,In_1795,In_129);
nand U1066 (N_1066,In_1435,In_510);
nor U1067 (N_1067,In_1519,In_1141);
or U1068 (N_1068,In_581,In_327);
or U1069 (N_1069,In_641,In_1254);
nor U1070 (N_1070,In_309,In_1805);
nand U1071 (N_1071,In_1411,In_1872);
or U1072 (N_1072,In_585,In_1004);
and U1073 (N_1073,In_1346,In_1854);
and U1074 (N_1074,In_440,In_1867);
and U1075 (N_1075,In_1527,In_489);
xnor U1076 (N_1076,In_726,In_1659);
or U1077 (N_1077,In_1985,In_574);
nand U1078 (N_1078,In_1024,In_1691);
or U1079 (N_1079,In_1443,In_1119);
nand U1080 (N_1080,In_739,In_617);
xnor U1081 (N_1081,In_1394,In_345);
and U1082 (N_1082,In_587,In_1832);
or U1083 (N_1083,In_1747,In_237);
nor U1084 (N_1084,In_1461,In_1663);
nand U1085 (N_1085,In_894,In_1233);
xor U1086 (N_1086,In_1389,In_537);
nor U1087 (N_1087,In_1688,In_1208);
nor U1088 (N_1088,In_1781,In_919);
nor U1089 (N_1089,In_1413,In_981);
and U1090 (N_1090,In_700,In_656);
nand U1091 (N_1091,In_363,In_1828);
or U1092 (N_1092,In_691,In_1223);
nand U1093 (N_1093,In_1873,In_619);
nor U1094 (N_1094,In_1821,In_392);
nand U1095 (N_1095,In_1826,In_1651);
or U1096 (N_1096,In_116,In_692);
and U1097 (N_1097,In_1085,In_1160);
or U1098 (N_1098,In_1766,In_1578);
or U1099 (N_1099,In_1598,In_870);
or U1100 (N_1100,In_98,In_1668);
or U1101 (N_1101,In_464,In_784);
and U1102 (N_1102,In_46,In_589);
or U1103 (N_1103,In_1662,In_1149);
and U1104 (N_1104,In_732,In_1868);
and U1105 (N_1105,In_446,In_1451);
nand U1106 (N_1106,In_325,In_1623);
or U1107 (N_1107,In_1880,In_1177);
nand U1108 (N_1108,In_241,In_11);
and U1109 (N_1109,In_1978,In_285);
and U1110 (N_1110,In_754,In_25);
nand U1111 (N_1111,In_125,In_1600);
or U1112 (N_1112,In_1859,In_569);
and U1113 (N_1113,In_1853,In_766);
or U1114 (N_1114,In_1446,In_750);
or U1115 (N_1115,In_1902,In_1958);
xor U1116 (N_1116,In_1198,In_323);
and U1117 (N_1117,In_1647,In_1765);
nor U1118 (N_1118,In_1227,In_104);
or U1119 (N_1119,In_1346,In_1545);
nor U1120 (N_1120,In_803,In_905);
and U1121 (N_1121,In_929,In_1971);
or U1122 (N_1122,In_26,In_1860);
and U1123 (N_1123,In_1001,In_798);
or U1124 (N_1124,In_1208,In_1800);
nor U1125 (N_1125,In_145,In_1110);
and U1126 (N_1126,In_1296,In_975);
nand U1127 (N_1127,In_1190,In_1465);
nor U1128 (N_1128,In_1036,In_136);
and U1129 (N_1129,In_205,In_1622);
nor U1130 (N_1130,In_1258,In_1407);
nor U1131 (N_1131,In_1873,In_552);
nor U1132 (N_1132,In_1822,In_1687);
nand U1133 (N_1133,In_790,In_654);
nor U1134 (N_1134,In_1360,In_1072);
nand U1135 (N_1135,In_1575,In_637);
xnor U1136 (N_1136,In_1540,In_1307);
or U1137 (N_1137,In_319,In_1505);
nor U1138 (N_1138,In_1999,In_229);
nor U1139 (N_1139,In_146,In_1997);
or U1140 (N_1140,In_1874,In_645);
and U1141 (N_1141,In_1484,In_1800);
and U1142 (N_1142,In_1059,In_308);
and U1143 (N_1143,In_411,In_178);
and U1144 (N_1144,In_529,In_159);
or U1145 (N_1145,In_1708,In_1260);
nor U1146 (N_1146,In_1526,In_162);
and U1147 (N_1147,In_507,In_1120);
and U1148 (N_1148,In_1117,In_81);
nand U1149 (N_1149,In_934,In_530);
nand U1150 (N_1150,In_560,In_490);
nand U1151 (N_1151,In_884,In_696);
or U1152 (N_1152,In_228,In_1756);
nor U1153 (N_1153,In_1654,In_1857);
and U1154 (N_1154,In_178,In_1431);
or U1155 (N_1155,In_817,In_1110);
nand U1156 (N_1156,In_1885,In_1042);
nor U1157 (N_1157,In_515,In_137);
nand U1158 (N_1158,In_887,In_1371);
nor U1159 (N_1159,In_780,In_593);
nor U1160 (N_1160,In_1693,In_1032);
or U1161 (N_1161,In_1158,In_988);
nand U1162 (N_1162,In_477,In_604);
nand U1163 (N_1163,In_1352,In_597);
nand U1164 (N_1164,In_1,In_1540);
or U1165 (N_1165,In_933,In_1347);
and U1166 (N_1166,In_1240,In_599);
and U1167 (N_1167,In_343,In_1311);
xnor U1168 (N_1168,In_254,In_1222);
nand U1169 (N_1169,In_1422,In_1798);
nand U1170 (N_1170,In_1366,In_990);
or U1171 (N_1171,In_381,In_999);
or U1172 (N_1172,In_886,In_14);
or U1173 (N_1173,In_1458,In_1542);
nand U1174 (N_1174,In_841,In_1292);
and U1175 (N_1175,In_1012,In_1815);
nand U1176 (N_1176,In_766,In_375);
nand U1177 (N_1177,In_579,In_1425);
nor U1178 (N_1178,In_926,In_1969);
nand U1179 (N_1179,In_996,In_1336);
and U1180 (N_1180,In_803,In_131);
xnor U1181 (N_1181,In_1325,In_1795);
nor U1182 (N_1182,In_512,In_527);
and U1183 (N_1183,In_1268,In_379);
nand U1184 (N_1184,In_81,In_1583);
nand U1185 (N_1185,In_1669,In_1088);
nor U1186 (N_1186,In_27,In_744);
or U1187 (N_1187,In_759,In_1799);
or U1188 (N_1188,In_1232,In_970);
and U1189 (N_1189,In_1697,In_170);
nor U1190 (N_1190,In_873,In_732);
and U1191 (N_1191,In_1971,In_474);
and U1192 (N_1192,In_618,In_1457);
nor U1193 (N_1193,In_504,In_509);
nand U1194 (N_1194,In_195,In_1419);
nor U1195 (N_1195,In_1967,In_126);
xor U1196 (N_1196,In_419,In_162);
nand U1197 (N_1197,In_1366,In_398);
and U1198 (N_1198,In_162,In_687);
and U1199 (N_1199,In_1405,In_1966);
or U1200 (N_1200,In_499,In_100);
and U1201 (N_1201,In_303,In_1995);
xor U1202 (N_1202,In_633,In_1441);
xnor U1203 (N_1203,In_1776,In_733);
nand U1204 (N_1204,In_1177,In_1686);
or U1205 (N_1205,In_1972,In_1004);
nor U1206 (N_1206,In_439,In_445);
or U1207 (N_1207,In_268,In_420);
nand U1208 (N_1208,In_979,In_433);
or U1209 (N_1209,In_1384,In_476);
nand U1210 (N_1210,In_237,In_1226);
nand U1211 (N_1211,In_1719,In_332);
nor U1212 (N_1212,In_1175,In_1339);
or U1213 (N_1213,In_1696,In_1490);
nor U1214 (N_1214,In_1552,In_1954);
and U1215 (N_1215,In_1777,In_1582);
xor U1216 (N_1216,In_1209,In_1528);
or U1217 (N_1217,In_519,In_234);
nor U1218 (N_1218,In_1435,In_1253);
and U1219 (N_1219,In_792,In_904);
and U1220 (N_1220,In_1013,In_114);
xor U1221 (N_1221,In_508,In_1764);
nand U1222 (N_1222,In_1966,In_1670);
nand U1223 (N_1223,In_1858,In_389);
nand U1224 (N_1224,In_1691,In_993);
nand U1225 (N_1225,In_944,In_1285);
or U1226 (N_1226,In_799,In_1115);
nor U1227 (N_1227,In_1098,In_899);
and U1228 (N_1228,In_524,In_0);
nor U1229 (N_1229,In_709,In_710);
nor U1230 (N_1230,In_1416,In_1385);
nor U1231 (N_1231,In_1628,In_1953);
nor U1232 (N_1232,In_1064,In_1488);
nor U1233 (N_1233,In_1698,In_59);
xor U1234 (N_1234,In_1520,In_54);
and U1235 (N_1235,In_62,In_1898);
nand U1236 (N_1236,In_247,In_206);
nand U1237 (N_1237,In_1114,In_1103);
or U1238 (N_1238,In_1037,In_1563);
nand U1239 (N_1239,In_1203,In_1833);
or U1240 (N_1240,In_1179,In_364);
nor U1241 (N_1241,In_29,In_729);
and U1242 (N_1242,In_1045,In_575);
nand U1243 (N_1243,In_1571,In_1589);
and U1244 (N_1244,In_1141,In_693);
nand U1245 (N_1245,In_968,In_361);
or U1246 (N_1246,In_1423,In_735);
nand U1247 (N_1247,In_739,In_1848);
and U1248 (N_1248,In_880,In_649);
nor U1249 (N_1249,In_372,In_1953);
nor U1250 (N_1250,In_1756,In_289);
nor U1251 (N_1251,In_1196,In_180);
xnor U1252 (N_1252,In_1255,In_1221);
xnor U1253 (N_1253,In_1939,In_290);
or U1254 (N_1254,In_720,In_742);
xor U1255 (N_1255,In_1864,In_26);
and U1256 (N_1256,In_1588,In_171);
and U1257 (N_1257,In_136,In_1345);
and U1258 (N_1258,In_1384,In_345);
and U1259 (N_1259,In_114,In_1106);
or U1260 (N_1260,In_237,In_1854);
xnor U1261 (N_1261,In_211,In_128);
nor U1262 (N_1262,In_1753,In_715);
nor U1263 (N_1263,In_1376,In_1739);
nor U1264 (N_1264,In_1148,In_75);
nor U1265 (N_1265,In_734,In_7);
nor U1266 (N_1266,In_1391,In_485);
nand U1267 (N_1267,In_1488,In_1629);
nor U1268 (N_1268,In_795,In_1493);
nor U1269 (N_1269,In_1230,In_1640);
nand U1270 (N_1270,In_1361,In_1823);
and U1271 (N_1271,In_1522,In_400);
and U1272 (N_1272,In_1682,In_660);
nor U1273 (N_1273,In_1798,In_783);
xnor U1274 (N_1274,In_728,In_458);
nand U1275 (N_1275,In_146,In_438);
nor U1276 (N_1276,In_660,In_1136);
nand U1277 (N_1277,In_1223,In_28);
nand U1278 (N_1278,In_1519,In_336);
or U1279 (N_1279,In_928,In_483);
nand U1280 (N_1280,In_1204,In_451);
xor U1281 (N_1281,In_1871,In_1878);
or U1282 (N_1282,In_1761,In_1196);
nand U1283 (N_1283,In_1230,In_1669);
nor U1284 (N_1284,In_303,In_882);
and U1285 (N_1285,In_152,In_1400);
nand U1286 (N_1286,In_1541,In_347);
nand U1287 (N_1287,In_243,In_108);
or U1288 (N_1288,In_1296,In_1906);
nor U1289 (N_1289,In_1896,In_340);
or U1290 (N_1290,In_1477,In_1372);
or U1291 (N_1291,In_1702,In_1299);
and U1292 (N_1292,In_248,In_1039);
nor U1293 (N_1293,In_356,In_1471);
nor U1294 (N_1294,In_1644,In_1296);
nor U1295 (N_1295,In_648,In_1946);
nor U1296 (N_1296,In_1676,In_1899);
xnor U1297 (N_1297,In_119,In_1363);
xnor U1298 (N_1298,In_1313,In_560);
and U1299 (N_1299,In_223,In_219);
and U1300 (N_1300,In_962,In_1417);
or U1301 (N_1301,In_1220,In_440);
and U1302 (N_1302,In_1170,In_1797);
nor U1303 (N_1303,In_1300,In_448);
and U1304 (N_1304,In_1006,In_1482);
or U1305 (N_1305,In_13,In_1375);
or U1306 (N_1306,In_174,In_232);
xnor U1307 (N_1307,In_1977,In_453);
or U1308 (N_1308,In_1525,In_52);
nor U1309 (N_1309,In_1289,In_1573);
nand U1310 (N_1310,In_1784,In_1783);
xor U1311 (N_1311,In_1449,In_925);
nand U1312 (N_1312,In_781,In_1912);
and U1313 (N_1313,In_101,In_352);
or U1314 (N_1314,In_849,In_564);
nand U1315 (N_1315,In_451,In_1222);
nor U1316 (N_1316,In_397,In_1385);
nand U1317 (N_1317,In_528,In_602);
and U1318 (N_1318,In_1693,In_771);
nand U1319 (N_1319,In_243,In_938);
nor U1320 (N_1320,In_806,In_299);
nor U1321 (N_1321,In_1965,In_271);
or U1322 (N_1322,In_957,In_831);
nor U1323 (N_1323,In_1191,In_1145);
xnor U1324 (N_1324,In_234,In_1858);
or U1325 (N_1325,In_1461,In_1813);
xnor U1326 (N_1326,In_1826,In_682);
and U1327 (N_1327,In_1126,In_1652);
nand U1328 (N_1328,In_72,In_923);
and U1329 (N_1329,In_1406,In_917);
nand U1330 (N_1330,In_1715,In_1516);
or U1331 (N_1331,In_671,In_1561);
and U1332 (N_1332,In_1023,In_572);
and U1333 (N_1333,In_1362,In_1031);
xor U1334 (N_1334,In_542,In_491);
or U1335 (N_1335,In_523,In_1648);
and U1336 (N_1336,In_1405,In_654);
nand U1337 (N_1337,In_1286,In_975);
nand U1338 (N_1338,In_335,In_1502);
nand U1339 (N_1339,In_1429,In_124);
and U1340 (N_1340,In_1182,In_1682);
and U1341 (N_1341,In_781,In_1819);
nor U1342 (N_1342,In_952,In_1236);
nor U1343 (N_1343,In_482,In_1821);
or U1344 (N_1344,In_829,In_1841);
xor U1345 (N_1345,In_814,In_731);
nor U1346 (N_1346,In_1039,In_711);
and U1347 (N_1347,In_586,In_490);
nand U1348 (N_1348,In_1311,In_619);
or U1349 (N_1349,In_880,In_736);
and U1350 (N_1350,In_390,In_1312);
nor U1351 (N_1351,In_1789,In_1669);
and U1352 (N_1352,In_1549,In_788);
nand U1353 (N_1353,In_1904,In_1238);
nor U1354 (N_1354,In_1613,In_88);
nor U1355 (N_1355,In_343,In_1341);
and U1356 (N_1356,In_96,In_931);
and U1357 (N_1357,In_1751,In_667);
nand U1358 (N_1358,In_1580,In_1150);
or U1359 (N_1359,In_1686,In_1423);
nand U1360 (N_1360,In_1074,In_158);
xor U1361 (N_1361,In_1573,In_1024);
or U1362 (N_1362,In_553,In_1203);
and U1363 (N_1363,In_1975,In_1796);
nor U1364 (N_1364,In_65,In_346);
and U1365 (N_1365,In_846,In_1885);
and U1366 (N_1366,In_722,In_749);
xor U1367 (N_1367,In_1261,In_127);
and U1368 (N_1368,In_784,In_832);
nor U1369 (N_1369,In_608,In_1528);
or U1370 (N_1370,In_752,In_1887);
nor U1371 (N_1371,In_1413,In_1902);
or U1372 (N_1372,In_1814,In_36);
nor U1373 (N_1373,In_284,In_218);
nor U1374 (N_1374,In_1933,In_1482);
nor U1375 (N_1375,In_385,In_466);
or U1376 (N_1376,In_167,In_1400);
nand U1377 (N_1377,In_25,In_780);
nand U1378 (N_1378,In_1915,In_438);
and U1379 (N_1379,In_1018,In_489);
and U1380 (N_1380,In_1569,In_629);
or U1381 (N_1381,In_351,In_224);
nand U1382 (N_1382,In_1568,In_299);
nand U1383 (N_1383,In_598,In_958);
nor U1384 (N_1384,In_1961,In_762);
or U1385 (N_1385,In_1690,In_1970);
nor U1386 (N_1386,In_347,In_189);
or U1387 (N_1387,In_1496,In_255);
or U1388 (N_1388,In_62,In_922);
nor U1389 (N_1389,In_323,In_1655);
and U1390 (N_1390,In_513,In_474);
and U1391 (N_1391,In_171,In_923);
nand U1392 (N_1392,In_1907,In_641);
nor U1393 (N_1393,In_1101,In_1159);
nor U1394 (N_1394,In_903,In_1731);
xnor U1395 (N_1395,In_1948,In_1977);
xnor U1396 (N_1396,In_285,In_195);
nand U1397 (N_1397,In_537,In_1273);
or U1398 (N_1398,In_1167,In_1450);
or U1399 (N_1399,In_701,In_185);
nand U1400 (N_1400,In_1902,In_1938);
or U1401 (N_1401,In_28,In_136);
or U1402 (N_1402,In_1042,In_1254);
nand U1403 (N_1403,In_1741,In_289);
xor U1404 (N_1404,In_116,In_1983);
xor U1405 (N_1405,In_1121,In_1058);
nand U1406 (N_1406,In_1591,In_1896);
or U1407 (N_1407,In_1013,In_753);
nand U1408 (N_1408,In_544,In_357);
and U1409 (N_1409,In_943,In_1817);
xnor U1410 (N_1410,In_528,In_92);
and U1411 (N_1411,In_717,In_1188);
and U1412 (N_1412,In_1037,In_474);
nand U1413 (N_1413,In_275,In_574);
nand U1414 (N_1414,In_1553,In_1120);
nand U1415 (N_1415,In_1584,In_977);
nor U1416 (N_1416,In_526,In_448);
xnor U1417 (N_1417,In_1323,In_255);
nor U1418 (N_1418,In_1097,In_569);
xnor U1419 (N_1419,In_894,In_1167);
and U1420 (N_1420,In_787,In_1976);
xnor U1421 (N_1421,In_1333,In_746);
or U1422 (N_1422,In_773,In_25);
or U1423 (N_1423,In_1751,In_932);
nor U1424 (N_1424,In_1702,In_977);
nand U1425 (N_1425,In_1545,In_263);
or U1426 (N_1426,In_654,In_560);
nand U1427 (N_1427,In_1884,In_1862);
nand U1428 (N_1428,In_1553,In_713);
nand U1429 (N_1429,In_1736,In_90);
xor U1430 (N_1430,In_280,In_1598);
and U1431 (N_1431,In_831,In_1673);
nand U1432 (N_1432,In_193,In_979);
or U1433 (N_1433,In_58,In_1946);
nor U1434 (N_1434,In_1461,In_1582);
nand U1435 (N_1435,In_31,In_938);
or U1436 (N_1436,In_1960,In_121);
nand U1437 (N_1437,In_234,In_1932);
and U1438 (N_1438,In_1231,In_548);
or U1439 (N_1439,In_1126,In_1088);
nor U1440 (N_1440,In_312,In_1131);
or U1441 (N_1441,In_1002,In_308);
and U1442 (N_1442,In_1335,In_1598);
and U1443 (N_1443,In_1184,In_1391);
nand U1444 (N_1444,In_1490,In_1876);
and U1445 (N_1445,In_1902,In_1113);
and U1446 (N_1446,In_1321,In_854);
or U1447 (N_1447,In_72,In_507);
nor U1448 (N_1448,In_1089,In_125);
or U1449 (N_1449,In_806,In_827);
nor U1450 (N_1450,In_1327,In_1042);
or U1451 (N_1451,In_1800,In_483);
or U1452 (N_1452,In_1334,In_1273);
and U1453 (N_1453,In_1145,In_367);
or U1454 (N_1454,In_75,In_88);
xnor U1455 (N_1455,In_1534,In_693);
nand U1456 (N_1456,In_1788,In_1550);
or U1457 (N_1457,In_1828,In_239);
nor U1458 (N_1458,In_1560,In_1353);
and U1459 (N_1459,In_1402,In_888);
and U1460 (N_1460,In_285,In_1454);
xor U1461 (N_1461,In_737,In_1543);
xnor U1462 (N_1462,In_448,In_105);
and U1463 (N_1463,In_122,In_843);
xor U1464 (N_1464,In_1841,In_1147);
nand U1465 (N_1465,In_74,In_1586);
xnor U1466 (N_1466,In_557,In_1743);
nor U1467 (N_1467,In_333,In_1074);
nand U1468 (N_1468,In_1337,In_255);
and U1469 (N_1469,In_58,In_1339);
nor U1470 (N_1470,In_1683,In_475);
nor U1471 (N_1471,In_44,In_642);
nand U1472 (N_1472,In_426,In_270);
or U1473 (N_1473,In_1627,In_542);
or U1474 (N_1474,In_459,In_1194);
nor U1475 (N_1475,In_327,In_1324);
or U1476 (N_1476,In_1247,In_211);
xnor U1477 (N_1477,In_1438,In_1845);
nor U1478 (N_1478,In_698,In_287);
nor U1479 (N_1479,In_177,In_389);
and U1480 (N_1480,In_841,In_730);
and U1481 (N_1481,In_414,In_124);
and U1482 (N_1482,In_325,In_779);
nor U1483 (N_1483,In_56,In_753);
nand U1484 (N_1484,In_138,In_1310);
and U1485 (N_1485,In_965,In_1136);
nand U1486 (N_1486,In_77,In_1851);
nor U1487 (N_1487,In_1116,In_326);
nor U1488 (N_1488,In_262,In_1981);
or U1489 (N_1489,In_1910,In_1410);
or U1490 (N_1490,In_389,In_59);
or U1491 (N_1491,In_648,In_1146);
or U1492 (N_1492,In_1656,In_301);
and U1493 (N_1493,In_66,In_708);
and U1494 (N_1494,In_1003,In_798);
nand U1495 (N_1495,In_891,In_1001);
nor U1496 (N_1496,In_346,In_234);
nor U1497 (N_1497,In_1736,In_1458);
nand U1498 (N_1498,In_435,In_1908);
nand U1499 (N_1499,In_208,In_1335);
and U1500 (N_1500,In_1687,In_627);
nor U1501 (N_1501,In_404,In_1029);
or U1502 (N_1502,In_432,In_1095);
nand U1503 (N_1503,In_915,In_579);
and U1504 (N_1504,In_887,In_520);
or U1505 (N_1505,In_1569,In_113);
nor U1506 (N_1506,In_1582,In_151);
nor U1507 (N_1507,In_1724,In_416);
and U1508 (N_1508,In_1196,In_351);
and U1509 (N_1509,In_324,In_1474);
nor U1510 (N_1510,In_1577,In_1816);
and U1511 (N_1511,In_33,In_496);
or U1512 (N_1512,In_887,In_17);
nor U1513 (N_1513,In_1335,In_1180);
nor U1514 (N_1514,In_324,In_917);
nand U1515 (N_1515,In_437,In_1084);
and U1516 (N_1516,In_1447,In_1698);
nor U1517 (N_1517,In_1317,In_864);
and U1518 (N_1518,In_1457,In_1772);
and U1519 (N_1519,In_252,In_765);
and U1520 (N_1520,In_1226,In_1996);
nand U1521 (N_1521,In_669,In_12);
nand U1522 (N_1522,In_349,In_1458);
nor U1523 (N_1523,In_877,In_1723);
and U1524 (N_1524,In_133,In_898);
and U1525 (N_1525,In_850,In_1280);
nor U1526 (N_1526,In_1219,In_365);
xnor U1527 (N_1527,In_1324,In_1109);
and U1528 (N_1528,In_1556,In_386);
nor U1529 (N_1529,In_248,In_353);
or U1530 (N_1530,In_1941,In_1251);
nor U1531 (N_1531,In_453,In_1076);
nand U1532 (N_1532,In_460,In_433);
or U1533 (N_1533,In_1830,In_1610);
and U1534 (N_1534,In_799,In_858);
nor U1535 (N_1535,In_1048,In_961);
or U1536 (N_1536,In_1189,In_92);
and U1537 (N_1537,In_1668,In_311);
or U1538 (N_1538,In_1251,In_214);
and U1539 (N_1539,In_1981,In_1205);
xor U1540 (N_1540,In_196,In_1220);
nor U1541 (N_1541,In_916,In_1396);
and U1542 (N_1542,In_646,In_1757);
or U1543 (N_1543,In_1565,In_1184);
or U1544 (N_1544,In_234,In_224);
nor U1545 (N_1545,In_1082,In_1773);
xnor U1546 (N_1546,In_501,In_1317);
or U1547 (N_1547,In_1331,In_1083);
nor U1548 (N_1548,In_466,In_1172);
nor U1549 (N_1549,In_312,In_1982);
nor U1550 (N_1550,In_8,In_784);
nor U1551 (N_1551,In_1917,In_1256);
nand U1552 (N_1552,In_273,In_887);
nor U1553 (N_1553,In_1632,In_746);
nor U1554 (N_1554,In_1716,In_386);
and U1555 (N_1555,In_1714,In_1770);
nor U1556 (N_1556,In_1963,In_1250);
nor U1557 (N_1557,In_945,In_517);
or U1558 (N_1558,In_57,In_663);
or U1559 (N_1559,In_1432,In_216);
and U1560 (N_1560,In_237,In_1384);
nand U1561 (N_1561,In_1644,In_268);
or U1562 (N_1562,In_488,In_1721);
nand U1563 (N_1563,In_1511,In_59);
nor U1564 (N_1564,In_1225,In_557);
nor U1565 (N_1565,In_1500,In_1773);
or U1566 (N_1566,In_736,In_1079);
or U1567 (N_1567,In_905,In_1585);
or U1568 (N_1568,In_754,In_845);
nand U1569 (N_1569,In_715,In_704);
and U1570 (N_1570,In_1238,In_1748);
and U1571 (N_1571,In_429,In_583);
and U1572 (N_1572,In_638,In_1433);
or U1573 (N_1573,In_1663,In_1025);
nand U1574 (N_1574,In_115,In_1680);
and U1575 (N_1575,In_1761,In_1356);
or U1576 (N_1576,In_1381,In_54);
nor U1577 (N_1577,In_346,In_82);
nand U1578 (N_1578,In_616,In_1867);
nand U1579 (N_1579,In_1319,In_1813);
or U1580 (N_1580,In_1269,In_1457);
nor U1581 (N_1581,In_598,In_1503);
nand U1582 (N_1582,In_898,In_582);
and U1583 (N_1583,In_795,In_1105);
nor U1584 (N_1584,In_725,In_1266);
and U1585 (N_1585,In_54,In_1460);
xnor U1586 (N_1586,In_1249,In_1473);
or U1587 (N_1587,In_1512,In_164);
nand U1588 (N_1588,In_350,In_430);
and U1589 (N_1589,In_233,In_1405);
nor U1590 (N_1590,In_767,In_1053);
and U1591 (N_1591,In_422,In_100);
and U1592 (N_1592,In_1651,In_208);
nand U1593 (N_1593,In_957,In_1291);
or U1594 (N_1594,In_1899,In_329);
nor U1595 (N_1595,In_74,In_1929);
and U1596 (N_1596,In_204,In_562);
or U1597 (N_1597,In_1111,In_1021);
xnor U1598 (N_1598,In_1962,In_389);
nand U1599 (N_1599,In_1265,In_1750);
or U1600 (N_1600,In_468,In_1260);
nor U1601 (N_1601,In_654,In_750);
and U1602 (N_1602,In_598,In_663);
or U1603 (N_1603,In_1414,In_1851);
and U1604 (N_1604,In_1563,In_54);
nand U1605 (N_1605,In_292,In_793);
nand U1606 (N_1606,In_1269,In_1364);
nand U1607 (N_1607,In_185,In_1752);
nor U1608 (N_1608,In_1901,In_1256);
or U1609 (N_1609,In_1880,In_1072);
nand U1610 (N_1610,In_26,In_805);
or U1611 (N_1611,In_916,In_1718);
nand U1612 (N_1612,In_710,In_1685);
xnor U1613 (N_1613,In_1298,In_877);
nor U1614 (N_1614,In_1912,In_1014);
nor U1615 (N_1615,In_1626,In_673);
and U1616 (N_1616,In_260,In_1923);
and U1617 (N_1617,In_1847,In_1983);
nor U1618 (N_1618,In_28,In_534);
nor U1619 (N_1619,In_95,In_803);
and U1620 (N_1620,In_929,In_1572);
nand U1621 (N_1621,In_643,In_1712);
or U1622 (N_1622,In_1432,In_1220);
nand U1623 (N_1623,In_870,In_1459);
nand U1624 (N_1624,In_249,In_830);
xnor U1625 (N_1625,In_353,In_1957);
nor U1626 (N_1626,In_1710,In_758);
nor U1627 (N_1627,In_1398,In_818);
nand U1628 (N_1628,In_332,In_1338);
nor U1629 (N_1629,In_1004,In_1186);
xnor U1630 (N_1630,In_889,In_937);
and U1631 (N_1631,In_1016,In_1567);
and U1632 (N_1632,In_735,In_703);
nand U1633 (N_1633,In_1586,In_1973);
and U1634 (N_1634,In_151,In_1043);
and U1635 (N_1635,In_430,In_1982);
nand U1636 (N_1636,In_587,In_248);
or U1637 (N_1637,In_307,In_1503);
nand U1638 (N_1638,In_1920,In_1816);
nand U1639 (N_1639,In_12,In_696);
nand U1640 (N_1640,In_1685,In_292);
nand U1641 (N_1641,In_551,In_792);
and U1642 (N_1642,In_150,In_1252);
nand U1643 (N_1643,In_938,In_1184);
nand U1644 (N_1644,In_224,In_883);
or U1645 (N_1645,In_1600,In_1852);
nor U1646 (N_1646,In_603,In_25);
nor U1647 (N_1647,In_825,In_686);
or U1648 (N_1648,In_792,In_81);
nand U1649 (N_1649,In_1957,In_1255);
or U1650 (N_1650,In_731,In_1101);
or U1651 (N_1651,In_767,In_592);
nor U1652 (N_1652,In_1688,In_175);
or U1653 (N_1653,In_1491,In_1725);
or U1654 (N_1654,In_1492,In_1123);
and U1655 (N_1655,In_1458,In_101);
or U1656 (N_1656,In_507,In_1858);
and U1657 (N_1657,In_13,In_1741);
or U1658 (N_1658,In_1069,In_490);
nor U1659 (N_1659,In_139,In_589);
xnor U1660 (N_1660,In_1750,In_638);
nor U1661 (N_1661,In_1839,In_612);
and U1662 (N_1662,In_1516,In_110);
xnor U1663 (N_1663,In_1685,In_1276);
or U1664 (N_1664,In_1012,In_1335);
nand U1665 (N_1665,In_679,In_820);
nor U1666 (N_1666,In_293,In_1786);
or U1667 (N_1667,In_1746,In_1008);
and U1668 (N_1668,In_657,In_714);
nand U1669 (N_1669,In_997,In_391);
or U1670 (N_1670,In_443,In_1143);
and U1671 (N_1671,In_343,In_381);
or U1672 (N_1672,In_885,In_1909);
nor U1673 (N_1673,In_607,In_609);
or U1674 (N_1674,In_1581,In_919);
nor U1675 (N_1675,In_1407,In_1003);
or U1676 (N_1676,In_206,In_1188);
or U1677 (N_1677,In_560,In_1564);
nand U1678 (N_1678,In_190,In_1501);
and U1679 (N_1679,In_211,In_1096);
or U1680 (N_1680,In_1557,In_788);
and U1681 (N_1681,In_296,In_1700);
xnor U1682 (N_1682,In_716,In_1007);
nand U1683 (N_1683,In_94,In_646);
nand U1684 (N_1684,In_256,In_1755);
nor U1685 (N_1685,In_1208,In_1951);
and U1686 (N_1686,In_533,In_1009);
nand U1687 (N_1687,In_552,In_1018);
nor U1688 (N_1688,In_1597,In_663);
or U1689 (N_1689,In_1572,In_80);
or U1690 (N_1690,In_1766,In_117);
nor U1691 (N_1691,In_502,In_480);
nor U1692 (N_1692,In_1511,In_851);
or U1693 (N_1693,In_1411,In_1974);
nor U1694 (N_1694,In_314,In_1581);
nand U1695 (N_1695,In_1054,In_66);
xnor U1696 (N_1696,In_1914,In_1064);
nand U1697 (N_1697,In_293,In_193);
nor U1698 (N_1698,In_314,In_1741);
nor U1699 (N_1699,In_1305,In_1085);
xor U1700 (N_1700,In_316,In_832);
or U1701 (N_1701,In_604,In_110);
or U1702 (N_1702,In_1322,In_410);
nor U1703 (N_1703,In_134,In_1100);
nand U1704 (N_1704,In_1519,In_579);
nand U1705 (N_1705,In_236,In_222);
xnor U1706 (N_1706,In_532,In_973);
or U1707 (N_1707,In_1856,In_412);
and U1708 (N_1708,In_1039,In_1717);
and U1709 (N_1709,In_1649,In_1973);
or U1710 (N_1710,In_399,In_824);
nand U1711 (N_1711,In_1687,In_91);
xnor U1712 (N_1712,In_285,In_54);
nor U1713 (N_1713,In_1292,In_1067);
and U1714 (N_1714,In_1885,In_1499);
or U1715 (N_1715,In_1627,In_1129);
nor U1716 (N_1716,In_1312,In_1466);
nor U1717 (N_1717,In_1949,In_338);
and U1718 (N_1718,In_1792,In_1451);
nor U1719 (N_1719,In_873,In_1000);
or U1720 (N_1720,In_1517,In_391);
and U1721 (N_1721,In_1322,In_423);
nor U1722 (N_1722,In_1029,In_141);
nor U1723 (N_1723,In_143,In_1279);
nor U1724 (N_1724,In_798,In_983);
or U1725 (N_1725,In_234,In_130);
nand U1726 (N_1726,In_1449,In_1582);
nor U1727 (N_1727,In_731,In_701);
nand U1728 (N_1728,In_807,In_1760);
nand U1729 (N_1729,In_1431,In_307);
nand U1730 (N_1730,In_1201,In_723);
nand U1731 (N_1731,In_1243,In_95);
and U1732 (N_1732,In_1705,In_1679);
nor U1733 (N_1733,In_1962,In_707);
nand U1734 (N_1734,In_1199,In_474);
and U1735 (N_1735,In_1035,In_1144);
or U1736 (N_1736,In_897,In_953);
nor U1737 (N_1737,In_1174,In_647);
nand U1738 (N_1738,In_842,In_1810);
nor U1739 (N_1739,In_1968,In_840);
or U1740 (N_1740,In_269,In_50);
and U1741 (N_1741,In_1512,In_870);
and U1742 (N_1742,In_117,In_338);
or U1743 (N_1743,In_1872,In_1998);
and U1744 (N_1744,In_57,In_872);
nor U1745 (N_1745,In_106,In_1905);
nor U1746 (N_1746,In_1594,In_1195);
nand U1747 (N_1747,In_190,In_1058);
nor U1748 (N_1748,In_1253,In_940);
and U1749 (N_1749,In_1226,In_1242);
or U1750 (N_1750,In_455,In_124);
and U1751 (N_1751,In_856,In_1567);
or U1752 (N_1752,In_824,In_1820);
nor U1753 (N_1753,In_776,In_1954);
nor U1754 (N_1754,In_1385,In_1462);
and U1755 (N_1755,In_687,In_1819);
nand U1756 (N_1756,In_1552,In_1332);
and U1757 (N_1757,In_1282,In_1706);
and U1758 (N_1758,In_283,In_713);
nor U1759 (N_1759,In_1741,In_504);
nor U1760 (N_1760,In_208,In_1588);
nand U1761 (N_1761,In_399,In_393);
nand U1762 (N_1762,In_322,In_995);
or U1763 (N_1763,In_1381,In_156);
nand U1764 (N_1764,In_308,In_1952);
and U1765 (N_1765,In_823,In_1453);
xor U1766 (N_1766,In_1368,In_349);
xnor U1767 (N_1767,In_1230,In_212);
nor U1768 (N_1768,In_1439,In_76);
or U1769 (N_1769,In_374,In_1625);
xnor U1770 (N_1770,In_1354,In_165);
xnor U1771 (N_1771,In_482,In_1938);
nor U1772 (N_1772,In_912,In_92);
or U1773 (N_1773,In_369,In_1967);
nor U1774 (N_1774,In_1414,In_1890);
or U1775 (N_1775,In_1302,In_1394);
or U1776 (N_1776,In_1774,In_981);
and U1777 (N_1777,In_1274,In_1162);
and U1778 (N_1778,In_1517,In_1008);
or U1779 (N_1779,In_1144,In_1899);
xor U1780 (N_1780,In_1728,In_1658);
or U1781 (N_1781,In_162,In_1157);
or U1782 (N_1782,In_586,In_1437);
nor U1783 (N_1783,In_1747,In_1337);
nand U1784 (N_1784,In_472,In_558);
nor U1785 (N_1785,In_344,In_1932);
or U1786 (N_1786,In_1905,In_1310);
and U1787 (N_1787,In_1231,In_1508);
nand U1788 (N_1788,In_157,In_877);
or U1789 (N_1789,In_115,In_1955);
nand U1790 (N_1790,In_1680,In_620);
nor U1791 (N_1791,In_328,In_1529);
nand U1792 (N_1792,In_344,In_987);
and U1793 (N_1793,In_833,In_1039);
and U1794 (N_1794,In_982,In_1857);
or U1795 (N_1795,In_1971,In_1333);
and U1796 (N_1796,In_1262,In_1270);
and U1797 (N_1797,In_1928,In_294);
or U1798 (N_1798,In_941,In_1409);
and U1799 (N_1799,In_1099,In_1097);
and U1800 (N_1800,In_184,In_609);
and U1801 (N_1801,In_1763,In_1823);
or U1802 (N_1802,In_1718,In_611);
and U1803 (N_1803,In_517,In_1959);
and U1804 (N_1804,In_1323,In_1146);
nor U1805 (N_1805,In_391,In_508);
nand U1806 (N_1806,In_1934,In_1972);
nand U1807 (N_1807,In_1190,In_890);
nor U1808 (N_1808,In_779,In_1624);
or U1809 (N_1809,In_1237,In_130);
or U1810 (N_1810,In_875,In_1515);
or U1811 (N_1811,In_1136,In_1107);
nor U1812 (N_1812,In_284,In_353);
nor U1813 (N_1813,In_1929,In_1722);
and U1814 (N_1814,In_1900,In_764);
and U1815 (N_1815,In_1016,In_1878);
xnor U1816 (N_1816,In_1930,In_1068);
or U1817 (N_1817,In_289,In_12);
and U1818 (N_1818,In_1702,In_1822);
and U1819 (N_1819,In_930,In_168);
nand U1820 (N_1820,In_119,In_684);
nor U1821 (N_1821,In_600,In_462);
nor U1822 (N_1822,In_944,In_1581);
or U1823 (N_1823,In_1639,In_615);
and U1824 (N_1824,In_1237,In_245);
or U1825 (N_1825,In_348,In_71);
xnor U1826 (N_1826,In_1921,In_1166);
or U1827 (N_1827,In_879,In_712);
nor U1828 (N_1828,In_1629,In_110);
or U1829 (N_1829,In_1303,In_1972);
and U1830 (N_1830,In_70,In_1677);
nand U1831 (N_1831,In_949,In_627);
or U1832 (N_1832,In_465,In_47);
nor U1833 (N_1833,In_1834,In_1309);
nor U1834 (N_1834,In_349,In_421);
xnor U1835 (N_1835,In_457,In_1617);
xnor U1836 (N_1836,In_1987,In_661);
xor U1837 (N_1837,In_626,In_1852);
or U1838 (N_1838,In_1780,In_795);
or U1839 (N_1839,In_918,In_44);
nand U1840 (N_1840,In_974,In_1896);
and U1841 (N_1841,In_197,In_81);
nand U1842 (N_1842,In_1526,In_1851);
xnor U1843 (N_1843,In_1604,In_499);
and U1844 (N_1844,In_1292,In_162);
nor U1845 (N_1845,In_1683,In_1147);
nand U1846 (N_1846,In_388,In_1017);
nand U1847 (N_1847,In_1690,In_999);
and U1848 (N_1848,In_1814,In_1810);
and U1849 (N_1849,In_1026,In_243);
or U1850 (N_1850,In_463,In_239);
nor U1851 (N_1851,In_57,In_1706);
or U1852 (N_1852,In_1038,In_909);
or U1853 (N_1853,In_1985,In_831);
nand U1854 (N_1854,In_180,In_1477);
or U1855 (N_1855,In_840,In_402);
nor U1856 (N_1856,In_1264,In_1034);
nand U1857 (N_1857,In_1281,In_1403);
nor U1858 (N_1858,In_186,In_1482);
nor U1859 (N_1859,In_1413,In_954);
xnor U1860 (N_1860,In_1440,In_1594);
or U1861 (N_1861,In_1226,In_903);
nor U1862 (N_1862,In_239,In_516);
or U1863 (N_1863,In_1336,In_526);
and U1864 (N_1864,In_1344,In_1153);
nor U1865 (N_1865,In_1297,In_1430);
nand U1866 (N_1866,In_1667,In_17);
or U1867 (N_1867,In_1147,In_1216);
or U1868 (N_1868,In_1994,In_1475);
and U1869 (N_1869,In_786,In_1698);
nand U1870 (N_1870,In_1264,In_274);
xor U1871 (N_1871,In_985,In_1825);
nor U1872 (N_1872,In_912,In_821);
nor U1873 (N_1873,In_1935,In_523);
and U1874 (N_1874,In_602,In_1170);
or U1875 (N_1875,In_410,In_174);
or U1876 (N_1876,In_520,In_604);
and U1877 (N_1877,In_812,In_1229);
and U1878 (N_1878,In_438,In_861);
and U1879 (N_1879,In_1009,In_88);
and U1880 (N_1880,In_1257,In_822);
nand U1881 (N_1881,In_1814,In_53);
and U1882 (N_1882,In_1363,In_1310);
nor U1883 (N_1883,In_554,In_1269);
and U1884 (N_1884,In_127,In_894);
nor U1885 (N_1885,In_370,In_1739);
nor U1886 (N_1886,In_556,In_576);
and U1887 (N_1887,In_1068,In_1874);
nand U1888 (N_1888,In_1318,In_48);
nor U1889 (N_1889,In_1010,In_1317);
nor U1890 (N_1890,In_1181,In_633);
and U1891 (N_1891,In_387,In_350);
nand U1892 (N_1892,In_1629,In_1361);
nor U1893 (N_1893,In_444,In_107);
xor U1894 (N_1894,In_1541,In_797);
xor U1895 (N_1895,In_445,In_930);
or U1896 (N_1896,In_425,In_1511);
nor U1897 (N_1897,In_1117,In_304);
or U1898 (N_1898,In_1992,In_959);
and U1899 (N_1899,In_540,In_1837);
nor U1900 (N_1900,In_183,In_1578);
or U1901 (N_1901,In_738,In_739);
nor U1902 (N_1902,In_297,In_1159);
or U1903 (N_1903,In_1875,In_1061);
and U1904 (N_1904,In_1162,In_1585);
and U1905 (N_1905,In_1331,In_1093);
or U1906 (N_1906,In_168,In_1541);
xor U1907 (N_1907,In_669,In_236);
nor U1908 (N_1908,In_939,In_5);
or U1909 (N_1909,In_883,In_846);
nor U1910 (N_1910,In_440,In_185);
nand U1911 (N_1911,In_1236,In_6);
xnor U1912 (N_1912,In_1045,In_461);
or U1913 (N_1913,In_745,In_1400);
and U1914 (N_1914,In_802,In_1418);
or U1915 (N_1915,In_1410,In_53);
nand U1916 (N_1916,In_1534,In_1237);
nand U1917 (N_1917,In_1464,In_1098);
and U1918 (N_1918,In_1678,In_507);
or U1919 (N_1919,In_333,In_1116);
or U1920 (N_1920,In_1582,In_1930);
and U1921 (N_1921,In_1270,In_350);
and U1922 (N_1922,In_56,In_1646);
nor U1923 (N_1923,In_498,In_1727);
or U1924 (N_1924,In_1562,In_785);
nand U1925 (N_1925,In_473,In_1261);
and U1926 (N_1926,In_33,In_1561);
nor U1927 (N_1927,In_438,In_1885);
or U1928 (N_1928,In_468,In_278);
and U1929 (N_1929,In_1398,In_225);
nor U1930 (N_1930,In_1872,In_166);
nor U1931 (N_1931,In_1499,In_912);
nand U1932 (N_1932,In_1192,In_31);
or U1933 (N_1933,In_594,In_1704);
or U1934 (N_1934,In_1498,In_1463);
nor U1935 (N_1935,In_1402,In_604);
nand U1936 (N_1936,In_673,In_40);
and U1937 (N_1937,In_1019,In_1273);
nand U1938 (N_1938,In_891,In_1358);
nand U1939 (N_1939,In_795,In_743);
nand U1940 (N_1940,In_783,In_428);
or U1941 (N_1941,In_1496,In_1685);
or U1942 (N_1942,In_618,In_863);
nand U1943 (N_1943,In_376,In_975);
and U1944 (N_1944,In_1773,In_1109);
or U1945 (N_1945,In_1649,In_305);
xor U1946 (N_1946,In_60,In_1208);
or U1947 (N_1947,In_929,In_1644);
nor U1948 (N_1948,In_42,In_953);
and U1949 (N_1949,In_73,In_534);
nand U1950 (N_1950,In_392,In_1108);
xor U1951 (N_1951,In_1656,In_173);
or U1952 (N_1952,In_907,In_597);
nand U1953 (N_1953,In_1319,In_1861);
or U1954 (N_1954,In_1235,In_1971);
xor U1955 (N_1955,In_1080,In_841);
nor U1956 (N_1956,In_1567,In_818);
or U1957 (N_1957,In_1514,In_901);
or U1958 (N_1958,In_899,In_680);
or U1959 (N_1959,In_1644,In_1625);
or U1960 (N_1960,In_97,In_1903);
xnor U1961 (N_1961,In_1461,In_867);
nor U1962 (N_1962,In_365,In_458);
xor U1963 (N_1963,In_108,In_1560);
and U1964 (N_1964,In_544,In_1130);
and U1965 (N_1965,In_1955,In_1536);
and U1966 (N_1966,In_1844,In_1352);
nor U1967 (N_1967,In_1783,In_1615);
or U1968 (N_1968,In_15,In_958);
nand U1969 (N_1969,In_1845,In_1004);
nor U1970 (N_1970,In_691,In_5);
nor U1971 (N_1971,In_1529,In_1987);
nor U1972 (N_1972,In_1496,In_271);
nand U1973 (N_1973,In_1037,In_1289);
nand U1974 (N_1974,In_65,In_445);
nor U1975 (N_1975,In_59,In_1800);
or U1976 (N_1976,In_473,In_58);
xnor U1977 (N_1977,In_446,In_1420);
or U1978 (N_1978,In_1109,In_796);
or U1979 (N_1979,In_79,In_1887);
nor U1980 (N_1980,In_404,In_756);
or U1981 (N_1981,In_1858,In_387);
or U1982 (N_1982,In_1912,In_1106);
nor U1983 (N_1983,In_609,In_1873);
or U1984 (N_1984,In_1074,In_9);
xnor U1985 (N_1985,In_1245,In_1011);
nand U1986 (N_1986,In_1743,In_1186);
and U1987 (N_1987,In_1225,In_619);
nand U1988 (N_1988,In_352,In_1921);
or U1989 (N_1989,In_535,In_1925);
nand U1990 (N_1990,In_1336,In_1799);
or U1991 (N_1991,In_719,In_157);
nor U1992 (N_1992,In_742,In_1376);
nor U1993 (N_1993,In_259,In_180);
xnor U1994 (N_1994,In_407,In_1539);
nor U1995 (N_1995,In_1835,In_1679);
nand U1996 (N_1996,In_1336,In_1125);
and U1997 (N_1997,In_1433,In_105);
and U1998 (N_1998,In_1119,In_1647);
nor U1999 (N_1999,In_709,In_1059);
xor U2000 (N_2000,In_1768,In_1628);
xor U2001 (N_2001,In_1365,In_376);
and U2002 (N_2002,In_1282,In_786);
or U2003 (N_2003,In_41,In_637);
nand U2004 (N_2004,In_1070,In_1230);
or U2005 (N_2005,In_886,In_505);
and U2006 (N_2006,In_1176,In_927);
nor U2007 (N_2007,In_989,In_1436);
and U2008 (N_2008,In_954,In_1914);
or U2009 (N_2009,In_49,In_1424);
nand U2010 (N_2010,In_1572,In_1763);
and U2011 (N_2011,In_387,In_951);
or U2012 (N_2012,In_947,In_286);
nor U2013 (N_2013,In_199,In_455);
nor U2014 (N_2014,In_1233,In_1490);
and U2015 (N_2015,In_988,In_1572);
nor U2016 (N_2016,In_450,In_1261);
nor U2017 (N_2017,In_1689,In_537);
nand U2018 (N_2018,In_1433,In_569);
nand U2019 (N_2019,In_1591,In_878);
nor U2020 (N_2020,In_1406,In_548);
nor U2021 (N_2021,In_106,In_1281);
nor U2022 (N_2022,In_1611,In_878);
nor U2023 (N_2023,In_251,In_1204);
xor U2024 (N_2024,In_1736,In_1623);
or U2025 (N_2025,In_128,In_1543);
nand U2026 (N_2026,In_483,In_1801);
nor U2027 (N_2027,In_1836,In_353);
and U2028 (N_2028,In_1944,In_1605);
nand U2029 (N_2029,In_1411,In_104);
or U2030 (N_2030,In_60,In_1878);
or U2031 (N_2031,In_1360,In_1116);
and U2032 (N_2032,In_1727,In_1265);
and U2033 (N_2033,In_500,In_1463);
nand U2034 (N_2034,In_1010,In_804);
or U2035 (N_2035,In_1520,In_631);
xnor U2036 (N_2036,In_1507,In_1828);
xnor U2037 (N_2037,In_660,In_1045);
or U2038 (N_2038,In_1046,In_512);
xor U2039 (N_2039,In_1457,In_1424);
nand U2040 (N_2040,In_95,In_283);
and U2041 (N_2041,In_225,In_1177);
nor U2042 (N_2042,In_74,In_1521);
or U2043 (N_2043,In_974,In_1464);
and U2044 (N_2044,In_934,In_1560);
and U2045 (N_2045,In_1891,In_602);
and U2046 (N_2046,In_1723,In_1560);
or U2047 (N_2047,In_1789,In_1995);
or U2048 (N_2048,In_1730,In_187);
or U2049 (N_2049,In_665,In_151);
or U2050 (N_2050,In_336,In_18);
and U2051 (N_2051,In_798,In_909);
or U2052 (N_2052,In_1285,In_608);
and U2053 (N_2053,In_550,In_1085);
nor U2054 (N_2054,In_555,In_284);
nor U2055 (N_2055,In_1317,In_931);
xor U2056 (N_2056,In_1797,In_1780);
xor U2057 (N_2057,In_224,In_1072);
nor U2058 (N_2058,In_1131,In_1870);
and U2059 (N_2059,In_713,In_1984);
and U2060 (N_2060,In_161,In_1324);
nor U2061 (N_2061,In_646,In_35);
nor U2062 (N_2062,In_6,In_1343);
xor U2063 (N_2063,In_1958,In_1082);
and U2064 (N_2064,In_1766,In_387);
xnor U2065 (N_2065,In_1659,In_1262);
nor U2066 (N_2066,In_376,In_438);
nor U2067 (N_2067,In_1571,In_926);
xnor U2068 (N_2068,In_1373,In_1876);
and U2069 (N_2069,In_465,In_361);
xnor U2070 (N_2070,In_283,In_1264);
and U2071 (N_2071,In_915,In_1211);
or U2072 (N_2072,In_1874,In_1173);
and U2073 (N_2073,In_812,In_1441);
or U2074 (N_2074,In_1455,In_1260);
nand U2075 (N_2075,In_1183,In_1503);
and U2076 (N_2076,In_747,In_1304);
nand U2077 (N_2077,In_404,In_1958);
nand U2078 (N_2078,In_1443,In_489);
nor U2079 (N_2079,In_1340,In_1319);
xnor U2080 (N_2080,In_1250,In_1534);
and U2081 (N_2081,In_740,In_113);
nand U2082 (N_2082,In_356,In_90);
nand U2083 (N_2083,In_433,In_1121);
and U2084 (N_2084,In_658,In_70);
nor U2085 (N_2085,In_1470,In_487);
and U2086 (N_2086,In_1371,In_399);
xor U2087 (N_2087,In_207,In_467);
nand U2088 (N_2088,In_1686,In_1365);
or U2089 (N_2089,In_1761,In_1430);
nor U2090 (N_2090,In_1513,In_1635);
nand U2091 (N_2091,In_107,In_1435);
nor U2092 (N_2092,In_59,In_92);
and U2093 (N_2093,In_1422,In_85);
nor U2094 (N_2094,In_1562,In_1476);
nand U2095 (N_2095,In_738,In_161);
and U2096 (N_2096,In_779,In_1947);
nor U2097 (N_2097,In_606,In_697);
or U2098 (N_2098,In_12,In_1041);
or U2099 (N_2099,In_193,In_1836);
and U2100 (N_2100,In_67,In_111);
nand U2101 (N_2101,In_794,In_1272);
xnor U2102 (N_2102,In_291,In_1909);
nor U2103 (N_2103,In_1284,In_1358);
nand U2104 (N_2104,In_888,In_1986);
nand U2105 (N_2105,In_1526,In_593);
or U2106 (N_2106,In_485,In_530);
nand U2107 (N_2107,In_952,In_1471);
or U2108 (N_2108,In_985,In_471);
nand U2109 (N_2109,In_1948,In_186);
nor U2110 (N_2110,In_438,In_1727);
nor U2111 (N_2111,In_1989,In_1336);
and U2112 (N_2112,In_1120,In_1493);
nor U2113 (N_2113,In_608,In_1589);
and U2114 (N_2114,In_1196,In_926);
nand U2115 (N_2115,In_988,In_424);
nand U2116 (N_2116,In_1448,In_188);
and U2117 (N_2117,In_124,In_166);
xnor U2118 (N_2118,In_535,In_1710);
and U2119 (N_2119,In_1506,In_1392);
nand U2120 (N_2120,In_1588,In_1393);
or U2121 (N_2121,In_264,In_994);
nand U2122 (N_2122,In_457,In_1065);
nand U2123 (N_2123,In_1414,In_1223);
nor U2124 (N_2124,In_937,In_1910);
nand U2125 (N_2125,In_1826,In_433);
and U2126 (N_2126,In_251,In_695);
xor U2127 (N_2127,In_1204,In_779);
xor U2128 (N_2128,In_1554,In_1967);
nand U2129 (N_2129,In_103,In_1208);
and U2130 (N_2130,In_845,In_715);
nor U2131 (N_2131,In_545,In_791);
and U2132 (N_2132,In_1054,In_554);
or U2133 (N_2133,In_1548,In_1813);
nor U2134 (N_2134,In_1179,In_766);
nand U2135 (N_2135,In_1235,In_1050);
and U2136 (N_2136,In_407,In_1206);
nor U2137 (N_2137,In_1491,In_1456);
nand U2138 (N_2138,In_1564,In_1368);
nand U2139 (N_2139,In_1972,In_683);
and U2140 (N_2140,In_358,In_970);
and U2141 (N_2141,In_897,In_512);
nand U2142 (N_2142,In_1193,In_500);
nor U2143 (N_2143,In_1359,In_1358);
xor U2144 (N_2144,In_1015,In_1304);
nor U2145 (N_2145,In_844,In_1333);
nor U2146 (N_2146,In_1093,In_1700);
and U2147 (N_2147,In_836,In_692);
xor U2148 (N_2148,In_45,In_1449);
or U2149 (N_2149,In_196,In_1152);
or U2150 (N_2150,In_91,In_1628);
nand U2151 (N_2151,In_1434,In_1370);
nand U2152 (N_2152,In_728,In_1187);
and U2153 (N_2153,In_1815,In_1480);
nand U2154 (N_2154,In_986,In_151);
nor U2155 (N_2155,In_1519,In_147);
or U2156 (N_2156,In_680,In_129);
or U2157 (N_2157,In_806,In_1864);
nand U2158 (N_2158,In_1450,In_1602);
and U2159 (N_2159,In_833,In_1738);
or U2160 (N_2160,In_341,In_27);
nand U2161 (N_2161,In_806,In_1487);
and U2162 (N_2162,In_1883,In_253);
or U2163 (N_2163,In_116,In_545);
or U2164 (N_2164,In_309,In_366);
nor U2165 (N_2165,In_1927,In_864);
xnor U2166 (N_2166,In_121,In_1156);
nor U2167 (N_2167,In_31,In_198);
or U2168 (N_2168,In_1873,In_451);
nor U2169 (N_2169,In_1740,In_1128);
nand U2170 (N_2170,In_1903,In_1260);
nor U2171 (N_2171,In_863,In_1616);
or U2172 (N_2172,In_934,In_618);
nor U2173 (N_2173,In_1162,In_660);
nor U2174 (N_2174,In_1415,In_1286);
or U2175 (N_2175,In_262,In_1776);
or U2176 (N_2176,In_9,In_178);
nand U2177 (N_2177,In_1065,In_1247);
and U2178 (N_2178,In_1130,In_360);
xor U2179 (N_2179,In_284,In_1511);
nor U2180 (N_2180,In_1386,In_1452);
nand U2181 (N_2181,In_1954,In_331);
and U2182 (N_2182,In_1941,In_1319);
and U2183 (N_2183,In_629,In_123);
nor U2184 (N_2184,In_1790,In_817);
nand U2185 (N_2185,In_911,In_1317);
nand U2186 (N_2186,In_1443,In_1878);
nand U2187 (N_2187,In_689,In_1604);
and U2188 (N_2188,In_1809,In_803);
xor U2189 (N_2189,In_999,In_88);
nand U2190 (N_2190,In_1693,In_1847);
and U2191 (N_2191,In_1600,In_1734);
nor U2192 (N_2192,In_1522,In_210);
or U2193 (N_2193,In_1471,In_282);
nand U2194 (N_2194,In_1263,In_242);
or U2195 (N_2195,In_267,In_1003);
and U2196 (N_2196,In_1170,In_1733);
nand U2197 (N_2197,In_1303,In_1249);
nand U2198 (N_2198,In_630,In_1211);
or U2199 (N_2199,In_1052,In_162);
or U2200 (N_2200,In_548,In_367);
nor U2201 (N_2201,In_845,In_541);
nand U2202 (N_2202,In_1245,In_148);
xnor U2203 (N_2203,In_1363,In_1083);
nor U2204 (N_2204,In_83,In_734);
and U2205 (N_2205,In_401,In_421);
xnor U2206 (N_2206,In_1965,In_1260);
nor U2207 (N_2207,In_1842,In_1783);
nor U2208 (N_2208,In_1130,In_954);
nand U2209 (N_2209,In_1001,In_183);
nand U2210 (N_2210,In_1301,In_1128);
xor U2211 (N_2211,In_874,In_1109);
or U2212 (N_2212,In_1340,In_864);
or U2213 (N_2213,In_412,In_697);
and U2214 (N_2214,In_172,In_1332);
nor U2215 (N_2215,In_1848,In_916);
or U2216 (N_2216,In_595,In_1933);
xor U2217 (N_2217,In_927,In_256);
nor U2218 (N_2218,In_1872,In_1853);
or U2219 (N_2219,In_845,In_865);
or U2220 (N_2220,In_1303,In_747);
nor U2221 (N_2221,In_1869,In_606);
nor U2222 (N_2222,In_1402,In_1547);
nor U2223 (N_2223,In_1966,In_1329);
nor U2224 (N_2224,In_1248,In_1588);
nor U2225 (N_2225,In_1002,In_1519);
and U2226 (N_2226,In_971,In_772);
nor U2227 (N_2227,In_853,In_1768);
nor U2228 (N_2228,In_341,In_1006);
nand U2229 (N_2229,In_1646,In_876);
nand U2230 (N_2230,In_238,In_604);
nand U2231 (N_2231,In_728,In_941);
and U2232 (N_2232,In_633,In_1417);
nor U2233 (N_2233,In_414,In_1711);
nor U2234 (N_2234,In_1209,In_204);
xor U2235 (N_2235,In_105,In_209);
nor U2236 (N_2236,In_1221,In_1094);
nor U2237 (N_2237,In_1653,In_210);
nand U2238 (N_2238,In_1254,In_202);
and U2239 (N_2239,In_933,In_1540);
nor U2240 (N_2240,In_1402,In_1976);
or U2241 (N_2241,In_587,In_1758);
nor U2242 (N_2242,In_590,In_1879);
and U2243 (N_2243,In_583,In_1833);
and U2244 (N_2244,In_976,In_3);
nand U2245 (N_2245,In_1566,In_1603);
or U2246 (N_2246,In_844,In_1267);
nor U2247 (N_2247,In_899,In_1025);
and U2248 (N_2248,In_754,In_211);
or U2249 (N_2249,In_133,In_1988);
xnor U2250 (N_2250,In_89,In_249);
nand U2251 (N_2251,In_1908,In_688);
and U2252 (N_2252,In_1837,In_1533);
nand U2253 (N_2253,In_1918,In_1980);
nand U2254 (N_2254,In_79,In_36);
and U2255 (N_2255,In_1481,In_1014);
or U2256 (N_2256,In_1696,In_1943);
nand U2257 (N_2257,In_267,In_852);
and U2258 (N_2258,In_1273,In_177);
and U2259 (N_2259,In_490,In_390);
nor U2260 (N_2260,In_760,In_1281);
and U2261 (N_2261,In_1604,In_1302);
or U2262 (N_2262,In_193,In_446);
nand U2263 (N_2263,In_1120,In_397);
xnor U2264 (N_2264,In_1968,In_1248);
nor U2265 (N_2265,In_330,In_541);
nor U2266 (N_2266,In_1557,In_1409);
and U2267 (N_2267,In_807,In_1144);
and U2268 (N_2268,In_193,In_1850);
and U2269 (N_2269,In_64,In_1577);
and U2270 (N_2270,In_1113,In_181);
xnor U2271 (N_2271,In_865,In_1646);
and U2272 (N_2272,In_1708,In_554);
and U2273 (N_2273,In_906,In_1573);
and U2274 (N_2274,In_450,In_1868);
nor U2275 (N_2275,In_570,In_255);
and U2276 (N_2276,In_453,In_1915);
nor U2277 (N_2277,In_1739,In_677);
nor U2278 (N_2278,In_118,In_1360);
nand U2279 (N_2279,In_624,In_1743);
and U2280 (N_2280,In_303,In_197);
or U2281 (N_2281,In_375,In_15);
nand U2282 (N_2282,In_1317,In_1395);
nor U2283 (N_2283,In_943,In_225);
nand U2284 (N_2284,In_770,In_677);
or U2285 (N_2285,In_1676,In_1289);
and U2286 (N_2286,In_143,In_500);
or U2287 (N_2287,In_1094,In_819);
or U2288 (N_2288,In_993,In_1352);
or U2289 (N_2289,In_1561,In_1005);
nand U2290 (N_2290,In_997,In_471);
nor U2291 (N_2291,In_232,In_1921);
and U2292 (N_2292,In_1,In_1673);
or U2293 (N_2293,In_1326,In_1837);
nand U2294 (N_2294,In_1769,In_970);
and U2295 (N_2295,In_1246,In_1531);
nor U2296 (N_2296,In_1921,In_91);
or U2297 (N_2297,In_1514,In_60);
nor U2298 (N_2298,In_639,In_318);
and U2299 (N_2299,In_113,In_1856);
and U2300 (N_2300,In_184,In_288);
or U2301 (N_2301,In_89,In_542);
and U2302 (N_2302,In_372,In_363);
nand U2303 (N_2303,In_1375,In_1010);
or U2304 (N_2304,In_215,In_1951);
nor U2305 (N_2305,In_288,In_413);
and U2306 (N_2306,In_1784,In_1732);
nor U2307 (N_2307,In_1611,In_110);
nand U2308 (N_2308,In_282,In_625);
xor U2309 (N_2309,In_1509,In_659);
xnor U2310 (N_2310,In_633,In_766);
nor U2311 (N_2311,In_1793,In_799);
or U2312 (N_2312,In_1405,In_175);
nor U2313 (N_2313,In_1797,In_604);
nand U2314 (N_2314,In_1565,In_501);
nor U2315 (N_2315,In_515,In_549);
nor U2316 (N_2316,In_1357,In_1400);
nand U2317 (N_2317,In_323,In_1129);
or U2318 (N_2318,In_875,In_594);
xnor U2319 (N_2319,In_1790,In_675);
xnor U2320 (N_2320,In_1811,In_1580);
or U2321 (N_2321,In_1219,In_352);
or U2322 (N_2322,In_1665,In_78);
xor U2323 (N_2323,In_922,In_49);
nor U2324 (N_2324,In_477,In_755);
or U2325 (N_2325,In_1800,In_1114);
nand U2326 (N_2326,In_784,In_715);
nor U2327 (N_2327,In_1717,In_576);
and U2328 (N_2328,In_664,In_130);
nand U2329 (N_2329,In_1426,In_1202);
and U2330 (N_2330,In_1644,In_517);
nor U2331 (N_2331,In_1310,In_1961);
nor U2332 (N_2332,In_1080,In_1107);
nand U2333 (N_2333,In_768,In_1942);
or U2334 (N_2334,In_965,In_1207);
nand U2335 (N_2335,In_1297,In_1065);
nand U2336 (N_2336,In_1595,In_1973);
or U2337 (N_2337,In_1277,In_1278);
nor U2338 (N_2338,In_258,In_1377);
or U2339 (N_2339,In_157,In_95);
xor U2340 (N_2340,In_673,In_1753);
and U2341 (N_2341,In_215,In_122);
or U2342 (N_2342,In_625,In_1846);
and U2343 (N_2343,In_849,In_1026);
nand U2344 (N_2344,In_683,In_757);
nand U2345 (N_2345,In_648,In_735);
nand U2346 (N_2346,In_1772,In_477);
nand U2347 (N_2347,In_343,In_1620);
and U2348 (N_2348,In_882,In_1196);
nor U2349 (N_2349,In_586,In_1141);
and U2350 (N_2350,In_1801,In_1116);
nand U2351 (N_2351,In_648,In_1804);
nand U2352 (N_2352,In_1826,In_54);
or U2353 (N_2353,In_1868,In_787);
nor U2354 (N_2354,In_1531,In_1965);
nand U2355 (N_2355,In_736,In_38);
nand U2356 (N_2356,In_380,In_1972);
nor U2357 (N_2357,In_1087,In_1411);
or U2358 (N_2358,In_323,In_108);
nand U2359 (N_2359,In_758,In_874);
and U2360 (N_2360,In_1529,In_591);
or U2361 (N_2361,In_1995,In_1709);
nor U2362 (N_2362,In_1920,In_1103);
and U2363 (N_2363,In_618,In_1161);
and U2364 (N_2364,In_1581,In_1765);
or U2365 (N_2365,In_1240,In_1598);
xor U2366 (N_2366,In_476,In_886);
or U2367 (N_2367,In_420,In_1233);
and U2368 (N_2368,In_407,In_1556);
nand U2369 (N_2369,In_1665,In_1945);
nor U2370 (N_2370,In_87,In_163);
nor U2371 (N_2371,In_673,In_1738);
xnor U2372 (N_2372,In_1256,In_576);
nand U2373 (N_2373,In_2,In_1066);
nand U2374 (N_2374,In_329,In_1726);
xnor U2375 (N_2375,In_274,In_588);
or U2376 (N_2376,In_1890,In_1120);
or U2377 (N_2377,In_1446,In_1195);
nand U2378 (N_2378,In_264,In_569);
and U2379 (N_2379,In_1956,In_1312);
nand U2380 (N_2380,In_1517,In_631);
or U2381 (N_2381,In_1310,In_1909);
or U2382 (N_2382,In_478,In_1817);
xor U2383 (N_2383,In_891,In_189);
or U2384 (N_2384,In_472,In_687);
nor U2385 (N_2385,In_38,In_1232);
and U2386 (N_2386,In_417,In_1587);
xor U2387 (N_2387,In_338,In_830);
or U2388 (N_2388,In_1349,In_1295);
nor U2389 (N_2389,In_1508,In_847);
or U2390 (N_2390,In_1221,In_1599);
and U2391 (N_2391,In_789,In_539);
nor U2392 (N_2392,In_667,In_21);
and U2393 (N_2393,In_1916,In_325);
or U2394 (N_2394,In_986,In_1248);
nor U2395 (N_2395,In_1121,In_229);
and U2396 (N_2396,In_539,In_889);
and U2397 (N_2397,In_561,In_1788);
or U2398 (N_2398,In_1136,In_998);
nor U2399 (N_2399,In_1835,In_1402);
xnor U2400 (N_2400,In_1936,In_754);
or U2401 (N_2401,In_977,In_567);
and U2402 (N_2402,In_1461,In_1098);
nor U2403 (N_2403,In_310,In_641);
and U2404 (N_2404,In_1335,In_675);
nand U2405 (N_2405,In_781,In_847);
or U2406 (N_2406,In_153,In_813);
or U2407 (N_2407,In_1108,In_1788);
xnor U2408 (N_2408,In_766,In_1053);
and U2409 (N_2409,In_1647,In_1052);
xnor U2410 (N_2410,In_179,In_1841);
xor U2411 (N_2411,In_1222,In_1939);
and U2412 (N_2412,In_184,In_1769);
and U2413 (N_2413,In_256,In_1060);
and U2414 (N_2414,In_835,In_19);
nor U2415 (N_2415,In_694,In_1256);
nand U2416 (N_2416,In_1366,In_1676);
nor U2417 (N_2417,In_969,In_1124);
or U2418 (N_2418,In_1878,In_1881);
nand U2419 (N_2419,In_230,In_1341);
or U2420 (N_2420,In_634,In_477);
and U2421 (N_2421,In_187,In_192);
and U2422 (N_2422,In_1724,In_330);
or U2423 (N_2423,In_1694,In_1253);
nand U2424 (N_2424,In_1,In_1748);
nand U2425 (N_2425,In_1152,In_510);
nand U2426 (N_2426,In_537,In_1791);
and U2427 (N_2427,In_1701,In_1674);
nand U2428 (N_2428,In_982,In_1862);
nor U2429 (N_2429,In_776,In_163);
nor U2430 (N_2430,In_1812,In_673);
nand U2431 (N_2431,In_1534,In_701);
or U2432 (N_2432,In_1537,In_1425);
and U2433 (N_2433,In_1740,In_543);
or U2434 (N_2434,In_934,In_1324);
nand U2435 (N_2435,In_1568,In_274);
xnor U2436 (N_2436,In_853,In_1620);
nand U2437 (N_2437,In_1355,In_1221);
nand U2438 (N_2438,In_310,In_1174);
and U2439 (N_2439,In_1273,In_98);
xor U2440 (N_2440,In_1878,In_300);
and U2441 (N_2441,In_1717,In_1007);
and U2442 (N_2442,In_1996,In_1669);
and U2443 (N_2443,In_588,In_965);
or U2444 (N_2444,In_540,In_765);
nand U2445 (N_2445,In_1389,In_253);
nor U2446 (N_2446,In_1400,In_1941);
and U2447 (N_2447,In_1801,In_1125);
xnor U2448 (N_2448,In_1005,In_917);
or U2449 (N_2449,In_795,In_325);
or U2450 (N_2450,In_1176,In_1952);
and U2451 (N_2451,In_1878,In_1228);
nand U2452 (N_2452,In_1476,In_1702);
nor U2453 (N_2453,In_1360,In_228);
nand U2454 (N_2454,In_488,In_914);
and U2455 (N_2455,In_213,In_1161);
and U2456 (N_2456,In_879,In_160);
nor U2457 (N_2457,In_1456,In_1175);
xor U2458 (N_2458,In_284,In_714);
or U2459 (N_2459,In_1275,In_1517);
and U2460 (N_2460,In_973,In_1162);
xnor U2461 (N_2461,In_941,In_1209);
and U2462 (N_2462,In_560,In_243);
xnor U2463 (N_2463,In_128,In_512);
nor U2464 (N_2464,In_1670,In_1329);
nor U2465 (N_2465,In_1836,In_405);
and U2466 (N_2466,In_878,In_406);
and U2467 (N_2467,In_1782,In_580);
and U2468 (N_2468,In_1181,In_1559);
and U2469 (N_2469,In_1019,In_625);
or U2470 (N_2470,In_118,In_1780);
xor U2471 (N_2471,In_46,In_1844);
nand U2472 (N_2472,In_698,In_1456);
or U2473 (N_2473,In_1389,In_216);
xnor U2474 (N_2474,In_819,In_543);
nand U2475 (N_2475,In_1736,In_421);
nand U2476 (N_2476,In_1125,In_1193);
nor U2477 (N_2477,In_931,In_918);
nand U2478 (N_2478,In_1538,In_1168);
xor U2479 (N_2479,In_633,In_1127);
nor U2480 (N_2480,In_1094,In_975);
nand U2481 (N_2481,In_244,In_1793);
xor U2482 (N_2482,In_970,In_417);
or U2483 (N_2483,In_1621,In_1881);
nand U2484 (N_2484,In_1587,In_190);
nor U2485 (N_2485,In_1289,In_1060);
and U2486 (N_2486,In_1456,In_1215);
and U2487 (N_2487,In_247,In_1490);
and U2488 (N_2488,In_883,In_401);
nor U2489 (N_2489,In_1123,In_20);
nand U2490 (N_2490,In_1130,In_1023);
and U2491 (N_2491,In_1033,In_1007);
or U2492 (N_2492,In_550,In_1541);
xnor U2493 (N_2493,In_1614,In_1879);
or U2494 (N_2494,In_162,In_1979);
and U2495 (N_2495,In_1070,In_485);
nor U2496 (N_2496,In_853,In_398);
nand U2497 (N_2497,In_666,In_514);
and U2498 (N_2498,In_233,In_1443);
or U2499 (N_2499,In_371,In_1683);
and U2500 (N_2500,In_1572,In_109);
and U2501 (N_2501,In_1690,In_60);
nand U2502 (N_2502,In_1038,In_559);
nor U2503 (N_2503,In_1316,In_343);
xnor U2504 (N_2504,In_331,In_9);
xnor U2505 (N_2505,In_662,In_243);
nand U2506 (N_2506,In_1186,In_1963);
xor U2507 (N_2507,In_1391,In_542);
nand U2508 (N_2508,In_438,In_1401);
nor U2509 (N_2509,In_812,In_1826);
nand U2510 (N_2510,In_532,In_1769);
and U2511 (N_2511,In_799,In_1129);
nand U2512 (N_2512,In_1871,In_846);
nor U2513 (N_2513,In_1283,In_1654);
and U2514 (N_2514,In_1902,In_450);
nor U2515 (N_2515,In_1712,In_253);
nand U2516 (N_2516,In_1143,In_950);
or U2517 (N_2517,In_360,In_727);
xnor U2518 (N_2518,In_386,In_1052);
nor U2519 (N_2519,In_1984,In_1105);
nand U2520 (N_2520,In_1916,In_1380);
xor U2521 (N_2521,In_65,In_898);
or U2522 (N_2522,In_1653,In_1203);
nor U2523 (N_2523,In_842,In_744);
or U2524 (N_2524,In_1141,In_20);
and U2525 (N_2525,In_1581,In_420);
or U2526 (N_2526,In_493,In_357);
or U2527 (N_2527,In_1555,In_657);
or U2528 (N_2528,In_897,In_1105);
or U2529 (N_2529,In_848,In_1950);
xnor U2530 (N_2530,In_949,In_466);
nor U2531 (N_2531,In_1456,In_1165);
nand U2532 (N_2532,In_980,In_188);
nor U2533 (N_2533,In_1956,In_674);
or U2534 (N_2534,In_1433,In_1810);
xor U2535 (N_2535,In_1228,In_367);
nand U2536 (N_2536,In_1047,In_266);
or U2537 (N_2537,In_492,In_1721);
or U2538 (N_2538,In_617,In_118);
and U2539 (N_2539,In_1154,In_588);
nand U2540 (N_2540,In_1109,In_1410);
or U2541 (N_2541,In_197,In_1809);
or U2542 (N_2542,In_46,In_285);
nor U2543 (N_2543,In_1529,In_1888);
and U2544 (N_2544,In_573,In_1480);
and U2545 (N_2545,In_1233,In_1629);
or U2546 (N_2546,In_1433,In_912);
nor U2547 (N_2547,In_1238,In_1373);
nor U2548 (N_2548,In_1442,In_1174);
and U2549 (N_2549,In_736,In_625);
nand U2550 (N_2550,In_1224,In_1526);
xnor U2551 (N_2551,In_702,In_328);
and U2552 (N_2552,In_1540,In_342);
and U2553 (N_2553,In_482,In_1936);
xor U2554 (N_2554,In_1721,In_1960);
xor U2555 (N_2555,In_1454,In_609);
and U2556 (N_2556,In_1026,In_218);
and U2557 (N_2557,In_1096,In_1357);
xnor U2558 (N_2558,In_1118,In_1515);
and U2559 (N_2559,In_964,In_1666);
nand U2560 (N_2560,In_1029,In_46);
nand U2561 (N_2561,In_689,In_711);
nor U2562 (N_2562,In_579,In_1688);
or U2563 (N_2563,In_315,In_463);
xnor U2564 (N_2564,In_1240,In_1513);
nand U2565 (N_2565,In_1617,In_1591);
nor U2566 (N_2566,In_811,In_601);
and U2567 (N_2567,In_317,In_970);
and U2568 (N_2568,In_459,In_1030);
or U2569 (N_2569,In_123,In_790);
or U2570 (N_2570,In_320,In_1670);
or U2571 (N_2571,In_1850,In_930);
and U2572 (N_2572,In_1056,In_19);
or U2573 (N_2573,In_306,In_361);
nand U2574 (N_2574,In_654,In_1978);
nand U2575 (N_2575,In_1475,In_1379);
nor U2576 (N_2576,In_1053,In_1668);
nor U2577 (N_2577,In_1541,In_267);
and U2578 (N_2578,In_662,In_972);
nand U2579 (N_2579,In_752,In_1443);
nor U2580 (N_2580,In_505,In_457);
or U2581 (N_2581,In_608,In_1216);
and U2582 (N_2582,In_639,In_1552);
or U2583 (N_2583,In_1876,In_1168);
or U2584 (N_2584,In_784,In_1194);
and U2585 (N_2585,In_214,In_553);
and U2586 (N_2586,In_1442,In_623);
nor U2587 (N_2587,In_1050,In_477);
nor U2588 (N_2588,In_1491,In_1404);
and U2589 (N_2589,In_988,In_523);
xnor U2590 (N_2590,In_77,In_134);
and U2591 (N_2591,In_1334,In_1162);
nand U2592 (N_2592,In_74,In_1741);
nand U2593 (N_2593,In_529,In_454);
or U2594 (N_2594,In_637,In_1699);
nand U2595 (N_2595,In_201,In_797);
and U2596 (N_2596,In_1214,In_1263);
nand U2597 (N_2597,In_580,In_66);
nor U2598 (N_2598,In_503,In_202);
nor U2599 (N_2599,In_293,In_133);
and U2600 (N_2600,In_1460,In_996);
or U2601 (N_2601,In_1138,In_679);
nor U2602 (N_2602,In_892,In_1085);
and U2603 (N_2603,In_681,In_1829);
and U2604 (N_2604,In_1706,In_800);
or U2605 (N_2605,In_1393,In_1310);
and U2606 (N_2606,In_1019,In_590);
and U2607 (N_2607,In_1254,In_1758);
nand U2608 (N_2608,In_420,In_1899);
nand U2609 (N_2609,In_1322,In_244);
or U2610 (N_2610,In_571,In_1667);
nand U2611 (N_2611,In_1056,In_983);
and U2612 (N_2612,In_1942,In_90);
nand U2613 (N_2613,In_774,In_1416);
or U2614 (N_2614,In_699,In_829);
nand U2615 (N_2615,In_1667,In_279);
nor U2616 (N_2616,In_456,In_1130);
and U2617 (N_2617,In_774,In_545);
nor U2618 (N_2618,In_373,In_1699);
nor U2619 (N_2619,In_1989,In_1330);
or U2620 (N_2620,In_1761,In_866);
or U2621 (N_2621,In_44,In_687);
nand U2622 (N_2622,In_43,In_457);
and U2623 (N_2623,In_1703,In_1375);
and U2624 (N_2624,In_1397,In_1666);
nand U2625 (N_2625,In_1701,In_1200);
or U2626 (N_2626,In_640,In_491);
and U2627 (N_2627,In_1909,In_1408);
or U2628 (N_2628,In_294,In_77);
and U2629 (N_2629,In_339,In_1880);
nand U2630 (N_2630,In_494,In_1688);
nor U2631 (N_2631,In_530,In_259);
and U2632 (N_2632,In_1665,In_989);
xor U2633 (N_2633,In_285,In_24);
and U2634 (N_2634,In_1678,In_1891);
nand U2635 (N_2635,In_251,In_1999);
and U2636 (N_2636,In_339,In_443);
nand U2637 (N_2637,In_812,In_588);
nor U2638 (N_2638,In_1791,In_1658);
and U2639 (N_2639,In_1516,In_222);
nand U2640 (N_2640,In_1608,In_1004);
and U2641 (N_2641,In_1971,In_165);
xor U2642 (N_2642,In_1151,In_795);
nand U2643 (N_2643,In_1782,In_1814);
and U2644 (N_2644,In_1013,In_1399);
nand U2645 (N_2645,In_651,In_204);
and U2646 (N_2646,In_495,In_1288);
nor U2647 (N_2647,In_1220,In_1009);
and U2648 (N_2648,In_1541,In_1817);
and U2649 (N_2649,In_1196,In_288);
nand U2650 (N_2650,In_585,In_109);
nand U2651 (N_2651,In_1745,In_864);
nand U2652 (N_2652,In_1571,In_549);
xnor U2653 (N_2653,In_1623,In_960);
and U2654 (N_2654,In_1986,In_669);
or U2655 (N_2655,In_1209,In_216);
and U2656 (N_2656,In_1325,In_1645);
and U2657 (N_2657,In_297,In_303);
and U2658 (N_2658,In_1360,In_406);
nor U2659 (N_2659,In_961,In_1373);
or U2660 (N_2660,In_1883,In_998);
xor U2661 (N_2661,In_656,In_405);
xnor U2662 (N_2662,In_1120,In_1207);
and U2663 (N_2663,In_1562,In_1361);
nor U2664 (N_2664,In_1742,In_1914);
nor U2665 (N_2665,In_1152,In_280);
and U2666 (N_2666,In_1192,In_559);
nand U2667 (N_2667,In_1521,In_410);
xnor U2668 (N_2668,In_29,In_616);
or U2669 (N_2669,In_1841,In_940);
and U2670 (N_2670,In_686,In_602);
nand U2671 (N_2671,In_1544,In_1905);
and U2672 (N_2672,In_1929,In_1441);
nand U2673 (N_2673,In_1370,In_561);
or U2674 (N_2674,In_1152,In_990);
xor U2675 (N_2675,In_1994,In_964);
nand U2676 (N_2676,In_397,In_596);
nor U2677 (N_2677,In_345,In_1376);
xnor U2678 (N_2678,In_204,In_1561);
or U2679 (N_2679,In_1060,In_1810);
nand U2680 (N_2680,In_807,In_1311);
xor U2681 (N_2681,In_1659,In_1472);
nand U2682 (N_2682,In_1409,In_1317);
and U2683 (N_2683,In_141,In_973);
or U2684 (N_2684,In_271,In_801);
and U2685 (N_2685,In_400,In_1810);
nor U2686 (N_2686,In_959,In_1593);
nor U2687 (N_2687,In_369,In_1697);
and U2688 (N_2688,In_551,In_432);
nor U2689 (N_2689,In_1490,In_481);
nand U2690 (N_2690,In_947,In_124);
or U2691 (N_2691,In_635,In_528);
xor U2692 (N_2692,In_846,In_209);
nand U2693 (N_2693,In_1629,In_1545);
and U2694 (N_2694,In_1893,In_1248);
nand U2695 (N_2695,In_221,In_968);
nand U2696 (N_2696,In_1562,In_426);
nand U2697 (N_2697,In_548,In_178);
nor U2698 (N_2698,In_1240,In_1419);
nor U2699 (N_2699,In_444,In_273);
nand U2700 (N_2700,In_1409,In_604);
or U2701 (N_2701,In_610,In_1849);
xor U2702 (N_2702,In_1068,In_1968);
or U2703 (N_2703,In_643,In_979);
nand U2704 (N_2704,In_985,In_1470);
nor U2705 (N_2705,In_1570,In_110);
nand U2706 (N_2706,In_561,In_1912);
xor U2707 (N_2707,In_1533,In_925);
nand U2708 (N_2708,In_1975,In_53);
or U2709 (N_2709,In_871,In_1327);
nand U2710 (N_2710,In_563,In_1953);
and U2711 (N_2711,In_264,In_481);
xnor U2712 (N_2712,In_1560,In_571);
nand U2713 (N_2713,In_281,In_828);
or U2714 (N_2714,In_1303,In_1193);
xnor U2715 (N_2715,In_519,In_113);
or U2716 (N_2716,In_762,In_1825);
or U2717 (N_2717,In_1994,In_826);
nand U2718 (N_2718,In_1407,In_981);
xor U2719 (N_2719,In_1857,In_1348);
or U2720 (N_2720,In_570,In_398);
xor U2721 (N_2721,In_1863,In_1131);
nor U2722 (N_2722,In_868,In_602);
nor U2723 (N_2723,In_669,In_959);
and U2724 (N_2724,In_186,In_902);
nor U2725 (N_2725,In_800,In_1227);
nor U2726 (N_2726,In_1491,In_6);
and U2727 (N_2727,In_1922,In_1925);
or U2728 (N_2728,In_1582,In_1528);
xor U2729 (N_2729,In_226,In_1709);
nor U2730 (N_2730,In_715,In_1053);
nand U2731 (N_2731,In_1093,In_1521);
or U2732 (N_2732,In_639,In_284);
nand U2733 (N_2733,In_679,In_1262);
nor U2734 (N_2734,In_338,In_192);
nand U2735 (N_2735,In_1066,In_1117);
or U2736 (N_2736,In_1095,In_1518);
or U2737 (N_2737,In_942,In_1997);
or U2738 (N_2738,In_657,In_791);
and U2739 (N_2739,In_93,In_1339);
nand U2740 (N_2740,In_695,In_1485);
nor U2741 (N_2741,In_1876,In_1090);
and U2742 (N_2742,In_1630,In_457);
or U2743 (N_2743,In_18,In_1822);
nand U2744 (N_2744,In_1123,In_1999);
or U2745 (N_2745,In_1741,In_460);
or U2746 (N_2746,In_1507,In_1027);
and U2747 (N_2747,In_713,In_1282);
nand U2748 (N_2748,In_625,In_1491);
or U2749 (N_2749,In_947,In_1662);
and U2750 (N_2750,In_1447,In_1075);
nand U2751 (N_2751,In_1218,In_68);
or U2752 (N_2752,In_760,In_881);
or U2753 (N_2753,In_733,In_979);
or U2754 (N_2754,In_1746,In_678);
and U2755 (N_2755,In_820,In_1810);
nor U2756 (N_2756,In_1420,In_1942);
xnor U2757 (N_2757,In_253,In_513);
nor U2758 (N_2758,In_1275,In_1526);
nor U2759 (N_2759,In_171,In_1227);
nor U2760 (N_2760,In_1196,In_1068);
and U2761 (N_2761,In_1868,In_1991);
and U2762 (N_2762,In_1515,In_1340);
nand U2763 (N_2763,In_583,In_1571);
or U2764 (N_2764,In_1616,In_1519);
nor U2765 (N_2765,In_1773,In_1089);
nor U2766 (N_2766,In_878,In_512);
and U2767 (N_2767,In_1212,In_180);
nor U2768 (N_2768,In_1804,In_1957);
nor U2769 (N_2769,In_1163,In_1663);
xor U2770 (N_2770,In_599,In_695);
nand U2771 (N_2771,In_804,In_1506);
nor U2772 (N_2772,In_1030,In_1660);
and U2773 (N_2773,In_202,In_1977);
and U2774 (N_2774,In_167,In_513);
xnor U2775 (N_2775,In_1469,In_251);
nor U2776 (N_2776,In_1892,In_528);
nor U2777 (N_2777,In_1345,In_992);
and U2778 (N_2778,In_464,In_1706);
nand U2779 (N_2779,In_353,In_1027);
and U2780 (N_2780,In_1156,In_1772);
nor U2781 (N_2781,In_1586,In_1576);
or U2782 (N_2782,In_655,In_1639);
and U2783 (N_2783,In_115,In_1734);
or U2784 (N_2784,In_1815,In_1921);
or U2785 (N_2785,In_687,In_998);
nor U2786 (N_2786,In_187,In_1387);
and U2787 (N_2787,In_936,In_255);
xor U2788 (N_2788,In_1238,In_998);
nor U2789 (N_2789,In_466,In_871);
or U2790 (N_2790,In_1703,In_1380);
nand U2791 (N_2791,In_1919,In_1737);
nor U2792 (N_2792,In_1676,In_172);
nor U2793 (N_2793,In_1478,In_1703);
xnor U2794 (N_2794,In_1663,In_1781);
nand U2795 (N_2795,In_1024,In_1145);
nor U2796 (N_2796,In_1170,In_1787);
nor U2797 (N_2797,In_1429,In_1067);
or U2798 (N_2798,In_768,In_790);
nand U2799 (N_2799,In_331,In_1794);
xor U2800 (N_2800,In_1701,In_637);
and U2801 (N_2801,In_58,In_553);
nand U2802 (N_2802,In_584,In_794);
nor U2803 (N_2803,In_114,In_1780);
nand U2804 (N_2804,In_902,In_785);
and U2805 (N_2805,In_900,In_1892);
and U2806 (N_2806,In_166,In_664);
or U2807 (N_2807,In_671,In_408);
nor U2808 (N_2808,In_334,In_1085);
or U2809 (N_2809,In_531,In_466);
nand U2810 (N_2810,In_692,In_818);
xor U2811 (N_2811,In_52,In_679);
or U2812 (N_2812,In_478,In_1348);
and U2813 (N_2813,In_1481,In_1339);
or U2814 (N_2814,In_1320,In_1999);
nand U2815 (N_2815,In_326,In_472);
nor U2816 (N_2816,In_1816,In_481);
or U2817 (N_2817,In_778,In_1310);
nand U2818 (N_2818,In_1399,In_250);
and U2819 (N_2819,In_707,In_1704);
and U2820 (N_2820,In_938,In_1443);
or U2821 (N_2821,In_1321,In_394);
nand U2822 (N_2822,In_1632,In_1775);
nor U2823 (N_2823,In_597,In_1180);
or U2824 (N_2824,In_1796,In_1402);
nor U2825 (N_2825,In_1495,In_1391);
or U2826 (N_2826,In_290,In_494);
and U2827 (N_2827,In_650,In_1758);
nand U2828 (N_2828,In_892,In_229);
or U2829 (N_2829,In_1622,In_1485);
nand U2830 (N_2830,In_1570,In_590);
and U2831 (N_2831,In_1858,In_945);
and U2832 (N_2832,In_161,In_1328);
nor U2833 (N_2833,In_950,In_869);
and U2834 (N_2834,In_1303,In_1214);
nor U2835 (N_2835,In_83,In_1088);
nor U2836 (N_2836,In_1708,In_842);
xnor U2837 (N_2837,In_427,In_717);
nand U2838 (N_2838,In_1684,In_961);
and U2839 (N_2839,In_1600,In_1264);
or U2840 (N_2840,In_1551,In_1022);
and U2841 (N_2841,In_1505,In_530);
and U2842 (N_2842,In_1016,In_1397);
or U2843 (N_2843,In_1525,In_847);
xnor U2844 (N_2844,In_134,In_1313);
nor U2845 (N_2845,In_1506,In_798);
or U2846 (N_2846,In_1744,In_426);
nand U2847 (N_2847,In_813,In_370);
nor U2848 (N_2848,In_1749,In_996);
or U2849 (N_2849,In_1247,In_342);
and U2850 (N_2850,In_777,In_1353);
nor U2851 (N_2851,In_318,In_1100);
nand U2852 (N_2852,In_1948,In_705);
or U2853 (N_2853,In_579,In_578);
nand U2854 (N_2854,In_740,In_634);
or U2855 (N_2855,In_1529,In_1297);
and U2856 (N_2856,In_484,In_154);
nor U2857 (N_2857,In_1285,In_574);
and U2858 (N_2858,In_267,In_1222);
or U2859 (N_2859,In_117,In_1967);
nand U2860 (N_2860,In_1751,In_1552);
and U2861 (N_2861,In_1479,In_1941);
nor U2862 (N_2862,In_1267,In_595);
nand U2863 (N_2863,In_786,In_237);
or U2864 (N_2864,In_522,In_1118);
nor U2865 (N_2865,In_1543,In_643);
and U2866 (N_2866,In_1049,In_1564);
nor U2867 (N_2867,In_1631,In_1345);
or U2868 (N_2868,In_1400,In_638);
nand U2869 (N_2869,In_1893,In_1496);
nand U2870 (N_2870,In_1507,In_62);
or U2871 (N_2871,In_1315,In_940);
xor U2872 (N_2872,In_229,In_1137);
nand U2873 (N_2873,In_1225,In_945);
or U2874 (N_2874,In_1301,In_1487);
nor U2875 (N_2875,In_1060,In_40);
nor U2876 (N_2876,In_1265,In_15);
nor U2877 (N_2877,In_545,In_1596);
nand U2878 (N_2878,In_183,In_835);
xor U2879 (N_2879,In_1279,In_1478);
nand U2880 (N_2880,In_76,In_211);
nand U2881 (N_2881,In_1770,In_1743);
nor U2882 (N_2882,In_779,In_1530);
nand U2883 (N_2883,In_404,In_826);
nand U2884 (N_2884,In_762,In_526);
nand U2885 (N_2885,In_1184,In_1873);
nand U2886 (N_2886,In_1212,In_269);
or U2887 (N_2887,In_138,In_484);
and U2888 (N_2888,In_1402,In_1872);
nand U2889 (N_2889,In_965,In_1930);
nor U2890 (N_2890,In_1798,In_125);
or U2891 (N_2891,In_1178,In_871);
or U2892 (N_2892,In_1692,In_1042);
xnor U2893 (N_2893,In_1274,In_90);
nor U2894 (N_2894,In_1603,In_1004);
or U2895 (N_2895,In_181,In_365);
nor U2896 (N_2896,In_674,In_1079);
nand U2897 (N_2897,In_1261,In_153);
nor U2898 (N_2898,In_778,In_835);
xor U2899 (N_2899,In_861,In_1714);
nand U2900 (N_2900,In_1582,In_238);
nand U2901 (N_2901,In_1969,In_1885);
nor U2902 (N_2902,In_686,In_720);
nor U2903 (N_2903,In_623,In_292);
nand U2904 (N_2904,In_1850,In_1368);
and U2905 (N_2905,In_1029,In_204);
or U2906 (N_2906,In_829,In_500);
and U2907 (N_2907,In_1344,In_731);
nand U2908 (N_2908,In_710,In_1612);
nand U2909 (N_2909,In_624,In_717);
nor U2910 (N_2910,In_915,In_1641);
nor U2911 (N_2911,In_442,In_680);
and U2912 (N_2912,In_1595,In_492);
or U2913 (N_2913,In_1173,In_1800);
nand U2914 (N_2914,In_613,In_1614);
nor U2915 (N_2915,In_1785,In_349);
nand U2916 (N_2916,In_1703,In_138);
or U2917 (N_2917,In_694,In_1848);
and U2918 (N_2918,In_1976,In_71);
nand U2919 (N_2919,In_314,In_493);
and U2920 (N_2920,In_812,In_1925);
or U2921 (N_2921,In_480,In_250);
nand U2922 (N_2922,In_266,In_1976);
xnor U2923 (N_2923,In_1485,In_1677);
or U2924 (N_2924,In_1295,In_991);
nor U2925 (N_2925,In_1221,In_879);
and U2926 (N_2926,In_917,In_1429);
nand U2927 (N_2927,In_1236,In_1174);
or U2928 (N_2928,In_105,In_1033);
nor U2929 (N_2929,In_920,In_1951);
or U2930 (N_2930,In_222,In_649);
and U2931 (N_2931,In_1498,In_1023);
nand U2932 (N_2932,In_772,In_1120);
nor U2933 (N_2933,In_746,In_1557);
and U2934 (N_2934,In_1956,In_1063);
nor U2935 (N_2935,In_953,In_1205);
nor U2936 (N_2936,In_1428,In_828);
nand U2937 (N_2937,In_11,In_1100);
and U2938 (N_2938,In_573,In_72);
nor U2939 (N_2939,In_1573,In_531);
or U2940 (N_2940,In_473,In_44);
nor U2941 (N_2941,In_82,In_1986);
and U2942 (N_2942,In_882,In_685);
xnor U2943 (N_2943,In_621,In_473);
nand U2944 (N_2944,In_1490,In_1638);
nand U2945 (N_2945,In_1213,In_1749);
and U2946 (N_2946,In_1966,In_848);
or U2947 (N_2947,In_515,In_100);
nand U2948 (N_2948,In_764,In_1215);
nor U2949 (N_2949,In_1633,In_533);
nand U2950 (N_2950,In_487,In_447);
and U2951 (N_2951,In_768,In_1884);
xor U2952 (N_2952,In_777,In_810);
nand U2953 (N_2953,In_1519,In_597);
and U2954 (N_2954,In_534,In_38);
nor U2955 (N_2955,In_111,In_992);
xor U2956 (N_2956,In_1535,In_91);
and U2957 (N_2957,In_1524,In_623);
nand U2958 (N_2958,In_1866,In_1962);
nand U2959 (N_2959,In_711,In_1564);
xor U2960 (N_2960,In_487,In_415);
or U2961 (N_2961,In_415,In_1011);
and U2962 (N_2962,In_906,In_729);
nand U2963 (N_2963,In_1309,In_1610);
nor U2964 (N_2964,In_1176,In_121);
nor U2965 (N_2965,In_1511,In_368);
or U2966 (N_2966,In_1711,In_568);
nand U2967 (N_2967,In_688,In_46);
nand U2968 (N_2968,In_808,In_918);
nor U2969 (N_2969,In_1723,In_551);
xor U2970 (N_2970,In_1780,In_1758);
nor U2971 (N_2971,In_1045,In_77);
nand U2972 (N_2972,In_1967,In_50);
nor U2973 (N_2973,In_404,In_653);
or U2974 (N_2974,In_94,In_583);
and U2975 (N_2975,In_201,In_398);
or U2976 (N_2976,In_115,In_1146);
xor U2977 (N_2977,In_1418,In_349);
or U2978 (N_2978,In_1088,In_1980);
nor U2979 (N_2979,In_1747,In_481);
nand U2980 (N_2980,In_1883,In_1965);
xor U2981 (N_2981,In_1709,In_1408);
nor U2982 (N_2982,In_723,In_96);
or U2983 (N_2983,In_865,In_892);
and U2984 (N_2984,In_1201,In_1622);
nor U2985 (N_2985,In_454,In_1737);
or U2986 (N_2986,In_173,In_432);
and U2987 (N_2987,In_1587,In_1198);
nor U2988 (N_2988,In_631,In_705);
nand U2989 (N_2989,In_1189,In_797);
or U2990 (N_2990,In_434,In_586);
nand U2991 (N_2991,In_1875,In_1364);
or U2992 (N_2992,In_1030,In_263);
nor U2993 (N_2993,In_363,In_1539);
or U2994 (N_2994,In_1787,In_340);
nand U2995 (N_2995,In_539,In_258);
nand U2996 (N_2996,In_1909,In_343);
nand U2997 (N_2997,In_883,In_928);
and U2998 (N_2998,In_1955,In_423);
nor U2999 (N_2999,In_597,In_1111);
or U3000 (N_3000,In_18,In_150);
or U3001 (N_3001,In_695,In_1514);
and U3002 (N_3002,In_1034,In_967);
nand U3003 (N_3003,In_1161,In_1236);
xnor U3004 (N_3004,In_896,In_68);
and U3005 (N_3005,In_105,In_1785);
and U3006 (N_3006,In_217,In_1003);
and U3007 (N_3007,In_1974,In_1322);
and U3008 (N_3008,In_185,In_1045);
xor U3009 (N_3009,In_357,In_943);
nor U3010 (N_3010,In_352,In_1899);
nand U3011 (N_3011,In_393,In_1714);
nand U3012 (N_3012,In_1620,In_1102);
xor U3013 (N_3013,In_891,In_1820);
or U3014 (N_3014,In_157,In_279);
xnor U3015 (N_3015,In_579,In_96);
nand U3016 (N_3016,In_1869,In_734);
or U3017 (N_3017,In_1417,In_637);
and U3018 (N_3018,In_1195,In_285);
or U3019 (N_3019,In_589,In_1634);
nand U3020 (N_3020,In_1750,In_1076);
nor U3021 (N_3021,In_534,In_1175);
xnor U3022 (N_3022,In_1997,In_1189);
nand U3023 (N_3023,In_1144,In_1293);
or U3024 (N_3024,In_1913,In_980);
nor U3025 (N_3025,In_1651,In_374);
nor U3026 (N_3026,In_766,In_1651);
nor U3027 (N_3027,In_198,In_1272);
nor U3028 (N_3028,In_1246,In_1867);
and U3029 (N_3029,In_1201,In_702);
xnor U3030 (N_3030,In_789,In_1556);
and U3031 (N_3031,In_1461,In_1334);
or U3032 (N_3032,In_1068,In_1430);
nor U3033 (N_3033,In_474,In_714);
xnor U3034 (N_3034,In_620,In_1406);
nand U3035 (N_3035,In_1090,In_1686);
or U3036 (N_3036,In_519,In_999);
and U3037 (N_3037,In_1007,In_1532);
nor U3038 (N_3038,In_885,In_1177);
nand U3039 (N_3039,In_1423,In_1721);
nor U3040 (N_3040,In_973,In_1795);
nand U3041 (N_3041,In_170,In_989);
nand U3042 (N_3042,In_1002,In_1028);
or U3043 (N_3043,In_892,In_1468);
nor U3044 (N_3044,In_370,In_9);
xor U3045 (N_3045,In_1458,In_720);
nor U3046 (N_3046,In_393,In_868);
nand U3047 (N_3047,In_1307,In_1113);
nand U3048 (N_3048,In_1131,In_396);
nor U3049 (N_3049,In_1323,In_1549);
nor U3050 (N_3050,In_1659,In_1696);
nor U3051 (N_3051,In_682,In_687);
nand U3052 (N_3052,In_1150,In_1853);
and U3053 (N_3053,In_99,In_439);
nand U3054 (N_3054,In_540,In_67);
and U3055 (N_3055,In_1037,In_1193);
or U3056 (N_3056,In_1037,In_1942);
and U3057 (N_3057,In_813,In_1020);
or U3058 (N_3058,In_1372,In_590);
nor U3059 (N_3059,In_500,In_501);
nor U3060 (N_3060,In_525,In_1787);
xnor U3061 (N_3061,In_255,In_1426);
nor U3062 (N_3062,In_1,In_795);
or U3063 (N_3063,In_1010,In_528);
or U3064 (N_3064,In_1261,In_1493);
and U3065 (N_3065,In_26,In_1156);
and U3066 (N_3066,In_1238,In_1160);
nand U3067 (N_3067,In_207,In_281);
nor U3068 (N_3068,In_408,In_1551);
or U3069 (N_3069,In_796,In_1701);
or U3070 (N_3070,In_60,In_511);
and U3071 (N_3071,In_352,In_170);
xnor U3072 (N_3072,In_717,In_775);
nand U3073 (N_3073,In_500,In_1848);
nor U3074 (N_3074,In_1618,In_1496);
xor U3075 (N_3075,In_128,In_271);
and U3076 (N_3076,In_175,In_1877);
and U3077 (N_3077,In_1297,In_1129);
or U3078 (N_3078,In_1720,In_931);
and U3079 (N_3079,In_1583,In_1050);
nand U3080 (N_3080,In_31,In_601);
nor U3081 (N_3081,In_1401,In_774);
and U3082 (N_3082,In_1127,In_1795);
nor U3083 (N_3083,In_1662,In_793);
nor U3084 (N_3084,In_1466,In_368);
nor U3085 (N_3085,In_1786,In_110);
nor U3086 (N_3086,In_1446,In_1328);
nor U3087 (N_3087,In_1263,In_1966);
and U3088 (N_3088,In_644,In_1336);
nor U3089 (N_3089,In_1247,In_1528);
nand U3090 (N_3090,In_1528,In_153);
nor U3091 (N_3091,In_394,In_1740);
or U3092 (N_3092,In_1309,In_365);
nand U3093 (N_3093,In_17,In_355);
xor U3094 (N_3094,In_981,In_438);
nor U3095 (N_3095,In_1763,In_1788);
nand U3096 (N_3096,In_1621,In_302);
xnor U3097 (N_3097,In_1842,In_1354);
and U3098 (N_3098,In_169,In_1501);
nor U3099 (N_3099,In_1137,In_460);
or U3100 (N_3100,In_1903,In_1507);
or U3101 (N_3101,In_1296,In_1863);
and U3102 (N_3102,In_1599,In_427);
nor U3103 (N_3103,In_1372,In_820);
nand U3104 (N_3104,In_68,In_656);
nor U3105 (N_3105,In_563,In_496);
nor U3106 (N_3106,In_1621,In_1594);
nand U3107 (N_3107,In_17,In_1321);
nor U3108 (N_3108,In_1871,In_1481);
xor U3109 (N_3109,In_270,In_1395);
and U3110 (N_3110,In_641,In_1112);
nor U3111 (N_3111,In_432,In_1475);
xnor U3112 (N_3112,In_681,In_628);
or U3113 (N_3113,In_152,In_474);
and U3114 (N_3114,In_1897,In_935);
nand U3115 (N_3115,In_615,In_363);
nor U3116 (N_3116,In_1261,In_223);
xnor U3117 (N_3117,In_203,In_883);
and U3118 (N_3118,In_1144,In_1667);
nor U3119 (N_3119,In_1283,In_1824);
nand U3120 (N_3120,In_1792,In_1957);
and U3121 (N_3121,In_1106,In_1742);
or U3122 (N_3122,In_1996,In_1912);
and U3123 (N_3123,In_1648,In_369);
or U3124 (N_3124,In_1948,In_1767);
or U3125 (N_3125,In_58,In_727);
and U3126 (N_3126,In_297,In_1650);
and U3127 (N_3127,In_83,In_1306);
or U3128 (N_3128,In_1648,In_1434);
and U3129 (N_3129,In_230,In_1058);
xor U3130 (N_3130,In_1157,In_1034);
xor U3131 (N_3131,In_994,In_1205);
and U3132 (N_3132,In_816,In_429);
and U3133 (N_3133,In_355,In_1415);
or U3134 (N_3134,In_751,In_182);
nor U3135 (N_3135,In_1835,In_980);
xor U3136 (N_3136,In_937,In_1662);
nand U3137 (N_3137,In_1229,In_1735);
or U3138 (N_3138,In_613,In_188);
or U3139 (N_3139,In_761,In_1492);
nor U3140 (N_3140,In_812,In_765);
nor U3141 (N_3141,In_905,In_866);
and U3142 (N_3142,In_1618,In_1252);
nand U3143 (N_3143,In_196,In_1667);
nor U3144 (N_3144,In_1903,In_382);
nor U3145 (N_3145,In_1389,In_761);
nand U3146 (N_3146,In_74,In_634);
and U3147 (N_3147,In_1812,In_927);
or U3148 (N_3148,In_1398,In_1117);
or U3149 (N_3149,In_1751,In_1832);
nor U3150 (N_3150,In_647,In_1324);
nor U3151 (N_3151,In_1448,In_560);
nor U3152 (N_3152,In_1736,In_1720);
nor U3153 (N_3153,In_690,In_840);
nor U3154 (N_3154,In_1267,In_106);
nor U3155 (N_3155,In_642,In_1488);
nor U3156 (N_3156,In_1656,In_64);
nor U3157 (N_3157,In_832,In_540);
and U3158 (N_3158,In_122,In_1671);
nor U3159 (N_3159,In_303,In_1071);
nor U3160 (N_3160,In_1050,In_792);
or U3161 (N_3161,In_1892,In_1478);
nand U3162 (N_3162,In_1029,In_1497);
xor U3163 (N_3163,In_684,In_114);
or U3164 (N_3164,In_195,In_337);
nand U3165 (N_3165,In_415,In_1217);
nand U3166 (N_3166,In_1932,In_94);
and U3167 (N_3167,In_1233,In_503);
nor U3168 (N_3168,In_7,In_1214);
nand U3169 (N_3169,In_230,In_241);
xor U3170 (N_3170,In_944,In_249);
nand U3171 (N_3171,In_514,In_644);
or U3172 (N_3172,In_605,In_14);
nor U3173 (N_3173,In_778,In_391);
nand U3174 (N_3174,In_1471,In_1142);
xnor U3175 (N_3175,In_1590,In_1734);
and U3176 (N_3176,In_1731,In_162);
xnor U3177 (N_3177,In_1055,In_972);
nand U3178 (N_3178,In_2,In_646);
nand U3179 (N_3179,In_1452,In_1895);
nor U3180 (N_3180,In_1974,In_1576);
nand U3181 (N_3181,In_1648,In_1338);
or U3182 (N_3182,In_363,In_1450);
or U3183 (N_3183,In_1822,In_81);
nand U3184 (N_3184,In_700,In_1100);
nor U3185 (N_3185,In_254,In_1368);
nand U3186 (N_3186,In_684,In_957);
xor U3187 (N_3187,In_925,In_1478);
and U3188 (N_3188,In_1485,In_669);
and U3189 (N_3189,In_522,In_901);
and U3190 (N_3190,In_1355,In_1164);
nand U3191 (N_3191,In_1534,In_1484);
nor U3192 (N_3192,In_1222,In_1917);
or U3193 (N_3193,In_387,In_1882);
or U3194 (N_3194,In_1716,In_1436);
nand U3195 (N_3195,In_1296,In_1085);
nor U3196 (N_3196,In_1046,In_1771);
nand U3197 (N_3197,In_377,In_1464);
xor U3198 (N_3198,In_106,In_413);
nor U3199 (N_3199,In_262,In_1525);
nor U3200 (N_3200,In_685,In_708);
nor U3201 (N_3201,In_1614,In_995);
nor U3202 (N_3202,In_1004,In_433);
or U3203 (N_3203,In_1451,In_781);
and U3204 (N_3204,In_1040,In_1704);
and U3205 (N_3205,In_278,In_30);
and U3206 (N_3206,In_1198,In_465);
and U3207 (N_3207,In_1151,In_1731);
nor U3208 (N_3208,In_1337,In_1830);
nand U3209 (N_3209,In_285,In_1788);
and U3210 (N_3210,In_1489,In_1137);
and U3211 (N_3211,In_1197,In_342);
nor U3212 (N_3212,In_1046,In_1870);
nor U3213 (N_3213,In_856,In_1223);
nand U3214 (N_3214,In_114,In_1295);
nand U3215 (N_3215,In_1510,In_1342);
or U3216 (N_3216,In_1428,In_1005);
and U3217 (N_3217,In_397,In_1865);
nand U3218 (N_3218,In_373,In_1041);
nand U3219 (N_3219,In_867,In_1251);
or U3220 (N_3220,In_1650,In_1216);
and U3221 (N_3221,In_1325,In_169);
nor U3222 (N_3222,In_19,In_1877);
or U3223 (N_3223,In_462,In_1953);
nor U3224 (N_3224,In_679,In_601);
nor U3225 (N_3225,In_506,In_775);
and U3226 (N_3226,In_1686,In_1765);
or U3227 (N_3227,In_713,In_908);
nand U3228 (N_3228,In_1197,In_1539);
or U3229 (N_3229,In_690,In_1531);
nor U3230 (N_3230,In_1137,In_1094);
nor U3231 (N_3231,In_151,In_97);
nor U3232 (N_3232,In_1750,In_1807);
xnor U3233 (N_3233,In_1657,In_1899);
nand U3234 (N_3234,In_1065,In_754);
nor U3235 (N_3235,In_1559,In_951);
xnor U3236 (N_3236,In_395,In_1343);
nor U3237 (N_3237,In_703,In_839);
xor U3238 (N_3238,In_1837,In_1949);
and U3239 (N_3239,In_1711,In_1989);
nand U3240 (N_3240,In_20,In_404);
or U3241 (N_3241,In_1486,In_555);
nor U3242 (N_3242,In_1972,In_1997);
nand U3243 (N_3243,In_1370,In_706);
xor U3244 (N_3244,In_1707,In_325);
nand U3245 (N_3245,In_1590,In_385);
nor U3246 (N_3246,In_303,In_565);
nor U3247 (N_3247,In_886,In_1673);
and U3248 (N_3248,In_1917,In_373);
or U3249 (N_3249,In_476,In_1377);
xor U3250 (N_3250,In_1856,In_263);
or U3251 (N_3251,In_254,In_1197);
nand U3252 (N_3252,In_1701,In_1940);
nand U3253 (N_3253,In_1784,In_15);
nor U3254 (N_3254,In_125,In_1394);
nor U3255 (N_3255,In_679,In_1954);
and U3256 (N_3256,In_526,In_1744);
nor U3257 (N_3257,In_257,In_1633);
nand U3258 (N_3258,In_764,In_921);
and U3259 (N_3259,In_454,In_1212);
nor U3260 (N_3260,In_1367,In_1532);
nor U3261 (N_3261,In_1903,In_673);
and U3262 (N_3262,In_563,In_139);
and U3263 (N_3263,In_659,In_1319);
nor U3264 (N_3264,In_1577,In_616);
or U3265 (N_3265,In_853,In_1123);
nor U3266 (N_3266,In_910,In_1997);
or U3267 (N_3267,In_655,In_1463);
and U3268 (N_3268,In_1631,In_1957);
or U3269 (N_3269,In_900,In_186);
nor U3270 (N_3270,In_1210,In_439);
nor U3271 (N_3271,In_137,In_1049);
nor U3272 (N_3272,In_1415,In_1251);
and U3273 (N_3273,In_1633,In_160);
nand U3274 (N_3274,In_1870,In_1176);
nor U3275 (N_3275,In_43,In_600);
or U3276 (N_3276,In_1084,In_648);
and U3277 (N_3277,In_1530,In_1623);
and U3278 (N_3278,In_149,In_569);
nor U3279 (N_3279,In_837,In_300);
xnor U3280 (N_3280,In_1950,In_1732);
nor U3281 (N_3281,In_1715,In_49);
or U3282 (N_3282,In_1687,In_1965);
nor U3283 (N_3283,In_98,In_309);
nand U3284 (N_3284,In_10,In_783);
nand U3285 (N_3285,In_1458,In_200);
and U3286 (N_3286,In_1574,In_1381);
or U3287 (N_3287,In_1486,In_1676);
and U3288 (N_3288,In_1425,In_1382);
xor U3289 (N_3289,In_1128,In_597);
and U3290 (N_3290,In_84,In_173);
nand U3291 (N_3291,In_1369,In_1163);
or U3292 (N_3292,In_589,In_599);
nor U3293 (N_3293,In_1016,In_56);
xor U3294 (N_3294,In_1508,In_846);
nand U3295 (N_3295,In_1942,In_1675);
nand U3296 (N_3296,In_1428,In_596);
nor U3297 (N_3297,In_695,In_1728);
or U3298 (N_3298,In_902,In_641);
xnor U3299 (N_3299,In_691,In_1704);
nand U3300 (N_3300,In_866,In_355);
nand U3301 (N_3301,In_1025,In_1330);
xor U3302 (N_3302,In_1156,In_984);
nand U3303 (N_3303,In_1453,In_1499);
or U3304 (N_3304,In_1363,In_480);
or U3305 (N_3305,In_389,In_885);
nor U3306 (N_3306,In_726,In_860);
nand U3307 (N_3307,In_31,In_1571);
and U3308 (N_3308,In_1583,In_1130);
nand U3309 (N_3309,In_1507,In_504);
xnor U3310 (N_3310,In_1083,In_87);
or U3311 (N_3311,In_1438,In_1926);
and U3312 (N_3312,In_378,In_1794);
and U3313 (N_3313,In_825,In_1366);
or U3314 (N_3314,In_607,In_1178);
and U3315 (N_3315,In_1514,In_1880);
or U3316 (N_3316,In_214,In_522);
or U3317 (N_3317,In_444,In_1979);
or U3318 (N_3318,In_532,In_1656);
or U3319 (N_3319,In_1602,In_937);
nor U3320 (N_3320,In_237,In_502);
nand U3321 (N_3321,In_1811,In_1479);
nor U3322 (N_3322,In_703,In_817);
or U3323 (N_3323,In_341,In_134);
and U3324 (N_3324,In_1825,In_1452);
or U3325 (N_3325,In_1854,In_1736);
xor U3326 (N_3326,In_1488,In_1037);
nor U3327 (N_3327,In_1932,In_1333);
nor U3328 (N_3328,In_1354,In_840);
nand U3329 (N_3329,In_350,In_1808);
or U3330 (N_3330,In_473,In_253);
or U3331 (N_3331,In_448,In_533);
and U3332 (N_3332,In_1449,In_8);
xor U3333 (N_3333,In_203,In_542);
and U3334 (N_3334,In_65,In_341);
or U3335 (N_3335,In_530,In_1049);
or U3336 (N_3336,In_1213,In_442);
nand U3337 (N_3337,In_272,In_9);
xor U3338 (N_3338,In_1291,In_628);
or U3339 (N_3339,In_1852,In_960);
and U3340 (N_3340,In_694,In_1816);
or U3341 (N_3341,In_597,In_1145);
or U3342 (N_3342,In_453,In_1650);
or U3343 (N_3343,In_1307,In_1998);
and U3344 (N_3344,In_351,In_1516);
nand U3345 (N_3345,In_111,In_622);
nor U3346 (N_3346,In_549,In_226);
nor U3347 (N_3347,In_1858,In_268);
nand U3348 (N_3348,In_1134,In_1949);
and U3349 (N_3349,In_1903,In_1578);
and U3350 (N_3350,In_75,In_1762);
nor U3351 (N_3351,In_173,In_485);
or U3352 (N_3352,In_1604,In_672);
nor U3353 (N_3353,In_242,In_828);
xor U3354 (N_3354,In_1485,In_276);
or U3355 (N_3355,In_1853,In_1586);
nand U3356 (N_3356,In_1500,In_1827);
and U3357 (N_3357,In_1305,In_1835);
and U3358 (N_3358,In_182,In_1872);
or U3359 (N_3359,In_1794,In_1138);
xnor U3360 (N_3360,In_1303,In_1107);
nand U3361 (N_3361,In_1358,In_1164);
nand U3362 (N_3362,In_257,In_925);
nor U3363 (N_3363,In_964,In_1113);
or U3364 (N_3364,In_1455,In_1909);
nor U3365 (N_3365,In_738,In_856);
nor U3366 (N_3366,In_551,In_258);
nand U3367 (N_3367,In_581,In_202);
and U3368 (N_3368,In_579,In_1313);
and U3369 (N_3369,In_1458,In_842);
and U3370 (N_3370,In_1363,In_1163);
nor U3371 (N_3371,In_1788,In_1605);
and U3372 (N_3372,In_1663,In_299);
nand U3373 (N_3373,In_1655,In_1842);
xor U3374 (N_3374,In_1426,In_476);
and U3375 (N_3375,In_823,In_1129);
and U3376 (N_3376,In_1962,In_1382);
or U3377 (N_3377,In_1768,In_1092);
nand U3378 (N_3378,In_1902,In_1223);
nor U3379 (N_3379,In_444,In_150);
xor U3380 (N_3380,In_1410,In_588);
nand U3381 (N_3381,In_1543,In_1817);
nor U3382 (N_3382,In_242,In_410);
and U3383 (N_3383,In_869,In_1954);
nand U3384 (N_3384,In_538,In_887);
nor U3385 (N_3385,In_408,In_1073);
and U3386 (N_3386,In_1404,In_1153);
nand U3387 (N_3387,In_1135,In_1524);
or U3388 (N_3388,In_969,In_1637);
or U3389 (N_3389,In_1719,In_1001);
nand U3390 (N_3390,In_1353,In_1840);
or U3391 (N_3391,In_424,In_1735);
xnor U3392 (N_3392,In_1104,In_1530);
nor U3393 (N_3393,In_1021,In_1626);
xor U3394 (N_3394,In_710,In_527);
xnor U3395 (N_3395,In_1069,In_1425);
nor U3396 (N_3396,In_1616,In_249);
and U3397 (N_3397,In_114,In_1261);
nor U3398 (N_3398,In_772,In_1921);
nor U3399 (N_3399,In_275,In_1803);
nor U3400 (N_3400,In_66,In_1835);
nor U3401 (N_3401,In_1490,In_556);
nor U3402 (N_3402,In_924,In_1959);
or U3403 (N_3403,In_1442,In_1744);
and U3404 (N_3404,In_1128,In_1225);
nand U3405 (N_3405,In_466,In_1868);
or U3406 (N_3406,In_681,In_1639);
nand U3407 (N_3407,In_1417,In_801);
and U3408 (N_3408,In_318,In_909);
nor U3409 (N_3409,In_1729,In_518);
or U3410 (N_3410,In_1235,In_1963);
and U3411 (N_3411,In_953,In_1710);
nand U3412 (N_3412,In_964,In_1481);
nor U3413 (N_3413,In_1041,In_524);
nand U3414 (N_3414,In_1505,In_1527);
nor U3415 (N_3415,In_1804,In_279);
nand U3416 (N_3416,In_1098,In_411);
or U3417 (N_3417,In_1640,In_296);
and U3418 (N_3418,In_1650,In_315);
nand U3419 (N_3419,In_1181,In_93);
xnor U3420 (N_3420,In_1080,In_489);
nand U3421 (N_3421,In_1392,In_892);
nor U3422 (N_3422,In_882,In_1573);
nand U3423 (N_3423,In_956,In_1287);
and U3424 (N_3424,In_124,In_429);
nor U3425 (N_3425,In_1688,In_1653);
nand U3426 (N_3426,In_1302,In_102);
or U3427 (N_3427,In_1882,In_1732);
and U3428 (N_3428,In_362,In_970);
nor U3429 (N_3429,In_1821,In_1364);
xor U3430 (N_3430,In_1641,In_212);
nor U3431 (N_3431,In_1025,In_1843);
nand U3432 (N_3432,In_924,In_446);
nor U3433 (N_3433,In_1077,In_769);
nand U3434 (N_3434,In_1737,In_649);
xnor U3435 (N_3435,In_251,In_1272);
or U3436 (N_3436,In_1726,In_1338);
and U3437 (N_3437,In_1002,In_1691);
nand U3438 (N_3438,In_382,In_1125);
and U3439 (N_3439,In_149,In_1853);
xor U3440 (N_3440,In_1463,In_1152);
and U3441 (N_3441,In_827,In_414);
nand U3442 (N_3442,In_481,In_963);
xor U3443 (N_3443,In_947,In_1137);
or U3444 (N_3444,In_630,In_32);
nand U3445 (N_3445,In_777,In_530);
and U3446 (N_3446,In_727,In_1200);
and U3447 (N_3447,In_636,In_1732);
and U3448 (N_3448,In_23,In_1325);
nand U3449 (N_3449,In_768,In_29);
nor U3450 (N_3450,In_1949,In_1290);
or U3451 (N_3451,In_1789,In_1743);
or U3452 (N_3452,In_1713,In_1325);
or U3453 (N_3453,In_1106,In_1035);
nand U3454 (N_3454,In_1423,In_1745);
nand U3455 (N_3455,In_170,In_407);
nand U3456 (N_3456,In_301,In_942);
xnor U3457 (N_3457,In_1205,In_1378);
nand U3458 (N_3458,In_1530,In_1424);
and U3459 (N_3459,In_1420,In_131);
nor U3460 (N_3460,In_498,In_349);
and U3461 (N_3461,In_399,In_1887);
nand U3462 (N_3462,In_687,In_935);
xnor U3463 (N_3463,In_1674,In_127);
nand U3464 (N_3464,In_734,In_1377);
xnor U3465 (N_3465,In_331,In_1490);
and U3466 (N_3466,In_1475,In_1035);
nor U3467 (N_3467,In_1107,In_814);
or U3468 (N_3468,In_1230,In_1921);
and U3469 (N_3469,In_696,In_1366);
nor U3470 (N_3470,In_1119,In_592);
or U3471 (N_3471,In_615,In_906);
or U3472 (N_3472,In_1541,In_570);
nand U3473 (N_3473,In_865,In_164);
or U3474 (N_3474,In_119,In_1233);
nor U3475 (N_3475,In_416,In_1955);
or U3476 (N_3476,In_720,In_1352);
or U3477 (N_3477,In_516,In_1515);
nand U3478 (N_3478,In_1697,In_63);
nand U3479 (N_3479,In_1498,In_1680);
and U3480 (N_3480,In_1356,In_1351);
nor U3481 (N_3481,In_209,In_446);
xor U3482 (N_3482,In_150,In_1304);
nor U3483 (N_3483,In_1239,In_927);
nor U3484 (N_3484,In_1406,In_207);
nand U3485 (N_3485,In_1678,In_1901);
and U3486 (N_3486,In_1491,In_1651);
nand U3487 (N_3487,In_27,In_445);
and U3488 (N_3488,In_758,In_1603);
or U3489 (N_3489,In_1587,In_1870);
nand U3490 (N_3490,In_912,In_80);
nand U3491 (N_3491,In_1428,In_939);
nand U3492 (N_3492,In_1798,In_1251);
nor U3493 (N_3493,In_181,In_33);
nand U3494 (N_3494,In_304,In_1865);
and U3495 (N_3495,In_26,In_1101);
xor U3496 (N_3496,In_1748,In_556);
or U3497 (N_3497,In_510,In_755);
xor U3498 (N_3498,In_301,In_332);
nand U3499 (N_3499,In_698,In_1100);
nand U3500 (N_3500,In_548,In_1083);
and U3501 (N_3501,In_1003,In_34);
nand U3502 (N_3502,In_443,In_874);
nand U3503 (N_3503,In_656,In_1733);
and U3504 (N_3504,In_356,In_696);
nand U3505 (N_3505,In_1828,In_277);
and U3506 (N_3506,In_1701,In_803);
nand U3507 (N_3507,In_1990,In_1811);
nand U3508 (N_3508,In_339,In_313);
nand U3509 (N_3509,In_262,In_1089);
and U3510 (N_3510,In_1297,In_802);
nand U3511 (N_3511,In_1362,In_187);
nand U3512 (N_3512,In_387,In_692);
or U3513 (N_3513,In_1192,In_1548);
xnor U3514 (N_3514,In_1476,In_47);
nand U3515 (N_3515,In_1609,In_384);
or U3516 (N_3516,In_109,In_1932);
or U3517 (N_3517,In_1469,In_71);
and U3518 (N_3518,In_1425,In_10);
or U3519 (N_3519,In_864,In_1936);
nand U3520 (N_3520,In_614,In_1209);
and U3521 (N_3521,In_1859,In_608);
or U3522 (N_3522,In_1135,In_68);
nand U3523 (N_3523,In_1858,In_125);
nand U3524 (N_3524,In_168,In_1903);
nor U3525 (N_3525,In_1342,In_272);
nand U3526 (N_3526,In_153,In_228);
and U3527 (N_3527,In_216,In_1763);
nor U3528 (N_3528,In_1644,In_1959);
and U3529 (N_3529,In_1793,In_411);
nand U3530 (N_3530,In_721,In_326);
or U3531 (N_3531,In_990,In_1909);
and U3532 (N_3532,In_1066,In_1021);
xnor U3533 (N_3533,In_1650,In_1771);
xor U3534 (N_3534,In_1424,In_1282);
nor U3535 (N_3535,In_1328,In_1295);
nor U3536 (N_3536,In_1256,In_964);
nor U3537 (N_3537,In_1134,In_1985);
nor U3538 (N_3538,In_1102,In_9);
nand U3539 (N_3539,In_381,In_409);
nor U3540 (N_3540,In_1910,In_1091);
xnor U3541 (N_3541,In_265,In_686);
or U3542 (N_3542,In_423,In_1945);
or U3543 (N_3543,In_702,In_888);
nor U3544 (N_3544,In_203,In_1513);
and U3545 (N_3545,In_359,In_1760);
and U3546 (N_3546,In_1723,In_536);
nor U3547 (N_3547,In_1839,In_1396);
nor U3548 (N_3548,In_1926,In_861);
nand U3549 (N_3549,In_398,In_324);
or U3550 (N_3550,In_59,In_1484);
nor U3551 (N_3551,In_1907,In_1121);
nand U3552 (N_3552,In_609,In_125);
and U3553 (N_3553,In_191,In_851);
nand U3554 (N_3554,In_1965,In_1917);
and U3555 (N_3555,In_815,In_249);
or U3556 (N_3556,In_1787,In_1144);
nand U3557 (N_3557,In_692,In_823);
nor U3558 (N_3558,In_533,In_391);
xnor U3559 (N_3559,In_1724,In_418);
nor U3560 (N_3560,In_1189,In_1065);
nand U3561 (N_3561,In_296,In_1617);
nand U3562 (N_3562,In_719,In_804);
or U3563 (N_3563,In_1504,In_332);
nor U3564 (N_3564,In_1918,In_836);
and U3565 (N_3565,In_1711,In_336);
or U3566 (N_3566,In_1176,In_1829);
and U3567 (N_3567,In_183,In_1703);
nor U3568 (N_3568,In_1549,In_1714);
nand U3569 (N_3569,In_322,In_913);
or U3570 (N_3570,In_1386,In_163);
and U3571 (N_3571,In_1842,In_1390);
and U3572 (N_3572,In_316,In_439);
nor U3573 (N_3573,In_1276,In_261);
nand U3574 (N_3574,In_827,In_1510);
nor U3575 (N_3575,In_194,In_1436);
nor U3576 (N_3576,In_250,In_752);
and U3577 (N_3577,In_144,In_1595);
nor U3578 (N_3578,In_1333,In_133);
nand U3579 (N_3579,In_1732,In_709);
nor U3580 (N_3580,In_1331,In_998);
and U3581 (N_3581,In_154,In_292);
xnor U3582 (N_3582,In_1200,In_1437);
and U3583 (N_3583,In_1215,In_445);
or U3584 (N_3584,In_700,In_765);
and U3585 (N_3585,In_926,In_520);
and U3586 (N_3586,In_332,In_1445);
nor U3587 (N_3587,In_655,In_971);
or U3588 (N_3588,In_1210,In_1475);
nor U3589 (N_3589,In_1039,In_1989);
or U3590 (N_3590,In_1022,In_1081);
or U3591 (N_3591,In_224,In_692);
nand U3592 (N_3592,In_983,In_291);
or U3593 (N_3593,In_874,In_1997);
or U3594 (N_3594,In_777,In_1539);
nand U3595 (N_3595,In_944,In_31);
nand U3596 (N_3596,In_1453,In_1340);
or U3597 (N_3597,In_579,In_1483);
nand U3598 (N_3598,In_643,In_1615);
and U3599 (N_3599,In_1596,In_1127);
nor U3600 (N_3600,In_1342,In_325);
or U3601 (N_3601,In_1953,In_89);
or U3602 (N_3602,In_1275,In_1509);
nand U3603 (N_3603,In_1869,In_735);
and U3604 (N_3604,In_618,In_1253);
nand U3605 (N_3605,In_902,In_274);
or U3606 (N_3606,In_1012,In_1314);
and U3607 (N_3607,In_746,In_286);
nand U3608 (N_3608,In_159,In_633);
or U3609 (N_3609,In_70,In_888);
nand U3610 (N_3610,In_1916,In_787);
nor U3611 (N_3611,In_1522,In_1910);
nand U3612 (N_3612,In_912,In_1810);
or U3613 (N_3613,In_597,In_785);
nand U3614 (N_3614,In_1825,In_1105);
xor U3615 (N_3615,In_984,In_1476);
xor U3616 (N_3616,In_95,In_101);
nor U3617 (N_3617,In_87,In_789);
nand U3618 (N_3618,In_401,In_1321);
and U3619 (N_3619,In_1303,In_1361);
nor U3620 (N_3620,In_1985,In_228);
nor U3621 (N_3621,In_1335,In_691);
and U3622 (N_3622,In_1962,In_1230);
nor U3623 (N_3623,In_595,In_388);
nor U3624 (N_3624,In_1633,In_256);
nand U3625 (N_3625,In_941,In_1251);
and U3626 (N_3626,In_656,In_135);
and U3627 (N_3627,In_1746,In_1968);
nor U3628 (N_3628,In_1919,In_1143);
or U3629 (N_3629,In_1427,In_1753);
nor U3630 (N_3630,In_706,In_1288);
or U3631 (N_3631,In_1872,In_596);
nor U3632 (N_3632,In_1080,In_1843);
nand U3633 (N_3633,In_967,In_834);
nand U3634 (N_3634,In_1938,In_1072);
xnor U3635 (N_3635,In_1566,In_327);
nand U3636 (N_3636,In_1721,In_1609);
and U3637 (N_3637,In_1622,In_952);
and U3638 (N_3638,In_1093,In_701);
or U3639 (N_3639,In_707,In_206);
or U3640 (N_3640,In_1762,In_904);
or U3641 (N_3641,In_1445,In_145);
or U3642 (N_3642,In_223,In_315);
and U3643 (N_3643,In_1226,In_782);
or U3644 (N_3644,In_1218,In_199);
or U3645 (N_3645,In_1807,In_1201);
nor U3646 (N_3646,In_1074,In_30);
nor U3647 (N_3647,In_1923,In_1476);
and U3648 (N_3648,In_1365,In_900);
xnor U3649 (N_3649,In_885,In_201);
or U3650 (N_3650,In_1358,In_1870);
and U3651 (N_3651,In_1736,In_971);
xnor U3652 (N_3652,In_359,In_1830);
nand U3653 (N_3653,In_1472,In_1773);
or U3654 (N_3654,In_996,In_1578);
nor U3655 (N_3655,In_584,In_403);
nor U3656 (N_3656,In_1561,In_774);
nor U3657 (N_3657,In_1227,In_1702);
nor U3658 (N_3658,In_1646,In_1493);
and U3659 (N_3659,In_918,In_455);
nand U3660 (N_3660,In_147,In_424);
xnor U3661 (N_3661,In_1210,In_1079);
nand U3662 (N_3662,In_576,In_586);
nand U3663 (N_3663,In_319,In_647);
nor U3664 (N_3664,In_1835,In_95);
nand U3665 (N_3665,In_1538,In_488);
or U3666 (N_3666,In_1059,In_1406);
and U3667 (N_3667,In_809,In_1083);
and U3668 (N_3668,In_1692,In_1412);
or U3669 (N_3669,In_1333,In_945);
and U3670 (N_3670,In_1137,In_727);
and U3671 (N_3671,In_929,In_542);
nor U3672 (N_3672,In_1885,In_269);
nor U3673 (N_3673,In_652,In_1274);
and U3674 (N_3674,In_494,In_1986);
or U3675 (N_3675,In_27,In_1557);
nand U3676 (N_3676,In_827,In_985);
and U3677 (N_3677,In_1392,In_1935);
xnor U3678 (N_3678,In_166,In_930);
nor U3679 (N_3679,In_981,In_1055);
or U3680 (N_3680,In_82,In_1337);
xor U3681 (N_3681,In_1923,In_1984);
nand U3682 (N_3682,In_1976,In_278);
nand U3683 (N_3683,In_1702,In_1383);
and U3684 (N_3684,In_527,In_1367);
nand U3685 (N_3685,In_1977,In_1326);
nand U3686 (N_3686,In_1600,In_387);
and U3687 (N_3687,In_1020,In_378);
or U3688 (N_3688,In_1975,In_1441);
nand U3689 (N_3689,In_1775,In_688);
xnor U3690 (N_3690,In_1132,In_421);
nor U3691 (N_3691,In_1699,In_1469);
nand U3692 (N_3692,In_1819,In_287);
nand U3693 (N_3693,In_1322,In_629);
and U3694 (N_3694,In_14,In_327);
or U3695 (N_3695,In_631,In_493);
and U3696 (N_3696,In_197,In_808);
and U3697 (N_3697,In_1033,In_1221);
nand U3698 (N_3698,In_1377,In_1453);
or U3699 (N_3699,In_1062,In_183);
nand U3700 (N_3700,In_1576,In_254);
or U3701 (N_3701,In_1083,In_793);
and U3702 (N_3702,In_38,In_447);
xor U3703 (N_3703,In_11,In_491);
and U3704 (N_3704,In_1157,In_1594);
xnor U3705 (N_3705,In_215,In_866);
and U3706 (N_3706,In_523,In_753);
nand U3707 (N_3707,In_1015,In_784);
nand U3708 (N_3708,In_1093,In_519);
or U3709 (N_3709,In_772,In_1893);
nand U3710 (N_3710,In_660,In_539);
nand U3711 (N_3711,In_1085,In_1168);
or U3712 (N_3712,In_1928,In_833);
xnor U3713 (N_3713,In_624,In_637);
nand U3714 (N_3714,In_1426,In_777);
or U3715 (N_3715,In_1818,In_1964);
nand U3716 (N_3716,In_1839,In_363);
nand U3717 (N_3717,In_1809,In_1135);
nor U3718 (N_3718,In_343,In_1250);
and U3719 (N_3719,In_72,In_570);
xnor U3720 (N_3720,In_56,In_320);
xnor U3721 (N_3721,In_1026,In_1935);
or U3722 (N_3722,In_660,In_747);
and U3723 (N_3723,In_899,In_1207);
or U3724 (N_3724,In_173,In_417);
xnor U3725 (N_3725,In_1729,In_165);
xor U3726 (N_3726,In_772,In_269);
nand U3727 (N_3727,In_871,In_342);
nor U3728 (N_3728,In_992,In_1953);
nor U3729 (N_3729,In_1279,In_489);
nand U3730 (N_3730,In_164,In_1504);
nand U3731 (N_3731,In_464,In_269);
and U3732 (N_3732,In_1497,In_1624);
or U3733 (N_3733,In_794,In_1476);
nor U3734 (N_3734,In_723,In_1679);
nand U3735 (N_3735,In_440,In_1656);
nand U3736 (N_3736,In_1526,In_168);
nand U3737 (N_3737,In_425,In_1922);
and U3738 (N_3738,In_866,In_1059);
and U3739 (N_3739,In_1294,In_1322);
and U3740 (N_3740,In_835,In_462);
nor U3741 (N_3741,In_1195,In_1085);
nor U3742 (N_3742,In_1075,In_1243);
xnor U3743 (N_3743,In_558,In_1213);
nor U3744 (N_3744,In_1116,In_474);
or U3745 (N_3745,In_1431,In_1284);
and U3746 (N_3746,In_1809,In_156);
xor U3747 (N_3747,In_1668,In_1491);
or U3748 (N_3748,In_778,In_1266);
nand U3749 (N_3749,In_1444,In_1926);
or U3750 (N_3750,In_967,In_218);
nand U3751 (N_3751,In_1967,In_120);
or U3752 (N_3752,In_296,In_234);
nand U3753 (N_3753,In_1872,In_1409);
xnor U3754 (N_3754,In_267,In_1516);
xnor U3755 (N_3755,In_915,In_839);
and U3756 (N_3756,In_1842,In_1400);
nand U3757 (N_3757,In_883,In_490);
nor U3758 (N_3758,In_1602,In_542);
nor U3759 (N_3759,In_1603,In_744);
nand U3760 (N_3760,In_1105,In_1388);
or U3761 (N_3761,In_1822,In_530);
nand U3762 (N_3762,In_1451,In_872);
or U3763 (N_3763,In_313,In_1760);
xnor U3764 (N_3764,In_128,In_177);
or U3765 (N_3765,In_816,In_133);
nor U3766 (N_3766,In_1952,In_1273);
nand U3767 (N_3767,In_1234,In_907);
nor U3768 (N_3768,In_1742,In_755);
nor U3769 (N_3769,In_1763,In_273);
xnor U3770 (N_3770,In_1460,In_444);
and U3771 (N_3771,In_1185,In_759);
nand U3772 (N_3772,In_1773,In_341);
nand U3773 (N_3773,In_614,In_1675);
and U3774 (N_3774,In_1559,In_1826);
nand U3775 (N_3775,In_1279,In_131);
or U3776 (N_3776,In_1851,In_952);
and U3777 (N_3777,In_730,In_527);
nor U3778 (N_3778,In_28,In_501);
or U3779 (N_3779,In_1351,In_1462);
and U3780 (N_3780,In_1083,In_1434);
nor U3781 (N_3781,In_1243,In_1822);
and U3782 (N_3782,In_1936,In_1084);
nand U3783 (N_3783,In_1425,In_950);
and U3784 (N_3784,In_1415,In_824);
nand U3785 (N_3785,In_425,In_1517);
or U3786 (N_3786,In_6,In_96);
nor U3787 (N_3787,In_875,In_654);
and U3788 (N_3788,In_1389,In_1552);
nand U3789 (N_3789,In_1340,In_1842);
nor U3790 (N_3790,In_751,In_812);
nor U3791 (N_3791,In_347,In_1218);
nand U3792 (N_3792,In_1422,In_990);
and U3793 (N_3793,In_1222,In_441);
nor U3794 (N_3794,In_1174,In_250);
nand U3795 (N_3795,In_668,In_682);
and U3796 (N_3796,In_1107,In_37);
or U3797 (N_3797,In_121,In_524);
nand U3798 (N_3798,In_759,In_260);
xnor U3799 (N_3799,In_1441,In_5);
xnor U3800 (N_3800,In_1731,In_713);
and U3801 (N_3801,In_1057,In_1244);
and U3802 (N_3802,In_1061,In_536);
and U3803 (N_3803,In_1798,In_928);
or U3804 (N_3804,In_787,In_1690);
or U3805 (N_3805,In_5,In_664);
or U3806 (N_3806,In_1205,In_1943);
xor U3807 (N_3807,In_443,In_1696);
nor U3808 (N_3808,In_1534,In_598);
nor U3809 (N_3809,In_433,In_1279);
or U3810 (N_3810,In_22,In_1561);
or U3811 (N_3811,In_1036,In_381);
nor U3812 (N_3812,In_453,In_1668);
nand U3813 (N_3813,In_533,In_1153);
nor U3814 (N_3814,In_455,In_1911);
and U3815 (N_3815,In_258,In_1938);
nand U3816 (N_3816,In_707,In_1186);
xor U3817 (N_3817,In_1347,In_919);
xor U3818 (N_3818,In_289,In_1769);
nor U3819 (N_3819,In_222,In_353);
nor U3820 (N_3820,In_562,In_1735);
and U3821 (N_3821,In_1247,In_1695);
xor U3822 (N_3822,In_93,In_150);
and U3823 (N_3823,In_650,In_245);
nor U3824 (N_3824,In_1695,In_935);
xor U3825 (N_3825,In_1305,In_859);
and U3826 (N_3826,In_1603,In_1983);
and U3827 (N_3827,In_560,In_1826);
nor U3828 (N_3828,In_823,In_1326);
nor U3829 (N_3829,In_1567,In_953);
xnor U3830 (N_3830,In_1445,In_1538);
nor U3831 (N_3831,In_1964,In_1402);
nor U3832 (N_3832,In_1319,In_1789);
and U3833 (N_3833,In_1007,In_909);
nor U3834 (N_3834,In_1201,In_582);
nand U3835 (N_3835,In_878,In_1060);
xnor U3836 (N_3836,In_745,In_22);
and U3837 (N_3837,In_1954,In_1799);
or U3838 (N_3838,In_1400,In_833);
nor U3839 (N_3839,In_1601,In_121);
and U3840 (N_3840,In_567,In_1271);
or U3841 (N_3841,In_1743,In_1868);
and U3842 (N_3842,In_81,In_604);
nand U3843 (N_3843,In_227,In_888);
xor U3844 (N_3844,In_1155,In_924);
or U3845 (N_3845,In_544,In_1672);
nand U3846 (N_3846,In_580,In_385);
or U3847 (N_3847,In_1556,In_463);
and U3848 (N_3848,In_693,In_1107);
or U3849 (N_3849,In_1466,In_883);
nand U3850 (N_3850,In_180,In_126);
or U3851 (N_3851,In_1967,In_1110);
nor U3852 (N_3852,In_1588,In_615);
xnor U3853 (N_3853,In_1077,In_377);
xor U3854 (N_3854,In_607,In_64);
and U3855 (N_3855,In_1352,In_657);
or U3856 (N_3856,In_492,In_1517);
or U3857 (N_3857,In_162,In_1668);
and U3858 (N_3858,In_127,In_319);
nor U3859 (N_3859,In_438,In_1214);
and U3860 (N_3860,In_583,In_134);
or U3861 (N_3861,In_918,In_495);
xnor U3862 (N_3862,In_1345,In_536);
nor U3863 (N_3863,In_325,In_1526);
nand U3864 (N_3864,In_714,In_1912);
nand U3865 (N_3865,In_1799,In_1756);
nor U3866 (N_3866,In_911,In_1280);
and U3867 (N_3867,In_1774,In_1486);
nor U3868 (N_3868,In_582,In_514);
or U3869 (N_3869,In_1700,In_631);
nand U3870 (N_3870,In_874,In_432);
nor U3871 (N_3871,In_1882,In_1272);
or U3872 (N_3872,In_277,In_640);
nand U3873 (N_3873,In_1655,In_506);
nand U3874 (N_3874,In_129,In_1236);
nor U3875 (N_3875,In_238,In_1844);
nand U3876 (N_3876,In_1457,In_327);
nand U3877 (N_3877,In_1199,In_914);
nand U3878 (N_3878,In_186,In_1867);
and U3879 (N_3879,In_868,In_1523);
nor U3880 (N_3880,In_1737,In_551);
nand U3881 (N_3881,In_1164,In_504);
xnor U3882 (N_3882,In_1334,In_788);
nor U3883 (N_3883,In_316,In_1458);
or U3884 (N_3884,In_1270,In_394);
or U3885 (N_3885,In_1572,In_332);
and U3886 (N_3886,In_109,In_1561);
nand U3887 (N_3887,In_1608,In_1567);
nand U3888 (N_3888,In_1176,In_743);
or U3889 (N_3889,In_378,In_999);
or U3890 (N_3890,In_634,In_1965);
nor U3891 (N_3891,In_574,In_1812);
xnor U3892 (N_3892,In_1687,In_168);
xnor U3893 (N_3893,In_1802,In_1043);
and U3894 (N_3894,In_609,In_548);
or U3895 (N_3895,In_256,In_215);
nor U3896 (N_3896,In_884,In_10);
nand U3897 (N_3897,In_415,In_764);
nor U3898 (N_3898,In_688,In_14);
nand U3899 (N_3899,In_219,In_98);
nor U3900 (N_3900,In_1902,In_65);
nor U3901 (N_3901,In_123,In_1419);
nand U3902 (N_3902,In_210,In_54);
nor U3903 (N_3903,In_1994,In_1730);
nor U3904 (N_3904,In_1528,In_1716);
or U3905 (N_3905,In_536,In_827);
and U3906 (N_3906,In_596,In_701);
nand U3907 (N_3907,In_526,In_1224);
nand U3908 (N_3908,In_178,In_435);
nor U3909 (N_3909,In_122,In_772);
nor U3910 (N_3910,In_138,In_1537);
xor U3911 (N_3911,In_1891,In_723);
xnor U3912 (N_3912,In_1024,In_1746);
or U3913 (N_3913,In_713,In_1548);
or U3914 (N_3914,In_858,In_1531);
or U3915 (N_3915,In_1300,In_201);
and U3916 (N_3916,In_718,In_1791);
nand U3917 (N_3917,In_1070,In_1346);
or U3918 (N_3918,In_463,In_1114);
nor U3919 (N_3919,In_825,In_334);
nand U3920 (N_3920,In_1861,In_829);
xor U3921 (N_3921,In_1703,In_1807);
and U3922 (N_3922,In_605,In_1171);
and U3923 (N_3923,In_799,In_1647);
nor U3924 (N_3924,In_110,In_812);
nor U3925 (N_3925,In_134,In_1686);
nand U3926 (N_3926,In_213,In_1932);
nor U3927 (N_3927,In_774,In_1876);
nor U3928 (N_3928,In_788,In_769);
or U3929 (N_3929,In_1304,In_890);
nor U3930 (N_3930,In_1007,In_617);
xnor U3931 (N_3931,In_1183,In_1565);
nor U3932 (N_3932,In_531,In_1377);
nand U3933 (N_3933,In_1015,In_1908);
xnor U3934 (N_3934,In_1748,In_1825);
nor U3935 (N_3935,In_1320,In_1938);
xor U3936 (N_3936,In_419,In_1719);
and U3937 (N_3937,In_346,In_1708);
or U3938 (N_3938,In_1828,In_1203);
or U3939 (N_3939,In_498,In_1120);
nor U3940 (N_3940,In_965,In_1589);
nor U3941 (N_3941,In_1993,In_651);
nand U3942 (N_3942,In_1110,In_990);
nand U3943 (N_3943,In_684,In_232);
nor U3944 (N_3944,In_912,In_435);
nor U3945 (N_3945,In_1887,In_240);
nand U3946 (N_3946,In_790,In_1533);
nand U3947 (N_3947,In_175,In_1307);
and U3948 (N_3948,In_231,In_273);
or U3949 (N_3949,In_56,In_1560);
xnor U3950 (N_3950,In_1812,In_34);
nor U3951 (N_3951,In_961,In_1182);
nand U3952 (N_3952,In_166,In_1035);
and U3953 (N_3953,In_105,In_1564);
or U3954 (N_3954,In_1775,In_707);
or U3955 (N_3955,In_71,In_1849);
nand U3956 (N_3956,In_1131,In_1903);
or U3957 (N_3957,In_1501,In_1869);
xnor U3958 (N_3958,In_750,In_1993);
nand U3959 (N_3959,In_731,In_1991);
nor U3960 (N_3960,In_1466,In_1189);
xnor U3961 (N_3961,In_1190,In_1671);
nor U3962 (N_3962,In_1666,In_1903);
or U3963 (N_3963,In_1504,In_75);
nor U3964 (N_3964,In_345,In_1509);
and U3965 (N_3965,In_1112,In_1441);
and U3966 (N_3966,In_1397,In_941);
and U3967 (N_3967,In_1077,In_834);
nand U3968 (N_3968,In_1941,In_757);
and U3969 (N_3969,In_1311,In_1168);
or U3970 (N_3970,In_240,In_1620);
and U3971 (N_3971,In_1568,In_1014);
or U3972 (N_3972,In_1178,In_1136);
nor U3973 (N_3973,In_1808,In_266);
nand U3974 (N_3974,In_1246,In_1984);
or U3975 (N_3975,In_1420,In_1752);
and U3976 (N_3976,In_636,In_714);
xnor U3977 (N_3977,In_1857,In_30);
nor U3978 (N_3978,In_1016,In_405);
nand U3979 (N_3979,In_906,In_742);
and U3980 (N_3980,In_704,In_1785);
or U3981 (N_3981,In_703,In_1018);
xnor U3982 (N_3982,In_1390,In_1397);
nor U3983 (N_3983,In_1247,In_255);
or U3984 (N_3984,In_967,In_731);
nor U3985 (N_3985,In_596,In_9);
nor U3986 (N_3986,In_433,In_1383);
or U3987 (N_3987,In_938,In_79);
and U3988 (N_3988,In_100,In_1216);
nor U3989 (N_3989,In_157,In_388);
and U3990 (N_3990,In_955,In_1758);
or U3991 (N_3991,In_336,In_942);
nor U3992 (N_3992,In_1520,In_133);
nor U3993 (N_3993,In_1813,In_866);
nor U3994 (N_3994,In_1677,In_1191);
and U3995 (N_3995,In_167,In_1671);
nor U3996 (N_3996,In_167,In_194);
or U3997 (N_3997,In_1835,In_1798);
or U3998 (N_3998,In_738,In_1578);
and U3999 (N_3999,In_573,In_1441);
xor U4000 (N_4000,N_2146,N_2528);
and U4001 (N_4001,N_456,N_2416);
nor U4002 (N_4002,N_1137,N_306);
nand U4003 (N_4003,N_2678,N_1939);
and U4004 (N_4004,N_214,N_3946);
xnor U4005 (N_4005,N_2210,N_3276);
nor U4006 (N_4006,N_2233,N_1722);
xnor U4007 (N_4007,N_3610,N_2921);
xor U4008 (N_4008,N_3599,N_1719);
or U4009 (N_4009,N_3872,N_3302);
or U4010 (N_4010,N_1111,N_2641);
and U4011 (N_4011,N_3836,N_1063);
or U4012 (N_4012,N_2190,N_3125);
or U4013 (N_4013,N_1817,N_1399);
or U4014 (N_4014,N_3981,N_3719);
nor U4015 (N_4015,N_3265,N_3029);
or U4016 (N_4016,N_2097,N_2972);
and U4017 (N_4017,N_2846,N_569);
and U4018 (N_4018,N_3631,N_3925);
and U4019 (N_4019,N_2005,N_3195);
xnor U4020 (N_4020,N_2477,N_1158);
nor U4021 (N_4021,N_136,N_1061);
and U4022 (N_4022,N_3950,N_86);
and U4023 (N_4023,N_2086,N_2610);
nand U4024 (N_4024,N_1733,N_3673);
or U4025 (N_4025,N_2742,N_2721);
and U4026 (N_4026,N_2628,N_958);
nand U4027 (N_4027,N_474,N_2926);
xor U4028 (N_4028,N_797,N_3198);
xor U4029 (N_4029,N_826,N_653);
or U4030 (N_4030,N_2383,N_230);
nor U4031 (N_4031,N_3965,N_768);
nor U4032 (N_4032,N_2163,N_3565);
nand U4033 (N_4033,N_528,N_1544);
or U4034 (N_4034,N_3654,N_130);
nor U4035 (N_4035,N_2540,N_3736);
nor U4036 (N_4036,N_3475,N_240);
nand U4037 (N_4037,N_2031,N_184);
xnor U4038 (N_4038,N_1262,N_1041);
nand U4039 (N_4039,N_2506,N_3114);
and U4040 (N_4040,N_2410,N_457);
xor U4041 (N_4041,N_767,N_2239);
nand U4042 (N_4042,N_3735,N_786);
or U4043 (N_4043,N_2343,N_1883);
nand U4044 (N_4044,N_1547,N_1049);
or U4045 (N_4045,N_1796,N_1223);
nor U4046 (N_4046,N_2384,N_175);
nand U4047 (N_4047,N_1365,N_281);
nand U4048 (N_4048,N_2437,N_3293);
nor U4049 (N_4049,N_720,N_1104);
or U4050 (N_4050,N_1983,N_3374);
xor U4051 (N_4051,N_58,N_3556);
xor U4052 (N_4052,N_100,N_2870);
nor U4053 (N_4053,N_3847,N_84);
nor U4054 (N_4054,N_2445,N_2228);
nand U4055 (N_4055,N_3839,N_2231);
and U4056 (N_4056,N_944,N_3510);
nor U4057 (N_4057,N_3319,N_341);
xor U4058 (N_4058,N_424,N_360);
and U4059 (N_4059,N_2762,N_1911);
nor U4060 (N_4060,N_2739,N_202);
and U4061 (N_4061,N_2668,N_3248);
or U4062 (N_4062,N_2254,N_1220);
or U4063 (N_4063,N_1383,N_2131);
and U4064 (N_4064,N_237,N_2130);
or U4065 (N_4065,N_3324,N_2043);
xnor U4066 (N_4066,N_2327,N_2861);
nand U4067 (N_4067,N_323,N_1283);
nand U4068 (N_4068,N_531,N_637);
nand U4069 (N_4069,N_1991,N_3030);
or U4070 (N_4070,N_3376,N_3746);
nand U4071 (N_4071,N_1357,N_254);
nand U4072 (N_4072,N_3653,N_579);
and U4073 (N_4073,N_1607,N_835);
or U4074 (N_4074,N_2838,N_3273);
nand U4075 (N_4075,N_3521,N_1067);
nand U4076 (N_4076,N_3009,N_3717);
nor U4077 (N_4077,N_2138,N_1336);
nand U4078 (N_4078,N_3795,N_2497);
or U4079 (N_4079,N_769,N_3621);
nand U4080 (N_4080,N_1881,N_1597);
nor U4081 (N_4081,N_3811,N_1844);
or U4082 (N_4082,N_745,N_1624);
xnor U4083 (N_4083,N_3512,N_3091);
nor U4084 (N_4084,N_556,N_3724);
nand U4085 (N_4085,N_3650,N_2457);
nand U4086 (N_4086,N_2105,N_978);
nor U4087 (N_4087,N_146,N_1350);
or U4088 (N_4088,N_2348,N_3691);
nor U4089 (N_4089,N_44,N_3874);
nor U4090 (N_4090,N_2609,N_1615);
or U4091 (N_4091,N_1435,N_1054);
nand U4092 (N_4092,N_2229,N_305);
or U4093 (N_4093,N_2554,N_1601);
and U4094 (N_4094,N_1484,N_1277);
and U4095 (N_4095,N_3220,N_664);
or U4096 (N_4096,N_2639,N_178);
and U4097 (N_4097,N_2749,N_3917);
nor U4098 (N_4098,N_1402,N_1211);
or U4099 (N_4099,N_477,N_918);
nor U4100 (N_4100,N_3619,N_2682);
and U4101 (N_4101,N_3812,N_3956);
xnor U4102 (N_4102,N_206,N_2605);
and U4103 (N_4103,N_1746,N_744);
xor U4104 (N_4104,N_2142,N_3860);
xnor U4105 (N_4105,N_3484,N_1929);
and U4106 (N_4106,N_296,N_1910);
and U4107 (N_4107,N_431,N_1860);
and U4108 (N_4108,N_2774,N_1015);
or U4109 (N_4109,N_45,N_1315);
nand U4110 (N_4110,N_1927,N_3543);
or U4111 (N_4111,N_1534,N_1055);
nand U4112 (N_4112,N_3715,N_1856);
nand U4113 (N_4113,N_2932,N_3012);
nor U4114 (N_4114,N_2746,N_1421);
or U4115 (N_4115,N_1135,N_3841);
and U4116 (N_4116,N_981,N_1393);
nand U4117 (N_4117,N_452,N_1821);
and U4118 (N_4118,N_3678,N_3122);
or U4119 (N_4119,N_1620,N_2355);
nor U4120 (N_4120,N_80,N_659);
or U4121 (N_4121,N_3323,N_2145);
or U4122 (N_4122,N_656,N_920);
or U4123 (N_4123,N_480,N_253);
xnor U4124 (N_4124,N_1070,N_954);
nand U4125 (N_4125,N_3140,N_2127);
or U4126 (N_4126,N_3796,N_3723);
or U4127 (N_4127,N_2614,N_1450);
nor U4128 (N_4128,N_3716,N_148);
or U4129 (N_4129,N_1784,N_3926);
nand U4130 (N_4130,N_1314,N_987);
or U4131 (N_4131,N_753,N_1014);
and U4132 (N_4132,N_875,N_1537);
or U4133 (N_4133,N_3077,N_1012);
or U4134 (N_4134,N_2096,N_2957);
and U4135 (N_4135,N_1605,N_3571);
nand U4136 (N_4136,N_1129,N_1596);
nor U4137 (N_4137,N_173,N_1662);
nand U4138 (N_4138,N_677,N_3005);
or U4139 (N_4139,N_1587,N_3267);
and U4140 (N_4140,N_646,N_370);
and U4141 (N_4141,N_2057,N_1665);
or U4142 (N_4142,N_1433,N_2652);
xnor U4143 (N_4143,N_1107,N_510);
nand U4144 (N_4144,N_1849,N_937);
and U4145 (N_4145,N_3883,N_3710);
nand U4146 (N_4146,N_3328,N_1275);
nor U4147 (N_4147,N_3632,N_3525);
or U4148 (N_4148,N_3279,N_1706);
and U4149 (N_4149,N_2322,N_1907);
or U4150 (N_4150,N_1338,N_3640);
and U4151 (N_4151,N_3814,N_668);
nand U4152 (N_4152,N_624,N_2435);
or U4153 (N_4153,N_3615,N_2430);
nor U4154 (N_4154,N_1294,N_3603);
and U4155 (N_4155,N_1538,N_427);
and U4156 (N_4156,N_640,N_1533);
and U4157 (N_4157,N_1021,N_3297);
or U4158 (N_4158,N_1467,N_3780);
nor U4159 (N_4159,N_1906,N_817);
or U4160 (N_4160,N_837,N_3730);
xnor U4161 (N_4161,N_549,N_1942);
nor U4162 (N_4162,N_3858,N_3407);
xor U4163 (N_4163,N_2001,N_1606);
or U4164 (N_4164,N_164,N_3851);
nand U4165 (N_4165,N_3581,N_550);
nor U4166 (N_4166,N_3585,N_1678);
xor U4167 (N_4167,N_662,N_2905);
nand U4168 (N_4168,N_1403,N_2177);
nor U4169 (N_4169,N_2770,N_772);
or U4170 (N_4170,N_3333,N_792);
and U4171 (N_4171,N_523,N_1663);
xnor U4172 (N_4172,N_3213,N_268);
and U4173 (N_4173,N_2321,N_911);
xnor U4174 (N_4174,N_1480,N_3771);
nand U4175 (N_4175,N_407,N_3164);
nor U4176 (N_4176,N_1398,N_2842);
nor U4177 (N_4177,N_2007,N_398);
nor U4178 (N_4178,N_1683,N_2829);
and U4179 (N_4179,N_1506,N_2387);
xor U4180 (N_4180,N_2029,N_1311);
and U4181 (N_4181,N_329,N_3762);
xor U4182 (N_4182,N_2629,N_2663);
or U4183 (N_4183,N_3306,N_2673);
xor U4184 (N_4184,N_3568,N_2850);
or U4185 (N_4185,N_3961,N_3313);
or U4186 (N_4186,N_3573,N_1236);
or U4187 (N_4187,N_1831,N_2755);
nor U4188 (N_4188,N_124,N_1751);
and U4189 (N_4189,N_3178,N_91);
nand U4190 (N_4190,N_2253,N_1859);
nor U4191 (N_4191,N_1951,N_2356);
nor U4192 (N_4192,N_3111,N_2169);
nor U4193 (N_4193,N_1543,N_3425);
nor U4194 (N_4194,N_1391,N_215);
nor U4195 (N_4195,N_983,N_3531);
or U4196 (N_4196,N_447,N_261);
nand U4197 (N_4197,N_2998,N_3873);
nand U4198 (N_4198,N_81,N_3238);
nor U4199 (N_4199,N_3138,N_2333);
or U4200 (N_4200,N_984,N_1224);
nor U4201 (N_4201,N_256,N_168);
and U4202 (N_4202,N_3576,N_3927);
nor U4203 (N_4203,N_1594,N_3738);
and U4204 (N_4204,N_1717,N_503);
xnor U4205 (N_4205,N_1572,N_2840);
and U4206 (N_4206,N_1657,N_3344);
nor U4207 (N_4207,N_2709,N_3522);
and U4208 (N_4208,N_2391,N_3509);
or U4209 (N_4209,N_3021,N_3907);
nor U4210 (N_4210,N_66,N_3101);
nand U4211 (N_4211,N_2699,N_3127);
nor U4212 (N_4212,N_2794,N_2808);
xnor U4213 (N_4213,N_3123,N_3642);
nor U4214 (N_4214,N_2273,N_2517);
xnor U4215 (N_4215,N_3897,N_1812);
nand U4216 (N_4216,N_2837,N_139);
nand U4217 (N_4217,N_2771,N_3283);
nand U4218 (N_4218,N_3161,N_2366);
nor U4219 (N_4219,N_1164,N_3998);
and U4220 (N_4220,N_2727,N_1968);
nand U4221 (N_4221,N_2452,N_2319);
and U4222 (N_4222,N_3758,N_1240);
nand U4223 (N_4223,N_2637,N_2519);
xnor U4224 (N_4224,N_227,N_1469);
or U4225 (N_4225,N_2582,N_2294);
nand U4226 (N_4226,N_904,N_1031);
nand U4227 (N_4227,N_1121,N_1271);
and U4228 (N_4228,N_3356,N_3886);
nand U4229 (N_4229,N_259,N_845);
nand U4230 (N_4230,N_2732,N_3815);
and U4231 (N_4231,N_2764,N_2286);
nand U4232 (N_4232,N_2157,N_2221);
nor U4233 (N_4233,N_3172,N_2607);
or U4234 (N_4234,N_3166,N_2378);
or U4235 (N_4235,N_2397,N_1380);
and U4236 (N_4236,N_1855,N_1837);
or U4237 (N_4237,N_383,N_538);
and U4238 (N_4238,N_1059,N_2351);
nor U4239 (N_4239,N_338,N_1892);
or U4240 (N_4240,N_3508,N_1950);
xnor U4241 (N_4241,N_3018,N_2219);
xor U4242 (N_4242,N_763,N_1475);
and U4243 (N_4243,N_1716,N_437);
and U4244 (N_4244,N_455,N_3613);
and U4245 (N_4245,N_3277,N_3084);
nand U4246 (N_4246,N_7,N_1081);
xor U4247 (N_4247,N_1161,N_881);
nor U4248 (N_4248,N_1612,N_243);
nand U4249 (N_4249,N_2274,N_3517);
nor U4250 (N_4250,N_1962,N_2234);
xor U4251 (N_4251,N_743,N_1576);
xor U4252 (N_4252,N_1813,N_2046);
nand U4253 (N_4253,N_3970,N_2396);
and U4254 (N_4254,N_2661,N_3402);
and U4255 (N_4255,N_2667,N_964);
nand U4256 (N_4256,N_3523,N_2217);
or U4257 (N_4257,N_1590,N_687);
nor U4258 (N_4258,N_2899,N_1546);
nand U4259 (N_4259,N_3808,N_2913);
xor U4260 (N_4260,N_69,N_843);
or U4261 (N_4261,N_1994,N_3821);
xor U4262 (N_4262,N_3035,N_318);
and U4263 (N_4263,N_3417,N_1191);
nand U4264 (N_4264,N_1351,N_2446);
or U4265 (N_4265,N_3931,N_2483);
or U4266 (N_4266,N_321,N_2792);
nor U4267 (N_4267,N_3414,N_315);
nand U4268 (N_4268,N_1173,N_176);
and U4269 (N_4269,N_1826,N_1006);
nor U4270 (N_4270,N_3726,N_3480);
nor U4271 (N_4271,N_3031,N_1861);
nand U4272 (N_4272,N_2866,N_3094);
or U4273 (N_4273,N_291,N_2750);
nor U4274 (N_4274,N_1263,N_2894);
or U4275 (N_4275,N_1375,N_610);
and U4276 (N_4276,N_585,N_2555);
and U4277 (N_4277,N_979,N_1470);
nor U4278 (N_4278,N_60,N_2928);
nor U4279 (N_4279,N_1267,N_224);
and U4280 (N_4280,N_339,N_1227);
or U4281 (N_4281,N_2363,N_1997);
nor U4282 (N_4282,N_1464,N_2971);
or U4283 (N_4283,N_3263,N_1858);
and U4284 (N_4284,N_1880,N_2059);
nor U4285 (N_4285,N_475,N_721);
nor U4286 (N_4286,N_2006,N_3545);
and U4287 (N_4287,N_2779,N_1875);
or U4288 (N_4288,N_438,N_409);
nor U4289 (N_4289,N_1639,N_811);
or U4290 (N_4290,N_3789,N_3281);
nor U4291 (N_4291,N_1047,N_3612);
and U4292 (N_4292,N_2980,N_3034);
and U4293 (N_4293,N_3079,N_2924);
nor U4294 (N_4294,N_1016,N_1769);
or U4295 (N_4295,N_2896,N_1975);
and U4296 (N_4296,N_3463,N_1183);
nand U4297 (N_4297,N_3835,N_2173);
nor U4298 (N_4298,N_3208,N_1102);
nor U4299 (N_4299,N_1025,N_1278);
nor U4300 (N_4300,N_694,N_3291);
nor U4301 (N_4301,N_369,N_22);
nand U4302 (N_4302,N_3353,N_3381);
nand U4303 (N_4303,N_1390,N_1149);
xnor U4304 (N_4304,N_3829,N_2979);
and U4305 (N_4305,N_2144,N_3148);
nand U4306 (N_4306,N_2686,N_1274);
nand U4307 (N_4307,N_462,N_2500);
and U4308 (N_4308,N_3027,N_933);
nand U4309 (N_4309,N_1553,N_2704);
or U4310 (N_4310,N_61,N_2115);
and U4311 (N_4311,N_924,N_2135);
nand U4312 (N_4312,N_1992,N_3819);
nand U4313 (N_4313,N_3329,N_3168);
or U4314 (N_4314,N_2608,N_3793);
and U4315 (N_4315,N_2561,N_1280);
nor U4316 (N_4316,N_1843,N_874);
nor U4317 (N_4317,N_3136,N_2224);
nand U4318 (N_4318,N_433,N_907);
nand U4319 (N_4319,N_2299,N_3434);
and U4320 (N_4320,N_2488,N_3274);
and U4321 (N_4321,N_1932,N_3877);
nor U4322 (N_4322,N_1082,N_660);
or U4323 (N_4323,N_1840,N_384);
xnor U4324 (N_4324,N_3008,N_1088);
or U4325 (N_4325,N_2479,N_1268);
nand U4326 (N_4326,N_78,N_2342);
nand U4327 (N_4327,N_109,N_1827);
nand U4328 (N_4328,N_2263,N_2855);
nand U4329 (N_4329,N_1783,N_1229);
nand U4330 (N_4330,N_162,N_2469);
xnor U4331 (N_4331,N_644,N_2474);
nor U4332 (N_4332,N_393,N_2986);
or U4333 (N_4333,N_3221,N_3994);
nand U4334 (N_4334,N_784,N_928);
nand U4335 (N_4335,N_1916,N_1957);
nand U4336 (N_4336,N_2906,N_1834);
nor U4337 (N_4337,N_2161,N_1528);
or U4338 (N_4338,N_541,N_1454);
nand U4339 (N_4339,N_3037,N_1027);
nor U4340 (N_4340,N_1857,N_2880);
or U4341 (N_4341,N_2613,N_862);
nor U4342 (N_4342,N_1002,N_1517);
or U4343 (N_4343,N_3044,N_2037);
or U4344 (N_4344,N_2298,N_965);
or U4345 (N_4345,N_104,N_257);
nor U4346 (N_4346,N_3714,N_3268);
or U4347 (N_4347,N_2507,N_2526);
and U4348 (N_4348,N_3209,N_1494);
nor U4349 (N_4349,N_3074,N_1257);
nor U4350 (N_4350,N_2015,N_876);
and U4351 (N_4351,N_1958,N_2915);
nor U4352 (N_4352,N_1175,N_212);
and U4353 (N_4353,N_1364,N_2431);
nand U4354 (N_4354,N_1451,N_1628);
nand U4355 (N_4355,N_2712,N_2152);
and U4356 (N_4356,N_3598,N_2753);
or U4357 (N_4357,N_779,N_2465);
or U4358 (N_4358,N_2615,N_1279);
or U4359 (N_4359,N_497,N_522);
and U4360 (N_4360,N_2741,N_3390);
nor U4361 (N_4361,N_736,N_1076);
nand U4362 (N_4362,N_3666,N_568);
or U4363 (N_4363,N_2955,N_851);
nand U4364 (N_4364,N_1136,N_1487);
nand U4365 (N_4365,N_1791,N_834);
nand U4366 (N_4366,N_3863,N_1923);
and U4367 (N_4367,N_1671,N_3862);
nor U4368 (N_4368,N_592,N_1947);
or U4369 (N_4369,N_187,N_3751);
nor U4370 (N_4370,N_337,N_2681);
and U4371 (N_4371,N_703,N_1655);
or U4372 (N_4372,N_1631,N_28);
nor U4373 (N_4373,N_181,N_3141);
nor U4374 (N_4374,N_1125,N_1795);
nor U4375 (N_4375,N_2133,N_1458);
nand U4376 (N_4376,N_820,N_3803);
nor U4377 (N_4377,N_2560,N_3117);
nor U4378 (N_4378,N_217,N_1281);
or U4379 (N_4379,N_3894,N_2751);
or U4380 (N_4380,N_1736,N_74);
or U4381 (N_4381,N_3708,N_103);
and U4382 (N_4382,N_714,N_1972);
nor U4383 (N_4383,N_2207,N_2245);
xor U4384 (N_4384,N_2977,N_2202);
or U4385 (N_4385,N_749,N_3093);
xnor U4386 (N_4386,N_2514,N_655);
nor U4387 (N_4387,N_2734,N_3483);
xor U4388 (N_4388,N_3126,N_3361);
nand U4389 (N_4389,N_894,N_3630);
and U4390 (N_4390,N_1591,N_2603);
or U4391 (N_4391,N_2111,N_389);
nor U4392 (N_4392,N_2344,N_685);
xnor U4393 (N_4393,N_1891,N_2244);
xor U4394 (N_4394,N_203,N_1297);
nand U4395 (N_4395,N_2864,N_1217);
nor U4396 (N_4396,N_1652,N_3661);
nor U4397 (N_4397,N_535,N_3954);
and U4398 (N_4398,N_939,N_3866);
or U4399 (N_4399,N_2028,N_2626);
and U4400 (N_4400,N_611,N_988);
and U4401 (N_4401,N_2511,N_3709);
xnor U4402 (N_4402,N_1273,N_156);
xnor U4403 (N_4403,N_2937,N_3199);
and U4404 (N_4404,N_1038,N_1674);
or U4405 (N_4405,N_2067,N_2339);
xor U4406 (N_4406,N_2197,N_676);
or U4407 (N_4407,N_3153,N_836);
and U4408 (N_4408,N_228,N_802);
and U4409 (N_4409,N_1512,N_882);
nor U4410 (N_4410,N_1805,N_1413);
nor U4411 (N_4411,N_413,N_1482);
nand U4412 (N_4412,N_1444,N_971);
nand U4413 (N_4413,N_142,N_3415);
nand U4414 (N_4414,N_1734,N_741);
and U4415 (N_4415,N_2951,N_3533);
and U4416 (N_4416,N_2576,N_3992);
nor U4417 (N_4417,N_1101,N_601);
nor U4418 (N_4418,N_1219,N_3753);
nand U4419 (N_4419,N_3888,N_1453);
or U4420 (N_4420,N_801,N_1699);
or U4421 (N_4421,N_500,N_83);
nand U4422 (N_4422,N_3875,N_1913);
nand U4423 (N_4423,N_3579,N_2571);
nand U4424 (N_4424,N_3949,N_252);
nor U4425 (N_4425,N_1684,N_35);
and U4426 (N_4426,N_1032,N_125);
nor U4427 (N_4427,N_950,N_3944);
or U4428 (N_4428,N_3103,N_1109);
and U4429 (N_4429,N_543,N_79);
nor U4430 (N_4430,N_1392,N_246);
nor U4431 (N_4431,N_3643,N_1965);
nor U4432 (N_4432,N_3014,N_3563);
xor U4433 (N_4433,N_2307,N_3955);
xnor U4434 (N_4434,N_3083,N_3748);
and U4435 (N_4435,N_3382,N_177);
nand U4436 (N_4436,N_1866,N_3270);
and U4437 (N_4437,N_328,N_960);
or U4438 (N_4438,N_2552,N_1171);
nor U4439 (N_4439,N_806,N_1354);
nor U4440 (N_4440,N_2941,N_2203);
xor U4441 (N_4441,N_1414,N_3520);
or U4442 (N_4442,N_3445,N_930);
or U4443 (N_4443,N_1847,N_412);
or U4444 (N_4444,N_459,N_1690);
nand U4445 (N_4445,N_548,N_1130);
xor U4446 (N_4446,N_3791,N_2482);
nor U4447 (N_4447,N_3745,N_1952);
nand U4448 (N_4448,N_3022,N_537);
xnor U4449 (N_4449,N_2337,N_2089);
and U4450 (N_4450,N_3660,N_2171);
nand U4451 (N_4451,N_1221,N_1260);
and U4452 (N_4452,N_1134,N_3278);
nor U4453 (N_4453,N_680,N_880);
nand U4454 (N_4454,N_2326,N_3868);
nand U4455 (N_4455,N_921,N_3947);
and U4456 (N_4456,N_3239,N_577);
nand U4457 (N_4457,N_2960,N_2009);
and U4458 (N_4458,N_2287,N_2021);
and U4459 (N_4459,N_3589,N_838);
nor U4460 (N_4460,N_3639,N_1308);
nand U4461 (N_4461,N_1835,N_1689);
and U4462 (N_4462,N_3658,N_3007);
and U4463 (N_4463,N_3592,N_1956);
xor U4464 (N_4464,N_1234,N_1064);
nand U4465 (N_4465,N_27,N_3179);
nand U4466 (N_4466,N_386,N_283);
xor U4467 (N_4467,N_3088,N_3655);
and U4468 (N_4468,N_2595,N_2486);
nor U4469 (N_4469,N_3932,N_2417);
or U4470 (N_4470,N_2853,N_701);
nor U4471 (N_4471,N_2565,N_356);
nor U4472 (N_4472,N_3432,N_762);
nor U4473 (N_4473,N_1304,N_3542);
nand U4474 (N_4474,N_3770,N_3902);
or U4475 (N_4475,N_165,N_1526);
xor U4476 (N_4476,N_1704,N_502);
and U4477 (N_4477,N_1419,N_3403);
nor U4478 (N_4478,N_2849,N_2470);
nor U4479 (N_4479,N_3775,N_1936);
nor U4480 (N_4480,N_863,N_2978);
nand U4481 (N_4481,N_3548,N_2525);
nand U4482 (N_4482,N_1651,N_3597);
xnor U4483 (N_4483,N_3401,N_2536);
nor U4484 (N_4484,N_776,N_2476);
or U4485 (N_4485,N_171,N_2257);
or U4486 (N_4486,N_2098,N_1409);
nand U4487 (N_4487,N_3880,N_674);
nor U4488 (N_4488,N_2534,N_1166);
nand U4489 (N_4489,N_3855,N_3211);
nor U4490 (N_4490,N_1818,N_814);
and U4491 (N_4491,N_2548,N_2748);
or U4492 (N_4492,N_373,N_526);
or U4493 (N_4493,N_1532,N_1708);
nor U4494 (N_4494,N_1442,N_596);
and U4495 (N_4495,N_2940,N_72);
nor U4496 (N_4496,N_3869,N_2461);
nand U4497 (N_4497,N_1204,N_1995);
nor U4498 (N_4498,N_1794,N_1718);
nand U4499 (N_4499,N_2578,N_3749);
or U4500 (N_4500,N_868,N_2523);
or U4501 (N_4501,N_3205,N_1112);
or U4502 (N_4502,N_1584,N_2400);
nand U4503 (N_4503,N_2093,N_1317);
nand U4504 (N_4504,N_3781,N_2041);
nor U4505 (N_4505,N_3514,N_1918);
nand U4506 (N_4506,N_1474,N_1810);
and U4507 (N_4507,N_3540,N_1226);
xor U4508 (N_4508,N_679,N_2104);
xor U4509 (N_4509,N_2967,N_1446);
or U4510 (N_4510,N_3076,N_2881);
and U4511 (N_4511,N_2532,N_231);
and U4512 (N_4512,N_1828,N_2107);
nand U4513 (N_4513,N_1524,N_2070);
nand U4514 (N_4514,N_489,N_2137);
nor U4515 (N_4515,N_739,N_968);
and U4516 (N_4516,N_1151,N_614);
or U4517 (N_4517,N_2053,N_129);
nand U4518 (N_4518,N_3269,N_2990);
nor U4519 (N_4519,N_421,N_3506);
or U4520 (N_4520,N_1197,N_1199);
or U4521 (N_4521,N_309,N_1156);
nor U4522 (N_4522,N_123,N_366);
and U4523 (N_4523,N_3647,N_1888);
or U4524 (N_4524,N_3922,N_2075);
and U4525 (N_4525,N_1300,N_1819);
nand U4526 (N_4526,N_1569,N_273);
xnor U4527 (N_4527,N_936,N_2311);
nor U4528 (N_4528,N_1894,N_1643);
nor U4529 (N_4529,N_2722,N_1299);
nand U4530 (N_4530,N_1626,N_2789);
nand U4531 (N_4531,N_558,N_2074);
xnor U4532 (N_4532,N_3999,N_2856);
or U4533 (N_4533,N_2892,N_670);
and U4534 (N_4534,N_1518,N_3554);
nor U4535 (N_4535,N_3192,N_1230);
and U4536 (N_4536,N_1730,N_1346);
and U4537 (N_4537,N_2587,N_3285);
nor U4538 (N_4538,N_355,N_3711);
and U4539 (N_4539,N_2766,N_1439);
nand U4540 (N_4540,N_2189,N_3108);
nand U4541 (N_4541,N_698,N_3259);
nand U4542 (N_4542,N_603,N_3082);
and U4543 (N_4543,N_3537,N_1988);
or U4544 (N_4544,N_625,N_1190);
nand U4545 (N_4545,N_1850,N_1945);
nor U4546 (N_4546,N_3487,N_3893);
and U4547 (N_4547,N_2964,N_1648);
nor U4548 (N_4548,N_3562,N_2220);
nor U4549 (N_4549,N_3912,N_2886);
or U4550 (N_4550,N_288,N_3825);
xnor U4551 (N_4551,N_951,N_234);
or U4552 (N_4552,N_2250,N_2035);
nor U4553 (N_4553,N_553,N_1558);
nor U4554 (N_4554,N_3713,N_3481);
nor U4555 (N_4555,N_1434,N_1138);
nor U4556 (N_4556,N_3150,N_1613);
and U4557 (N_4557,N_3242,N_1187);
nor U4558 (N_4558,N_2249,N_1396);
nand U4559 (N_4559,N_3092,N_691);
and U4560 (N_4560,N_1259,N_390);
and U4561 (N_4561,N_2081,N_3060);
and U4562 (N_4562,N_3134,N_1989);
or U4563 (N_4563,N_3942,N_530);
nand U4564 (N_4564,N_3983,N_172);
nand U4565 (N_4565,N_2063,N_3561);
or U4566 (N_4566,N_1307,N_1157);
nor U4567 (N_4567,N_3885,N_1585);
or U4568 (N_4568,N_3372,N_1960);
xnor U4569 (N_4569,N_1209,N_2570);
nand U4570 (N_4570,N_3634,N_738);
and U4571 (N_4571,N_766,N_333);
or U4572 (N_4572,N_551,N_2073);
and U4573 (N_4573,N_199,N_717);
nand U4574 (N_4574,N_3915,N_491);
nor U4575 (N_4575,N_352,N_1324);
nor U4576 (N_4576,N_3951,N_919);
or U4577 (N_4577,N_899,N_2775);
nand U4578 (N_4578,N_3526,N_3958);
xnor U4579 (N_4579,N_3507,N_1944);
nor U4580 (N_4580,N_2275,N_41);
nor U4581 (N_4581,N_2423,N_1374);
and U4582 (N_4582,N_3025,N_63);
nand U4583 (N_4583,N_235,N_2455);
nor U4584 (N_4584,N_3431,N_3045);
nor U4585 (N_4585,N_3305,N_3373);
nor U4586 (N_4586,N_3913,N_841);
nor U4587 (N_4587,N_2281,N_1491);
nor U4588 (N_4588,N_2559,N_3890);
or U4589 (N_4589,N_2651,N_2769);
nand U4590 (N_4590,N_3096,N_1384);
nor U4591 (N_4591,N_2087,N_3937);
nand U4592 (N_4592,N_994,N_1401);
nor U4593 (N_4593,N_320,N_3679);
or U4594 (N_4594,N_1979,N_730);
xor U4595 (N_4595,N_2504,N_2697);
nor U4596 (N_4596,N_2736,N_3410);
nand U4597 (N_4597,N_3347,N_1552);
and U4598 (N_4598,N_56,N_2424);
nand U4599 (N_4599,N_3413,N_2562);
and U4600 (N_4600,N_3809,N_3491);
nand U4601 (N_4601,N_842,N_3498);
and U4602 (N_4602,N_1499,N_3154);
and U4603 (N_4603,N_1431,N_1029);
xnor U4604 (N_4604,N_3594,N_2688);
or U4605 (N_4605,N_2922,N_1438);
and U4606 (N_4606,N_3360,N_1367);
xor U4607 (N_4607,N_326,N_3620);
xnor U4608 (N_4608,N_3002,N_2255);
or U4609 (N_4609,N_357,N_1940);
nor U4610 (N_4610,N_1202,N_367);
and U4611 (N_4611,N_2014,N_1666);
nand U4612 (N_4612,N_756,N_1614);
nor U4613 (N_4613,N_2215,N_3217);
or U4614 (N_4614,N_3707,N_334);
nor U4615 (N_4615,N_3290,N_2412);
nand U4616 (N_4616,N_2933,N_3455);
and U4617 (N_4617,N_138,N_2974);
nor U4618 (N_4618,N_914,N_2791);
nor U4619 (N_4619,N_1170,N_3881);
and U4620 (N_4620,N_651,N_3457);
nor U4621 (N_4621,N_702,N_3804);
or U4622 (N_4622,N_71,N_3544);
xnor U4623 (N_4623,N_2592,N_615);
and U4624 (N_4624,N_1195,N_2090);
nand U4625 (N_4625,N_1249,N_3964);
or U4626 (N_4626,N_1243,N_2314);
nor U4627 (N_4627,N_445,N_14);
nor U4628 (N_4628,N_1776,N_3387);
xnor U4629 (N_4629,N_2017,N_1087);
xor U4630 (N_4630,N_3176,N_883);
nand U4631 (N_4631,N_313,N_1050);
xnor U4632 (N_4632,N_3249,N_1186);
nor U4633 (N_4633,N_3020,N_1286);
or U4634 (N_4634,N_419,N_2016);
nand U4635 (N_4635,N_3182,N_877);
nor U4636 (N_4636,N_2404,N_2372);
nor U4637 (N_4637,N_2900,N_3112);
and U4638 (N_4638,N_428,N_2332);
or U4639 (N_4639,N_207,N_2108);
nand U4640 (N_4640,N_2044,N_3446);
and U4641 (N_4641,N_3078,N_816);
or U4642 (N_4642,N_2306,N_276);
nand U4643 (N_4643,N_2349,N_1637);
nand U4644 (N_4644,N_1803,N_351);
nor U4645 (N_4645,N_3870,N_3696);
or U4646 (N_4646,N_2917,N_3160);
or U4647 (N_4647,N_628,N_2442);
nand U4648 (N_4648,N_2887,N_3760);
nor U4649 (N_4649,N_76,N_2718);
nor U4650 (N_4650,N_740,N_3423);
and U4651 (N_4651,N_2062,N_1348);
nor U4652 (N_4652,N_38,N_3566);
or U4653 (N_4653,N_2335,N_3019);
or U4654 (N_4654,N_461,N_3941);
or U4655 (N_4655,N_897,N_2374);
nor U4656 (N_4656,N_529,N_2247);
and U4657 (N_4657,N_1040,N_1424);
or U4658 (N_4658,N_3584,N_1020);
xor U4659 (N_4659,N_2328,N_1382);
nor U4660 (N_4660,N_3929,N_3681);
or U4661 (N_4661,N_1098,N_975);
xor U4662 (N_4662,N_3940,N_761);
or U4663 (N_4663,N_1756,N_448);
nand U4664 (N_4664,N_3527,N_706);
xnor U4665 (N_4665,N_1340,N_1181);
and U4666 (N_4666,N_1679,N_2158);
or U4667 (N_4667,N_388,N_2839);
and U4668 (N_4668,N_1058,N_1747);
nor U4669 (N_4669,N_2061,N_2591);
nand U4670 (N_4670,N_2395,N_3933);
and U4671 (N_4671,N_2585,N_716);
or U4672 (N_4672,N_3739,N_3604);
or U4673 (N_4673,N_3493,N_1400);
and U4674 (N_4674,N_2176,N_2795);
nand U4675 (N_4675,N_1562,N_2654);
nor U4676 (N_4676,N_2577,N_3519);
and U4677 (N_4677,N_866,N_2003);
nand U4678 (N_4678,N_1228,N_2487);
and U4679 (N_4679,N_2499,N_3788);
and U4680 (N_4680,N_1327,N_3472);
nand U4681 (N_4681,N_1608,N_116);
and U4682 (N_4682,N_3722,N_3538);
and U4683 (N_4683,N_2226,N_3474);
nand U4684 (N_4684,N_909,N_67);
and U4685 (N_4685,N_2804,N_2586);
nand U4686 (N_4686,N_211,N_343);
or U4687 (N_4687,N_3229,N_3436);
and U4688 (N_4688,N_382,N_993);
nand U4689 (N_4689,N_822,N_3861);
xnor U4690 (N_4690,N_1978,N_97);
nand U4691 (N_4691,N_2623,N_1853);
and U4692 (N_4692,N_2865,N_3422);
or U4693 (N_4693,N_194,N_2389);
or U4694 (N_4694,N_2401,N_3222);
or U4695 (N_4695,N_1969,N_1632);
nand U4696 (N_4696,N_2828,N_2222);
xor U4697 (N_4697,N_1005,N_330);
or U4698 (N_4698,N_295,N_1200);
xnor U4699 (N_4699,N_2944,N_2538);
nor U4700 (N_4700,N_684,N_2381);
and U4701 (N_4701,N_1877,N_2744);
and U4702 (N_4702,N_303,N_1807);
or U4703 (N_4703,N_3120,N_3663);
and U4704 (N_4704,N_105,N_2821);
and U4705 (N_4705,N_3204,N_2634);
nand U4706 (N_4706,N_1201,N_967);
or U4707 (N_4707,N_2811,N_2502);
nor U4708 (N_4708,N_3638,N_152);
and U4709 (N_4709,N_2292,N_2958);
or U4710 (N_4710,N_1692,N_3732);
nand U4711 (N_4711,N_891,N_3212);
nor U4712 (N_4712,N_3948,N_608);
xor U4713 (N_4713,N_2975,N_3938);
and U4714 (N_4714,N_3840,N_3974);
or U4715 (N_4715,N_3656,N_3185);
nor U4716 (N_4716,N_885,N_117);
nor U4717 (N_4717,N_3464,N_3617);
nand U4718 (N_4718,N_3989,N_98);
xor U4719 (N_4719,N_2494,N_3755);
nor U4720 (N_4720,N_3366,N_2758);
and U4721 (N_4721,N_2945,N_322);
nor U4722 (N_4722,N_141,N_467);
nor U4723 (N_4723,N_2812,N_3201);
and U4724 (N_4724,N_2223,N_985);
and U4725 (N_4725,N_3032,N_255);
nor U4726 (N_4726,N_3023,N_1077);
nor U4727 (N_4727,N_2466,N_3476);
nand U4728 (N_4728,N_3024,N_747);
nand U4729 (N_4729,N_375,N_2347);
nor U4730 (N_4730,N_2813,N_2918);
or U4731 (N_4731,N_2375,N_3799);
nand U4732 (N_4732,N_931,N_1998);
nand U4733 (N_4733,N_3262,N_2365);
nand U4734 (N_4734,N_2781,N_195);
nand U4735 (N_4735,N_3657,N_1019);
nand U4736 (N_4736,N_1009,N_2020);
or U4737 (N_4737,N_632,N_3536);
or U4738 (N_4738,N_3501,N_3810);
nand U4739 (N_4739,N_618,N_1824);
nand U4740 (N_4740,N_3137,N_2759);
nor U4741 (N_4741,N_1500,N_2696);
nor U4742 (N_4742,N_752,N_414);
xor U4743 (N_4743,N_1700,N_208);
and U4744 (N_4744,N_2999,N_3671);
xor U4745 (N_4745,N_1845,N_2034);
nor U4746 (N_4746,N_2359,N_3827);
and U4747 (N_4747,N_2475,N_1440);
and U4748 (N_4748,N_2725,N_1865);
nor U4749 (N_4749,N_755,N_3695);
nor U4750 (N_4750,N_1481,N_287);
nor U4751 (N_4751,N_2777,N_1742);
or U4752 (N_4752,N_3,N_3129);
xor U4753 (N_4753,N_2700,N_3859);
or U4754 (N_4754,N_672,N_3499);
nand U4755 (N_4755,N_2495,N_657);
nand U4756 (N_4756,N_576,N_986);
or U4757 (N_4757,N_128,N_1922);
nor U4758 (N_4758,N_892,N_1143);
and U4759 (N_4759,N_1764,N_3266);
and U4760 (N_4760,N_602,N_1508);
nor U4761 (N_4761,N_589,N_1092);
nor U4762 (N_4762,N_2183,N_3190);
xnor U4763 (N_4763,N_3857,N_1711);
nand U4764 (N_4764,N_2632,N_1389);
or U4765 (N_4765,N_785,N_451);
nor U4766 (N_4766,N_1574,N_3555);
or U4767 (N_4767,N_1695,N_153);
nand U4768 (N_4768,N_3143,N_884);
or U4769 (N_4769,N_2735,N_115);
and U4770 (N_4770,N_3596,N_1640);
or U4771 (N_4771,N_2656,N_3602);
nand U4772 (N_4772,N_2290,N_2065);
and U4773 (N_4773,N_2132,N_2246);
xnor U4774 (N_4774,N_2588,N_2180);
or U4775 (N_4775,N_1344,N_1677);
nor U4776 (N_4776,N_2295,N_299);
nand U4777 (N_4777,N_1017,N_1593);
and U4778 (N_4778,N_1036,N_411);
and U4779 (N_4779,N_3528,N_2206);
or U4780 (N_4780,N_430,N_1310);
nand U4781 (N_4781,N_3330,N_2841);
or U4782 (N_4782,N_3105,N_1724);
and U4783 (N_4783,N_1768,N_87);
and U4784 (N_4784,N_536,N_1106);
and U4785 (N_4785,N_715,N_3332);
xor U4786 (N_4786,N_2126,N_121);
or U4787 (N_4787,N_1337,N_2039);
nand U4788 (N_4788,N_2754,N_1176);
nor U4789 (N_4789,N_3769,N_953);
nor U4790 (N_4790,N_794,N_3685);
or U4791 (N_4791,N_3971,N_1964);
or U4792 (N_4792,N_1545,N_2278);
xor U4793 (N_4793,N_345,N_9);
or U4794 (N_4794,N_922,N_1529);
nor U4795 (N_4795,N_641,N_3288);
nor U4796 (N_4796,N_1361,N_2622);
or U4797 (N_4797,N_2545,N_2195);
and U4798 (N_4798,N_3041,N_1970);
or U4799 (N_4799,N_946,N_2618);
and U4800 (N_4800,N_3485,N_1493);
nand U4801 (N_4801,N_3340,N_1496);
nand U4802 (N_4802,N_2513,N_1447);
or U4803 (N_4803,N_3240,N_722);
nor U4804 (N_4804,N_2052,N_3174);
nand U4805 (N_4805,N_925,N_2405);
nor U4806 (N_4806,N_1429,N_861);
nand U4807 (N_4807,N_1869,N_3337);
nor U4808 (N_4808,N_760,N_1985);
and U4809 (N_4809,N_1588,N_2630);
nor U4810 (N_4810,N_1428,N_1550);
nor U4811 (N_4811,N_2419,N_249);
nand U4812 (N_4812,N_3375,N_3790);
or U4813 (N_4813,N_1515,N_2205);
and U4814 (N_4814,N_1046,N_3962);
and U4815 (N_4815,N_307,N_423);
nand U4816 (N_4816,N_2129,N_3320);
or U4817 (N_4817,N_590,N_1802);
nand U4818 (N_4818,N_3038,N_3648);
nand U4819 (N_4819,N_1462,N_3767);
and U4820 (N_4820,N_3420,N_3659);
and U4821 (N_4821,N_2172,N_612);
nand U4822 (N_4822,N_135,N_1852);
and U4823 (N_4823,N_1455,N_1086);
nor U4824 (N_4824,N_3072,N_483);
nand U4825 (N_4825,N_3672,N_1667);
and U4826 (N_4826,N_3574,N_540);
nand U4827 (N_4827,N_1037,N_3826);
or U4828 (N_4828,N_633,N_3924);
and U4829 (N_4829,N_1293,N_3429);
nor U4830 (N_4830,N_196,N_2201);
or U4831 (N_4831,N_190,N_1312);
xor U4832 (N_4832,N_350,N_494);
nor U4833 (N_4833,N_1285,N_2251);
nand U4834 (N_4834,N_1232,N_2248);
and U4835 (N_4835,N_2019,N_3100);
nor U4836 (N_4836,N_397,N_102);
nand U4837 (N_4837,N_2316,N_2179);
nand U4838 (N_4838,N_604,N_3818);
and U4839 (N_4839,N_1519,N_917);
nand U4840 (N_4840,N_2790,N_2054);
nand U4841 (N_4841,N_1238,N_1426);
xor U4842 (N_4842,N_1437,N_3003);
nor U4843 (N_4843,N_65,N_3513);
nand U4844 (N_4844,N_353,N_3066);
or U4845 (N_4845,N_1152,N_2503);
and U4846 (N_4846,N_2312,N_2490);
and U4847 (N_4847,N_1241,N_439);
nand U4848 (N_4848,N_1980,N_1782);
nand U4849 (N_4849,N_112,N_759);
xor U4850 (N_4850,N_468,N_754);
nor U4851 (N_4851,N_469,N_2353);
nand U4852 (N_4852,N_85,N_3349);
or U4853 (N_4853,N_2168,N_101);
or U4854 (N_4854,N_3688,N_1598);
nor U4855 (N_4855,N_110,N_2443);
and U4856 (N_4856,N_2141,N_3419);
nor U4857 (N_4857,N_54,N_2048);
nand U4858 (N_4858,N_1902,N_170);
and U4859 (N_4859,N_2027,N_460);
nor U4860 (N_4860,N_133,N_3687);
nor U4861 (N_4861,N_464,N_2574);
or U4862 (N_4862,N_2324,N_1905);
nor U4863 (N_4863,N_2134,N_732);
nand U4864 (N_4864,N_947,N_533);
or U4865 (N_4865,N_495,N_3652);
and U4866 (N_4866,N_645,N_2810);
nor U4867 (N_4867,N_3059,N_1903);
and U4868 (N_4868,N_201,N_847);
nor U4869 (N_4869,N_2350,N_2376);
or U4870 (N_4870,N_887,N_3055);
or U4871 (N_4871,N_2551,N_3384);
nand U4872 (N_4872,N_1410,N_2648);
nand U4873 (N_4873,N_3535,N_2371);
nand U4874 (N_4874,N_3131,N_2649);
or U4875 (N_4875,N_1811,N_2154);
nand U4876 (N_4876,N_2976,N_3995);
nor U4877 (N_4877,N_1305,N_1416);
or U4878 (N_4878,N_839,N_1971);
nor U4879 (N_4879,N_301,N_3435);
nor U4880 (N_4880,N_3593,N_1514);
or U4881 (N_4881,N_2757,N_570);
and U4882 (N_4882,N_3251,N_247);
nand U4883 (N_4883,N_2106,N_1694);
or U4884 (N_4884,N_2852,N_1977);
nand U4885 (N_4885,N_3460,N_158);
or U4886 (N_4886,N_3233,N_1313);
or U4887 (N_4887,N_465,N_2091);
nor U4888 (N_4888,N_2518,N_150);
nor U4889 (N_4889,N_2491,N_2993);
and U4890 (N_4890,N_789,N_812);
and U4891 (N_4891,N_2535,N_580);
nand U4892 (N_4892,N_2282,N_945);
or U4893 (N_4893,N_88,N_970);
and U4894 (N_4894,N_1258,N_1261);
nor U4895 (N_4895,N_623,N_482);
nor U4896 (N_4896,N_2863,N_1345);
and U4897 (N_4897,N_3939,N_2313);
nor U4898 (N_4898,N_1664,N_2800);
and U4899 (N_4899,N_3095,N_3430);
nor U4900 (N_4900,N_1713,N_2296);
nand U4901 (N_4901,N_3834,N_3705);
nand U4902 (N_4902,N_1654,N_2261);
nand U4903 (N_4903,N_3416,N_2149);
nand U4904 (N_4904,N_62,N_1895);
or U4905 (N_4905,N_1333,N_765);
or U4906 (N_4906,N_2320,N_561);
or U4907 (N_4907,N_2539,N_1938);
nor U4908 (N_4908,N_2910,N_2309);
nor U4909 (N_4909,N_3570,N_1625);
nor U4910 (N_4910,N_3467,N_3909);
nor U4911 (N_4911,N_1530,N_3468);
nor U4912 (N_4912,N_731,N_2032);
or U4913 (N_4913,N_1319,N_3550);
nor U4914 (N_4914,N_1043,N_385);
and U4915 (N_4915,N_594,N_2952);
xnor U4916 (N_4916,N_2123,N_392);
or U4917 (N_4917,N_1459,N_1996);
nor U4918 (N_4918,N_3000,N_3316);
nor U4919 (N_4919,N_3646,N_3896);
nor U4920 (N_4920,N_2954,N_3345);
xor U4921 (N_4921,N_3689,N_1288);
and U4922 (N_4922,N_2959,N_1119);
nor U4923 (N_4923,N_626,N_3737);
and U4924 (N_4924,N_3346,N_1255);
or U4925 (N_4925,N_3412,N_2929);
nand U4926 (N_4926,N_1656,N_3049);
nor U4927 (N_4927,N_2833,N_1115);
or U4928 (N_4928,N_1172,N_2235);
or U4929 (N_4929,N_1642,N_1342);
and U4930 (N_4930,N_3186,N_2981);
or U4931 (N_4931,N_3081,N_3569);
xnor U4932 (N_4932,N_2598,N_2155);
nor U4933 (N_4933,N_1071,N_1488);
nand U4934 (N_4934,N_2653,N_2399);
nand U4935 (N_4935,N_2860,N_991);
or U4936 (N_4936,N_2912,N_2283);
and U4937 (N_4937,N_867,N_1417);
and U4938 (N_4938,N_3371,N_1490);
nand U4939 (N_4939,N_2666,N_2047);
xor U4940 (N_4940,N_1180,N_807);
nor U4941 (N_4941,N_1177,N_163);
nor U4942 (N_4942,N_3004,N_709);
nor U4943 (N_4943,N_362,N_3532);
and U4944 (N_4944,N_2450,N_1887);
nor U4945 (N_4945,N_504,N_572);
and U4946 (N_4946,N_3547,N_1207);
nand U4947 (N_4947,N_2665,N_380);
and U4948 (N_4948,N_1218,N_1766);
nor U4949 (N_4949,N_2867,N_1189);
and U4950 (N_4950,N_1815,N_1531);
or U4951 (N_4951,N_1658,N_1253);
or U4952 (N_4952,N_2723,N_1460);
nand U4953 (N_4953,N_2018,N_2684);
xor U4954 (N_4954,N_2816,N_2266);
nand U4955 (N_4955,N_166,N_3181);
and U4956 (N_4956,N_1302,N_3171);
nor U4957 (N_4957,N_517,N_1254);
nand U4958 (N_4958,N_2293,N_3189);
nor U4959 (N_4959,N_271,N_53);
nor U4960 (N_4960,N_2481,N_869);
nand U4961 (N_4961,N_2270,N_1729);
or U4962 (N_4962,N_118,N_1318);
or U4963 (N_4963,N_3149,N_3057);
and U4964 (N_4964,N_16,N_368);
or U4965 (N_4965,N_2453,N_1194);
nor U4966 (N_4966,N_2420,N_3703);
nand U4967 (N_4967,N_3047,N_248);
and U4968 (N_4968,N_977,N_1926);
nor U4969 (N_4969,N_3231,N_1247);
nand U4970 (N_4970,N_3783,N_1925);
or U4971 (N_4971,N_2773,N_3828);
nor U4972 (N_4972,N_1069,N_3797);
and U4973 (N_4973,N_1266,N_3452);
nand U4974 (N_4974,N_1406,N_3606);
nand U4975 (N_4975,N_2768,N_511);
xnor U4976 (N_4976,N_1296,N_844);
nor U4977 (N_4977,N_1322,N_1867);
and U4978 (N_4978,N_1485,N_2635);
or U4979 (N_4979,N_2724,N_3500);
or U4980 (N_4980,N_3173,N_1145);
xor U4981 (N_4981,N_3121,N_2857);
nor U4982 (N_4982,N_1430,N_3080);
nand U4983 (N_4983,N_3918,N_3742);
or U4984 (N_4984,N_2042,N_2064);
nand U4985 (N_4985,N_3697,N_17);
or U4986 (N_4986,N_1042,N_219);
nand U4987 (N_4987,N_2984,N_2024);
nor U4988 (N_4988,N_1685,N_1178);
and U4989 (N_4989,N_1505,N_267);
or U4990 (N_4990,N_864,N_2767);
or U4991 (N_4991,N_3359,N_2835);
and U4992 (N_4992,N_134,N_1443);
and U4993 (N_4993,N_962,N_2785);
and U4994 (N_4994,N_311,N_1339);
and U4995 (N_4995,N_2080,N_3608);
nand U4996 (N_4996,N_2038,N_1966);
nor U4997 (N_4997,N_2788,N_3441);
nand U4998 (N_4998,N_3163,N_481);
nand U4999 (N_4999,N_3985,N_3086);
nor U5000 (N_5000,N_3601,N_2966);
or U5001 (N_5001,N_3930,N_2672);
xnor U5002 (N_5002,N_3089,N_3756);
nor U5003 (N_5003,N_2346,N_2690);
nand U5004 (N_5004,N_1720,N_3605);
nand U5005 (N_5005,N_3010,N_748);
xnor U5006 (N_5006,N_805,N_1235);
or U5007 (N_5007,N_1726,N_1456);
and U5008 (N_5008,N_1618,N_888);
nor U5009 (N_5009,N_3454,N_3591);
and U5010 (N_5010,N_2471,N_1551);
nand U5011 (N_5011,N_3264,N_1486);
or U5012 (N_5012,N_3062,N_1105);
xnor U5013 (N_5013,N_2701,N_2644);
nand U5014 (N_5014,N_25,N_1330);
nor U5015 (N_5015,N_2473,N_225);
nor U5016 (N_5016,N_3794,N_1301);
nand U5017 (N_5017,N_2498,N_2165);
or U5018 (N_5018,N_2413,N_1159);
nand U5019 (N_5019,N_2802,N_2891);
and U5020 (N_5020,N_1884,N_827);
or U5021 (N_5021,N_1898,N_1252);
nor U5022 (N_5022,N_1797,N_2557);
nand U5023 (N_5023,N_1882,N_15);
or U5024 (N_5024,N_3124,N_132);
nor U5025 (N_5025,N_3177,N_2364);
or U5026 (N_5026,N_1250,N_3629);
or U5027 (N_5027,N_1703,N_3625);
and U5028 (N_5028,N_2143,N_1737);
or U5029 (N_5029,N_699,N_1825);
nand U5030 (N_5030,N_2872,N_3752);
and U5031 (N_5031,N_1934,N_524);
nand U5032 (N_5032,N_2695,N_2660);
nand U5033 (N_5033,N_1697,N_2991);
or U5034 (N_5034,N_3132,N_1193);
or U5035 (N_5035,N_3050,N_2604);
nand U5036 (N_5036,N_2782,N_582);
nor U5037 (N_5037,N_3017,N_3700);
or U5038 (N_5038,N_3286,N_220);
or U5039 (N_5039,N_3056,N_1179);
nor U5040 (N_5040,N_893,N_2071);
and U5041 (N_5041,N_697,N_332);
or U5042 (N_5042,N_21,N_1244);
and U5043 (N_5043,N_189,N_1775);
or U5044 (N_5044,N_2898,N_2969);
xnor U5045 (N_5045,N_1323,N_2527);
nand U5046 (N_5046,N_2830,N_263);
nand U5047 (N_5047,N_1316,N_2178);
or U5048 (N_5048,N_31,N_1185);
and U5049 (N_5049,N_3115,N_2713);
nand U5050 (N_5050,N_1117,N_2406);
and U5051 (N_5051,N_2433,N_3351);
nand U5052 (N_5052,N_1723,N_89);
nor U5053 (N_5053,N_484,N_1627);
nor U5054 (N_5054,N_2264,N_2638);
nor U5055 (N_5055,N_2580,N_3257);
and U5056 (N_5056,N_3284,N_3734);
nand U5057 (N_5057,N_3986,N_929);
and U5058 (N_5058,N_1623,N_2428);
and U5059 (N_5059,N_3187,N_270);
nor U5060 (N_5060,N_2601,N_1332);
nand U5061 (N_5061,N_938,N_2702);
nand U5062 (N_5062,N_1793,N_3459);
nand U5063 (N_5063,N_2531,N_1868);
xor U5064 (N_5064,N_3334,N_3295);
nor U5065 (N_5065,N_2728,N_2807);
xnor U5066 (N_5066,N_3001,N_1291);
nor U5067 (N_5067,N_3391,N_365);
and U5068 (N_5068,N_2920,N_2095);
nor U5069 (N_5069,N_3183,N_896);
nand U5070 (N_5070,N_2094,N_298);
nor U5071 (N_5071,N_508,N_833);
or U5072 (N_5072,N_1208,N_1993);
nand U5073 (N_5073,N_3743,N_3787);
and U5074 (N_5074,N_2068,N_780);
nor U5075 (N_5075,N_2809,N_2243);
or U5076 (N_5076,N_1921,N_3097);
and U5077 (N_5077,N_1800,N_1676);
and U5078 (N_5078,N_1904,N_3479);
nand U5079 (N_5079,N_3307,N_3128);
and U5080 (N_5080,N_3935,N_943);
and U5081 (N_5081,N_2939,N_1981);
nor U5082 (N_5082,N_3645,N_588);
xor U5083 (N_5083,N_3497,N_3968);
nor U5084 (N_5084,N_3733,N_238);
nand U5085 (N_5085,N_3256,N_1830);
xnor U5086 (N_5086,N_2040,N_1931);
and U5087 (N_5087,N_1660,N_3358);
or U5088 (N_5088,N_29,N_2780);
nand U5089 (N_5089,N_3478,N_1535);
nor U5090 (N_5090,N_2719,N_1816);
nand U5091 (N_5091,N_3824,N_209);
nor U5092 (N_5092,N_586,N_3443);
nor U5093 (N_5093,N_30,N_401);
and U5094 (N_5094,N_300,N_1889);
nand U5095 (N_5095,N_2200,N_3772);
or U5096 (N_5096,N_2738,N_205);
or U5097 (N_5097,N_2670,N_1355);
and U5098 (N_5098,N_1140,N_2418);
xnor U5099 (N_5099,N_635,N_450);
nand U5100 (N_5100,N_2218,N_2459);
nand U5101 (N_5101,N_1147,N_1999);
and U5102 (N_5102,N_2429,N_3792);
and U5103 (N_5103,N_3175,N_2646);
xnor U5104 (N_5104,N_1483,N_3426);
or U5105 (N_5105,N_94,N_2012);
nand U5106 (N_5106,N_3823,N_3310);
and U5107 (N_5107,N_3469,N_1743);
and U5108 (N_5108,N_3139,N_179);
and U5109 (N_5109,N_42,N_2546);
nand U5110 (N_5110,N_2213,N_2241);
nand U5111 (N_5111,N_2564,N_1554);
or U5112 (N_5112,N_2441,N_1833);
xnor U5113 (N_5113,N_3747,N_2671);
and U5114 (N_5114,N_1044,N_2756);
xor U5115 (N_5115,N_1003,N_3618);
nand U5116 (N_5116,N_1377,N_186);
and U5117 (N_5117,N_2166,N_3766);
and U5118 (N_5118,N_2680,N_3151);
nand U5119 (N_5119,N_788,N_3357);
and U5120 (N_5120,N_1893,N_501);
nor U5121 (N_5121,N_2033,N_403);
nand U5122 (N_5122,N_1205,N_2022);
nand U5123 (N_5123,N_713,N_3223);
xnor U5124 (N_5124,N_2868,N_3516);
xnor U5125 (N_5125,N_1846,N_1463);
nor U5126 (N_5126,N_2890,N_2302);
or U5127 (N_5127,N_2462,N_425);
or U5128 (N_5128,N_3878,N_3225);
nor U5129 (N_5129,N_2117,N_3194);
or U5130 (N_5130,N_813,N_2092);
nor U5131 (N_5131,N_2985,N_4);
nand U5132 (N_5132,N_773,N_1820);
or U5133 (N_5133,N_1686,N_3558);
nor U5134 (N_5134,N_2447,N_3011);
and U5135 (N_5135,N_265,N_3304);
or U5136 (N_5136,N_663,N_2543);
nand U5137 (N_5137,N_2566,N_595);
or U5138 (N_5138,N_1162,N_1213);
nand U5139 (N_5139,N_59,N_3102);
or U5140 (N_5140,N_2170,N_949);
xnor U5141 (N_5141,N_886,N_1610);
nand U5142 (N_5142,N_3379,N_2411);
nand U5143 (N_5143,N_3383,N_1386);
nor U5144 (N_5144,N_473,N_1765);
and U5145 (N_5145,N_3214,N_2889);
or U5146 (N_5146,N_3162,N_1418);
and U5147 (N_5147,N_3440,N_294);
nand U5148 (N_5148,N_1078,N_2076);
nand U5149 (N_5149,N_2569,N_509);
or U5150 (N_5150,N_621,N_70);
nand U5151 (N_5151,N_1080,N_941);
nand U5152 (N_5152,N_1110,N_440);
nand U5153 (N_5153,N_2110,N_3069);
nand U5154 (N_5154,N_1008,N_683);
and U5155 (N_5155,N_2186,N_3853);
nor U5156 (N_5156,N_1629,N_3637);
xor U5157 (N_5157,N_3871,N_151);
or U5158 (N_5158,N_2198,N_1872);
xnor U5159 (N_5159,N_616,N_2493);
nor U5160 (N_5160,N_2386,N_3043);
and U5161 (N_5161,N_3904,N_2820);
and U5162 (N_5162,N_1139,N_1372);
nand U5163 (N_5163,N_223,N_310);
or U5164 (N_5164,N_1376,N_145);
and U5165 (N_5165,N_796,N_1210);
xor U5166 (N_5166,N_2584,N_1876);
or U5167 (N_5167,N_2834,N_3993);
nor U5168 (N_5168,N_180,N_3252);
xor U5169 (N_5169,N_1465,N_3165);
and U5170 (N_5170,N_2995,N_3776);
nand U5171 (N_5171,N_1264,N_18);
and U5172 (N_5172,N_492,N_3765);
and U5173 (N_5173,N_1750,N_3773);
nand U5174 (N_5174,N_2209,N_2515);
or U5175 (N_5175,N_2426,N_3130);
nor U5176 (N_5176,N_441,N_3919);
or U5177 (N_5177,N_830,N_593);
nand U5178 (N_5178,N_1953,N_708);
nor U5179 (N_5179,N_2943,N_3905);
or U5180 (N_5180,N_415,N_955);
nor U5181 (N_5181,N_169,N_1095);
and U5182 (N_5182,N_3990,N_3317);
nand U5183 (N_5183,N_3979,N_236);
or U5184 (N_5184,N_1854,N_790);
and U5185 (N_5185,N_1513,N_1321);
nor U5186 (N_5186,N_1789,N_1368);
xor U5187 (N_5187,N_358,N_3590);
or U5188 (N_5188,N_1548,N_2388);
nor U5189 (N_5189,N_1669,N_562);
nor U5190 (N_5190,N_3427,N_3350);
nor U5191 (N_5191,N_3482,N_3075);
or U5192 (N_5192,N_2987,N_2216);
xnor U5193 (N_5193,N_992,N_2765);
or U5194 (N_5194,N_2492,N_2522);
and U5195 (N_5195,N_1216,N_3530);
or U5196 (N_5196,N_3699,N_3830);
nand U5197 (N_5197,N_2291,N_251);
nand U5198 (N_5198,N_3169,N_1919);
nand U5199 (N_5199,N_327,N_742);
or U5200 (N_5200,N_2256,N_1668);
and U5201 (N_5201,N_391,N_1917);
or U5202 (N_5202,N_2509,N_1072);
or U5203 (N_5203,N_1461,N_848);
and U5204 (N_5204,N_2496,N_213);
nor U5205 (N_5205,N_479,N_3987);
and U5206 (N_5206,N_3622,N_2510);
or U5207 (N_5207,N_1001,N_2589);
or U5208 (N_5208,N_1707,N_800);
and U5209 (N_5209,N_2633,N_1987);
or U5210 (N_5210,N_2705,N_1899);
and U5211 (N_5211,N_3054,N_934);
nor U5212 (N_5212,N_3466,N_913);
nor U5213 (N_5213,N_1871,N_689);
nand U5214 (N_5214,N_1497,N_471);
and U5215 (N_5215,N_316,N_463);
and U5216 (N_5216,N_2645,N_3098);
and U5217 (N_5217,N_1928,N_2403);
nand U5218 (N_5218,N_3235,N_707);
xnor U5219 (N_5219,N_905,N_3757);
nand U5220 (N_5220,N_2315,N_1549);
or U5221 (N_5221,N_2708,N_600);
nor U5222 (N_5222,N_3439,N_1026);
nand U5223 (N_5223,N_518,N_2711);
xor U5224 (N_5224,N_2893,N_222);
nand U5225 (N_5225,N_3116,N_901);
and U5226 (N_5226,N_764,N_2516);
nand U5227 (N_5227,N_2269,N_167);
nor U5228 (N_5228,N_2590,N_1760);
xnor U5229 (N_5229,N_157,N_3099);
nor U5230 (N_5230,N_2113,N_2147);
and U5231 (N_5231,N_516,N_997);
or U5232 (N_5232,N_1862,N_3611);
nor U5233 (N_5233,N_3063,N_2859);
nor U5234 (N_5234,N_3322,N_2079);
or U5235 (N_5235,N_916,N_2340);
or U5236 (N_5236,N_1583,N_1182);
and U5237 (N_5237,N_48,N_2911);
xnor U5238 (N_5238,N_2458,N_377);
xnor U5239 (N_5239,N_182,N_3367);
nand U5240 (N_5240,N_1347,N_1269);
nand U5241 (N_5241,N_2731,N_3816);
and U5242 (N_5242,N_2478,N_654);
or U5243 (N_5243,N_1874,N_2692);
nand U5244 (N_5244,N_3144,N_111);
nand U5245 (N_5245,N_2300,N_3502);
nor U5246 (N_5246,N_1511,N_1359);
nand U5247 (N_5247,N_3750,N_274);
nor U5248 (N_5248,N_3838,N_3184);
nand U5249 (N_5249,N_3813,N_432);
nor U5250 (N_5250,N_3806,N_2640);
or U5251 (N_5251,N_3729,N_2826);
nand U5252 (N_5252,N_2191,N_2803);
nand U5253 (N_5253,N_2112,N_514);
or U5254 (N_5254,N_3110,N_1540);
nand U5255 (N_5255,N_2193,N_2675);
nand U5256 (N_5256,N_2687,N_3071);
nor U5257 (N_5257,N_3343,N_39);
and U5258 (N_5258,N_1661,N_3583);
xnor U5259 (N_5259,N_972,N_314);
and U5260 (N_5260,N_3399,N_1225);
nand U5261 (N_5261,N_3633,N_560);
nor U5262 (N_5262,N_1522,N_3627);
or U5263 (N_5263,N_3559,N_193);
or U5264 (N_5264,N_2377,N_290);
nor U5265 (N_5265,N_2125,N_1556);
or U5266 (N_5266,N_3348,N_3674);
xor U5267 (N_5267,N_1099,N_1941);
nand U5268 (N_5268,N_617,N_3312);
or U5269 (N_5269,N_2060,N_1806);
xnor U5270 (N_5270,N_2827,N_3411);
nand U5271 (N_5271,N_108,N_1141);
or U5272 (N_5272,N_1873,N_3215);
nor U5273 (N_5273,N_2927,N_3575);
or U5274 (N_5274,N_3856,N_3761);
and U5275 (N_5275,N_2023,N_2318);
nor U5276 (N_5276,N_1498,N_1369);
nor U5277 (N_5277,N_3963,N_3028);
or U5278 (N_5278,N_2553,N_2888);
and U5279 (N_5279,N_2390,N_2730);
nor U5280 (N_5280,N_47,N_2875);
xor U5281 (N_5281,N_1381,N_3996);
nor U5282 (N_5282,N_798,N_3843);
nand U5283 (N_5283,N_1479,N_1955);
and U5284 (N_5284,N_3026,N_1974);
nand U5285 (N_5285,N_2621,N_515);
nand U5286 (N_5286,N_3247,N_2101);
nor U5287 (N_5287,N_513,N_3113);
and U5288 (N_5288,N_3311,N_829);
xnor U5289 (N_5289,N_2961,N_3219);
xnor U5290 (N_5290,N_3503,N_2677);
or U5291 (N_5291,N_131,N_3899);
or U5292 (N_5292,N_272,N_1214);
nand U5293 (N_5293,N_1842,N_1272);
nand U5294 (N_5294,N_3064,N_3641);
and U5295 (N_5295,N_751,N_68);
nand U5296 (N_5296,N_719,N_2547);
xor U5297 (N_5297,N_3586,N_669);
or U5298 (N_5298,N_1023,N_840);
or U5299 (N_5299,N_1395,N_2973);
or U5300 (N_5300,N_2331,N_3303);
nor U5301 (N_5301,N_2118,N_1520);
nor U5302 (N_5302,N_363,N_704);
nand U5303 (N_5303,N_454,N_1449);
nor U5304 (N_5304,N_1986,N_325);
nand U5305 (N_5305,N_3053,N_50);
and U5306 (N_5306,N_436,N_2715);
and U5307 (N_5307,N_1829,N_192);
and U5308 (N_5308,N_11,N_539);
nor U5309 (N_5309,N_324,N_3250);
or U5310 (N_5310,N_2181,N_1502);
nor U5311 (N_5311,N_2679,N_2572);
nor U5312 (N_5312,N_113,N_2805);
nand U5313 (N_5313,N_2352,N_2763);
xor U5314 (N_5314,N_1798,N_2851);
xor U5315 (N_5315,N_1525,N_46);
and U5316 (N_5316,N_1075,N_2520);
or U5317 (N_5317,N_3364,N_1982);
or U5318 (N_5318,N_3976,N_3227);
and U5319 (N_5319,N_3068,N_2354);
nor U5320 (N_5320,N_278,N_3147);
nand U5321 (N_5321,N_2994,N_3433);
or U5322 (N_5322,N_3015,N_1329);
nor U5323 (N_5323,N_818,N_2211);
xor U5324 (N_5324,N_1908,N_591);
or U5325 (N_5325,N_3354,N_1265);
nand U5326 (N_5326,N_3690,N_2124);
and U5327 (N_5327,N_2563,N_3698);
or U5328 (N_5328,N_2914,N_910);
nand U5329 (N_5329,N_1555,N_2078);
xnor U5330 (N_5330,N_2432,N_3578);
or U5331 (N_5331,N_371,N_3662);
or U5332 (N_5332,N_2116,N_1085);
xnor U5333 (N_5333,N_791,N_1644);
and U5334 (N_5334,N_2636,N_1471);
nor U5335 (N_5335,N_781,N_3694);
nor U5336 (N_5336,N_2823,N_1018);
and U5337 (N_5337,N_1473,N_915);
or U5338 (N_5338,N_1804,N_746);
xor U5339 (N_5339,N_859,N_1388);
nand U5340 (N_5340,N_3731,N_2772);
and U5341 (N_5341,N_405,N_1638);
and U5342 (N_5342,N_2505,N_783);
and U5343 (N_5343,N_485,N_1060);
or U5344 (N_5344,N_1039,N_2847);
or U5345 (N_5345,N_1363,N_1890);
nor U5346 (N_5346,N_2930,N_2953);
xor U5347 (N_5347,N_2600,N_2357);
nor U5348 (N_5348,N_2208,N_1809);
or U5349 (N_5349,N_3759,N_3778);
nor U5350 (N_5350,N_2694,N_458);
or U5351 (N_5351,N_3261,N_1174);
nor U5352 (N_5352,N_3444,N_2260);
or U5353 (N_5353,N_1680,N_3560);
nand U5354 (N_5354,N_1937,N_809);
xor U5355 (N_5355,N_1303,N_1066);
xor U5356 (N_5356,N_2310,N_1153);
or U5357 (N_5357,N_1146,N_3980);
xor U5358 (N_5358,N_2549,N_1949);
and U5359 (N_5359,N_1673,N_2877);
and U5360 (N_5360,N_2237,N_966);
and U5361 (N_5361,N_803,N_2529);
xnor U5362 (N_5362,N_774,N_2693);
nor U5363 (N_5363,N_2533,N_1477);
nor U5364 (N_5364,N_1290,N_2935);
or U5365 (N_5365,N_1476,N_1780);
or U5366 (N_5366,N_3253,N_3470);
or U5367 (N_5367,N_2360,N_2597);
and U5368 (N_5368,N_342,N_3271);
nor U5369 (N_5369,N_3626,N_3385);
and U5370 (N_5370,N_1289,N_2279);
xor U5371 (N_5371,N_1577,N_3567);
xor U5372 (N_5372,N_1599,N_289);
nor U5373 (N_5373,N_394,N_2422);
nand U5374 (N_5374,N_982,N_2392);
xor U5375 (N_5375,N_2289,N_718);
and U5376 (N_5376,N_2594,N_3720);
and U5377 (N_5377,N_2151,N_269);
and U5378 (N_5378,N_903,N_665);
and U5379 (N_5379,N_3967,N_902);
and U5380 (N_5380,N_3036,N_3180);
or U5381 (N_5381,N_2258,N_1633);
nand U5382 (N_5382,N_1343,N_643);
and U5383 (N_5383,N_3636,N_1885);
nor U5384 (N_5384,N_2464,N_1778);
or U5385 (N_5385,N_331,N_1116);
nand U5386 (N_5386,N_1838,N_3202);
and U5387 (N_5387,N_682,N_1759);
or U5388 (N_5388,N_3398,N_2308);
nor U5389 (N_5389,N_1132,N_1103);
or U5390 (N_5390,N_3534,N_2415);
or U5391 (N_5391,N_1035,N_1131);
or U5392 (N_5392,N_1507,N_354);
nand U5393 (N_5393,N_1752,N_2204);
nor U5394 (N_5394,N_285,N_2382);
nand U5395 (N_5395,N_404,N_2824);
and U5396 (N_5396,N_1617,N_3206);
or U5397 (N_5397,N_2801,N_770);
nor U5398 (N_5398,N_3196,N_823);
nand U5399 (N_5399,N_638,N_174);
and U5400 (N_5400,N_3109,N_726);
or U5401 (N_5401,N_2776,N_607);
xnor U5402 (N_5402,N_3292,N_2212);
nor U5403 (N_5403,N_2451,N_6);
or U5404 (N_5404,N_1963,N_2088);
nand U5405 (N_5405,N_0,N_3362);
xor U5406 (N_5406,N_2002,N_1864);
and U5407 (N_5407,N_1154,N_2901);
or U5408 (N_5408,N_1912,N_2114);
or U5409 (N_5409,N_2871,N_378);
nand U5410 (N_5410,N_1647,N_2970);
xnor U5411 (N_5411,N_695,N_2524);
nor U5412 (N_5412,N_2066,N_2650);
nand U5413 (N_5413,N_364,N_3495);
nand U5414 (N_5414,N_1212,N_3651);
or U5415 (N_5415,N_302,N_443);
and U5416 (N_5416,N_396,N_387);
nand U5417 (N_5417,N_712,N_3712);
nor U5418 (N_5418,N_1814,N_2521);
or U5419 (N_5419,N_2272,N_825);
and U5420 (N_5420,N_1622,N_1787);
and U5421 (N_5421,N_609,N_2402);
or U5422 (N_5422,N_3040,N_3988);
or U5423 (N_5423,N_999,N_3203);
nand U5424 (N_5424,N_700,N_2573);
nand U5425 (N_5425,N_3051,N_312);
nor U5426 (N_5426,N_3518,N_1328);
and U5427 (N_5427,N_1510,N_1387);
nand U5428 (N_5428,N_3397,N_527);
nand U5429 (N_5429,N_2745,N_3237);
and U5430 (N_5430,N_3852,N_3275);
and U5431 (N_5431,N_19,N_1030);
nor U5432 (N_5432,N_3107,N_2167);
nor U5433 (N_5433,N_2271,N_292);
nor U5434 (N_5434,N_2139,N_5);
nand U5435 (N_5435,N_2691,N_3230);
and U5436 (N_5436,N_681,N_1832);
nor U5437 (N_5437,N_57,N_3865);
nor U5438 (N_5438,N_2956,N_3342);
nor U5439 (N_5439,N_149,N_1732);
nor U5440 (N_5440,N_1851,N_2717);
and U5441 (N_5441,N_2140,N_973);
nor U5442 (N_5442,N_1468,N_3718);
nand U5443 (N_5443,N_3309,N_3740);
or U5444 (N_5444,N_666,N_2798);
nor U5445 (N_5445,N_1466,N_3070);
and U5446 (N_5446,N_520,N_2056);
nor U5447 (N_5447,N_3492,N_990);
and U5448 (N_5448,N_346,N_758);
nand U5449 (N_5449,N_571,N_3644);
nor U5450 (N_5450,N_3675,N_348);
or U5451 (N_5451,N_232,N_3764);
nand U5452 (N_5452,N_581,N_3458);
xor U5453 (N_5453,N_854,N_2156);
nor U5454 (N_5454,N_2454,N_3298);
nand U5455 (N_5455,N_2049,N_10);
or U5456 (N_5456,N_1541,N_2501);
nor U5457 (N_5457,N_2227,N_1568);
xnor U5458 (N_5458,N_2862,N_73);
and U5459 (N_5459,N_1051,N_1792);
nand U5460 (N_5460,N_96,N_1160);
nor U5461 (N_5461,N_2184,N_3910);
and U5462 (N_5462,N_1659,N_2182);
or U5463 (N_5463,N_1245,N_2947);
nor U5464 (N_5464,N_82,N_1248);
and U5465 (N_5465,N_3193,N_952);
and U5466 (N_5466,N_3210,N_996);
or U5467 (N_5467,N_470,N_3289);
and U5468 (N_5468,N_2083,N_2620);
and U5469 (N_5469,N_2036,N_1011);
nor U5470 (N_5470,N_2611,N_566);
nor U5471 (N_5471,N_3321,N_2025);
nor U5472 (N_5472,N_2988,N_878);
and U5473 (N_5473,N_1065,N_3395);
and U5474 (N_5474,N_410,N_2581);
nand U5475 (N_5475,N_667,N_1841);
and U5476 (N_5476,N_831,N_1165);
or U5477 (N_5477,N_2669,N_3546);
or U5478 (N_5478,N_2369,N_1222);
xor U5479 (N_5479,N_2747,N_1356);
and U5480 (N_5480,N_1757,N_293);
nor U5481 (N_5481,N_1582,N_2903);
and U5482 (N_5482,N_1168,N_3280);
or U5483 (N_5483,N_399,N_2370);
nor U5484 (N_5484,N_1360,N_2285);
or U5485 (N_5485,N_381,N_957);
and U5486 (N_5486,N_3006,N_372);
or U5487 (N_5487,N_3489,N_64);
and U5488 (N_5488,N_3085,N_599);
nand U5489 (N_5489,N_1571,N_3609);
nor U5490 (N_5490,N_3580,N_233);
nor U5491 (N_5491,N_1799,N_161);
and U5492 (N_5492,N_2436,N_956);
and U5493 (N_5493,N_2737,N_1284);
and U5494 (N_5494,N_544,N_3335);
nand U5495 (N_5495,N_995,N_1298);
and U5496 (N_5496,N_693,N_1761);
xnor U5497 (N_5497,N_1731,N_1206);
nor U5498 (N_5498,N_3515,N_1745);
or U5499 (N_5499,N_3582,N_804);
or U5500 (N_5500,N_1687,N_787);
and U5501 (N_5501,N_3997,N_3396);
or U5502 (N_5502,N_2815,N_2128);
xor U5503 (N_5503,N_3449,N_245);
or U5504 (N_5504,N_1521,N_1251);
nor U5505 (N_5505,N_2119,N_2480);
nand U5506 (N_5506,N_376,N_1758);
nand U5507 (N_5507,N_2602,N_2844);
nand U5508 (N_5508,N_3725,N_1650);
nor U5509 (N_5509,N_1420,N_3287);
or U5510 (N_5510,N_2619,N_671);
or U5511 (N_5511,N_3451,N_1239);
xor U5512 (N_5512,N_1196,N_1693);
nor U5513 (N_5513,N_3669,N_532);
nand U5514 (N_5514,N_3272,N_2393);
xnor U5515 (N_5515,N_55,N_2818);
and U5516 (N_5516,N_3142,N_1646);
nand U5517 (N_5517,N_241,N_3046);
and U5518 (N_5518,N_3891,N_1503);
nand U5519 (N_5519,N_1641,N_2407);
nor U5520 (N_5520,N_160,N_3786);
and U5521 (N_5521,N_1609,N_2472);
nand U5522 (N_5522,N_242,N_1823);
or U5523 (N_5523,N_810,N_1563);
or U5524 (N_5524,N_2026,N_1094);
or U5525 (N_5525,N_710,N_1309);
nand U5526 (N_5526,N_2642,N_873);
nor U5527 (N_5527,N_107,N_2362);
or U5528 (N_5528,N_3232,N_2907);
nand U5529 (N_5529,N_3246,N_2942);
or U5530 (N_5530,N_3418,N_1781);
nor U5531 (N_5531,N_969,N_3301);
nand U5532 (N_5532,N_3744,N_2361);
and U5533 (N_5533,N_3864,N_3754);
nand U5534 (N_5534,N_43,N_3966);
and U5535 (N_5535,N_2822,N_3505);
nor U5536 (N_5536,N_3991,N_3016);
and U5537 (N_5537,N_3706,N_2884);
nand U5538 (N_5538,N_534,N_2948);
nor U5539 (N_5539,N_1785,N_282);
nor U5540 (N_5540,N_1523,N_1744);
nand U5541 (N_5541,N_2467,N_2280);
or U5542 (N_5542,N_2004,N_2262);
nand U5543 (N_5543,N_856,N_3511);
xor U5544 (N_5544,N_2148,N_3442);
nor U5545 (N_5545,N_446,N_2194);
or U5546 (N_5546,N_3409,N_3331);
xor U5547 (N_5547,N_286,N_871);
and U5548 (N_5548,N_2008,N_2936);
nand U5549 (N_5549,N_3923,N_737);
nor U5550 (N_5550,N_2904,N_2240);
nand U5551 (N_5551,N_2192,N_155);
nand U5552 (N_5552,N_2664,N_2879);
nor U5553 (N_5553,N_1405,N_3721);
nand U5554 (N_5554,N_1404,N_3377);
and U5555 (N_5555,N_3106,N_2874);
nand U5556 (N_5556,N_2303,N_2878);
nand U5557 (N_5557,N_1739,N_2726);
xnor U5558 (N_5558,N_1007,N_2787);
xnor U5559 (N_5559,N_2277,N_648);
and U5560 (N_5560,N_559,N_2729);
nand U5561 (N_5561,N_297,N_631);
nand U5562 (N_5562,N_828,N_1341);
nor U5563 (N_5563,N_734,N_2463);
nand U5564 (N_5564,N_2885,N_1100);
and U5565 (N_5565,N_3067,N_1422);
nor U5566 (N_5566,N_2259,N_275);
or U5567 (N_5567,N_3541,N_989);
or U5568 (N_5568,N_563,N_2556);
nor U5569 (N_5569,N_711,N_2544);
xor U5570 (N_5570,N_2806,N_3614);
and U5571 (N_5571,N_3405,N_2843);
nor U5572 (N_5572,N_1943,N_3146);
nor U5573 (N_5573,N_1062,N_2334);
nor U5574 (N_5574,N_486,N_852);
xor U5575 (N_5575,N_2575,N_976);
or U5576 (N_5576,N_1863,N_3884);
xor U5577 (N_5577,N_3300,N_2341);
nand U5578 (N_5578,N_855,N_429);
xor U5579 (N_5579,N_1114,N_3368);
or U5580 (N_5580,N_244,N_2380);
or U5581 (N_5581,N_3953,N_2895);
xor U5582 (N_5582,N_573,N_2902);
or U5583 (N_5583,N_1188,N_1097);
nor U5584 (N_5584,N_361,N_1113);
nand U5585 (N_5585,N_1184,N_13);
or U5586 (N_5586,N_127,N_2055);
and U5587 (N_5587,N_567,N_2997);
nor U5588 (N_5588,N_565,N_2409);
and U5589 (N_5589,N_2345,N_453);
and U5590 (N_5590,N_1714,N_2983);
xor U5591 (N_5591,N_574,N_724);
nor U5592 (N_5592,N_1148,N_1586);
nand U5593 (N_5593,N_1801,N_8);
nor U5594 (N_5594,N_3197,N_1203);
and U5595 (N_5595,N_2460,N_2836);
nand U5596 (N_5596,N_1976,N_1349);
nand U5597 (N_5597,N_3159,N_552);
nand U5598 (N_5598,N_3529,N_2150);
nor U5599 (N_5599,N_1231,N_1385);
nor U5600 (N_5600,N_2485,N_143);
or U5601 (N_5601,N_34,N_1320);
or U5602 (N_5602,N_185,N_1);
or U5603 (N_5603,N_2962,N_2305);
and U5604 (N_5604,N_2102,N_3846);
or U5605 (N_5605,N_1457,N_3820);
nand U5606 (N_5606,N_1048,N_99);
or U5607 (N_5607,N_3052,N_1774);
nor U5608 (N_5608,N_374,N_188);
nor U5609 (N_5609,N_729,N_3369);
xnor U5610 (N_5610,N_1118,N_2882);
nor U5611 (N_5611,N_1068,N_1536);
or U5612 (N_5612,N_1427,N_1725);
nor U5613 (N_5613,N_1127,N_3727);
nand U5614 (N_5614,N_974,N_319);
and U5615 (N_5615,N_466,N_3595);
and U5616 (N_5616,N_1691,N_3978);
or U5617 (N_5617,N_2082,N_889);
or U5618 (N_5618,N_23,N_137);
or U5619 (N_5619,N_1705,N_3844);
xnor U5620 (N_5620,N_3973,N_3133);
nor U5621 (N_5621,N_3245,N_3447);
and U5622 (N_5622,N_2164,N_3975);
nor U5623 (N_5623,N_2845,N_2109);
or U5624 (N_5624,N_1748,N_1353);
xor U5625 (N_5625,N_487,N_3552);
nor U5626 (N_5626,N_3428,N_554);
or U5627 (N_5627,N_434,N_279);
and U5628 (N_5628,N_119,N_3920);
nor U5629 (N_5629,N_1150,N_2136);
and U5630 (N_5630,N_935,N_33);
xor U5631 (N_5631,N_3341,N_1771);
nor U5632 (N_5632,N_2013,N_12);
and U5633 (N_5633,N_1635,N_2103);
and U5634 (N_5634,N_3921,N_2778);
nand U5635 (N_5635,N_2456,N_782);
or U5636 (N_5636,N_1379,N_3832);
nand U5637 (N_5637,N_850,N_2963);
nand U5638 (N_5638,N_3914,N_1848);
nand U5639 (N_5639,N_3299,N_1045);
and U5640 (N_5640,N_1133,N_3982);
nor U5641 (N_5641,N_2077,N_2185);
or U5642 (N_5642,N_1727,N_3216);
and U5643 (N_5643,N_1741,N_277);
nand U5644 (N_5644,N_948,N_1448);
nand U5645 (N_5645,N_980,N_1896);
and U5646 (N_5646,N_3254,N_2297);
nor U5647 (N_5647,N_3911,N_2616);
xor U5648 (N_5648,N_2793,N_2225);
and U5649 (N_5649,N_583,N_2550);
and U5650 (N_5650,N_3404,N_1754);
xor U5651 (N_5651,N_2599,N_2338);
or U5652 (N_5652,N_3437,N_3577);
nor U5653 (N_5653,N_750,N_1169);
xnor U5654 (N_5654,N_3972,N_1057);
nor U5655 (N_5655,N_2232,N_2230);
and U5656 (N_5656,N_2238,N_2643);
nand U5657 (N_5657,N_1670,N_1378);
and U5658 (N_5658,N_940,N_3226);
nor U5659 (N_5659,N_2439,N_416);
or U5660 (N_5660,N_2010,N_3282);
nor U5661 (N_5661,N_92,N_3296);
and U5662 (N_5662,N_3587,N_832);
xor U5663 (N_5663,N_1331,N_3616);
and U5664 (N_5664,N_1370,N_2703);
or U5665 (N_5665,N_3854,N_3462);
and U5666 (N_5666,N_3876,N_1192);
nor U5667 (N_5667,N_2199,N_3207);
nor U5668 (N_5668,N_2323,N_649);
or U5669 (N_5669,N_3665,N_1542);
nand U5670 (N_5670,N_650,N_2358);
xnor U5671 (N_5671,N_2760,N_1010);
xor U5672 (N_5672,N_2949,N_3822);
or U5673 (N_5673,N_3845,N_3380);
and U5674 (N_5674,N_3465,N_250);
xnor U5675 (N_5675,N_3600,N_1362);
nand U5676 (N_5676,N_493,N_1933);
nand U5677 (N_5677,N_1425,N_2489);
nor U5678 (N_5678,N_3255,N_3087);
or U5679 (N_5679,N_1595,N_686);
nand U5680 (N_5680,N_705,N_1142);
or U5681 (N_5681,N_2558,N_1645);
and U5682 (N_5682,N_2689,N_3461);
nand U5683 (N_5683,N_1083,N_725);
nor U5684 (N_5684,N_506,N_2085);
or U5685 (N_5685,N_1616,N_1740);
nand U5686 (N_5686,N_1930,N_37);
nand U5687 (N_5687,N_3667,N_1539);
xnor U5688 (N_5688,N_2288,N_3900);
and U5689 (N_5689,N_3188,N_1636);
or U5690 (N_5690,N_3549,N_2743);
or U5691 (N_5691,N_793,N_2121);
or U5692 (N_5692,N_3945,N_3061);
nand U5693 (N_5693,N_1415,N_2706);
and U5694 (N_5694,N_926,N_3833);
nor U5695 (N_5695,N_3524,N_2175);
and U5696 (N_5696,N_735,N_144);
and U5697 (N_5697,N_3228,N_2698);
and U5698 (N_5698,N_2819,N_778);
nor U5699 (N_5699,N_2301,N_3807);
and U5700 (N_5700,N_3801,N_2659);
or U5701 (N_5701,N_1715,N_1215);
nor U5702 (N_5702,N_1325,N_1935);
nor U5703 (N_5703,N_1600,N_3895);
nor U5704 (N_5704,N_3802,N_239);
or U5705 (N_5705,N_545,N_512);
nor U5706 (N_5706,N_1052,N_3984);
and U5707 (N_5707,N_547,N_24);
nand U5708 (N_5708,N_3477,N_1592);
nand U5709 (N_5709,N_3389,N_183);
and U5710 (N_5710,N_3628,N_3943);
nand U5711 (N_5711,N_3959,N_860);
nor U5712 (N_5712,N_1681,N_1777);
xnor U5713 (N_5713,N_3013,N_1527);
nor U5714 (N_5714,N_658,N_3934);
or U5715 (N_5715,N_1033,N_197);
nand U5716 (N_5716,N_3393,N_3308);
nor U5717 (N_5717,N_1621,N_1559);
nand U5718 (N_5718,N_3158,N_619);
and U5719 (N_5719,N_555,N_870);
or U5720 (N_5720,N_3352,N_1024);
and U5721 (N_5721,N_1710,N_2897);
nor U5722 (N_5722,N_2000,N_3798);
nand U5723 (N_5723,N_1589,N_2425);
or U5724 (N_5724,N_2925,N_3906);
or U5725 (N_5725,N_3119,N_3167);
nand U5726 (N_5726,N_3471,N_3889);
xnor U5727 (N_5727,N_3701,N_1767);
nor U5728 (N_5728,N_1649,N_1056);
or U5729 (N_5729,N_1013,N_3624);
and U5730 (N_5730,N_846,N_2909);
xor U5731 (N_5731,N_1702,N_1790);
or U5732 (N_5732,N_2242,N_2761);
and U5733 (N_5733,N_3339,N_1163);
or U5734 (N_5734,N_1504,N_2568);
and U5735 (N_5735,N_3378,N_2252);
nand U5736 (N_5736,N_673,N_584);
or U5737 (N_5737,N_3867,N_1786);
or U5738 (N_5738,N_49,N_507);
nand U5739 (N_5739,N_890,N_1870);
nor U5740 (N_5740,N_3692,N_3557);
nor U5741 (N_5741,N_613,N_1436);
nand U5742 (N_5742,N_3191,N_3496);
nor U5743 (N_5743,N_2783,N_3649);
and U5744 (N_5744,N_2448,N_733);
or U5745 (N_5745,N_3849,N_1728);
nand U5746 (N_5746,N_2733,N_3224);
or U5747 (N_5747,N_3258,N_642);
nand U5748 (N_5748,N_2050,N_1123);
and U5749 (N_5749,N_2440,N_3438);
or U5750 (N_5750,N_2,N_2427);
and U5751 (N_5751,N_3135,N_1237);
nor U5752 (N_5752,N_1478,N_262);
nand U5753 (N_5753,N_1028,N_1808);
and U5754 (N_5754,N_488,N_3363);
nand U5755 (N_5755,N_1292,N_525);
nor U5756 (N_5756,N_344,N_3916);
nand U5757 (N_5757,N_3936,N_723);
nor U5758 (N_5758,N_3784,N_260);
or U5759 (N_5759,N_696,N_1408);
or U5760 (N_5760,N_1570,N_853);
nand U5761 (N_5761,N_2385,N_2051);
nor U5762 (N_5762,N_3635,N_1701);
and U5763 (N_5763,N_1034,N_620);
and U5764 (N_5764,N_1580,N_1074);
nand U5765 (N_5765,N_420,N_1961);
nand U5766 (N_5766,N_1836,N_2267);
xnor U5767 (N_5767,N_221,N_2946);
nand U5768 (N_5768,N_2214,N_728);
or U5769 (N_5769,N_3490,N_606);
nor U5770 (N_5770,N_2606,N_1753);
and U5771 (N_5771,N_1712,N_218);
or U5772 (N_5772,N_498,N_819);
nor U5773 (N_5773,N_2716,N_3702);
or U5774 (N_5774,N_2799,N_496);
nor U5775 (N_5775,N_3170,N_2160);
xor U5776 (N_5776,N_2284,N_3145);
or U5777 (N_5777,N_777,N_1373);
xor U5778 (N_5778,N_26,N_1495);
nor U5779 (N_5779,N_688,N_2583);
and U5780 (N_5780,N_3424,N_258);
and U5781 (N_5781,N_36,N_3392);
nor U5782 (N_5782,N_1565,N_1120);
and U5783 (N_5783,N_2982,N_2720);
and U5784 (N_5784,N_2187,N_2832);
nor U5785 (N_5785,N_1879,N_2444);
and U5786 (N_5786,N_2196,N_1423);
or U5787 (N_5787,N_634,N_1167);
xor U5788 (N_5788,N_2814,N_1721);
and U5789 (N_5789,N_2394,N_1276);
and U5790 (N_5790,N_2468,N_3782);
and U5791 (N_5791,N_3850,N_2379);
and U5792 (N_5792,N_1079,N_1394);
nor U5793 (N_5793,N_587,N_690);
xnor U5794 (N_5794,N_2449,N_2317);
or U5795 (N_5795,N_1575,N_3048);
and U5796 (N_5796,N_3779,N_284);
or U5797 (N_5797,N_2398,N_3073);
xnor U5798 (N_5798,N_191,N_675);
or U5799 (N_5799,N_159,N_3365);
nand U5800 (N_5800,N_3370,N_95);
nand U5801 (N_5801,N_3774,N_1920);
or U5802 (N_5802,N_106,N_1611);
xor U5803 (N_5803,N_490,N_3564);
and U5804 (N_5804,N_1770,N_1509);
and U5805 (N_5805,N_3763,N_2923);
and U5806 (N_5806,N_3218,N_1352);
xor U5807 (N_5807,N_449,N_2265);
nand U5808 (N_5808,N_3157,N_1022);
nand U5809 (N_5809,N_2848,N_2740);
nor U5810 (N_5810,N_3314,N_3805);
nor U5811 (N_5811,N_2236,N_476);
nor U5812 (N_5812,N_3668,N_120);
or U5813 (N_5813,N_1604,N_1738);
xor U5814 (N_5814,N_2325,N_1755);
nand U5815 (N_5815,N_379,N_198);
nor U5816 (N_5816,N_3969,N_406);
nand U5817 (N_5817,N_1900,N_2714);
xor U5818 (N_5818,N_2512,N_598);
nand U5819 (N_5819,N_1564,N_418);
and U5820 (N_5820,N_3676,N_1560);
and U5821 (N_5821,N_359,N_1566);
nand U5822 (N_5822,N_32,N_1924);
or U5823 (N_5823,N_652,N_77);
nand U5824 (N_5824,N_1561,N_417);
nor U5825 (N_5825,N_317,N_2655);
or U5826 (N_5826,N_1909,N_2883);
nor U5827 (N_5827,N_3104,N_2657);
nor U5828 (N_5828,N_3315,N_2934);
nor U5829 (N_5829,N_799,N_900);
xor U5830 (N_5830,N_2989,N_335);
nor U5831 (N_5831,N_3848,N_1959);
nor U5832 (N_5832,N_1672,N_3039);
or U5833 (N_5833,N_519,N_1108);
or U5834 (N_5834,N_963,N_630);
or U5835 (N_5835,N_2542,N_336);
and U5836 (N_5836,N_3892,N_3450);
nand U5837 (N_5837,N_1256,N_1282);
and U5838 (N_5838,N_2784,N_1619);
nor U5839 (N_5839,N_1334,N_1128);
nand U5840 (N_5840,N_3260,N_2631);
or U5841 (N_5841,N_3325,N_1093);
or U5842 (N_5842,N_3338,N_3421);
nor U5843 (N_5843,N_3090,N_3553);
nor U5844 (N_5844,N_2069,N_1779);
or U5845 (N_5845,N_3898,N_895);
xor U5846 (N_5846,N_154,N_1412);
xor U5847 (N_5847,N_2950,N_2996);
and U5848 (N_5848,N_3494,N_1233);
and U5849 (N_5849,N_578,N_1773);
nor U5850 (N_5850,N_771,N_1573);
or U5851 (N_5851,N_2876,N_2438);
nand U5852 (N_5852,N_147,N_923);
xnor U5853 (N_5853,N_3394,N_2797);
and U5854 (N_5854,N_3607,N_349);
nor U5855 (N_5855,N_266,N_2931);
or U5856 (N_5856,N_824,N_1306);
or U5857 (N_5857,N_821,N_2188);
nand U5858 (N_5858,N_757,N_1501);
and U5859 (N_5859,N_114,N_1698);
xor U5860 (N_5860,N_3879,N_499);
nand U5861 (N_5861,N_3842,N_3486);
nor U5862 (N_5862,N_1878,N_1472);
or U5863 (N_5863,N_122,N_1366);
nand U5864 (N_5864,N_1696,N_1915);
xnor U5865 (N_5865,N_2045,N_2579);
nor U5866 (N_5866,N_2919,N_3588);
xnor U5867 (N_5867,N_557,N_3887);
nand U5868 (N_5868,N_912,N_858);
xor U5869 (N_5869,N_2159,N_1411);
and U5870 (N_5870,N_998,N_444);
or U5871 (N_5871,N_3406,N_629);
or U5872 (N_5872,N_1489,N_2541);
or U5873 (N_5873,N_435,N_2854);
and U5874 (N_5874,N_3326,N_1578);
xor U5875 (N_5875,N_1516,N_3156);
or U5876 (N_5876,N_3977,N_1096);
and U5877 (N_5877,N_2817,N_1772);
xnor U5878 (N_5878,N_3244,N_3903);
nor U5879 (N_5879,N_2596,N_2916);
nor U5880 (N_5880,N_2869,N_3680);
nor U5881 (N_5881,N_542,N_2908);
xor U5882 (N_5882,N_815,N_3686);
and U5883 (N_5883,N_2268,N_1630);
nand U5884 (N_5884,N_2658,N_2153);
nand U5885 (N_5885,N_1124,N_1822);
nor U5886 (N_5886,N_472,N_2873);
xnor U5887 (N_5887,N_1948,N_3033);
and U5888 (N_5888,N_3684,N_1445);
nor U5889 (N_5889,N_75,N_521);
and U5890 (N_5890,N_3388,N_2162);
nand U5891 (N_5891,N_3473,N_1688);
or U5892 (N_5892,N_3355,N_3728);
and U5893 (N_5893,N_2625,N_727);
nor U5894 (N_5894,N_2858,N_3572);
nor U5895 (N_5895,N_408,N_927);
or U5896 (N_5896,N_3551,N_3704);
nand U5897 (N_5897,N_1914,N_1709);
nand U5898 (N_5898,N_3952,N_1090);
nand U5899 (N_5899,N_564,N_1089);
xnor U5900 (N_5900,N_3741,N_1557);
or U5901 (N_5901,N_605,N_1603);
or U5902 (N_5902,N_1762,N_1371);
and U5903 (N_5903,N_140,N_2685);
nor U5904 (N_5904,N_1155,N_3777);
nor U5905 (N_5905,N_1897,N_865);
nor U5906 (N_5906,N_3682,N_226);
and U5907 (N_5907,N_2992,N_505);
nand U5908 (N_5908,N_1735,N_627);
nand U5909 (N_5909,N_1946,N_2965);
nor U5910 (N_5910,N_3504,N_1749);
xor U5911 (N_5911,N_1634,N_2011);
nand U5912 (N_5912,N_426,N_546);
and U5913 (N_5913,N_2408,N_3236);
and U5914 (N_5914,N_1295,N_2647);
and U5915 (N_5915,N_280,N_3928);
nor U5916 (N_5916,N_3785,N_2662);
nand U5917 (N_5917,N_304,N_3664);
or U5918 (N_5918,N_3327,N_2796);
or U5919 (N_5919,N_1073,N_90);
nand U5920 (N_5920,N_898,N_1335);
nor U5921 (N_5921,N_1901,N_932);
nand U5922 (N_5922,N_2683,N_1084);
and U5923 (N_5923,N_2825,N_2831);
and U5924 (N_5924,N_2674,N_639);
and U5925 (N_5925,N_1788,N_2567);
nor U5926 (N_5926,N_216,N_2537);
and U5927 (N_5927,N_2084,N_2072);
or U5928 (N_5928,N_1122,N_3386);
or U5929 (N_5929,N_1326,N_2414);
or U5930 (N_5930,N_3831,N_3539);
nor U5931 (N_5931,N_2100,N_2120);
nand U5932 (N_5932,N_1091,N_3241);
xor U5933 (N_5933,N_2030,N_1675);
nor U5934 (N_5934,N_1581,N_808);
xor U5935 (N_5935,N_1144,N_2434);
nor U5936 (N_5936,N_1990,N_2676);
or U5937 (N_5937,N_1441,N_20);
xnor U5938 (N_5938,N_93,N_395);
nor U5939 (N_5939,N_2752,N_3960);
and U5940 (N_5940,N_2058,N_1984);
and U5941 (N_5941,N_2938,N_3677);
nand U5942 (N_5942,N_2368,N_2336);
nor U5943 (N_5943,N_661,N_3908);
nor U5944 (N_5944,N_3901,N_3837);
nand U5945 (N_5945,N_2593,N_2330);
nor U5946 (N_5946,N_1579,N_775);
nor U5947 (N_5947,N_2508,N_1452);
and U5948 (N_5948,N_3336,N_3118);
nor U5949 (N_5949,N_2530,N_3294);
or U5950 (N_5950,N_2421,N_3623);
or U5951 (N_5951,N_678,N_2099);
nor U5952 (N_5952,N_400,N_1567);
nand U5953 (N_5953,N_3768,N_308);
nor U5954 (N_5954,N_402,N_1198);
or U5955 (N_5955,N_3456,N_2373);
or U5956 (N_5956,N_3453,N_2367);
and U5957 (N_5957,N_478,N_2786);
or U5958 (N_5958,N_2276,N_126);
or U5959 (N_5959,N_1653,N_647);
nor U5960 (N_5960,N_1242,N_1886);
nand U5961 (N_5961,N_1432,N_264);
nor U5962 (N_5962,N_795,N_3400);
nor U5963 (N_5963,N_2617,N_3488);
nand U5964 (N_5964,N_3243,N_40);
nand U5965 (N_5965,N_422,N_692);
nor U5966 (N_5966,N_3065,N_597);
nand U5967 (N_5967,N_1839,N_229);
and U5968 (N_5968,N_1004,N_204);
nor U5969 (N_5969,N_51,N_622);
nand U5970 (N_5970,N_2304,N_1967);
or U5971 (N_5971,N_3670,N_879);
xnor U5972 (N_5972,N_3408,N_3058);
or U5973 (N_5973,N_857,N_942);
nand U5974 (N_5974,N_210,N_1602);
nor U5975 (N_5975,N_1246,N_1954);
nand U5976 (N_5976,N_2707,N_1763);
nor U5977 (N_5977,N_1973,N_636);
or U5978 (N_5978,N_1000,N_908);
and U5979 (N_5979,N_1492,N_2329);
nor U5980 (N_5980,N_52,N_1397);
nand U5981 (N_5981,N_2122,N_200);
nor U5982 (N_5982,N_906,N_1053);
and U5983 (N_5983,N_1358,N_3200);
nand U5984 (N_5984,N_1407,N_1287);
nor U5985 (N_5985,N_1126,N_3683);
nand U5986 (N_5986,N_3882,N_3152);
or U5987 (N_5987,N_2612,N_340);
nand U5988 (N_5988,N_3817,N_3318);
or U5989 (N_5989,N_3800,N_2627);
or U5990 (N_5990,N_575,N_2968);
or U5991 (N_5991,N_872,N_3693);
or U5992 (N_5992,N_3957,N_442);
nand U5993 (N_5993,N_3234,N_1270);
or U5994 (N_5994,N_849,N_3042);
nand U5995 (N_5995,N_3448,N_2174);
xor U5996 (N_5996,N_2624,N_959);
xor U5997 (N_5997,N_347,N_1682);
and U5998 (N_5998,N_961,N_3155);
nor U5999 (N_5999,N_2484,N_2710);
nor U6000 (N_6000,N_216,N_2946);
nor U6001 (N_6001,N_3524,N_3538);
nor U6002 (N_6002,N_2159,N_2071);
or U6003 (N_6003,N_2428,N_3937);
and U6004 (N_6004,N_739,N_3855);
nand U6005 (N_6005,N_2795,N_1038);
and U6006 (N_6006,N_73,N_3566);
and U6007 (N_6007,N_2700,N_3657);
nand U6008 (N_6008,N_3674,N_585);
or U6009 (N_6009,N_2406,N_3245);
and U6010 (N_6010,N_2720,N_3262);
and U6011 (N_6011,N_1691,N_2035);
and U6012 (N_6012,N_338,N_255);
nand U6013 (N_6013,N_2155,N_3549);
or U6014 (N_6014,N_3194,N_3412);
xnor U6015 (N_6015,N_3379,N_302);
nand U6016 (N_6016,N_338,N_3271);
or U6017 (N_6017,N_2090,N_2639);
nand U6018 (N_6018,N_1022,N_1138);
nor U6019 (N_6019,N_97,N_579);
and U6020 (N_6020,N_3427,N_1293);
nand U6021 (N_6021,N_367,N_1109);
or U6022 (N_6022,N_962,N_684);
and U6023 (N_6023,N_1467,N_1213);
and U6024 (N_6024,N_3891,N_300);
and U6025 (N_6025,N_3972,N_2139);
and U6026 (N_6026,N_1767,N_501);
and U6027 (N_6027,N_3205,N_2674);
and U6028 (N_6028,N_373,N_160);
nand U6029 (N_6029,N_1744,N_3385);
and U6030 (N_6030,N_2262,N_3602);
or U6031 (N_6031,N_467,N_2584);
nand U6032 (N_6032,N_3559,N_99);
or U6033 (N_6033,N_1184,N_3505);
or U6034 (N_6034,N_3864,N_76);
and U6035 (N_6035,N_963,N_2233);
nand U6036 (N_6036,N_3940,N_1929);
or U6037 (N_6037,N_285,N_2323);
and U6038 (N_6038,N_1357,N_511);
nor U6039 (N_6039,N_2741,N_1916);
nor U6040 (N_6040,N_353,N_1767);
nor U6041 (N_6041,N_442,N_3548);
and U6042 (N_6042,N_835,N_172);
nor U6043 (N_6043,N_340,N_3335);
nand U6044 (N_6044,N_3265,N_3406);
or U6045 (N_6045,N_2777,N_2224);
and U6046 (N_6046,N_3139,N_2083);
nand U6047 (N_6047,N_2455,N_3050);
xor U6048 (N_6048,N_3546,N_3265);
nor U6049 (N_6049,N_3472,N_961);
nand U6050 (N_6050,N_203,N_2929);
nor U6051 (N_6051,N_3426,N_579);
or U6052 (N_6052,N_2059,N_2899);
nor U6053 (N_6053,N_214,N_759);
nand U6054 (N_6054,N_874,N_2734);
xnor U6055 (N_6055,N_282,N_2850);
nand U6056 (N_6056,N_506,N_2074);
nand U6057 (N_6057,N_3982,N_2379);
nor U6058 (N_6058,N_1457,N_3570);
nor U6059 (N_6059,N_2139,N_16);
and U6060 (N_6060,N_1997,N_1137);
nor U6061 (N_6061,N_2230,N_3816);
or U6062 (N_6062,N_2495,N_1550);
nor U6063 (N_6063,N_1612,N_2504);
nor U6064 (N_6064,N_1141,N_1401);
nand U6065 (N_6065,N_2780,N_2843);
nor U6066 (N_6066,N_2272,N_1761);
nand U6067 (N_6067,N_3538,N_1332);
nor U6068 (N_6068,N_3745,N_297);
nor U6069 (N_6069,N_1206,N_1634);
or U6070 (N_6070,N_2506,N_72);
or U6071 (N_6071,N_1292,N_286);
nor U6072 (N_6072,N_3954,N_1944);
nor U6073 (N_6073,N_3500,N_336);
nand U6074 (N_6074,N_884,N_939);
nand U6075 (N_6075,N_3576,N_3570);
and U6076 (N_6076,N_3005,N_2476);
nor U6077 (N_6077,N_2908,N_1919);
xnor U6078 (N_6078,N_652,N_2779);
and U6079 (N_6079,N_2502,N_2193);
nand U6080 (N_6080,N_1247,N_1828);
nand U6081 (N_6081,N_3687,N_2710);
nor U6082 (N_6082,N_2039,N_2636);
and U6083 (N_6083,N_3079,N_3119);
nor U6084 (N_6084,N_2210,N_3875);
nand U6085 (N_6085,N_2036,N_1260);
xnor U6086 (N_6086,N_3024,N_2210);
xnor U6087 (N_6087,N_71,N_2764);
nor U6088 (N_6088,N_3619,N_1245);
and U6089 (N_6089,N_2855,N_1917);
and U6090 (N_6090,N_3291,N_3524);
nand U6091 (N_6091,N_1419,N_784);
nor U6092 (N_6092,N_2664,N_1517);
nor U6093 (N_6093,N_676,N_380);
and U6094 (N_6094,N_259,N_954);
or U6095 (N_6095,N_1347,N_2298);
nor U6096 (N_6096,N_1258,N_1992);
or U6097 (N_6097,N_3435,N_3222);
xor U6098 (N_6098,N_596,N_604);
or U6099 (N_6099,N_614,N_2748);
nand U6100 (N_6100,N_58,N_3761);
xor U6101 (N_6101,N_3479,N_3262);
nor U6102 (N_6102,N_298,N_1016);
nand U6103 (N_6103,N_2897,N_3332);
or U6104 (N_6104,N_794,N_1566);
and U6105 (N_6105,N_3883,N_3152);
nor U6106 (N_6106,N_2099,N_3162);
and U6107 (N_6107,N_2111,N_2863);
or U6108 (N_6108,N_300,N_66);
or U6109 (N_6109,N_498,N_3153);
and U6110 (N_6110,N_3933,N_1088);
or U6111 (N_6111,N_2458,N_1397);
and U6112 (N_6112,N_1972,N_1729);
and U6113 (N_6113,N_527,N_2578);
nor U6114 (N_6114,N_658,N_2377);
nand U6115 (N_6115,N_3106,N_3005);
or U6116 (N_6116,N_403,N_1864);
nand U6117 (N_6117,N_2758,N_91);
or U6118 (N_6118,N_3359,N_3757);
nor U6119 (N_6119,N_3887,N_3853);
nor U6120 (N_6120,N_687,N_3291);
xor U6121 (N_6121,N_3624,N_2445);
nor U6122 (N_6122,N_3679,N_1717);
and U6123 (N_6123,N_3037,N_808);
or U6124 (N_6124,N_1816,N_2541);
nand U6125 (N_6125,N_537,N_2172);
xor U6126 (N_6126,N_3663,N_3212);
nand U6127 (N_6127,N_1874,N_3334);
or U6128 (N_6128,N_630,N_1673);
xnor U6129 (N_6129,N_349,N_652);
and U6130 (N_6130,N_2675,N_1998);
and U6131 (N_6131,N_2709,N_3850);
nor U6132 (N_6132,N_2646,N_2447);
nand U6133 (N_6133,N_2151,N_2728);
nor U6134 (N_6134,N_607,N_3488);
and U6135 (N_6135,N_1253,N_2918);
nand U6136 (N_6136,N_1954,N_1728);
or U6137 (N_6137,N_1035,N_3838);
and U6138 (N_6138,N_3649,N_59);
xnor U6139 (N_6139,N_601,N_3792);
or U6140 (N_6140,N_2875,N_3100);
or U6141 (N_6141,N_1260,N_3477);
nor U6142 (N_6142,N_886,N_3046);
nor U6143 (N_6143,N_849,N_2390);
or U6144 (N_6144,N_3312,N_730);
nor U6145 (N_6145,N_238,N_2799);
xor U6146 (N_6146,N_3719,N_502);
and U6147 (N_6147,N_2619,N_83);
or U6148 (N_6148,N_96,N_2501);
and U6149 (N_6149,N_1138,N_3757);
nand U6150 (N_6150,N_2510,N_388);
nor U6151 (N_6151,N_3429,N_2233);
and U6152 (N_6152,N_902,N_3660);
nand U6153 (N_6153,N_1441,N_672);
nor U6154 (N_6154,N_3623,N_690);
nand U6155 (N_6155,N_3305,N_3945);
nand U6156 (N_6156,N_1624,N_3939);
nor U6157 (N_6157,N_1912,N_1736);
nand U6158 (N_6158,N_109,N_1212);
and U6159 (N_6159,N_2048,N_1493);
xor U6160 (N_6160,N_3963,N_1114);
nor U6161 (N_6161,N_2011,N_2146);
or U6162 (N_6162,N_3727,N_1640);
or U6163 (N_6163,N_21,N_1233);
or U6164 (N_6164,N_1867,N_2243);
xor U6165 (N_6165,N_1364,N_200);
nor U6166 (N_6166,N_746,N_2307);
nor U6167 (N_6167,N_1787,N_3155);
or U6168 (N_6168,N_2452,N_2578);
or U6169 (N_6169,N_1146,N_942);
nand U6170 (N_6170,N_1617,N_3163);
xor U6171 (N_6171,N_2632,N_237);
nor U6172 (N_6172,N_2169,N_1613);
nand U6173 (N_6173,N_3999,N_1680);
nand U6174 (N_6174,N_3910,N_746);
nand U6175 (N_6175,N_1721,N_1718);
xor U6176 (N_6176,N_2873,N_3396);
or U6177 (N_6177,N_573,N_1082);
xor U6178 (N_6178,N_978,N_745);
nor U6179 (N_6179,N_3858,N_3083);
xor U6180 (N_6180,N_1910,N_3027);
and U6181 (N_6181,N_792,N_2870);
or U6182 (N_6182,N_1966,N_2765);
and U6183 (N_6183,N_714,N_871);
or U6184 (N_6184,N_1916,N_2420);
xor U6185 (N_6185,N_3799,N_3480);
nand U6186 (N_6186,N_2055,N_2376);
nand U6187 (N_6187,N_2522,N_2461);
or U6188 (N_6188,N_470,N_1076);
or U6189 (N_6189,N_1944,N_1015);
nor U6190 (N_6190,N_3866,N_218);
nand U6191 (N_6191,N_3848,N_1158);
or U6192 (N_6192,N_3971,N_2304);
and U6193 (N_6193,N_531,N_211);
nor U6194 (N_6194,N_3996,N_1036);
xor U6195 (N_6195,N_2010,N_3495);
and U6196 (N_6196,N_340,N_1574);
xnor U6197 (N_6197,N_1453,N_2973);
nor U6198 (N_6198,N_3858,N_276);
and U6199 (N_6199,N_2841,N_659);
nand U6200 (N_6200,N_1337,N_951);
nand U6201 (N_6201,N_448,N_1788);
nand U6202 (N_6202,N_780,N_2324);
nand U6203 (N_6203,N_3727,N_2036);
nand U6204 (N_6204,N_747,N_2013);
nand U6205 (N_6205,N_2665,N_1200);
or U6206 (N_6206,N_216,N_2486);
nor U6207 (N_6207,N_3613,N_814);
nand U6208 (N_6208,N_1200,N_696);
and U6209 (N_6209,N_3187,N_636);
or U6210 (N_6210,N_1502,N_3926);
nor U6211 (N_6211,N_2226,N_3818);
and U6212 (N_6212,N_3087,N_2928);
nand U6213 (N_6213,N_2992,N_317);
nand U6214 (N_6214,N_2969,N_3377);
nor U6215 (N_6215,N_1159,N_1293);
xor U6216 (N_6216,N_3305,N_3897);
or U6217 (N_6217,N_32,N_244);
or U6218 (N_6218,N_3020,N_775);
nand U6219 (N_6219,N_3651,N_955);
or U6220 (N_6220,N_2262,N_108);
and U6221 (N_6221,N_2631,N_1610);
nand U6222 (N_6222,N_3062,N_2509);
nand U6223 (N_6223,N_1922,N_1555);
nand U6224 (N_6224,N_65,N_1536);
or U6225 (N_6225,N_3738,N_191);
and U6226 (N_6226,N_3327,N_1);
nand U6227 (N_6227,N_2198,N_1102);
xor U6228 (N_6228,N_920,N_1450);
nand U6229 (N_6229,N_3299,N_2870);
and U6230 (N_6230,N_1958,N_2399);
nor U6231 (N_6231,N_3520,N_2254);
or U6232 (N_6232,N_2578,N_3419);
nor U6233 (N_6233,N_706,N_2490);
nand U6234 (N_6234,N_1657,N_3873);
nor U6235 (N_6235,N_1250,N_2771);
nand U6236 (N_6236,N_3828,N_2846);
or U6237 (N_6237,N_3645,N_2500);
nor U6238 (N_6238,N_2914,N_3865);
nand U6239 (N_6239,N_2614,N_1618);
xnor U6240 (N_6240,N_2816,N_48);
xnor U6241 (N_6241,N_2933,N_168);
and U6242 (N_6242,N_3316,N_792);
xor U6243 (N_6243,N_1470,N_3124);
and U6244 (N_6244,N_548,N_2320);
nor U6245 (N_6245,N_3796,N_3721);
or U6246 (N_6246,N_3182,N_3698);
nand U6247 (N_6247,N_989,N_294);
and U6248 (N_6248,N_2132,N_929);
or U6249 (N_6249,N_2154,N_2462);
or U6250 (N_6250,N_309,N_723);
nor U6251 (N_6251,N_2385,N_550);
nand U6252 (N_6252,N_3030,N_487);
or U6253 (N_6253,N_1185,N_63);
or U6254 (N_6254,N_2481,N_104);
nor U6255 (N_6255,N_2732,N_595);
nand U6256 (N_6256,N_209,N_3582);
or U6257 (N_6257,N_3846,N_1615);
xnor U6258 (N_6258,N_1247,N_264);
nor U6259 (N_6259,N_3261,N_1824);
xor U6260 (N_6260,N_1158,N_3487);
nor U6261 (N_6261,N_263,N_317);
nor U6262 (N_6262,N_3622,N_3242);
or U6263 (N_6263,N_1191,N_876);
nand U6264 (N_6264,N_3887,N_1591);
nor U6265 (N_6265,N_233,N_3724);
and U6266 (N_6266,N_2691,N_2934);
nand U6267 (N_6267,N_2441,N_1555);
nor U6268 (N_6268,N_2651,N_1809);
nand U6269 (N_6269,N_519,N_937);
nand U6270 (N_6270,N_2823,N_1256);
nand U6271 (N_6271,N_3246,N_2778);
or U6272 (N_6272,N_3825,N_1510);
or U6273 (N_6273,N_2024,N_3713);
nand U6274 (N_6274,N_3581,N_3392);
nand U6275 (N_6275,N_1940,N_1052);
nor U6276 (N_6276,N_2486,N_3369);
nor U6277 (N_6277,N_1513,N_2412);
or U6278 (N_6278,N_3361,N_2904);
xor U6279 (N_6279,N_2064,N_1328);
nor U6280 (N_6280,N_3703,N_1544);
nor U6281 (N_6281,N_1956,N_464);
nor U6282 (N_6282,N_3308,N_571);
nand U6283 (N_6283,N_3500,N_241);
or U6284 (N_6284,N_2920,N_3268);
nand U6285 (N_6285,N_2013,N_1667);
nand U6286 (N_6286,N_3036,N_304);
or U6287 (N_6287,N_721,N_2717);
or U6288 (N_6288,N_3508,N_2489);
nor U6289 (N_6289,N_1721,N_1086);
and U6290 (N_6290,N_255,N_1942);
and U6291 (N_6291,N_527,N_722);
xor U6292 (N_6292,N_1175,N_1947);
nand U6293 (N_6293,N_1740,N_2032);
nand U6294 (N_6294,N_2880,N_1437);
or U6295 (N_6295,N_3411,N_2753);
xor U6296 (N_6296,N_180,N_1107);
or U6297 (N_6297,N_1539,N_204);
nand U6298 (N_6298,N_2988,N_1930);
xnor U6299 (N_6299,N_3672,N_93);
xor U6300 (N_6300,N_3723,N_1503);
or U6301 (N_6301,N_2132,N_2225);
and U6302 (N_6302,N_3815,N_2621);
and U6303 (N_6303,N_3515,N_2956);
and U6304 (N_6304,N_2542,N_2136);
and U6305 (N_6305,N_759,N_2034);
nor U6306 (N_6306,N_1945,N_2061);
and U6307 (N_6307,N_216,N_2285);
or U6308 (N_6308,N_2900,N_258);
nand U6309 (N_6309,N_3615,N_2647);
nor U6310 (N_6310,N_388,N_1023);
nor U6311 (N_6311,N_487,N_2642);
or U6312 (N_6312,N_2619,N_2606);
nand U6313 (N_6313,N_926,N_2965);
or U6314 (N_6314,N_3776,N_2356);
xnor U6315 (N_6315,N_3665,N_1648);
nand U6316 (N_6316,N_2398,N_2436);
nor U6317 (N_6317,N_1836,N_3186);
and U6318 (N_6318,N_2720,N_1715);
nor U6319 (N_6319,N_2083,N_3735);
and U6320 (N_6320,N_522,N_2742);
and U6321 (N_6321,N_1312,N_932);
xor U6322 (N_6322,N_2261,N_302);
nor U6323 (N_6323,N_2492,N_1206);
or U6324 (N_6324,N_3034,N_3387);
and U6325 (N_6325,N_3995,N_3498);
xnor U6326 (N_6326,N_2764,N_2246);
nor U6327 (N_6327,N_2839,N_653);
nand U6328 (N_6328,N_1909,N_551);
nand U6329 (N_6329,N_1199,N_2037);
nand U6330 (N_6330,N_3014,N_3553);
and U6331 (N_6331,N_1358,N_2671);
or U6332 (N_6332,N_2480,N_2942);
nand U6333 (N_6333,N_2632,N_1503);
and U6334 (N_6334,N_2346,N_1147);
nor U6335 (N_6335,N_2301,N_3873);
nand U6336 (N_6336,N_1100,N_1306);
or U6337 (N_6337,N_1890,N_1894);
nand U6338 (N_6338,N_3257,N_561);
nor U6339 (N_6339,N_2641,N_2185);
or U6340 (N_6340,N_3324,N_214);
or U6341 (N_6341,N_2625,N_73);
xnor U6342 (N_6342,N_1599,N_1375);
or U6343 (N_6343,N_1690,N_559);
nand U6344 (N_6344,N_1497,N_1039);
nand U6345 (N_6345,N_2138,N_1058);
or U6346 (N_6346,N_2389,N_2922);
nand U6347 (N_6347,N_1719,N_3401);
nand U6348 (N_6348,N_3588,N_3022);
and U6349 (N_6349,N_1442,N_3514);
and U6350 (N_6350,N_1369,N_515);
and U6351 (N_6351,N_2044,N_2904);
nand U6352 (N_6352,N_2758,N_3164);
or U6353 (N_6353,N_844,N_1439);
nor U6354 (N_6354,N_2024,N_678);
nand U6355 (N_6355,N_2934,N_644);
and U6356 (N_6356,N_1329,N_1019);
nand U6357 (N_6357,N_3633,N_3738);
or U6358 (N_6358,N_3111,N_995);
nor U6359 (N_6359,N_591,N_3044);
nor U6360 (N_6360,N_3561,N_2727);
and U6361 (N_6361,N_3978,N_2366);
nand U6362 (N_6362,N_1579,N_2628);
nand U6363 (N_6363,N_1838,N_2982);
nor U6364 (N_6364,N_1761,N_245);
and U6365 (N_6365,N_1440,N_1566);
nand U6366 (N_6366,N_794,N_1162);
and U6367 (N_6367,N_3203,N_3589);
nor U6368 (N_6368,N_3858,N_1028);
or U6369 (N_6369,N_3081,N_959);
and U6370 (N_6370,N_1568,N_1606);
xnor U6371 (N_6371,N_3869,N_3642);
nand U6372 (N_6372,N_2719,N_1900);
nor U6373 (N_6373,N_3751,N_1840);
nor U6374 (N_6374,N_642,N_1020);
or U6375 (N_6375,N_3678,N_824);
or U6376 (N_6376,N_3940,N_2466);
or U6377 (N_6377,N_200,N_1553);
and U6378 (N_6378,N_1017,N_3296);
nor U6379 (N_6379,N_2155,N_1910);
and U6380 (N_6380,N_2766,N_3859);
nor U6381 (N_6381,N_1669,N_2259);
xnor U6382 (N_6382,N_167,N_3347);
nor U6383 (N_6383,N_3050,N_3647);
nand U6384 (N_6384,N_3427,N_3487);
nand U6385 (N_6385,N_2287,N_2173);
and U6386 (N_6386,N_3924,N_438);
nor U6387 (N_6387,N_2480,N_1459);
or U6388 (N_6388,N_1366,N_592);
or U6389 (N_6389,N_1787,N_1444);
nor U6390 (N_6390,N_3911,N_2685);
and U6391 (N_6391,N_1359,N_2407);
nand U6392 (N_6392,N_903,N_3565);
and U6393 (N_6393,N_1093,N_1169);
and U6394 (N_6394,N_3091,N_2963);
or U6395 (N_6395,N_178,N_2525);
or U6396 (N_6396,N_65,N_3747);
nand U6397 (N_6397,N_3626,N_978);
and U6398 (N_6398,N_2865,N_722);
and U6399 (N_6399,N_781,N_2918);
or U6400 (N_6400,N_2057,N_1515);
nor U6401 (N_6401,N_2878,N_53);
or U6402 (N_6402,N_1426,N_2475);
or U6403 (N_6403,N_2347,N_2518);
and U6404 (N_6404,N_1471,N_2114);
nand U6405 (N_6405,N_816,N_2173);
and U6406 (N_6406,N_1131,N_3252);
xor U6407 (N_6407,N_1102,N_2435);
xnor U6408 (N_6408,N_2116,N_118);
and U6409 (N_6409,N_788,N_2819);
nor U6410 (N_6410,N_3457,N_1187);
nor U6411 (N_6411,N_1498,N_2983);
nor U6412 (N_6412,N_146,N_2818);
nand U6413 (N_6413,N_3125,N_3142);
or U6414 (N_6414,N_937,N_723);
xnor U6415 (N_6415,N_1925,N_2964);
or U6416 (N_6416,N_644,N_3027);
xor U6417 (N_6417,N_3921,N_3317);
or U6418 (N_6418,N_2775,N_1312);
or U6419 (N_6419,N_319,N_3131);
and U6420 (N_6420,N_3754,N_3392);
xor U6421 (N_6421,N_3554,N_1424);
nand U6422 (N_6422,N_2624,N_3240);
nand U6423 (N_6423,N_3874,N_886);
nand U6424 (N_6424,N_1617,N_1780);
or U6425 (N_6425,N_435,N_3708);
or U6426 (N_6426,N_3050,N_3843);
nor U6427 (N_6427,N_364,N_3037);
or U6428 (N_6428,N_1307,N_319);
and U6429 (N_6429,N_1328,N_191);
and U6430 (N_6430,N_2269,N_554);
nor U6431 (N_6431,N_2060,N_3900);
nor U6432 (N_6432,N_1559,N_1511);
xnor U6433 (N_6433,N_1336,N_187);
and U6434 (N_6434,N_3303,N_3627);
nand U6435 (N_6435,N_99,N_2763);
or U6436 (N_6436,N_3963,N_2498);
nand U6437 (N_6437,N_898,N_800);
nor U6438 (N_6438,N_875,N_3922);
and U6439 (N_6439,N_2098,N_884);
or U6440 (N_6440,N_1469,N_1916);
nand U6441 (N_6441,N_2316,N_684);
and U6442 (N_6442,N_1765,N_2003);
and U6443 (N_6443,N_3530,N_571);
or U6444 (N_6444,N_3345,N_1354);
nor U6445 (N_6445,N_2137,N_3281);
or U6446 (N_6446,N_1862,N_2227);
nor U6447 (N_6447,N_3282,N_244);
and U6448 (N_6448,N_1569,N_1386);
nor U6449 (N_6449,N_2346,N_1629);
and U6450 (N_6450,N_2276,N_2215);
and U6451 (N_6451,N_18,N_1658);
and U6452 (N_6452,N_3895,N_2623);
or U6453 (N_6453,N_2920,N_965);
nand U6454 (N_6454,N_3723,N_2940);
or U6455 (N_6455,N_983,N_1943);
nor U6456 (N_6456,N_3921,N_2614);
or U6457 (N_6457,N_2976,N_408);
and U6458 (N_6458,N_2385,N_1516);
or U6459 (N_6459,N_3392,N_1315);
or U6460 (N_6460,N_2446,N_2888);
nor U6461 (N_6461,N_305,N_3451);
and U6462 (N_6462,N_3695,N_1985);
and U6463 (N_6463,N_1252,N_36);
and U6464 (N_6464,N_1483,N_1348);
or U6465 (N_6465,N_3988,N_2211);
nand U6466 (N_6466,N_239,N_2430);
and U6467 (N_6467,N_3003,N_3961);
nand U6468 (N_6468,N_1126,N_3731);
or U6469 (N_6469,N_1349,N_1425);
and U6470 (N_6470,N_2555,N_1825);
or U6471 (N_6471,N_2740,N_716);
nor U6472 (N_6472,N_60,N_394);
xor U6473 (N_6473,N_2476,N_429);
and U6474 (N_6474,N_2731,N_7);
or U6475 (N_6475,N_1445,N_1070);
nand U6476 (N_6476,N_2427,N_3339);
nor U6477 (N_6477,N_773,N_1965);
nor U6478 (N_6478,N_33,N_1038);
nand U6479 (N_6479,N_980,N_1337);
nand U6480 (N_6480,N_2212,N_2186);
nor U6481 (N_6481,N_2696,N_2243);
or U6482 (N_6482,N_1331,N_2342);
and U6483 (N_6483,N_3209,N_825);
and U6484 (N_6484,N_1004,N_2377);
and U6485 (N_6485,N_310,N_2235);
nand U6486 (N_6486,N_3290,N_3830);
nand U6487 (N_6487,N_520,N_2123);
xor U6488 (N_6488,N_207,N_2222);
nand U6489 (N_6489,N_2896,N_1439);
or U6490 (N_6490,N_2840,N_2852);
xnor U6491 (N_6491,N_2764,N_1033);
nor U6492 (N_6492,N_201,N_641);
and U6493 (N_6493,N_336,N_2471);
and U6494 (N_6494,N_2963,N_3916);
nand U6495 (N_6495,N_2110,N_3559);
nor U6496 (N_6496,N_1096,N_1117);
and U6497 (N_6497,N_1564,N_1875);
and U6498 (N_6498,N_612,N_607);
nand U6499 (N_6499,N_60,N_1478);
or U6500 (N_6500,N_337,N_1095);
and U6501 (N_6501,N_3872,N_3283);
and U6502 (N_6502,N_2625,N_452);
xor U6503 (N_6503,N_1773,N_2377);
and U6504 (N_6504,N_1533,N_3215);
nand U6505 (N_6505,N_2752,N_259);
nand U6506 (N_6506,N_392,N_1422);
nand U6507 (N_6507,N_3574,N_1180);
nor U6508 (N_6508,N_3350,N_1159);
nor U6509 (N_6509,N_2624,N_3150);
nor U6510 (N_6510,N_1502,N_2806);
xor U6511 (N_6511,N_2013,N_2020);
nor U6512 (N_6512,N_1542,N_3252);
nor U6513 (N_6513,N_1853,N_123);
or U6514 (N_6514,N_1685,N_3181);
and U6515 (N_6515,N_1336,N_3123);
nor U6516 (N_6516,N_2724,N_2638);
or U6517 (N_6517,N_2098,N_962);
and U6518 (N_6518,N_3021,N_3020);
or U6519 (N_6519,N_1854,N_2661);
nand U6520 (N_6520,N_2478,N_931);
or U6521 (N_6521,N_2268,N_892);
nor U6522 (N_6522,N_1401,N_1424);
nand U6523 (N_6523,N_1410,N_2627);
or U6524 (N_6524,N_3064,N_382);
or U6525 (N_6525,N_2434,N_2887);
or U6526 (N_6526,N_2742,N_1559);
nand U6527 (N_6527,N_3897,N_1737);
and U6528 (N_6528,N_872,N_3891);
or U6529 (N_6529,N_2489,N_3745);
or U6530 (N_6530,N_920,N_364);
nor U6531 (N_6531,N_3543,N_2163);
and U6532 (N_6532,N_3928,N_2545);
xor U6533 (N_6533,N_516,N_2857);
nand U6534 (N_6534,N_167,N_1108);
nor U6535 (N_6535,N_338,N_3255);
or U6536 (N_6536,N_3291,N_2306);
and U6537 (N_6537,N_2859,N_2086);
and U6538 (N_6538,N_3375,N_2413);
nor U6539 (N_6539,N_3954,N_3710);
nor U6540 (N_6540,N_1521,N_3295);
or U6541 (N_6541,N_1240,N_966);
nand U6542 (N_6542,N_411,N_92);
or U6543 (N_6543,N_822,N_3665);
xor U6544 (N_6544,N_891,N_2882);
nand U6545 (N_6545,N_2457,N_3714);
nor U6546 (N_6546,N_70,N_3923);
and U6547 (N_6547,N_2579,N_1864);
nor U6548 (N_6548,N_3119,N_3186);
or U6549 (N_6549,N_888,N_1192);
nor U6550 (N_6550,N_1036,N_970);
nor U6551 (N_6551,N_1153,N_2193);
nor U6552 (N_6552,N_2424,N_2344);
and U6553 (N_6553,N_703,N_1340);
nor U6554 (N_6554,N_2921,N_3185);
nor U6555 (N_6555,N_1629,N_1886);
xnor U6556 (N_6556,N_1490,N_1262);
xnor U6557 (N_6557,N_443,N_2158);
nand U6558 (N_6558,N_3708,N_1236);
or U6559 (N_6559,N_1984,N_2280);
nor U6560 (N_6560,N_261,N_1342);
and U6561 (N_6561,N_2189,N_2990);
or U6562 (N_6562,N_1753,N_3003);
xor U6563 (N_6563,N_2345,N_12);
or U6564 (N_6564,N_3897,N_1389);
nand U6565 (N_6565,N_1821,N_1379);
and U6566 (N_6566,N_953,N_3183);
nor U6567 (N_6567,N_52,N_2206);
and U6568 (N_6568,N_3605,N_3595);
or U6569 (N_6569,N_3974,N_700);
nand U6570 (N_6570,N_2251,N_1131);
xnor U6571 (N_6571,N_1739,N_3835);
or U6572 (N_6572,N_1255,N_2414);
nor U6573 (N_6573,N_2889,N_1805);
or U6574 (N_6574,N_2827,N_343);
nand U6575 (N_6575,N_1240,N_3919);
or U6576 (N_6576,N_1324,N_1402);
or U6577 (N_6577,N_3118,N_2699);
nand U6578 (N_6578,N_617,N_3498);
and U6579 (N_6579,N_953,N_1414);
nand U6580 (N_6580,N_2993,N_3006);
nor U6581 (N_6581,N_3944,N_3927);
nand U6582 (N_6582,N_3733,N_697);
nand U6583 (N_6583,N_91,N_7);
nand U6584 (N_6584,N_566,N_3560);
xor U6585 (N_6585,N_227,N_1633);
nand U6586 (N_6586,N_600,N_1562);
nand U6587 (N_6587,N_506,N_2416);
nor U6588 (N_6588,N_1719,N_708);
nor U6589 (N_6589,N_3286,N_589);
nor U6590 (N_6590,N_214,N_913);
nor U6591 (N_6591,N_1294,N_2658);
nor U6592 (N_6592,N_3690,N_7);
or U6593 (N_6593,N_835,N_954);
nand U6594 (N_6594,N_1523,N_1877);
or U6595 (N_6595,N_2050,N_2250);
nor U6596 (N_6596,N_2155,N_2563);
nor U6597 (N_6597,N_3164,N_960);
or U6598 (N_6598,N_874,N_869);
or U6599 (N_6599,N_634,N_3724);
and U6600 (N_6600,N_3700,N_328);
xor U6601 (N_6601,N_1643,N_1054);
nand U6602 (N_6602,N_3695,N_1016);
or U6603 (N_6603,N_2166,N_2034);
nor U6604 (N_6604,N_1470,N_150);
nor U6605 (N_6605,N_2731,N_3519);
nor U6606 (N_6606,N_1893,N_3518);
nand U6607 (N_6607,N_1295,N_1323);
xnor U6608 (N_6608,N_2943,N_2465);
and U6609 (N_6609,N_598,N_878);
nor U6610 (N_6610,N_3026,N_3038);
and U6611 (N_6611,N_3150,N_1219);
xnor U6612 (N_6612,N_3265,N_330);
or U6613 (N_6613,N_200,N_399);
xor U6614 (N_6614,N_2146,N_903);
or U6615 (N_6615,N_1694,N_1473);
or U6616 (N_6616,N_940,N_1424);
nand U6617 (N_6617,N_13,N_835);
and U6618 (N_6618,N_1284,N_3752);
or U6619 (N_6619,N_1534,N_3360);
and U6620 (N_6620,N_794,N_2890);
and U6621 (N_6621,N_260,N_1609);
xor U6622 (N_6622,N_2717,N_2455);
and U6623 (N_6623,N_1715,N_3595);
nand U6624 (N_6624,N_1535,N_2691);
nor U6625 (N_6625,N_2173,N_873);
nand U6626 (N_6626,N_2851,N_2648);
nand U6627 (N_6627,N_1450,N_2406);
or U6628 (N_6628,N_2796,N_65);
nor U6629 (N_6629,N_2935,N_2643);
nor U6630 (N_6630,N_2650,N_1399);
or U6631 (N_6631,N_2371,N_1437);
nand U6632 (N_6632,N_2202,N_241);
nor U6633 (N_6633,N_1125,N_3398);
or U6634 (N_6634,N_797,N_1560);
and U6635 (N_6635,N_432,N_673);
nor U6636 (N_6636,N_1148,N_1078);
nand U6637 (N_6637,N_1986,N_1247);
nand U6638 (N_6638,N_2396,N_1592);
or U6639 (N_6639,N_3121,N_1826);
and U6640 (N_6640,N_3999,N_1612);
nor U6641 (N_6641,N_3141,N_2523);
nand U6642 (N_6642,N_2010,N_958);
nand U6643 (N_6643,N_1937,N_3430);
nand U6644 (N_6644,N_2558,N_3038);
nor U6645 (N_6645,N_1003,N_3379);
nor U6646 (N_6646,N_3195,N_2838);
nand U6647 (N_6647,N_3922,N_2586);
and U6648 (N_6648,N_1431,N_548);
nand U6649 (N_6649,N_2994,N_1146);
nand U6650 (N_6650,N_3716,N_2266);
nand U6651 (N_6651,N_1979,N_272);
nand U6652 (N_6652,N_2605,N_1620);
nand U6653 (N_6653,N_543,N_3359);
nor U6654 (N_6654,N_632,N_423);
and U6655 (N_6655,N_1532,N_1720);
nor U6656 (N_6656,N_1308,N_959);
or U6657 (N_6657,N_3340,N_1230);
nand U6658 (N_6658,N_964,N_1463);
or U6659 (N_6659,N_2642,N_1292);
nand U6660 (N_6660,N_2201,N_737);
nand U6661 (N_6661,N_2815,N_3181);
nor U6662 (N_6662,N_1925,N_1725);
or U6663 (N_6663,N_1452,N_1361);
nand U6664 (N_6664,N_3383,N_1185);
nand U6665 (N_6665,N_1966,N_486);
nand U6666 (N_6666,N_3116,N_508);
xor U6667 (N_6667,N_2306,N_3968);
nor U6668 (N_6668,N_813,N_2828);
and U6669 (N_6669,N_2381,N_455);
nor U6670 (N_6670,N_3290,N_2007);
nand U6671 (N_6671,N_2726,N_3170);
or U6672 (N_6672,N_3331,N_1515);
nand U6673 (N_6673,N_1050,N_2689);
or U6674 (N_6674,N_1225,N_1523);
or U6675 (N_6675,N_2136,N_1433);
and U6676 (N_6676,N_714,N_1659);
nor U6677 (N_6677,N_2141,N_1735);
xnor U6678 (N_6678,N_2522,N_2690);
or U6679 (N_6679,N_1037,N_88);
nand U6680 (N_6680,N_94,N_3381);
or U6681 (N_6681,N_3116,N_3363);
nor U6682 (N_6682,N_464,N_2719);
xor U6683 (N_6683,N_2730,N_3521);
nand U6684 (N_6684,N_3749,N_3316);
and U6685 (N_6685,N_730,N_882);
nor U6686 (N_6686,N_1381,N_3683);
or U6687 (N_6687,N_643,N_485);
or U6688 (N_6688,N_3331,N_1880);
nor U6689 (N_6689,N_1200,N_749);
nor U6690 (N_6690,N_2561,N_1224);
and U6691 (N_6691,N_2882,N_3891);
or U6692 (N_6692,N_231,N_2549);
nand U6693 (N_6693,N_2775,N_480);
and U6694 (N_6694,N_3409,N_3519);
nand U6695 (N_6695,N_1754,N_2543);
nor U6696 (N_6696,N_1391,N_2464);
and U6697 (N_6697,N_2872,N_1057);
nor U6698 (N_6698,N_1258,N_3589);
nand U6699 (N_6699,N_3800,N_2151);
or U6700 (N_6700,N_1244,N_721);
nand U6701 (N_6701,N_38,N_2405);
nand U6702 (N_6702,N_2231,N_1605);
nand U6703 (N_6703,N_2717,N_651);
and U6704 (N_6704,N_881,N_2783);
nor U6705 (N_6705,N_1642,N_1442);
or U6706 (N_6706,N_1785,N_1144);
and U6707 (N_6707,N_256,N_3577);
and U6708 (N_6708,N_2359,N_1357);
or U6709 (N_6709,N_564,N_3517);
xor U6710 (N_6710,N_1604,N_3910);
xnor U6711 (N_6711,N_3558,N_1898);
or U6712 (N_6712,N_3763,N_3452);
nand U6713 (N_6713,N_1217,N_2739);
nor U6714 (N_6714,N_1298,N_1684);
nand U6715 (N_6715,N_94,N_538);
xnor U6716 (N_6716,N_1825,N_2853);
nor U6717 (N_6717,N_3567,N_327);
nor U6718 (N_6718,N_1329,N_997);
nor U6719 (N_6719,N_3842,N_3444);
nor U6720 (N_6720,N_2837,N_3906);
nand U6721 (N_6721,N_3863,N_12);
nand U6722 (N_6722,N_2518,N_1732);
nor U6723 (N_6723,N_3242,N_507);
or U6724 (N_6724,N_2408,N_2076);
nor U6725 (N_6725,N_3759,N_1691);
and U6726 (N_6726,N_2443,N_1880);
and U6727 (N_6727,N_1401,N_1156);
or U6728 (N_6728,N_3392,N_1066);
and U6729 (N_6729,N_959,N_3015);
and U6730 (N_6730,N_1496,N_2011);
and U6731 (N_6731,N_3593,N_2836);
or U6732 (N_6732,N_1330,N_1336);
nor U6733 (N_6733,N_1776,N_3689);
xnor U6734 (N_6734,N_74,N_293);
nand U6735 (N_6735,N_2725,N_353);
nand U6736 (N_6736,N_934,N_3399);
nor U6737 (N_6737,N_376,N_852);
and U6738 (N_6738,N_723,N_3456);
nand U6739 (N_6739,N_1215,N_960);
and U6740 (N_6740,N_62,N_2415);
nor U6741 (N_6741,N_2666,N_699);
nor U6742 (N_6742,N_3053,N_423);
nand U6743 (N_6743,N_3214,N_2025);
and U6744 (N_6744,N_3996,N_562);
or U6745 (N_6745,N_2052,N_3856);
nor U6746 (N_6746,N_3807,N_3554);
and U6747 (N_6747,N_2473,N_2426);
nand U6748 (N_6748,N_3988,N_3600);
and U6749 (N_6749,N_849,N_1396);
or U6750 (N_6750,N_601,N_2288);
nand U6751 (N_6751,N_966,N_1199);
or U6752 (N_6752,N_3395,N_3599);
and U6753 (N_6753,N_1864,N_3778);
or U6754 (N_6754,N_2277,N_3493);
xnor U6755 (N_6755,N_2627,N_2715);
and U6756 (N_6756,N_3966,N_1643);
nor U6757 (N_6757,N_1847,N_3939);
nor U6758 (N_6758,N_1544,N_1068);
or U6759 (N_6759,N_2975,N_3575);
or U6760 (N_6760,N_3041,N_1170);
nor U6761 (N_6761,N_1678,N_3285);
nor U6762 (N_6762,N_1467,N_334);
xor U6763 (N_6763,N_374,N_3192);
and U6764 (N_6764,N_119,N_1998);
and U6765 (N_6765,N_2460,N_3998);
and U6766 (N_6766,N_3921,N_3455);
nand U6767 (N_6767,N_2461,N_3333);
or U6768 (N_6768,N_2868,N_2350);
nand U6769 (N_6769,N_1393,N_964);
and U6770 (N_6770,N_850,N_1506);
and U6771 (N_6771,N_928,N_2441);
and U6772 (N_6772,N_690,N_614);
nor U6773 (N_6773,N_1593,N_3061);
and U6774 (N_6774,N_1858,N_894);
and U6775 (N_6775,N_3818,N_2779);
nor U6776 (N_6776,N_1936,N_2815);
nor U6777 (N_6777,N_1875,N_636);
nor U6778 (N_6778,N_875,N_3771);
and U6779 (N_6779,N_2499,N_998);
xnor U6780 (N_6780,N_2172,N_2042);
nand U6781 (N_6781,N_2818,N_2271);
or U6782 (N_6782,N_3420,N_1074);
xor U6783 (N_6783,N_722,N_3430);
nor U6784 (N_6784,N_2988,N_3302);
or U6785 (N_6785,N_1352,N_557);
and U6786 (N_6786,N_3463,N_1972);
nand U6787 (N_6787,N_3188,N_2348);
and U6788 (N_6788,N_1054,N_3569);
nor U6789 (N_6789,N_432,N_2523);
nor U6790 (N_6790,N_3071,N_3504);
nor U6791 (N_6791,N_3276,N_1554);
or U6792 (N_6792,N_1977,N_3742);
or U6793 (N_6793,N_3203,N_107);
nand U6794 (N_6794,N_40,N_3325);
or U6795 (N_6795,N_3557,N_2960);
nand U6796 (N_6796,N_744,N_1996);
and U6797 (N_6797,N_3249,N_1144);
and U6798 (N_6798,N_2399,N_1308);
or U6799 (N_6799,N_3061,N_1837);
or U6800 (N_6800,N_2584,N_2904);
nor U6801 (N_6801,N_3214,N_3938);
and U6802 (N_6802,N_2203,N_1793);
or U6803 (N_6803,N_1019,N_2282);
or U6804 (N_6804,N_2329,N_1212);
or U6805 (N_6805,N_711,N_2702);
and U6806 (N_6806,N_3447,N_931);
xor U6807 (N_6807,N_3375,N_3954);
or U6808 (N_6808,N_2517,N_523);
and U6809 (N_6809,N_1034,N_2993);
or U6810 (N_6810,N_2304,N_1374);
nand U6811 (N_6811,N_2420,N_1937);
nor U6812 (N_6812,N_1904,N_1649);
and U6813 (N_6813,N_3201,N_2553);
nand U6814 (N_6814,N_3904,N_1177);
or U6815 (N_6815,N_1623,N_3023);
xor U6816 (N_6816,N_2741,N_2324);
and U6817 (N_6817,N_1637,N_1428);
nand U6818 (N_6818,N_2872,N_222);
nor U6819 (N_6819,N_2050,N_3981);
nand U6820 (N_6820,N_2112,N_2302);
or U6821 (N_6821,N_1503,N_3583);
and U6822 (N_6822,N_393,N_935);
nand U6823 (N_6823,N_1731,N_699);
nand U6824 (N_6824,N_1264,N_3039);
or U6825 (N_6825,N_2680,N_2165);
xor U6826 (N_6826,N_665,N_2341);
or U6827 (N_6827,N_854,N_1678);
or U6828 (N_6828,N_372,N_1687);
xor U6829 (N_6829,N_752,N_947);
or U6830 (N_6830,N_702,N_1608);
or U6831 (N_6831,N_3560,N_690);
or U6832 (N_6832,N_2317,N_1603);
nor U6833 (N_6833,N_2837,N_2316);
or U6834 (N_6834,N_3300,N_1894);
nor U6835 (N_6835,N_2921,N_995);
or U6836 (N_6836,N_2243,N_3079);
nor U6837 (N_6837,N_3088,N_3841);
nor U6838 (N_6838,N_938,N_3497);
and U6839 (N_6839,N_2276,N_3607);
nor U6840 (N_6840,N_1444,N_1763);
xor U6841 (N_6841,N_2782,N_1841);
and U6842 (N_6842,N_3425,N_1415);
or U6843 (N_6843,N_3063,N_3601);
nor U6844 (N_6844,N_1000,N_1260);
nand U6845 (N_6845,N_2831,N_1427);
nor U6846 (N_6846,N_3475,N_693);
nor U6847 (N_6847,N_1080,N_156);
nand U6848 (N_6848,N_2258,N_739);
and U6849 (N_6849,N_3863,N_109);
nand U6850 (N_6850,N_3077,N_3912);
xnor U6851 (N_6851,N_900,N_1668);
or U6852 (N_6852,N_361,N_3136);
nand U6853 (N_6853,N_706,N_1142);
nor U6854 (N_6854,N_809,N_3138);
and U6855 (N_6855,N_888,N_199);
nand U6856 (N_6856,N_2457,N_1538);
nor U6857 (N_6857,N_366,N_77);
or U6858 (N_6858,N_483,N_751);
and U6859 (N_6859,N_2056,N_2588);
or U6860 (N_6860,N_3554,N_2209);
nor U6861 (N_6861,N_1178,N_3979);
nor U6862 (N_6862,N_76,N_2235);
and U6863 (N_6863,N_935,N_3225);
nand U6864 (N_6864,N_1160,N_3022);
or U6865 (N_6865,N_3865,N_415);
or U6866 (N_6866,N_458,N_775);
xor U6867 (N_6867,N_3621,N_2832);
nor U6868 (N_6868,N_3655,N_1176);
nand U6869 (N_6869,N_3668,N_2696);
and U6870 (N_6870,N_3695,N_99);
and U6871 (N_6871,N_1778,N_2776);
nor U6872 (N_6872,N_3160,N_3445);
nand U6873 (N_6873,N_314,N_211);
and U6874 (N_6874,N_185,N_443);
nand U6875 (N_6875,N_3704,N_2638);
and U6876 (N_6876,N_2897,N_2096);
or U6877 (N_6877,N_3212,N_1350);
nor U6878 (N_6878,N_1761,N_3390);
nand U6879 (N_6879,N_170,N_3591);
xor U6880 (N_6880,N_405,N_846);
or U6881 (N_6881,N_452,N_124);
or U6882 (N_6882,N_1690,N_1357);
nor U6883 (N_6883,N_1519,N_163);
xnor U6884 (N_6884,N_2004,N_51);
and U6885 (N_6885,N_336,N_350);
and U6886 (N_6886,N_1323,N_1794);
nor U6887 (N_6887,N_2200,N_2852);
or U6888 (N_6888,N_3241,N_2269);
and U6889 (N_6889,N_3798,N_2676);
nor U6890 (N_6890,N_349,N_2390);
or U6891 (N_6891,N_3755,N_926);
nand U6892 (N_6892,N_3338,N_2065);
and U6893 (N_6893,N_1687,N_154);
and U6894 (N_6894,N_2080,N_3791);
and U6895 (N_6895,N_3166,N_2869);
xor U6896 (N_6896,N_3100,N_2771);
or U6897 (N_6897,N_896,N_3056);
or U6898 (N_6898,N_980,N_3857);
nor U6899 (N_6899,N_2268,N_250);
or U6900 (N_6900,N_1027,N_3173);
nand U6901 (N_6901,N_652,N_1066);
nor U6902 (N_6902,N_3615,N_3060);
nor U6903 (N_6903,N_785,N_3990);
and U6904 (N_6904,N_1411,N_1833);
nand U6905 (N_6905,N_1076,N_480);
nor U6906 (N_6906,N_3556,N_573);
nor U6907 (N_6907,N_31,N_455);
or U6908 (N_6908,N_2366,N_1032);
or U6909 (N_6909,N_138,N_153);
nand U6910 (N_6910,N_434,N_1420);
nor U6911 (N_6911,N_3030,N_2869);
xnor U6912 (N_6912,N_406,N_3686);
or U6913 (N_6913,N_3668,N_1054);
and U6914 (N_6914,N_2102,N_737);
xor U6915 (N_6915,N_452,N_3407);
nand U6916 (N_6916,N_2181,N_3860);
xnor U6917 (N_6917,N_2421,N_3431);
and U6918 (N_6918,N_2271,N_2904);
nor U6919 (N_6919,N_2564,N_460);
and U6920 (N_6920,N_835,N_2039);
and U6921 (N_6921,N_3422,N_827);
nor U6922 (N_6922,N_2709,N_86);
nand U6923 (N_6923,N_3844,N_1680);
or U6924 (N_6924,N_3573,N_1276);
xnor U6925 (N_6925,N_952,N_2414);
xnor U6926 (N_6926,N_3792,N_193);
nor U6927 (N_6927,N_3068,N_3617);
nor U6928 (N_6928,N_2471,N_3421);
nor U6929 (N_6929,N_3655,N_781);
and U6930 (N_6930,N_2119,N_1923);
nand U6931 (N_6931,N_3693,N_673);
nand U6932 (N_6932,N_2759,N_3814);
xor U6933 (N_6933,N_3602,N_2976);
nor U6934 (N_6934,N_867,N_438);
nand U6935 (N_6935,N_2502,N_2631);
nor U6936 (N_6936,N_3264,N_104);
or U6937 (N_6937,N_6,N_2068);
and U6938 (N_6938,N_321,N_2190);
nand U6939 (N_6939,N_3523,N_7);
nor U6940 (N_6940,N_712,N_1265);
nor U6941 (N_6941,N_2131,N_413);
or U6942 (N_6942,N_491,N_714);
nand U6943 (N_6943,N_3753,N_1524);
or U6944 (N_6944,N_2196,N_169);
or U6945 (N_6945,N_3420,N_3423);
and U6946 (N_6946,N_2813,N_345);
or U6947 (N_6947,N_1362,N_3707);
and U6948 (N_6948,N_964,N_3624);
nor U6949 (N_6949,N_249,N_1742);
nor U6950 (N_6950,N_865,N_1937);
or U6951 (N_6951,N_3808,N_2964);
nand U6952 (N_6952,N_3414,N_1945);
or U6953 (N_6953,N_887,N_1809);
or U6954 (N_6954,N_3603,N_718);
or U6955 (N_6955,N_823,N_854);
or U6956 (N_6956,N_1293,N_3187);
and U6957 (N_6957,N_2893,N_2085);
and U6958 (N_6958,N_2477,N_1485);
and U6959 (N_6959,N_2344,N_1233);
and U6960 (N_6960,N_2714,N_1262);
xor U6961 (N_6961,N_3359,N_3373);
or U6962 (N_6962,N_3353,N_2983);
nor U6963 (N_6963,N_2218,N_2003);
or U6964 (N_6964,N_603,N_431);
or U6965 (N_6965,N_1280,N_994);
nand U6966 (N_6966,N_2917,N_3131);
or U6967 (N_6967,N_2873,N_1187);
nor U6968 (N_6968,N_1978,N_3450);
or U6969 (N_6969,N_2028,N_3880);
nor U6970 (N_6970,N_1139,N_2214);
nor U6971 (N_6971,N_1085,N_2333);
and U6972 (N_6972,N_999,N_2901);
or U6973 (N_6973,N_200,N_2549);
and U6974 (N_6974,N_1769,N_1138);
nor U6975 (N_6975,N_3614,N_2419);
nor U6976 (N_6976,N_1939,N_1558);
or U6977 (N_6977,N_593,N_2552);
or U6978 (N_6978,N_3444,N_1576);
nor U6979 (N_6979,N_2105,N_2858);
nor U6980 (N_6980,N_3248,N_743);
nor U6981 (N_6981,N_2747,N_3432);
nand U6982 (N_6982,N_3217,N_2765);
or U6983 (N_6983,N_1085,N_240);
xnor U6984 (N_6984,N_1929,N_422);
and U6985 (N_6985,N_1603,N_1866);
or U6986 (N_6986,N_3606,N_1860);
or U6987 (N_6987,N_2454,N_1013);
and U6988 (N_6988,N_1119,N_3450);
nand U6989 (N_6989,N_3916,N_2209);
and U6990 (N_6990,N_1339,N_2909);
and U6991 (N_6991,N_1225,N_3196);
and U6992 (N_6992,N_681,N_764);
nand U6993 (N_6993,N_1273,N_2);
and U6994 (N_6994,N_970,N_3887);
and U6995 (N_6995,N_677,N_178);
and U6996 (N_6996,N_2920,N_3231);
nor U6997 (N_6997,N_1794,N_2037);
or U6998 (N_6998,N_2660,N_796);
and U6999 (N_6999,N_2340,N_353);
nand U7000 (N_7000,N_747,N_1093);
or U7001 (N_7001,N_2892,N_833);
nor U7002 (N_7002,N_1667,N_843);
nand U7003 (N_7003,N_670,N_2731);
nand U7004 (N_7004,N_2985,N_275);
or U7005 (N_7005,N_3254,N_2312);
or U7006 (N_7006,N_3411,N_3349);
nand U7007 (N_7007,N_21,N_1264);
and U7008 (N_7008,N_1869,N_2527);
or U7009 (N_7009,N_3302,N_374);
or U7010 (N_7010,N_3812,N_2851);
and U7011 (N_7011,N_2622,N_3023);
nand U7012 (N_7012,N_3613,N_3065);
nand U7013 (N_7013,N_3220,N_595);
or U7014 (N_7014,N_3339,N_799);
nor U7015 (N_7015,N_1542,N_1407);
nor U7016 (N_7016,N_1891,N_1570);
xnor U7017 (N_7017,N_2649,N_1857);
nor U7018 (N_7018,N_3070,N_2691);
and U7019 (N_7019,N_170,N_161);
nand U7020 (N_7020,N_2520,N_1843);
nand U7021 (N_7021,N_39,N_1711);
and U7022 (N_7022,N_1937,N_706);
nand U7023 (N_7023,N_3374,N_976);
nand U7024 (N_7024,N_608,N_124);
and U7025 (N_7025,N_3239,N_2137);
or U7026 (N_7026,N_3314,N_3694);
nor U7027 (N_7027,N_791,N_2121);
nand U7028 (N_7028,N_625,N_1028);
nor U7029 (N_7029,N_2854,N_3920);
or U7030 (N_7030,N_1002,N_3721);
nand U7031 (N_7031,N_357,N_2741);
nor U7032 (N_7032,N_2684,N_2486);
nand U7033 (N_7033,N_1344,N_2357);
xnor U7034 (N_7034,N_2164,N_2513);
and U7035 (N_7035,N_1735,N_2348);
xnor U7036 (N_7036,N_2928,N_2445);
nand U7037 (N_7037,N_2,N_3672);
or U7038 (N_7038,N_3661,N_2383);
nor U7039 (N_7039,N_248,N_131);
and U7040 (N_7040,N_3566,N_2693);
xnor U7041 (N_7041,N_2564,N_574);
nor U7042 (N_7042,N_1730,N_1299);
and U7043 (N_7043,N_3030,N_544);
or U7044 (N_7044,N_2378,N_2626);
xor U7045 (N_7045,N_3565,N_1050);
xnor U7046 (N_7046,N_401,N_3629);
or U7047 (N_7047,N_2738,N_695);
or U7048 (N_7048,N_3613,N_2714);
nand U7049 (N_7049,N_2545,N_3105);
or U7050 (N_7050,N_2733,N_2945);
or U7051 (N_7051,N_1791,N_2893);
nor U7052 (N_7052,N_1083,N_3751);
and U7053 (N_7053,N_103,N_1436);
nand U7054 (N_7054,N_942,N_1804);
or U7055 (N_7055,N_880,N_635);
xor U7056 (N_7056,N_534,N_2349);
or U7057 (N_7057,N_1116,N_3620);
or U7058 (N_7058,N_2345,N_2943);
nor U7059 (N_7059,N_1208,N_3340);
and U7060 (N_7060,N_742,N_1764);
nand U7061 (N_7061,N_1359,N_2467);
and U7062 (N_7062,N_1784,N_2937);
xor U7063 (N_7063,N_1124,N_3071);
xor U7064 (N_7064,N_3670,N_343);
nand U7065 (N_7065,N_3629,N_2512);
nand U7066 (N_7066,N_1892,N_1090);
xor U7067 (N_7067,N_3161,N_2874);
and U7068 (N_7068,N_2004,N_1260);
xor U7069 (N_7069,N_3663,N_1636);
nor U7070 (N_7070,N_1520,N_3899);
nand U7071 (N_7071,N_278,N_416);
and U7072 (N_7072,N_1894,N_1502);
nand U7073 (N_7073,N_2045,N_2126);
xnor U7074 (N_7074,N_325,N_1535);
or U7075 (N_7075,N_2021,N_3919);
nand U7076 (N_7076,N_3192,N_1508);
and U7077 (N_7077,N_2005,N_406);
and U7078 (N_7078,N_2726,N_2922);
nand U7079 (N_7079,N_2187,N_1203);
or U7080 (N_7080,N_702,N_3884);
xnor U7081 (N_7081,N_3975,N_2807);
and U7082 (N_7082,N_2504,N_3938);
or U7083 (N_7083,N_791,N_1447);
and U7084 (N_7084,N_3931,N_886);
nor U7085 (N_7085,N_95,N_2426);
and U7086 (N_7086,N_797,N_3627);
and U7087 (N_7087,N_1835,N_1160);
xor U7088 (N_7088,N_873,N_909);
and U7089 (N_7089,N_3077,N_1887);
or U7090 (N_7090,N_2742,N_721);
nand U7091 (N_7091,N_1952,N_164);
and U7092 (N_7092,N_1966,N_1793);
nand U7093 (N_7093,N_1017,N_2168);
xor U7094 (N_7094,N_3543,N_3115);
or U7095 (N_7095,N_3859,N_3363);
xnor U7096 (N_7096,N_20,N_887);
nor U7097 (N_7097,N_2334,N_2579);
nand U7098 (N_7098,N_2072,N_1946);
nor U7099 (N_7099,N_178,N_574);
nor U7100 (N_7100,N_1459,N_1484);
and U7101 (N_7101,N_3988,N_262);
nand U7102 (N_7102,N_3636,N_3841);
nand U7103 (N_7103,N_2016,N_797);
or U7104 (N_7104,N_897,N_2794);
and U7105 (N_7105,N_731,N_3280);
nand U7106 (N_7106,N_748,N_249);
and U7107 (N_7107,N_372,N_551);
xor U7108 (N_7108,N_2605,N_820);
nor U7109 (N_7109,N_1135,N_918);
nand U7110 (N_7110,N_2159,N_3821);
nor U7111 (N_7111,N_3960,N_229);
nor U7112 (N_7112,N_3136,N_1734);
nand U7113 (N_7113,N_379,N_3148);
nand U7114 (N_7114,N_137,N_2688);
or U7115 (N_7115,N_2171,N_1110);
nor U7116 (N_7116,N_3813,N_161);
nand U7117 (N_7117,N_2061,N_2622);
nor U7118 (N_7118,N_1565,N_1559);
nor U7119 (N_7119,N_3979,N_1735);
or U7120 (N_7120,N_519,N_3701);
nor U7121 (N_7121,N_2881,N_3861);
nor U7122 (N_7122,N_747,N_3725);
nor U7123 (N_7123,N_2482,N_1006);
nand U7124 (N_7124,N_506,N_324);
and U7125 (N_7125,N_1614,N_1642);
or U7126 (N_7126,N_1074,N_885);
and U7127 (N_7127,N_720,N_2395);
or U7128 (N_7128,N_2499,N_986);
and U7129 (N_7129,N_2281,N_1219);
or U7130 (N_7130,N_3906,N_962);
or U7131 (N_7131,N_3153,N_925);
xor U7132 (N_7132,N_3901,N_141);
or U7133 (N_7133,N_2299,N_1837);
nand U7134 (N_7134,N_3150,N_2139);
nor U7135 (N_7135,N_1250,N_1413);
or U7136 (N_7136,N_2425,N_3863);
nor U7137 (N_7137,N_2761,N_584);
and U7138 (N_7138,N_2723,N_1629);
nor U7139 (N_7139,N_814,N_3633);
nand U7140 (N_7140,N_3681,N_3125);
nor U7141 (N_7141,N_2154,N_291);
nand U7142 (N_7142,N_37,N_415);
nor U7143 (N_7143,N_3134,N_494);
xor U7144 (N_7144,N_443,N_3955);
nand U7145 (N_7145,N_2931,N_3454);
or U7146 (N_7146,N_1844,N_695);
nor U7147 (N_7147,N_2113,N_3524);
nand U7148 (N_7148,N_3472,N_3623);
or U7149 (N_7149,N_2781,N_1760);
or U7150 (N_7150,N_136,N_316);
xnor U7151 (N_7151,N_342,N_1966);
and U7152 (N_7152,N_2059,N_3720);
nor U7153 (N_7153,N_3704,N_198);
xnor U7154 (N_7154,N_1290,N_1619);
nor U7155 (N_7155,N_316,N_21);
nand U7156 (N_7156,N_2714,N_1594);
and U7157 (N_7157,N_3881,N_1714);
nand U7158 (N_7158,N_3530,N_3282);
and U7159 (N_7159,N_85,N_2958);
nand U7160 (N_7160,N_2819,N_3347);
nor U7161 (N_7161,N_1237,N_1685);
nor U7162 (N_7162,N_3711,N_2166);
xnor U7163 (N_7163,N_1710,N_1705);
nand U7164 (N_7164,N_861,N_3855);
or U7165 (N_7165,N_2205,N_730);
or U7166 (N_7166,N_3955,N_317);
and U7167 (N_7167,N_2208,N_3207);
nand U7168 (N_7168,N_2249,N_14);
nor U7169 (N_7169,N_3246,N_2965);
nand U7170 (N_7170,N_541,N_2266);
or U7171 (N_7171,N_1312,N_2314);
nand U7172 (N_7172,N_1205,N_3468);
or U7173 (N_7173,N_3798,N_1423);
and U7174 (N_7174,N_1037,N_2269);
xnor U7175 (N_7175,N_2744,N_585);
nand U7176 (N_7176,N_2823,N_1960);
nand U7177 (N_7177,N_592,N_3587);
nand U7178 (N_7178,N_2206,N_3889);
nand U7179 (N_7179,N_560,N_1761);
nor U7180 (N_7180,N_2562,N_917);
nand U7181 (N_7181,N_3479,N_1368);
nor U7182 (N_7182,N_3301,N_449);
nand U7183 (N_7183,N_3575,N_973);
nand U7184 (N_7184,N_1580,N_890);
xor U7185 (N_7185,N_761,N_3466);
and U7186 (N_7186,N_805,N_333);
nor U7187 (N_7187,N_103,N_2281);
or U7188 (N_7188,N_2262,N_626);
and U7189 (N_7189,N_2004,N_1173);
nand U7190 (N_7190,N_692,N_3032);
and U7191 (N_7191,N_52,N_3393);
nor U7192 (N_7192,N_1144,N_3183);
nand U7193 (N_7193,N_2622,N_2255);
or U7194 (N_7194,N_1927,N_3456);
nor U7195 (N_7195,N_3828,N_312);
nor U7196 (N_7196,N_2067,N_3007);
xor U7197 (N_7197,N_3619,N_3881);
nor U7198 (N_7198,N_179,N_2885);
or U7199 (N_7199,N_2898,N_3001);
and U7200 (N_7200,N_242,N_1365);
xor U7201 (N_7201,N_239,N_2557);
nor U7202 (N_7202,N_1098,N_2055);
or U7203 (N_7203,N_2140,N_1445);
nand U7204 (N_7204,N_40,N_1385);
or U7205 (N_7205,N_2225,N_2644);
and U7206 (N_7206,N_2005,N_1664);
nor U7207 (N_7207,N_3177,N_3257);
xor U7208 (N_7208,N_765,N_1003);
or U7209 (N_7209,N_2227,N_3579);
xnor U7210 (N_7210,N_448,N_752);
or U7211 (N_7211,N_2172,N_2318);
nand U7212 (N_7212,N_3844,N_3458);
nand U7213 (N_7213,N_1802,N_535);
and U7214 (N_7214,N_63,N_1512);
xnor U7215 (N_7215,N_2457,N_3707);
and U7216 (N_7216,N_1952,N_987);
nor U7217 (N_7217,N_3470,N_3571);
and U7218 (N_7218,N_899,N_1802);
and U7219 (N_7219,N_2326,N_3133);
and U7220 (N_7220,N_2688,N_604);
nor U7221 (N_7221,N_2932,N_3938);
or U7222 (N_7222,N_1945,N_2455);
nor U7223 (N_7223,N_26,N_174);
xnor U7224 (N_7224,N_3721,N_3834);
nand U7225 (N_7225,N_3642,N_3481);
nor U7226 (N_7226,N_874,N_1589);
nand U7227 (N_7227,N_2210,N_2627);
or U7228 (N_7228,N_935,N_1741);
nand U7229 (N_7229,N_1976,N_2775);
nor U7230 (N_7230,N_1674,N_169);
xnor U7231 (N_7231,N_2387,N_2453);
or U7232 (N_7232,N_3510,N_3980);
or U7233 (N_7233,N_2581,N_3810);
and U7234 (N_7234,N_1022,N_695);
or U7235 (N_7235,N_2071,N_2408);
nor U7236 (N_7236,N_1359,N_3160);
and U7237 (N_7237,N_1529,N_221);
or U7238 (N_7238,N_3871,N_3325);
nor U7239 (N_7239,N_2186,N_1659);
or U7240 (N_7240,N_2152,N_496);
nand U7241 (N_7241,N_1219,N_3191);
nor U7242 (N_7242,N_3788,N_1276);
and U7243 (N_7243,N_1216,N_3848);
nand U7244 (N_7244,N_3293,N_1286);
nor U7245 (N_7245,N_1842,N_187);
xnor U7246 (N_7246,N_2421,N_307);
xor U7247 (N_7247,N_1105,N_71);
xor U7248 (N_7248,N_3099,N_3470);
or U7249 (N_7249,N_3086,N_1741);
nand U7250 (N_7250,N_2346,N_649);
or U7251 (N_7251,N_2880,N_3952);
nand U7252 (N_7252,N_2341,N_3970);
nand U7253 (N_7253,N_2431,N_2326);
nand U7254 (N_7254,N_3667,N_2896);
or U7255 (N_7255,N_652,N_917);
nand U7256 (N_7256,N_1357,N_666);
and U7257 (N_7257,N_1334,N_1593);
or U7258 (N_7258,N_211,N_1220);
and U7259 (N_7259,N_286,N_755);
or U7260 (N_7260,N_2493,N_2595);
nand U7261 (N_7261,N_3051,N_2254);
xor U7262 (N_7262,N_2916,N_2888);
nor U7263 (N_7263,N_2674,N_1594);
nor U7264 (N_7264,N_1641,N_3625);
and U7265 (N_7265,N_920,N_3444);
nor U7266 (N_7266,N_3625,N_1325);
nand U7267 (N_7267,N_2583,N_1575);
nor U7268 (N_7268,N_1123,N_3350);
xnor U7269 (N_7269,N_3639,N_2929);
or U7270 (N_7270,N_2716,N_3612);
nand U7271 (N_7271,N_2529,N_2132);
nand U7272 (N_7272,N_3633,N_66);
and U7273 (N_7273,N_1265,N_1246);
and U7274 (N_7274,N_758,N_573);
nand U7275 (N_7275,N_3304,N_3429);
xor U7276 (N_7276,N_2207,N_98);
nand U7277 (N_7277,N_60,N_3162);
nor U7278 (N_7278,N_702,N_2537);
nand U7279 (N_7279,N_1063,N_1470);
nor U7280 (N_7280,N_1374,N_3179);
nand U7281 (N_7281,N_3769,N_2357);
and U7282 (N_7282,N_2547,N_3852);
or U7283 (N_7283,N_2014,N_240);
or U7284 (N_7284,N_1429,N_2128);
or U7285 (N_7285,N_2301,N_2785);
and U7286 (N_7286,N_691,N_165);
and U7287 (N_7287,N_2228,N_2922);
nor U7288 (N_7288,N_3354,N_1384);
nand U7289 (N_7289,N_435,N_205);
or U7290 (N_7290,N_829,N_3865);
and U7291 (N_7291,N_3185,N_2649);
nand U7292 (N_7292,N_412,N_2738);
and U7293 (N_7293,N_1727,N_1686);
or U7294 (N_7294,N_3417,N_1862);
or U7295 (N_7295,N_387,N_2486);
nor U7296 (N_7296,N_2473,N_3225);
nor U7297 (N_7297,N_900,N_2817);
xnor U7298 (N_7298,N_1464,N_923);
and U7299 (N_7299,N_847,N_195);
nor U7300 (N_7300,N_3192,N_3586);
nor U7301 (N_7301,N_1722,N_2161);
and U7302 (N_7302,N_416,N_3035);
xnor U7303 (N_7303,N_1545,N_2023);
nor U7304 (N_7304,N_1446,N_2798);
or U7305 (N_7305,N_3589,N_957);
nor U7306 (N_7306,N_638,N_1942);
or U7307 (N_7307,N_270,N_3524);
nor U7308 (N_7308,N_867,N_3211);
or U7309 (N_7309,N_3055,N_2644);
or U7310 (N_7310,N_534,N_3248);
xor U7311 (N_7311,N_2232,N_2698);
or U7312 (N_7312,N_833,N_2883);
nand U7313 (N_7313,N_1458,N_3696);
and U7314 (N_7314,N_749,N_2193);
nand U7315 (N_7315,N_3994,N_2555);
nor U7316 (N_7316,N_1531,N_1510);
nand U7317 (N_7317,N_1806,N_3680);
nor U7318 (N_7318,N_3953,N_1038);
or U7319 (N_7319,N_899,N_931);
nor U7320 (N_7320,N_2697,N_2985);
or U7321 (N_7321,N_772,N_3347);
xor U7322 (N_7322,N_167,N_864);
or U7323 (N_7323,N_1020,N_3135);
or U7324 (N_7324,N_3628,N_359);
and U7325 (N_7325,N_1644,N_3459);
and U7326 (N_7326,N_2402,N_3192);
nand U7327 (N_7327,N_3603,N_3659);
and U7328 (N_7328,N_1801,N_3805);
xnor U7329 (N_7329,N_444,N_2710);
or U7330 (N_7330,N_393,N_1437);
and U7331 (N_7331,N_2409,N_1420);
and U7332 (N_7332,N_545,N_2243);
or U7333 (N_7333,N_2578,N_2290);
nand U7334 (N_7334,N_80,N_49);
or U7335 (N_7335,N_375,N_37);
xor U7336 (N_7336,N_438,N_2318);
or U7337 (N_7337,N_1876,N_2880);
xnor U7338 (N_7338,N_1780,N_3036);
nor U7339 (N_7339,N_3324,N_3996);
xor U7340 (N_7340,N_1922,N_268);
or U7341 (N_7341,N_236,N_504);
nand U7342 (N_7342,N_206,N_1979);
nor U7343 (N_7343,N_2284,N_415);
nor U7344 (N_7344,N_3647,N_2042);
and U7345 (N_7345,N_1641,N_1243);
or U7346 (N_7346,N_2416,N_3042);
nor U7347 (N_7347,N_2327,N_1594);
and U7348 (N_7348,N_2066,N_2602);
or U7349 (N_7349,N_2848,N_185);
nand U7350 (N_7350,N_1671,N_2886);
nand U7351 (N_7351,N_2571,N_2110);
or U7352 (N_7352,N_3314,N_369);
or U7353 (N_7353,N_3483,N_334);
nor U7354 (N_7354,N_3031,N_768);
nor U7355 (N_7355,N_402,N_3339);
nor U7356 (N_7356,N_1394,N_125);
and U7357 (N_7357,N_2510,N_142);
and U7358 (N_7358,N_985,N_1660);
nand U7359 (N_7359,N_2277,N_2912);
and U7360 (N_7360,N_815,N_2961);
nand U7361 (N_7361,N_1352,N_275);
nand U7362 (N_7362,N_2734,N_3257);
nand U7363 (N_7363,N_3520,N_832);
and U7364 (N_7364,N_2986,N_2628);
nand U7365 (N_7365,N_2712,N_742);
nand U7366 (N_7366,N_3299,N_2091);
and U7367 (N_7367,N_125,N_2540);
xor U7368 (N_7368,N_2171,N_3757);
or U7369 (N_7369,N_691,N_76);
and U7370 (N_7370,N_3714,N_1061);
nand U7371 (N_7371,N_1422,N_915);
xor U7372 (N_7372,N_370,N_3845);
nand U7373 (N_7373,N_1894,N_392);
or U7374 (N_7374,N_3923,N_2047);
nand U7375 (N_7375,N_956,N_1979);
nand U7376 (N_7376,N_459,N_1334);
nand U7377 (N_7377,N_2669,N_1161);
xor U7378 (N_7378,N_3579,N_2868);
nor U7379 (N_7379,N_1601,N_3093);
and U7380 (N_7380,N_2811,N_1738);
or U7381 (N_7381,N_3466,N_611);
and U7382 (N_7382,N_1100,N_2195);
and U7383 (N_7383,N_305,N_2372);
or U7384 (N_7384,N_2925,N_32);
or U7385 (N_7385,N_3758,N_2253);
or U7386 (N_7386,N_1681,N_993);
or U7387 (N_7387,N_2543,N_2727);
xnor U7388 (N_7388,N_2258,N_2710);
or U7389 (N_7389,N_1062,N_2669);
nor U7390 (N_7390,N_595,N_1739);
or U7391 (N_7391,N_2465,N_3735);
or U7392 (N_7392,N_1670,N_548);
or U7393 (N_7393,N_55,N_3281);
and U7394 (N_7394,N_1589,N_1313);
or U7395 (N_7395,N_508,N_1894);
and U7396 (N_7396,N_1584,N_3060);
nand U7397 (N_7397,N_3610,N_36);
and U7398 (N_7398,N_2496,N_1154);
xnor U7399 (N_7399,N_572,N_1523);
and U7400 (N_7400,N_2333,N_3771);
nor U7401 (N_7401,N_1428,N_3277);
nor U7402 (N_7402,N_150,N_1511);
and U7403 (N_7403,N_854,N_2082);
nand U7404 (N_7404,N_561,N_96);
nor U7405 (N_7405,N_1504,N_2574);
xor U7406 (N_7406,N_168,N_2715);
nor U7407 (N_7407,N_2371,N_1432);
xnor U7408 (N_7408,N_1792,N_2591);
or U7409 (N_7409,N_2312,N_232);
and U7410 (N_7410,N_2560,N_1490);
nor U7411 (N_7411,N_220,N_460);
nand U7412 (N_7412,N_3866,N_2794);
or U7413 (N_7413,N_303,N_2634);
nand U7414 (N_7414,N_3910,N_3590);
nor U7415 (N_7415,N_2267,N_1208);
or U7416 (N_7416,N_2473,N_308);
and U7417 (N_7417,N_172,N_1273);
nor U7418 (N_7418,N_892,N_671);
nor U7419 (N_7419,N_649,N_1408);
and U7420 (N_7420,N_2729,N_3174);
and U7421 (N_7421,N_1665,N_599);
or U7422 (N_7422,N_3126,N_991);
or U7423 (N_7423,N_3719,N_3817);
and U7424 (N_7424,N_3847,N_1800);
nand U7425 (N_7425,N_1003,N_1185);
nor U7426 (N_7426,N_1421,N_3913);
nor U7427 (N_7427,N_1603,N_3417);
or U7428 (N_7428,N_3910,N_3558);
or U7429 (N_7429,N_2088,N_467);
and U7430 (N_7430,N_9,N_2441);
or U7431 (N_7431,N_3406,N_2460);
xnor U7432 (N_7432,N_2223,N_2205);
nand U7433 (N_7433,N_355,N_389);
nand U7434 (N_7434,N_740,N_88);
nand U7435 (N_7435,N_353,N_2699);
nor U7436 (N_7436,N_934,N_2000);
xor U7437 (N_7437,N_306,N_603);
nand U7438 (N_7438,N_2322,N_2473);
nor U7439 (N_7439,N_3352,N_1662);
xor U7440 (N_7440,N_1074,N_171);
or U7441 (N_7441,N_2193,N_2772);
and U7442 (N_7442,N_2765,N_2156);
and U7443 (N_7443,N_2973,N_2932);
nor U7444 (N_7444,N_1684,N_1696);
or U7445 (N_7445,N_3283,N_2334);
nand U7446 (N_7446,N_3531,N_3881);
nor U7447 (N_7447,N_1162,N_1198);
and U7448 (N_7448,N_2762,N_3694);
nor U7449 (N_7449,N_2573,N_3326);
or U7450 (N_7450,N_552,N_1051);
nor U7451 (N_7451,N_2246,N_1160);
nor U7452 (N_7452,N_803,N_2338);
nor U7453 (N_7453,N_1576,N_186);
xnor U7454 (N_7454,N_2281,N_1027);
or U7455 (N_7455,N_2029,N_2289);
nand U7456 (N_7456,N_1769,N_1533);
xor U7457 (N_7457,N_1857,N_2026);
xor U7458 (N_7458,N_1534,N_2115);
nand U7459 (N_7459,N_1980,N_3128);
nand U7460 (N_7460,N_1351,N_2094);
and U7461 (N_7461,N_2048,N_921);
xor U7462 (N_7462,N_1141,N_1602);
nor U7463 (N_7463,N_3208,N_1114);
and U7464 (N_7464,N_107,N_2189);
nor U7465 (N_7465,N_385,N_3383);
nor U7466 (N_7466,N_2120,N_1822);
nand U7467 (N_7467,N_3047,N_2697);
nor U7468 (N_7468,N_2233,N_117);
and U7469 (N_7469,N_1889,N_3260);
nor U7470 (N_7470,N_1881,N_966);
xor U7471 (N_7471,N_2420,N_602);
and U7472 (N_7472,N_2896,N_635);
and U7473 (N_7473,N_1652,N_3750);
and U7474 (N_7474,N_3286,N_2556);
and U7475 (N_7475,N_2319,N_1082);
xnor U7476 (N_7476,N_2563,N_287);
and U7477 (N_7477,N_3129,N_2361);
nor U7478 (N_7478,N_1603,N_2187);
nand U7479 (N_7479,N_556,N_1385);
and U7480 (N_7480,N_1664,N_1467);
nand U7481 (N_7481,N_2210,N_3242);
or U7482 (N_7482,N_939,N_1571);
xnor U7483 (N_7483,N_2982,N_212);
and U7484 (N_7484,N_1061,N_899);
and U7485 (N_7485,N_2165,N_1392);
and U7486 (N_7486,N_2397,N_2489);
nor U7487 (N_7487,N_3706,N_1209);
nor U7488 (N_7488,N_507,N_2124);
and U7489 (N_7489,N_390,N_479);
and U7490 (N_7490,N_348,N_3969);
nand U7491 (N_7491,N_1740,N_775);
and U7492 (N_7492,N_1969,N_2785);
nor U7493 (N_7493,N_705,N_2399);
nand U7494 (N_7494,N_1199,N_2065);
and U7495 (N_7495,N_2814,N_3049);
nand U7496 (N_7496,N_971,N_3404);
or U7497 (N_7497,N_2440,N_3418);
nor U7498 (N_7498,N_12,N_2735);
and U7499 (N_7499,N_1166,N_1824);
nand U7500 (N_7500,N_3945,N_2250);
or U7501 (N_7501,N_2590,N_1887);
or U7502 (N_7502,N_2466,N_2219);
or U7503 (N_7503,N_3960,N_1711);
nor U7504 (N_7504,N_1342,N_3539);
nor U7505 (N_7505,N_3063,N_2714);
xor U7506 (N_7506,N_3912,N_3197);
and U7507 (N_7507,N_1470,N_3507);
nand U7508 (N_7508,N_3350,N_1870);
and U7509 (N_7509,N_956,N_1756);
nand U7510 (N_7510,N_403,N_3739);
and U7511 (N_7511,N_2455,N_1029);
and U7512 (N_7512,N_2074,N_2894);
or U7513 (N_7513,N_3780,N_3682);
xor U7514 (N_7514,N_954,N_1309);
xnor U7515 (N_7515,N_2283,N_2975);
or U7516 (N_7516,N_3087,N_1313);
nand U7517 (N_7517,N_1075,N_1465);
nor U7518 (N_7518,N_2286,N_342);
nor U7519 (N_7519,N_2076,N_3889);
nor U7520 (N_7520,N_3669,N_1638);
nand U7521 (N_7521,N_2881,N_3521);
nand U7522 (N_7522,N_2921,N_2621);
nor U7523 (N_7523,N_2705,N_120);
xor U7524 (N_7524,N_99,N_2534);
xor U7525 (N_7525,N_3656,N_3239);
nand U7526 (N_7526,N_2017,N_3993);
nor U7527 (N_7527,N_2683,N_708);
or U7528 (N_7528,N_1870,N_654);
xor U7529 (N_7529,N_1964,N_1729);
or U7530 (N_7530,N_1112,N_255);
and U7531 (N_7531,N_1853,N_1523);
nand U7532 (N_7532,N_3426,N_333);
nand U7533 (N_7533,N_1566,N_3523);
and U7534 (N_7534,N_3641,N_571);
and U7535 (N_7535,N_1152,N_2536);
nor U7536 (N_7536,N_2776,N_2752);
and U7537 (N_7537,N_50,N_2783);
and U7538 (N_7538,N_2980,N_314);
nand U7539 (N_7539,N_1783,N_2304);
nor U7540 (N_7540,N_3806,N_2416);
nand U7541 (N_7541,N_955,N_850);
xor U7542 (N_7542,N_3048,N_1041);
nor U7543 (N_7543,N_2810,N_2780);
nand U7544 (N_7544,N_1835,N_1505);
nand U7545 (N_7545,N_2515,N_1588);
nor U7546 (N_7546,N_2227,N_1479);
nor U7547 (N_7547,N_998,N_857);
and U7548 (N_7548,N_1710,N_211);
nand U7549 (N_7549,N_1831,N_659);
nor U7550 (N_7550,N_3204,N_594);
nor U7551 (N_7551,N_40,N_2836);
nand U7552 (N_7552,N_3401,N_1106);
nand U7553 (N_7553,N_3663,N_2872);
or U7554 (N_7554,N_92,N_2019);
and U7555 (N_7555,N_3374,N_622);
nand U7556 (N_7556,N_774,N_2814);
nor U7557 (N_7557,N_318,N_1805);
or U7558 (N_7558,N_1522,N_3474);
nand U7559 (N_7559,N_3847,N_1777);
nand U7560 (N_7560,N_2522,N_1895);
and U7561 (N_7561,N_852,N_1874);
or U7562 (N_7562,N_2418,N_560);
and U7563 (N_7563,N_3093,N_2102);
nor U7564 (N_7564,N_2777,N_3344);
nor U7565 (N_7565,N_657,N_621);
nor U7566 (N_7566,N_2029,N_1841);
or U7567 (N_7567,N_165,N_569);
or U7568 (N_7568,N_1538,N_2466);
xnor U7569 (N_7569,N_2058,N_2753);
or U7570 (N_7570,N_3053,N_2756);
nor U7571 (N_7571,N_1324,N_1226);
nor U7572 (N_7572,N_1780,N_3329);
or U7573 (N_7573,N_3220,N_323);
nand U7574 (N_7574,N_3660,N_1684);
and U7575 (N_7575,N_906,N_1497);
nand U7576 (N_7576,N_1181,N_294);
and U7577 (N_7577,N_3841,N_3495);
and U7578 (N_7578,N_1783,N_3437);
or U7579 (N_7579,N_1894,N_88);
nand U7580 (N_7580,N_1461,N_2891);
xor U7581 (N_7581,N_3099,N_3542);
nand U7582 (N_7582,N_1393,N_870);
and U7583 (N_7583,N_1600,N_1016);
and U7584 (N_7584,N_727,N_786);
nor U7585 (N_7585,N_3677,N_1797);
nor U7586 (N_7586,N_1711,N_894);
or U7587 (N_7587,N_3309,N_3104);
nand U7588 (N_7588,N_2612,N_1837);
or U7589 (N_7589,N_1202,N_1368);
nor U7590 (N_7590,N_2491,N_1317);
and U7591 (N_7591,N_2877,N_1155);
and U7592 (N_7592,N_2935,N_3658);
xor U7593 (N_7593,N_1480,N_2342);
and U7594 (N_7594,N_2558,N_1985);
nor U7595 (N_7595,N_1051,N_585);
and U7596 (N_7596,N_3292,N_1206);
nand U7597 (N_7597,N_2509,N_3712);
nand U7598 (N_7598,N_3732,N_767);
and U7599 (N_7599,N_1653,N_3267);
or U7600 (N_7600,N_2929,N_2731);
or U7601 (N_7601,N_620,N_2228);
nor U7602 (N_7602,N_551,N_1521);
or U7603 (N_7603,N_1954,N_3345);
nor U7604 (N_7604,N_1659,N_1066);
nor U7605 (N_7605,N_1251,N_1764);
nor U7606 (N_7606,N_509,N_1571);
nor U7607 (N_7607,N_2803,N_2344);
or U7608 (N_7608,N_2664,N_3546);
nor U7609 (N_7609,N_2345,N_2268);
nand U7610 (N_7610,N_2927,N_59);
and U7611 (N_7611,N_67,N_3899);
nor U7612 (N_7612,N_1841,N_2604);
or U7613 (N_7613,N_2580,N_2170);
and U7614 (N_7614,N_2336,N_1127);
nor U7615 (N_7615,N_3807,N_3484);
or U7616 (N_7616,N_52,N_1141);
and U7617 (N_7617,N_3362,N_3097);
nand U7618 (N_7618,N_1168,N_1942);
or U7619 (N_7619,N_1341,N_2073);
or U7620 (N_7620,N_728,N_27);
and U7621 (N_7621,N_2245,N_2639);
and U7622 (N_7622,N_1321,N_3261);
and U7623 (N_7623,N_3994,N_2368);
nand U7624 (N_7624,N_305,N_203);
xnor U7625 (N_7625,N_2460,N_2841);
and U7626 (N_7626,N_2807,N_616);
xnor U7627 (N_7627,N_1080,N_3140);
nor U7628 (N_7628,N_1205,N_512);
xnor U7629 (N_7629,N_1186,N_1710);
xor U7630 (N_7630,N_2931,N_462);
xor U7631 (N_7631,N_1066,N_2014);
nor U7632 (N_7632,N_2368,N_3902);
and U7633 (N_7633,N_855,N_3606);
nor U7634 (N_7634,N_1093,N_1331);
or U7635 (N_7635,N_2959,N_288);
or U7636 (N_7636,N_3704,N_1355);
and U7637 (N_7637,N_1034,N_3433);
or U7638 (N_7638,N_294,N_2535);
nor U7639 (N_7639,N_3750,N_3234);
and U7640 (N_7640,N_3487,N_2537);
nor U7641 (N_7641,N_910,N_3563);
and U7642 (N_7642,N_1862,N_3709);
nor U7643 (N_7643,N_2009,N_1908);
nand U7644 (N_7644,N_3144,N_249);
nand U7645 (N_7645,N_2471,N_1087);
nor U7646 (N_7646,N_940,N_783);
and U7647 (N_7647,N_2834,N_3794);
nand U7648 (N_7648,N_3634,N_195);
or U7649 (N_7649,N_2477,N_3072);
or U7650 (N_7650,N_1350,N_2827);
nand U7651 (N_7651,N_1907,N_932);
or U7652 (N_7652,N_892,N_3194);
and U7653 (N_7653,N_3225,N_1560);
or U7654 (N_7654,N_3526,N_3036);
and U7655 (N_7655,N_3507,N_1346);
and U7656 (N_7656,N_2,N_3299);
nand U7657 (N_7657,N_2449,N_2903);
nor U7658 (N_7658,N_1616,N_1986);
nor U7659 (N_7659,N_2635,N_1033);
nor U7660 (N_7660,N_3334,N_3504);
or U7661 (N_7661,N_1354,N_1185);
or U7662 (N_7662,N_2984,N_2919);
and U7663 (N_7663,N_3673,N_1163);
nor U7664 (N_7664,N_256,N_2659);
nand U7665 (N_7665,N_464,N_1254);
or U7666 (N_7666,N_1490,N_2765);
and U7667 (N_7667,N_3445,N_2871);
nand U7668 (N_7668,N_3152,N_1838);
nand U7669 (N_7669,N_2851,N_2439);
or U7670 (N_7670,N_1268,N_2371);
or U7671 (N_7671,N_2131,N_54);
and U7672 (N_7672,N_175,N_799);
nor U7673 (N_7673,N_2348,N_397);
nor U7674 (N_7674,N_2904,N_1644);
nand U7675 (N_7675,N_1225,N_3561);
or U7676 (N_7676,N_1915,N_1752);
nand U7677 (N_7677,N_2865,N_867);
and U7678 (N_7678,N_2608,N_1053);
and U7679 (N_7679,N_3160,N_368);
xor U7680 (N_7680,N_2165,N_2599);
and U7681 (N_7681,N_177,N_1582);
and U7682 (N_7682,N_2578,N_1682);
or U7683 (N_7683,N_3655,N_2472);
xor U7684 (N_7684,N_1963,N_2067);
nand U7685 (N_7685,N_2878,N_1);
and U7686 (N_7686,N_488,N_1677);
and U7687 (N_7687,N_1243,N_336);
nand U7688 (N_7688,N_1045,N_1987);
or U7689 (N_7689,N_3130,N_1864);
and U7690 (N_7690,N_313,N_3562);
nor U7691 (N_7691,N_1659,N_2352);
xor U7692 (N_7692,N_215,N_2891);
and U7693 (N_7693,N_2896,N_1598);
and U7694 (N_7694,N_391,N_3201);
and U7695 (N_7695,N_678,N_1873);
nand U7696 (N_7696,N_1418,N_1176);
nand U7697 (N_7697,N_3487,N_848);
and U7698 (N_7698,N_2936,N_2448);
and U7699 (N_7699,N_1645,N_1674);
or U7700 (N_7700,N_2769,N_2301);
nor U7701 (N_7701,N_3912,N_1879);
nor U7702 (N_7702,N_87,N_3204);
and U7703 (N_7703,N_3016,N_147);
nor U7704 (N_7704,N_1250,N_1260);
xor U7705 (N_7705,N_3572,N_3494);
nand U7706 (N_7706,N_47,N_3448);
nand U7707 (N_7707,N_3124,N_920);
or U7708 (N_7708,N_514,N_1411);
nor U7709 (N_7709,N_3116,N_3725);
nor U7710 (N_7710,N_1224,N_1143);
or U7711 (N_7711,N_1464,N_525);
nor U7712 (N_7712,N_841,N_281);
nor U7713 (N_7713,N_3221,N_2305);
and U7714 (N_7714,N_1721,N_2888);
xor U7715 (N_7715,N_1396,N_309);
nand U7716 (N_7716,N_2505,N_62);
and U7717 (N_7717,N_504,N_3781);
nor U7718 (N_7718,N_1089,N_3435);
and U7719 (N_7719,N_3431,N_3880);
nor U7720 (N_7720,N_2596,N_500);
nand U7721 (N_7721,N_3586,N_2151);
nor U7722 (N_7722,N_2801,N_3280);
nor U7723 (N_7723,N_1064,N_279);
nor U7724 (N_7724,N_50,N_2342);
and U7725 (N_7725,N_1912,N_3289);
and U7726 (N_7726,N_1542,N_3504);
or U7727 (N_7727,N_1141,N_469);
and U7728 (N_7728,N_1540,N_1317);
and U7729 (N_7729,N_3533,N_3397);
nor U7730 (N_7730,N_1285,N_1646);
xnor U7731 (N_7731,N_804,N_2190);
nor U7732 (N_7732,N_3754,N_1194);
or U7733 (N_7733,N_1360,N_2675);
and U7734 (N_7734,N_908,N_2678);
or U7735 (N_7735,N_2811,N_3588);
nand U7736 (N_7736,N_1315,N_2426);
nand U7737 (N_7737,N_2481,N_3649);
and U7738 (N_7738,N_59,N_1555);
and U7739 (N_7739,N_2020,N_3307);
nand U7740 (N_7740,N_2084,N_2508);
and U7741 (N_7741,N_2301,N_692);
xnor U7742 (N_7742,N_1099,N_551);
or U7743 (N_7743,N_1419,N_358);
xor U7744 (N_7744,N_2602,N_2958);
and U7745 (N_7745,N_617,N_2090);
and U7746 (N_7746,N_976,N_2448);
and U7747 (N_7747,N_3957,N_1657);
nor U7748 (N_7748,N_2209,N_636);
or U7749 (N_7749,N_1723,N_1032);
and U7750 (N_7750,N_1218,N_1125);
nand U7751 (N_7751,N_3022,N_3408);
nand U7752 (N_7752,N_945,N_3243);
nand U7753 (N_7753,N_3340,N_447);
xor U7754 (N_7754,N_831,N_1529);
nand U7755 (N_7755,N_508,N_1227);
or U7756 (N_7756,N_2768,N_1973);
xor U7757 (N_7757,N_875,N_2677);
nor U7758 (N_7758,N_2374,N_389);
or U7759 (N_7759,N_583,N_1177);
and U7760 (N_7760,N_1976,N_2509);
or U7761 (N_7761,N_1765,N_1404);
nand U7762 (N_7762,N_2098,N_2401);
or U7763 (N_7763,N_236,N_352);
or U7764 (N_7764,N_1184,N_2186);
and U7765 (N_7765,N_2066,N_2537);
or U7766 (N_7766,N_2121,N_3307);
or U7767 (N_7767,N_278,N_2797);
or U7768 (N_7768,N_820,N_1209);
nor U7769 (N_7769,N_468,N_3605);
nor U7770 (N_7770,N_842,N_2274);
and U7771 (N_7771,N_711,N_1694);
nand U7772 (N_7772,N_624,N_3932);
nor U7773 (N_7773,N_2174,N_846);
xnor U7774 (N_7774,N_1618,N_262);
nand U7775 (N_7775,N_1160,N_2804);
nand U7776 (N_7776,N_1360,N_1041);
xnor U7777 (N_7777,N_231,N_2485);
nor U7778 (N_7778,N_3814,N_2612);
nor U7779 (N_7779,N_975,N_2622);
nor U7780 (N_7780,N_1586,N_3276);
or U7781 (N_7781,N_2031,N_1478);
nand U7782 (N_7782,N_2858,N_1308);
nor U7783 (N_7783,N_2268,N_2289);
nand U7784 (N_7784,N_100,N_37);
nor U7785 (N_7785,N_3884,N_1452);
nor U7786 (N_7786,N_2213,N_1305);
xnor U7787 (N_7787,N_3368,N_3322);
xnor U7788 (N_7788,N_2725,N_2646);
nor U7789 (N_7789,N_1128,N_916);
xor U7790 (N_7790,N_1400,N_1164);
and U7791 (N_7791,N_2097,N_3722);
or U7792 (N_7792,N_462,N_3751);
nor U7793 (N_7793,N_3153,N_1563);
nand U7794 (N_7794,N_2659,N_2186);
nand U7795 (N_7795,N_1371,N_3765);
nand U7796 (N_7796,N_1547,N_1999);
xor U7797 (N_7797,N_3661,N_2432);
xnor U7798 (N_7798,N_2323,N_34);
nor U7799 (N_7799,N_339,N_432);
nor U7800 (N_7800,N_858,N_1628);
and U7801 (N_7801,N_2124,N_1378);
nor U7802 (N_7802,N_2498,N_369);
and U7803 (N_7803,N_363,N_1427);
nor U7804 (N_7804,N_488,N_2653);
nor U7805 (N_7805,N_275,N_2193);
and U7806 (N_7806,N_3980,N_1356);
or U7807 (N_7807,N_25,N_1850);
xnor U7808 (N_7808,N_55,N_912);
xnor U7809 (N_7809,N_3378,N_2452);
or U7810 (N_7810,N_1954,N_2899);
or U7811 (N_7811,N_2778,N_2501);
xnor U7812 (N_7812,N_2623,N_179);
or U7813 (N_7813,N_1539,N_3968);
nor U7814 (N_7814,N_564,N_174);
nor U7815 (N_7815,N_676,N_2466);
xnor U7816 (N_7816,N_1073,N_1637);
xnor U7817 (N_7817,N_332,N_727);
or U7818 (N_7818,N_752,N_144);
or U7819 (N_7819,N_2812,N_1255);
nor U7820 (N_7820,N_1844,N_2004);
nor U7821 (N_7821,N_3489,N_848);
xor U7822 (N_7822,N_703,N_3494);
nand U7823 (N_7823,N_330,N_1853);
or U7824 (N_7824,N_2325,N_3057);
xnor U7825 (N_7825,N_329,N_3933);
and U7826 (N_7826,N_1687,N_3936);
nand U7827 (N_7827,N_306,N_2477);
nand U7828 (N_7828,N_2905,N_1937);
xnor U7829 (N_7829,N_3557,N_278);
and U7830 (N_7830,N_2127,N_12);
or U7831 (N_7831,N_1217,N_3528);
nand U7832 (N_7832,N_3706,N_1613);
nand U7833 (N_7833,N_620,N_225);
nor U7834 (N_7834,N_2221,N_3609);
nor U7835 (N_7835,N_123,N_2663);
or U7836 (N_7836,N_3706,N_2429);
nor U7837 (N_7837,N_877,N_3269);
nor U7838 (N_7838,N_3336,N_828);
xor U7839 (N_7839,N_1885,N_3905);
nand U7840 (N_7840,N_3481,N_2188);
or U7841 (N_7841,N_2007,N_2168);
nand U7842 (N_7842,N_1977,N_1375);
or U7843 (N_7843,N_3257,N_2429);
nand U7844 (N_7844,N_3831,N_2035);
and U7845 (N_7845,N_2625,N_625);
nand U7846 (N_7846,N_1969,N_2071);
and U7847 (N_7847,N_2612,N_2483);
and U7848 (N_7848,N_814,N_3738);
nand U7849 (N_7849,N_3481,N_1008);
nor U7850 (N_7850,N_839,N_2198);
nand U7851 (N_7851,N_1284,N_3044);
xor U7852 (N_7852,N_2972,N_3051);
or U7853 (N_7853,N_80,N_1249);
nor U7854 (N_7854,N_2621,N_952);
and U7855 (N_7855,N_1935,N_3884);
xnor U7856 (N_7856,N_2835,N_3961);
xnor U7857 (N_7857,N_581,N_1922);
nand U7858 (N_7858,N_981,N_2507);
or U7859 (N_7859,N_234,N_2935);
or U7860 (N_7860,N_3869,N_1622);
nand U7861 (N_7861,N_963,N_1612);
nand U7862 (N_7862,N_589,N_3774);
nor U7863 (N_7863,N_620,N_1925);
and U7864 (N_7864,N_3496,N_1947);
and U7865 (N_7865,N_2273,N_472);
nand U7866 (N_7866,N_3729,N_448);
nand U7867 (N_7867,N_2372,N_2710);
and U7868 (N_7868,N_2473,N_1277);
or U7869 (N_7869,N_939,N_3321);
or U7870 (N_7870,N_3428,N_2816);
nand U7871 (N_7871,N_2953,N_3982);
nand U7872 (N_7872,N_3714,N_1823);
or U7873 (N_7873,N_2489,N_1021);
or U7874 (N_7874,N_1525,N_1591);
and U7875 (N_7875,N_2127,N_3225);
or U7876 (N_7876,N_656,N_593);
nand U7877 (N_7877,N_1999,N_1393);
and U7878 (N_7878,N_2293,N_3593);
and U7879 (N_7879,N_2695,N_2178);
or U7880 (N_7880,N_3013,N_1806);
or U7881 (N_7881,N_298,N_3689);
and U7882 (N_7882,N_2549,N_1811);
nand U7883 (N_7883,N_3566,N_1404);
and U7884 (N_7884,N_2195,N_3697);
or U7885 (N_7885,N_3634,N_559);
or U7886 (N_7886,N_384,N_3301);
nand U7887 (N_7887,N_2645,N_3296);
xor U7888 (N_7888,N_3386,N_3218);
and U7889 (N_7889,N_892,N_3461);
and U7890 (N_7890,N_563,N_2863);
nor U7891 (N_7891,N_3111,N_79);
xor U7892 (N_7892,N_2877,N_1399);
nand U7893 (N_7893,N_2132,N_930);
and U7894 (N_7894,N_2342,N_2226);
or U7895 (N_7895,N_610,N_2118);
nand U7896 (N_7896,N_1732,N_44);
and U7897 (N_7897,N_3444,N_328);
xnor U7898 (N_7898,N_1215,N_1489);
nand U7899 (N_7899,N_3065,N_1724);
nor U7900 (N_7900,N_1172,N_3288);
or U7901 (N_7901,N_982,N_3698);
nand U7902 (N_7902,N_2682,N_440);
nand U7903 (N_7903,N_723,N_2074);
nor U7904 (N_7904,N_669,N_941);
or U7905 (N_7905,N_3745,N_3432);
nand U7906 (N_7906,N_1649,N_1640);
nor U7907 (N_7907,N_1336,N_1226);
or U7908 (N_7908,N_592,N_2800);
nor U7909 (N_7909,N_1763,N_872);
or U7910 (N_7910,N_3837,N_2677);
or U7911 (N_7911,N_1923,N_354);
nor U7912 (N_7912,N_283,N_268);
and U7913 (N_7913,N_3428,N_219);
or U7914 (N_7914,N_713,N_1365);
nand U7915 (N_7915,N_3880,N_3681);
xnor U7916 (N_7916,N_2648,N_552);
and U7917 (N_7917,N_3886,N_1709);
nand U7918 (N_7918,N_2793,N_3252);
and U7919 (N_7919,N_1570,N_3939);
and U7920 (N_7920,N_3764,N_485);
and U7921 (N_7921,N_598,N_1173);
and U7922 (N_7922,N_1233,N_1929);
nand U7923 (N_7923,N_603,N_3971);
or U7924 (N_7924,N_3847,N_3625);
nand U7925 (N_7925,N_3682,N_1968);
and U7926 (N_7926,N_218,N_1381);
nor U7927 (N_7927,N_990,N_349);
nor U7928 (N_7928,N_1329,N_2798);
nor U7929 (N_7929,N_3441,N_1233);
nand U7930 (N_7930,N_1431,N_347);
nand U7931 (N_7931,N_1444,N_3135);
xnor U7932 (N_7932,N_3621,N_836);
or U7933 (N_7933,N_2752,N_3668);
or U7934 (N_7934,N_1336,N_2898);
or U7935 (N_7935,N_1247,N_2678);
nor U7936 (N_7936,N_3680,N_233);
or U7937 (N_7937,N_1074,N_1878);
or U7938 (N_7938,N_3409,N_1005);
nor U7939 (N_7939,N_1023,N_1792);
nor U7940 (N_7940,N_3580,N_2620);
nand U7941 (N_7941,N_462,N_246);
and U7942 (N_7942,N_1245,N_95);
and U7943 (N_7943,N_3257,N_146);
or U7944 (N_7944,N_3050,N_527);
and U7945 (N_7945,N_1137,N_1204);
xnor U7946 (N_7946,N_571,N_3787);
nand U7947 (N_7947,N_242,N_1591);
nor U7948 (N_7948,N_3746,N_3334);
nand U7949 (N_7949,N_2572,N_432);
or U7950 (N_7950,N_1078,N_390);
nand U7951 (N_7951,N_833,N_2510);
and U7952 (N_7952,N_2447,N_2356);
xor U7953 (N_7953,N_1563,N_3140);
nor U7954 (N_7954,N_1405,N_3339);
or U7955 (N_7955,N_1065,N_3065);
nand U7956 (N_7956,N_858,N_943);
and U7957 (N_7957,N_3216,N_1163);
nand U7958 (N_7958,N_3840,N_1055);
nand U7959 (N_7959,N_4,N_1006);
nand U7960 (N_7960,N_2622,N_2644);
nand U7961 (N_7961,N_3212,N_863);
nand U7962 (N_7962,N_1878,N_87);
nand U7963 (N_7963,N_1677,N_3043);
or U7964 (N_7964,N_182,N_2008);
or U7965 (N_7965,N_12,N_45);
or U7966 (N_7966,N_1360,N_2921);
and U7967 (N_7967,N_1191,N_1173);
and U7968 (N_7968,N_3899,N_2361);
and U7969 (N_7969,N_3809,N_909);
and U7970 (N_7970,N_2254,N_764);
nand U7971 (N_7971,N_3499,N_2336);
or U7972 (N_7972,N_2406,N_2822);
and U7973 (N_7973,N_569,N_1333);
and U7974 (N_7974,N_3272,N_2838);
and U7975 (N_7975,N_877,N_1644);
nor U7976 (N_7976,N_1339,N_2433);
nor U7977 (N_7977,N_2956,N_3659);
and U7978 (N_7978,N_185,N_3502);
and U7979 (N_7979,N_663,N_2098);
nor U7980 (N_7980,N_3745,N_1478);
nor U7981 (N_7981,N_1216,N_3579);
and U7982 (N_7982,N_2173,N_3449);
nor U7983 (N_7983,N_2558,N_956);
nor U7984 (N_7984,N_3792,N_2585);
or U7985 (N_7985,N_1738,N_1449);
nand U7986 (N_7986,N_2758,N_3131);
and U7987 (N_7987,N_311,N_3932);
and U7988 (N_7988,N_1128,N_1754);
xor U7989 (N_7989,N_953,N_370);
and U7990 (N_7990,N_375,N_3146);
or U7991 (N_7991,N_1247,N_1216);
nand U7992 (N_7992,N_3863,N_1290);
xnor U7993 (N_7993,N_3367,N_1236);
and U7994 (N_7994,N_2279,N_1471);
nand U7995 (N_7995,N_574,N_1151);
or U7996 (N_7996,N_2719,N_1708);
nand U7997 (N_7997,N_38,N_1963);
or U7998 (N_7998,N_2373,N_650);
nand U7999 (N_7999,N_3099,N_269);
and U8000 (N_8000,N_4977,N_4271);
and U8001 (N_8001,N_6992,N_6839);
or U8002 (N_8002,N_7914,N_7792);
and U8003 (N_8003,N_7292,N_4036);
or U8004 (N_8004,N_5537,N_7529);
nand U8005 (N_8005,N_7653,N_5275);
and U8006 (N_8006,N_4479,N_7420);
and U8007 (N_8007,N_7394,N_4264);
or U8008 (N_8008,N_6500,N_5533);
nand U8009 (N_8009,N_4139,N_4591);
or U8010 (N_8010,N_5729,N_6808);
nor U8011 (N_8011,N_4365,N_6843);
or U8012 (N_8012,N_7576,N_5828);
nor U8013 (N_8013,N_5498,N_5393);
and U8014 (N_8014,N_5089,N_6665);
or U8015 (N_8015,N_5176,N_7213);
xnor U8016 (N_8016,N_4832,N_4802);
and U8017 (N_8017,N_7030,N_5338);
or U8018 (N_8018,N_5316,N_5640);
and U8019 (N_8019,N_6383,N_4649);
and U8020 (N_8020,N_6260,N_7434);
and U8021 (N_8021,N_7722,N_7528);
and U8022 (N_8022,N_7675,N_7437);
nand U8023 (N_8023,N_5630,N_5797);
nor U8024 (N_8024,N_6675,N_5831);
nor U8025 (N_8025,N_5981,N_7823);
or U8026 (N_8026,N_5241,N_5815);
and U8027 (N_8027,N_4637,N_5890);
nor U8028 (N_8028,N_4806,N_6540);
nor U8029 (N_8029,N_6418,N_7808);
or U8030 (N_8030,N_4237,N_5078);
or U8031 (N_8031,N_6167,N_6371);
and U8032 (N_8032,N_7705,N_6460);
and U8033 (N_8033,N_7926,N_6049);
nand U8034 (N_8034,N_7215,N_4339);
nor U8035 (N_8035,N_7759,N_7524);
nor U8036 (N_8036,N_5020,N_4896);
nand U8037 (N_8037,N_4048,N_7659);
nand U8038 (N_8038,N_4951,N_5614);
nand U8039 (N_8039,N_7028,N_4984);
or U8040 (N_8040,N_6569,N_6374);
nand U8041 (N_8041,N_5723,N_6150);
nand U8042 (N_8042,N_6325,N_4699);
and U8043 (N_8043,N_7970,N_4549);
or U8044 (N_8044,N_4269,N_4097);
or U8045 (N_8045,N_4386,N_6180);
or U8046 (N_8046,N_7344,N_7731);
or U8047 (N_8047,N_7170,N_7564);
or U8048 (N_8048,N_4650,N_6246);
nor U8049 (N_8049,N_6193,N_5520);
nor U8050 (N_8050,N_4065,N_5497);
and U8051 (N_8051,N_6161,N_5691);
xnor U8052 (N_8052,N_6506,N_4535);
and U8053 (N_8053,N_7060,N_5978);
nand U8054 (N_8054,N_4162,N_5915);
nor U8055 (N_8055,N_7253,N_4175);
or U8056 (N_8056,N_7007,N_4983);
nor U8057 (N_8057,N_6596,N_7645);
nor U8058 (N_8058,N_7918,N_4192);
nand U8059 (N_8059,N_7136,N_7508);
or U8060 (N_8060,N_5342,N_6566);
nand U8061 (N_8061,N_7967,N_6057);
nand U8062 (N_8062,N_4800,N_5866);
or U8063 (N_8063,N_7198,N_5598);
nand U8064 (N_8064,N_6767,N_7015);
and U8065 (N_8065,N_6893,N_5127);
nand U8066 (N_8066,N_4655,N_4739);
nor U8067 (N_8067,N_4556,N_4058);
and U8068 (N_8068,N_5642,N_4672);
and U8069 (N_8069,N_7257,N_7486);
or U8070 (N_8070,N_5024,N_5790);
or U8071 (N_8071,N_5712,N_5119);
and U8072 (N_8072,N_5715,N_5561);
and U8073 (N_8073,N_5923,N_7336);
nor U8074 (N_8074,N_6457,N_7484);
nand U8075 (N_8075,N_6414,N_7747);
nand U8076 (N_8076,N_4747,N_7280);
and U8077 (N_8077,N_4706,N_5986);
nand U8078 (N_8078,N_7848,N_7948);
or U8079 (N_8079,N_7322,N_4403);
nand U8080 (N_8080,N_6033,N_7507);
xor U8081 (N_8081,N_7575,N_6858);
xnor U8082 (N_8082,N_4457,N_5171);
and U8083 (N_8083,N_7372,N_7021);
nor U8084 (N_8084,N_5179,N_5971);
and U8085 (N_8085,N_5679,N_6873);
and U8086 (N_8086,N_5752,N_5268);
or U8087 (N_8087,N_6668,N_5002);
xor U8088 (N_8088,N_5294,N_5508);
nor U8089 (N_8089,N_7511,N_7699);
nand U8090 (N_8090,N_5647,N_4049);
and U8091 (N_8091,N_4679,N_5433);
nand U8092 (N_8092,N_6357,N_4309);
and U8093 (N_8093,N_4647,N_6101);
or U8094 (N_8094,N_5129,N_7019);
and U8095 (N_8095,N_6170,N_7519);
nand U8096 (N_8096,N_4117,N_6689);
or U8097 (N_8097,N_5776,N_6078);
nand U8098 (N_8098,N_6929,N_7192);
and U8099 (N_8099,N_6548,N_7742);
and U8100 (N_8100,N_5746,N_6127);
or U8101 (N_8101,N_7798,N_5962);
nand U8102 (N_8102,N_6313,N_4427);
and U8103 (N_8103,N_5237,N_7563);
or U8104 (N_8104,N_7211,N_5800);
and U8105 (N_8105,N_6226,N_7230);
nand U8106 (N_8106,N_7724,N_4718);
and U8107 (N_8107,N_7728,N_5466);
nand U8108 (N_8108,N_4456,N_6289);
nand U8109 (N_8109,N_5845,N_7039);
nor U8110 (N_8110,N_7812,N_6177);
nand U8111 (N_8111,N_5054,N_4317);
or U8112 (N_8112,N_7342,N_5391);
nand U8113 (N_8113,N_7713,N_6716);
nor U8114 (N_8114,N_7913,N_5034);
nor U8115 (N_8115,N_5827,N_4367);
or U8116 (N_8116,N_4858,N_4203);
or U8117 (N_8117,N_5768,N_4540);
and U8118 (N_8118,N_4410,N_4771);
xnor U8119 (N_8119,N_5190,N_4939);
or U8120 (N_8120,N_6221,N_4823);
nand U8121 (N_8121,N_6205,N_7591);
nor U8122 (N_8122,N_4232,N_6681);
nor U8123 (N_8123,N_5101,N_5091);
or U8124 (N_8124,N_5577,N_7071);
nor U8125 (N_8125,N_5925,N_6484);
nand U8126 (N_8126,N_7923,N_6467);
nor U8127 (N_8127,N_4153,N_7952);
nor U8128 (N_8128,N_4093,N_5567);
nand U8129 (N_8129,N_4357,N_6222);
nand U8130 (N_8130,N_4736,N_5726);
and U8131 (N_8131,N_4653,N_4876);
or U8132 (N_8132,N_5629,N_4678);
and U8133 (N_8133,N_4099,N_4111);
or U8134 (N_8134,N_7741,N_6669);
nor U8135 (N_8135,N_7387,N_5059);
or U8136 (N_8136,N_4543,N_4319);
or U8137 (N_8137,N_7629,N_5450);
and U8138 (N_8138,N_6069,N_5330);
nor U8139 (N_8139,N_5596,N_7890);
nand U8140 (N_8140,N_7116,N_5370);
xnor U8141 (N_8141,N_7580,N_4283);
or U8142 (N_8142,N_6288,N_5114);
and U8143 (N_8143,N_5215,N_4483);
or U8144 (N_8144,N_5998,N_7963);
or U8145 (N_8145,N_7882,N_6585);
nand U8146 (N_8146,N_5161,N_5501);
nand U8147 (N_8147,N_4826,N_5810);
and U8148 (N_8148,N_4711,N_6666);
or U8149 (N_8149,N_6030,N_7047);
nor U8150 (N_8150,N_6744,N_7026);
and U8151 (N_8151,N_4617,N_5397);
or U8152 (N_8152,N_7202,N_5584);
and U8153 (N_8153,N_6159,N_7604);
or U8154 (N_8154,N_4859,N_5731);
nor U8155 (N_8155,N_7538,N_7837);
nor U8156 (N_8156,N_4918,N_4805);
nand U8157 (N_8157,N_4392,N_5774);
nand U8158 (N_8158,N_7874,N_6541);
or U8159 (N_8159,N_5053,N_4866);
nor U8160 (N_8160,N_4369,N_4752);
and U8161 (N_8161,N_5755,N_7103);
or U8162 (N_8162,N_5112,N_5488);
or U8163 (N_8163,N_5126,N_5489);
nor U8164 (N_8164,N_6395,N_5144);
nand U8165 (N_8165,N_7270,N_5136);
and U8166 (N_8166,N_5359,N_6187);
nor U8167 (N_8167,N_5884,N_6268);
or U8168 (N_8168,N_6577,N_6447);
nand U8169 (N_8169,N_5337,N_6622);
or U8170 (N_8170,N_7842,N_6904);
nand U8171 (N_8171,N_5992,N_4627);
nor U8172 (N_8172,N_6185,N_4495);
nand U8173 (N_8173,N_5673,N_4172);
xnor U8174 (N_8174,N_4976,N_7343);
nand U8175 (N_8175,N_5867,N_7481);
xor U8176 (N_8176,N_6199,N_7818);
or U8177 (N_8177,N_7536,N_6113);
or U8178 (N_8178,N_5902,N_4467);
xnor U8179 (N_8179,N_5582,N_4725);
nand U8180 (N_8180,N_5667,N_4697);
nor U8181 (N_8181,N_7717,N_4925);
or U8182 (N_8182,N_6864,N_7618);
xnor U8183 (N_8183,N_5722,N_7477);
nor U8184 (N_8184,N_6483,N_6774);
nor U8185 (N_8185,N_5764,N_7846);
or U8186 (N_8186,N_4384,N_6836);
or U8187 (N_8187,N_6311,N_5261);
or U8188 (N_8188,N_5977,N_4607);
xnor U8189 (N_8189,N_6018,N_7549);
and U8190 (N_8190,N_6935,N_7543);
or U8191 (N_8191,N_7735,N_7700);
and U8192 (N_8192,N_4121,N_7912);
nor U8193 (N_8193,N_7844,N_7694);
xor U8194 (N_8194,N_4792,N_7256);
nand U8195 (N_8195,N_7302,N_7303);
and U8196 (N_8196,N_7318,N_7858);
nand U8197 (N_8197,N_7402,N_7853);
and U8198 (N_8198,N_4374,N_4767);
nor U8199 (N_8199,N_4790,N_6280);
and U8200 (N_8200,N_7405,N_4251);
and U8201 (N_8201,N_5278,N_5321);
nor U8202 (N_8202,N_6820,N_4406);
or U8203 (N_8203,N_6857,N_5872);
nor U8204 (N_8204,N_7693,N_4590);
or U8205 (N_8205,N_7241,N_6146);
nand U8206 (N_8206,N_5514,N_5988);
and U8207 (N_8207,N_7894,N_4003);
xor U8208 (N_8208,N_7815,N_4020);
or U8209 (N_8209,N_7445,N_5188);
and U8210 (N_8210,N_4361,N_4994);
or U8211 (N_8211,N_7287,N_4959);
and U8212 (N_8212,N_6007,N_5841);
or U8213 (N_8213,N_7781,N_6564);
and U8214 (N_8214,N_4713,N_4052);
nand U8215 (N_8215,N_7867,N_5661);
and U8216 (N_8216,N_7570,N_6570);
or U8217 (N_8217,N_7165,N_6446);
or U8218 (N_8218,N_4614,N_5648);
nor U8219 (N_8219,N_4033,N_6402);
xnor U8220 (N_8220,N_5784,N_5331);
nor U8221 (N_8221,N_7355,N_6777);
or U8222 (N_8222,N_6776,N_5315);
nand U8223 (N_8223,N_5181,N_4334);
nand U8224 (N_8224,N_4997,N_6501);
or U8225 (N_8225,N_7623,N_4761);
nor U8226 (N_8226,N_5571,N_7692);
nand U8227 (N_8227,N_7573,N_5960);
nor U8228 (N_8228,N_4423,N_7951);
nand U8229 (N_8229,N_7064,N_7690);
and U8230 (N_8230,N_4030,N_7817);
nand U8231 (N_8231,N_7606,N_5506);
nor U8232 (N_8232,N_5502,N_6971);
xor U8233 (N_8233,N_7525,N_7955);
or U8234 (N_8234,N_5684,N_4195);
nor U8235 (N_8235,N_4857,N_5756);
and U8236 (N_8236,N_7979,N_6064);
or U8237 (N_8237,N_5157,N_7650);
xnor U8238 (N_8238,N_6378,N_4814);
or U8239 (N_8239,N_4810,N_6201);
nor U8240 (N_8240,N_6735,N_6215);
and U8241 (N_8241,N_7440,N_5682);
or U8242 (N_8242,N_5467,N_5895);
nand U8243 (N_8243,N_6551,N_6968);
nor U8244 (N_8244,N_7162,N_7857);
or U8245 (N_8245,N_7959,N_4504);
or U8246 (N_8246,N_4273,N_5137);
nor U8247 (N_8247,N_4663,N_4008);
and U8248 (N_8248,N_6923,N_7058);
nor U8249 (N_8249,N_7369,N_5754);
and U8250 (N_8250,N_4990,N_4769);
nor U8251 (N_8251,N_7225,N_5930);
nor U8252 (N_8252,N_4444,N_5415);
or U8253 (N_8253,N_6136,N_6137);
nand U8254 (N_8254,N_4538,N_5523);
or U8255 (N_8255,N_7736,N_7093);
and U8256 (N_8256,N_5468,N_6287);
nand U8257 (N_8257,N_5973,N_4873);
and U8258 (N_8258,N_6191,N_4945);
xnor U8259 (N_8259,N_6542,N_6334);
and U8260 (N_8260,N_7422,N_6041);
nand U8261 (N_8261,N_4480,N_6419);
nand U8262 (N_8262,N_7467,N_7803);
and U8263 (N_8263,N_6658,N_6629);
and U8264 (N_8264,N_5894,N_4773);
and U8265 (N_8265,N_4865,N_6111);
and U8266 (N_8266,N_6677,N_6497);
nor U8267 (N_8267,N_4408,N_7682);
xnor U8268 (N_8268,N_5837,N_4569);
xor U8269 (N_8269,N_5750,N_5896);
xor U8270 (N_8270,N_7930,N_4615);
nor U8271 (N_8271,N_4503,N_4530);
and U8272 (N_8272,N_5234,N_7092);
nand U8273 (N_8273,N_4078,N_4106);
nor U8274 (N_8274,N_4345,N_6135);
nand U8275 (N_8275,N_6937,N_4807);
nand U8276 (N_8276,N_7991,N_6801);
nor U8277 (N_8277,N_6595,N_5135);
xnor U8278 (N_8278,N_5027,N_6789);
nor U8279 (N_8279,N_4528,N_4952);
nor U8280 (N_8280,N_6795,N_5263);
and U8281 (N_8281,N_6295,N_7012);
and U8282 (N_8282,N_6763,N_5233);
or U8283 (N_8283,N_5505,N_7626);
or U8284 (N_8284,N_6386,N_7904);
and U8285 (N_8285,N_5128,N_5562);
and U8286 (N_8286,N_7607,N_5107);
or U8287 (N_8287,N_4331,N_4312);
xor U8288 (N_8288,N_5371,N_7960);
xor U8289 (N_8289,N_5649,N_4947);
nand U8290 (N_8290,N_5859,N_4766);
and U8291 (N_8291,N_5772,N_7022);
or U8292 (N_8292,N_4562,N_7181);
nand U8293 (N_8293,N_6593,N_5441);
and U8294 (N_8294,N_5641,N_5373);
xor U8295 (N_8295,N_6163,N_5938);
and U8296 (N_8296,N_6095,N_6473);
and U8297 (N_8297,N_4222,N_4573);
or U8298 (N_8298,N_7578,N_7943);
xnor U8299 (N_8299,N_5516,N_5888);
or U8300 (N_8300,N_5568,N_6526);
nor U8301 (N_8301,N_5352,N_5258);
and U8302 (N_8302,N_6967,N_7997);
nor U8303 (N_8303,N_5914,N_6942);
and U8304 (N_8304,N_6648,N_4991);
xnor U8305 (N_8305,N_7295,N_5404);
or U8306 (N_8306,N_7373,N_6976);
and U8307 (N_8307,N_6911,N_4354);
nand U8308 (N_8308,N_4491,N_7680);
and U8309 (N_8309,N_6365,N_4608);
or U8310 (N_8310,N_5623,N_6863);
nand U8311 (N_8311,N_6579,N_7050);
and U8312 (N_8312,N_7245,N_7456);
nor U8313 (N_8313,N_5317,N_4624);
nor U8314 (N_8314,N_7586,N_4574);
xnor U8315 (N_8315,N_7655,N_6425);
or U8316 (N_8316,N_4130,N_4629);
and U8317 (N_8317,N_4693,N_5830);
nor U8318 (N_8318,N_5558,N_4870);
and U8319 (N_8319,N_4750,N_5392);
or U8320 (N_8320,N_4522,N_7868);
xnor U8321 (N_8321,N_6074,N_6933);
or U8322 (N_8322,N_4332,N_4698);
xor U8323 (N_8323,N_7249,N_7768);
nor U8324 (N_8324,N_7567,N_7893);
nor U8325 (N_8325,N_6026,N_4801);
nor U8326 (N_8326,N_6584,N_6055);
nor U8327 (N_8327,N_4335,N_7319);
or U8328 (N_8328,N_5133,N_7721);
and U8329 (N_8329,N_6745,N_4791);
and U8330 (N_8330,N_7632,N_6458);
nor U8331 (N_8331,N_6443,N_6508);
or U8332 (N_8332,N_7239,N_7104);
nor U8333 (N_8333,N_7631,N_5536);
or U8334 (N_8334,N_5248,N_6775);
nor U8335 (N_8335,N_7832,N_7449);
xnor U8336 (N_8336,N_6384,N_5442);
and U8337 (N_8337,N_7587,N_4245);
nand U8338 (N_8338,N_5987,N_6979);
xnor U8339 (N_8339,N_7118,N_6981);
nor U8340 (N_8340,N_4027,N_6004);
or U8341 (N_8341,N_6552,N_7880);
and U8342 (N_8342,N_6633,N_6248);
nor U8343 (N_8343,N_6673,N_6950);
nand U8344 (N_8344,N_4128,N_7431);
nor U8345 (N_8345,N_4073,N_5551);
nand U8346 (N_8346,N_7708,N_7497);
or U8347 (N_8347,N_6387,N_6263);
and U8348 (N_8348,N_7221,N_4905);
nor U8349 (N_8349,N_5111,N_4440);
or U8350 (N_8350,N_6915,N_7423);
and U8351 (N_8351,N_5728,N_4889);
nand U8352 (N_8352,N_6752,N_7246);
nand U8353 (N_8353,N_4975,N_6613);
nand U8354 (N_8354,N_6943,N_4723);
nand U8355 (N_8355,N_4306,N_4936);
nor U8356 (N_8356,N_4916,N_7097);
nor U8357 (N_8357,N_6547,N_4372);
nor U8358 (N_8358,N_6277,N_4643);
nor U8359 (N_8359,N_4555,N_4547);
and U8360 (N_8360,N_6054,N_4064);
or U8361 (N_8361,N_5001,N_7333);
or U8362 (N_8362,N_7496,N_5663);
and U8363 (N_8363,N_6875,N_7679);
xnor U8364 (N_8364,N_5909,N_5249);
and U8365 (N_8365,N_6385,N_6035);
nor U8366 (N_8366,N_5105,N_4531);
nand U8367 (N_8367,N_4518,N_6082);
and U8368 (N_8368,N_7539,N_6164);
and U8369 (N_8369,N_7516,N_7131);
and U8370 (N_8370,N_4145,N_7856);
nand U8371 (N_8371,N_7622,N_6867);
nand U8372 (N_8372,N_6835,N_5819);
xor U8373 (N_8373,N_4690,N_7711);
and U8374 (N_8374,N_5677,N_4062);
nor U8375 (N_8375,N_4011,N_7363);
nand U8376 (N_8376,N_7083,N_4907);
nand U8377 (N_8377,N_4709,N_7727);
nand U8378 (N_8378,N_7800,N_4450);
and U8379 (N_8379,N_7461,N_7770);
nor U8380 (N_8380,N_7608,N_7351);
nor U8381 (N_8381,N_4044,N_7977);
nand U8382 (N_8382,N_7610,N_5069);
nor U8383 (N_8383,N_6530,N_6424);
xor U8384 (N_8384,N_7809,N_5250);
nor U8385 (N_8385,N_6048,N_5386);
xnor U8386 (N_8386,N_5918,N_4681);
xor U8387 (N_8387,N_4968,N_5019);
and U8388 (N_8388,N_5021,N_6335);
and U8389 (N_8389,N_5660,N_5443);
and U8390 (N_8390,N_4586,N_5319);
or U8391 (N_8391,N_5378,N_4327);
nor U8392 (N_8392,N_7732,N_5060);
nor U8393 (N_8393,N_4305,N_6223);
xnor U8394 (N_8394,N_5363,N_4532);
and U8395 (N_8395,N_5995,N_5327);
nand U8396 (N_8396,N_5238,N_5786);
nand U8397 (N_8397,N_4735,N_4376);
and U8398 (N_8398,N_4887,N_6102);
nand U8399 (N_8399,N_5480,N_5569);
nor U8400 (N_8400,N_7316,N_6079);
nand U8401 (N_8401,N_4834,N_6961);
nor U8402 (N_8402,N_7276,N_5897);
nand U8403 (N_8403,N_7320,N_5878);
nand U8404 (N_8404,N_6022,N_7234);
nor U8405 (N_8405,N_4088,N_5022);
nand U8406 (N_8406,N_6451,N_4728);
and U8407 (N_8407,N_4851,N_6509);
nor U8408 (N_8408,N_5984,N_7377);
and U8409 (N_8409,N_7521,N_6825);
or U8410 (N_8410,N_6370,N_6412);
and U8411 (N_8411,N_6283,N_7040);
nor U8412 (N_8412,N_5381,N_7767);
or U8413 (N_8413,N_4032,N_6105);
nand U8414 (N_8414,N_4017,N_7714);
nand U8415 (N_8415,N_5184,N_7008);
nand U8416 (N_8416,N_5891,N_5149);
or U8417 (N_8417,N_4705,N_5085);
nand U8418 (N_8418,N_4007,N_5300);
and U8419 (N_8419,N_7775,N_5796);
and U8420 (N_8420,N_4177,N_6369);
and U8421 (N_8421,N_4929,N_6156);
nand U8422 (N_8422,N_4911,N_7485);
nand U8423 (N_8423,N_5740,N_5622);
nor U8424 (N_8424,N_5518,N_4004);
nand U8425 (N_8425,N_5997,N_6852);
xnor U8426 (N_8426,N_5879,N_4508);
xor U8427 (N_8427,N_7370,N_4740);
nor U8428 (N_8428,N_4398,N_5871);
or U8429 (N_8429,N_5616,N_7474);
or U8430 (N_8430,N_5375,N_7443);
or U8431 (N_8431,N_4388,N_7148);
or U8432 (N_8432,N_7795,N_7637);
nor U8433 (N_8433,N_4466,N_6225);
nand U8434 (N_8434,N_5196,N_7099);
and U8435 (N_8435,N_5376,N_5175);
nand U8436 (N_8436,N_7900,N_7765);
and U8437 (N_8437,N_5645,N_4425);
and U8438 (N_8438,N_4119,N_7448);
or U8439 (N_8439,N_4566,N_7003);
nand U8440 (N_8440,N_5298,N_7805);
nand U8441 (N_8441,N_7349,N_4470);
or U8442 (N_8442,N_6408,N_7673);
nor U8443 (N_8443,N_4437,N_4259);
nor U8444 (N_8444,N_6594,N_5482);
nor U8445 (N_8445,N_5760,N_6993);
nor U8446 (N_8446,N_5766,N_7180);
xor U8447 (N_8447,N_5010,N_5326);
nor U8448 (N_8448,N_5881,N_5855);
nand U8449 (N_8449,N_4459,N_4443);
nor U8450 (N_8450,N_4218,N_5820);
and U8451 (N_8451,N_6192,N_7086);
or U8452 (N_8452,N_6855,N_5314);
or U8453 (N_8453,N_4136,N_6618);
nand U8454 (N_8454,N_5980,N_7460);
xor U8455 (N_8455,N_4108,N_7175);
and U8456 (N_8456,N_7866,N_4176);
and U8457 (N_8457,N_7176,N_6736);
and U8458 (N_8458,N_7688,N_7354);
nand U8459 (N_8459,N_7324,N_4321);
and U8460 (N_8460,N_5949,N_4730);
nor U8461 (N_8461,N_4726,N_7044);
or U8462 (N_8462,N_6884,N_4090);
xnor U8463 (N_8463,N_4901,N_6067);
nand U8464 (N_8464,N_7523,N_6362);
nor U8465 (N_8465,N_7400,N_7163);
or U8466 (N_8466,N_7757,N_4318);
and U8467 (N_8467,N_7327,N_7184);
or U8468 (N_8468,N_5491,N_6667);
nor U8469 (N_8469,N_6821,N_7419);
nor U8470 (N_8470,N_6607,N_4915);
and U8471 (N_8471,N_6328,N_7429);
or U8472 (N_8472,N_4804,N_5852);
or U8473 (N_8473,N_4417,N_6065);
and U8474 (N_8474,N_5038,N_5599);
nor U8475 (N_8475,N_4580,N_6053);
or U8476 (N_8476,N_5767,N_6573);
nand U8477 (N_8477,N_7671,N_7123);
and U8478 (N_8478,N_4342,N_6107);
and U8479 (N_8479,N_6214,N_6771);
or U8480 (N_8480,N_6112,N_4979);
xnor U8481 (N_8481,N_7408,N_6028);
nand U8482 (N_8482,N_4359,N_4040);
nand U8483 (N_8483,N_5213,N_6360);
nor U8484 (N_8484,N_6986,N_5704);
and U8485 (N_8485,N_7738,N_5945);
and U8486 (N_8486,N_5098,N_7228);
and U8487 (N_8487,N_5472,N_5075);
or U8488 (N_8488,N_4107,N_7487);
nand U8489 (N_8489,N_5727,N_6117);
nand U8490 (N_8490,N_7861,N_6612);
nor U8491 (N_8491,N_5325,N_5037);
or U8492 (N_8492,N_5628,N_4515);
and U8493 (N_8493,N_7666,N_6417);
nor U8494 (N_8494,N_7965,N_5322);
nor U8495 (N_8495,N_5564,N_7976);
nor U8496 (N_8496,N_5874,N_4928);
and U8497 (N_8497,N_6020,N_7686);
nor U8498 (N_8498,N_6931,N_7799);
or U8499 (N_8499,N_7678,N_5192);
nand U8500 (N_8500,N_5202,N_4213);
or U8501 (N_8501,N_5301,N_5398);
and U8502 (N_8502,N_6606,N_6298);
nand U8503 (N_8503,N_5910,N_4184);
nor U8504 (N_8504,N_4146,N_6238);
or U8505 (N_8505,N_7944,N_5601);
nor U8506 (N_8506,N_5479,N_5547);
nor U8507 (N_8507,N_6638,N_7338);
nand U8508 (N_8508,N_7648,N_7469);
nand U8509 (N_8509,N_4131,N_4856);
and U8510 (N_8510,N_5769,N_6727);
nor U8511 (N_8511,N_7617,N_7389);
nor U8512 (N_8512,N_4182,N_7196);
and U8513 (N_8513,N_5426,N_5173);
and U8514 (N_8514,N_7540,N_4161);
or U8515 (N_8515,N_5221,N_4824);
or U8516 (N_8516,N_7672,N_5849);
nor U8517 (N_8517,N_7052,N_7642);
nand U8518 (N_8518,N_4405,N_6907);
xor U8519 (N_8519,N_7042,N_5917);
and U8520 (N_8520,N_7031,N_6645);
nor U8521 (N_8521,N_6045,N_6879);
or U8522 (N_8522,N_6440,N_6255);
or U8523 (N_8523,N_5036,N_4821);
nand U8524 (N_8524,N_5676,N_7207);
nor U8525 (N_8525,N_6901,N_4967);
or U8526 (N_8526,N_7219,N_4461);
and U8527 (N_8527,N_7371,N_7401);
nand U8528 (N_8528,N_6546,N_4287);
or U8529 (N_8529,N_4370,N_7661);
or U8530 (N_8530,N_5446,N_4567);
and U8531 (N_8531,N_5634,N_5452);
and U8532 (N_8532,N_4770,N_6732);
and U8533 (N_8533,N_4534,N_6188);
nor U8534 (N_8534,N_5267,N_5035);
nand U8535 (N_8535,N_4024,N_6433);
nand U8536 (N_8536,N_5688,N_5924);
nor U8537 (N_8537,N_4018,N_4105);
xor U8538 (N_8538,N_6351,N_5965);
nor U8539 (N_8539,N_5850,N_5383);
nand U8540 (N_8540,N_4133,N_7584);
nor U8541 (N_8541,N_5364,N_4611);
and U8542 (N_8542,N_6162,N_6881);
nand U8543 (N_8543,N_4668,N_6529);
nor U8544 (N_8544,N_4551,N_7114);
nand U8545 (N_8545,N_6352,N_7399);
nand U8546 (N_8546,N_6160,N_7820);
xnor U8547 (N_8547,N_5374,N_6897);
and U8548 (N_8548,N_5887,N_6896);
or U8549 (N_8549,N_7518,N_4778);
nand U8550 (N_8550,N_6920,N_5490);
and U8551 (N_8551,N_7953,N_7932);
and U8552 (N_8552,N_4005,N_4526);
nor U8553 (N_8553,N_6837,N_4575);
and U8554 (N_8554,N_5710,N_4311);
or U8555 (N_8555,N_4496,N_4719);
and U8556 (N_8556,N_6050,N_5526);
or U8557 (N_8557,N_5606,N_6922);
nor U8558 (N_8558,N_6410,N_4514);
and U8559 (N_8559,N_6476,N_5055);
and U8560 (N_8560,N_6493,N_7649);
and U8561 (N_8561,N_5736,N_4618);
nand U8562 (N_8562,N_4243,N_7447);
nor U8563 (N_8563,N_7901,N_5771);
and U8564 (N_8564,N_4842,N_7544);
or U8565 (N_8565,N_7962,N_7082);
nand U8566 (N_8566,N_5559,N_4396);
nand U8567 (N_8567,N_4158,N_7532);
and U8568 (N_8568,N_4358,N_4558);
nand U8569 (N_8569,N_6058,N_7178);
nor U8570 (N_8570,N_7220,N_7685);
and U8571 (N_8571,N_6831,N_4971);
nand U8572 (N_8572,N_7300,N_6559);
or U8573 (N_8573,N_6989,N_7186);
nor U8574 (N_8574,N_5347,N_4277);
xor U8575 (N_8575,N_7365,N_5719);
nand U8576 (N_8576,N_4734,N_7048);
or U8577 (N_8577,N_4654,N_5372);
or U8578 (N_8578,N_6537,N_6141);
or U8579 (N_8579,N_7024,N_5230);
xnor U8580 (N_8580,N_4098,N_5826);
or U8581 (N_8581,N_7067,N_4211);
and U8582 (N_8582,N_7899,N_5651);
nand U8583 (N_8583,N_6657,N_5507);
nand U8584 (N_8584,N_5937,N_4812);
or U8585 (N_8585,N_4338,N_7433);
or U8586 (N_8586,N_6039,N_7902);
and U8587 (N_8587,N_6494,N_5836);
and U8588 (N_8588,N_5993,N_5023);
or U8589 (N_8589,N_5063,N_6142);
nor U8590 (N_8590,N_6347,N_7701);
nand U8591 (N_8591,N_7096,N_5072);
and U8592 (N_8592,N_6331,N_7226);
nand U8593 (N_8593,N_5099,N_7251);
or U8594 (N_8594,N_7223,N_5389);
nand U8595 (N_8595,N_5690,N_4042);
xor U8596 (N_8596,N_6822,N_6730);
xnor U8597 (N_8597,N_5758,N_4853);
and U8598 (N_8598,N_7950,N_4059);
nand U8599 (N_8599,N_5280,N_6025);
xnor U8600 (N_8600,N_4502,N_5410);
or U8601 (N_8601,N_4490,N_4541);
nor U8602 (N_8602,N_4825,N_5702);
and U8603 (N_8603,N_6243,N_5927);
xnor U8604 (N_8604,N_5459,N_6980);
or U8605 (N_8605,N_4696,N_7283);
or U8606 (N_8606,N_4848,N_6722);
xnor U8607 (N_8607,N_6084,N_4841);
nor U8608 (N_8608,N_5256,N_4238);
nor U8609 (N_8609,N_5394,N_6525);
and U8610 (N_8610,N_4096,N_7810);
nand U8611 (N_8611,N_6571,N_6524);
nor U8612 (N_8612,N_7939,N_7928);
nand U8613 (N_8613,N_4879,N_4230);
and U8614 (N_8614,N_6528,N_4442);
nand U8615 (N_8615,N_6038,N_4675);
nor U8616 (N_8616,N_5117,N_4383);
nand U8617 (N_8617,N_6872,N_4346);
nor U8618 (N_8618,N_6533,N_7752);
or U8619 (N_8619,N_5799,N_4464);
xor U8620 (N_8620,N_7013,N_4676);
nor U8621 (N_8621,N_4308,N_6023);
or U8622 (N_8622,N_5975,N_6659);
xnor U8623 (N_8623,N_7146,N_5164);
xor U8624 (N_8624,N_7398,N_4949);
or U8625 (N_8625,N_4006,N_5286);
and U8626 (N_8626,N_5773,N_4171);
nor U8627 (N_8627,N_7020,N_4958);
and U8628 (N_8628,N_6765,N_7368);
or U8629 (N_8629,N_4811,N_5088);
nand U8630 (N_8630,N_6216,N_5735);
nor U8631 (N_8631,N_4395,N_5700);
nand U8632 (N_8632,N_5817,N_6389);
xor U8633 (N_8633,N_5926,N_6726);
and U8634 (N_8634,N_7035,N_7876);
xor U8635 (N_8635,N_7006,N_5150);
xor U8636 (N_8636,N_5400,N_7462);
nand U8637 (N_8637,N_7478,N_7231);
and U8638 (N_8638,N_6235,N_5552);
nor U8639 (N_8639,N_6505,N_7233);
nor U8640 (N_8640,N_4249,N_5658);
nor U8641 (N_8641,N_5223,N_5496);
and U8642 (N_8642,N_4955,N_5209);
or U8643 (N_8643,N_7309,N_5777);
or U8644 (N_8644,N_7274,N_5193);
and U8645 (N_8645,N_6344,N_4478);
and U8646 (N_8646,N_6866,N_4212);
or U8647 (N_8647,N_7613,N_7126);
or U8648 (N_8648,N_5328,N_7509);
or U8649 (N_8649,N_6034,N_4781);
or U8650 (N_8650,N_5589,N_5485);
nand U8651 (N_8651,N_5985,N_7358);
nand U8652 (N_8652,N_4685,N_6381);
nand U8653 (N_8653,N_6543,N_4688);
nor U8654 (N_8654,N_4831,N_4701);
and U8655 (N_8655,N_4737,N_5116);
and U8656 (N_8656,N_7829,N_4326);
or U8657 (N_8657,N_7384,N_4209);
or U8658 (N_8658,N_7845,N_5048);
and U8659 (N_8659,N_5793,N_7933);
or U8660 (N_8660,N_5070,N_6687);
nor U8661 (N_8661,N_7865,N_5385);
or U8662 (N_8662,N_7113,N_4127);
nand U8663 (N_8663,N_4570,N_7503);
xor U8664 (N_8664,N_6760,N_4600);
or U8665 (N_8665,N_4616,N_7189);
nor U8666 (N_8666,N_7515,N_6535);
and U8667 (N_8667,N_5487,N_7142);
xor U8668 (N_8668,N_6655,N_4149);
nor U8669 (N_8669,N_7978,N_6326);
or U8670 (N_8670,N_5904,N_6532);
or U8671 (N_8671,N_5259,N_5382);
nand U8672 (N_8672,N_5293,N_7964);
and U8673 (N_8673,N_5204,N_7760);
nor U8674 (N_8674,N_6734,N_7641);
or U8675 (N_8675,N_4659,N_7468);
nand U8676 (N_8676,N_7657,N_7773);
nor U8677 (N_8677,N_7392,N_7784);
nor U8678 (N_8678,N_7315,N_6338);
nand U8679 (N_8679,N_4179,N_5229);
and U8680 (N_8680,N_4867,N_4188);
or U8681 (N_8681,N_6487,N_4930);
xnor U8682 (N_8682,N_5231,N_6781);
and U8683 (N_8683,N_6877,N_6415);
nand U8684 (N_8684,N_6725,N_5620);
nand U8685 (N_8685,N_4956,N_7243);
nand U8686 (N_8686,N_4102,N_6027);
and U8687 (N_8687,N_5104,N_6891);
and U8688 (N_8688,N_4095,N_4639);
xor U8689 (N_8689,N_6008,N_4267);
or U8690 (N_8690,N_7739,N_6145);
nand U8691 (N_8691,N_6060,N_6206);
and U8692 (N_8692,N_5207,N_7438);
xor U8693 (N_8693,N_4343,N_4509);
and U8694 (N_8694,N_7506,N_6405);
and U8695 (N_8695,N_5211,N_7885);
and U8696 (N_8696,N_7201,N_4430);
and U8697 (N_8697,N_4075,N_4733);
nand U8698 (N_8698,N_6605,N_5310);
nor U8699 (N_8699,N_7137,N_5168);
nand U8700 (N_8700,N_5578,N_6842);
or U8701 (N_8701,N_6522,N_6108);
or U8702 (N_8702,N_4571,N_7080);
xnor U8703 (N_8703,N_4579,N_7763);
xor U8704 (N_8704,N_5585,N_6849);
nor U8705 (N_8705,N_4234,N_4274);
xor U8706 (N_8706,N_5545,N_7229);
and U8707 (N_8707,N_6581,N_5304);
or U8708 (N_8708,N_6557,N_7288);
and U8709 (N_8709,N_7592,N_4988);
xor U8710 (N_8710,N_7664,N_6181);
nand U8711 (N_8711,N_6951,N_5465);
or U8712 (N_8712,N_5721,N_7410);
and U8713 (N_8713,N_7154,N_4498);
and U8714 (N_8714,N_7827,N_6109);
and U8715 (N_8715,N_4112,N_4009);
or U8716 (N_8716,N_5781,N_5946);
nor U8717 (N_8717,N_4416,N_4585);
nor U8718 (N_8718,N_5579,N_4068);
xnor U8719 (N_8719,N_7149,N_7143);
xnor U8720 (N_8720,N_4113,N_7260);
nand U8721 (N_8721,N_6454,N_7985);
and U8722 (N_8722,N_6834,N_5605);
xnor U8723 (N_8723,N_4640,N_4664);
nor U8724 (N_8724,N_6969,N_6106);
and U8725 (N_8725,N_5447,N_4536);
nand U8726 (N_8726,N_4224,N_4642);
or U8727 (N_8727,N_4471,N_7758);
and U8728 (N_8728,N_4151,N_5635);
and U8729 (N_8729,N_7611,N_7317);
nor U8730 (N_8730,N_6892,N_6005);
or U8731 (N_8731,N_5575,N_5549);
xor U8732 (N_8732,N_4246,N_5543);
or U8733 (N_8733,N_7279,N_7884);
nor U8734 (N_8734,N_5939,N_7574);
nand U8735 (N_8735,N_6800,N_4749);
nor U8736 (N_8736,N_6413,N_4019);
or U8737 (N_8737,N_7329,N_6492);
and U8738 (N_8738,N_4293,N_6231);
nand U8739 (N_8739,N_5739,N_7761);
or U8740 (N_8740,N_4072,N_7797);
or U8741 (N_8741,N_4140,N_6699);
nor U8742 (N_8742,N_7205,N_4307);
nand U8743 (N_8743,N_5254,N_6523);
xnor U8744 (N_8744,N_7925,N_4265);
and U8745 (N_8745,N_7624,N_4758);
or U8746 (N_8746,N_5524,N_5706);
nand U8747 (N_8747,N_6827,N_6118);
nor U8748 (N_8748,N_6983,N_4160);
or U8749 (N_8749,N_5816,N_5839);
nor U8750 (N_8750,N_5039,N_6816);
or U8751 (N_8751,N_5932,N_5182);
or U8752 (N_8752,N_7597,N_6224);
nor U8753 (N_8753,N_7066,N_4985);
nor U8754 (N_8754,N_6286,N_7594);
nand U8755 (N_8755,N_5186,N_5440);
and U8756 (N_8756,N_6723,N_5698);
nor U8757 (N_8757,N_6829,N_7454);
nand U8758 (N_8758,N_4795,N_5451);
nand U8759 (N_8759,N_5743,N_5138);
nor U8760 (N_8760,N_7915,N_5659);
nand U8761 (N_8761,N_6154,N_7150);
or U8762 (N_8762,N_6480,N_5948);
nor U8763 (N_8763,N_4666,N_7078);
and U8764 (N_8764,N_6218,N_5041);
or U8765 (N_8765,N_7749,N_6847);
nor U8766 (N_8766,N_5503,N_7345);
or U8767 (N_8767,N_4609,N_7984);
and U8768 (N_8768,N_7566,N_7822);
xor U8769 (N_8769,N_5950,N_6649);
xor U8770 (N_8770,N_5619,N_4025);
nand U8771 (N_8771,N_4835,N_4204);
or U8772 (N_8772,N_4772,N_5809);
or U8773 (N_8773,N_4137,N_5812);
or U8774 (N_8774,N_5066,N_6174);
nand U8775 (N_8775,N_7390,N_4481);
and U8776 (N_8776,N_5848,N_6538);
or U8777 (N_8777,N_6985,N_5228);
and U8778 (N_8778,N_7062,N_5666);
nor U8779 (N_8779,N_5808,N_7439);
nand U8780 (N_8780,N_4282,N_5428);
or U8781 (N_8781,N_6220,N_7621);
xnor U8782 (N_8782,N_7299,N_6741);
nor U8783 (N_8783,N_4050,N_7609);
or U8784 (N_8784,N_4843,N_4485);
nand U8785 (N_8785,N_4546,N_7643);
nor U8786 (N_8786,N_6211,N_7426);
nor U8787 (N_8787,N_5349,N_7101);
nor U8788 (N_8788,N_5077,N_7197);
or U8789 (N_8789,N_6061,N_5043);
or U8790 (N_8790,N_4404,N_5892);
nand U8791 (N_8791,N_4519,N_4239);
nand U8792 (N_8792,N_6828,N_4784);
and U8793 (N_8793,N_4215,N_5668);
xor U8794 (N_8794,N_4284,N_6043);
nand U8795 (N_8795,N_4315,N_7167);
and U8796 (N_8796,N_5643,N_5051);
nor U8797 (N_8797,N_6390,N_7051);
nand U8798 (N_8798,N_4301,N_7341);
nand U8799 (N_8799,N_6407,N_7558);
nand U8800 (N_8800,N_7891,N_5738);
nor U8801 (N_8801,N_6780,N_6183);
or U8802 (N_8802,N_4798,N_7862);
and U8803 (N_8803,N_5593,N_4082);
or U8804 (N_8804,N_7297,N_7730);
and U8805 (N_8805,N_7847,N_7109);
nor U8806 (N_8806,N_7938,N_6660);
nand U8807 (N_8807,N_7428,N_7886);
or U8808 (N_8808,N_5832,N_4366);
nand U8809 (N_8809,N_6545,N_5004);
xor U8810 (N_8810,N_5174,N_5813);
nand U8811 (N_8811,N_6823,N_4296);
or U8812 (N_8812,N_7087,N_4330);
xor U8813 (N_8813,N_5664,N_6275);
and U8814 (N_8814,N_5336,N_4753);
nand U8815 (N_8815,N_6797,N_4599);
or U8816 (N_8816,N_5194,N_7920);
or U8817 (N_8817,N_4297,N_5109);
nor U8818 (N_8818,N_7911,N_5445);
or U8819 (N_8819,N_6832,N_6278);
or U8820 (N_8820,N_5102,N_6544);
nand U8821 (N_8821,N_4167,N_5411);
and U8822 (N_8822,N_6482,N_4511);
and U8823 (N_8823,N_4844,N_7424);
nor U8824 (N_8824,N_7772,N_7640);
and U8825 (N_8825,N_4356,N_5899);
nor U8826 (N_8826,N_6282,N_6303);
or U8827 (N_8827,N_4187,N_4438);
or U8828 (N_8828,N_4118,N_6450);
nand U8829 (N_8829,N_5476,N_7596);
nor U8830 (N_8830,N_7380,N_4435);
or U8831 (N_8831,N_5499,N_6104);
nand U8832 (N_8832,N_6032,N_5463);
or U8833 (N_8833,N_5513,N_7628);
or U8834 (N_8834,N_4029,N_4623);
nand U8835 (N_8835,N_7480,N_4612);
and U8836 (N_8836,N_6468,N_4605);
and U8837 (N_8837,N_4288,N_5139);
nor U8838 (N_8838,N_6076,N_6330);
or U8839 (N_8839,N_5646,N_5044);
nor U8840 (N_8840,N_4104,N_4494);
or U8841 (N_8841,N_6748,N_5573);
nand U8842 (N_8842,N_7413,N_6941);
nand U8843 (N_8843,N_7185,N_5763);
nor U8844 (N_8844,N_6116,N_6549);
and U8845 (N_8845,N_6910,N_5818);
nor U8846 (N_8846,N_5106,N_5947);
nor U8847 (N_8847,N_4755,N_4644);
nor U8848 (N_8848,N_6854,N_7111);
and U8849 (N_8849,N_5877,N_6554);
or U8850 (N_8850,N_7425,N_4746);
xnor U8851 (N_8851,N_6754,N_6514);
or U8852 (N_8852,N_7956,N_7106);
nor U8853 (N_8853,N_7053,N_6380);
nand U8854 (N_8854,N_6179,N_7045);
xor U8855 (N_8855,N_4923,N_6322);
and U8856 (N_8856,N_6906,N_4482);
xor U8857 (N_8857,N_4933,N_4071);
nand U8858 (N_8858,N_6228,N_6886);
xor U8859 (N_8859,N_6740,N_6376);
and U8860 (N_8860,N_4762,N_5172);
nor U8861 (N_8861,N_4077,N_4402);
or U8862 (N_8862,N_5835,N_4902);
xor U8863 (N_8863,N_4721,N_4512);
and U8864 (N_8864,N_4016,N_6802);
nand U8865 (N_8865,N_4813,N_5913);
and U8866 (N_8866,N_4576,N_6343);
and U8867 (N_8867,N_7135,N_6462);
nor U8868 (N_8868,N_4170,N_4375);
nand U8869 (N_8869,N_5989,N_7879);
nor U8870 (N_8870,N_7555,N_4950);
nand U8871 (N_8871,N_7998,N_4954);
and U8872 (N_8872,N_5414,N_5951);
and U8873 (N_8873,N_6833,N_5431);
or U8874 (N_8874,N_5297,N_6096);
or U8875 (N_8875,N_6799,N_6870);
nor U8876 (N_8876,N_4587,N_5288);
nor U8877 (N_8877,N_6044,N_6636);
nand U8878 (N_8878,N_7286,N_4201);
xor U8879 (N_8879,N_4156,N_4557);
or U8880 (N_8880,N_4254,N_5421);
nor U8881 (N_8881,N_6792,N_6155);
and U8882 (N_8882,N_6240,N_4860);
or U8883 (N_8883,N_4553,N_6046);
or U8884 (N_8884,N_4671,N_6373);
and U8885 (N_8885,N_4424,N_6251);
and U8886 (N_8886,N_7703,N_7883);
nor U8887 (N_8887,N_5065,N_7614);
nor U8888 (N_8888,N_4981,N_4217);
or U8889 (N_8889,N_6253,N_7482);
or U8890 (N_8890,N_5699,N_4420);
nor U8891 (N_8891,N_4839,N_5588);
and U8892 (N_8892,N_5638,N_6168);
xnor U8893 (N_8893,N_5206,N_7210);
and U8894 (N_8894,N_4240,N_4268);
and U8895 (N_8895,N_4002,N_5017);
nand U8896 (N_8896,N_6749,N_5683);
xor U8897 (N_8897,N_5097,N_5592);
or U8898 (N_8898,N_4115,N_7553);
nand U8899 (N_8899,N_5717,N_5198);
or U8900 (N_8900,N_6456,N_6688);
nor U8901 (N_8901,N_5863,N_5994);
or U8902 (N_8902,N_6956,N_6959);
nor U8903 (N_8903,N_6826,N_5996);
nand U8904 (N_8904,N_6599,N_7084);
or U8905 (N_8905,N_7903,N_5765);
or U8906 (N_8906,N_5000,N_5145);
and U8907 (N_8907,N_5032,N_7929);
and U8908 (N_8908,N_5200,N_6790);
nand U8909 (N_8909,N_6813,N_7307);
nor U8910 (N_8910,N_6994,N_6404);
and U8911 (N_8911,N_4799,N_5554);
nand U8912 (N_8912,N_7004,N_7605);
or U8913 (N_8913,N_6731,N_5607);
or U8914 (N_8914,N_7718,N_5083);
nor U8915 (N_8915,N_5885,N_5071);
nand U8916 (N_8916,N_5615,N_6936);
nor U8917 (N_8917,N_5709,N_7191);
nor U8918 (N_8918,N_6368,N_6444);
or U8919 (N_8919,N_7183,N_4888);
nor U8920 (N_8920,N_4669,N_4776);
and U8921 (N_8921,N_7835,N_7931);
or U8922 (N_8922,N_6262,N_7870);
nand U8923 (N_8923,N_4320,N_6764);
nor U8924 (N_8924,N_4381,N_5006);
nand U8925 (N_8925,N_6345,N_6747);
xor U8926 (N_8926,N_6305,N_5435);
or U8927 (N_8927,N_4499,N_7391);
and U8928 (N_8928,N_6341,N_5550);
and U8929 (N_8929,N_4763,N_6083);
and U8930 (N_8930,N_7188,N_4595);
xor U8931 (N_8931,N_6324,N_4066);
and U8932 (N_8932,N_4589,N_5281);
and U8933 (N_8933,N_5464,N_7689);
or U8934 (N_8934,N_6361,N_7466);
or U8935 (N_8935,N_4079,N_6196);
or U8936 (N_8936,N_5031,N_7887);
and U8937 (N_8937,N_6320,N_7572);
nand U8938 (N_8938,N_7743,N_6213);
nor U8939 (N_8939,N_4389,N_4242);
nor U8940 (N_8940,N_6406,N_4622);
xnor U8941 (N_8941,N_5225,N_6758);
and U8942 (N_8942,N_4076,N_5295);
nor U8943 (N_8943,N_7382,N_6683);
nand U8944 (N_8944,N_4303,N_6428);
nand U8945 (N_8945,N_5477,N_4436);
nand U8946 (N_8946,N_7108,N_6290);
and U8947 (N_8947,N_4148,N_4092);
xor U8948 (N_8948,N_6739,N_6656);
and U8949 (N_8949,N_4362,N_4694);
nand U8950 (N_8950,N_7565,N_5705);
or U8951 (N_8951,N_7560,N_5675);
or U8952 (N_8952,N_5444,N_4081);
nor U8953 (N_8953,N_4926,N_5334);
nand U8954 (N_8954,N_6300,N_6435);
nor U8955 (N_8955,N_6682,N_7494);
nor U8956 (N_8956,N_4552,N_7282);
nor U8957 (N_8957,N_4015,N_4120);
and U8958 (N_8958,N_4797,N_4626);
nand U8959 (N_8959,N_6469,N_5742);
nor U8960 (N_8960,N_6477,N_6960);
nor U8961 (N_8961,N_5030,N_5205);
and U8962 (N_8962,N_7707,N_7301);
xnor U8963 (N_8963,N_7041,N_5954);
nand U8964 (N_8964,N_5500,N_4854);
nor U8965 (N_8965,N_5942,N_7125);
and U8966 (N_8966,N_6899,N_7107);
nand U8967 (N_8967,N_6988,N_6952);
nand U8968 (N_8968,N_6485,N_5292);
nand U8969 (N_8969,N_6641,N_4584);
and U8970 (N_8970,N_7616,N_7259);
or U8971 (N_8971,N_4310,N_5574);
nor U8972 (N_8972,N_5076,N_4074);
nand U8973 (N_8973,N_5586,N_5656);
xor U8974 (N_8974,N_5061,N_7266);
nand U8975 (N_8975,N_6133,N_5320);
nand U8976 (N_8976,N_7836,N_6563);
nor U8977 (N_8977,N_6264,N_6449);
nand U8978 (N_8978,N_7556,N_6807);
nor U8979 (N_8979,N_6249,N_5576);
and U8980 (N_8980,N_7036,N_7357);
nand U8981 (N_8981,N_6210,N_6153);
and U8982 (N_8982,N_7973,N_4328);
or U8983 (N_8983,N_4178,N_6171);
nand U8984 (N_8984,N_4891,N_7335);
or U8985 (N_8985,N_4892,N_4921);
and U8986 (N_8986,N_7855,N_5759);
xor U8987 (N_8987,N_6919,N_5695);
or U8988 (N_8988,N_4493,N_5794);
nor U8989 (N_8989,N_6474,N_7023);
and U8990 (N_8990,N_6583,N_6818);
nand U8991 (N_8991,N_4159,N_7755);
and U8992 (N_8992,N_4913,N_7495);
nor U8993 (N_8993,N_7252,N_5113);
nor U8994 (N_8994,N_7871,N_7917);
and U8995 (N_8995,N_6743,N_4809);
and U8996 (N_8996,N_5040,N_4324);
and U8997 (N_8997,N_4426,N_6695);
or U8998 (N_8998,N_4469,N_6488);
xnor U8999 (N_8999,N_4745,N_4409);
and U9000 (N_9000,N_7961,N_6787);
nor U9001 (N_9001,N_7273,N_5876);
or U9002 (N_9002,N_5348,N_4904);
xor U9003 (N_9003,N_6513,N_4260);
nor U9004 (N_9004,N_6114,N_6592);
nor U9005 (N_9005,N_6561,N_5057);
nand U9006 (N_9006,N_6340,N_5637);
nor U9007 (N_9007,N_6770,N_7638);
nor U9008 (N_9008,N_7254,N_7174);
nor U9009 (N_9009,N_7100,N_5457);
nand U9010 (N_9010,N_6694,N_5242);
and U9011 (N_9011,N_7311,N_6713);
and U9012 (N_9012,N_4298,N_5227);
nand U9013 (N_9013,N_4166,N_4604);
or U9014 (N_9014,N_6437,N_4818);
nand U9015 (N_9015,N_4602,N_4080);
nand U9016 (N_9016,N_7791,N_4110);
and U9017 (N_9017,N_7937,N_6087);
nand U9018 (N_9018,N_5408,N_4295);
nand U9019 (N_9019,N_7811,N_6503);
nor U9020 (N_9020,N_7038,N_6189);
nor U9021 (N_9021,N_6299,N_4827);
xor U9022 (N_9022,N_7446,N_6186);
nor U9023 (N_9023,N_7547,N_4715);
or U9024 (N_9024,N_4980,N_6597);
xor U9025 (N_9025,N_4200,N_6778);
or U9026 (N_9026,N_5271,N_7824);
or U9027 (N_9027,N_4881,N_4053);
and U9028 (N_9028,N_6000,N_4141);
xor U9029 (N_9029,N_5413,N_7542);
nor U9030 (N_9030,N_6144,N_4210);
nor U9031 (N_9031,N_6031,N_6811);
nor U9032 (N_9032,N_4665,N_4987);
nor U9033 (N_9033,N_5449,N_4228);
xor U9034 (N_9034,N_7813,N_4194);
and U9035 (N_9035,N_6591,N_4035);
or U9036 (N_9036,N_4419,N_5806);
and U9037 (N_9037,N_7284,N_4995);
or U9038 (N_9038,N_4765,N_7550);
and U9039 (N_9039,N_6720,N_7630);
xor U9040 (N_9040,N_4173,N_5339);
or U9041 (N_9041,N_6916,N_7662);
nor U9042 (N_9042,N_6182,N_5911);
nand U9043 (N_9043,N_6686,N_5279);
nand U9044 (N_9044,N_7079,N_7947);
or U9045 (N_9045,N_4592,N_4229);
nand U9046 (N_9046,N_7941,N_6394);
xnor U9047 (N_9047,N_6401,N_5889);
nor U9048 (N_9048,N_6954,N_5714);
and U9049 (N_9049,N_7451,N_4501);
or U9050 (N_9050,N_7388,N_4236);
nor U9051 (N_9051,N_7852,N_4191);
nand U9052 (N_9052,N_4817,N_7043);
and U9053 (N_9053,N_6489,N_7599);
xnor U9054 (N_9054,N_6851,N_5921);
nand U9055 (N_9055,N_5708,N_6276);
or U9056 (N_9056,N_4023,N_4815);
or U9057 (N_9057,N_7132,N_6560);
and U9058 (N_9058,N_4061,N_7285);
or U9059 (N_9059,N_5438,N_5343);
xor U9060 (N_9060,N_7806,N_4169);
nor U9061 (N_9061,N_4290,N_5045);
nand U9062 (N_9062,N_4731,N_5685);
nor U9063 (N_9063,N_4561,N_6623);
nand U9064 (N_9064,N_7393,N_6784);
or U9065 (N_9065,N_5395,N_4154);
or U9066 (N_9066,N_7667,N_4692);
xor U9067 (N_9067,N_7881,N_5716);
xnor U9068 (N_9068,N_7061,N_4394);
or U9069 (N_9069,N_6364,N_7488);
nand U9070 (N_9070,N_5388,N_6887);
and U9071 (N_9071,N_4418,N_6042);
nor U9072 (N_9072,N_4683,N_6148);
nor U9073 (N_9073,N_4695,N_6871);
nor U9074 (N_9074,N_6353,N_6572);
and U9075 (N_9075,N_4658,N_7427);
and U9076 (N_9076,N_4401,N_4189);
nand U9077 (N_9077,N_4316,N_6982);
xnor U9078 (N_9078,N_6958,N_5252);
or U9079 (N_9079,N_4322,N_7945);
and U9080 (N_9080,N_6093,N_6372);
or U9081 (N_9081,N_5761,N_7133);
nand U9082 (N_9082,N_4407,N_4434);
nor U9083 (N_9083,N_5180,N_6336);
or U9084 (N_9084,N_4941,N_6319);
xnor U9085 (N_9085,N_7909,N_4012);
nand U9086 (N_9086,N_6219,N_7416);
and U9087 (N_9087,N_7395,N_4462);
and U9088 (N_9088,N_6601,N_5340);
xnor U9089 (N_9089,N_5311,N_4542);
nor U9090 (N_9090,N_5846,N_6429);
or U9091 (N_9091,N_7330,N_5453);
nor U9092 (N_9092,N_7305,N_6698);
nand U9093 (N_9093,N_5825,N_7409);
or U9094 (N_9094,N_6644,N_6321);
or U9095 (N_9095,N_5529,N_6690);
nor U9096 (N_9096,N_4645,N_6865);
nand U9097 (N_9097,N_4894,N_7552);
and U9098 (N_9098,N_7145,N_7077);
and U9099 (N_9099,N_5670,N_7014);
and U9100 (N_9100,N_4488,N_4957);
nand U9101 (N_9101,N_5399,N_4344);
nand U9102 (N_9102,N_4026,N_6755);
nand U9103 (N_9103,N_4124,N_4351);
or U9104 (N_9104,N_5847,N_4619);
xor U9105 (N_9105,N_4577,N_5454);
nand U9106 (N_9106,N_4056,N_7366);
nor U9107 (N_9107,N_4261,N_6120);
nand U9108 (N_9108,N_6463,N_4864);
and U9109 (N_9109,N_5341,N_7589);
nor U9110 (N_9110,N_7212,N_5687);
or U9111 (N_9111,N_4452,N_5302);
or U9112 (N_9112,N_6869,N_6925);
nor U9113 (N_9113,N_6712,N_5594);
nand U9114 (N_9114,N_6692,N_4010);
xnor U9115 (N_9115,N_5264,N_5944);
and U9116 (N_9116,N_7982,N_7634);
nand U9117 (N_9117,N_7501,N_7522);
nand U9118 (N_9118,N_5284,N_4181);
and U9119 (N_9119,N_7802,N_6230);
or U9120 (N_9120,N_4830,N_7140);
and U9121 (N_9121,N_4768,N_7147);
nand U9122 (N_9122,N_4914,N_7729);
or U9123 (N_9123,N_7247,N_4621);
xnor U9124 (N_9124,N_7236,N_4729);
xor U9125 (N_9125,N_7290,N_7352);
and U9126 (N_9126,N_7161,N_6070);
nand U9127 (N_9127,N_5560,N_4400);
or U9128 (N_9128,N_6701,N_5838);
xor U9129 (N_9129,N_4634,N_7313);
and U9130 (N_9130,N_6466,N_7794);
nor U9131 (N_9131,N_4572,N_7737);
nand U9132 (N_9132,N_4083,N_7411);
nand U9133 (N_9133,N_7244,N_5448);
nor U9134 (N_9134,N_4651,N_6578);
or U9135 (N_9135,N_7922,N_6081);
or U9136 (N_9136,N_5701,N_4682);
xnor U9137 (N_9137,N_5541,N_5357);
nand U9138 (N_9138,N_5266,N_5843);
nor U9139 (N_9139,N_7987,N_4114);
nand U9140 (N_9140,N_4034,N_7182);
and U9141 (N_9141,N_4231,N_6890);
nand U9142 (N_9142,N_5669,N_4638);
nand U9143 (N_9143,N_7646,N_7242);
or U9144 (N_9144,N_7924,N_4898);
or U9145 (N_9145,N_5901,N_6702);
or U9146 (N_9146,N_4353,N_7312);
and U9147 (N_9147,N_4661,N_7206);
and U9148 (N_9148,N_4379,N_7010);
nor U9149 (N_9149,N_4691,N_5833);
or U9150 (N_9150,N_5905,N_4855);
or U9151 (N_9151,N_5026,N_7293);
nor U9152 (N_9152,N_6921,N_6090);
nor U9153 (N_9153,N_7850,N_6555);
nand U9154 (N_9154,N_4054,N_7988);
and U9155 (N_9155,N_7533,N_7085);
nor U9156 (N_9156,N_6737,N_4474);
or U9157 (N_9157,N_4754,N_4869);
nor U9158 (N_9158,N_7321,N_7081);
and U9159 (N_9159,N_7379,N_7152);
nor U9160 (N_9160,N_6323,N_4820);
nand U9161 (N_9161,N_7706,N_6966);
or U9162 (N_9162,N_6520,N_7790);
or U9163 (N_9163,N_6292,N_4447);
and U9164 (N_9164,N_5792,N_6588);
and U9165 (N_9165,N_5474,N_4961);
nand U9166 (N_9166,N_5384,N_6254);
nand U9167 (N_9167,N_4861,N_4031);
nand U9168 (N_9168,N_4185,N_5290);
nand U9169 (N_9169,N_5572,N_5922);
or U9170 (N_9170,N_5864,N_5920);
nor U9171 (N_9171,N_7783,N_7619);
nor U9172 (N_9172,N_4960,N_6759);
or U9173 (N_9173,N_6676,N_4885);
and U9174 (N_9174,N_7750,N_7788);
nand U9175 (N_9175,N_6092,N_5287);
nand U9176 (N_9176,N_7561,N_5653);
nand U9177 (N_9177,N_4510,N_7069);
or U9178 (N_9178,N_4122,N_4944);
xnor U9179 (N_9179,N_7908,N_6175);
or U9180 (N_9180,N_7177,N_4742);
xor U9181 (N_9181,N_5527,N_5624);
and U9182 (N_9182,N_5417,N_7888);
or U9183 (N_9183,N_7374,N_6926);
and U9184 (N_9184,N_4142,N_4686);
or U9185 (N_9185,N_7656,N_6453);
nand U9186 (N_9186,N_4196,N_7216);
nor U9187 (N_9187,N_6129,N_6426);
or U9188 (N_9188,N_7238,N_7825);
nor U9189 (N_9189,N_6719,N_7860);
xnor U9190 (N_9190,N_6442,N_6333);
nand U9191 (N_9191,N_7227,N_4822);
or U9192 (N_9192,N_5240,N_6889);
or U9193 (N_9193,N_5329,N_4662);
nand U9194 (N_9194,N_5531,N_7089);
nor U9195 (N_9195,N_4593,N_6195);
nand U9196 (N_9196,N_5217,N_7278);
nand U9197 (N_9197,N_4109,N_7074);
nor U9198 (N_9198,N_4103,N_4221);
and U9199 (N_9199,N_6608,N_6256);
nor U9200 (N_9200,N_4847,N_4055);
and U9201 (N_9201,N_5003,N_4390);
nand U9202 (N_9202,N_7777,N_5553);
or U9203 (N_9203,N_5842,N_5618);
nand U9204 (N_9204,N_5062,N_7972);
nor U9205 (N_9205,N_6245,N_6208);
xor U9206 (N_9206,N_5522,N_7778);
and U9207 (N_9207,N_6930,N_6475);
and U9208 (N_9208,N_7514,N_4337);
xor U9209 (N_9209,N_5402,N_6001);
or U9210 (N_9210,N_5246,N_6269);
or U9211 (N_9211,N_5958,N_7430);
nor U9212 (N_9212,N_7435,N_5405);
nand U9213 (N_9213,N_5191,N_7115);
nand U9214 (N_9214,N_7579,N_6377);
xnor U9215 (N_9215,N_5694,N_7989);
nand U9216 (N_9216,N_7187,N_5303);
or U9217 (N_9217,N_6803,N_6502);
nor U9218 (N_9218,N_4506,N_7217);
nand U9219 (N_9219,N_4833,N_6198);
nor U9220 (N_9220,N_7491,N_6997);
or U9221 (N_9221,N_7873,N_5439);
nor U9222 (N_9222,N_6422,N_5166);
and U9223 (N_9223,N_7208,N_4712);
nor U9224 (N_9224,N_7072,N_7404);
nand U9225 (N_9225,N_5693,N_4630);
nand U9226 (N_9226,N_7633,N_4777);
or U9227 (N_9227,N_5216,N_4155);
nor U9228 (N_9228,N_7725,N_7159);
nand U9229 (N_9229,N_6318,N_6068);
xnor U9230 (N_9230,N_4060,N_4606);
xnor U9231 (N_9231,N_4940,N_5580);
and U9232 (N_9232,N_4247,N_7766);
and U9233 (N_9233,N_7016,N_7980);
or U9234 (N_9234,N_4816,N_7789);
or U9235 (N_9235,N_5697,N_4673);
nor U9236 (N_9236,N_7595,N_5081);
or U9237 (N_9237,N_5469,N_5880);
nand U9238 (N_9238,N_5613,N_4387);
or U9239 (N_9239,N_7748,N_6565);
nor U9240 (N_9240,N_5158,N_6089);
nand U9241 (N_9241,N_4601,N_7002);
and U9242 (N_9242,N_7194,N_5556);
nor U9243 (N_9243,N_7780,N_5730);
nor U9244 (N_9244,N_7179,N_5870);
nor U9245 (N_9245,N_5805,N_7715);
nand U9246 (N_9246,N_7171,N_6738);
nand U9247 (N_9247,N_4724,N_7457);
and U9248 (N_9248,N_6271,N_4085);
or U9249 (N_9249,N_7262,N_4917);
nor U9250 (N_9250,N_5566,N_7669);
nor U9251 (N_9251,N_6392,N_7472);
nand U9252 (N_9252,N_4281,N_7453);
or U9253 (N_9253,N_7872,N_5047);
and U9254 (N_9254,N_5563,N_4472);
and U9255 (N_9255,N_6710,N_6878);
nor U9256 (N_9256,N_6949,N_6628);
nand U9257 (N_9257,N_6815,N_6126);
xnor U9258 (N_9258,N_6086,N_5530);
or U9259 (N_9259,N_7691,N_6709);
or U9260 (N_9260,N_7442,N_5080);
nand U9261 (N_9261,N_7601,N_7088);
and U9262 (N_9262,N_6938,N_6367);
nor U9263 (N_9263,N_4710,N_7562);
nand U9264 (N_9264,N_4043,N_6707);
or U9265 (N_9265,N_4684,N_4527);
or U9266 (N_9266,N_4492,N_4186);
nor U9267 (N_9267,N_4646,N_7222);
nor U9268 (N_9268,N_7475,N_4299);
and U9269 (N_9269,N_7905,N_5929);
nor U9270 (N_9270,N_4703,N_5718);
nor U9271 (N_9271,N_6432,N_7971);
nand U9272 (N_9272,N_6810,N_6486);
nor U9273 (N_9273,N_4744,N_6308);
xor U9274 (N_9274,N_7600,N_7328);
and U9275 (N_9275,N_6841,N_6471);
xor U9276 (N_9276,N_6598,N_4702);
or U9277 (N_9277,N_6970,N_4441);
nor U9278 (N_9278,N_5203,N_6495);
nand U9279 (N_9279,N_4964,N_5822);
and U9280 (N_9280,N_6363,N_6169);
nor U9281 (N_9281,N_6346,N_6661);
or U9282 (N_9282,N_7033,N_7756);
nand U9283 (N_9283,N_6804,N_7935);
and U9284 (N_9284,N_5068,N_4505);
and U9285 (N_9285,N_7385,N_7340);
nor U9286 (N_9286,N_6642,N_4455);
and U9287 (N_9287,N_4610,N_5955);
nand U9288 (N_9288,N_4292,N_7049);
and U9289 (N_9289,N_7751,N_4038);
or U9290 (N_9290,N_4743,N_6498);
nand U9291 (N_9291,N_4895,N_7582);
and U9292 (N_9292,N_4164,N_4523);
nor U9293 (N_9293,N_6512,N_5935);
nor U9294 (N_9294,N_4421,N_5094);
and U9295 (N_9295,N_7954,N_7898);
nand U9296 (N_9296,N_5377,N_4764);
nand U9297 (N_9297,N_6427,N_7863);
and U9298 (N_9298,N_5125,N_5657);
nand U9299 (N_9299,N_4760,N_7498);
or U9300 (N_9300,N_5548,N_5757);
xor U9301 (N_9301,N_6779,N_7683);
xnor U9302 (N_9302,N_6507,N_5644);
and U9303 (N_9303,N_4978,N_7375);
xnor U9304 (N_9304,N_5956,N_5626);
nand U9305 (N_9305,N_6274,N_4874);
nor U9306 (N_9306,N_6806,N_7493);
and U9307 (N_9307,N_4906,N_7660);
and U9308 (N_9308,N_5437,N_7826);
or U9309 (N_9309,N_5791,N_6769);
and U9310 (N_9310,N_7554,N_4465);
and U9311 (N_9311,N_4890,N_5131);
xnor U9312 (N_9312,N_4525,N_6908);
or U9313 (N_9313,N_6962,N_5612);
or U9314 (N_9314,N_5461,N_6349);
and U9315 (N_9315,N_5222,N_6237);
nor U9316 (N_9316,N_6059,N_6998);
nor U9317 (N_9317,N_5475,N_6423);
nand U9318 (N_9318,N_5652,N_7864);
nor U9319 (N_9319,N_6809,N_5515);
and U9320 (N_9320,N_5115,N_5253);
nand U9321 (N_9321,N_4620,N_6678);
or U9322 (N_9322,N_5762,N_7534);
nand U9323 (N_9323,N_6197,N_4270);
nand U9324 (N_9324,N_5632,N_4796);
and U9325 (N_9325,N_6637,N_6539);
and U9326 (N_9326,N_4877,N_6388);
nor U9327 (N_9327,N_6172,N_6717);
nor U9328 (N_9328,N_4937,N_7248);
nand U9329 (N_9329,N_4722,N_6684);
nand U9330 (N_9330,N_6817,N_4829);
nor U9331 (N_9331,N_5814,N_7999);
and U9332 (N_9332,N_7712,N_4207);
nor U9333 (N_9333,N_7403,N_7627);
xor U9334 (N_9334,N_5387,N_6696);
nand U9335 (N_9335,N_5255,N_5154);
nand U9336 (N_9336,N_5733,N_6382);
nand U9337 (N_9337,N_5854,N_6991);
xor U9338 (N_9338,N_5581,N_7009);
and U9339 (N_9339,N_7255,N_7551);
and U9340 (N_9340,N_5873,N_4300);
and U9341 (N_9341,N_6693,N_6972);
nand U9342 (N_9342,N_7158,N_5178);
nor U9343 (N_9343,N_5011,N_7500);
nor U9344 (N_9344,N_4989,N_5597);
nor U9345 (N_9345,N_5857,N_7687);
nand U9346 (N_9346,N_7169,N_5108);
or U9347 (N_9347,N_4837,N_4687);
nand U9348 (N_9348,N_5591,N_6073);
nor U9349 (N_9349,N_5432,N_7834);
and U9350 (N_9350,N_5093,N_7541);
or U9351 (N_9351,N_6266,N_6119);
and U9352 (N_9352,N_5087,N_5681);
nand U9353 (N_9353,N_5963,N_7875);
nor U9354 (N_9354,N_6024,N_4094);
and U9355 (N_9355,N_7470,N_4280);
xnor U9356 (N_9356,N_7127,N_7889);
xor U9357 (N_9357,N_6234,N_7139);
and U9358 (N_9358,N_5356,N_6448);
and U9359 (N_9359,N_5672,N_6284);
or U9360 (N_9360,N_6496,N_4399);
and U9361 (N_9361,N_4963,N_7235);
and U9362 (N_9362,N_5219,N_6314);
nand U9363 (N_9363,N_7698,N_5434);
nand U9364 (N_9364,N_5565,N_6452);
nor U9365 (N_9365,N_4278,N_7740);
or U9366 (N_9366,N_4717,N_4513);
nor U9367 (N_9367,N_5737,N_4432);
nand U9368 (N_9368,N_4581,N_6088);
xnor U9369 (N_9369,N_6603,N_7314);
xor U9370 (N_9370,N_4924,N_6244);
and U9371 (N_9371,N_5420,N_5013);
nand U9372 (N_9372,N_7588,N_6575);
nand U9373 (N_9373,N_5521,N_7585);
and U9374 (N_9374,N_5510,N_4689);
nor U9375 (N_9375,N_7271,N_7709);
nand U9376 (N_9376,N_6332,N_5285);
xor U9377 (N_9377,N_7644,N_6121);
nor U9378 (N_9378,N_5495,N_6327);
xor U9379 (N_9379,N_7492,N_4325);
or U9380 (N_9380,N_5118,N_6531);
or U9381 (N_9381,N_4487,N_6987);
xor U9382 (N_9382,N_4225,N_5163);
nor U9383 (N_9383,N_5539,N_7155);
and U9384 (N_9384,N_5074,N_6125);
nor U9385 (N_9385,N_5140,N_6632);
or U9386 (N_9386,N_6015,N_4594);
and U9387 (N_9387,N_6672,N_5195);
xnor U9388 (N_9388,N_7936,N_6261);
nand U9389 (N_9389,N_4013,N_5197);
and U9390 (N_9390,N_7526,N_6099);
nor U9391 (N_9391,N_4084,N_7334);
or U9392 (N_9392,N_7094,N_4803);
or U9393 (N_9393,N_6194,N_4453);
or U9394 (N_9394,N_5165,N_5090);
nor U9395 (N_9395,N_6143,N_4206);
xor U9396 (N_9396,N_5155,N_6845);
nor U9397 (N_9397,N_4333,N_6705);
nand U9398 (N_9398,N_4350,N_6151);
nand U9399 (N_9399,N_7723,N_4037);
nand U9400 (N_9400,N_4787,N_5308);
nor U9401 (N_9401,N_6953,N_7769);
nor U9402 (N_9402,N_4727,N_5306);
and U9403 (N_9403,N_5396,N_4468);
nand U9404 (N_9404,N_4908,N_6464);
or U9405 (N_9405,N_4448,N_7326);
nand U9406 (N_9406,N_7471,N_4845);
and U9407 (N_9407,N_6166,N_6296);
xor U9408 (N_9408,N_6900,N_7577);
or U9409 (N_9409,N_5460,N_7117);
nor U9410 (N_9410,N_6903,N_5957);
or U9411 (N_9411,N_6640,N_6830);
nor U9412 (N_9412,N_7940,N_6576);
nand U9413 (N_9413,N_4828,N_7957);
or U9414 (N_9414,N_4636,N_4100);
xnor U9415 (N_9415,N_5050,N_5346);
nand U9416 (N_9416,N_5535,N_6643);
nor U9417 (N_9417,N_4349,N_4497);
or U9418 (N_9418,N_5875,N_6948);
nand U9419 (N_9419,N_6647,N_4041);
and U9420 (N_9420,N_6624,N_4486);
nand U9421 (N_9421,N_4347,N_7992);
xnor U9422 (N_9422,N_4233,N_6098);
nor U9423 (N_9423,N_5636,N_4289);
xnor U9424 (N_9424,N_5983,N_5538);
and U9425 (N_9425,N_7782,N_6130);
or U9426 (N_9426,N_6252,N_6178);
xnor U9427 (N_9427,N_5807,N_4886);
or U9428 (N_9428,N_4880,N_6706);
and U9429 (N_9429,N_4578,N_7464);
nor U9430 (N_9430,N_7172,N_7378);
nand U9431 (N_9431,N_4197,N_6037);
nor U9432 (N_9432,N_4275,N_5570);
and U9433 (N_9433,N_5313,N_4341);
nand U9434 (N_9434,N_6147,N_5860);
or U9435 (N_9435,N_7261,N_5858);
or U9436 (N_9436,N_6281,N_7250);
nand U9437 (N_9437,N_6786,N_4973);
nand U9438 (N_9438,N_5276,N_5966);
or U9439 (N_9439,N_7583,N_7804);
xnor U9440 (N_9440,N_6010,N_4871);
and U9441 (N_9441,N_4974,N_5121);
nand U9442 (N_9442,N_7130,N_6400);
nor U9443 (N_9443,N_6625,N_4286);
or U9444 (N_9444,N_5224,N_7258);
nor U9445 (N_9445,N_5367,N_5602);
xnor U9446 (N_9446,N_6519,N_4143);
nor U9447 (N_9447,N_5273,N_7787);
and U9448 (N_9448,N_7527,N_6134);
and U9449 (N_9449,N_4439,N_6128);
or U9450 (N_9450,N_5344,N_4263);
and U9451 (N_9451,N_5143,N_5029);
nand U9452 (N_9452,N_7075,N_5122);
or U9453 (N_9453,N_5358,N_4223);
nand U9454 (N_9454,N_6957,N_5928);
nand U9455 (N_9455,N_4932,N_7489);
nor U9456 (N_9456,N_7744,N_6553);
nor U9457 (N_9457,N_5251,N_5033);
nand U9458 (N_9458,N_6974,N_4202);
xor U9459 (N_9459,N_6366,N_4919);
nor U9460 (N_9460,N_7625,N_6354);
nor U9461 (N_9461,N_5907,N_5018);
or U9462 (N_9462,N_6751,N_4544);
nor U9463 (N_9463,N_5745,N_5265);
or U9464 (N_9464,N_7164,N_6302);
nor U9465 (N_9465,N_4539,N_5422);
nand U9466 (N_9466,N_7674,N_6590);
and U9467 (N_9467,N_7530,N_7733);
nand U9468 (N_9468,N_6139,N_6013);
and U9469 (N_9469,N_4368,N_6587);
and U9470 (N_9470,N_4927,N_5780);
xor U9471 (N_9471,N_6934,N_4836);
nand U9472 (N_9472,N_5236,N_6293);
or U9473 (N_9473,N_7057,N_4147);
nor U9474 (N_9474,N_4603,N_6876);
xor U9475 (N_9475,N_7843,N_4596);
or U9476 (N_9476,N_7173,N_6490);
xnor U9477 (N_9477,N_4875,N_4935);
or U9478 (N_9478,N_4454,N_4415);
and U9479 (N_9479,N_4632,N_6270);
or U9480 (N_9480,N_4373,N_4789);
nor U9481 (N_9481,N_5751,N_7946);
and U9482 (N_9482,N_6409,N_5692);
nor U9483 (N_9483,N_6416,N_6568);
and U9484 (N_9484,N_7981,N_5734);
nor U9485 (N_9485,N_4329,N_7919);
nor U9486 (N_9486,N_6762,N_6733);
and U9487 (N_9487,N_7281,N_7786);
and U9488 (N_9488,N_7339,N_5862);
nor U9489 (N_9489,N_5959,N_4808);
xor U9490 (N_9490,N_6782,N_4992);
and U9491 (N_9491,N_7990,N_7559);
or U9492 (N_9492,N_7350,N_6616);
or U9493 (N_9493,N_7415,N_5214);
or U9494 (N_9494,N_4872,N_6600);
nor U9495 (N_9495,N_5906,N_4788);
or U9496 (N_9496,N_4716,N_5156);
nor U9497 (N_9497,N_6511,N_5177);
and U9498 (N_9498,N_6517,N_4910);
or U9499 (N_9499,N_6885,N_4377);
xor U9500 (N_9500,N_6441,N_6627);
or U9501 (N_9501,N_5390,N_7027);
nor U9502 (N_9502,N_7232,N_7362);
and U9503 (N_9503,N_6227,N_6895);
nand U9504 (N_9504,N_5470,N_5789);
or U9505 (N_9505,N_4674,N_7499);
nand U9506 (N_9506,N_7665,N_6066);
xor U9507 (N_9507,N_4893,N_5187);
nand U9508 (N_9508,N_7272,N_7195);
or U9509 (N_9509,N_6756,N_4458);
nand U9510 (N_9510,N_5770,N_4294);
nand U9511 (N_9511,N_6272,N_4352);
or U9512 (N_9512,N_7450,N_5943);
nor U9513 (N_9513,N_4428,N_5603);
and U9514 (N_9514,N_6461,N_4628);
or U9515 (N_9515,N_6247,N_4134);
nor U9516 (N_9516,N_7676,N_5801);
and U9517 (N_9517,N_6924,N_5483);
or U9518 (N_9518,N_6620,N_6309);
or U9519 (N_9519,N_6819,N_7571);
and U9520 (N_9520,N_4216,N_4782);
nor U9521 (N_9521,N_7590,N_5147);
or U9522 (N_9522,N_7546,N_6527);
nand U9523 (N_9523,N_7854,N_6859);
and U9524 (N_9524,N_6621,N_7310);
nor U9525 (N_9525,N_7537,N_7840);
nor U9526 (N_9526,N_6567,N_5244);
nor U9527 (N_9527,N_5788,N_7277);
nor U9528 (N_9528,N_6630,N_4214);
nor U9529 (N_9529,N_6411,N_7347);
xnor U9530 (N_9530,N_6431,N_6798);
nor U9531 (N_9531,N_6674,N_5124);
nand U9532 (N_9532,N_4970,N_5703);
xnor U9533 (N_9533,N_6984,N_7720);
nand U9534 (N_9534,N_6459,N_6995);
and U9535 (N_9535,N_4449,N_4838);
and U9536 (N_9536,N_7531,N_5365);
or U9537 (N_9537,N_7828,N_4786);
or U9538 (N_9538,N_7793,N_5748);
or U9539 (N_9539,N_7465,N_6510);
xnor U9540 (N_9540,N_6610,N_4500);
and U9541 (N_9541,N_5282,N_6304);
and U9542 (N_9542,N_4597,N_4086);
or U9543 (N_9543,N_5517,N_6310);
nor U9544 (N_9544,N_6051,N_5471);
or U9545 (N_9545,N_4946,N_5351);
nand U9546 (N_9546,N_5546,N_7214);
nor U9547 (N_9547,N_6680,N_4067);
nand U9548 (N_9548,N_5096,N_6653);
xnor U9549 (N_9549,N_6202,N_5120);
or U9550 (N_9550,N_4138,N_7569);
xnor U9551 (N_9551,N_7361,N_7037);
or U9552 (N_9552,N_5380,N_7776);
and U9553 (N_9553,N_7289,N_7849);
nand U9554 (N_9554,N_6862,N_5834);
nor U9555 (N_9555,N_6472,N_5724);
xor U9556 (N_9556,N_6761,N_4336);
or U9557 (N_9557,N_4756,N_7418);
and U9558 (N_9558,N_7710,N_5972);
nor U9559 (N_9559,N_5416,N_7325);
or U9560 (N_9560,N_6019,N_7612);
nand U9561 (N_9561,N_7993,N_7063);
xnor U9562 (N_9562,N_6097,N_4548);
and U9563 (N_9563,N_6329,N_5028);
nand U9564 (N_9564,N_7651,N_7520);
and U9565 (N_9565,N_6853,N_5430);
or U9566 (N_9566,N_7073,N_7218);
nor U9567 (N_9567,N_6996,N_7859);
xnor U9568 (N_9568,N_7203,N_6439);
nor U9569 (N_9569,N_6615,N_7018);
and U9570 (N_9570,N_6420,N_5555);
or U9571 (N_9571,N_7838,N_5153);
nand U9572 (N_9572,N_6550,N_5609);
or U9573 (N_9573,N_5970,N_4707);
or U9574 (N_9574,N_5084,N_4360);
or U9575 (N_9575,N_6742,N_7568);
or U9576 (N_9576,N_5103,N_4475);
nor U9577 (N_9577,N_5412,N_6611);
nand U9578 (N_9578,N_4657,N_4463);
nand U9579 (N_9579,N_6814,N_7983);
nor U9580 (N_9580,N_6356,N_5067);
nor U9581 (N_9581,N_5142,N_5528);
and U9582 (N_9582,N_7105,N_7323);
xor U9583 (N_9583,N_6558,N_6880);
or U9584 (N_9584,N_4554,N_5519);
or U9585 (N_9585,N_5844,N_7771);
nor U9586 (N_9586,N_4774,N_4253);
xor U9587 (N_9587,N_4846,N_5610);
nor U9588 (N_9588,N_5484,N_6868);
nor U9589 (N_9589,N_7414,N_7119);
and U9590 (N_9590,N_5407,N_6052);
nor U9591 (N_9591,N_5189,N_6236);
nand U9592 (N_9592,N_7942,N_5804);
and U9593 (N_9593,N_6975,N_5900);
or U9594 (N_9594,N_5005,N_6047);
nand U9595 (N_9595,N_4938,N_7545);
and U9596 (N_9596,N_7091,N_5611);
nor U9597 (N_9597,N_7603,N_5608);
nor U9598 (N_9598,N_7153,N_7141);
or U9599 (N_9599,N_6071,N_4986);
nand U9600 (N_9600,N_6209,N_7745);
nand U9601 (N_9601,N_4741,N_6626);
xor U9602 (N_9602,N_5865,N_4862);
nor U9603 (N_9603,N_4996,N_4759);
nand U9604 (N_9604,N_7306,N_5824);
nor U9605 (N_9605,N_7684,N_5893);
nor U9606 (N_9606,N_4545,N_4255);
nor U9607 (N_9607,N_5110,N_6375);
nand U9608 (N_9608,N_6124,N_6703);
nor U9609 (N_9609,N_6339,N_7065);
or U9610 (N_9610,N_6791,N_7193);
or U9611 (N_9611,N_7332,N_7986);
and U9612 (N_9612,N_7264,N_5183);
or U9613 (N_9613,N_6312,N_4257);
nand U9614 (N_9614,N_7265,N_4180);
nor U9615 (N_9615,N_6504,N_6965);
nor U9616 (N_9616,N_5262,N_4429);
nor U9617 (N_9617,N_5713,N_4227);
and U9618 (N_9618,N_6947,N_7291);
and U9619 (N_9619,N_5886,N_7070);
or U9620 (N_9620,N_5350,N_6306);
or U9621 (N_9621,N_5525,N_7878);
nor U9622 (N_9622,N_5291,N_6233);
nor U9623 (N_9623,N_5095,N_4900);
and U9624 (N_9624,N_4720,N_4943);
or U9625 (N_9625,N_4965,N_5534);
nor U9626 (N_9626,N_5058,N_5366);
or U9627 (N_9627,N_6006,N_4070);
or U9628 (N_9628,N_6631,N_5423);
nor U9629 (N_9629,N_5856,N_5654);
and U9630 (N_9630,N_5462,N_7346);
nor U9631 (N_9631,N_5680,N_6840);
or U9632 (N_9632,N_4708,N_6337);
xor U9633 (N_9633,N_5868,N_7237);
nor U9634 (N_9634,N_4385,N_5478);
or U9635 (N_9635,N_4413,N_5968);
and U9636 (N_9636,N_5146,N_4507);
nand U9637 (N_9637,N_6103,N_6072);
and U9638 (N_9638,N_4568,N_5092);
xnor U9639 (N_9639,N_7819,N_6750);
nor U9640 (N_9640,N_6646,N_6165);
and U9641 (N_9641,N_4116,N_5689);
xnor U9642 (N_9642,N_4028,N_7090);
and U9643 (N_9643,N_6824,N_5239);
nor U9644 (N_9644,N_5243,N_4537);
and U9645 (N_9645,N_6909,N_7452);
nand U9646 (N_9646,N_6157,N_4314);
nor U9647 (N_9647,N_6679,N_6515);
nor U9648 (N_9648,N_5795,N_4903);
or U9649 (N_9649,N_4087,N_6259);
nand U9650 (N_9650,N_6397,N_6315);
nor U9651 (N_9651,N_5650,N_4899);
nor U9652 (N_9652,N_5512,N_7677);
nand U9653 (N_9653,N_6604,N_6715);
nand U9654 (N_9654,N_7557,N_6708);
and U9655 (N_9655,N_4244,N_4779);
xor U9656 (N_9656,N_7138,N_4393);
or U9657 (N_9657,N_6436,N_4126);
nor U9658 (N_9658,N_7121,N_7011);
or U9659 (N_9659,N_6883,N_5332);
or U9660 (N_9660,N_4878,N_5982);
xor U9661 (N_9661,N_7000,N_5232);
or U9662 (N_9662,N_7459,N_5908);
nor U9663 (N_9663,N_6110,N_6671);
nor U9664 (N_9664,N_6239,N_4794);
and U9665 (N_9665,N_4445,N_6455);
and U9666 (N_9666,N_5583,N_4340);
nor U9667 (N_9667,N_5368,N_7240);
nor U9668 (N_9668,N_7110,N_5270);
and U9669 (N_9669,N_6635,N_6711);
and U9670 (N_9670,N_6700,N_5655);
or U9671 (N_9671,N_4063,N_5312);
or U9672 (N_9672,N_7927,N_6131);
nor U9673 (N_9673,N_7156,N_6003);
nand U9674 (N_9674,N_5015,N_4993);
or U9675 (N_9675,N_4850,N_6294);
nand U9676 (N_9676,N_7128,N_5779);
or U9677 (N_9677,N_4667,N_6123);
nand U9678 (N_9678,N_7005,N_6946);
or U9679 (N_9679,N_4909,N_5401);
or U9680 (N_9680,N_4738,N_6257);
or U9681 (N_9681,N_5941,N_4235);
nand U9682 (N_9682,N_6358,N_6582);
and U9683 (N_9683,N_5604,N_6860);
and U9684 (N_9684,N_4631,N_5335);
and U9685 (N_9685,N_4920,N_4391);
or U9686 (N_9686,N_5934,N_5260);
nand U9687 (N_9687,N_7696,N_6939);
or U9688 (N_9688,N_5952,N_6014);
or U9689 (N_9689,N_6691,N_5152);
nand U9690 (N_9690,N_7663,N_4132);
nand U9691 (N_9691,N_5882,N_4014);
or U9692 (N_9692,N_6173,N_4226);
nor U9693 (N_9693,N_5720,N_6491);
or U9694 (N_9694,N_4641,N_5811);
nand U9695 (N_9695,N_5903,N_7831);
and U9696 (N_9696,N_6927,N_4560);
or U9697 (N_9697,N_5345,N_7098);
nor U9698 (N_9698,N_7668,N_6307);
xor U9699 (N_9699,N_5665,N_4422);
xnor U9700 (N_9700,N_7032,N_4258);
nor U9701 (N_9701,N_5353,N_6753);
or U9702 (N_9702,N_6438,N_5199);
and U9703 (N_9703,N_6342,N_6379);
or U9704 (N_9704,N_7046,N_7670);
xor U9705 (N_9705,N_6977,N_7406);
nor U9706 (N_9706,N_6963,N_5829);
or U9707 (N_9707,N_6094,N_7490);
or U9708 (N_9708,N_4780,N_4446);
and U9709 (N_9709,N_7479,N_6140);
and U9710 (N_9710,N_5362,N_5933);
nand U9711 (N_9711,N_5361,N_7966);
nand U9712 (N_9712,N_6241,N_7774);
and U9713 (N_9713,N_4150,N_5744);
xnor U9714 (N_9714,N_7190,N_5418);
nor U9715 (N_9715,N_7548,N_7417);
nand U9716 (N_9716,N_6650,N_6662);
nand U9717 (N_9717,N_5557,N_6012);
xnor U9718 (N_9718,N_5979,N_6721);
xnor U9719 (N_9719,N_7779,N_5775);
or U9720 (N_9720,N_6685,N_4193);
xnor U9721 (N_9721,N_6932,N_4266);
nor U9722 (N_9722,N_5425,N_5778);
and U9723 (N_9723,N_6085,N_5821);
nor U9724 (N_9724,N_6016,N_5631);
xnor U9725 (N_9725,N_6728,N_7337);
and U9726 (N_9726,N_5883,N_5042);
nand U9727 (N_9727,N_5967,N_5212);
and U9728 (N_9728,N_4793,N_5782);
or U9729 (N_9729,N_7263,N_4999);
or U9730 (N_9730,N_6664,N_7455);
xor U9731 (N_9731,N_4144,N_6316);
or U9732 (N_9732,N_4460,N_6945);
nand U9733 (N_9733,N_4840,N_7331);
nand U9734 (N_9734,N_7168,N_6200);
nor U9735 (N_9735,N_6964,N_4785);
or U9736 (N_9736,N_6838,N_4313);
nor U9737 (N_9737,N_6856,N_6882);
nor U9738 (N_9738,N_5436,N_7432);
or U9739 (N_9739,N_6445,N_6955);
nand U9740 (N_9740,N_5277,N_6729);
and U9741 (N_9741,N_7593,N_4039);
nand U9742 (N_9742,N_4524,N_5159);
nand U9743 (N_9743,N_7017,N_7615);
or U9744 (N_9744,N_7639,N_5333);
nand U9745 (N_9745,N_6229,N_4168);
or U9746 (N_9746,N_4001,N_6499);
and U9747 (N_9747,N_6783,N_5936);
nor U9748 (N_9748,N_4069,N_4125);
nand U9749 (N_9749,N_7636,N_4412);
nor U9750 (N_9750,N_4046,N_7785);
nor U9751 (N_9751,N_6430,N_4451);
xnor U9752 (N_9752,N_7969,N_7275);
nor U9753 (N_9753,N_6651,N_5309);
or U9754 (N_9754,N_6479,N_4931);
nand U9755 (N_9755,N_4414,N_6091);
or U9756 (N_9756,N_5621,N_5235);
or U9757 (N_9757,N_6796,N_4047);
and U9758 (N_9758,N_6773,N_4101);
and U9759 (N_9759,N_6396,N_7517);
nand U9760 (N_9760,N_7975,N_4431);
nand U9761 (N_9761,N_6056,N_7029);
or U9762 (N_9762,N_6011,N_4000);
and U9763 (N_9763,N_5696,N_4198);
xnor U9764 (N_9764,N_4304,N_5869);
nor U9765 (N_9765,N_7124,N_4157);
nor U9766 (N_9766,N_5732,N_5170);
xor U9767 (N_9767,N_6652,N_6518);
nor U9768 (N_9768,N_5257,N_7995);
or U9769 (N_9769,N_6184,N_4484);
nand U9770 (N_9770,N_5851,N_6724);
or U9771 (N_9771,N_5486,N_7209);
and U9772 (N_9772,N_6697,N_4135);
and U9773 (N_9773,N_6100,N_4250);
and U9774 (N_9774,N_4582,N_7144);
xnor U9775 (N_9775,N_5749,N_4953);
nor U9776 (N_9776,N_7654,N_4635);
and U9777 (N_9777,N_5916,N_4529);
nor U9778 (N_9778,N_6393,N_6176);
or U9779 (N_9779,N_6978,N_7746);
or U9780 (N_9780,N_4045,N_5100);
and U9781 (N_9781,N_5940,N_5590);
nand U9782 (N_9782,N_7968,N_4380);
or U9783 (N_9783,N_7598,N_6609);
or U9784 (N_9784,N_5481,N_6063);
or U9785 (N_9785,N_4670,N_5662);
xnor U9786 (N_9786,N_6021,N_5898);
nand U9787 (N_9787,N_6279,N_4057);
or U9788 (N_9788,N_7647,N_5627);
nand U9789 (N_9789,N_7535,N_4285);
or U9790 (N_9790,N_6258,N_4190);
nor U9791 (N_9791,N_4677,N_4922);
nand U9792 (N_9792,N_5274,N_4219);
or U9793 (N_9793,N_5148,N_6232);
nand U9794 (N_9794,N_4411,N_5185);
and U9795 (N_9795,N_5964,N_4966);
or U9796 (N_9796,N_7054,N_6080);
or U9797 (N_9797,N_5151,N_5511);
nand U9798 (N_9798,N_4378,N_5424);
or U9799 (N_9799,N_6670,N_4783);
and U9800 (N_9800,N_6614,N_5082);
xor U9801 (N_9801,N_6918,N_5674);
or U9802 (N_9802,N_7055,N_5379);
and U9803 (N_9803,N_7994,N_7421);
or U9804 (N_9804,N_6190,N_6619);
nor U9805 (N_9805,N_5974,N_6898);
nand U9806 (N_9806,N_7762,N_5639);
and U9807 (N_9807,N_6138,N_7367);
or U9808 (N_9808,N_4550,N_7396);
nor U9809 (N_9809,N_6291,N_5678);
nor U9810 (N_9810,N_5747,N_4364);
and U9811 (N_9811,N_7120,N_4433);
or U9812 (N_9812,N_6212,N_5999);
and U9813 (N_9813,N_5861,N_4700);
and U9814 (N_9814,N_6639,N_6894);
and U9815 (N_9815,N_7697,N_5931);
nand U9816 (N_9816,N_5052,N_5167);
nor U9817 (N_9817,N_5269,N_5707);
or U9818 (N_9818,N_7025,N_7602);
nor U9819 (N_9819,N_6846,N_7476);
or U9820 (N_9820,N_6399,N_4948);
nand U9821 (N_9821,N_5355,N_6844);
or U9822 (N_9822,N_4934,N_4477);
nand U9823 (N_9823,N_4279,N_7830);
nor U9824 (N_9824,N_5990,N_6036);
nor U9825 (N_9825,N_4942,N_4633);
and U9826 (N_9826,N_6746,N_4884);
nand U9827 (N_9827,N_6203,N_7907);
or U9828 (N_9828,N_4972,N_5132);
or U9829 (N_9829,N_5953,N_7877);
or U9830 (N_9830,N_4868,N_6850);
and U9831 (N_9831,N_7381,N_7841);
and U9832 (N_9832,N_5307,N_6521);
and U9833 (N_9833,N_6403,N_7958);
or U9834 (N_9834,N_6556,N_4819);
or U9835 (N_9835,N_6273,N_5725);
nor U9836 (N_9836,N_7916,N_5840);
nand U9837 (N_9837,N_4323,N_4248);
or U9838 (N_9838,N_5012,N_6250);
nand U9839 (N_9839,N_5633,N_6928);
or U9840 (N_9840,N_7304,N_4613);
and U9841 (N_9841,N_5064,N_7895);
or U9842 (N_9842,N_5969,N_7444);
xnor U9843 (N_9843,N_6029,N_6785);
nand U9844 (N_9844,N_7129,N_5123);
nand U9845 (N_9845,N_5823,N_4371);
and U9846 (N_9846,N_4363,N_7839);
and U9847 (N_9847,N_5494,N_7359);
and U9848 (N_9848,N_5671,N_7581);
or U9849 (N_9849,N_5783,N_4564);
nand U9850 (N_9850,N_6562,N_6149);
or U9851 (N_9851,N_5162,N_4883);
nor U9852 (N_9852,N_7504,N_6481);
nand U9853 (N_9853,N_5991,N_7386);
and U9854 (N_9854,N_6888,N_6348);
nand U9855 (N_9855,N_4982,N_4382);
and U9856 (N_9856,N_5785,N_7681);
nor U9857 (N_9857,N_5009,N_6115);
nor U9858 (N_9858,N_6040,N_7376);
nor U9859 (N_9859,N_6766,N_5299);
or U9860 (N_9860,N_7199,N_7726);
and U9861 (N_9861,N_7076,N_6704);
nand U9862 (N_9862,N_4521,N_6391);
or U9863 (N_9863,N_7360,N_5220);
or U9864 (N_9864,N_7869,N_6940);
or U9865 (N_9865,N_7348,N_5210);
nand U9866 (N_9866,N_6075,N_7298);
nand U9867 (N_9867,N_7157,N_4563);
and U9868 (N_9868,N_5912,N_7949);
xor U9869 (N_9869,N_7068,N_6574);
and U9870 (N_9870,N_7056,N_5283);
and U9871 (N_9871,N_5245,N_5625);
and U9872 (N_9872,N_4051,N_7412);
nand U9873 (N_9873,N_4252,N_7151);
or U9874 (N_9874,N_7716,N_6359);
nor U9875 (N_9875,N_5409,N_4397);
and U9876 (N_9876,N_5056,N_5025);
or U9877 (N_9877,N_5141,N_7267);
nand U9878 (N_9878,N_6285,N_6990);
nand U9879 (N_9879,N_7102,N_6793);
and U9880 (N_9880,N_6077,N_5803);
and U9881 (N_9881,N_7658,N_7095);
nor U9882 (N_9882,N_4882,N_7134);
or U9883 (N_9883,N_5419,N_6478);
or U9884 (N_9884,N_7719,N_5046);
nand U9885 (N_9885,N_7764,N_6580);
nand U9886 (N_9886,N_4775,N_7833);
xor U9887 (N_9887,N_4849,N_6912);
and U9888 (N_9888,N_5493,N_7364);
or U9889 (N_9889,N_4680,N_6534);
and U9890 (N_9890,N_6465,N_4533);
nand U9891 (N_9891,N_6772,N_7483);
nand U9892 (N_9892,N_6973,N_7458);
or U9893 (N_9893,N_5007,N_5544);
xnor U9894 (N_9894,N_7897,N_4473);
or U9895 (N_9895,N_5008,N_7512);
and U9896 (N_9896,N_6355,N_6398);
nor U9897 (N_9897,N_5134,N_4129);
nand U9898 (N_9898,N_7166,N_5504);
and U9899 (N_9899,N_6421,N_4998);
xor U9900 (N_9900,N_4220,N_7620);
or U9901 (N_9901,N_6714,N_4022);
or U9902 (N_9902,N_5160,N_7160);
nand U9903 (N_9903,N_4272,N_4199);
or U9904 (N_9904,N_6617,N_7473);
nand U9905 (N_9905,N_6663,N_5289);
nor U9906 (N_9906,N_7383,N_7821);
nand U9907 (N_9907,N_5540,N_7034);
or U9908 (N_9908,N_7224,N_6297);
nor U9909 (N_9909,N_4912,N_7814);
or U9910 (N_9910,N_7801,N_4516);
or U9911 (N_9911,N_6848,N_5324);
nor U9912 (N_9912,N_6158,N_5079);
and U9913 (N_9913,N_5600,N_4165);
nor U9914 (N_9914,N_7502,N_5323);
nor U9915 (N_9915,N_5016,N_5049);
nand U9916 (N_9916,N_5587,N_7906);
nor U9917 (N_9917,N_6768,N_4704);
or U9918 (N_9918,N_6999,N_7510);
and U9919 (N_9919,N_7296,N_7934);
or U9920 (N_9920,N_7269,N_6132);
nor U9921 (N_9921,N_6718,N_4241);
nor U9922 (N_9922,N_4969,N_4583);
nor U9923 (N_9923,N_6902,N_5686);
xnor U9924 (N_9924,N_7734,N_6009);
xnor U9925 (N_9925,N_5961,N_4183);
nand U9926 (N_9926,N_6350,N_4648);
nor U9927 (N_9927,N_5509,N_6242);
nor U9928 (N_9928,N_4163,N_6017);
nand U9929 (N_9929,N_4291,N_7996);
nand U9930 (N_9930,N_4276,N_5014);
nand U9931 (N_9931,N_4355,N_6654);
nor U9932 (N_9932,N_7796,N_7807);
nor U9933 (N_9933,N_4489,N_5429);
nand U9934 (N_9934,N_7122,N_5455);
and U9935 (N_9935,N_6152,N_4302);
or U9936 (N_9936,N_6207,N_7702);
or U9937 (N_9937,N_7974,N_4091);
nand U9938 (N_9938,N_7505,N_7695);
and U9939 (N_9939,N_7704,N_6434);
nand U9940 (N_9940,N_7892,N_4897);
xor U9941 (N_9941,N_5208,N_7441);
nor U9942 (N_9942,N_5492,N_6122);
or U9943 (N_9943,N_4962,N_4476);
nor U9944 (N_9944,N_5787,N_7204);
and U9945 (N_9945,N_7816,N_4652);
or U9946 (N_9946,N_7513,N_7753);
nor U9947 (N_9947,N_6002,N_5741);
or U9948 (N_9948,N_5595,N_7921);
nand U9949 (N_9949,N_4714,N_4174);
nor U9950 (N_9950,N_5473,N_4152);
nand U9951 (N_9951,N_4588,N_7896);
nand U9952 (N_9952,N_4863,N_7294);
nor U9953 (N_9953,N_6217,N_7353);
or U9954 (N_9954,N_4598,N_6794);
nor U9955 (N_9955,N_6301,N_6634);
and U9956 (N_9956,N_5919,N_4656);
nor U9957 (N_9957,N_7356,N_6267);
nand U9958 (N_9958,N_5542,N_6589);
or U9959 (N_9959,N_6874,N_4520);
and U9960 (N_9960,N_4517,N_7652);
nand U9961 (N_9961,N_5617,N_6470);
nand U9962 (N_9962,N_6917,N_4208);
and U9963 (N_9963,N_5976,N_5853);
nor U9964 (N_9964,N_7112,N_6944);
nor U9965 (N_9965,N_5218,N_5247);
nor U9966 (N_9966,N_7397,N_4751);
nand U9967 (N_9967,N_6317,N_6516);
nand U9968 (N_9968,N_7268,N_5369);
nand U9969 (N_9969,N_4262,N_6861);
nand U9970 (N_9970,N_7001,N_5798);
or U9971 (N_9971,N_6812,N_4625);
nand U9972 (N_9972,N_5086,N_4565);
nand U9973 (N_9973,N_5073,N_6757);
and U9974 (N_9974,N_5354,N_7463);
nand U9975 (N_9975,N_4123,N_4852);
nand U9976 (N_9976,N_4021,N_5169);
and U9977 (N_9977,N_5427,N_6913);
and U9978 (N_9978,N_5318,N_7910);
nor U9979 (N_9979,N_7851,N_6536);
or U9980 (N_9980,N_6788,N_6062);
and U9981 (N_9981,N_4256,N_5456);
nand U9982 (N_9982,N_5296,N_5532);
and U9983 (N_9983,N_5802,N_4757);
nor U9984 (N_9984,N_5226,N_4748);
or U9985 (N_9985,N_5201,N_5458);
nor U9986 (N_9986,N_5272,N_7754);
or U9987 (N_9987,N_5130,N_4660);
or U9988 (N_9988,N_7200,N_5753);
nand U9989 (N_9989,N_6805,N_5406);
nand U9990 (N_9990,N_6204,N_4205);
and U9991 (N_9991,N_6914,N_4732);
or U9992 (N_9992,N_7407,N_4559);
nor U9993 (N_9993,N_6586,N_5403);
and U9994 (N_9994,N_7635,N_5360);
nor U9995 (N_9995,N_7308,N_5305);
or U9996 (N_9996,N_7436,N_4348);
nand U9997 (N_9997,N_5711,N_6602);
or U9998 (N_9998,N_4089,N_7059);
and U9999 (N_9999,N_6905,N_6265);
nor U10000 (N_10000,N_6692,N_7258);
and U10001 (N_10001,N_6510,N_7389);
nand U10002 (N_10002,N_6720,N_7464);
nand U10003 (N_10003,N_7928,N_6377);
xor U10004 (N_10004,N_6994,N_4739);
nor U10005 (N_10005,N_6324,N_6815);
nand U10006 (N_10006,N_5993,N_6126);
and U10007 (N_10007,N_6854,N_4081);
nand U10008 (N_10008,N_7210,N_4314);
xor U10009 (N_10009,N_4869,N_4835);
or U10010 (N_10010,N_7681,N_4375);
and U10011 (N_10011,N_6890,N_7481);
and U10012 (N_10012,N_5358,N_6560);
nor U10013 (N_10013,N_6334,N_6480);
nand U10014 (N_10014,N_5503,N_5398);
and U10015 (N_10015,N_4013,N_4387);
xnor U10016 (N_10016,N_4141,N_7288);
nor U10017 (N_10017,N_4828,N_7793);
and U10018 (N_10018,N_5065,N_7621);
xnor U10019 (N_10019,N_7118,N_6536);
or U10020 (N_10020,N_6616,N_6007);
or U10021 (N_10021,N_5318,N_6560);
nand U10022 (N_10022,N_6967,N_6656);
nand U10023 (N_10023,N_6263,N_6434);
xor U10024 (N_10024,N_5041,N_6341);
nor U10025 (N_10025,N_6473,N_5166);
nor U10026 (N_10026,N_5728,N_6122);
nor U10027 (N_10027,N_7315,N_7392);
nor U10028 (N_10028,N_4821,N_4336);
nand U10029 (N_10029,N_4463,N_5538);
or U10030 (N_10030,N_7074,N_4167);
or U10031 (N_10031,N_4188,N_6199);
or U10032 (N_10032,N_6573,N_5014);
nand U10033 (N_10033,N_6890,N_4206);
nand U10034 (N_10034,N_6206,N_5074);
nor U10035 (N_10035,N_7155,N_6301);
or U10036 (N_10036,N_5907,N_6838);
nand U10037 (N_10037,N_6367,N_6491);
and U10038 (N_10038,N_6523,N_7433);
xor U10039 (N_10039,N_4129,N_5681);
nor U10040 (N_10040,N_5973,N_5634);
nor U10041 (N_10041,N_7428,N_6494);
and U10042 (N_10042,N_6298,N_6487);
or U10043 (N_10043,N_6801,N_7313);
nand U10044 (N_10044,N_5649,N_5622);
or U10045 (N_10045,N_5589,N_5199);
and U10046 (N_10046,N_6854,N_6172);
nor U10047 (N_10047,N_5813,N_6670);
or U10048 (N_10048,N_4424,N_5134);
xnor U10049 (N_10049,N_5272,N_7747);
nor U10050 (N_10050,N_5065,N_5638);
or U10051 (N_10051,N_5261,N_4857);
nor U10052 (N_10052,N_6526,N_4627);
and U10053 (N_10053,N_4272,N_7704);
and U10054 (N_10054,N_4724,N_4699);
and U10055 (N_10055,N_7724,N_6592);
and U10056 (N_10056,N_5317,N_6520);
and U10057 (N_10057,N_5077,N_6770);
nand U10058 (N_10058,N_7794,N_7368);
nand U10059 (N_10059,N_5965,N_4534);
or U10060 (N_10060,N_7516,N_4901);
or U10061 (N_10061,N_5645,N_6242);
nand U10062 (N_10062,N_5473,N_7573);
and U10063 (N_10063,N_4924,N_6989);
or U10064 (N_10064,N_4453,N_6800);
and U10065 (N_10065,N_6661,N_5844);
nor U10066 (N_10066,N_4032,N_4196);
and U10067 (N_10067,N_4833,N_6824);
and U10068 (N_10068,N_6370,N_4490);
nor U10069 (N_10069,N_5906,N_6114);
and U10070 (N_10070,N_6988,N_4707);
nand U10071 (N_10071,N_5717,N_5754);
nand U10072 (N_10072,N_6593,N_7004);
nor U10073 (N_10073,N_6024,N_6823);
or U10074 (N_10074,N_7893,N_4283);
xnor U10075 (N_10075,N_4587,N_7415);
or U10076 (N_10076,N_6949,N_6627);
and U10077 (N_10077,N_4466,N_4574);
nor U10078 (N_10078,N_6492,N_7745);
nor U10079 (N_10079,N_4807,N_4065);
or U10080 (N_10080,N_4682,N_5244);
nand U10081 (N_10081,N_6653,N_7631);
nor U10082 (N_10082,N_6693,N_6143);
nand U10083 (N_10083,N_4832,N_7212);
and U10084 (N_10084,N_4038,N_4342);
xor U10085 (N_10085,N_6694,N_4377);
nand U10086 (N_10086,N_5007,N_6877);
xnor U10087 (N_10087,N_5885,N_4794);
or U10088 (N_10088,N_6989,N_7446);
or U10089 (N_10089,N_5674,N_5741);
nor U10090 (N_10090,N_7016,N_7752);
or U10091 (N_10091,N_6773,N_4307);
nor U10092 (N_10092,N_5652,N_5012);
or U10093 (N_10093,N_5302,N_4345);
nand U10094 (N_10094,N_4699,N_4975);
nand U10095 (N_10095,N_6496,N_6714);
and U10096 (N_10096,N_4349,N_7511);
and U10097 (N_10097,N_4064,N_5563);
xor U10098 (N_10098,N_6719,N_6229);
and U10099 (N_10099,N_6512,N_4852);
nand U10100 (N_10100,N_7009,N_6226);
and U10101 (N_10101,N_7083,N_5935);
or U10102 (N_10102,N_5356,N_7529);
or U10103 (N_10103,N_6484,N_6041);
and U10104 (N_10104,N_6998,N_6316);
nand U10105 (N_10105,N_7934,N_5072);
nor U10106 (N_10106,N_6123,N_4500);
nand U10107 (N_10107,N_6511,N_6533);
nor U10108 (N_10108,N_5093,N_6247);
xnor U10109 (N_10109,N_5551,N_5902);
or U10110 (N_10110,N_7708,N_6671);
and U10111 (N_10111,N_4117,N_5056);
nor U10112 (N_10112,N_5808,N_6353);
xor U10113 (N_10113,N_5676,N_6500);
nor U10114 (N_10114,N_6172,N_7744);
nor U10115 (N_10115,N_4017,N_5429);
nor U10116 (N_10116,N_6426,N_7976);
xnor U10117 (N_10117,N_6441,N_4062);
or U10118 (N_10118,N_7342,N_6443);
or U10119 (N_10119,N_6243,N_7240);
and U10120 (N_10120,N_7063,N_7620);
or U10121 (N_10121,N_5665,N_6685);
or U10122 (N_10122,N_4153,N_4253);
nand U10123 (N_10123,N_5297,N_7938);
or U10124 (N_10124,N_5413,N_5775);
nor U10125 (N_10125,N_6416,N_7347);
nand U10126 (N_10126,N_4995,N_6745);
nand U10127 (N_10127,N_6685,N_6385);
or U10128 (N_10128,N_7275,N_6990);
nor U10129 (N_10129,N_5371,N_6868);
nand U10130 (N_10130,N_4281,N_7589);
and U10131 (N_10131,N_6340,N_7632);
nand U10132 (N_10132,N_7917,N_5989);
xor U10133 (N_10133,N_4503,N_4080);
and U10134 (N_10134,N_6558,N_4521);
and U10135 (N_10135,N_7795,N_6069);
nand U10136 (N_10136,N_6183,N_5153);
or U10137 (N_10137,N_4988,N_5729);
and U10138 (N_10138,N_7897,N_5741);
and U10139 (N_10139,N_7805,N_7150);
and U10140 (N_10140,N_4677,N_4998);
or U10141 (N_10141,N_7641,N_7236);
or U10142 (N_10142,N_6878,N_5945);
nor U10143 (N_10143,N_4678,N_4161);
nand U10144 (N_10144,N_7635,N_5897);
nand U10145 (N_10145,N_4813,N_4703);
or U10146 (N_10146,N_7514,N_5211);
nor U10147 (N_10147,N_4270,N_5385);
and U10148 (N_10148,N_7295,N_6203);
or U10149 (N_10149,N_7568,N_5851);
nor U10150 (N_10150,N_5650,N_5239);
nand U10151 (N_10151,N_7350,N_7324);
nand U10152 (N_10152,N_4819,N_5457);
or U10153 (N_10153,N_7558,N_4711);
or U10154 (N_10154,N_5796,N_6132);
and U10155 (N_10155,N_5265,N_6328);
or U10156 (N_10156,N_4395,N_6674);
and U10157 (N_10157,N_7864,N_5747);
xor U10158 (N_10158,N_5639,N_7511);
xor U10159 (N_10159,N_7835,N_6991);
nand U10160 (N_10160,N_4402,N_7644);
nor U10161 (N_10161,N_5970,N_5039);
and U10162 (N_10162,N_4467,N_6380);
or U10163 (N_10163,N_7025,N_7738);
nor U10164 (N_10164,N_6112,N_6494);
or U10165 (N_10165,N_6660,N_6369);
or U10166 (N_10166,N_4268,N_4325);
nand U10167 (N_10167,N_6868,N_4756);
nand U10168 (N_10168,N_5125,N_6993);
nand U10169 (N_10169,N_4339,N_5556);
nor U10170 (N_10170,N_7250,N_6847);
nand U10171 (N_10171,N_6880,N_6553);
nand U10172 (N_10172,N_6307,N_5298);
xor U10173 (N_10173,N_7975,N_5298);
and U10174 (N_10174,N_4182,N_7496);
xnor U10175 (N_10175,N_5932,N_4947);
and U10176 (N_10176,N_5833,N_6898);
or U10177 (N_10177,N_5332,N_6628);
xnor U10178 (N_10178,N_7451,N_6837);
and U10179 (N_10179,N_7829,N_4013);
nand U10180 (N_10180,N_4888,N_4007);
or U10181 (N_10181,N_6335,N_4491);
and U10182 (N_10182,N_6170,N_7521);
nand U10183 (N_10183,N_6807,N_7985);
nand U10184 (N_10184,N_7507,N_4190);
nor U10185 (N_10185,N_6641,N_7386);
nor U10186 (N_10186,N_6193,N_6229);
and U10187 (N_10187,N_7994,N_6509);
and U10188 (N_10188,N_4484,N_4815);
and U10189 (N_10189,N_7385,N_7262);
and U10190 (N_10190,N_7993,N_6974);
xor U10191 (N_10191,N_5036,N_5904);
nor U10192 (N_10192,N_6449,N_7158);
nand U10193 (N_10193,N_5441,N_6622);
xor U10194 (N_10194,N_6110,N_7060);
and U10195 (N_10195,N_6113,N_7697);
and U10196 (N_10196,N_5197,N_4828);
nor U10197 (N_10197,N_6240,N_5791);
nor U10198 (N_10198,N_4332,N_6423);
xnor U10199 (N_10199,N_4200,N_4590);
or U10200 (N_10200,N_4081,N_6018);
and U10201 (N_10201,N_6158,N_4398);
nor U10202 (N_10202,N_4483,N_7324);
nor U10203 (N_10203,N_7837,N_7349);
and U10204 (N_10204,N_7556,N_4349);
nand U10205 (N_10205,N_6477,N_4828);
nor U10206 (N_10206,N_7759,N_4179);
nor U10207 (N_10207,N_6778,N_6244);
nand U10208 (N_10208,N_4010,N_6761);
and U10209 (N_10209,N_4735,N_6387);
or U10210 (N_10210,N_7317,N_7603);
or U10211 (N_10211,N_4055,N_6081);
nor U10212 (N_10212,N_4023,N_6948);
and U10213 (N_10213,N_7826,N_4907);
or U10214 (N_10214,N_6866,N_5495);
and U10215 (N_10215,N_5998,N_5928);
nand U10216 (N_10216,N_7775,N_5199);
and U10217 (N_10217,N_7429,N_5385);
or U10218 (N_10218,N_5036,N_6960);
xor U10219 (N_10219,N_4978,N_4619);
or U10220 (N_10220,N_5634,N_6916);
nand U10221 (N_10221,N_7772,N_5245);
nand U10222 (N_10222,N_5791,N_6250);
xnor U10223 (N_10223,N_7982,N_4316);
or U10224 (N_10224,N_5507,N_4145);
nor U10225 (N_10225,N_6932,N_7403);
xnor U10226 (N_10226,N_7280,N_6742);
nand U10227 (N_10227,N_5768,N_7276);
nor U10228 (N_10228,N_5455,N_7996);
and U10229 (N_10229,N_5779,N_5089);
or U10230 (N_10230,N_4752,N_7145);
nor U10231 (N_10231,N_6903,N_4905);
and U10232 (N_10232,N_6190,N_5192);
nand U10233 (N_10233,N_5038,N_6730);
nand U10234 (N_10234,N_7159,N_5691);
nor U10235 (N_10235,N_4564,N_5263);
or U10236 (N_10236,N_5083,N_6516);
nand U10237 (N_10237,N_7246,N_6848);
nor U10238 (N_10238,N_6213,N_6416);
nor U10239 (N_10239,N_4537,N_4705);
and U10240 (N_10240,N_4889,N_6803);
or U10241 (N_10241,N_6721,N_7150);
and U10242 (N_10242,N_5607,N_6970);
and U10243 (N_10243,N_7547,N_6943);
or U10244 (N_10244,N_5383,N_5452);
nand U10245 (N_10245,N_4442,N_7550);
nor U10246 (N_10246,N_7223,N_4769);
xnor U10247 (N_10247,N_6377,N_6895);
or U10248 (N_10248,N_6841,N_5252);
and U10249 (N_10249,N_5714,N_7210);
nand U10250 (N_10250,N_7813,N_4610);
nand U10251 (N_10251,N_5475,N_5680);
xor U10252 (N_10252,N_6896,N_5223);
and U10253 (N_10253,N_6365,N_5437);
and U10254 (N_10254,N_6664,N_6138);
nand U10255 (N_10255,N_7663,N_6845);
and U10256 (N_10256,N_7086,N_6214);
or U10257 (N_10257,N_7803,N_4988);
or U10258 (N_10258,N_5749,N_6680);
nor U10259 (N_10259,N_6438,N_4782);
or U10260 (N_10260,N_6377,N_7958);
nand U10261 (N_10261,N_4860,N_6120);
or U10262 (N_10262,N_5299,N_7846);
xnor U10263 (N_10263,N_4590,N_4970);
nand U10264 (N_10264,N_6383,N_5408);
nand U10265 (N_10265,N_4782,N_5154);
xor U10266 (N_10266,N_7599,N_4733);
nand U10267 (N_10267,N_5110,N_5066);
nand U10268 (N_10268,N_5063,N_7102);
nand U10269 (N_10269,N_5724,N_7181);
or U10270 (N_10270,N_7926,N_4655);
or U10271 (N_10271,N_6948,N_6988);
and U10272 (N_10272,N_4267,N_7134);
and U10273 (N_10273,N_7846,N_7866);
nand U10274 (N_10274,N_6938,N_5423);
nand U10275 (N_10275,N_7048,N_5390);
or U10276 (N_10276,N_5319,N_4851);
nand U10277 (N_10277,N_7065,N_4397);
or U10278 (N_10278,N_4948,N_4383);
or U10279 (N_10279,N_6632,N_4880);
nand U10280 (N_10280,N_5476,N_4949);
and U10281 (N_10281,N_6079,N_7483);
nand U10282 (N_10282,N_7510,N_6817);
and U10283 (N_10283,N_6511,N_5378);
nand U10284 (N_10284,N_4391,N_7423);
nor U10285 (N_10285,N_6756,N_4127);
and U10286 (N_10286,N_7909,N_4252);
nand U10287 (N_10287,N_7891,N_5385);
or U10288 (N_10288,N_7943,N_7978);
and U10289 (N_10289,N_4398,N_7549);
nor U10290 (N_10290,N_4449,N_6338);
nor U10291 (N_10291,N_5442,N_7645);
or U10292 (N_10292,N_6440,N_4543);
nor U10293 (N_10293,N_5489,N_7257);
or U10294 (N_10294,N_7528,N_7514);
nor U10295 (N_10295,N_4921,N_5705);
or U10296 (N_10296,N_4641,N_4930);
nor U10297 (N_10297,N_5879,N_7825);
and U10298 (N_10298,N_6922,N_7006);
nor U10299 (N_10299,N_5360,N_6802);
nor U10300 (N_10300,N_6825,N_5434);
and U10301 (N_10301,N_4532,N_6229);
nor U10302 (N_10302,N_7777,N_4447);
nand U10303 (N_10303,N_6645,N_4207);
and U10304 (N_10304,N_7097,N_7758);
or U10305 (N_10305,N_4204,N_7797);
nor U10306 (N_10306,N_4152,N_7410);
or U10307 (N_10307,N_4348,N_5721);
and U10308 (N_10308,N_4672,N_5520);
nand U10309 (N_10309,N_6768,N_6654);
nor U10310 (N_10310,N_6145,N_4597);
xnor U10311 (N_10311,N_4963,N_4133);
and U10312 (N_10312,N_6927,N_5198);
and U10313 (N_10313,N_4630,N_6741);
or U10314 (N_10314,N_5995,N_5346);
or U10315 (N_10315,N_6808,N_6514);
or U10316 (N_10316,N_7337,N_7190);
nor U10317 (N_10317,N_7775,N_5836);
nand U10318 (N_10318,N_6881,N_5703);
xor U10319 (N_10319,N_5160,N_4584);
and U10320 (N_10320,N_4929,N_7012);
nand U10321 (N_10321,N_6117,N_7961);
nor U10322 (N_10322,N_5653,N_5174);
nand U10323 (N_10323,N_6325,N_7480);
nand U10324 (N_10324,N_6243,N_4393);
xor U10325 (N_10325,N_4302,N_5601);
or U10326 (N_10326,N_5727,N_6448);
nand U10327 (N_10327,N_6725,N_6734);
or U10328 (N_10328,N_6436,N_7265);
nand U10329 (N_10329,N_6534,N_5382);
and U10330 (N_10330,N_5222,N_4918);
or U10331 (N_10331,N_7844,N_4602);
nor U10332 (N_10332,N_4861,N_6754);
xor U10333 (N_10333,N_6930,N_6088);
nor U10334 (N_10334,N_4797,N_7469);
and U10335 (N_10335,N_5457,N_7216);
or U10336 (N_10336,N_7150,N_6474);
xor U10337 (N_10337,N_4747,N_6802);
and U10338 (N_10338,N_5220,N_6360);
nand U10339 (N_10339,N_5181,N_5802);
and U10340 (N_10340,N_4641,N_5312);
or U10341 (N_10341,N_4413,N_4827);
nor U10342 (N_10342,N_7786,N_4697);
and U10343 (N_10343,N_4525,N_7228);
and U10344 (N_10344,N_6250,N_4844);
and U10345 (N_10345,N_4638,N_6868);
and U10346 (N_10346,N_7183,N_5288);
or U10347 (N_10347,N_4640,N_5351);
or U10348 (N_10348,N_7570,N_4948);
or U10349 (N_10349,N_6560,N_6194);
xnor U10350 (N_10350,N_4330,N_6844);
nor U10351 (N_10351,N_5924,N_4260);
xnor U10352 (N_10352,N_5843,N_6514);
or U10353 (N_10353,N_7835,N_6183);
or U10354 (N_10354,N_5378,N_6700);
nand U10355 (N_10355,N_7961,N_7469);
and U10356 (N_10356,N_7895,N_7914);
xor U10357 (N_10357,N_6068,N_5869);
and U10358 (N_10358,N_7444,N_6504);
or U10359 (N_10359,N_5111,N_4793);
and U10360 (N_10360,N_6136,N_6812);
and U10361 (N_10361,N_7733,N_6400);
and U10362 (N_10362,N_4006,N_4920);
nor U10363 (N_10363,N_5593,N_5486);
and U10364 (N_10364,N_7506,N_5200);
or U10365 (N_10365,N_5924,N_7082);
and U10366 (N_10366,N_6056,N_4060);
and U10367 (N_10367,N_7999,N_4890);
xor U10368 (N_10368,N_5607,N_7260);
nor U10369 (N_10369,N_7332,N_6565);
nand U10370 (N_10370,N_7189,N_5746);
nor U10371 (N_10371,N_5464,N_5988);
and U10372 (N_10372,N_4153,N_6722);
or U10373 (N_10373,N_7230,N_6798);
nand U10374 (N_10374,N_6305,N_5642);
and U10375 (N_10375,N_6633,N_6886);
and U10376 (N_10376,N_7215,N_4411);
nand U10377 (N_10377,N_4665,N_4011);
or U10378 (N_10378,N_4880,N_7614);
nand U10379 (N_10379,N_7110,N_7539);
or U10380 (N_10380,N_6850,N_7347);
nor U10381 (N_10381,N_4455,N_7123);
and U10382 (N_10382,N_5664,N_5922);
or U10383 (N_10383,N_5016,N_5584);
or U10384 (N_10384,N_4229,N_7708);
nand U10385 (N_10385,N_5458,N_4159);
and U10386 (N_10386,N_7777,N_5717);
or U10387 (N_10387,N_6513,N_6747);
or U10388 (N_10388,N_4488,N_4716);
or U10389 (N_10389,N_4608,N_5440);
and U10390 (N_10390,N_5737,N_7675);
nor U10391 (N_10391,N_7004,N_6951);
and U10392 (N_10392,N_5513,N_6805);
or U10393 (N_10393,N_6577,N_5176);
xnor U10394 (N_10394,N_4323,N_4107);
nand U10395 (N_10395,N_5258,N_6644);
nand U10396 (N_10396,N_7591,N_7582);
nor U10397 (N_10397,N_5074,N_4005);
and U10398 (N_10398,N_6077,N_4053);
nor U10399 (N_10399,N_5358,N_7006);
nor U10400 (N_10400,N_6915,N_6634);
or U10401 (N_10401,N_7472,N_6209);
or U10402 (N_10402,N_7364,N_4096);
nor U10403 (N_10403,N_4615,N_4191);
and U10404 (N_10404,N_6442,N_4338);
nor U10405 (N_10405,N_6884,N_7063);
and U10406 (N_10406,N_6145,N_6331);
and U10407 (N_10407,N_5969,N_5274);
xnor U10408 (N_10408,N_5841,N_7893);
nor U10409 (N_10409,N_7143,N_6473);
and U10410 (N_10410,N_7445,N_6127);
nand U10411 (N_10411,N_6463,N_4794);
and U10412 (N_10412,N_5614,N_4284);
nor U10413 (N_10413,N_6502,N_6815);
and U10414 (N_10414,N_6194,N_7389);
or U10415 (N_10415,N_5106,N_4441);
nor U10416 (N_10416,N_7908,N_7907);
nand U10417 (N_10417,N_6986,N_4197);
or U10418 (N_10418,N_4820,N_6624);
nor U10419 (N_10419,N_4468,N_4077);
nor U10420 (N_10420,N_6369,N_7324);
or U10421 (N_10421,N_6576,N_4403);
nand U10422 (N_10422,N_7663,N_4789);
nor U10423 (N_10423,N_6767,N_5075);
or U10424 (N_10424,N_4450,N_7358);
and U10425 (N_10425,N_5726,N_4472);
and U10426 (N_10426,N_4296,N_6783);
and U10427 (N_10427,N_4502,N_7915);
or U10428 (N_10428,N_6717,N_7425);
or U10429 (N_10429,N_4934,N_7813);
nor U10430 (N_10430,N_4048,N_5202);
nor U10431 (N_10431,N_6714,N_6808);
xnor U10432 (N_10432,N_6049,N_5061);
nor U10433 (N_10433,N_4969,N_7919);
nand U10434 (N_10434,N_5977,N_7357);
or U10435 (N_10435,N_5836,N_6785);
or U10436 (N_10436,N_7351,N_7639);
and U10437 (N_10437,N_6493,N_4812);
and U10438 (N_10438,N_5522,N_5428);
nand U10439 (N_10439,N_7880,N_4777);
and U10440 (N_10440,N_7816,N_6990);
nor U10441 (N_10441,N_7048,N_6682);
or U10442 (N_10442,N_7467,N_7722);
xnor U10443 (N_10443,N_7723,N_5357);
or U10444 (N_10444,N_5723,N_4007);
and U10445 (N_10445,N_6654,N_7556);
nor U10446 (N_10446,N_7221,N_6634);
and U10447 (N_10447,N_5113,N_5364);
and U10448 (N_10448,N_7848,N_5408);
and U10449 (N_10449,N_5401,N_4516);
and U10450 (N_10450,N_4583,N_4757);
nand U10451 (N_10451,N_6979,N_6336);
and U10452 (N_10452,N_5844,N_7793);
nand U10453 (N_10453,N_4520,N_5343);
nand U10454 (N_10454,N_5428,N_6650);
and U10455 (N_10455,N_5097,N_4765);
nor U10456 (N_10456,N_7150,N_4972);
nand U10457 (N_10457,N_5586,N_6430);
nand U10458 (N_10458,N_7802,N_5076);
and U10459 (N_10459,N_4496,N_5304);
or U10460 (N_10460,N_6087,N_5771);
xor U10461 (N_10461,N_7708,N_6540);
and U10462 (N_10462,N_4815,N_4609);
xor U10463 (N_10463,N_4212,N_6364);
and U10464 (N_10464,N_5397,N_7593);
nor U10465 (N_10465,N_7740,N_5286);
nand U10466 (N_10466,N_7443,N_5963);
or U10467 (N_10467,N_5222,N_7014);
or U10468 (N_10468,N_4242,N_6482);
nand U10469 (N_10469,N_6787,N_4294);
and U10470 (N_10470,N_7753,N_4959);
nor U10471 (N_10471,N_6081,N_7170);
nand U10472 (N_10472,N_5351,N_5983);
nand U10473 (N_10473,N_5468,N_4566);
nor U10474 (N_10474,N_4282,N_5923);
nor U10475 (N_10475,N_7750,N_4692);
or U10476 (N_10476,N_4166,N_4678);
or U10477 (N_10477,N_5896,N_7497);
and U10478 (N_10478,N_6185,N_6343);
nor U10479 (N_10479,N_7753,N_6617);
and U10480 (N_10480,N_7023,N_4201);
nor U10481 (N_10481,N_5091,N_7372);
and U10482 (N_10482,N_6036,N_4275);
xor U10483 (N_10483,N_6953,N_6803);
nand U10484 (N_10484,N_5219,N_5777);
nand U10485 (N_10485,N_6583,N_6413);
xnor U10486 (N_10486,N_4558,N_7748);
nand U10487 (N_10487,N_5235,N_5254);
xnor U10488 (N_10488,N_5836,N_6617);
nor U10489 (N_10489,N_5824,N_7391);
nor U10490 (N_10490,N_4352,N_6476);
and U10491 (N_10491,N_5164,N_7120);
nand U10492 (N_10492,N_5277,N_4582);
nor U10493 (N_10493,N_7878,N_7305);
nand U10494 (N_10494,N_7066,N_6167);
and U10495 (N_10495,N_4248,N_5817);
nor U10496 (N_10496,N_4059,N_6235);
and U10497 (N_10497,N_6775,N_4004);
nand U10498 (N_10498,N_7621,N_4841);
nand U10499 (N_10499,N_4349,N_5210);
nor U10500 (N_10500,N_4723,N_4772);
and U10501 (N_10501,N_5918,N_6022);
and U10502 (N_10502,N_5285,N_4246);
nand U10503 (N_10503,N_6036,N_5867);
or U10504 (N_10504,N_5130,N_5411);
nand U10505 (N_10505,N_4929,N_6322);
and U10506 (N_10506,N_4519,N_5874);
nand U10507 (N_10507,N_5553,N_7516);
nand U10508 (N_10508,N_7680,N_5807);
nor U10509 (N_10509,N_4707,N_7064);
nand U10510 (N_10510,N_5638,N_6700);
xnor U10511 (N_10511,N_6245,N_7879);
and U10512 (N_10512,N_5708,N_7979);
or U10513 (N_10513,N_5418,N_7524);
or U10514 (N_10514,N_4818,N_6110);
nand U10515 (N_10515,N_7825,N_4978);
or U10516 (N_10516,N_5592,N_6764);
or U10517 (N_10517,N_6598,N_5263);
and U10518 (N_10518,N_5650,N_6595);
nand U10519 (N_10519,N_5969,N_5093);
or U10520 (N_10520,N_5359,N_4879);
and U10521 (N_10521,N_5615,N_7447);
nand U10522 (N_10522,N_7163,N_4502);
xor U10523 (N_10523,N_4534,N_5467);
and U10524 (N_10524,N_4485,N_7485);
and U10525 (N_10525,N_7504,N_5365);
or U10526 (N_10526,N_5418,N_4738);
or U10527 (N_10527,N_7108,N_4507);
nor U10528 (N_10528,N_6873,N_5995);
and U10529 (N_10529,N_4498,N_5865);
or U10530 (N_10530,N_6784,N_5499);
xor U10531 (N_10531,N_7068,N_7800);
and U10532 (N_10532,N_7153,N_6084);
and U10533 (N_10533,N_4160,N_6121);
or U10534 (N_10534,N_4891,N_5150);
and U10535 (N_10535,N_4189,N_5761);
and U10536 (N_10536,N_6962,N_7294);
and U10537 (N_10537,N_5294,N_4928);
nand U10538 (N_10538,N_5030,N_7865);
or U10539 (N_10539,N_5842,N_7817);
xnor U10540 (N_10540,N_7467,N_4143);
or U10541 (N_10541,N_5520,N_4641);
nand U10542 (N_10542,N_6311,N_5042);
and U10543 (N_10543,N_5204,N_4746);
or U10544 (N_10544,N_6997,N_5223);
xor U10545 (N_10545,N_7785,N_4279);
and U10546 (N_10546,N_7974,N_7138);
or U10547 (N_10547,N_5373,N_5619);
and U10548 (N_10548,N_7846,N_6157);
and U10549 (N_10549,N_4032,N_6212);
and U10550 (N_10550,N_6736,N_7652);
and U10551 (N_10551,N_7051,N_5851);
nand U10552 (N_10552,N_7944,N_5846);
nand U10553 (N_10553,N_6627,N_7299);
and U10554 (N_10554,N_6312,N_6554);
or U10555 (N_10555,N_7017,N_4669);
nor U10556 (N_10556,N_6232,N_4446);
and U10557 (N_10557,N_6145,N_4489);
nand U10558 (N_10558,N_7687,N_5864);
or U10559 (N_10559,N_6580,N_7789);
xnor U10560 (N_10560,N_4871,N_5102);
nand U10561 (N_10561,N_7409,N_6937);
nor U10562 (N_10562,N_7930,N_4316);
nor U10563 (N_10563,N_6772,N_7956);
or U10564 (N_10564,N_7788,N_5354);
nand U10565 (N_10565,N_6758,N_5624);
and U10566 (N_10566,N_4386,N_7743);
or U10567 (N_10567,N_7721,N_5687);
nor U10568 (N_10568,N_6961,N_6690);
and U10569 (N_10569,N_7047,N_4009);
nor U10570 (N_10570,N_4629,N_4062);
and U10571 (N_10571,N_6513,N_7533);
nor U10572 (N_10572,N_7416,N_7995);
nand U10573 (N_10573,N_7557,N_7603);
nand U10574 (N_10574,N_6470,N_5888);
nor U10575 (N_10575,N_5599,N_4911);
nand U10576 (N_10576,N_6268,N_4258);
or U10577 (N_10577,N_6926,N_5999);
nand U10578 (N_10578,N_4575,N_5603);
nor U10579 (N_10579,N_6343,N_6646);
nor U10580 (N_10580,N_6759,N_7677);
and U10581 (N_10581,N_4200,N_4909);
or U10582 (N_10582,N_5874,N_7248);
or U10583 (N_10583,N_7344,N_7134);
nand U10584 (N_10584,N_5726,N_5808);
xor U10585 (N_10585,N_4118,N_7386);
and U10586 (N_10586,N_4678,N_7551);
nand U10587 (N_10587,N_5315,N_6963);
or U10588 (N_10588,N_5093,N_7260);
nor U10589 (N_10589,N_6378,N_6676);
nand U10590 (N_10590,N_6470,N_6879);
nand U10591 (N_10591,N_6717,N_4028);
or U10592 (N_10592,N_6157,N_6677);
and U10593 (N_10593,N_4587,N_5842);
nand U10594 (N_10594,N_5352,N_4015);
xor U10595 (N_10595,N_4651,N_4452);
nand U10596 (N_10596,N_6872,N_7509);
nor U10597 (N_10597,N_6773,N_6726);
or U10598 (N_10598,N_7843,N_5342);
and U10599 (N_10599,N_6909,N_7004);
nor U10600 (N_10600,N_4782,N_4030);
or U10601 (N_10601,N_5487,N_4012);
and U10602 (N_10602,N_6655,N_7046);
nor U10603 (N_10603,N_5612,N_6847);
nand U10604 (N_10604,N_6623,N_4761);
nand U10605 (N_10605,N_6069,N_5381);
xnor U10606 (N_10606,N_7683,N_5991);
or U10607 (N_10607,N_5983,N_7895);
nand U10608 (N_10608,N_5449,N_6404);
nand U10609 (N_10609,N_7395,N_7508);
or U10610 (N_10610,N_6771,N_6976);
nand U10611 (N_10611,N_4473,N_4359);
and U10612 (N_10612,N_6240,N_5954);
nand U10613 (N_10613,N_6280,N_4099);
nor U10614 (N_10614,N_7645,N_6842);
and U10615 (N_10615,N_6683,N_7446);
and U10616 (N_10616,N_4761,N_7591);
nor U10617 (N_10617,N_7444,N_7022);
xor U10618 (N_10618,N_7504,N_6770);
xnor U10619 (N_10619,N_7681,N_5733);
nor U10620 (N_10620,N_7063,N_6278);
nor U10621 (N_10621,N_4010,N_5922);
nor U10622 (N_10622,N_7113,N_7756);
or U10623 (N_10623,N_4749,N_6875);
xnor U10624 (N_10624,N_6962,N_4810);
and U10625 (N_10625,N_7432,N_7740);
and U10626 (N_10626,N_6081,N_5636);
nand U10627 (N_10627,N_5001,N_4556);
and U10628 (N_10628,N_7201,N_7871);
and U10629 (N_10629,N_5325,N_6643);
nand U10630 (N_10630,N_6438,N_7015);
nor U10631 (N_10631,N_6993,N_5253);
and U10632 (N_10632,N_5056,N_6914);
nand U10633 (N_10633,N_6737,N_4240);
or U10634 (N_10634,N_5636,N_7927);
nand U10635 (N_10635,N_5754,N_6214);
or U10636 (N_10636,N_5082,N_7009);
and U10637 (N_10637,N_6398,N_5466);
nand U10638 (N_10638,N_7044,N_5929);
and U10639 (N_10639,N_5124,N_6015);
or U10640 (N_10640,N_5986,N_7690);
nand U10641 (N_10641,N_7422,N_4944);
or U10642 (N_10642,N_4790,N_4114);
nor U10643 (N_10643,N_5935,N_4745);
nand U10644 (N_10644,N_7825,N_6422);
nand U10645 (N_10645,N_5854,N_5300);
nand U10646 (N_10646,N_5824,N_4821);
or U10647 (N_10647,N_7878,N_7659);
nand U10648 (N_10648,N_7507,N_4613);
and U10649 (N_10649,N_5214,N_4328);
nor U10650 (N_10650,N_7237,N_5627);
nor U10651 (N_10651,N_4948,N_4893);
or U10652 (N_10652,N_6304,N_7366);
or U10653 (N_10653,N_4328,N_6318);
nand U10654 (N_10654,N_5320,N_6445);
nand U10655 (N_10655,N_7749,N_7664);
nor U10656 (N_10656,N_5167,N_7963);
and U10657 (N_10657,N_6888,N_4078);
or U10658 (N_10658,N_6698,N_4736);
xor U10659 (N_10659,N_5537,N_7517);
and U10660 (N_10660,N_4875,N_5370);
nand U10661 (N_10661,N_5604,N_6179);
nor U10662 (N_10662,N_5988,N_4212);
or U10663 (N_10663,N_5708,N_6479);
and U10664 (N_10664,N_4937,N_4161);
nand U10665 (N_10665,N_7365,N_4248);
nand U10666 (N_10666,N_7291,N_4871);
and U10667 (N_10667,N_7242,N_6974);
nor U10668 (N_10668,N_7389,N_6111);
nor U10669 (N_10669,N_4637,N_6784);
nand U10670 (N_10670,N_6927,N_6402);
nand U10671 (N_10671,N_5268,N_4984);
nor U10672 (N_10672,N_5581,N_5253);
nor U10673 (N_10673,N_7232,N_4357);
and U10674 (N_10674,N_5306,N_4272);
nor U10675 (N_10675,N_5458,N_7355);
nor U10676 (N_10676,N_6218,N_6755);
and U10677 (N_10677,N_6879,N_6166);
and U10678 (N_10678,N_5134,N_7485);
and U10679 (N_10679,N_4440,N_6885);
nand U10680 (N_10680,N_6964,N_7865);
or U10681 (N_10681,N_5446,N_7998);
xor U10682 (N_10682,N_6707,N_5439);
xnor U10683 (N_10683,N_5000,N_4514);
xnor U10684 (N_10684,N_5855,N_6354);
xnor U10685 (N_10685,N_4675,N_4457);
or U10686 (N_10686,N_5936,N_6672);
xor U10687 (N_10687,N_4723,N_7212);
and U10688 (N_10688,N_5009,N_7784);
nor U10689 (N_10689,N_4943,N_4904);
nand U10690 (N_10690,N_4192,N_5918);
xnor U10691 (N_10691,N_6493,N_4378);
nor U10692 (N_10692,N_6341,N_6715);
nand U10693 (N_10693,N_6431,N_7633);
or U10694 (N_10694,N_4693,N_4145);
and U10695 (N_10695,N_5361,N_7299);
or U10696 (N_10696,N_6978,N_4993);
or U10697 (N_10697,N_7148,N_6947);
xor U10698 (N_10698,N_6885,N_4450);
xor U10699 (N_10699,N_5381,N_7715);
and U10700 (N_10700,N_6168,N_6200);
or U10701 (N_10701,N_5211,N_6739);
and U10702 (N_10702,N_5522,N_6760);
nor U10703 (N_10703,N_7992,N_4063);
nand U10704 (N_10704,N_7980,N_6596);
nand U10705 (N_10705,N_7931,N_6021);
or U10706 (N_10706,N_6030,N_7220);
or U10707 (N_10707,N_5848,N_7877);
or U10708 (N_10708,N_4185,N_7044);
and U10709 (N_10709,N_4879,N_5372);
nand U10710 (N_10710,N_6538,N_5262);
nor U10711 (N_10711,N_4468,N_6694);
nand U10712 (N_10712,N_5568,N_6361);
or U10713 (N_10713,N_5233,N_6898);
and U10714 (N_10714,N_5993,N_7621);
or U10715 (N_10715,N_5787,N_4441);
nor U10716 (N_10716,N_5349,N_6868);
or U10717 (N_10717,N_6430,N_5155);
nand U10718 (N_10718,N_4546,N_4649);
and U10719 (N_10719,N_5786,N_4045);
nor U10720 (N_10720,N_7486,N_5751);
and U10721 (N_10721,N_7205,N_7350);
nor U10722 (N_10722,N_4840,N_7402);
nor U10723 (N_10723,N_5343,N_5692);
nor U10724 (N_10724,N_7835,N_7755);
nand U10725 (N_10725,N_7826,N_6967);
nor U10726 (N_10726,N_6814,N_6506);
nand U10727 (N_10727,N_6280,N_7720);
and U10728 (N_10728,N_7440,N_6824);
or U10729 (N_10729,N_5314,N_4994);
nor U10730 (N_10730,N_4617,N_6882);
nor U10731 (N_10731,N_5948,N_7813);
nand U10732 (N_10732,N_6456,N_7810);
and U10733 (N_10733,N_5826,N_7773);
nand U10734 (N_10734,N_7047,N_5629);
xor U10735 (N_10735,N_7796,N_5122);
and U10736 (N_10736,N_7028,N_7900);
and U10737 (N_10737,N_6348,N_6148);
nand U10738 (N_10738,N_7462,N_5721);
nand U10739 (N_10739,N_5022,N_6156);
xor U10740 (N_10740,N_7693,N_5224);
nand U10741 (N_10741,N_4459,N_4802);
nor U10742 (N_10742,N_6061,N_5499);
nand U10743 (N_10743,N_7567,N_5933);
nand U10744 (N_10744,N_7823,N_5824);
and U10745 (N_10745,N_7132,N_6964);
or U10746 (N_10746,N_6435,N_7277);
and U10747 (N_10747,N_5613,N_6063);
nand U10748 (N_10748,N_5849,N_4839);
or U10749 (N_10749,N_5994,N_6534);
and U10750 (N_10750,N_7048,N_7098);
nor U10751 (N_10751,N_7825,N_7030);
and U10752 (N_10752,N_4506,N_6778);
nor U10753 (N_10753,N_6025,N_6685);
nor U10754 (N_10754,N_4113,N_7752);
and U10755 (N_10755,N_4353,N_4169);
and U10756 (N_10756,N_6714,N_7258);
nor U10757 (N_10757,N_7914,N_4827);
nand U10758 (N_10758,N_4756,N_4542);
nand U10759 (N_10759,N_4166,N_5794);
nor U10760 (N_10760,N_6761,N_7640);
xnor U10761 (N_10761,N_7170,N_4142);
nand U10762 (N_10762,N_4923,N_6693);
or U10763 (N_10763,N_7551,N_6169);
nor U10764 (N_10764,N_5812,N_6575);
and U10765 (N_10765,N_7241,N_6440);
and U10766 (N_10766,N_6530,N_6113);
xnor U10767 (N_10767,N_6462,N_7816);
and U10768 (N_10768,N_5615,N_4530);
and U10769 (N_10769,N_7625,N_5396);
xnor U10770 (N_10770,N_6640,N_4037);
or U10771 (N_10771,N_6941,N_4345);
nor U10772 (N_10772,N_7386,N_7622);
or U10773 (N_10773,N_4074,N_6726);
or U10774 (N_10774,N_5442,N_5283);
or U10775 (N_10775,N_4966,N_6443);
nand U10776 (N_10776,N_4561,N_4906);
or U10777 (N_10777,N_6793,N_6576);
nand U10778 (N_10778,N_4591,N_6638);
or U10779 (N_10779,N_5118,N_5502);
and U10780 (N_10780,N_7031,N_4940);
nand U10781 (N_10781,N_4013,N_6655);
and U10782 (N_10782,N_5583,N_4023);
xor U10783 (N_10783,N_6568,N_5749);
and U10784 (N_10784,N_4073,N_7091);
nand U10785 (N_10785,N_6186,N_4773);
nor U10786 (N_10786,N_4454,N_5428);
nor U10787 (N_10787,N_5916,N_5474);
nor U10788 (N_10788,N_5328,N_6947);
xnor U10789 (N_10789,N_6949,N_5976);
and U10790 (N_10790,N_5648,N_7168);
xor U10791 (N_10791,N_7370,N_4570);
nand U10792 (N_10792,N_4674,N_7173);
nor U10793 (N_10793,N_4955,N_5129);
xor U10794 (N_10794,N_7590,N_5438);
xnor U10795 (N_10795,N_7233,N_6048);
or U10796 (N_10796,N_5702,N_5666);
or U10797 (N_10797,N_4546,N_5293);
or U10798 (N_10798,N_5333,N_5634);
and U10799 (N_10799,N_7831,N_5795);
or U10800 (N_10800,N_6464,N_5742);
nand U10801 (N_10801,N_4604,N_4941);
nor U10802 (N_10802,N_7174,N_4179);
nand U10803 (N_10803,N_6794,N_5306);
and U10804 (N_10804,N_7281,N_6726);
nand U10805 (N_10805,N_4992,N_7384);
or U10806 (N_10806,N_7804,N_6508);
xor U10807 (N_10807,N_6947,N_7087);
or U10808 (N_10808,N_7811,N_4531);
nand U10809 (N_10809,N_7412,N_7767);
nand U10810 (N_10810,N_5408,N_4983);
or U10811 (N_10811,N_5299,N_7519);
nor U10812 (N_10812,N_6529,N_7357);
and U10813 (N_10813,N_4540,N_7227);
and U10814 (N_10814,N_7713,N_7036);
or U10815 (N_10815,N_5307,N_4105);
and U10816 (N_10816,N_5090,N_4623);
xnor U10817 (N_10817,N_6066,N_6121);
nor U10818 (N_10818,N_7337,N_7466);
xor U10819 (N_10819,N_4602,N_4769);
nor U10820 (N_10820,N_7917,N_7524);
xnor U10821 (N_10821,N_7329,N_5542);
nor U10822 (N_10822,N_7320,N_7988);
and U10823 (N_10823,N_7876,N_6392);
xor U10824 (N_10824,N_4740,N_7093);
nand U10825 (N_10825,N_5536,N_7559);
or U10826 (N_10826,N_4815,N_4751);
xor U10827 (N_10827,N_7510,N_4022);
or U10828 (N_10828,N_5796,N_7164);
xor U10829 (N_10829,N_7027,N_4023);
and U10830 (N_10830,N_6347,N_4891);
xnor U10831 (N_10831,N_5185,N_6581);
and U10832 (N_10832,N_7800,N_7873);
nand U10833 (N_10833,N_6378,N_6995);
nand U10834 (N_10834,N_5051,N_7446);
and U10835 (N_10835,N_7083,N_4119);
nor U10836 (N_10836,N_5162,N_6208);
nor U10837 (N_10837,N_4938,N_7458);
nand U10838 (N_10838,N_4801,N_7082);
nand U10839 (N_10839,N_5123,N_4783);
nor U10840 (N_10840,N_5796,N_4057);
nand U10841 (N_10841,N_4759,N_5439);
nand U10842 (N_10842,N_4812,N_7121);
or U10843 (N_10843,N_5047,N_5910);
and U10844 (N_10844,N_7351,N_6393);
nand U10845 (N_10845,N_6424,N_7474);
or U10846 (N_10846,N_5081,N_4724);
nand U10847 (N_10847,N_6098,N_4052);
nor U10848 (N_10848,N_7278,N_5918);
or U10849 (N_10849,N_6254,N_6756);
and U10850 (N_10850,N_7747,N_4660);
and U10851 (N_10851,N_4459,N_4066);
nand U10852 (N_10852,N_5931,N_7020);
nor U10853 (N_10853,N_5245,N_4078);
nor U10854 (N_10854,N_4995,N_4604);
nand U10855 (N_10855,N_7128,N_6662);
or U10856 (N_10856,N_5000,N_6956);
nand U10857 (N_10857,N_6867,N_6476);
and U10858 (N_10858,N_5620,N_5659);
or U10859 (N_10859,N_7105,N_5238);
nand U10860 (N_10860,N_4122,N_6159);
nand U10861 (N_10861,N_4064,N_6850);
xnor U10862 (N_10862,N_6389,N_5033);
nand U10863 (N_10863,N_4004,N_4675);
xor U10864 (N_10864,N_7990,N_4555);
xor U10865 (N_10865,N_5866,N_5031);
or U10866 (N_10866,N_5646,N_5027);
nor U10867 (N_10867,N_4443,N_6134);
and U10868 (N_10868,N_5817,N_6966);
or U10869 (N_10869,N_6733,N_4251);
nand U10870 (N_10870,N_6871,N_4216);
xnor U10871 (N_10871,N_7978,N_6380);
nand U10872 (N_10872,N_7784,N_6833);
or U10873 (N_10873,N_5157,N_4049);
or U10874 (N_10874,N_5214,N_4111);
nand U10875 (N_10875,N_5424,N_5107);
or U10876 (N_10876,N_7571,N_4722);
nand U10877 (N_10877,N_5748,N_6121);
nor U10878 (N_10878,N_6458,N_7306);
nor U10879 (N_10879,N_7756,N_4914);
xnor U10880 (N_10880,N_7769,N_6488);
nor U10881 (N_10881,N_4397,N_5304);
nor U10882 (N_10882,N_5529,N_7473);
nor U10883 (N_10883,N_5149,N_5914);
or U10884 (N_10884,N_4501,N_7866);
nand U10885 (N_10885,N_5115,N_5615);
and U10886 (N_10886,N_6822,N_4779);
nand U10887 (N_10887,N_7341,N_4312);
nor U10888 (N_10888,N_5344,N_6135);
nand U10889 (N_10889,N_7688,N_6584);
and U10890 (N_10890,N_7708,N_4997);
nor U10891 (N_10891,N_4447,N_5291);
and U10892 (N_10892,N_4829,N_6205);
or U10893 (N_10893,N_7387,N_5389);
or U10894 (N_10894,N_5280,N_6041);
or U10895 (N_10895,N_4996,N_4865);
or U10896 (N_10896,N_7273,N_4887);
or U10897 (N_10897,N_5037,N_7454);
xnor U10898 (N_10898,N_4869,N_5424);
nor U10899 (N_10899,N_4425,N_4157);
and U10900 (N_10900,N_7183,N_6286);
or U10901 (N_10901,N_6731,N_4281);
nor U10902 (N_10902,N_6578,N_4301);
nor U10903 (N_10903,N_7070,N_7682);
xnor U10904 (N_10904,N_5444,N_6636);
xor U10905 (N_10905,N_5570,N_4902);
and U10906 (N_10906,N_5710,N_7059);
and U10907 (N_10907,N_4844,N_4190);
and U10908 (N_10908,N_7911,N_5447);
and U10909 (N_10909,N_7694,N_5106);
nand U10910 (N_10910,N_4900,N_6574);
nor U10911 (N_10911,N_6473,N_7630);
or U10912 (N_10912,N_7232,N_4400);
and U10913 (N_10913,N_6681,N_4687);
and U10914 (N_10914,N_4106,N_6433);
xor U10915 (N_10915,N_7195,N_4908);
nand U10916 (N_10916,N_4141,N_4987);
or U10917 (N_10917,N_4704,N_6393);
nor U10918 (N_10918,N_6743,N_6276);
or U10919 (N_10919,N_7433,N_7127);
and U10920 (N_10920,N_6782,N_4532);
or U10921 (N_10921,N_5695,N_7664);
xnor U10922 (N_10922,N_4178,N_7957);
or U10923 (N_10923,N_5271,N_6554);
xor U10924 (N_10924,N_4910,N_5275);
and U10925 (N_10925,N_6369,N_7503);
or U10926 (N_10926,N_7821,N_5531);
nand U10927 (N_10927,N_4316,N_5245);
nor U10928 (N_10928,N_4031,N_5839);
xnor U10929 (N_10929,N_6583,N_4786);
nand U10930 (N_10930,N_7860,N_7987);
or U10931 (N_10931,N_7182,N_4771);
nor U10932 (N_10932,N_6800,N_6124);
xor U10933 (N_10933,N_5135,N_6606);
and U10934 (N_10934,N_4179,N_7490);
or U10935 (N_10935,N_6730,N_5149);
or U10936 (N_10936,N_4970,N_6376);
or U10937 (N_10937,N_4320,N_6951);
or U10938 (N_10938,N_6109,N_4794);
and U10939 (N_10939,N_6205,N_5173);
nor U10940 (N_10940,N_4956,N_6297);
nand U10941 (N_10941,N_7686,N_7509);
and U10942 (N_10942,N_6675,N_6256);
nand U10943 (N_10943,N_5265,N_4399);
xnor U10944 (N_10944,N_5973,N_7604);
or U10945 (N_10945,N_5629,N_6557);
or U10946 (N_10946,N_6778,N_6729);
xnor U10947 (N_10947,N_4675,N_4107);
nor U10948 (N_10948,N_5200,N_5768);
and U10949 (N_10949,N_4928,N_5975);
nand U10950 (N_10950,N_5237,N_4701);
or U10951 (N_10951,N_4958,N_4029);
nand U10952 (N_10952,N_5014,N_5989);
nor U10953 (N_10953,N_6334,N_4348);
nor U10954 (N_10954,N_7322,N_5477);
xor U10955 (N_10955,N_5913,N_5500);
nor U10956 (N_10956,N_4948,N_6030);
nor U10957 (N_10957,N_5123,N_5700);
nand U10958 (N_10958,N_7288,N_5532);
nor U10959 (N_10959,N_4307,N_6431);
nor U10960 (N_10960,N_6845,N_5285);
nand U10961 (N_10961,N_7152,N_4207);
nor U10962 (N_10962,N_6847,N_6540);
nand U10963 (N_10963,N_4268,N_7903);
nor U10964 (N_10964,N_6299,N_5566);
nor U10965 (N_10965,N_7435,N_7424);
nand U10966 (N_10966,N_7453,N_5632);
nand U10967 (N_10967,N_4040,N_5942);
nand U10968 (N_10968,N_4245,N_4644);
or U10969 (N_10969,N_4609,N_7594);
or U10970 (N_10970,N_6492,N_6528);
or U10971 (N_10971,N_6732,N_6179);
nor U10972 (N_10972,N_6706,N_7590);
and U10973 (N_10973,N_7012,N_6151);
nor U10974 (N_10974,N_4021,N_7900);
nor U10975 (N_10975,N_4613,N_7374);
nor U10976 (N_10976,N_6592,N_6442);
nand U10977 (N_10977,N_5262,N_5195);
and U10978 (N_10978,N_4418,N_5972);
or U10979 (N_10979,N_7489,N_5145);
nand U10980 (N_10980,N_4173,N_6027);
nor U10981 (N_10981,N_7018,N_5778);
nor U10982 (N_10982,N_4623,N_4689);
nor U10983 (N_10983,N_7275,N_7182);
and U10984 (N_10984,N_4384,N_6013);
or U10985 (N_10985,N_6366,N_4567);
and U10986 (N_10986,N_4727,N_4964);
or U10987 (N_10987,N_5663,N_5413);
or U10988 (N_10988,N_4176,N_7799);
nand U10989 (N_10989,N_7241,N_7410);
nand U10990 (N_10990,N_5007,N_7581);
nor U10991 (N_10991,N_4818,N_5482);
and U10992 (N_10992,N_7330,N_6194);
or U10993 (N_10993,N_4843,N_7409);
or U10994 (N_10994,N_5697,N_4993);
nor U10995 (N_10995,N_6958,N_4002);
and U10996 (N_10996,N_5378,N_4475);
xor U10997 (N_10997,N_6949,N_4088);
or U10998 (N_10998,N_6950,N_6562);
or U10999 (N_10999,N_7055,N_4026);
nor U11000 (N_11000,N_4646,N_5094);
nor U11001 (N_11001,N_4851,N_4700);
nor U11002 (N_11002,N_7563,N_7504);
or U11003 (N_11003,N_5999,N_4797);
and U11004 (N_11004,N_5023,N_6986);
or U11005 (N_11005,N_6759,N_6899);
and U11006 (N_11006,N_7929,N_7953);
nor U11007 (N_11007,N_6524,N_5452);
and U11008 (N_11008,N_4881,N_6694);
nand U11009 (N_11009,N_6614,N_7776);
or U11010 (N_11010,N_6513,N_4822);
xor U11011 (N_11011,N_7201,N_6915);
or U11012 (N_11012,N_5587,N_6791);
and U11013 (N_11013,N_5008,N_5976);
nor U11014 (N_11014,N_4954,N_7612);
nand U11015 (N_11015,N_7086,N_4920);
nand U11016 (N_11016,N_7635,N_5905);
or U11017 (N_11017,N_5866,N_4905);
and U11018 (N_11018,N_5606,N_4818);
nor U11019 (N_11019,N_4959,N_4665);
or U11020 (N_11020,N_5523,N_5318);
xnor U11021 (N_11021,N_4576,N_4736);
or U11022 (N_11022,N_6284,N_6170);
xnor U11023 (N_11023,N_6546,N_6519);
nand U11024 (N_11024,N_5978,N_4316);
and U11025 (N_11025,N_6577,N_5395);
or U11026 (N_11026,N_4274,N_7815);
or U11027 (N_11027,N_7259,N_5266);
or U11028 (N_11028,N_4708,N_6027);
or U11029 (N_11029,N_6239,N_4535);
and U11030 (N_11030,N_6856,N_5570);
nor U11031 (N_11031,N_4552,N_4511);
nor U11032 (N_11032,N_6857,N_4098);
nand U11033 (N_11033,N_6118,N_7918);
or U11034 (N_11034,N_7145,N_6759);
nand U11035 (N_11035,N_6169,N_6073);
or U11036 (N_11036,N_5065,N_4708);
nor U11037 (N_11037,N_4679,N_7068);
or U11038 (N_11038,N_6734,N_7694);
or U11039 (N_11039,N_4091,N_4731);
nand U11040 (N_11040,N_6924,N_4776);
or U11041 (N_11041,N_7890,N_7306);
nand U11042 (N_11042,N_7968,N_7361);
nand U11043 (N_11043,N_4723,N_5664);
or U11044 (N_11044,N_7451,N_6535);
or U11045 (N_11045,N_7641,N_4440);
or U11046 (N_11046,N_7913,N_4538);
nand U11047 (N_11047,N_6543,N_6834);
and U11048 (N_11048,N_4723,N_6777);
or U11049 (N_11049,N_4608,N_4784);
or U11050 (N_11050,N_5259,N_7607);
nand U11051 (N_11051,N_6317,N_5322);
nand U11052 (N_11052,N_5800,N_4577);
and U11053 (N_11053,N_6866,N_7956);
nor U11054 (N_11054,N_5954,N_4093);
xnor U11055 (N_11055,N_6915,N_5013);
nor U11056 (N_11056,N_7405,N_4105);
nor U11057 (N_11057,N_6798,N_4338);
nor U11058 (N_11058,N_5229,N_4673);
nand U11059 (N_11059,N_7423,N_6995);
nand U11060 (N_11060,N_7630,N_4312);
nor U11061 (N_11061,N_4521,N_7670);
or U11062 (N_11062,N_7463,N_7568);
nand U11063 (N_11063,N_4297,N_4267);
or U11064 (N_11064,N_6800,N_5929);
nand U11065 (N_11065,N_7104,N_5521);
nand U11066 (N_11066,N_4872,N_5250);
nand U11067 (N_11067,N_4283,N_5476);
and U11068 (N_11068,N_5661,N_4174);
and U11069 (N_11069,N_5003,N_5727);
nor U11070 (N_11070,N_6193,N_5869);
nor U11071 (N_11071,N_5930,N_6217);
xnor U11072 (N_11072,N_6479,N_4698);
nand U11073 (N_11073,N_6475,N_5035);
and U11074 (N_11074,N_7091,N_6985);
and U11075 (N_11075,N_4052,N_7335);
nor U11076 (N_11076,N_4962,N_5690);
nand U11077 (N_11077,N_7929,N_4904);
nor U11078 (N_11078,N_4265,N_6180);
and U11079 (N_11079,N_7657,N_7852);
nor U11080 (N_11080,N_6193,N_7541);
and U11081 (N_11081,N_6509,N_7440);
nand U11082 (N_11082,N_5910,N_5644);
and U11083 (N_11083,N_7944,N_7001);
or U11084 (N_11084,N_6048,N_7877);
or U11085 (N_11085,N_7583,N_6850);
nor U11086 (N_11086,N_7225,N_4511);
or U11087 (N_11087,N_5911,N_5792);
or U11088 (N_11088,N_5003,N_4937);
nor U11089 (N_11089,N_7985,N_5621);
nor U11090 (N_11090,N_7866,N_6482);
and U11091 (N_11091,N_7200,N_7703);
xnor U11092 (N_11092,N_6545,N_5453);
nand U11093 (N_11093,N_4792,N_4556);
xor U11094 (N_11094,N_6759,N_5556);
nor U11095 (N_11095,N_7123,N_6970);
nand U11096 (N_11096,N_7810,N_5462);
or U11097 (N_11097,N_6588,N_7229);
nor U11098 (N_11098,N_5070,N_5541);
nand U11099 (N_11099,N_7843,N_7015);
or U11100 (N_11100,N_6975,N_6174);
xnor U11101 (N_11101,N_4240,N_6812);
nor U11102 (N_11102,N_4171,N_6494);
or U11103 (N_11103,N_6063,N_4758);
nand U11104 (N_11104,N_6788,N_6793);
or U11105 (N_11105,N_5292,N_4648);
or U11106 (N_11106,N_5184,N_4742);
and U11107 (N_11107,N_6431,N_5049);
or U11108 (N_11108,N_5265,N_4975);
nor U11109 (N_11109,N_7275,N_7466);
nor U11110 (N_11110,N_4702,N_6974);
nand U11111 (N_11111,N_5218,N_6219);
nor U11112 (N_11112,N_4251,N_7021);
or U11113 (N_11113,N_7292,N_4822);
or U11114 (N_11114,N_4182,N_4812);
nor U11115 (N_11115,N_6983,N_4778);
or U11116 (N_11116,N_7587,N_7522);
nand U11117 (N_11117,N_6557,N_5514);
or U11118 (N_11118,N_5782,N_7679);
nand U11119 (N_11119,N_5858,N_6362);
nand U11120 (N_11120,N_4563,N_5525);
or U11121 (N_11121,N_7757,N_4600);
nor U11122 (N_11122,N_5138,N_5866);
nand U11123 (N_11123,N_6646,N_5271);
nor U11124 (N_11124,N_6088,N_5325);
xnor U11125 (N_11125,N_7210,N_5679);
and U11126 (N_11126,N_4186,N_4996);
or U11127 (N_11127,N_6485,N_6497);
or U11128 (N_11128,N_7411,N_4423);
and U11129 (N_11129,N_5263,N_5949);
xor U11130 (N_11130,N_5354,N_6193);
and U11131 (N_11131,N_5431,N_6277);
or U11132 (N_11132,N_6666,N_6814);
and U11133 (N_11133,N_4879,N_6512);
nand U11134 (N_11134,N_7596,N_7534);
or U11135 (N_11135,N_4005,N_4783);
nand U11136 (N_11136,N_5863,N_7766);
and U11137 (N_11137,N_4328,N_5614);
and U11138 (N_11138,N_5814,N_7907);
nand U11139 (N_11139,N_7983,N_5487);
nor U11140 (N_11140,N_4073,N_5048);
and U11141 (N_11141,N_4197,N_6964);
or U11142 (N_11142,N_5239,N_7076);
or U11143 (N_11143,N_6081,N_7143);
or U11144 (N_11144,N_5475,N_7548);
nand U11145 (N_11145,N_6206,N_5923);
and U11146 (N_11146,N_7663,N_5589);
nand U11147 (N_11147,N_7806,N_5189);
nand U11148 (N_11148,N_4927,N_7893);
xnor U11149 (N_11149,N_5472,N_7333);
nor U11150 (N_11150,N_5178,N_5962);
xor U11151 (N_11151,N_6280,N_5734);
nor U11152 (N_11152,N_7893,N_6570);
nor U11153 (N_11153,N_4538,N_4406);
or U11154 (N_11154,N_7180,N_4753);
xor U11155 (N_11155,N_5474,N_7130);
nand U11156 (N_11156,N_7686,N_6188);
and U11157 (N_11157,N_4812,N_5224);
nor U11158 (N_11158,N_6162,N_7401);
and U11159 (N_11159,N_5648,N_7500);
or U11160 (N_11160,N_5164,N_4665);
nand U11161 (N_11161,N_4696,N_5511);
nand U11162 (N_11162,N_6624,N_4699);
nor U11163 (N_11163,N_4212,N_5103);
or U11164 (N_11164,N_5124,N_7892);
nor U11165 (N_11165,N_5845,N_6702);
nor U11166 (N_11166,N_7731,N_6806);
and U11167 (N_11167,N_5811,N_4369);
and U11168 (N_11168,N_5886,N_5195);
nor U11169 (N_11169,N_7362,N_6776);
or U11170 (N_11170,N_4674,N_5340);
and U11171 (N_11171,N_7612,N_7266);
and U11172 (N_11172,N_5259,N_7208);
xnor U11173 (N_11173,N_7666,N_5858);
or U11174 (N_11174,N_7614,N_5441);
nor U11175 (N_11175,N_4325,N_7068);
nand U11176 (N_11176,N_4893,N_4468);
or U11177 (N_11177,N_6456,N_4149);
nand U11178 (N_11178,N_6080,N_4765);
nor U11179 (N_11179,N_7488,N_4747);
or U11180 (N_11180,N_7524,N_7491);
or U11181 (N_11181,N_5409,N_7711);
and U11182 (N_11182,N_4420,N_4506);
or U11183 (N_11183,N_4691,N_5778);
nor U11184 (N_11184,N_5894,N_4672);
and U11185 (N_11185,N_5102,N_4549);
nor U11186 (N_11186,N_6509,N_5695);
or U11187 (N_11187,N_7649,N_4844);
nor U11188 (N_11188,N_6985,N_4206);
nand U11189 (N_11189,N_7023,N_5944);
nor U11190 (N_11190,N_6416,N_5864);
nor U11191 (N_11191,N_4690,N_6913);
and U11192 (N_11192,N_5508,N_7915);
or U11193 (N_11193,N_4080,N_4589);
or U11194 (N_11194,N_7189,N_6493);
xnor U11195 (N_11195,N_5795,N_4881);
nand U11196 (N_11196,N_7898,N_6213);
and U11197 (N_11197,N_4177,N_6863);
and U11198 (N_11198,N_5271,N_5213);
xnor U11199 (N_11199,N_4997,N_4628);
xor U11200 (N_11200,N_4118,N_5699);
or U11201 (N_11201,N_4500,N_4993);
nand U11202 (N_11202,N_7037,N_7179);
nor U11203 (N_11203,N_5183,N_7006);
nor U11204 (N_11204,N_6530,N_4694);
nand U11205 (N_11205,N_6703,N_6739);
and U11206 (N_11206,N_6818,N_5778);
and U11207 (N_11207,N_4369,N_4048);
or U11208 (N_11208,N_6810,N_5039);
or U11209 (N_11209,N_6002,N_4715);
or U11210 (N_11210,N_4803,N_7677);
and U11211 (N_11211,N_4824,N_5683);
nand U11212 (N_11212,N_6909,N_6756);
nand U11213 (N_11213,N_5788,N_4937);
or U11214 (N_11214,N_7145,N_6937);
nand U11215 (N_11215,N_7110,N_5373);
and U11216 (N_11216,N_5340,N_4798);
and U11217 (N_11217,N_5611,N_7452);
xor U11218 (N_11218,N_5997,N_6106);
xnor U11219 (N_11219,N_7757,N_4067);
or U11220 (N_11220,N_7073,N_5323);
nand U11221 (N_11221,N_4921,N_6945);
and U11222 (N_11222,N_7367,N_7810);
xor U11223 (N_11223,N_7225,N_7667);
and U11224 (N_11224,N_4355,N_5676);
and U11225 (N_11225,N_7089,N_6959);
nor U11226 (N_11226,N_5300,N_4357);
and U11227 (N_11227,N_4649,N_5686);
or U11228 (N_11228,N_7722,N_5381);
nor U11229 (N_11229,N_6595,N_4330);
nand U11230 (N_11230,N_6646,N_6173);
or U11231 (N_11231,N_6123,N_6135);
nand U11232 (N_11232,N_7782,N_6731);
nand U11233 (N_11233,N_7707,N_6123);
or U11234 (N_11234,N_7344,N_5115);
and U11235 (N_11235,N_4037,N_7030);
xor U11236 (N_11236,N_4125,N_7791);
xnor U11237 (N_11237,N_4158,N_5143);
or U11238 (N_11238,N_4829,N_4621);
nor U11239 (N_11239,N_4750,N_7935);
or U11240 (N_11240,N_6706,N_7494);
or U11241 (N_11241,N_4841,N_7360);
or U11242 (N_11242,N_4182,N_6326);
nor U11243 (N_11243,N_4212,N_7608);
nand U11244 (N_11244,N_6939,N_6869);
nor U11245 (N_11245,N_7278,N_7980);
xnor U11246 (N_11246,N_6211,N_6236);
and U11247 (N_11247,N_7470,N_4663);
nand U11248 (N_11248,N_4748,N_6059);
and U11249 (N_11249,N_7805,N_5708);
and U11250 (N_11250,N_4099,N_5071);
and U11251 (N_11251,N_5100,N_6393);
nor U11252 (N_11252,N_4933,N_6421);
xor U11253 (N_11253,N_7565,N_5414);
and U11254 (N_11254,N_4892,N_4101);
nor U11255 (N_11255,N_4128,N_5913);
nor U11256 (N_11256,N_5703,N_5714);
nor U11257 (N_11257,N_4775,N_5382);
and U11258 (N_11258,N_5375,N_7932);
and U11259 (N_11259,N_5285,N_4604);
nor U11260 (N_11260,N_7338,N_6636);
and U11261 (N_11261,N_4076,N_4812);
nand U11262 (N_11262,N_7433,N_6204);
nand U11263 (N_11263,N_6298,N_7655);
nor U11264 (N_11264,N_5987,N_6721);
and U11265 (N_11265,N_7442,N_6533);
nand U11266 (N_11266,N_4318,N_4015);
nand U11267 (N_11267,N_5670,N_6165);
nand U11268 (N_11268,N_6906,N_7057);
nand U11269 (N_11269,N_6463,N_7634);
and U11270 (N_11270,N_4067,N_6092);
and U11271 (N_11271,N_5577,N_7613);
or U11272 (N_11272,N_4813,N_4377);
nand U11273 (N_11273,N_6405,N_4828);
and U11274 (N_11274,N_6694,N_4738);
nand U11275 (N_11275,N_5682,N_7564);
and U11276 (N_11276,N_7928,N_4026);
and U11277 (N_11277,N_6108,N_5104);
or U11278 (N_11278,N_6025,N_5641);
or U11279 (N_11279,N_7515,N_7076);
and U11280 (N_11280,N_4488,N_5725);
or U11281 (N_11281,N_6843,N_5235);
nor U11282 (N_11282,N_4960,N_6651);
and U11283 (N_11283,N_6548,N_5688);
xnor U11284 (N_11284,N_5170,N_7831);
nor U11285 (N_11285,N_4333,N_7562);
xnor U11286 (N_11286,N_4118,N_4138);
nand U11287 (N_11287,N_5855,N_6381);
and U11288 (N_11288,N_4509,N_7621);
nor U11289 (N_11289,N_6484,N_6307);
nor U11290 (N_11290,N_5707,N_6723);
or U11291 (N_11291,N_6148,N_7712);
and U11292 (N_11292,N_6511,N_5188);
nand U11293 (N_11293,N_4084,N_6942);
nor U11294 (N_11294,N_4312,N_4287);
nor U11295 (N_11295,N_6340,N_5374);
or U11296 (N_11296,N_6222,N_4442);
or U11297 (N_11297,N_5346,N_6321);
and U11298 (N_11298,N_7935,N_6788);
and U11299 (N_11299,N_4598,N_7708);
nor U11300 (N_11300,N_5530,N_5843);
and U11301 (N_11301,N_6710,N_4467);
nor U11302 (N_11302,N_5725,N_5269);
nor U11303 (N_11303,N_6017,N_6744);
nand U11304 (N_11304,N_6586,N_4720);
and U11305 (N_11305,N_7183,N_5569);
or U11306 (N_11306,N_7961,N_7883);
nand U11307 (N_11307,N_5385,N_5340);
or U11308 (N_11308,N_7466,N_7583);
or U11309 (N_11309,N_6452,N_4824);
and U11310 (N_11310,N_4033,N_6113);
nor U11311 (N_11311,N_7822,N_6728);
nand U11312 (N_11312,N_7538,N_4473);
or U11313 (N_11313,N_6404,N_6681);
or U11314 (N_11314,N_7568,N_7484);
nor U11315 (N_11315,N_4226,N_4020);
or U11316 (N_11316,N_4624,N_4984);
nor U11317 (N_11317,N_4356,N_6752);
nand U11318 (N_11318,N_7060,N_7446);
nor U11319 (N_11319,N_5712,N_7316);
nor U11320 (N_11320,N_6091,N_4889);
nand U11321 (N_11321,N_4184,N_7243);
nand U11322 (N_11322,N_5579,N_5212);
or U11323 (N_11323,N_6303,N_4164);
xnor U11324 (N_11324,N_6984,N_4776);
nand U11325 (N_11325,N_6312,N_7788);
nand U11326 (N_11326,N_7596,N_7227);
nand U11327 (N_11327,N_4079,N_5558);
nor U11328 (N_11328,N_5530,N_4491);
or U11329 (N_11329,N_5788,N_7757);
and U11330 (N_11330,N_6657,N_4770);
nor U11331 (N_11331,N_6887,N_6404);
or U11332 (N_11332,N_4475,N_6539);
or U11333 (N_11333,N_5508,N_4636);
nor U11334 (N_11334,N_6058,N_5536);
xor U11335 (N_11335,N_7294,N_4718);
or U11336 (N_11336,N_7663,N_7737);
or U11337 (N_11337,N_5352,N_5948);
nand U11338 (N_11338,N_7160,N_6948);
nor U11339 (N_11339,N_5282,N_5923);
or U11340 (N_11340,N_7992,N_6813);
nand U11341 (N_11341,N_5608,N_7410);
nand U11342 (N_11342,N_7897,N_5581);
nand U11343 (N_11343,N_7329,N_5207);
nand U11344 (N_11344,N_6617,N_6878);
nand U11345 (N_11345,N_4934,N_6195);
or U11346 (N_11346,N_7298,N_5776);
or U11347 (N_11347,N_7413,N_5983);
nand U11348 (N_11348,N_7597,N_4686);
nor U11349 (N_11349,N_5640,N_4167);
nor U11350 (N_11350,N_4238,N_5505);
nand U11351 (N_11351,N_4903,N_7937);
xnor U11352 (N_11352,N_6525,N_5859);
and U11353 (N_11353,N_7258,N_5879);
nor U11354 (N_11354,N_6133,N_4867);
nand U11355 (N_11355,N_5946,N_4010);
nand U11356 (N_11356,N_7464,N_6184);
or U11357 (N_11357,N_5910,N_4895);
or U11358 (N_11358,N_6328,N_7306);
nor U11359 (N_11359,N_6665,N_5890);
or U11360 (N_11360,N_6859,N_4244);
and U11361 (N_11361,N_6110,N_5548);
xnor U11362 (N_11362,N_4775,N_7162);
or U11363 (N_11363,N_4764,N_5291);
and U11364 (N_11364,N_6471,N_4307);
or U11365 (N_11365,N_6845,N_7769);
nor U11366 (N_11366,N_5541,N_7277);
and U11367 (N_11367,N_5996,N_7327);
and U11368 (N_11368,N_7242,N_6131);
and U11369 (N_11369,N_4241,N_5735);
nor U11370 (N_11370,N_6457,N_5078);
and U11371 (N_11371,N_7154,N_6319);
or U11372 (N_11372,N_7981,N_6097);
and U11373 (N_11373,N_7271,N_4902);
nand U11374 (N_11374,N_5028,N_7712);
xnor U11375 (N_11375,N_5601,N_5023);
nand U11376 (N_11376,N_6403,N_4235);
nor U11377 (N_11377,N_6456,N_5787);
nor U11378 (N_11378,N_7687,N_7346);
or U11379 (N_11379,N_6405,N_5759);
and U11380 (N_11380,N_4879,N_6482);
and U11381 (N_11381,N_6775,N_6365);
or U11382 (N_11382,N_6861,N_4145);
nor U11383 (N_11383,N_4235,N_7777);
or U11384 (N_11384,N_7351,N_4501);
nand U11385 (N_11385,N_7110,N_6161);
nand U11386 (N_11386,N_5692,N_4386);
or U11387 (N_11387,N_5553,N_6846);
nor U11388 (N_11388,N_7295,N_7428);
or U11389 (N_11389,N_7330,N_7064);
xnor U11390 (N_11390,N_7571,N_4879);
and U11391 (N_11391,N_5029,N_5787);
nor U11392 (N_11392,N_6587,N_6793);
nand U11393 (N_11393,N_4313,N_7680);
nor U11394 (N_11394,N_6566,N_5497);
nor U11395 (N_11395,N_6024,N_7204);
nor U11396 (N_11396,N_5398,N_4760);
nor U11397 (N_11397,N_4002,N_7019);
xor U11398 (N_11398,N_5417,N_4826);
nor U11399 (N_11399,N_7729,N_4505);
nand U11400 (N_11400,N_7251,N_5668);
and U11401 (N_11401,N_6565,N_5380);
and U11402 (N_11402,N_7424,N_4268);
and U11403 (N_11403,N_5038,N_7055);
and U11404 (N_11404,N_6978,N_4446);
nor U11405 (N_11405,N_6544,N_5700);
nand U11406 (N_11406,N_5698,N_5533);
or U11407 (N_11407,N_5639,N_6140);
nor U11408 (N_11408,N_4342,N_5775);
or U11409 (N_11409,N_6192,N_6304);
nor U11410 (N_11410,N_7632,N_4675);
nand U11411 (N_11411,N_6269,N_5192);
or U11412 (N_11412,N_4583,N_5344);
nand U11413 (N_11413,N_5443,N_7635);
or U11414 (N_11414,N_6485,N_5733);
or U11415 (N_11415,N_7435,N_5159);
nand U11416 (N_11416,N_5399,N_7984);
nand U11417 (N_11417,N_4446,N_6901);
or U11418 (N_11418,N_4150,N_7471);
or U11419 (N_11419,N_5339,N_7197);
or U11420 (N_11420,N_5578,N_6738);
and U11421 (N_11421,N_4626,N_6969);
and U11422 (N_11422,N_6307,N_6767);
nor U11423 (N_11423,N_6200,N_4834);
and U11424 (N_11424,N_7876,N_7522);
or U11425 (N_11425,N_6516,N_4140);
or U11426 (N_11426,N_4594,N_7068);
and U11427 (N_11427,N_6211,N_4217);
and U11428 (N_11428,N_6967,N_5712);
or U11429 (N_11429,N_5011,N_5425);
and U11430 (N_11430,N_4137,N_5305);
or U11431 (N_11431,N_4164,N_5607);
or U11432 (N_11432,N_4075,N_5870);
nor U11433 (N_11433,N_7981,N_6199);
nand U11434 (N_11434,N_4659,N_4703);
or U11435 (N_11435,N_5490,N_7522);
nand U11436 (N_11436,N_4006,N_6527);
nand U11437 (N_11437,N_5524,N_4849);
or U11438 (N_11438,N_5221,N_5625);
and U11439 (N_11439,N_6762,N_6381);
nor U11440 (N_11440,N_6767,N_6335);
or U11441 (N_11441,N_4122,N_7826);
nor U11442 (N_11442,N_7535,N_7906);
or U11443 (N_11443,N_4654,N_5292);
nor U11444 (N_11444,N_7389,N_4873);
or U11445 (N_11445,N_6134,N_6449);
and U11446 (N_11446,N_5399,N_7031);
nand U11447 (N_11447,N_7752,N_4051);
and U11448 (N_11448,N_5956,N_7005);
xor U11449 (N_11449,N_4369,N_4300);
nand U11450 (N_11450,N_6369,N_4017);
and U11451 (N_11451,N_5495,N_5001);
xnor U11452 (N_11452,N_4236,N_7879);
nand U11453 (N_11453,N_4248,N_7992);
and U11454 (N_11454,N_4333,N_5203);
or U11455 (N_11455,N_5712,N_5917);
xor U11456 (N_11456,N_5588,N_6257);
nor U11457 (N_11457,N_6910,N_5236);
nand U11458 (N_11458,N_7534,N_7759);
nor U11459 (N_11459,N_5618,N_4248);
nand U11460 (N_11460,N_5350,N_5700);
xor U11461 (N_11461,N_6919,N_6359);
nand U11462 (N_11462,N_7516,N_7168);
nand U11463 (N_11463,N_5665,N_6250);
nor U11464 (N_11464,N_6663,N_4198);
nor U11465 (N_11465,N_7909,N_5784);
nor U11466 (N_11466,N_6256,N_6605);
xnor U11467 (N_11467,N_7089,N_6415);
and U11468 (N_11468,N_5647,N_6869);
and U11469 (N_11469,N_5940,N_7179);
and U11470 (N_11470,N_7503,N_4613);
or U11471 (N_11471,N_6425,N_7315);
nor U11472 (N_11472,N_7643,N_6753);
or U11473 (N_11473,N_5121,N_7356);
nand U11474 (N_11474,N_6791,N_5901);
nor U11475 (N_11475,N_6288,N_6686);
xor U11476 (N_11476,N_6178,N_7003);
nand U11477 (N_11477,N_6832,N_4852);
or U11478 (N_11478,N_5385,N_5346);
nand U11479 (N_11479,N_5662,N_4608);
or U11480 (N_11480,N_7311,N_4181);
or U11481 (N_11481,N_7320,N_5832);
nor U11482 (N_11482,N_5370,N_6769);
nor U11483 (N_11483,N_5148,N_6201);
or U11484 (N_11484,N_4121,N_6975);
or U11485 (N_11485,N_4989,N_5805);
and U11486 (N_11486,N_5068,N_4855);
and U11487 (N_11487,N_5216,N_4865);
or U11488 (N_11488,N_5067,N_4413);
and U11489 (N_11489,N_4969,N_6956);
xnor U11490 (N_11490,N_5752,N_5379);
or U11491 (N_11491,N_6453,N_7086);
nor U11492 (N_11492,N_7851,N_6293);
or U11493 (N_11493,N_6745,N_4051);
and U11494 (N_11494,N_4328,N_4411);
or U11495 (N_11495,N_6769,N_4739);
nand U11496 (N_11496,N_4837,N_7876);
and U11497 (N_11497,N_6564,N_5126);
nand U11498 (N_11498,N_5879,N_7439);
or U11499 (N_11499,N_5189,N_7197);
nor U11500 (N_11500,N_4657,N_4725);
and U11501 (N_11501,N_6902,N_5631);
and U11502 (N_11502,N_5672,N_4310);
nor U11503 (N_11503,N_4445,N_7816);
xor U11504 (N_11504,N_6617,N_4072);
nand U11505 (N_11505,N_4931,N_4108);
nor U11506 (N_11506,N_5111,N_4613);
nand U11507 (N_11507,N_7556,N_5975);
or U11508 (N_11508,N_7575,N_6773);
nand U11509 (N_11509,N_4608,N_6884);
and U11510 (N_11510,N_7983,N_4619);
nand U11511 (N_11511,N_7384,N_5626);
nor U11512 (N_11512,N_4766,N_5604);
nor U11513 (N_11513,N_4991,N_5963);
nor U11514 (N_11514,N_7931,N_4024);
nand U11515 (N_11515,N_6128,N_6931);
or U11516 (N_11516,N_4475,N_6826);
nor U11517 (N_11517,N_7715,N_6095);
nor U11518 (N_11518,N_5496,N_6887);
nor U11519 (N_11519,N_5955,N_6400);
or U11520 (N_11520,N_6631,N_6050);
xnor U11521 (N_11521,N_5437,N_6992);
xor U11522 (N_11522,N_4257,N_6808);
nor U11523 (N_11523,N_6728,N_7004);
and U11524 (N_11524,N_7849,N_6583);
nor U11525 (N_11525,N_4437,N_5274);
xor U11526 (N_11526,N_6460,N_5401);
nor U11527 (N_11527,N_7739,N_7384);
nand U11528 (N_11528,N_5947,N_6652);
xor U11529 (N_11529,N_6768,N_7610);
nand U11530 (N_11530,N_6569,N_5094);
nand U11531 (N_11531,N_4044,N_5665);
nor U11532 (N_11532,N_5405,N_5801);
nand U11533 (N_11533,N_5421,N_5098);
and U11534 (N_11534,N_4998,N_4770);
nor U11535 (N_11535,N_4132,N_5252);
nand U11536 (N_11536,N_5426,N_4681);
nand U11537 (N_11537,N_5614,N_7718);
or U11538 (N_11538,N_5999,N_7936);
and U11539 (N_11539,N_6782,N_6261);
nor U11540 (N_11540,N_7981,N_7074);
or U11541 (N_11541,N_4645,N_7984);
or U11542 (N_11542,N_6275,N_5400);
or U11543 (N_11543,N_4117,N_6876);
xor U11544 (N_11544,N_6890,N_4621);
nand U11545 (N_11545,N_7592,N_6728);
xor U11546 (N_11546,N_6825,N_6782);
and U11547 (N_11547,N_7862,N_5848);
or U11548 (N_11548,N_4547,N_7169);
nor U11549 (N_11549,N_7246,N_5546);
nor U11550 (N_11550,N_4528,N_4546);
xnor U11551 (N_11551,N_4220,N_7925);
nor U11552 (N_11552,N_4412,N_7429);
nand U11553 (N_11553,N_5532,N_5654);
and U11554 (N_11554,N_6345,N_5013);
nor U11555 (N_11555,N_5255,N_5711);
or U11556 (N_11556,N_4712,N_4152);
or U11557 (N_11557,N_6561,N_7172);
and U11558 (N_11558,N_5537,N_6956);
nor U11559 (N_11559,N_5972,N_7401);
nor U11560 (N_11560,N_7523,N_6536);
nand U11561 (N_11561,N_4237,N_6634);
or U11562 (N_11562,N_7720,N_7824);
or U11563 (N_11563,N_6348,N_5706);
nand U11564 (N_11564,N_6200,N_7356);
nor U11565 (N_11565,N_6471,N_4376);
nor U11566 (N_11566,N_4921,N_6420);
nand U11567 (N_11567,N_7525,N_5549);
nor U11568 (N_11568,N_5010,N_4672);
nand U11569 (N_11569,N_5309,N_6221);
and U11570 (N_11570,N_6361,N_6969);
xnor U11571 (N_11571,N_6712,N_5035);
nor U11572 (N_11572,N_5203,N_5841);
and U11573 (N_11573,N_5458,N_5927);
and U11574 (N_11574,N_7892,N_4771);
nor U11575 (N_11575,N_5505,N_6467);
and U11576 (N_11576,N_6934,N_7412);
and U11577 (N_11577,N_5025,N_4493);
nand U11578 (N_11578,N_6139,N_5406);
and U11579 (N_11579,N_6579,N_5331);
nor U11580 (N_11580,N_4704,N_7637);
nor U11581 (N_11581,N_5769,N_4214);
and U11582 (N_11582,N_5306,N_5258);
or U11583 (N_11583,N_6819,N_6142);
and U11584 (N_11584,N_7283,N_6295);
and U11585 (N_11585,N_7056,N_6223);
or U11586 (N_11586,N_6260,N_4754);
or U11587 (N_11587,N_4337,N_7292);
nand U11588 (N_11588,N_4274,N_7858);
nand U11589 (N_11589,N_7630,N_4445);
and U11590 (N_11590,N_6722,N_4026);
nand U11591 (N_11591,N_7468,N_4765);
and U11592 (N_11592,N_7404,N_6773);
xor U11593 (N_11593,N_6461,N_5159);
nor U11594 (N_11594,N_5691,N_6223);
or U11595 (N_11595,N_7620,N_6573);
and U11596 (N_11596,N_4027,N_6211);
nand U11597 (N_11597,N_6378,N_4525);
xor U11598 (N_11598,N_5906,N_7698);
nor U11599 (N_11599,N_4316,N_4683);
nor U11600 (N_11600,N_4163,N_7354);
nand U11601 (N_11601,N_7311,N_7761);
and U11602 (N_11602,N_4977,N_7622);
and U11603 (N_11603,N_7593,N_6959);
nand U11604 (N_11604,N_4713,N_4764);
nor U11605 (N_11605,N_6574,N_7716);
nor U11606 (N_11606,N_5564,N_7695);
nor U11607 (N_11607,N_4094,N_7958);
xnor U11608 (N_11608,N_5997,N_5164);
or U11609 (N_11609,N_6322,N_4295);
and U11610 (N_11610,N_4546,N_6032);
xor U11611 (N_11611,N_7861,N_7748);
xnor U11612 (N_11612,N_7680,N_6232);
or U11613 (N_11613,N_5614,N_7763);
nor U11614 (N_11614,N_5499,N_7414);
nor U11615 (N_11615,N_5129,N_7575);
nand U11616 (N_11616,N_4067,N_7589);
nor U11617 (N_11617,N_4295,N_5387);
nor U11618 (N_11618,N_7083,N_4060);
xnor U11619 (N_11619,N_4674,N_4444);
or U11620 (N_11620,N_6512,N_6821);
or U11621 (N_11621,N_5515,N_5482);
nor U11622 (N_11622,N_7475,N_6495);
and U11623 (N_11623,N_4943,N_6908);
or U11624 (N_11624,N_4022,N_5116);
nand U11625 (N_11625,N_7595,N_5612);
or U11626 (N_11626,N_6233,N_6606);
and U11627 (N_11627,N_4770,N_6987);
or U11628 (N_11628,N_5343,N_7012);
and U11629 (N_11629,N_7751,N_5970);
and U11630 (N_11630,N_5531,N_4225);
xor U11631 (N_11631,N_5296,N_4841);
xor U11632 (N_11632,N_7743,N_4566);
xnor U11633 (N_11633,N_4761,N_4537);
nand U11634 (N_11634,N_4719,N_7405);
nand U11635 (N_11635,N_5381,N_6514);
or U11636 (N_11636,N_6890,N_6142);
and U11637 (N_11637,N_5681,N_6286);
or U11638 (N_11638,N_5386,N_4439);
and U11639 (N_11639,N_4334,N_7987);
nor U11640 (N_11640,N_6858,N_4738);
nor U11641 (N_11641,N_7247,N_4263);
nand U11642 (N_11642,N_7852,N_4337);
xor U11643 (N_11643,N_7384,N_6165);
nor U11644 (N_11644,N_6489,N_4743);
or U11645 (N_11645,N_7928,N_7434);
nor U11646 (N_11646,N_7355,N_4100);
nand U11647 (N_11647,N_7236,N_5228);
nand U11648 (N_11648,N_5957,N_6458);
or U11649 (N_11649,N_4094,N_7069);
or U11650 (N_11650,N_6763,N_4467);
and U11651 (N_11651,N_4364,N_6550);
and U11652 (N_11652,N_4704,N_5337);
xor U11653 (N_11653,N_6302,N_7581);
nor U11654 (N_11654,N_4971,N_6815);
nor U11655 (N_11655,N_5431,N_6615);
nor U11656 (N_11656,N_4600,N_7988);
nor U11657 (N_11657,N_6920,N_5406);
nand U11658 (N_11658,N_5213,N_6975);
nor U11659 (N_11659,N_5189,N_7363);
nand U11660 (N_11660,N_6986,N_7027);
nand U11661 (N_11661,N_6315,N_7013);
or U11662 (N_11662,N_4322,N_6417);
nor U11663 (N_11663,N_5700,N_6712);
nand U11664 (N_11664,N_6560,N_4278);
and U11665 (N_11665,N_7270,N_4801);
and U11666 (N_11666,N_5333,N_4330);
nor U11667 (N_11667,N_7218,N_5587);
xor U11668 (N_11668,N_5125,N_5097);
or U11669 (N_11669,N_4456,N_6130);
nor U11670 (N_11670,N_6723,N_6372);
nor U11671 (N_11671,N_4384,N_4722);
nor U11672 (N_11672,N_4218,N_4252);
nand U11673 (N_11673,N_6083,N_7666);
xnor U11674 (N_11674,N_7625,N_6637);
or U11675 (N_11675,N_5609,N_4780);
or U11676 (N_11676,N_6279,N_5334);
and U11677 (N_11677,N_4307,N_5731);
nand U11678 (N_11678,N_4614,N_5369);
nand U11679 (N_11679,N_5215,N_5176);
or U11680 (N_11680,N_6261,N_4285);
and U11681 (N_11681,N_5116,N_7053);
nor U11682 (N_11682,N_4335,N_6884);
nand U11683 (N_11683,N_6663,N_7488);
nand U11684 (N_11684,N_7953,N_6495);
nor U11685 (N_11685,N_7376,N_5080);
or U11686 (N_11686,N_4474,N_7524);
nor U11687 (N_11687,N_4997,N_5950);
and U11688 (N_11688,N_4356,N_4392);
nor U11689 (N_11689,N_4764,N_5965);
and U11690 (N_11690,N_4129,N_6325);
and U11691 (N_11691,N_6362,N_4883);
and U11692 (N_11692,N_5190,N_7184);
and U11693 (N_11693,N_6091,N_5691);
nor U11694 (N_11694,N_6693,N_7614);
nand U11695 (N_11695,N_5618,N_7341);
nand U11696 (N_11696,N_6420,N_6918);
nand U11697 (N_11697,N_4600,N_5327);
nand U11698 (N_11698,N_4508,N_4444);
nand U11699 (N_11699,N_6652,N_7256);
nor U11700 (N_11700,N_6814,N_5614);
nor U11701 (N_11701,N_4817,N_7780);
or U11702 (N_11702,N_5661,N_7983);
or U11703 (N_11703,N_6824,N_5912);
nor U11704 (N_11704,N_6550,N_6517);
nor U11705 (N_11705,N_6415,N_6859);
and U11706 (N_11706,N_5834,N_5391);
or U11707 (N_11707,N_6562,N_6120);
and U11708 (N_11708,N_5152,N_4068);
or U11709 (N_11709,N_7189,N_5576);
and U11710 (N_11710,N_7912,N_7050);
or U11711 (N_11711,N_5773,N_4866);
or U11712 (N_11712,N_5528,N_4199);
or U11713 (N_11713,N_6112,N_4250);
or U11714 (N_11714,N_6568,N_4885);
nand U11715 (N_11715,N_4372,N_4278);
nand U11716 (N_11716,N_4001,N_6997);
nor U11717 (N_11717,N_4014,N_5690);
or U11718 (N_11718,N_5409,N_5020);
nor U11719 (N_11719,N_6944,N_5907);
or U11720 (N_11720,N_6686,N_7844);
xor U11721 (N_11721,N_7376,N_5402);
nand U11722 (N_11722,N_5575,N_4411);
nand U11723 (N_11723,N_6927,N_5743);
nor U11724 (N_11724,N_7393,N_4332);
nand U11725 (N_11725,N_7968,N_7426);
xnor U11726 (N_11726,N_5221,N_5728);
nand U11727 (N_11727,N_5396,N_7584);
or U11728 (N_11728,N_4497,N_4026);
nor U11729 (N_11729,N_7030,N_5537);
nand U11730 (N_11730,N_6764,N_4235);
nand U11731 (N_11731,N_7677,N_5179);
nand U11732 (N_11732,N_4846,N_4484);
or U11733 (N_11733,N_5384,N_6736);
and U11734 (N_11734,N_4986,N_5540);
or U11735 (N_11735,N_4866,N_6802);
nand U11736 (N_11736,N_5544,N_4332);
or U11737 (N_11737,N_7353,N_5034);
nor U11738 (N_11738,N_5211,N_4992);
nand U11739 (N_11739,N_5405,N_7052);
and U11740 (N_11740,N_5691,N_5097);
or U11741 (N_11741,N_7084,N_4062);
or U11742 (N_11742,N_4340,N_6583);
nand U11743 (N_11743,N_7854,N_6310);
and U11744 (N_11744,N_6940,N_7101);
nand U11745 (N_11745,N_5329,N_6587);
and U11746 (N_11746,N_7776,N_6217);
and U11747 (N_11747,N_5388,N_7670);
nor U11748 (N_11748,N_5024,N_5471);
or U11749 (N_11749,N_4978,N_5780);
or U11750 (N_11750,N_7803,N_5288);
or U11751 (N_11751,N_7843,N_6665);
nor U11752 (N_11752,N_4706,N_4409);
nand U11753 (N_11753,N_5398,N_5716);
and U11754 (N_11754,N_6688,N_5348);
xnor U11755 (N_11755,N_7627,N_4606);
and U11756 (N_11756,N_7699,N_4661);
or U11757 (N_11757,N_5271,N_5073);
nand U11758 (N_11758,N_5250,N_7762);
xnor U11759 (N_11759,N_6857,N_4000);
nand U11760 (N_11760,N_7147,N_4591);
nand U11761 (N_11761,N_6775,N_7310);
and U11762 (N_11762,N_7438,N_4152);
xor U11763 (N_11763,N_7518,N_4219);
or U11764 (N_11764,N_4545,N_5255);
or U11765 (N_11765,N_5256,N_7987);
nand U11766 (N_11766,N_5646,N_7134);
and U11767 (N_11767,N_6358,N_7577);
nand U11768 (N_11768,N_5686,N_5363);
nand U11769 (N_11769,N_7670,N_4366);
nor U11770 (N_11770,N_7882,N_4002);
nand U11771 (N_11771,N_6672,N_4905);
and U11772 (N_11772,N_5429,N_4875);
nor U11773 (N_11773,N_7551,N_5603);
and U11774 (N_11774,N_4121,N_6194);
or U11775 (N_11775,N_6767,N_6067);
nand U11776 (N_11776,N_7999,N_7251);
nand U11777 (N_11777,N_6479,N_5745);
or U11778 (N_11778,N_6255,N_5321);
nand U11779 (N_11779,N_5418,N_4901);
nand U11780 (N_11780,N_6345,N_6434);
nand U11781 (N_11781,N_6405,N_6106);
or U11782 (N_11782,N_6711,N_7256);
or U11783 (N_11783,N_7521,N_7771);
or U11784 (N_11784,N_6941,N_6061);
nor U11785 (N_11785,N_5503,N_4866);
nor U11786 (N_11786,N_4561,N_4854);
or U11787 (N_11787,N_6071,N_5131);
or U11788 (N_11788,N_7570,N_6946);
xnor U11789 (N_11789,N_5869,N_6229);
nand U11790 (N_11790,N_4604,N_6499);
or U11791 (N_11791,N_6777,N_7603);
nand U11792 (N_11792,N_4468,N_7359);
or U11793 (N_11793,N_4954,N_7963);
nand U11794 (N_11794,N_4935,N_4270);
nor U11795 (N_11795,N_6020,N_5697);
nand U11796 (N_11796,N_5201,N_7646);
nor U11797 (N_11797,N_7330,N_4683);
or U11798 (N_11798,N_4187,N_4337);
nor U11799 (N_11799,N_6164,N_6647);
or U11800 (N_11800,N_4200,N_7366);
and U11801 (N_11801,N_6139,N_7649);
or U11802 (N_11802,N_6511,N_5311);
nor U11803 (N_11803,N_4488,N_6730);
nor U11804 (N_11804,N_6680,N_6216);
nor U11805 (N_11805,N_7280,N_7856);
and U11806 (N_11806,N_6931,N_5613);
or U11807 (N_11807,N_7237,N_4776);
nor U11808 (N_11808,N_4106,N_6915);
nand U11809 (N_11809,N_4652,N_5436);
or U11810 (N_11810,N_6798,N_6697);
or U11811 (N_11811,N_7370,N_4896);
and U11812 (N_11812,N_6650,N_4824);
or U11813 (N_11813,N_4746,N_6524);
nor U11814 (N_11814,N_4983,N_5941);
nand U11815 (N_11815,N_7380,N_5046);
and U11816 (N_11816,N_5791,N_5227);
or U11817 (N_11817,N_7195,N_7412);
nor U11818 (N_11818,N_5017,N_5319);
or U11819 (N_11819,N_7263,N_7176);
nor U11820 (N_11820,N_6180,N_7166);
nand U11821 (N_11821,N_4464,N_7013);
or U11822 (N_11822,N_6075,N_5195);
or U11823 (N_11823,N_7571,N_7851);
and U11824 (N_11824,N_7024,N_4221);
nor U11825 (N_11825,N_7993,N_7567);
nand U11826 (N_11826,N_4333,N_6601);
nor U11827 (N_11827,N_4607,N_6157);
nor U11828 (N_11828,N_4723,N_5838);
xnor U11829 (N_11829,N_7810,N_7709);
and U11830 (N_11830,N_7540,N_5397);
xnor U11831 (N_11831,N_7474,N_6765);
or U11832 (N_11832,N_5266,N_7985);
xor U11833 (N_11833,N_7800,N_7650);
and U11834 (N_11834,N_4841,N_4550);
nor U11835 (N_11835,N_7435,N_4873);
nor U11836 (N_11836,N_5327,N_4332);
and U11837 (N_11837,N_6850,N_7359);
and U11838 (N_11838,N_4637,N_4246);
nand U11839 (N_11839,N_5420,N_7704);
nor U11840 (N_11840,N_6574,N_5861);
xor U11841 (N_11841,N_6091,N_4598);
and U11842 (N_11842,N_7242,N_5097);
xnor U11843 (N_11843,N_6012,N_7815);
nand U11844 (N_11844,N_7217,N_4700);
nand U11845 (N_11845,N_4365,N_5143);
and U11846 (N_11846,N_5891,N_7825);
or U11847 (N_11847,N_4653,N_6739);
nor U11848 (N_11848,N_4590,N_6236);
nor U11849 (N_11849,N_6025,N_5193);
xnor U11850 (N_11850,N_4343,N_6787);
or U11851 (N_11851,N_5817,N_6388);
nand U11852 (N_11852,N_6560,N_7681);
or U11853 (N_11853,N_6526,N_6068);
or U11854 (N_11854,N_6156,N_4775);
nand U11855 (N_11855,N_7618,N_5269);
xnor U11856 (N_11856,N_7978,N_5862);
nor U11857 (N_11857,N_7772,N_6163);
or U11858 (N_11858,N_6118,N_5613);
nor U11859 (N_11859,N_4853,N_4635);
nand U11860 (N_11860,N_5408,N_6361);
and U11861 (N_11861,N_6270,N_5993);
or U11862 (N_11862,N_6965,N_5898);
or U11863 (N_11863,N_5018,N_6752);
xnor U11864 (N_11864,N_7765,N_5737);
nor U11865 (N_11865,N_4877,N_5007);
nor U11866 (N_11866,N_5423,N_5075);
nand U11867 (N_11867,N_6259,N_4789);
nor U11868 (N_11868,N_4454,N_6440);
nand U11869 (N_11869,N_6911,N_7162);
or U11870 (N_11870,N_4232,N_4968);
nand U11871 (N_11871,N_6229,N_6891);
nor U11872 (N_11872,N_6298,N_5704);
or U11873 (N_11873,N_5024,N_4740);
and U11874 (N_11874,N_7149,N_4343);
nor U11875 (N_11875,N_7584,N_6190);
nand U11876 (N_11876,N_5833,N_6138);
nand U11877 (N_11877,N_5331,N_7639);
nand U11878 (N_11878,N_5356,N_6551);
nand U11879 (N_11879,N_6129,N_7482);
nand U11880 (N_11880,N_7003,N_7108);
and U11881 (N_11881,N_7995,N_4693);
nor U11882 (N_11882,N_6236,N_4671);
nor U11883 (N_11883,N_5197,N_4741);
nand U11884 (N_11884,N_6602,N_7475);
and U11885 (N_11885,N_7407,N_7210);
and U11886 (N_11886,N_7250,N_6594);
and U11887 (N_11887,N_6885,N_6058);
nor U11888 (N_11888,N_6715,N_5929);
or U11889 (N_11889,N_4371,N_7361);
and U11890 (N_11890,N_6207,N_4454);
and U11891 (N_11891,N_7254,N_4153);
nor U11892 (N_11892,N_6801,N_7849);
xor U11893 (N_11893,N_5264,N_5478);
and U11894 (N_11894,N_7352,N_4247);
nor U11895 (N_11895,N_5841,N_4666);
and U11896 (N_11896,N_5128,N_6765);
and U11897 (N_11897,N_6317,N_6204);
and U11898 (N_11898,N_7424,N_6855);
and U11899 (N_11899,N_6434,N_7568);
and U11900 (N_11900,N_5747,N_5453);
or U11901 (N_11901,N_5563,N_6235);
nand U11902 (N_11902,N_7333,N_6979);
nand U11903 (N_11903,N_7763,N_4909);
or U11904 (N_11904,N_5017,N_7435);
nor U11905 (N_11905,N_7305,N_5251);
or U11906 (N_11906,N_7995,N_4461);
nor U11907 (N_11907,N_5056,N_7937);
or U11908 (N_11908,N_7872,N_5828);
nor U11909 (N_11909,N_5878,N_6047);
or U11910 (N_11910,N_6830,N_4811);
xnor U11911 (N_11911,N_5787,N_6734);
or U11912 (N_11912,N_7186,N_5187);
and U11913 (N_11913,N_5753,N_5576);
nor U11914 (N_11914,N_4651,N_5549);
and U11915 (N_11915,N_4884,N_6470);
xnor U11916 (N_11916,N_4127,N_7243);
nor U11917 (N_11917,N_6699,N_4006);
and U11918 (N_11918,N_6467,N_7730);
and U11919 (N_11919,N_5026,N_5127);
nand U11920 (N_11920,N_5552,N_5318);
nand U11921 (N_11921,N_6667,N_4449);
xor U11922 (N_11922,N_4363,N_4506);
nand U11923 (N_11923,N_7597,N_4659);
and U11924 (N_11924,N_4247,N_4773);
and U11925 (N_11925,N_4499,N_7567);
nor U11926 (N_11926,N_5299,N_5837);
and U11927 (N_11927,N_6468,N_5142);
nor U11928 (N_11928,N_5888,N_4486);
nand U11929 (N_11929,N_6927,N_4987);
and U11930 (N_11930,N_4862,N_4113);
nor U11931 (N_11931,N_4229,N_6899);
nor U11932 (N_11932,N_6070,N_6474);
and U11933 (N_11933,N_5906,N_5894);
nand U11934 (N_11934,N_5414,N_6013);
or U11935 (N_11935,N_7915,N_6834);
xor U11936 (N_11936,N_5754,N_5152);
xnor U11937 (N_11937,N_6626,N_6384);
nand U11938 (N_11938,N_4366,N_7740);
nor U11939 (N_11939,N_7909,N_5695);
nor U11940 (N_11940,N_7499,N_5306);
nand U11941 (N_11941,N_6693,N_6425);
nor U11942 (N_11942,N_4407,N_6338);
or U11943 (N_11943,N_4659,N_6061);
nor U11944 (N_11944,N_6068,N_4139);
or U11945 (N_11945,N_4433,N_4522);
and U11946 (N_11946,N_7024,N_5278);
or U11947 (N_11947,N_5609,N_7490);
or U11948 (N_11948,N_4848,N_5145);
nor U11949 (N_11949,N_6051,N_5438);
or U11950 (N_11950,N_7027,N_5559);
or U11951 (N_11951,N_7432,N_7794);
nand U11952 (N_11952,N_4274,N_5299);
and U11953 (N_11953,N_4823,N_5589);
or U11954 (N_11954,N_7255,N_5166);
and U11955 (N_11955,N_6139,N_4794);
nor U11956 (N_11956,N_7878,N_4383);
and U11957 (N_11957,N_4272,N_4586);
nand U11958 (N_11958,N_4867,N_4254);
or U11959 (N_11959,N_5948,N_6245);
nor U11960 (N_11960,N_4796,N_5012);
nand U11961 (N_11961,N_4912,N_6507);
xnor U11962 (N_11962,N_6932,N_4210);
xnor U11963 (N_11963,N_4850,N_6012);
nand U11964 (N_11964,N_4334,N_7446);
nor U11965 (N_11965,N_6392,N_5731);
nor U11966 (N_11966,N_7369,N_6012);
nand U11967 (N_11967,N_7056,N_5567);
nor U11968 (N_11968,N_4925,N_4888);
nor U11969 (N_11969,N_6028,N_4280);
xnor U11970 (N_11970,N_6762,N_5843);
nor U11971 (N_11971,N_6714,N_6293);
nor U11972 (N_11972,N_4185,N_6968);
nor U11973 (N_11973,N_6117,N_4172);
or U11974 (N_11974,N_4681,N_5948);
or U11975 (N_11975,N_7973,N_7353);
nor U11976 (N_11976,N_4944,N_4562);
nor U11977 (N_11977,N_4965,N_4843);
nor U11978 (N_11978,N_7997,N_4333);
nand U11979 (N_11979,N_7290,N_6262);
nor U11980 (N_11980,N_5036,N_6798);
nor U11981 (N_11981,N_6473,N_7294);
or U11982 (N_11982,N_7736,N_6813);
nor U11983 (N_11983,N_6163,N_5770);
nor U11984 (N_11984,N_7020,N_7705);
or U11985 (N_11985,N_6197,N_4053);
xor U11986 (N_11986,N_5508,N_5024);
nand U11987 (N_11987,N_4549,N_7772);
or U11988 (N_11988,N_7513,N_6675);
and U11989 (N_11989,N_5817,N_7603);
or U11990 (N_11990,N_6517,N_5554);
xnor U11991 (N_11991,N_5711,N_4325);
nor U11992 (N_11992,N_5339,N_5774);
and U11993 (N_11993,N_7906,N_4612);
nor U11994 (N_11994,N_6293,N_6042);
nor U11995 (N_11995,N_5099,N_5226);
nor U11996 (N_11996,N_7419,N_7050);
or U11997 (N_11997,N_7667,N_4711);
nor U11998 (N_11998,N_6074,N_4519);
and U11999 (N_11999,N_6096,N_4210);
nand U12000 (N_12000,N_10752,N_9640);
nand U12001 (N_12001,N_9387,N_9773);
or U12002 (N_12002,N_10683,N_11419);
nand U12003 (N_12003,N_8431,N_9541);
xnor U12004 (N_12004,N_8244,N_11086);
nand U12005 (N_12005,N_9627,N_10237);
or U12006 (N_12006,N_8580,N_9732);
nand U12007 (N_12007,N_8281,N_10125);
xnor U12008 (N_12008,N_8837,N_11626);
and U12009 (N_12009,N_10588,N_10368);
xor U12010 (N_12010,N_8475,N_11065);
nand U12011 (N_12011,N_10478,N_9235);
or U12012 (N_12012,N_9139,N_11237);
nand U12013 (N_12013,N_10000,N_10124);
or U12014 (N_12014,N_11830,N_8752);
or U12015 (N_12015,N_10476,N_10099);
and U12016 (N_12016,N_10185,N_9319);
and U12017 (N_12017,N_10038,N_8730);
xnor U12018 (N_12018,N_10204,N_11159);
nand U12019 (N_12019,N_8455,N_11598);
and U12020 (N_12020,N_9934,N_11232);
and U12021 (N_12021,N_8635,N_8458);
nand U12022 (N_12022,N_10266,N_11037);
nand U12023 (N_12023,N_8710,N_9098);
and U12024 (N_12024,N_9320,N_10540);
nand U12025 (N_12025,N_8848,N_9920);
xor U12026 (N_12026,N_10777,N_9129);
and U12027 (N_12027,N_10570,N_10695);
nor U12028 (N_12028,N_9563,N_11718);
nand U12029 (N_12029,N_10286,N_11593);
nor U12030 (N_12030,N_11643,N_8792);
or U12031 (N_12031,N_11653,N_8563);
and U12032 (N_12032,N_10801,N_11901);
xor U12033 (N_12033,N_9717,N_8107);
and U12034 (N_12034,N_8644,N_10451);
xor U12035 (N_12035,N_10456,N_9980);
and U12036 (N_12036,N_10883,N_9799);
or U12037 (N_12037,N_9629,N_11807);
nor U12038 (N_12038,N_9205,N_10437);
nor U12039 (N_12039,N_10200,N_11640);
or U12040 (N_12040,N_8985,N_11912);
nor U12041 (N_12041,N_9008,N_9577);
nand U12042 (N_12042,N_8062,N_10575);
nand U12043 (N_12043,N_9957,N_10130);
nor U12044 (N_12044,N_11535,N_10968);
nand U12045 (N_12045,N_9306,N_11781);
nand U12046 (N_12046,N_10958,N_10094);
or U12047 (N_12047,N_10720,N_8116);
or U12048 (N_12048,N_8591,N_11141);
or U12049 (N_12049,N_8777,N_11767);
or U12050 (N_12050,N_10264,N_9156);
nand U12051 (N_12051,N_10747,N_10372);
and U12052 (N_12052,N_11569,N_10195);
or U12053 (N_12053,N_9927,N_8690);
xor U12054 (N_12054,N_8226,N_11456);
nor U12055 (N_12055,N_11424,N_11841);
or U12056 (N_12056,N_10894,N_8781);
nand U12057 (N_12057,N_9995,N_10671);
or U12058 (N_12058,N_9258,N_9068);
nand U12059 (N_12059,N_8542,N_9051);
nor U12060 (N_12060,N_11461,N_10736);
nor U12061 (N_12061,N_10392,N_11246);
or U12062 (N_12062,N_8725,N_10091);
nor U12063 (N_12063,N_8682,N_8467);
or U12064 (N_12064,N_10089,N_11746);
nand U12065 (N_12065,N_9789,N_11394);
nor U12066 (N_12066,N_9349,N_11112);
nand U12067 (N_12067,N_8368,N_9095);
or U12068 (N_12068,N_10233,N_11624);
nand U12069 (N_12069,N_10098,N_9428);
and U12070 (N_12070,N_10627,N_8469);
nor U12071 (N_12071,N_8233,N_9027);
nand U12072 (N_12072,N_8262,N_9551);
xnor U12073 (N_12073,N_11639,N_9815);
xor U12074 (N_12074,N_11976,N_9979);
nand U12075 (N_12075,N_11450,N_9619);
xnor U12076 (N_12076,N_9612,N_10730);
nand U12077 (N_12077,N_11557,N_10250);
or U12078 (N_12078,N_9291,N_9321);
nor U12079 (N_12079,N_11114,N_9723);
xnor U12080 (N_12080,N_10406,N_8780);
and U12081 (N_12081,N_10263,N_8979);
or U12082 (N_12082,N_8847,N_10737);
nor U12083 (N_12083,N_11978,N_10892);
and U12084 (N_12084,N_10203,N_9521);
nand U12085 (N_12085,N_11292,N_11966);
nor U12086 (N_12086,N_11417,N_11730);
or U12087 (N_12087,N_10510,N_8810);
or U12088 (N_12088,N_10506,N_10316);
xnor U12089 (N_12089,N_11791,N_9648);
or U12090 (N_12090,N_11370,N_11464);
or U12091 (N_12091,N_9896,N_9249);
nand U12092 (N_12092,N_9292,N_9193);
nor U12093 (N_12093,N_8053,N_9378);
and U12094 (N_12094,N_10624,N_10234);
nand U12095 (N_12095,N_9173,N_10218);
nor U12096 (N_12096,N_10839,N_11062);
and U12097 (N_12097,N_11465,N_8842);
nor U12098 (N_12098,N_11705,N_9794);
nand U12099 (N_12099,N_9881,N_9337);
and U12100 (N_12100,N_9391,N_9816);
nand U12101 (N_12101,N_10044,N_10703);
or U12102 (N_12102,N_10032,N_10379);
nand U12103 (N_12103,N_8027,N_9342);
and U12104 (N_12104,N_9631,N_9854);
nand U12105 (N_12105,N_8779,N_8066);
nor U12106 (N_12106,N_9454,N_9088);
nor U12107 (N_12107,N_11646,N_9308);
or U12108 (N_12108,N_8172,N_10533);
and U12109 (N_12109,N_10600,N_10981);
nand U12110 (N_12110,N_11356,N_11310);
or U12111 (N_12111,N_11704,N_8503);
and U12112 (N_12112,N_8277,N_10536);
and U12113 (N_12113,N_8917,N_10093);
and U12114 (N_12114,N_9346,N_9059);
xor U12115 (N_12115,N_10542,N_8023);
nor U12116 (N_12116,N_11388,N_8140);
nand U12117 (N_12117,N_9586,N_11234);
and U12118 (N_12118,N_9519,N_9138);
and U12119 (N_12119,N_10776,N_11027);
nand U12120 (N_12120,N_11793,N_9668);
or U12121 (N_12121,N_11230,N_9607);
and U12122 (N_12122,N_8742,N_9626);
and U12123 (N_12123,N_11466,N_8190);
and U12124 (N_12124,N_10483,N_10873);
and U12125 (N_12125,N_8894,N_10256);
nand U12126 (N_12126,N_11383,N_11127);
nor U12127 (N_12127,N_11601,N_9818);
or U12128 (N_12128,N_11253,N_10722);
nor U12129 (N_12129,N_9774,N_8605);
and U12130 (N_12130,N_11856,N_9116);
and U12131 (N_12131,N_11533,N_9322);
nand U12132 (N_12132,N_10914,N_8218);
xor U12133 (N_12133,N_8174,N_10210);
and U12134 (N_12134,N_8912,N_10447);
xnor U12135 (N_12135,N_11085,N_8869);
nand U12136 (N_12136,N_8035,N_8575);
nand U12137 (N_12137,N_9667,N_8106);
nand U12138 (N_12138,N_8112,N_9264);
nand U12139 (N_12139,N_11615,N_11642);
nand U12140 (N_12140,N_9123,N_8138);
and U12141 (N_12141,N_10459,N_9561);
or U12142 (N_12142,N_11932,N_9753);
and U12143 (N_12143,N_10698,N_9420);
nor U12144 (N_12144,N_8483,N_8685);
nand U12145 (N_12145,N_9000,N_11679);
nor U12146 (N_12146,N_10658,N_10283);
and U12147 (N_12147,N_11252,N_10319);
nor U12148 (N_12148,N_9108,N_9417);
nor U12149 (N_12149,N_9950,N_10423);
or U12150 (N_12150,N_11373,N_9520);
xor U12151 (N_12151,N_10708,N_9733);
or U12152 (N_12152,N_8599,N_11335);
or U12153 (N_12153,N_10844,N_9903);
and U12154 (N_12154,N_8430,N_8378);
nor U12155 (N_12155,N_11962,N_10933);
nand U12156 (N_12156,N_8724,N_11291);
nand U12157 (N_12157,N_10076,N_10582);
xor U12158 (N_12158,N_9537,N_10211);
and U12159 (N_12159,N_9189,N_11503);
nor U12160 (N_12160,N_10718,N_8992);
nor U12161 (N_12161,N_10384,N_9099);
xor U12162 (N_12162,N_8427,N_9140);
nor U12163 (N_12163,N_11838,N_10896);
and U12164 (N_12164,N_8625,N_11104);
nand U12165 (N_12165,N_9429,N_11866);
nor U12166 (N_12166,N_11371,N_11621);
and U12167 (N_12167,N_10449,N_10854);
and U12168 (N_12168,N_11697,N_9048);
and U12169 (N_12169,N_8373,N_9097);
or U12170 (N_12170,N_9623,N_8868);
and U12171 (N_12171,N_11648,N_10630);
or U12172 (N_12172,N_9225,N_8829);
and U12173 (N_12173,N_11053,N_10388);
or U12174 (N_12174,N_11025,N_8069);
or U12175 (N_12175,N_8183,N_9826);
or U12176 (N_12176,N_11622,N_9295);
and U12177 (N_12177,N_11000,N_8684);
nand U12178 (N_12178,N_9355,N_9608);
xnor U12179 (N_12179,N_8026,N_9535);
or U12180 (N_12180,N_8885,N_10407);
nor U12181 (N_12181,N_11735,N_9599);
nand U12182 (N_12182,N_8288,N_8549);
nand U12183 (N_12183,N_9849,N_10174);
and U12184 (N_12184,N_8996,N_9237);
xor U12185 (N_12185,N_8231,N_9560);
nand U12186 (N_12186,N_9567,N_9795);
xnor U12187 (N_12187,N_10434,N_10011);
nor U12188 (N_12188,N_11307,N_8594);
nor U12189 (N_12189,N_11880,N_10706);
nor U12190 (N_12190,N_11766,N_8672);
or U12191 (N_12191,N_8778,N_10635);
and U12192 (N_12192,N_11493,N_9688);
or U12193 (N_12193,N_10490,N_8411);
and U12194 (N_12194,N_8477,N_9268);
or U12195 (N_12195,N_11109,N_9504);
nand U12196 (N_12196,N_11606,N_8002);
and U12197 (N_12197,N_9426,N_8993);
nor U12198 (N_12198,N_8068,N_8816);
and U12199 (N_12199,N_10908,N_10984);
or U12200 (N_12200,N_9054,N_10673);
nand U12201 (N_12201,N_9506,N_9461);
nor U12202 (N_12202,N_10727,N_9202);
nor U12203 (N_12203,N_11119,N_9239);
xor U12204 (N_12204,N_9945,N_11729);
or U12205 (N_12205,N_10340,N_9061);
nor U12206 (N_12206,N_10520,N_10620);
xnor U12207 (N_12207,N_10564,N_10178);
and U12208 (N_12208,N_10811,N_10429);
and U12209 (N_12209,N_9164,N_8474);
xnor U12210 (N_12210,N_9827,N_9588);
or U12211 (N_12211,N_9634,N_9356);
and U12212 (N_12212,N_9968,N_11055);
nand U12213 (N_12213,N_11251,N_10357);
nand U12214 (N_12214,N_10999,N_8279);
and U12215 (N_12215,N_8963,N_8852);
xor U12216 (N_12216,N_10663,N_10106);
or U12217 (N_12217,N_10045,N_11130);
or U12218 (N_12218,N_8711,N_11713);
nor U12219 (N_12219,N_10834,N_10608);
nor U12220 (N_12220,N_9282,N_10660);
or U12221 (N_12221,N_11478,N_11519);
xor U12222 (N_12222,N_10833,N_10962);
or U12223 (N_12223,N_9141,N_10581);
or U12224 (N_12224,N_10553,N_10767);
nor U12225 (N_12225,N_10640,N_9999);
xor U12226 (N_12226,N_10383,N_10487);
nor U12227 (N_12227,N_9833,N_10590);
or U12228 (N_12228,N_11675,N_9214);
or U12229 (N_12229,N_8751,N_9340);
or U12230 (N_12230,N_8924,N_9365);
nand U12231 (N_12231,N_8299,N_10924);
xor U12232 (N_12232,N_11341,N_11980);
nand U12233 (N_12233,N_8929,N_11798);
nor U12234 (N_12234,N_8891,N_10002);
nor U12235 (N_12235,N_8903,N_10554);
xor U12236 (N_12236,N_9070,N_8433);
nand U12237 (N_12237,N_8389,N_11459);
nor U12238 (N_12238,N_9079,N_9037);
nand U12239 (N_12239,N_11574,N_9817);
nand U12240 (N_12240,N_9593,N_11512);
nand U12241 (N_12241,N_10010,N_8346);
or U12242 (N_12242,N_11967,N_9332);
or U12243 (N_12243,N_9357,N_8569);
and U12244 (N_12244,N_10444,N_11579);
nand U12245 (N_12245,N_8001,N_8223);
nand U12246 (N_12246,N_10146,N_9559);
nand U12247 (N_12247,N_10589,N_10289);
and U12248 (N_12248,N_9451,N_11451);
xnor U12249 (N_12249,N_8480,N_11403);
xnor U12250 (N_12250,N_8079,N_8444);
or U12251 (N_12251,N_8214,N_9911);
nor U12252 (N_12252,N_10438,N_8128);
and U12253 (N_12253,N_10988,N_8524);
and U12254 (N_12254,N_8339,N_11182);
or U12255 (N_12255,N_11347,N_11360);
and U12256 (N_12256,N_8384,N_9065);
nor U12257 (N_12257,N_9408,N_11080);
nand U12258 (N_12258,N_9720,N_9962);
xnor U12259 (N_12259,N_8385,N_9836);
nor U12260 (N_12260,N_11337,N_10657);
xor U12261 (N_12261,N_11379,N_11799);
or U12262 (N_12262,N_10493,N_11655);
and U12263 (N_12263,N_8876,N_11514);
nand U12264 (N_12264,N_10293,N_9403);
xor U12265 (N_12265,N_8399,N_8228);
nand U12266 (N_12266,N_11985,N_10659);
nand U12267 (N_12267,N_11524,N_11368);
nor U12268 (N_12268,N_11874,N_11496);
nor U12269 (N_12269,N_11212,N_8061);
nand U12270 (N_12270,N_10973,N_11391);
nor U12271 (N_12271,N_11092,N_10682);
or U12272 (N_12272,N_10466,N_8489);
nor U12273 (N_12273,N_11765,N_8950);
xor U12274 (N_12274,N_8877,N_8000);
and U12275 (N_12275,N_9958,N_11158);
and U12276 (N_12276,N_9587,N_10820);
nor U12277 (N_12277,N_9310,N_9296);
or U12278 (N_12278,N_8611,N_11777);
xor U12279 (N_12279,N_10742,N_8381);
nand U12280 (N_12280,N_11521,N_9829);
and U12281 (N_12281,N_9807,N_8292);
xor U12282 (N_12282,N_11894,N_10842);
nand U12283 (N_12283,N_9693,N_8939);
and U12284 (N_12284,N_9499,N_8956);
xor U12285 (N_12285,N_10381,N_9662);
or U12286 (N_12286,N_8793,N_9677);
nand U12287 (N_12287,N_8920,N_9146);
nand U12288 (N_12288,N_10016,N_11229);
nand U12289 (N_12289,N_11007,N_8731);
or U12290 (N_12290,N_9183,N_10157);
xor U12291 (N_12291,N_10020,N_10546);
and U12292 (N_12292,N_9137,N_11952);
nand U12293 (N_12293,N_10005,N_10893);
nand U12294 (N_12294,N_9477,N_11869);
or U12295 (N_12295,N_11612,N_8864);
nor U12296 (N_12296,N_11986,N_10315);
nand U12297 (N_12297,N_8666,N_9240);
nor U12298 (N_12298,N_10403,N_9476);
and U12299 (N_12299,N_9393,N_11162);
nand U12300 (N_12300,N_10351,N_8916);
nand U12301 (N_12301,N_8817,N_10312);
nand U12302 (N_12302,N_11336,N_9121);
or U12303 (N_12303,N_11448,N_8067);
and U12304 (N_12304,N_9769,N_11430);
nor U12305 (N_12305,N_8688,N_11170);
or U12306 (N_12306,N_9280,N_8139);
nand U12307 (N_12307,N_8042,N_11800);
nand U12308 (N_12308,N_8372,N_11329);
nor U12309 (N_12309,N_8045,N_8986);
nor U12310 (N_12310,N_10966,N_8219);
and U12311 (N_12311,N_8783,N_9207);
and U12312 (N_12312,N_11604,N_11994);
nand U12313 (N_12313,N_10069,N_10543);
nor U12314 (N_12314,N_9916,N_11222);
xor U12315 (N_12315,N_8153,N_10639);
nand U12316 (N_12316,N_9557,N_11725);
or U12317 (N_12317,N_8994,N_11823);
nand U12318 (N_12318,N_9707,N_9734);
or U12319 (N_12319,N_8670,N_10674);
or U12320 (N_12320,N_10514,N_8377);
and U12321 (N_12321,N_10051,N_9921);
or U12322 (N_12322,N_11256,N_10859);
nor U12323 (N_12323,N_10775,N_11836);
nand U12324 (N_12324,N_9431,N_8391);
xnor U12325 (N_12325,N_10342,N_11124);
nor U12326 (N_12326,N_10052,N_9542);
and U12327 (N_12327,N_11500,N_10969);
and U12328 (N_12328,N_8721,N_8613);
nor U12329 (N_12329,N_11721,N_8495);
and U12330 (N_12330,N_10860,N_10486);
nand U12331 (N_12331,N_9242,N_11010);
nor U12332 (N_12332,N_9380,N_9007);
or U12333 (N_12333,N_11803,N_8785);
or U12334 (N_12334,N_8487,N_11043);
nand U12335 (N_12335,N_8154,N_10279);
and U12336 (N_12336,N_10992,N_8418);
or U12337 (N_12337,N_10864,N_11516);
or U12338 (N_12338,N_8784,N_10667);
and U12339 (N_12339,N_10039,N_10135);
nor U12340 (N_12340,N_11077,N_10549);
xnor U12341 (N_12341,N_11400,N_10762);
and U12342 (N_12342,N_10184,N_9107);
or U12343 (N_12343,N_10602,N_10205);
and U12344 (N_12344,N_8705,N_11619);
xor U12345 (N_12345,N_8831,N_9887);
nand U12346 (N_12346,N_11892,N_11283);
or U12347 (N_12347,N_9248,N_9851);
and U12348 (N_12348,N_10503,N_11281);
and U12349 (N_12349,N_11833,N_9166);
nand U12350 (N_12350,N_10081,N_8421);
and U12351 (N_12351,N_9569,N_11021);
nor U12352 (N_12352,N_10920,N_10793);
and U12353 (N_12353,N_9238,N_11979);
nor U12354 (N_12354,N_10729,N_11174);
and U12355 (N_12355,N_11431,N_11607);
or U12356 (N_12356,N_10910,N_9768);
xor U12357 (N_12357,N_10199,N_11304);
and U12358 (N_12358,N_11804,N_8738);
and U12359 (N_12359,N_11399,N_9370);
nand U12360 (N_12360,N_11198,N_9969);
nand U12361 (N_12361,N_11770,N_11790);
nor U12362 (N_12362,N_9122,N_9160);
or U12363 (N_12363,N_9632,N_10194);
or U12364 (N_12364,N_11469,N_10348);
nand U12365 (N_12365,N_8247,N_8732);
nor U12366 (N_12366,N_11227,N_10937);
or U12367 (N_12367,N_11282,N_10037);
nand U12368 (N_12368,N_9771,N_11947);
and U12369 (N_12369,N_9498,N_9191);
nor U12370 (N_12370,N_11270,N_8317);
or U12371 (N_12371,N_9201,N_8576);
nor U12372 (N_12372,N_10904,N_9034);
nand U12373 (N_12373,N_10042,N_10522);
or U12374 (N_12374,N_10367,N_10905);
nor U12375 (N_12375,N_11523,N_10055);
nand U12376 (N_12376,N_10886,N_9379);
nand U12377 (N_12377,N_11492,N_10685);
and U12378 (N_12378,N_10358,N_9917);
xor U12379 (N_12379,N_10723,N_11364);
nor U12380 (N_12380,N_8207,N_8692);
and U12381 (N_12381,N_8072,N_11595);
xor U12382 (N_12382,N_10862,N_9650);
nor U12383 (N_12383,N_10151,N_9610);
or U12384 (N_12384,N_9805,N_8006);
and U12385 (N_12385,N_9119,N_8124);
nor U12386 (N_12386,N_9185,N_9044);
nor U12387 (N_12387,N_10559,N_11690);
nand U12388 (N_12388,N_11207,N_8445);
or U12389 (N_12389,N_8163,N_11999);
and U12390 (N_12390,N_11047,N_10259);
nand U12391 (N_12391,N_9215,N_9184);
nand U12392 (N_12392,N_8225,N_8661);
nor U12393 (N_12393,N_10013,N_10725);
nor U12394 (N_12394,N_11998,N_8886);
nor U12395 (N_12395,N_11775,N_10949);
nor U12396 (N_12396,N_11069,N_8862);
or U12397 (N_12397,N_11795,N_10356);
or U12398 (N_12398,N_9605,N_11155);
xnor U12399 (N_12399,N_11949,N_8872);
and U12400 (N_12400,N_11250,N_9919);
xnor U12401 (N_12401,N_11989,N_8913);
or U12402 (N_12402,N_10191,N_11299);
nor U12403 (N_12403,N_10394,N_10030);
and U12404 (N_12404,N_9446,N_11651);
or U12405 (N_12405,N_11498,N_10555);
xor U12406 (N_12406,N_11020,N_9870);
nor U12407 (N_12407,N_8047,N_8806);
nand U12408 (N_12408,N_11847,N_9444);
nor U12409 (N_12409,N_11996,N_10127);
and U12410 (N_12410,N_8498,N_9012);
nand U12411 (N_12411,N_9689,N_11378);
nor U12412 (N_12412,N_11285,N_8313);
nand U12413 (N_12413,N_9411,N_10623);
and U12414 (N_12414,N_10524,N_11206);
nand U12415 (N_12415,N_9077,N_10552);
nand U12416 (N_12416,N_8125,N_9656);
nor U12417 (N_12417,N_8131,N_10505);
nor U12418 (N_12418,N_9368,N_8374);
and U12419 (N_12419,N_10754,N_9820);
nand U12420 (N_12420,N_8536,N_10025);
and U12421 (N_12421,N_11779,N_8960);
and U12422 (N_12422,N_10414,N_10939);
and U12423 (N_12423,N_10251,N_11477);
or U12424 (N_12424,N_9318,N_10017);
nor U12425 (N_12425,N_10782,N_10397);
nand U12426 (N_12426,N_8169,N_8961);
nor U12427 (N_12427,N_9948,N_9433);
and U12428 (N_12428,N_8865,N_10298);
and U12429 (N_12429,N_8130,N_8533);
xor U12430 (N_12430,N_11046,N_10338);
nor U12431 (N_12431,N_8323,N_11520);
nand U12432 (N_12432,N_8155,N_9133);
nor U12433 (N_12433,N_10376,N_9482);
and U12434 (N_12434,N_8320,N_8895);
and U12435 (N_12435,N_9495,N_11151);
or U12436 (N_12436,N_11916,N_11078);
nand U12437 (N_12437,N_11375,N_9302);
nor U12438 (N_12438,N_10391,N_9155);
and U12439 (N_12439,N_9947,N_11241);
or U12440 (N_12440,N_9149,N_10335);
nand U12441 (N_12441,N_10196,N_9294);
nor U12442 (N_12442,N_9327,N_10171);
and U12443 (N_12443,N_9930,N_8795);
and U12444 (N_12444,N_10529,N_11035);
xor U12445 (N_12445,N_11889,N_9289);
or U12446 (N_12446,N_9840,N_11290);
and U12447 (N_12447,N_8904,N_9544);
and U12448 (N_12448,N_9157,N_8973);
or U12449 (N_12449,N_9102,N_11497);
and U12450 (N_12450,N_9404,N_10728);
or U12451 (N_12451,N_8025,N_11121);
nor U12452 (N_12452,N_9271,N_11458);
nor U12453 (N_12453,N_9230,N_11472);
nor U12454 (N_12454,N_11580,N_8702);
and U12455 (N_12455,N_9330,N_9045);
xnor U12456 (N_12456,N_11481,N_10295);
nand U12457 (N_12457,N_10462,N_9348);
or U12458 (N_12458,N_10008,N_9430);
nor U12459 (N_12459,N_8159,N_8592);
nand U12460 (N_12460,N_9316,N_9313);
and U12461 (N_12461,N_9530,N_10960);
nand U12462 (N_12462,N_8941,N_10726);
or U12463 (N_12463,N_8350,N_10410);
nand U12464 (N_12464,N_10079,N_9491);
and U12465 (N_12465,N_8091,N_11991);
xor U12466 (N_12466,N_10912,N_9719);
nor U12467 (N_12467,N_8241,N_10852);
nand U12468 (N_12468,N_11553,N_11848);
or U12469 (N_12469,N_8254,N_9243);
or U12470 (N_12470,N_9011,N_9669);
or U12471 (N_12471,N_10700,N_8028);
and U12472 (N_12472,N_9017,N_9860);
nor U12473 (N_12473,N_10360,N_10713);
or U12474 (N_12474,N_9664,N_8925);
nor U12475 (N_12475,N_9407,N_8735);
or U12476 (N_12476,N_10225,N_10018);
nor U12477 (N_12477,N_9203,N_11969);
or U12478 (N_12478,N_10927,N_8796);
nand U12479 (N_12479,N_11029,N_9522);
and U12480 (N_12480,N_9010,N_8623);
and U12481 (N_12481,N_9712,N_11395);
nand U12482 (N_12482,N_10669,N_8016);
nor U12483 (N_12483,N_10764,N_9582);
nand U12484 (N_12484,N_10027,N_11576);
xnor U12485 (N_12485,N_10741,N_8302);
or U12486 (N_12486,N_10783,N_10572);
or U12487 (N_12487,N_10666,N_11594);
nand U12488 (N_12488,N_10967,N_11657);
nand U12489 (N_12489,N_11540,N_8543);
and U12490 (N_12490,N_10080,N_11636);
nand U12491 (N_12491,N_10240,N_10154);
nand U12492 (N_12492,N_11181,N_9305);
nand U12493 (N_12493,N_8791,N_10442);
and U12494 (N_12494,N_9661,N_10441);
and U12495 (N_12495,N_11148,N_8539);
nand U12496 (N_12496,N_10566,N_11832);
xnor U12497 (N_12497,N_11720,N_9726);
xnor U12498 (N_12498,N_9862,N_9671);
xnor U12499 (N_12499,N_8659,N_11177);
xor U12500 (N_12500,N_8734,N_9351);
and U12501 (N_12501,N_11968,N_9786);
nand U12502 (N_12502,N_9596,N_10048);
nor U12503 (N_12503,N_9063,N_10799);
xnor U12504 (N_12504,N_8641,N_8935);
or U12505 (N_12505,N_9480,N_9939);
and U12506 (N_12506,N_9991,N_11363);
and U12507 (N_12507,N_9219,N_9955);
nor U12508 (N_12508,N_10686,N_9244);
or U12509 (N_12509,N_8609,N_11686);
and U12510 (N_12510,N_11526,N_10735);
nor U12511 (N_12511,N_10647,N_8843);
xnor U12512 (N_12512,N_10761,N_10343);
or U12513 (N_12513,N_11278,N_8127);
and U12514 (N_12514,N_10788,N_9449);
and U12515 (N_12515,N_8311,N_11739);
nand U12516 (N_12516,N_11990,N_9206);
or U12517 (N_12517,N_8099,N_9811);
nand U12518 (N_12518,N_8270,N_11167);
nor U12519 (N_12519,N_9039,N_9485);
and U12520 (N_12520,N_11573,N_10574);
nor U12521 (N_12521,N_9513,N_8621);
nand U12522 (N_12522,N_9724,N_11249);
or U12523 (N_12523,N_11871,N_11042);
and U12524 (N_12524,N_9301,N_10498);
or U12525 (N_12525,N_10477,N_8434);
or U12526 (N_12526,N_10113,N_8517);
nor U12527 (N_12527,N_9566,N_8420);
and U12528 (N_12528,N_8040,N_9467);
nor U12529 (N_12529,N_9819,N_11462);
nor U12530 (N_12530,N_9960,N_11864);
nand U12531 (N_12531,N_9679,N_8541);
or U12532 (N_12532,N_8931,N_9038);
and U12533 (N_12533,N_8665,N_9128);
or U12534 (N_12534,N_8998,N_10954);
nor U12535 (N_12535,N_11974,N_8454);
nor U12536 (N_12536,N_8607,N_10134);
nand U12537 (N_12537,N_8020,N_8646);
nand U12538 (N_12538,N_10347,N_11122);
nor U12539 (N_12539,N_8014,N_11937);
nor U12540 (N_12540,N_8030,N_10915);
xor U12541 (N_12541,N_10314,N_8769);
nor U12542 (N_12542,N_10463,N_10758);
nand U12543 (N_12543,N_11584,N_9580);
xnor U12544 (N_12544,N_9680,N_10616);
nand U12545 (N_12545,N_8376,N_10492);
and U12546 (N_12546,N_10796,N_8460);
nor U12547 (N_12547,N_9423,N_9260);
or U12548 (N_12548,N_10304,N_11175);
nor U12549 (N_12549,N_8686,N_11457);
and U12550 (N_12550,N_8388,N_8287);
or U12551 (N_12551,N_11327,N_8953);
or U12552 (N_12552,N_8152,N_8149);
nor U12553 (N_12553,N_11171,N_8194);
and U12554 (N_12554,N_10861,N_8120);
nand U12555 (N_12555,N_11263,N_11247);
or U12556 (N_12556,N_8122,N_11529);
nand U12557 (N_12557,N_10231,N_10690);
and U12558 (N_12558,N_9001,N_9456);
xor U12559 (N_12559,N_11742,N_11614);
or U12560 (N_12560,N_8959,N_11076);
nand U12561 (N_12561,N_11782,N_10148);
and U12562 (N_12562,N_11658,N_10637);
or U12563 (N_12563,N_11072,N_11353);
or U12564 (N_12564,N_8798,N_9255);
or U12565 (N_12565,N_8584,N_8451);
and U12566 (N_12566,N_8259,N_10095);
and U12567 (N_12567,N_11928,N_9067);
and U12568 (N_12568,N_8039,N_11096);
nand U12569 (N_12569,N_9441,N_8371);
nor U12570 (N_12570,N_10070,N_10997);
nor U12571 (N_12571,N_8619,N_11248);
or U12572 (N_12572,N_10857,N_8273);
or U12573 (N_12573,N_8823,N_9787);
nor U12574 (N_12574,N_10409,N_11216);
xor U12575 (N_12575,N_10800,N_11189);
nor U12576 (N_12576,N_8095,N_9762);
nand U12577 (N_12577,N_11097,N_9159);
or U12578 (N_12578,N_10596,N_9145);
or U12579 (N_12579,N_9642,N_10323);
nor U12580 (N_12580,N_11139,N_8165);
nand U12581 (N_12581,N_8522,N_10161);
nand U12582 (N_12582,N_8182,N_9466);
nor U12583 (N_12583,N_11164,N_10961);
nand U12584 (N_12584,N_11397,N_11088);
nor U12585 (N_12585,N_9180,N_10846);
and U12586 (N_12586,N_11693,N_11199);
or U12587 (N_12587,N_8761,N_10644);
nand U12588 (N_12588,N_11757,N_10665);
xnor U12589 (N_12589,N_10712,N_10748);
nand U12590 (N_12590,N_8456,N_11144);
or U12591 (N_12591,N_11405,N_11054);
nor U12592 (N_12592,N_9841,N_9150);
and U12593 (N_12593,N_8177,N_9400);
or U12594 (N_12594,N_9965,N_10819);
or U12595 (N_12595,N_11333,N_10103);
xor U12596 (N_12596,N_9217,N_10643);
nand U12597 (N_12597,N_10525,N_11887);
nor U12598 (N_12598,N_11239,N_8056);
nand U12599 (N_12599,N_11362,N_9638);
nor U12600 (N_12600,N_9442,N_8747);
and U12601 (N_12601,N_10561,N_8867);
nor U12602 (N_12602,N_11446,N_8740);
nor U12603 (N_12603,N_11572,N_8077);
nand U12604 (N_12604,N_9142,N_11752);
nor U12605 (N_12605,N_10101,N_8975);
or U12606 (N_12606,N_11971,N_10202);
nand U12607 (N_12607,N_8509,N_11703);
or U12608 (N_12608,N_9646,N_9912);
nand U12609 (N_12609,N_10638,N_9178);
xor U12610 (N_12610,N_9785,N_8799);
xnor U12611 (N_12611,N_11664,N_8321);
or U12612 (N_12612,N_8708,N_11958);
or U12613 (N_12613,N_11599,N_11975);
nor U12614 (N_12614,N_9872,N_9548);
nand U12615 (N_12615,N_11600,N_10744);
nor U12616 (N_12616,N_9825,N_8046);
nand U12617 (N_12617,N_8361,N_9236);
and U12618 (N_12618,N_9928,N_10271);
nand U12619 (N_12619,N_10865,N_11414);
xor U12620 (N_12620,N_10517,N_8628);
nor U12621 (N_12621,N_9481,N_11138);
nor U12622 (N_12622,N_11411,N_9698);
xnor U12623 (N_12623,N_8386,N_8370);
xor U12624 (N_12624,N_8200,N_11039);
nand U12625 (N_12625,N_8111,N_10268);
nor U12626 (N_12626,N_10100,N_11835);
or U12627 (N_12627,N_9307,N_8422);
nand U12628 (N_12628,N_10497,N_8583);
or U12629 (N_12629,N_8243,N_10355);
xor U12630 (N_12630,N_8176,N_8720);
nor U12631 (N_12631,N_10511,N_8074);
and U12632 (N_12632,N_11567,N_10925);
or U12633 (N_12633,N_9975,N_11374);
nand U12634 (N_12634,N_11495,N_9761);
nor U12635 (N_12635,N_8531,N_11499);
or U12636 (N_12636,N_9625,N_8133);
or U12637 (N_12637,N_11441,N_11126);
and U12638 (N_12638,N_10064,N_9453);
and U12639 (N_12639,N_11809,N_8492);
or U12640 (N_12640,N_10119,N_11896);
nor U12641 (N_12641,N_11432,N_10244);
nor U12642 (N_12642,N_9022,N_9532);
xnor U12643 (N_12643,N_10179,N_11410);
xor U12644 (N_12644,N_10189,N_8090);
and U12645 (N_12645,N_11925,N_11691);
nor U12646 (N_12646,N_11862,N_9448);
nor U12647 (N_12647,N_9055,N_11111);
or U12648 (N_12648,N_11217,N_11760);
xnor U12649 (N_12649,N_11785,N_10214);
and U12650 (N_12650,N_8019,N_11209);
and U12651 (N_12651,N_8261,N_9286);
and U12652 (N_12652,N_8351,N_9501);
xnor U12653 (N_12653,N_9372,N_11277);
nand U12654 (N_12654,N_8699,N_8424);
and U12655 (N_12655,N_11632,N_10473);
nand U12656 (N_12656,N_10837,N_11300);
nand U12657 (N_12657,N_10353,N_9932);
xnor U12658 (N_12658,N_9756,N_10166);
and U12659 (N_12659,N_9822,N_9529);
nand U12660 (N_12660,N_10512,N_8545);
xnor U12661 (N_12661,N_10303,N_10110);
xnor U12662 (N_12662,N_10895,N_10273);
or U12663 (N_12663,N_10023,N_11647);
nand U12664 (N_12664,N_10705,N_10550);
nand U12665 (N_12665,N_9345,N_11981);
nand U12666 (N_12666,N_11873,N_10972);
nand U12667 (N_12667,N_9959,N_10900);
and U12668 (N_12668,N_9279,N_10646);
xor U12669 (N_12669,N_11620,N_11831);
nor U12670 (N_12670,N_11289,N_9565);
nand U12671 (N_12671,N_11101,N_10285);
nand U12672 (N_12672,N_9683,N_10021);
xnor U12673 (N_12673,N_11471,N_11810);
nand U12674 (N_12674,N_8827,N_9040);
and U12675 (N_12675,N_9125,N_9888);
or U12676 (N_12676,N_8830,N_9174);
and U12677 (N_12677,N_8196,N_9035);
and U12678 (N_12678,N_8278,N_9266);
nand U12679 (N_12679,N_9933,N_11628);
nor U12680 (N_12680,N_8396,N_8870);
nand U12681 (N_12681,N_8485,N_10721);
or U12682 (N_12682,N_8071,N_11191);
or U12683 (N_12683,N_10216,N_8633);
and U12684 (N_12684,N_11786,N_8240);
nand U12685 (N_12685,N_9708,N_9853);
and U12686 (N_12686,N_8008,N_9283);
nand U12687 (N_12687,N_9360,N_10082);
xnor U12688 (N_12688,N_11185,N_9194);
nand U12689 (N_12689,N_11988,N_10369);
xor U12690 (N_12690,N_9033,N_8818);
or U12691 (N_12691,N_9066,N_10711);
or U12692 (N_12692,N_9578,N_9177);
nand U12693 (N_12693,N_9171,N_10334);
nand U12694 (N_12694,N_11749,N_9584);
nor U12695 (N_12695,N_11233,N_9198);
xnor U12696 (N_12696,N_10794,N_9452);
nor U12697 (N_12697,N_10494,N_8168);
nor U12698 (N_12698,N_11930,N_9470);
nor U12699 (N_12699,N_9894,N_8770);
nand U12700 (N_12700,N_11806,N_11190);
and U12701 (N_12701,N_11812,N_9434);
or U12702 (N_12702,N_9262,N_10991);
nand U12703 (N_12703,N_10948,N_9858);
and U12704 (N_12704,N_10613,N_9437);
nand U12705 (N_12705,N_10152,N_10617);
or U12706 (N_12706,N_8652,N_10870);
nand U12707 (N_12707,N_10399,N_8728);
or U12708 (N_12708,N_9743,N_10707);
and U12709 (N_12709,N_8540,N_10963);
nand U12710 (N_12710,N_11433,N_10702);
and U12711 (N_12711,N_10569,N_8343);
nand U12712 (N_12712,N_9190,N_8119);
nand U12713 (N_12713,N_9304,N_8296);
nor U12714 (N_12714,N_8275,N_9270);
nor U12715 (N_12715,N_10330,N_10693);
nor U12716 (N_12716,N_8971,N_11107);
nand U12717 (N_12717,N_10701,N_9410);
xnor U12718 (N_12718,N_8693,N_10142);
or U12719 (N_12719,N_9914,N_9893);
and U12720 (N_12720,N_11429,N_9425);
nor U12721 (N_12721,N_9490,N_9649);
nand U12722 (N_12722,N_9830,N_10474);
nor U12723 (N_12723,N_9808,N_10491);
nor U12724 (N_12724,N_10114,N_9186);
nor U12725 (N_12725,N_8358,N_9030);
nor U12726 (N_12726,N_8972,N_9523);
or U12727 (N_12727,N_9143,N_10714);
nand U12728 (N_12728,N_9702,N_8353);
nor U12729 (N_12729,N_9151,N_8640);
or U12730 (N_12730,N_11566,N_8570);
nor U12731 (N_12731,N_10253,N_11261);
or U12732 (N_12732,N_9367,N_11452);
and U12733 (N_12733,N_11276,N_10416);
xnor U12734 (N_12734,N_8146,N_11977);
and U12735 (N_12735,N_9676,N_11902);
nand U12736 (N_12736,N_9074,N_11596);
nand U12737 (N_12737,N_9665,N_10929);
or U12738 (N_12738,N_8562,N_8824);
nand U12739 (N_12739,N_8974,N_8115);
and U12740 (N_12740,N_8589,N_10916);
and U12741 (N_12741,N_9538,N_10221);
and U12742 (N_12742,N_9531,N_11293);
nand U12743 (N_12743,N_9697,N_11473);
nand U12744 (N_12744,N_9435,N_10940);
or U12745 (N_12745,N_8076,N_11339);
or U12746 (N_12746,N_10996,N_8566);
nor U12747 (N_12747,N_8630,N_8737);
nor U12748 (N_12748,N_9211,N_9828);
xnor U12749 (N_12749,N_11681,N_9622);
nor U12750 (N_12750,N_11011,N_8809);
nor U12751 (N_12751,N_8560,N_9613);
nand U12752 (N_12752,N_11186,N_9502);
nor U12753 (N_12753,N_8683,N_11305);
and U12754 (N_12754,N_9842,N_10598);
or U12755 (N_12755,N_10294,N_11402);
nand U12756 (N_12756,N_11157,N_11100);
nor U12757 (N_12757,N_8304,N_10919);
or U12758 (N_12758,N_8404,N_8013);
and U12759 (N_12759,N_11071,N_10502);
or U12760 (N_12760,N_8631,N_11868);
or U12761 (N_12761,N_9124,N_10584);
nor U12762 (N_12762,N_9793,N_11517);
nand U12763 (N_12763,N_9892,N_10547);
nand U12764 (N_12764,N_9136,N_10242);
xor U12765 (N_12765,N_8579,N_8064);
nand U12766 (N_12766,N_10457,N_9748);
nand U12767 (N_12767,N_9091,N_8216);
and U12768 (N_12768,N_11406,N_9009);
and U12769 (N_12769,N_11683,N_10120);
nand U12770 (N_12770,N_8861,N_10802);
xnor U12771 (N_12771,N_11015,N_8849);
or U12772 (N_12772,N_10245,N_10901);
or U12773 (N_12773,N_9806,N_9273);
nand U12774 (N_12774,N_10634,N_11331);
xnor U12775 (N_12775,N_8191,N_11922);
or U12776 (N_12776,N_9483,N_11001);
or U12777 (N_12777,N_10906,N_10580);
nor U12778 (N_12778,N_8716,N_10519);
or U12779 (N_12779,N_11161,N_8400);
nand U12780 (N_12780,N_10978,N_11708);
and U12781 (N_12781,N_11002,N_10281);
or U12782 (N_12782,N_10257,N_8948);
nand U12783 (N_12783,N_9254,N_11545);
nor U12784 (N_12784,N_10654,N_9674);
nand U12785 (N_12785,N_11816,N_8426);
nor U12786 (N_12786,N_9722,N_10352);
nand U12787 (N_12787,N_9658,N_9331);
nor U12788 (N_12788,N_10255,N_8181);
and U12789 (N_12789,N_9090,N_11794);
and U12790 (N_12790,N_9639,N_10633);
and U12791 (N_12791,N_8552,N_11568);
nand U12792 (N_12792,N_11808,N_9197);
and U12793 (N_12793,N_9616,N_11324);
or U12794 (N_12794,N_8638,N_11878);
nor U12795 (N_12795,N_9314,N_8463);
nor U12796 (N_12796,N_10578,N_10432);
nand U12797 (N_12797,N_8601,N_9790);
nand U12798 (N_12798,N_9015,N_10156);
and U12799 (N_12799,N_8554,N_11137);
xor U12800 (N_12800,N_10935,N_9633);
and U12801 (N_12801,N_8417,N_11727);
nand U12802 (N_12802,N_8344,N_8516);
nand U12803 (N_12803,N_8104,N_8983);
nand U12804 (N_12804,N_8429,N_11407);
nand U12805 (N_12805,N_10931,N_9120);
nand U12806 (N_12806,N_9620,N_11041);
or U12807 (N_12807,N_11413,N_10612);
xnor U12808 (N_12808,N_11954,N_10460);
nor U12809 (N_12809,N_8018,N_11259);
nand U12810 (N_12810,N_10215,N_8844);
nor U12811 (N_12811,N_8882,N_9637);
or U12812 (N_12812,N_9210,N_8887);
nor U12813 (N_12813,N_10428,N_10740);
nand U12814 (N_12814,N_10986,N_8797);
and U12815 (N_12815,N_11425,N_10296);
nand U12816 (N_12816,N_11387,N_11294);
and U12817 (N_12817,N_9574,N_9025);
or U12818 (N_12818,N_8380,N_11480);
and U12819 (N_12819,N_8186,N_11505);
and U12820 (N_12820,N_8585,N_8551);
and U12821 (N_12821,N_11719,N_8011);
or U12822 (N_12822,N_9488,N_11822);
nand U12823 (N_12823,N_9152,N_11426);
nor U12824 (N_12824,N_11817,N_10453);
and U12825 (N_12825,N_11048,N_11771);
and U12826 (N_12826,N_10467,N_11311);
nand U12827 (N_12827,N_11287,N_10535);
nor U12828 (N_12828,N_10987,N_9175);
or U12829 (N_12829,N_11677,N_11591);
and U12830 (N_12830,N_8412,N_9213);
xnor U12831 (N_12831,N_10385,N_10789);
xnor U12832 (N_12832,N_8906,N_9187);
and U12833 (N_12833,N_10699,N_9555);
or U12834 (N_12834,N_10567,N_10848);
and U12835 (N_12835,N_8349,N_11941);
and U12836 (N_12836,N_11556,N_8274);
nand U12837 (N_12837,N_9422,N_8464);
and U12838 (N_12838,N_8326,N_8999);
nand U12839 (N_12839,N_8359,N_10274);
nor U12840 (N_12840,N_9427,N_11260);
or U12841 (N_12841,N_11936,N_11829);
nor U12842 (N_12842,N_8893,N_9343);
xnor U12843 (N_12843,N_8884,N_10359);
and U12844 (N_12844,N_10828,N_8970);
nor U12845 (N_12845,N_9901,N_9750);
nand U12846 (N_12846,N_9961,N_11706);
xnor U12847 (N_12847,N_8413,N_8896);
nor U12848 (N_12848,N_8245,N_11638);
nor U12849 (N_12849,N_9867,N_10054);
or U12850 (N_12850,N_8845,N_10446);
nor U12851 (N_12851,N_8835,N_10405);
or U12852 (N_12852,N_11169,N_10576);
xnor U12853 (N_12853,N_9371,N_11861);
nand U12854 (N_12854,N_9281,N_10258);
nand U12855 (N_12855,N_9005,N_10309);
nor U12856 (N_12856,N_9227,N_11345);
or U12857 (N_12857,N_8397,N_10733);
xnor U12858 (N_12858,N_9963,N_11898);
or U12859 (N_12859,N_10504,N_9475);
and U12860 (N_12860,N_11662,N_8851);
nand U12861 (N_12861,N_11231,N_11330);
and U12862 (N_12862,N_9381,N_8504);
nand U12863 (N_12863,N_9598,N_11343);
nor U12864 (N_12864,N_9234,N_8832);
or U12865 (N_12865,N_11712,N_9660);
and U12866 (N_12866,N_11026,N_8572);
or U12867 (N_12867,N_10565,N_9317);
nor U12868 (N_12868,N_9218,N_8494);
xor U12869 (N_12869,N_11460,N_8488);
nor U12870 (N_12870,N_10648,N_8087);
xnor U12871 (N_12871,N_10063,N_8415);
nor U12872 (N_12872,N_9096,N_10807);
nor U12873 (N_12873,N_8208,N_8537);
nor U12874 (N_12874,N_9844,N_10836);
and U12875 (N_12875,N_10950,N_8969);
nand U12876 (N_12876,N_10183,N_10326);
nand U12877 (N_12877,N_10944,N_11396);
and U12878 (N_12878,N_8523,N_8329);
and U12879 (N_12879,N_11352,N_10035);
nand U12880 (N_12880,N_10252,N_9739);
or U12881 (N_12881,N_8340,N_8298);
nor U12882 (N_12882,N_10170,N_10661);
nand U12883 (N_12883,N_8910,N_9611);
nor U12884 (N_12884,N_8902,N_9363);
nand U12885 (N_12885,N_8457,N_10689);
or U12886 (N_12886,N_9884,N_9985);
nand U12887 (N_12887,N_11006,N_8235);
and U12888 (N_12888,N_10509,N_10175);
and U12889 (N_12889,N_11711,N_10138);
xor U12890 (N_12890,N_9725,N_11188);
and U12891 (N_12891,N_8059,N_10508);
and U12892 (N_12892,N_11984,N_8697);
nand U12893 (N_12893,N_11269,N_8529);
or U12894 (N_12894,N_9412,N_9223);
nand U12895 (N_12895,N_10096,N_10167);
nor U12896 (N_12896,N_9558,N_10626);
nor U12897 (N_12897,N_9109,N_10874);
and U12898 (N_12898,N_11993,N_11117);
and U12899 (N_12899,N_8185,N_9486);
and U12900 (N_12900,N_9500,N_8102);
nand U12901 (N_12901,N_9792,N_10930);
and U12902 (N_12902,N_11682,N_8871);
and U12903 (N_12903,N_10856,N_8526);
nand U12904 (N_12904,N_8324,N_9776);
or U12905 (N_12905,N_8535,N_10022);
xor U12906 (N_12906,N_8765,N_11592);
or U12907 (N_12907,N_11858,N_10875);
and U12908 (N_12908,N_10426,N_9259);
nor U12909 (N_12909,N_11081,N_8143);
xnor U12910 (N_12910,N_11698,N_8300);
and U12911 (N_12911,N_11783,N_10817);
or U12912 (N_12912,N_10102,N_9915);
or U12913 (N_12913,N_11688,N_9373);
nand U12914 (N_12914,N_11602,N_11273);
nor U12915 (N_12915,N_8905,N_8530);
xnor U12916 (N_12916,N_8980,N_9859);
or U12917 (N_12917,N_11959,N_10795);
and U12918 (N_12918,N_9003,N_10945);
or U12919 (N_12919,N_11582,N_10619);
or U12920 (N_12920,N_11134,N_9744);
or U12921 (N_12921,N_8269,N_11625);
nor U12922 (N_12922,N_8648,N_9976);
or U12923 (N_12923,N_8577,N_11197);
xor U12924 (N_12924,N_8898,N_9713);
nor U12925 (N_12925,N_11955,N_9204);
nor U12926 (N_12926,N_9986,N_10308);
and U12927 (N_12927,N_9908,N_10207);
nor U12928 (N_12928,N_9873,N_9031);
nand U12929 (N_12929,N_9384,N_11631);
and U12930 (N_12930,N_10209,N_8671);
and U12931 (N_12931,N_9199,N_11732);
nand U12932 (N_12932,N_10607,N_9988);
or U12933 (N_12933,N_10056,N_11738);
and U12934 (N_12934,N_8875,N_11187);
or U12935 (N_12935,N_11205,N_10248);
or U12936 (N_12936,N_10162,N_10213);
and U12937 (N_12937,N_8677,N_11257);
or U12938 (N_12938,N_11860,N_9974);
or U12939 (N_12939,N_11494,N_11562);
and U12940 (N_12940,N_8878,N_9857);
and U12941 (N_12941,N_10386,N_10123);
or U12942 (N_12942,N_11764,N_8109);
nand U12943 (N_12943,N_10880,N_11412);
or U12944 (N_12944,N_10953,N_9964);
or U12945 (N_12945,N_9685,N_8364);
and U12946 (N_12946,N_8197,N_8555);
nor U12947 (N_12947,N_9315,N_8990);
and U12948 (N_12948,N_8436,N_10957);
nand U12949 (N_12949,N_11142,N_8305);
xor U12950 (N_12950,N_8315,N_11934);
nand U12951 (N_12951,N_8822,N_8309);
nand U12952 (N_12952,N_11438,N_8556);
and U12953 (N_12953,N_10557,N_8813);
and U12954 (N_12954,N_9742,N_9751);
nand U12955 (N_12955,N_9886,N_11825);
and U12956 (N_12956,N_8239,N_11877);
xor U12957 (N_12957,N_8198,N_8739);
xnor U12958 (N_12958,N_8057,N_9376);
nor U12959 (N_12959,N_8667,N_9525);
nor U12960 (N_12960,N_11774,N_10709);
xor U12961 (N_12961,N_9755,N_9791);
nor U12962 (N_12962,N_10239,N_11235);
nand U12963 (N_12963,N_11555,N_8936);
and U12964 (N_12964,N_9983,N_9624);
nor U12965 (N_12965,N_10041,N_11153);
nand U12966 (N_12966,N_11737,N_11073);
or U12967 (N_12967,N_8880,N_10219);
xnor U12968 (N_12968,N_8676,N_8134);
and U12969 (N_12969,N_8653,N_8874);
nand U12970 (N_12970,N_8407,N_11824);
nor U12971 (N_12971,N_10755,N_11578);
nor U12972 (N_12972,N_9600,N_8354);
and U12973 (N_12973,N_8227,N_11717);
nand U12974 (N_12974,N_8678,N_10813);
nand U12975 (N_12975,N_10760,N_8550);
and U12976 (N_12976,N_8478,N_10551);
nand U12977 (N_12977,N_10845,N_9468);
or U12978 (N_12978,N_8922,N_8615);
xnor U12979 (N_12979,N_11527,N_9325);
nand U12980 (N_12980,N_9850,N_8007);
nor U12981 (N_12981,N_10374,N_10579);
nand U12982 (N_12982,N_10375,N_8213);
nor U12983 (N_12983,N_11013,N_11882);
and U12984 (N_12984,N_9564,N_10075);
nand U12985 (N_12985,N_9952,N_8435);
nand U12986 (N_12986,N_10625,N_11610);
xor U12987 (N_12987,N_11763,N_9450);
nand U12988 (N_12988,N_11911,N_10872);
and U12989 (N_12989,N_9104,N_9545);
and U12990 (N_12990,N_9246,N_11268);
nand U12991 (N_12991,N_9154,N_11487);
and U12992 (N_12992,N_10400,N_11613);
nand U12993 (N_12993,N_10632,N_9505);
xor U12994 (N_12994,N_9832,N_9700);
nand U12995 (N_12995,N_11223,N_8856);
and U12996 (N_12996,N_9706,N_8933);
nand U12997 (N_12997,N_8423,N_8760);
and U12998 (N_12998,N_11361,N_9265);
and U12999 (N_12999,N_11813,N_11577);
nor U13000 (N_13000,N_11332,N_9899);
nor U13001 (N_13001,N_8468,N_11132);
nor U13002 (N_13002,N_9126,N_11255);
and U13003 (N_13003,N_9267,N_10804);
nand U13004 (N_13004,N_8081,N_11641);
nor U13005 (N_13005,N_9907,N_11597);
nor U13006 (N_13006,N_8160,N_9909);
xnor U13007 (N_13007,N_11099,N_8357);
xor U13008 (N_13008,N_8890,N_8930);
nand U13009 (N_13009,N_11534,N_8425);
and U13010 (N_13010,N_9018,N_9344);
nor U13011 (N_13011,N_9399,N_9663);
nand U13012 (N_13012,N_9871,N_11537);
and U13013 (N_13013,N_11178,N_10322);
or U13014 (N_13014,N_8005,N_8808);
and U13015 (N_13015,N_8286,N_9937);
or U13016 (N_13016,N_11609,N_10004);
and U13017 (N_13017,N_9643,N_10475);
or U13018 (N_13018,N_11245,N_11059);
xor U13019 (N_13019,N_9594,N_9796);
and U13020 (N_13020,N_11546,N_10222);
or U13021 (N_13021,N_9510,N_9383);
nand U13022 (N_13022,N_11909,N_10029);
or U13023 (N_13023,N_9162,N_8255);
nor U13024 (N_13024,N_10126,N_11891);
nand U13025 (N_13025,N_11802,N_8100);
nor U13026 (N_13026,N_10815,N_9478);
or U13027 (N_13027,N_9977,N_8775);
and U13028 (N_13028,N_11295,N_11328);
or U13029 (N_13029,N_9016,N_8419);
and U13030 (N_13030,N_8754,N_9782);
and U13031 (N_13031,N_8147,N_10262);
or U13032 (N_13032,N_8282,N_11953);
nor U13033 (N_13033,N_11468,N_10421);
nor U13034 (N_13034,N_10515,N_8821);
and U13035 (N_13035,N_8360,N_10172);
nor U13036 (N_13036,N_10746,N_10398);
nand U13037 (N_13037,N_8486,N_10046);
nand U13038 (N_13038,N_8889,N_9951);
nor U13039 (N_13039,N_9382,N_11313);
nand U13040 (N_13040,N_8568,N_9636);
nand U13041 (N_13041,N_10768,N_9705);
and U13042 (N_13042,N_11089,N_10147);
nor U13043 (N_13043,N_9721,N_10464);
and U13044 (N_13044,N_11772,N_9115);
nor U13045 (N_13045,N_10628,N_9457);
nand U13046 (N_13046,N_10371,N_10452);
xnor U13047 (N_13047,N_11886,N_11128);
nor U13048 (N_13048,N_10946,N_9880);
or U13049 (N_13049,N_9445,N_8297);
and U13050 (N_13050,N_11743,N_9402);
and U13051 (N_13051,N_9868,N_8518);
and U13052 (N_13052,N_9992,N_9944);
or U13053 (N_13053,N_11550,N_8833);
nand U13054 (N_13054,N_9539,N_10176);
xnor U13055 (N_13055,N_8501,N_8022);
nor U13056 (N_13056,N_11416,N_9278);
nor U13057 (N_13057,N_8546,N_11734);
nand U13058 (N_13058,N_11068,N_9970);
or U13059 (N_13059,N_9875,N_8318);
nor U13060 (N_13060,N_10790,N_9338);
nand U13061 (N_13061,N_10823,N_11842);
nor U13062 (N_13062,N_10670,N_11918);
and U13063 (N_13063,N_8083,N_10346);
or U13064 (N_13064,N_11511,N_8639);
and U13065 (N_13065,N_8689,N_8263);
and U13066 (N_13066,N_9573,N_11208);
nor U13067 (N_13067,N_9615,N_11927);
nand U13068 (N_13068,N_8547,N_11951);
nor U13069 (N_13069,N_10363,N_11945);
nand U13070 (N_13070,N_11837,N_9002);
or U13071 (N_13071,N_10585,N_9080);
nand U13072 (N_13072,N_9984,N_10797);
nor U13073 (N_13073,N_11365,N_8333);
nand U13074 (N_13074,N_9889,N_11890);
or U13075 (N_13075,N_11689,N_10922);
nor U13076 (N_13076,N_9856,N_9982);
nand U13077 (N_13077,N_9020,N_8319);
nor U13078 (N_13078,N_8280,N_9783);
nand U13079 (N_13079,N_8352,N_11637);
or U13080 (N_13080,N_11778,N_8506);
xor U13081 (N_13081,N_8508,N_8669);
or U13082 (N_13082,N_8749,N_8794);
or U13083 (N_13083,N_10378,N_8499);
nor U13084 (N_13084,N_9526,N_11325);
xor U13085 (N_13085,N_8180,N_9747);
xnor U13086 (N_13086,N_11544,N_8544);
nor U13087 (N_13087,N_10482,N_11074);
and U13088 (N_13088,N_9024,N_11420);
nand U13089 (N_13089,N_9364,N_11956);
xor U13090 (N_13090,N_9581,N_8610);
and U13091 (N_13091,N_11853,N_9192);
xnor U13092 (N_13092,N_10073,N_11744);
or U13093 (N_13093,N_8070,N_9354);
nand U13094 (N_13094,N_11740,N_8937);
nand U13095 (N_13095,N_11156,N_10521);
or U13096 (N_13096,N_10332,N_10443);
nand U13097 (N_13097,N_8723,N_9524);
and U13098 (N_13098,N_10662,N_11929);
xnor U13099 (N_13099,N_9455,N_9418);
and U13100 (N_13100,N_9777,N_10544);
or U13101 (N_13101,N_8126,N_10532);
nor U13102 (N_13102,N_10853,N_8573);
nand U13103 (N_13103,N_8137,N_8713);
and U13104 (N_13104,N_8588,N_9132);
nor U13105 (N_13105,N_8471,N_8663);
and U13106 (N_13106,N_9069,N_8968);
or U13107 (N_13107,N_8341,N_11279);
nor U13108 (N_13108,N_9512,N_11017);
and U13109 (N_13109,N_10320,N_11762);
xor U13110 (N_13110,N_8306,N_11851);
nor U13111 (N_13111,N_8049,N_10028);
or U13112 (N_13112,N_9323,N_11372);
and U13113 (N_13113,N_9339,N_8617);
and U13114 (N_13114,N_10193,N_11501);
or U13115 (N_13115,N_10445,N_9220);
and U13116 (N_13116,N_10786,N_8819);
or U13117 (N_13117,N_9272,N_8170);
nor U13118 (N_13118,N_8114,N_8271);
nand U13119 (N_13119,N_8838,N_8586);
or U13120 (N_13120,N_9052,N_10879);
nand U13121 (N_13121,N_9703,N_10306);
nand U13122 (N_13122,N_10676,N_11665);
xor U13123 (N_13123,N_10349,N_9134);
nor U13124 (N_13124,N_10696,N_8957);
or U13125 (N_13125,N_9728,N_10324);
or U13126 (N_13126,N_11536,N_11200);
nor U13127 (N_13127,N_8502,N_10774);
and U13128 (N_13128,N_11484,N_11885);
nor U13129 (N_13129,N_8800,N_9941);
and U13130 (N_13130,N_11821,N_10192);
or U13131 (N_13131,N_11805,N_11707);
nor U13132 (N_13132,N_9647,N_10336);
or U13133 (N_13133,N_9670,N_8771);
nor U13134 (N_13134,N_11845,N_8332);
nand U13135 (N_13135,N_11666,N_8512);
nand U13136 (N_13136,N_10902,N_11064);
or U13137 (N_13137,N_8238,N_9772);
nand U13138 (N_13138,N_11709,N_8987);
or U13139 (N_13139,N_8199,N_9879);
or U13140 (N_13140,N_10006,N_9897);
and U13141 (N_13141,N_11611,N_9474);
and U13142 (N_13142,N_8105,N_10932);
nor U13143 (N_13143,N_10065,N_9672);
or U13144 (N_13144,N_9759,N_10743);
or U13145 (N_13145,N_11987,N_9026);
xor U13146 (N_13146,N_9967,N_11203);
nor U13147 (N_13147,N_9414,N_8528);
and U13148 (N_13148,N_11312,N_10530);
or U13149 (N_13149,N_9458,N_9906);
and U13150 (N_13150,N_9250,N_11061);
xor U13151 (N_13151,N_8314,N_11005);
and U13152 (N_13152,N_9553,N_8253);
or U13153 (N_13153,N_11483,N_8637);
nor U13154 (N_13154,N_9989,N_11321);
xnor U13155 (N_13155,N_11242,N_9374);
nor U13156 (N_13156,N_9398,N_10238);
or U13157 (N_13157,N_10809,N_10450);
nand U13158 (N_13158,N_11384,N_10603);
or U13159 (N_13159,N_8029,N_9053);
nand U13160 (N_13160,N_10061,N_9049);
nand U13161 (N_13161,N_11635,N_10899);
and U13162 (N_13162,N_8733,N_10220);
nor U13163 (N_13163,N_9071,N_10419);
xor U13164 (N_13164,N_11296,N_8596);
xnor U13165 (N_13165,N_8345,N_10928);
or U13166 (N_13166,N_9591,N_9745);
or U13167 (N_13167,N_8755,N_8312);
or U13168 (N_13168,N_8860,N_11654);
nor U13169 (N_13169,N_9336,N_9686);
nor U13170 (N_13170,N_10433,N_9212);
nor U13171 (N_13171,N_9595,N_11913);
and U13172 (N_13172,N_9508,N_10548);
xor U13173 (N_13173,N_8561,N_9032);
nand U13174 (N_13174,N_8293,N_9814);
nand U13175 (N_13175,N_8472,N_9746);
nand U13176 (N_13176,N_10526,N_11587);
nand U13177 (N_13177,N_8402,N_8221);
nand U13178 (N_13178,N_9287,N_8717);
nand U13179 (N_13179,N_8803,N_9737);
nand U13180 (N_13180,N_10499,N_10448);
and U13181 (N_13181,N_9023,N_11904);
nand U13182 (N_13182,N_11103,N_9131);
nor U13183 (N_13183,N_8301,N_8727);
or U13184 (N_13184,N_9900,N_11133);
and U13185 (N_13185,N_8212,N_8217);
xor U13186 (N_13186,N_10380,N_11140);
or U13187 (N_13187,N_8883,N_10382);
xor U13188 (N_13188,N_10977,N_10333);
nor U13189 (N_13189,N_11113,N_8405);
and U13190 (N_13190,N_10724,N_10926);
or U13191 (N_13191,N_10704,N_8051);
and U13192 (N_13192,N_9101,N_11563);
nand U13193 (N_13193,N_9803,N_10610);
or U13194 (N_13194,N_8097,N_8322);
nor U13195 (N_13195,N_8634,N_9076);
or U13196 (N_13196,N_11220,N_10757);
nor U13197 (N_13197,N_9047,N_11933);
nor U13198 (N_13198,N_10938,N_11548);
and U13199 (N_13199,N_11673,N_10539);
or U13200 (N_13200,N_10260,N_9232);
nor U13201 (N_13201,N_9247,N_9117);
and U13202 (N_13202,N_8272,N_9925);
nand U13203 (N_13203,N_11942,N_10889);
and U13204 (N_13204,N_11058,N_10144);
nor U13205 (N_13205,N_10876,N_9757);
and U13206 (N_13206,N_9516,N_10034);
or U13207 (N_13207,N_11008,N_8907);
nand U13208 (N_13208,N_11895,N_11663);
nor U13209 (N_13209,N_9261,N_10049);
and U13210 (N_13210,N_9845,N_8291);
and U13211 (N_13211,N_9087,N_8003);
or U13212 (N_13212,N_11585,N_11115);
xnor U13213 (N_13213,N_10974,N_8598);
xnor U13214 (N_13214,N_8952,N_8203);
nand U13215 (N_13215,N_10655,N_9176);
nor U13216 (N_13216,N_9484,N_9692);
xor U13217 (N_13217,N_8926,N_8726);
nand U13218 (N_13218,N_11627,N_11940);
nand U13219 (N_13219,N_8582,N_11485);
nand U13220 (N_13220,N_8338,N_8117);
and U13221 (N_13221,N_10642,N_10128);
or U13222 (N_13222,N_11939,N_9885);
and U13223 (N_13223,N_11995,N_11789);
nor U13224 (N_13224,N_10943,N_9515);
and U13225 (N_13225,N_10111,N_9929);
and U13226 (N_13226,N_11528,N_9727);
nand U13227 (N_13227,N_10855,N_11850);
nand U13228 (N_13228,N_9866,N_11258);
xnor U13229 (N_13229,N_9810,N_8249);
and U13230 (N_13230,N_11172,N_10792);
and U13231 (N_13231,N_10007,N_10843);
nor U13232 (N_13232,N_8010,N_11454);
nand U13233 (N_13233,N_10489,N_10305);
or U13234 (N_13234,N_8709,N_10354);
nor U13235 (N_13235,N_9763,N_9738);
xnor U13236 (N_13236,N_9396,N_9303);
and U13237 (N_13237,N_10653,N_10345);
nand U13238 (N_13238,N_10604,N_10664);
or U13239 (N_13239,N_9375,N_11667);
or U13240 (N_13240,N_11965,N_11271);
nor U13241 (N_13241,N_8187,N_9019);
nand U13242 (N_13242,N_11254,N_10594);
or U13243 (N_13243,N_10066,N_11715);
nand U13244 (N_13244,N_11154,N_11150);
nand U13245 (N_13245,N_9678,N_8232);
nand U13246 (N_13246,N_8215,N_9111);
nand U13247 (N_13247,N_10877,N_11676);
and U13248 (N_13248,N_10424,N_10440);
or U13249 (N_13249,N_8567,N_9993);
nand U13250 (N_13250,N_8995,N_10523);
and U13251 (N_13251,N_10249,N_10278);
and U13252 (N_13252,N_9274,N_9533);
nor U13253 (N_13253,N_8899,N_10187);
nor U13254 (N_13254,N_8043,N_11415);
and U13255 (N_13255,N_11262,N_10302);
and U13256 (N_13256,N_9029,N_8078);
or U13257 (N_13257,N_11957,N_8222);
nand U13258 (N_13258,N_9824,N_10177);
and U13259 (N_13259,N_9571,N_11660);
and U13260 (N_13260,N_10241,N_9931);
or U13261 (N_13261,N_9543,N_10970);
nor U13262 (N_13262,N_8201,N_9245);
and U13263 (N_13263,N_11087,N_11016);
or U13264 (N_13264,N_10697,N_11306);
and U13265 (N_13265,N_10168,N_11525);
nand U13266 (N_13266,N_8394,N_8009);
nor U13267 (N_13267,N_11486,N_9848);
or U13268 (N_13268,N_11948,N_10393);
nor U13269 (N_13269,N_10083,N_9439);
and U13270 (N_13270,N_9299,N_11702);
nand U13271 (N_13271,N_10745,N_8976);
xor U13272 (N_13272,N_11539,N_8674);
and U13273 (N_13273,N_8167,N_8643);
and U13274 (N_13274,N_8021,N_10501);
or U13275 (N_13275,N_8964,N_8395);
nand U13276 (N_13276,N_8136,N_8938);
or U13277 (N_13277,N_11303,N_10012);
nor U13278 (N_13278,N_8166,N_11098);
and U13279 (N_13279,N_8151,N_11409);
or U13280 (N_13280,N_8597,N_8658);
nand U13281 (N_13281,N_11349,N_10847);
or U13282 (N_13282,N_9924,N_9990);
or U13283 (N_13283,N_11298,N_11120);
or U13284 (N_13284,N_8363,N_9300);
or U13285 (N_13285,N_9329,N_11340);
nand U13286 (N_13286,N_11820,N_10112);
nor U13287 (N_13287,N_11131,N_8466);
nand U13288 (N_13288,N_9874,N_11870);
nand U13289 (N_13289,N_10387,N_9797);
or U13290 (N_13290,N_11854,N_8015);
or U13291 (N_13291,N_10092,N_8863);
nor U13292 (N_13292,N_9397,N_11192);
or U13293 (N_13293,N_11575,N_8336);
nor U13294 (N_13294,N_9709,N_11316);
nor U13295 (N_13295,N_9493,N_9347);
nor U13296 (N_13296,N_8250,N_11056);
xnor U13297 (N_13297,N_9731,N_11439);
and U13298 (N_13298,N_8559,N_11926);
and U13299 (N_13299,N_9082,N_8908);
nand U13300 (N_13300,N_8171,N_8289);
or U13301 (N_13301,N_11973,N_10479);
nor U13302 (N_13302,N_8764,N_11166);
and U13303 (N_13303,N_11863,N_9334);
xnor U13304 (N_13304,N_9949,N_10759);
nor U13305 (N_13305,N_9890,N_10390);
and U13306 (N_13306,N_11747,N_8164);
nand U13307 (N_13307,N_10155,N_8041);
nor U13308 (N_13308,N_9041,N_8707);
nor U13309 (N_13309,N_10750,N_10329);
or U13310 (N_13310,N_8909,N_10921);
nand U13311 (N_13311,N_8654,N_8691);
xor U13312 (N_13312,N_9754,N_10229);
nor U13313 (N_13313,N_11421,N_9086);
nor U13314 (N_13314,N_8295,N_10976);
xnor U13315 (N_13315,N_8629,N_8657);
nand U13316 (N_13316,N_10631,N_8651);
or U13317 (N_13317,N_10024,N_10272);
and U13318 (N_13318,N_9182,N_9388);
nor U13319 (N_13319,N_11386,N_9666);
and U13320 (N_13320,N_10913,N_8706);
and U13321 (N_13321,N_9971,N_10599);
or U13322 (N_13322,N_10731,N_9130);
and U13323 (N_13323,N_10672,N_8989);
or U13324 (N_13324,N_10337,N_9341);
and U13325 (N_13325,N_11780,N_8675);
nor U13326 (N_13326,N_8205,N_11146);
and U13327 (N_13327,N_10145,N_8017);
and U13328 (N_13328,N_10292,N_8773);
and U13329 (N_13329,N_11694,N_9226);
or U13330 (N_13330,N_11423,N_9046);
nand U13331 (N_13331,N_8132,N_8743);
nor U13332 (N_13332,N_9276,N_11796);
nor U13333 (N_13333,N_9935,N_10556);
nor U13334 (N_13334,N_10078,N_10267);
and U13335 (N_13335,N_9093,N_9127);
xnor U13336 (N_13336,N_11769,N_9293);
and U13337 (N_13337,N_8034,N_9865);
nand U13338 (N_13338,N_8897,N_11570);
and U13339 (N_13339,N_9147,N_9554);
nor U13340 (N_13340,N_9195,N_9972);
nand U13341 (N_13341,N_8624,N_11652);
xnor U13342 (N_13342,N_10275,N_10982);
and U13343 (N_13343,N_11811,N_10838);
and U13344 (N_13344,N_11320,N_10226);
or U13345 (N_13345,N_8038,N_8158);
or U13346 (N_13346,N_11083,N_11301);
and U13347 (N_13347,N_9883,N_9718);
nand U13348 (N_13348,N_8148,N_9312);
and U13349 (N_13349,N_10611,N_8065);
nand U13350 (N_13350,N_8966,N_9216);
or U13351 (N_13351,N_10299,N_11756);
xnor U13352 (N_13352,N_8612,N_9459);
xor U13353 (N_13353,N_10116,N_9395);
and U13354 (N_13354,N_10062,N_8447);
or U13355 (N_13355,N_10136,N_9081);
and U13356 (N_13356,N_11455,N_10867);
and U13357 (N_13357,N_11338,N_9469);
or U13358 (N_13358,N_8465,N_11479);
nand U13359 (N_13359,N_11915,N_11963);
and U13360 (N_13360,N_11389,N_10985);
and U13361 (N_13361,N_11102,N_8788);
xor U13362 (N_13362,N_11924,N_9257);
nor U13363 (N_13363,N_11106,N_9179);
or U13364 (N_13364,N_8355,N_8303);
and U13365 (N_13365,N_11359,N_8054);
nor U13366 (N_13366,N_8406,N_9394);
nand U13367 (N_13367,N_11014,N_11040);
or U13368 (N_13368,N_11669,N_11280);
nor U13369 (N_13369,N_8521,N_10362);
nand U13370 (N_13370,N_11274,N_11275);
nand U13371 (N_13371,N_11826,N_10781);
nor U13372 (N_13372,N_8955,N_10656);
nand U13373 (N_13373,N_11992,N_10538);
xor U13374 (N_13374,N_10871,N_9802);
and U13375 (N_13375,N_11921,N_11297);
nand U13376 (N_13376,N_11228,N_10313);
nand U13377 (N_13377,N_10150,N_10224);
and U13378 (N_13378,N_8701,N_10835);
or U13379 (N_13379,N_10105,N_10751);
nor U13380 (N_13380,N_10545,N_8500);
nor U13381 (N_13381,N_9114,N_9438);
nor U13382 (N_13382,N_9590,N_8032);
and U13383 (N_13383,N_9413,N_9311);
or U13384 (N_13384,N_10803,N_8932);
nand U13385 (N_13385,N_9135,N_10942);
xnor U13386 (N_13386,N_11938,N_11549);
nor U13387 (N_13387,N_9256,N_8729);
xnor U13388 (N_13388,N_10201,N_8943);
xnor U13389 (N_13389,N_11852,N_8846);
nand U13390 (N_13390,N_11488,N_10365);
or U13391 (N_13391,N_11447,N_11267);
nor U13392 (N_13392,N_10307,N_11700);
nor U13393 (N_13393,N_10825,N_9652);
or U13394 (N_13394,N_9855,N_8188);
xor U13395 (N_13395,N_8759,N_9775);
or U13396 (N_13396,N_8944,N_8284);
nand U13397 (N_13397,N_8919,N_8310);
or U13398 (N_13398,N_10137,N_10153);
nor U13399 (N_13399,N_11745,N_11696);
and U13400 (N_13400,N_11265,N_11196);
and U13401 (N_13401,N_11355,N_11193);
or U13402 (N_13402,N_11272,N_8050);
and U13403 (N_13403,N_10321,N_11033);
nand U13404 (N_13404,N_9798,N_8450);
nand U13405 (N_13405,N_10085,N_8772);
nor U13406 (N_13406,N_10636,N_11463);
and U13407 (N_13407,N_9006,N_10587);
xnor U13408 (N_13408,N_8696,N_10691);
nor U13409 (N_13409,N_10411,N_9072);
or U13410 (N_13410,N_8763,N_10173);
and U13411 (N_13411,N_10769,N_10677);
and U13412 (N_13412,N_11728,N_9966);
and U13413 (N_13413,N_9576,N_8758);
nor U13414 (N_13414,N_11908,N_11888);
nand U13415 (N_13415,N_9736,N_8782);
xor U13416 (N_13416,N_11067,N_8392);
xnor U13417 (N_13417,N_10810,N_11369);
nand U13418 (N_13418,N_8438,N_10821);
or U13419 (N_13419,N_10067,N_11091);
and U13420 (N_13420,N_10965,N_10395);
nor U13421 (N_13421,N_11692,N_11680);
nor U13422 (N_13422,N_9056,N_10773);
or U13423 (N_13423,N_9172,N_11358);
and U13424 (N_13424,N_11819,N_11761);
and U13425 (N_13425,N_11094,N_8900);
nand U13426 (N_13426,N_10787,N_8954);
nor U13427 (N_13427,N_11788,N_8403);
or U13428 (N_13428,N_10350,N_10480);
or U13429 (N_13429,N_9847,N_10592);
xor U13430 (N_13430,N_10164,N_10606);
or U13431 (N_13431,N_8285,N_9895);
nor U13432 (N_13432,N_8248,N_10805);
and U13433 (N_13433,N_11509,N_9696);
nor U13434 (N_13434,N_9297,N_9392);
nand U13435 (N_13435,N_9788,N_8055);
or U13436 (N_13436,N_8283,N_8616);
nor U13437 (N_13437,N_9801,N_10139);
nand U13438 (N_13438,N_10327,N_10280);
nand U13439 (N_13439,N_9043,N_11581);
nor U13440 (N_13440,N_8080,N_8622);
and U13441 (N_13441,N_8600,N_11759);
or U13442 (N_13442,N_8700,N_8714);
or U13443 (N_13443,N_11558,N_11884);
or U13444 (N_13444,N_10622,N_10197);
nor U13445 (N_13445,N_10983,N_8211);
xnor U13446 (N_13446,N_10998,N_11518);
and U13447 (N_13447,N_11867,N_8704);
and U13448 (N_13448,N_9361,N_8220);
or U13449 (N_13449,N_8811,N_9419);
nor U13450 (N_13450,N_11066,N_8266);
or U13451 (N_13451,N_8553,N_10404);
or U13452 (N_13452,N_8790,N_11108);
or U13453 (N_13453,N_10217,N_9877);
or U13454 (N_13454,N_8921,N_8719);
nand U13455 (N_13455,N_10824,N_8012);
or U13456 (N_13456,N_10766,N_11490);
xor U13457 (N_13457,N_11726,N_11961);
nand U13458 (N_13458,N_8534,N_10756);
nand U13459 (N_13459,N_9760,N_9153);
or U13460 (N_13460,N_10439,N_11049);
nand U13461 (N_13461,N_10019,N_8325);
nor U13462 (N_13462,N_9752,N_8382);
nand U13463 (N_13463,N_8058,N_9421);
nor U13464 (N_13464,N_8209,N_11427);
or U13465 (N_13465,N_11238,N_10830);
nor U13466 (N_13466,N_10361,N_8470);
nand U13467 (N_13467,N_8977,N_8787);
nor U13468 (N_13468,N_10422,N_10408);
xor U13469 (N_13469,N_9028,N_11476);
or U13470 (N_13470,N_9592,N_10541);
and U13471 (N_13471,N_9839,N_11418);
nand U13472 (N_13472,N_8145,N_9876);
nor U13473 (N_13473,N_10868,N_9440);
and U13474 (N_13474,N_9926,N_10614);
and U13475 (N_13475,N_8768,N_8698);
and U13476 (N_13476,N_9284,N_8230);
and U13477 (N_13477,N_8914,N_10047);
or U13478 (N_13478,N_10115,N_8490);
nand U13479 (N_13479,N_10163,N_8118);
or U13480 (N_13480,N_11670,N_10531);
or U13481 (N_13481,N_8981,N_11554);
xor U13482 (N_13482,N_9585,N_10562);
nor U13483 (N_13483,N_8157,N_8393);
nor U13484 (N_13484,N_8650,N_8767);
or U13485 (N_13485,N_11768,N_11741);
and U13486 (N_13486,N_8915,N_10328);
nor U13487 (N_13487,N_9106,N_8037);
and U13488 (N_13488,N_8252,N_8951);
or U13489 (N_13489,N_8416,N_8826);
nor U13490 (N_13490,N_11571,N_11036);
nor U13491 (N_13491,N_9540,N_9570);
or U13492 (N_13492,N_8988,N_8812);
nand U13493 (N_13493,N_10832,N_8497);
and U13494 (N_13494,N_10107,N_9042);
nand U13495 (N_13495,N_11435,N_11408);
and U13496 (N_13496,N_11565,N_10734);
and U13497 (N_13497,N_9635,N_11145);
xor U13498 (N_13498,N_10121,N_9252);
nor U13499 (N_13499,N_8204,N_10715);
and U13500 (N_13500,N_10500,N_8854);
xnor U13501 (N_13501,N_10869,N_11213);
nand U13502 (N_13502,N_11801,N_8834);
nor U13503 (N_13503,N_11914,N_10318);
and U13504 (N_13504,N_10140,N_9231);
nand U13505 (N_13505,N_8408,N_11489);
and U13506 (N_13506,N_11552,N_11547);
nor U13507 (N_13507,N_11583,N_8337);
and U13508 (N_13508,N_8258,N_10841);
or U13509 (N_13509,N_9575,N_9740);
and U13510 (N_13510,N_10851,N_9335);
nor U13511 (N_13511,N_11225,N_10528);
nor U13512 (N_13512,N_11308,N_8982);
nor U13513 (N_13513,N_10808,N_8202);
and U13514 (N_13514,N_9489,N_11723);
nand U13515 (N_13515,N_11240,N_11872);
and U13516 (N_13516,N_8496,N_8075);
and U13517 (N_13517,N_10401,N_8356);
nand U13518 (N_13518,N_8195,N_11392);
nor U13519 (N_13519,N_9655,N_11393);
and U13520 (N_13520,N_8330,N_10577);
and U13521 (N_13521,N_11724,N_10181);
and U13522 (N_13522,N_8459,N_10688);
nor U13523 (N_13523,N_8557,N_11204);
or U13524 (N_13524,N_8327,N_11398);
and U13525 (N_13525,N_11943,N_9366);
or U13526 (N_13526,N_11284,N_9473);
nor U13527 (N_13527,N_9084,N_10435);
or U13528 (N_13528,N_10301,N_10087);
and U13529 (N_13529,N_10235,N_8265);
or U13530 (N_13530,N_10650,N_10160);
nor U13531 (N_13531,N_9735,N_10850);
and U13532 (N_13532,N_11603,N_10816);
or U13533 (N_13533,N_10890,N_11350);
nand U13534 (N_13534,N_8092,N_10822);
or U13535 (N_13535,N_10680,N_11515);
nor U13536 (N_13536,N_11202,N_9263);
nand U13537 (N_13537,N_8173,N_10681);
nor U13538 (N_13538,N_11093,N_10344);
and U13539 (N_13539,N_10165,N_10033);
nor U13540 (N_13540,N_11899,N_11618);
or U13541 (N_13541,N_10586,N_11510);
nor U13542 (N_13542,N_8260,N_9641);
and U13543 (N_13543,N_9659,N_11314);
and U13544 (N_13544,N_9715,N_10270);
nand U13545 (N_13545,N_8449,N_10074);
nor U13546 (N_13546,N_11357,N_10692);
and U13547 (N_13547,N_11532,N_10818);
nand U13548 (N_13548,N_11401,N_9165);
and U13549 (N_13549,N_8660,N_10277);
xnor U13550 (N_13550,N_11022,N_11589);
and U13551 (N_13551,N_9409,N_10088);
and U13552 (N_13552,N_11051,N_11748);
and U13553 (N_13553,N_9779,N_10104);
and U13554 (N_13554,N_11176,N_9359);
and U13555 (N_13555,N_8267,N_10247);
nand U13556 (N_13556,N_11843,N_10907);
and U13557 (N_13557,N_10300,N_11440);
xor U13558 (N_13558,N_11382,N_11684);
and U13559 (N_13559,N_9309,N_11201);
and U13560 (N_13560,N_8121,N_10923);
and U13561 (N_13561,N_9910,N_9645);
nand U13562 (N_13562,N_11179,N_10188);
or U13563 (N_13563,N_11903,N_8664);
nand U13564 (N_13564,N_10485,N_11019);
or U13565 (N_13565,N_9556,N_10568);
and U13566 (N_13566,N_10118,N_9113);
and U13567 (N_13567,N_8694,N_11143);
or U13568 (N_13568,N_8103,N_8063);
nand U13569 (N_13569,N_9654,N_9479);
nand U13570 (N_13570,N_10765,N_8744);
nor U13571 (N_13571,N_9835,N_8965);
or U13572 (N_13572,N_11504,N_8479);
nand U13573 (N_13573,N_10488,N_8484);
nor U13574 (N_13574,N_9324,N_11960);
nand U13575 (N_13575,N_11964,N_9487);
or U13576 (N_13576,N_8367,N_11367);
and U13577 (N_13577,N_8206,N_9075);
xnor U13578 (N_13578,N_10436,N_11334);
and U13579 (N_13579,N_9514,N_11090);
nand U13580 (N_13580,N_8662,N_10881);
nor U13581 (N_13581,N_10829,N_11215);
xor U13582 (N_13582,N_10558,N_8141);
nand U13583 (N_13583,N_8647,N_8614);
or U13584 (N_13584,N_11815,N_9681);
nor U13585 (N_13585,N_9902,N_11045);
nand U13586 (N_13586,N_8855,N_10427);
or U13587 (N_13587,N_11118,N_8410);
nand U13588 (N_13588,N_9784,N_8210);
nand U13589 (N_13589,N_8841,N_8850);
and U13590 (N_13590,N_8036,N_9549);
or U13591 (N_13591,N_11060,N_8603);
xnor U13592 (N_13592,N_9673,N_8162);
nor U13593 (N_13593,N_9800,N_10325);
or U13594 (N_13594,N_9882,N_8462);
xnor U13595 (N_13595,N_10236,N_8587);
nor U13596 (N_13596,N_8123,N_9170);
or U13597 (N_13597,N_8608,N_11616);
nor U13598 (N_13598,N_10537,N_8476);
or U13599 (N_13599,N_8680,N_8762);
nand U13600 (N_13600,N_11226,N_9085);
and U13601 (N_13601,N_9406,N_11758);
nand U13602 (N_13602,N_11129,N_8439);
nor U13603 (N_13603,N_10287,N_8086);
nand U13604 (N_13604,N_8096,N_11586);
or U13605 (N_13605,N_10389,N_8234);
nor U13606 (N_13606,N_8237,N_8256);
xor U13607 (N_13607,N_11070,N_9831);
xnor U13608 (N_13608,N_8082,N_10265);
nor U13609 (N_13609,N_11160,N_10863);
and U13610 (N_13610,N_10050,N_8888);
xor U13611 (N_13611,N_10785,N_10971);
nand U13612 (N_13612,N_11004,N_9699);
and U13613 (N_13613,N_8681,N_9188);
xor U13614 (N_13614,N_8606,N_9583);
and U13615 (N_13615,N_8101,N_9765);
and U13616 (N_13616,N_11920,N_11135);
and U13617 (N_13617,N_9416,N_10717);
and U13618 (N_13618,N_11445,N_9509);
and U13619 (N_13619,N_10903,N_10694);
and U13620 (N_13620,N_8746,N_10771);
nor U13621 (N_13621,N_10678,N_11659);
or U13622 (N_13622,N_10471,N_11678);
nor U13623 (N_13623,N_9465,N_10952);
or U13624 (N_13624,N_10043,N_11997);
and U13625 (N_13625,N_10605,N_9144);
xnor U13626 (N_13626,N_8527,N_9690);
nand U13627 (N_13627,N_9973,N_9534);
xnor U13628 (N_13628,N_10516,N_9630);
or U13629 (N_13629,N_10827,N_11630);
or U13630 (N_13630,N_8150,N_11288);
nand U13631 (N_13631,N_11123,N_8632);
or U13632 (N_13632,N_10143,N_10716);
or U13633 (N_13633,N_10645,N_9073);
nand U13634 (N_13634,N_10364,N_11475);
or U13635 (N_13635,N_11787,N_8307);
nor U13636 (N_13636,N_8911,N_10513);
or U13637 (N_13637,N_11538,N_11266);
xnor U13638 (N_13638,N_9864,N_11075);
or U13639 (N_13639,N_11318,N_9589);
nand U13640 (N_13640,N_8687,N_8515);
nand U13641 (N_13641,N_9804,N_10009);
or U13642 (N_13642,N_8110,N_9978);
and U13643 (N_13643,N_10097,N_10812);
and U13644 (N_13644,N_10959,N_11970);
or U13645 (N_13645,N_10951,N_11828);
or U13646 (N_13646,N_10560,N_10484);
or U13647 (N_13647,N_11317,N_8401);
or U13648 (N_13648,N_10186,N_8642);
nand U13649 (N_13649,N_8331,N_10772);
or U13650 (N_13650,N_9922,N_8161);
or U13651 (N_13651,N_11645,N_8748);
nand U13652 (N_13652,N_11136,N_9710);
and U13653 (N_13653,N_8836,N_11034);
nand U13654 (N_13654,N_10071,N_8532);
or U13655 (N_13655,N_10015,N_10887);
or U13656 (N_13656,N_8649,N_9809);
xnor U13657 (N_13657,N_9507,N_11701);
nor U13658 (N_13658,N_11881,N_10208);
xor U13659 (N_13659,N_8934,N_10036);
or U13660 (N_13660,N_11194,N_8574);
nand U13661 (N_13661,N_9714,N_9222);
or U13662 (N_13662,N_8453,N_9251);
nand U13663 (N_13663,N_10001,N_10415);
nor U13664 (N_13664,N_9424,N_8940);
and U13665 (N_13665,N_8264,N_10885);
nor U13666 (N_13666,N_11380,N_10778);
or U13667 (N_13667,N_11063,N_8178);
and U13668 (N_13668,N_11531,N_8581);
or U13669 (N_13669,N_11434,N_11859);
nand U13670 (N_13670,N_9603,N_8695);
nand U13671 (N_13671,N_11541,N_11219);
nor U13672 (N_13672,N_11032,N_10909);
or U13673 (N_13673,N_9653,N_11753);
and U13674 (N_13674,N_10858,N_10831);
nor U13675 (N_13675,N_9579,N_11183);
or U13676 (N_13676,N_11385,N_11346);
or U13677 (N_13677,N_11079,N_10518);
and U13678 (N_13678,N_10461,N_9389);
xor U13679 (N_13679,N_11542,N_10840);
nand U13680 (N_13680,N_8369,N_8276);
xnor U13681 (N_13681,N_8246,N_9277);
or U13682 (N_13682,N_10826,N_9675);
nor U13683 (N_13683,N_9021,N_8441);
nand U13684 (N_13684,N_8505,N_11530);
and U13685 (N_13685,N_10169,N_9333);
and U13686 (N_13686,N_10331,N_9353);
nor U13687 (N_13687,N_11470,N_9517);
xor U13688 (N_13688,N_10770,N_11617);
and U13689 (N_13689,N_8858,N_9168);
and U13690 (N_13690,N_11522,N_11422);
or U13691 (N_13691,N_10182,N_10591);
and U13692 (N_13692,N_9158,N_8362);
nor U13693 (N_13693,N_10117,N_10276);
xnor U13694 (N_13694,N_10975,N_9601);
nor U13695 (N_13695,N_11844,N_10223);
and U13696 (N_13696,N_9644,N_8129);
or U13697 (N_13697,N_8807,N_11286);
nor U13698 (N_13698,N_8892,N_9572);
and U13699 (N_13699,N_10057,N_11982);
nand U13700 (N_13700,N_10878,N_11038);
or U13701 (N_13701,N_10068,N_9778);
nand U13702 (N_13702,N_9463,N_8923);
nor U13703 (N_13703,N_9228,N_8094);
nor U13704 (N_13704,N_10291,N_11221);
xnor U13705 (N_13705,N_9036,N_11633);
and U13706 (N_13706,N_10141,N_9253);
and U13707 (N_13707,N_9604,N_8491);
or U13708 (N_13708,N_10888,N_9758);
and U13709 (N_13709,N_8443,N_8766);
or U13710 (N_13710,N_9943,N_10866);
nand U13711 (N_13711,N_8626,N_11855);
and U13712 (N_13712,N_9918,N_9503);
nor U13713 (N_13713,N_11163,N_8398);
or U13714 (N_13714,N_11184,N_9614);
and U13715 (N_13715,N_9711,N_11560);
nand U13716 (N_13716,N_10651,N_8801);
nand U13717 (N_13717,N_10947,N_8538);
xnor U13718 (N_13718,N_8390,N_8828);
or U13719 (N_13719,N_10527,N_10060);
nand U13720 (N_13720,N_9386,N_10084);
and U13721 (N_13721,N_10955,N_10341);
and U13722 (N_13722,N_10339,N_10470);
and U13723 (N_13723,N_11875,N_9462);
and U13724 (N_13724,N_8604,N_8776);
and U13725 (N_13725,N_8715,N_8945);
nand U13726 (N_13726,N_10026,N_10882);
or U13727 (N_13727,N_9350,N_9161);
nor U13728 (N_13728,N_10618,N_11502);
nand U13729 (N_13729,N_9229,N_11917);
nand U13730 (N_13730,N_11052,N_11428);
or U13731 (N_13731,N_11687,N_8958);
nand U13732 (N_13732,N_11722,N_11983);
and U13733 (N_13733,N_8437,N_11716);
nand U13734 (N_13734,N_10979,N_11224);
or U13735 (N_13735,N_9362,N_9385);
nand U13736 (N_13736,N_9695,N_9716);
nor U13737 (N_13737,N_9094,N_9861);
nor U13738 (N_13738,N_10431,N_9730);
or U13739 (N_13739,N_10621,N_11376);
and U13740 (N_13740,N_8446,N_8365);
xnor U13741 (N_13741,N_8565,N_8928);
nor U13742 (N_13742,N_10583,N_10396);
nor U13743 (N_13743,N_11309,N_9208);
or U13744 (N_13744,N_11342,N_9956);
and U13745 (N_13745,N_11236,N_10675);
nand U13746 (N_13746,N_10481,N_11755);
nand U13747 (N_13747,N_9497,N_9405);
xor U13748 (N_13748,N_11009,N_8052);
xnor U13749 (N_13749,N_11095,N_10058);
or U13750 (N_13750,N_8387,N_11674);
xnor U13751 (N_13751,N_10897,N_8525);
nor U13752 (N_13752,N_10684,N_10791);
nor U13753 (N_13753,N_11195,N_8636);
xor U13754 (N_13754,N_10377,N_11003);
nand U13755 (N_13755,N_9290,N_8942);
or U13756 (N_13756,N_11784,N_9869);
xnor U13757 (N_13757,N_8753,N_10090);
xnor U13758 (N_13758,N_9105,N_10458);
nor U13759 (N_13759,N_8290,N_11024);
or U13760 (N_13760,N_10290,N_8268);
xor U13761 (N_13761,N_9167,N_9694);
and U13762 (N_13762,N_10269,N_10190);
xnor U13763 (N_13763,N_11354,N_10687);
or U13764 (N_13764,N_10571,N_10652);
nand U13765 (N_13765,N_11590,N_8736);
nand U13766 (N_13766,N_10072,N_8375);
nor U13767 (N_13767,N_11323,N_9527);
xnor U13768 (N_13768,N_11264,N_11588);
xnor U13769 (N_13769,N_8493,N_10641);
and U13770 (N_13770,N_9701,N_8440);
nor U13771 (N_13771,N_8618,N_8144);
or U13772 (N_13772,N_11147,N_9358);
and U13773 (N_13773,N_9812,N_8949);
nand U13774 (N_13774,N_10212,N_10132);
or U13775 (N_13775,N_8620,N_11773);
and U13776 (N_13776,N_10317,N_8668);
xnor U13777 (N_13777,N_8108,N_8175);
nor U13778 (N_13778,N_9004,N_10891);
xnor U13779 (N_13779,N_9729,N_8135);
xor U13780 (N_13780,N_11879,N_11482);
xor U13781 (N_13781,N_10918,N_11672);
and U13782 (N_13782,N_9691,N_11390);
nand U13783 (N_13783,N_9233,N_8745);
or U13784 (N_13784,N_11906,N_10149);
xnor U13785 (N_13785,N_8593,N_8033);
and U13786 (N_13786,N_10232,N_8093);
or U13787 (N_13787,N_11634,N_11865);
nor U13788 (N_13788,N_9704,N_11564);
nor U13789 (N_13789,N_11436,N_11028);
nand U13790 (N_13790,N_9987,N_9997);
nand U13791 (N_13791,N_11559,N_8840);
nand U13792 (N_13792,N_10609,N_8189);
and U13793 (N_13793,N_10898,N_10749);
nand U13794 (N_13794,N_9415,N_8461);
nand U13795 (N_13795,N_11827,N_8786);
or U13796 (N_13796,N_9492,N_9432);
nor U13797 (N_13797,N_8558,N_8428);
and U13798 (N_13798,N_10053,N_9103);
or U13799 (N_13799,N_9471,N_10597);
xnor U13800 (N_13800,N_11168,N_8179);
and U13801 (N_13801,N_11404,N_11031);
nor U13802 (N_13802,N_9472,N_11629);
or U13803 (N_13803,N_8805,N_8347);
nor U13804 (N_13804,N_10413,N_10284);
or U13805 (N_13805,N_11733,N_10615);
and U13806 (N_13806,N_11661,N_8656);
or U13807 (N_13807,N_11814,N_8348);
or U13808 (N_13808,N_9547,N_11508);
nor U13809 (N_13809,N_9298,N_9241);
nand U13810 (N_13810,N_8967,N_9994);
nand U13811 (N_13811,N_9209,N_11381);
or U13812 (N_13812,N_11776,N_11714);
and U13813 (N_13813,N_11857,N_9940);
nand U13814 (N_13814,N_10311,N_9953);
nor U13815 (N_13815,N_8825,N_9891);
and U13816 (N_13816,N_10014,N_9221);
nor U13817 (N_13817,N_8718,N_8513);
and U13818 (N_13818,N_11437,N_9390);
or U13819 (N_13819,N_10261,N_9200);
nand U13820 (N_13820,N_8085,N_9898);
or U13821 (N_13821,N_9781,N_8750);
nand U13822 (N_13822,N_9058,N_10158);
or U13823 (N_13823,N_8156,N_9169);
and U13824 (N_13824,N_8947,N_11608);
xor U13825 (N_13825,N_11326,N_10763);
xor U13826 (N_13826,N_10917,N_9913);
nor U13827 (N_13827,N_11656,N_9436);
and U13828 (N_13828,N_10031,N_11849);
or U13829 (N_13829,N_9062,N_9904);
nand U13830 (N_13830,N_8184,N_8571);
nand U13831 (N_13831,N_11218,N_9834);
and U13832 (N_13832,N_8519,N_8084);
or U13833 (N_13833,N_9089,N_11057);
xnor U13834 (N_13834,N_8984,N_8627);
or U13835 (N_13835,N_8442,N_10495);
nand U13836 (N_13836,N_10994,N_11444);
nand U13837 (N_13837,N_8578,N_9464);
xor U13838 (N_13838,N_10373,N_11211);
nand U13839 (N_13839,N_11513,N_10468);
and U13840 (N_13840,N_11944,N_11243);
and U13841 (N_13841,N_9905,N_10814);
nor U13842 (N_13842,N_9837,N_9092);
and U13843 (N_13843,N_11442,N_9923);
nor U13844 (N_13844,N_11905,N_10956);
and U13845 (N_13845,N_10679,N_9060);
and U13846 (N_13846,N_10593,N_10934);
nor U13847 (N_13847,N_8089,N_10849);
xnor U13848 (N_13848,N_10370,N_11605);
xor U13849 (N_13849,N_11210,N_11649);
nor U13850 (N_13850,N_8814,N_9766);
and U13851 (N_13851,N_11453,N_11893);
nand U13852 (N_13852,N_10131,N_10739);
nor U13853 (N_13853,N_10732,N_8703);
and U13854 (N_13854,N_11449,N_11149);
and U13855 (N_13855,N_9377,N_11946);
nor U13856 (N_13856,N_9110,N_8514);
and U13857 (N_13857,N_9998,N_8379);
nor U13858 (N_13858,N_10109,N_9617);
or U13859 (N_13859,N_11467,N_9597);
nor U13860 (N_13860,N_11919,N_9050);
and U13861 (N_13861,N_11322,N_9494);
nor U13862 (N_13862,N_11543,N_8294);
xor U13863 (N_13863,N_11897,N_9780);
and U13864 (N_13864,N_11840,N_8251);
or U13865 (N_13865,N_8366,N_9118);
nand U13866 (N_13866,N_11623,N_9767);
and U13867 (N_13867,N_9657,N_11377);
nand U13868 (N_13868,N_10995,N_10710);
nor U13869 (N_13869,N_10595,N_10534);
nor U13870 (N_13870,N_9606,N_8857);
xor U13871 (N_13871,N_9770,N_11474);
or U13872 (N_13872,N_10282,N_8409);
xor U13873 (N_13873,N_10198,N_10472);
or U13874 (N_13874,N_11834,N_8962);
nor U13875 (N_13875,N_8859,N_8236);
xnor U13876 (N_13876,N_8991,N_9621);
or U13877 (N_13877,N_8060,N_9562);
nand U13878 (N_13878,N_9528,N_11551);
nand U13879 (N_13879,N_8334,N_11931);
or U13880 (N_13880,N_8088,N_10108);
nand U13881 (N_13881,N_10454,N_11012);
nand U13882 (N_13882,N_10993,N_10496);
and U13883 (N_13883,N_8335,N_8997);
or U13884 (N_13884,N_11030,N_10254);
nand U13885 (N_13885,N_9163,N_9942);
or U13886 (N_13886,N_11116,N_10573);
nor U13887 (N_13887,N_11344,N_9352);
nand U13888 (N_13888,N_9852,N_11883);
or U13889 (N_13889,N_8679,N_11876);
nand U13890 (N_13890,N_8712,N_10059);
nand U13891 (N_13891,N_11910,N_9682);
nand U13892 (N_13892,N_10964,N_9846);
or U13893 (N_13893,N_11839,N_11084);
or U13894 (N_13894,N_9878,N_9181);
or U13895 (N_13895,N_11935,N_9288);
xor U13896 (N_13896,N_11710,N_8595);
nand U13897 (N_13897,N_8452,N_10417);
nand U13898 (N_13898,N_8048,N_8590);
or U13899 (N_13899,N_8655,N_8741);
or U13900 (N_13900,N_8432,N_10310);
nand U13901 (N_13901,N_11846,N_11315);
or U13902 (N_13902,N_9938,N_8098);
and U13903 (N_13903,N_11699,N_11900);
or U13904 (N_13904,N_8673,N_8511);
or U13905 (N_13905,N_8802,N_11650);
and U13906 (N_13906,N_8004,N_8073);
nor U13907 (N_13907,N_8774,N_8978);
nand U13908 (N_13908,N_10629,N_11244);
nand U13909 (N_13909,N_9609,N_8473);
nand U13910 (N_13910,N_11685,N_10133);
or U13911 (N_13911,N_9328,N_11507);
xor U13912 (N_13912,N_8242,N_11671);
nand U13913 (N_13913,N_8853,N_9014);
nand U13914 (N_13914,N_9546,N_10206);
nor U13915 (N_13915,N_10412,N_11302);
and U13916 (N_13916,N_8192,N_11165);
nor U13917 (N_13917,N_9369,N_11366);
or U13918 (N_13918,N_11348,N_8510);
and U13919 (N_13919,N_8722,N_10230);
and U13920 (N_13920,N_8383,N_11023);
nor U13921 (N_13921,N_10122,N_9057);
nand U13922 (N_13922,N_9821,N_10649);
nand U13923 (N_13923,N_11754,N_8224);
and U13924 (N_13924,N_9100,N_8564);
nand U13925 (N_13925,N_10668,N_9602);
nor U13926 (N_13926,N_11319,N_11923);
or U13927 (N_13927,N_8839,N_9447);
or U13928 (N_13928,N_8482,N_8757);
or U13929 (N_13929,N_8308,N_8328);
or U13930 (N_13930,N_8866,N_10563);
nand U13931 (N_13931,N_11044,N_11695);
or U13932 (N_13932,N_10297,N_9083);
nand U13933 (N_13933,N_9764,N_11351);
nand U13934 (N_13934,N_9443,N_8520);
nand U13935 (N_13935,N_11792,N_9552);
nor U13936 (N_13936,N_10430,N_10086);
nand U13937 (N_13937,N_9936,N_8481);
nor U13938 (N_13938,N_10228,N_10936);
nor U13939 (N_13939,N_9741,N_11050);
nand U13940 (N_13940,N_10941,N_10989);
nor U13941 (N_13941,N_10465,N_11110);
or U13942 (N_13942,N_9618,N_11173);
nor U13943 (N_13943,N_11105,N_10601);
xnor U13944 (N_13944,N_8602,N_10003);
xor U13945 (N_13945,N_10246,N_9863);
and U13946 (N_13946,N_8113,N_11907);
and U13947 (N_13947,N_9326,N_9224);
xnor U13948 (N_13948,N_9511,N_11731);
xor U13949 (N_13949,N_8645,N_10753);
nand U13950 (N_13950,N_10798,N_8414);
or U13951 (N_13951,N_10402,N_9687);
or U13952 (N_13952,N_10159,N_8024);
nand U13953 (N_13953,N_11950,N_9496);
nor U13954 (N_13954,N_11018,N_11125);
nand U13955 (N_13955,N_9460,N_8804);
and U13956 (N_13956,N_10784,N_8193);
nand U13957 (N_13957,N_11972,N_8257);
or U13958 (N_13958,N_9078,N_10420);
nor U13959 (N_13959,N_8031,N_10243);
nor U13960 (N_13960,N_11443,N_9401);
nor U13961 (N_13961,N_9749,N_10884);
or U13962 (N_13962,N_10779,N_8820);
nor U13963 (N_13963,N_9651,N_9196);
nor U13964 (N_13964,N_9275,N_8946);
xnor U13965 (N_13965,N_9112,N_10366);
or U13966 (N_13966,N_8901,N_9946);
nand U13967 (N_13967,N_9550,N_8873);
nand U13968 (N_13968,N_11561,N_10455);
nand U13969 (N_13969,N_8316,N_9813);
nand U13970 (N_13970,N_11491,N_11797);
and U13971 (N_13971,N_10418,N_9269);
nand U13972 (N_13972,N_9148,N_11180);
nor U13973 (N_13973,N_9285,N_10806);
and U13974 (N_13974,N_11736,N_9838);
or U13975 (N_13975,N_9628,N_8342);
nand U13976 (N_13976,N_11818,N_9013);
or U13977 (N_13977,N_8756,N_10911);
nand U13978 (N_13978,N_9684,N_8448);
or U13979 (N_13979,N_9843,N_8548);
and U13980 (N_13980,N_10719,N_10040);
or U13981 (N_13981,N_10990,N_9518);
nor U13982 (N_13982,N_10469,N_11668);
nor U13983 (N_13983,N_10780,N_8815);
or U13984 (N_13984,N_9996,N_8789);
nor U13985 (N_13985,N_11214,N_10980);
xor U13986 (N_13986,N_8142,N_10227);
or U13987 (N_13987,N_9981,N_8879);
or U13988 (N_13988,N_11751,N_11750);
nand U13989 (N_13989,N_10180,N_11506);
nand U13990 (N_13990,N_9064,N_9823);
nor U13991 (N_13991,N_10077,N_10425);
nand U13992 (N_13992,N_8918,N_8927);
or U13993 (N_13993,N_9954,N_8507);
or U13994 (N_13994,N_11152,N_10288);
xnor U13995 (N_13995,N_8881,N_11082);
and U13996 (N_13996,N_8229,N_8044);
nand U13997 (N_13997,N_9536,N_10129);
or U13998 (N_13998,N_9568,N_11644);
and U13999 (N_13999,N_10507,N_10738);
and U14000 (N_14000,N_11997,N_8244);
nor U14001 (N_14001,N_10687,N_9705);
nand U14002 (N_14002,N_8254,N_8970);
and U14003 (N_14003,N_9765,N_8061);
nand U14004 (N_14004,N_11542,N_9784);
or U14005 (N_14005,N_10546,N_10181);
and U14006 (N_14006,N_8919,N_11621);
nand U14007 (N_14007,N_9300,N_11895);
nor U14008 (N_14008,N_10685,N_9124);
nand U14009 (N_14009,N_8518,N_9296);
or U14010 (N_14010,N_8917,N_9376);
nor U14011 (N_14011,N_9786,N_9351);
nor U14012 (N_14012,N_8476,N_9324);
nand U14013 (N_14013,N_9062,N_10564);
or U14014 (N_14014,N_11875,N_9647);
or U14015 (N_14015,N_10576,N_8674);
and U14016 (N_14016,N_11180,N_9684);
and U14017 (N_14017,N_8205,N_11570);
nand U14018 (N_14018,N_8878,N_9205);
and U14019 (N_14019,N_10098,N_8701);
nand U14020 (N_14020,N_8293,N_10344);
nor U14021 (N_14021,N_8523,N_8656);
nand U14022 (N_14022,N_11509,N_9171);
or U14023 (N_14023,N_11555,N_11796);
xor U14024 (N_14024,N_10000,N_8481);
nand U14025 (N_14025,N_9770,N_8373);
nand U14026 (N_14026,N_9070,N_10536);
or U14027 (N_14027,N_9477,N_10189);
nor U14028 (N_14028,N_11948,N_10275);
nand U14029 (N_14029,N_9624,N_10545);
or U14030 (N_14030,N_8327,N_9828);
and U14031 (N_14031,N_10507,N_10635);
nand U14032 (N_14032,N_10052,N_8799);
nor U14033 (N_14033,N_10191,N_9325);
and U14034 (N_14034,N_11586,N_10342);
and U14035 (N_14035,N_8715,N_11119);
or U14036 (N_14036,N_9277,N_10516);
nor U14037 (N_14037,N_8388,N_11548);
nor U14038 (N_14038,N_8988,N_11178);
nand U14039 (N_14039,N_11578,N_9840);
nand U14040 (N_14040,N_11847,N_8178);
xnor U14041 (N_14041,N_11162,N_10792);
and U14042 (N_14042,N_9314,N_11349);
xnor U14043 (N_14043,N_9605,N_8147);
or U14044 (N_14044,N_8322,N_11402);
xnor U14045 (N_14045,N_9320,N_10752);
and U14046 (N_14046,N_8883,N_10774);
and U14047 (N_14047,N_11568,N_10120);
nand U14048 (N_14048,N_10600,N_10471);
nand U14049 (N_14049,N_11427,N_11139);
nor U14050 (N_14050,N_11407,N_8759);
or U14051 (N_14051,N_8490,N_10137);
and U14052 (N_14052,N_10995,N_9409);
nand U14053 (N_14053,N_11203,N_9609);
nand U14054 (N_14054,N_10231,N_8121);
nor U14055 (N_14055,N_11058,N_11984);
or U14056 (N_14056,N_8239,N_10273);
nand U14057 (N_14057,N_10591,N_11381);
and U14058 (N_14058,N_11491,N_11974);
nand U14059 (N_14059,N_10095,N_9640);
nand U14060 (N_14060,N_10701,N_10297);
nor U14061 (N_14061,N_8456,N_9619);
or U14062 (N_14062,N_8291,N_8980);
or U14063 (N_14063,N_8419,N_10744);
and U14064 (N_14064,N_11942,N_10916);
nor U14065 (N_14065,N_8202,N_11600);
xnor U14066 (N_14066,N_8642,N_11191);
xnor U14067 (N_14067,N_8974,N_8679);
nand U14068 (N_14068,N_9921,N_11434);
and U14069 (N_14069,N_11498,N_10651);
nor U14070 (N_14070,N_9242,N_9408);
and U14071 (N_14071,N_11213,N_9614);
nand U14072 (N_14072,N_11199,N_10605);
nand U14073 (N_14073,N_11042,N_11105);
nor U14074 (N_14074,N_11743,N_10182);
nand U14075 (N_14075,N_9653,N_8207);
and U14076 (N_14076,N_9536,N_11315);
or U14077 (N_14077,N_10032,N_8645);
nand U14078 (N_14078,N_8408,N_9177);
nand U14079 (N_14079,N_9224,N_9448);
nand U14080 (N_14080,N_11653,N_10192);
xnor U14081 (N_14081,N_11833,N_8186);
nor U14082 (N_14082,N_8173,N_11208);
or U14083 (N_14083,N_8566,N_11579);
nand U14084 (N_14084,N_11661,N_9736);
or U14085 (N_14085,N_10992,N_9294);
nor U14086 (N_14086,N_8830,N_11298);
nand U14087 (N_14087,N_10394,N_8974);
or U14088 (N_14088,N_11127,N_8609);
nor U14089 (N_14089,N_8975,N_8320);
nor U14090 (N_14090,N_10134,N_10864);
nor U14091 (N_14091,N_9591,N_8640);
nor U14092 (N_14092,N_9298,N_10221);
or U14093 (N_14093,N_9988,N_9564);
nor U14094 (N_14094,N_9388,N_11412);
or U14095 (N_14095,N_11125,N_10008);
nand U14096 (N_14096,N_10409,N_8330);
or U14097 (N_14097,N_10129,N_11858);
nand U14098 (N_14098,N_11069,N_10408);
nor U14099 (N_14099,N_8203,N_8620);
nand U14100 (N_14100,N_8437,N_10208);
or U14101 (N_14101,N_11601,N_11850);
nand U14102 (N_14102,N_9243,N_10558);
nand U14103 (N_14103,N_8836,N_8211);
nor U14104 (N_14104,N_8676,N_10067);
nand U14105 (N_14105,N_9687,N_11432);
and U14106 (N_14106,N_9680,N_10143);
or U14107 (N_14107,N_10036,N_8111);
and U14108 (N_14108,N_8462,N_11635);
or U14109 (N_14109,N_10839,N_11342);
or U14110 (N_14110,N_10866,N_10186);
nor U14111 (N_14111,N_8770,N_8796);
or U14112 (N_14112,N_11744,N_10515);
nor U14113 (N_14113,N_9762,N_9592);
or U14114 (N_14114,N_8213,N_9476);
and U14115 (N_14115,N_8876,N_9207);
nand U14116 (N_14116,N_9696,N_9282);
nand U14117 (N_14117,N_8547,N_10072);
nand U14118 (N_14118,N_11328,N_11517);
and U14119 (N_14119,N_10597,N_10474);
xor U14120 (N_14120,N_8392,N_9690);
nand U14121 (N_14121,N_10680,N_11805);
nor U14122 (N_14122,N_10393,N_10056);
nand U14123 (N_14123,N_10140,N_10443);
and U14124 (N_14124,N_8462,N_9545);
or U14125 (N_14125,N_11917,N_9644);
or U14126 (N_14126,N_10058,N_9487);
nor U14127 (N_14127,N_8911,N_8889);
nand U14128 (N_14128,N_8151,N_11536);
or U14129 (N_14129,N_8485,N_9331);
nand U14130 (N_14130,N_11025,N_10402);
and U14131 (N_14131,N_11436,N_11567);
nand U14132 (N_14132,N_9596,N_11172);
nand U14133 (N_14133,N_10171,N_10558);
nor U14134 (N_14134,N_10185,N_11800);
nand U14135 (N_14135,N_8366,N_10027);
nor U14136 (N_14136,N_10219,N_9031);
nor U14137 (N_14137,N_11282,N_9505);
nand U14138 (N_14138,N_9781,N_10873);
and U14139 (N_14139,N_11311,N_10131);
nand U14140 (N_14140,N_8201,N_8864);
and U14141 (N_14141,N_11823,N_11762);
nand U14142 (N_14142,N_8269,N_9807);
or U14143 (N_14143,N_10248,N_10171);
and U14144 (N_14144,N_11923,N_11991);
and U14145 (N_14145,N_11039,N_9015);
nor U14146 (N_14146,N_10945,N_10510);
and U14147 (N_14147,N_9701,N_9867);
and U14148 (N_14148,N_10573,N_8009);
and U14149 (N_14149,N_9641,N_11976);
or U14150 (N_14150,N_11226,N_8800);
and U14151 (N_14151,N_10556,N_9054);
nor U14152 (N_14152,N_11559,N_8946);
nor U14153 (N_14153,N_9303,N_10590);
nor U14154 (N_14154,N_8582,N_11752);
nand U14155 (N_14155,N_9375,N_10942);
or U14156 (N_14156,N_8990,N_11662);
nand U14157 (N_14157,N_11485,N_8365);
and U14158 (N_14158,N_10373,N_8304);
nand U14159 (N_14159,N_10100,N_9900);
xnor U14160 (N_14160,N_9173,N_8793);
or U14161 (N_14161,N_10989,N_9192);
nor U14162 (N_14162,N_10471,N_10280);
nor U14163 (N_14163,N_11798,N_9002);
or U14164 (N_14164,N_9114,N_9675);
nand U14165 (N_14165,N_9678,N_11525);
nor U14166 (N_14166,N_8309,N_11738);
nor U14167 (N_14167,N_10593,N_10611);
nand U14168 (N_14168,N_11751,N_8639);
xor U14169 (N_14169,N_10669,N_10951);
nand U14170 (N_14170,N_11558,N_11089);
or U14171 (N_14171,N_8512,N_10662);
and U14172 (N_14172,N_10577,N_10624);
nand U14173 (N_14173,N_8812,N_11858);
and U14174 (N_14174,N_9958,N_11846);
nor U14175 (N_14175,N_11546,N_11079);
or U14176 (N_14176,N_9698,N_9958);
nand U14177 (N_14177,N_10693,N_11511);
nor U14178 (N_14178,N_11204,N_9118);
nor U14179 (N_14179,N_11449,N_10685);
nor U14180 (N_14180,N_11804,N_8105);
nor U14181 (N_14181,N_9733,N_9395);
and U14182 (N_14182,N_10785,N_10285);
and U14183 (N_14183,N_10979,N_8975);
xor U14184 (N_14184,N_10249,N_10226);
nor U14185 (N_14185,N_8013,N_9993);
nor U14186 (N_14186,N_11772,N_8449);
nand U14187 (N_14187,N_11154,N_9722);
xnor U14188 (N_14188,N_10441,N_11697);
or U14189 (N_14189,N_10852,N_9661);
and U14190 (N_14190,N_10440,N_10464);
and U14191 (N_14191,N_10623,N_9475);
nand U14192 (N_14192,N_10957,N_9213);
and U14193 (N_14193,N_8147,N_10631);
or U14194 (N_14194,N_10124,N_11469);
xnor U14195 (N_14195,N_11803,N_11790);
and U14196 (N_14196,N_11551,N_10554);
nor U14197 (N_14197,N_9367,N_8317);
xor U14198 (N_14198,N_9292,N_8536);
xnor U14199 (N_14199,N_10198,N_11909);
and U14200 (N_14200,N_9263,N_8780);
or U14201 (N_14201,N_10319,N_11353);
nand U14202 (N_14202,N_10564,N_11589);
or U14203 (N_14203,N_11527,N_11624);
or U14204 (N_14204,N_10727,N_11295);
nor U14205 (N_14205,N_8454,N_9138);
or U14206 (N_14206,N_9640,N_11195);
nand U14207 (N_14207,N_9094,N_9626);
xnor U14208 (N_14208,N_10743,N_9300);
xor U14209 (N_14209,N_9349,N_11801);
nand U14210 (N_14210,N_11074,N_9629);
nor U14211 (N_14211,N_8116,N_10725);
or U14212 (N_14212,N_11597,N_9668);
nor U14213 (N_14213,N_9799,N_11350);
nor U14214 (N_14214,N_11142,N_8572);
nand U14215 (N_14215,N_9506,N_9215);
nand U14216 (N_14216,N_9746,N_11096);
or U14217 (N_14217,N_9544,N_9258);
nor U14218 (N_14218,N_11294,N_11045);
xnor U14219 (N_14219,N_11531,N_10999);
nor U14220 (N_14220,N_10077,N_8946);
nand U14221 (N_14221,N_10341,N_10572);
or U14222 (N_14222,N_8330,N_11654);
and U14223 (N_14223,N_11891,N_8388);
nand U14224 (N_14224,N_8364,N_10932);
xnor U14225 (N_14225,N_10272,N_8920);
nand U14226 (N_14226,N_9611,N_10421);
nor U14227 (N_14227,N_9906,N_10809);
and U14228 (N_14228,N_10690,N_10857);
and U14229 (N_14229,N_11203,N_8868);
xnor U14230 (N_14230,N_10384,N_8154);
nand U14231 (N_14231,N_10251,N_9123);
nand U14232 (N_14232,N_10450,N_10945);
nor U14233 (N_14233,N_11839,N_8431);
nor U14234 (N_14234,N_10953,N_8698);
nand U14235 (N_14235,N_8396,N_9833);
nand U14236 (N_14236,N_10433,N_10951);
nand U14237 (N_14237,N_8902,N_11065);
or U14238 (N_14238,N_9158,N_8567);
xor U14239 (N_14239,N_9974,N_9215);
or U14240 (N_14240,N_11051,N_9138);
nand U14241 (N_14241,N_10407,N_10258);
and U14242 (N_14242,N_10067,N_9009);
nand U14243 (N_14243,N_10555,N_8503);
or U14244 (N_14244,N_8156,N_9595);
nand U14245 (N_14245,N_11073,N_11594);
and U14246 (N_14246,N_11038,N_8527);
nand U14247 (N_14247,N_8717,N_10832);
and U14248 (N_14248,N_11556,N_10181);
and U14249 (N_14249,N_10618,N_10821);
and U14250 (N_14250,N_9013,N_10814);
or U14251 (N_14251,N_11212,N_10028);
or U14252 (N_14252,N_8441,N_9530);
xor U14253 (N_14253,N_8762,N_8989);
or U14254 (N_14254,N_11143,N_11837);
and U14255 (N_14255,N_10392,N_8828);
nor U14256 (N_14256,N_9720,N_9386);
and U14257 (N_14257,N_8092,N_10671);
nor U14258 (N_14258,N_9781,N_10426);
and U14259 (N_14259,N_8021,N_10102);
or U14260 (N_14260,N_11390,N_10055);
and U14261 (N_14261,N_9786,N_9896);
and U14262 (N_14262,N_9653,N_11033);
nand U14263 (N_14263,N_9926,N_8768);
nand U14264 (N_14264,N_8841,N_8918);
xor U14265 (N_14265,N_11818,N_8076);
or U14266 (N_14266,N_10961,N_11084);
nor U14267 (N_14267,N_11185,N_11938);
nor U14268 (N_14268,N_9519,N_8551);
and U14269 (N_14269,N_10812,N_10187);
nand U14270 (N_14270,N_9205,N_11195);
nor U14271 (N_14271,N_10592,N_10310);
nand U14272 (N_14272,N_10579,N_8728);
nand U14273 (N_14273,N_11170,N_10781);
xnor U14274 (N_14274,N_8632,N_8675);
and U14275 (N_14275,N_10703,N_8584);
nand U14276 (N_14276,N_8536,N_11432);
nor U14277 (N_14277,N_10647,N_10806);
nor U14278 (N_14278,N_10467,N_11568);
nor U14279 (N_14279,N_10031,N_9102);
nor U14280 (N_14280,N_11367,N_9445);
or U14281 (N_14281,N_10140,N_9555);
and U14282 (N_14282,N_11265,N_9931);
nor U14283 (N_14283,N_11108,N_11026);
or U14284 (N_14284,N_8729,N_10208);
or U14285 (N_14285,N_10322,N_8022);
xor U14286 (N_14286,N_9173,N_11229);
or U14287 (N_14287,N_8372,N_11733);
nand U14288 (N_14288,N_10040,N_9603);
and U14289 (N_14289,N_11732,N_9207);
nor U14290 (N_14290,N_9571,N_10407);
nor U14291 (N_14291,N_9854,N_9882);
or U14292 (N_14292,N_11899,N_9105);
and U14293 (N_14293,N_8171,N_10977);
xor U14294 (N_14294,N_11965,N_9087);
and U14295 (N_14295,N_10676,N_11348);
nand U14296 (N_14296,N_9733,N_8371);
and U14297 (N_14297,N_8187,N_11234);
and U14298 (N_14298,N_10498,N_10153);
nor U14299 (N_14299,N_10851,N_10091);
xor U14300 (N_14300,N_9983,N_9443);
nor U14301 (N_14301,N_11215,N_8292);
or U14302 (N_14302,N_10880,N_8259);
or U14303 (N_14303,N_11607,N_11573);
xor U14304 (N_14304,N_9078,N_10486);
or U14305 (N_14305,N_8351,N_9428);
or U14306 (N_14306,N_10728,N_10004);
xor U14307 (N_14307,N_11355,N_9951);
nand U14308 (N_14308,N_8318,N_10530);
nand U14309 (N_14309,N_8212,N_8219);
and U14310 (N_14310,N_11398,N_8094);
nor U14311 (N_14311,N_9847,N_9929);
or U14312 (N_14312,N_10337,N_11271);
and U14313 (N_14313,N_11146,N_8003);
xnor U14314 (N_14314,N_11108,N_8969);
nor U14315 (N_14315,N_8154,N_11196);
or U14316 (N_14316,N_11958,N_11681);
nor U14317 (N_14317,N_9858,N_9047);
nor U14318 (N_14318,N_8546,N_10999);
and U14319 (N_14319,N_11491,N_10315);
xor U14320 (N_14320,N_10389,N_11059);
or U14321 (N_14321,N_8799,N_8095);
nor U14322 (N_14322,N_9104,N_9117);
nor U14323 (N_14323,N_11185,N_8878);
nand U14324 (N_14324,N_8118,N_8382);
and U14325 (N_14325,N_11969,N_11824);
or U14326 (N_14326,N_8549,N_8317);
nand U14327 (N_14327,N_10245,N_8424);
nand U14328 (N_14328,N_10648,N_11771);
nor U14329 (N_14329,N_10617,N_9157);
nor U14330 (N_14330,N_11304,N_11945);
and U14331 (N_14331,N_8457,N_8928);
nand U14332 (N_14332,N_11284,N_11331);
nor U14333 (N_14333,N_9821,N_8284);
nand U14334 (N_14334,N_10474,N_10944);
or U14335 (N_14335,N_10207,N_9109);
nand U14336 (N_14336,N_8426,N_8803);
nand U14337 (N_14337,N_10952,N_8073);
or U14338 (N_14338,N_10224,N_8616);
nand U14339 (N_14339,N_11349,N_9422);
xor U14340 (N_14340,N_10691,N_10720);
xnor U14341 (N_14341,N_9868,N_10081);
or U14342 (N_14342,N_10211,N_8068);
and U14343 (N_14343,N_9628,N_11891);
nor U14344 (N_14344,N_10781,N_9144);
nand U14345 (N_14345,N_11712,N_11957);
nand U14346 (N_14346,N_8893,N_9388);
and U14347 (N_14347,N_8386,N_11796);
xor U14348 (N_14348,N_8153,N_11960);
or U14349 (N_14349,N_11564,N_11403);
nor U14350 (N_14350,N_11880,N_10171);
nand U14351 (N_14351,N_8970,N_11108);
nand U14352 (N_14352,N_9993,N_8863);
nor U14353 (N_14353,N_10913,N_8113);
or U14354 (N_14354,N_9500,N_9808);
nand U14355 (N_14355,N_11220,N_11641);
nand U14356 (N_14356,N_10240,N_8192);
nand U14357 (N_14357,N_9311,N_9010);
nor U14358 (N_14358,N_9710,N_11661);
nor U14359 (N_14359,N_11021,N_8328);
or U14360 (N_14360,N_11290,N_9282);
nor U14361 (N_14361,N_10113,N_8855);
nand U14362 (N_14362,N_9914,N_8850);
or U14363 (N_14363,N_8548,N_11128);
xnor U14364 (N_14364,N_10179,N_9140);
and U14365 (N_14365,N_10894,N_9389);
and U14366 (N_14366,N_9803,N_10351);
nand U14367 (N_14367,N_9763,N_9434);
nor U14368 (N_14368,N_8375,N_9437);
and U14369 (N_14369,N_10753,N_11857);
or U14370 (N_14370,N_8417,N_10987);
or U14371 (N_14371,N_10490,N_9077);
nand U14372 (N_14372,N_10885,N_11340);
xnor U14373 (N_14373,N_10565,N_8590);
nand U14374 (N_14374,N_10854,N_8096);
and U14375 (N_14375,N_11421,N_10146);
and U14376 (N_14376,N_11419,N_10653);
and U14377 (N_14377,N_8444,N_9490);
nor U14378 (N_14378,N_8673,N_8233);
and U14379 (N_14379,N_11890,N_10641);
or U14380 (N_14380,N_9297,N_10727);
xor U14381 (N_14381,N_9352,N_11816);
or U14382 (N_14382,N_10098,N_10879);
or U14383 (N_14383,N_8405,N_11534);
and U14384 (N_14384,N_10986,N_11041);
or U14385 (N_14385,N_10918,N_10434);
nand U14386 (N_14386,N_9444,N_11555);
nor U14387 (N_14387,N_11104,N_9526);
nand U14388 (N_14388,N_9860,N_10071);
and U14389 (N_14389,N_9007,N_11953);
or U14390 (N_14390,N_11514,N_10423);
nand U14391 (N_14391,N_11766,N_8378);
xnor U14392 (N_14392,N_11453,N_9476);
or U14393 (N_14393,N_9736,N_9314);
nor U14394 (N_14394,N_11849,N_9284);
nor U14395 (N_14395,N_11139,N_11944);
nand U14396 (N_14396,N_8703,N_9947);
nor U14397 (N_14397,N_10602,N_10935);
nor U14398 (N_14398,N_8964,N_8051);
and U14399 (N_14399,N_8918,N_8413);
nand U14400 (N_14400,N_10203,N_10018);
nand U14401 (N_14401,N_10156,N_9875);
or U14402 (N_14402,N_11125,N_10712);
and U14403 (N_14403,N_9800,N_9690);
nor U14404 (N_14404,N_8133,N_11299);
nand U14405 (N_14405,N_8696,N_10425);
nand U14406 (N_14406,N_10621,N_11526);
or U14407 (N_14407,N_10055,N_8890);
or U14408 (N_14408,N_9961,N_8445);
nand U14409 (N_14409,N_11037,N_9765);
nor U14410 (N_14410,N_8331,N_10559);
or U14411 (N_14411,N_8414,N_8654);
or U14412 (N_14412,N_9230,N_11419);
nor U14413 (N_14413,N_11778,N_11733);
and U14414 (N_14414,N_8519,N_11170);
xnor U14415 (N_14415,N_10514,N_10885);
and U14416 (N_14416,N_8001,N_10172);
and U14417 (N_14417,N_9065,N_11171);
nor U14418 (N_14418,N_10355,N_9720);
and U14419 (N_14419,N_11633,N_9127);
nor U14420 (N_14420,N_8406,N_9981);
nor U14421 (N_14421,N_8062,N_11734);
and U14422 (N_14422,N_9637,N_11562);
nor U14423 (N_14423,N_10114,N_11065);
and U14424 (N_14424,N_9594,N_8697);
or U14425 (N_14425,N_10189,N_11781);
and U14426 (N_14426,N_9279,N_11441);
nor U14427 (N_14427,N_9563,N_8054);
nor U14428 (N_14428,N_9539,N_10611);
and U14429 (N_14429,N_10238,N_11171);
nor U14430 (N_14430,N_9415,N_9998);
nor U14431 (N_14431,N_10034,N_9836);
nand U14432 (N_14432,N_11470,N_9133);
or U14433 (N_14433,N_10022,N_10448);
or U14434 (N_14434,N_10541,N_10088);
and U14435 (N_14435,N_8682,N_10754);
nand U14436 (N_14436,N_9044,N_8691);
nand U14437 (N_14437,N_10131,N_11228);
and U14438 (N_14438,N_11052,N_10082);
nor U14439 (N_14439,N_11964,N_9055);
nor U14440 (N_14440,N_8069,N_8627);
nor U14441 (N_14441,N_9321,N_10760);
nor U14442 (N_14442,N_8961,N_10530);
nor U14443 (N_14443,N_9627,N_8318);
nor U14444 (N_14444,N_10667,N_9489);
and U14445 (N_14445,N_8365,N_10098);
nor U14446 (N_14446,N_8701,N_11161);
nor U14447 (N_14447,N_9064,N_8337);
and U14448 (N_14448,N_10723,N_10828);
or U14449 (N_14449,N_8988,N_8679);
and U14450 (N_14450,N_9827,N_8942);
and U14451 (N_14451,N_10396,N_11950);
nand U14452 (N_14452,N_11324,N_9351);
nor U14453 (N_14453,N_11304,N_11616);
nor U14454 (N_14454,N_11501,N_10233);
or U14455 (N_14455,N_9055,N_10985);
xnor U14456 (N_14456,N_10387,N_11901);
nand U14457 (N_14457,N_10727,N_11656);
nor U14458 (N_14458,N_10989,N_9846);
or U14459 (N_14459,N_10650,N_10472);
nand U14460 (N_14460,N_8177,N_9059);
or U14461 (N_14461,N_8424,N_9490);
nand U14462 (N_14462,N_10027,N_11931);
or U14463 (N_14463,N_11831,N_8293);
nand U14464 (N_14464,N_8496,N_8732);
or U14465 (N_14465,N_9645,N_11539);
or U14466 (N_14466,N_9453,N_9972);
and U14467 (N_14467,N_11285,N_9694);
nand U14468 (N_14468,N_9464,N_11125);
or U14469 (N_14469,N_10256,N_8328);
and U14470 (N_14470,N_11168,N_8796);
nand U14471 (N_14471,N_10313,N_9658);
and U14472 (N_14472,N_8309,N_10605);
and U14473 (N_14473,N_9391,N_11893);
nor U14474 (N_14474,N_9664,N_10575);
nand U14475 (N_14475,N_11093,N_11177);
and U14476 (N_14476,N_11730,N_8921);
or U14477 (N_14477,N_10394,N_8773);
xnor U14478 (N_14478,N_10655,N_8837);
nand U14479 (N_14479,N_9925,N_9378);
or U14480 (N_14480,N_9826,N_10428);
nor U14481 (N_14481,N_11066,N_9858);
xnor U14482 (N_14482,N_9445,N_8249);
nand U14483 (N_14483,N_11953,N_10218);
nor U14484 (N_14484,N_10403,N_9223);
nor U14485 (N_14485,N_10172,N_9886);
nand U14486 (N_14486,N_11304,N_11267);
and U14487 (N_14487,N_10653,N_9293);
or U14488 (N_14488,N_11690,N_10991);
xor U14489 (N_14489,N_10776,N_9763);
or U14490 (N_14490,N_9597,N_10312);
nand U14491 (N_14491,N_11615,N_11543);
nand U14492 (N_14492,N_8379,N_11351);
nand U14493 (N_14493,N_11051,N_10418);
nand U14494 (N_14494,N_9731,N_11074);
or U14495 (N_14495,N_9783,N_10397);
nand U14496 (N_14496,N_11535,N_11838);
and U14497 (N_14497,N_11585,N_9190);
nor U14498 (N_14498,N_10705,N_9933);
nor U14499 (N_14499,N_11122,N_11952);
nor U14500 (N_14500,N_10548,N_9428);
nor U14501 (N_14501,N_9769,N_11626);
and U14502 (N_14502,N_10739,N_9430);
nor U14503 (N_14503,N_8778,N_9759);
and U14504 (N_14504,N_10364,N_11845);
nor U14505 (N_14505,N_8824,N_8890);
or U14506 (N_14506,N_11851,N_8130);
nor U14507 (N_14507,N_11614,N_8404);
or U14508 (N_14508,N_10502,N_10317);
xnor U14509 (N_14509,N_10009,N_8753);
nor U14510 (N_14510,N_10545,N_11041);
nand U14511 (N_14511,N_11044,N_8952);
or U14512 (N_14512,N_9363,N_8801);
xor U14513 (N_14513,N_10391,N_11633);
nor U14514 (N_14514,N_10187,N_10512);
or U14515 (N_14515,N_10906,N_8965);
and U14516 (N_14516,N_8214,N_11480);
xnor U14517 (N_14517,N_11525,N_10420);
and U14518 (N_14518,N_9492,N_10729);
nand U14519 (N_14519,N_10545,N_8605);
nand U14520 (N_14520,N_11969,N_11737);
nor U14521 (N_14521,N_8103,N_11685);
and U14522 (N_14522,N_8722,N_10579);
nor U14523 (N_14523,N_11870,N_10856);
nor U14524 (N_14524,N_9478,N_8866);
and U14525 (N_14525,N_10661,N_10277);
or U14526 (N_14526,N_11469,N_9556);
or U14527 (N_14527,N_8167,N_10923);
nand U14528 (N_14528,N_11794,N_10058);
nor U14529 (N_14529,N_10841,N_11115);
and U14530 (N_14530,N_10586,N_11083);
or U14531 (N_14531,N_11964,N_11093);
nand U14532 (N_14532,N_8157,N_10180);
or U14533 (N_14533,N_10351,N_11984);
xnor U14534 (N_14534,N_10195,N_10843);
nor U14535 (N_14535,N_11708,N_10040);
xnor U14536 (N_14536,N_8716,N_10436);
nor U14537 (N_14537,N_10937,N_11006);
nor U14538 (N_14538,N_8512,N_9858);
and U14539 (N_14539,N_10733,N_10152);
and U14540 (N_14540,N_9138,N_8666);
nor U14541 (N_14541,N_10408,N_11677);
or U14542 (N_14542,N_10968,N_9147);
nand U14543 (N_14543,N_11316,N_8431);
or U14544 (N_14544,N_8862,N_10438);
nor U14545 (N_14545,N_8890,N_9365);
and U14546 (N_14546,N_11466,N_11318);
nor U14547 (N_14547,N_11344,N_10394);
or U14548 (N_14548,N_10840,N_11471);
and U14549 (N_14549,N_9446,N_11537);
nand U14550 (N_14550,N_8319,N_11880);
nor U14551 (N_14551,N_11133,N_11686);
xor U14552 (N_14552,N_11927,N_10190);
nand U14553 (N_14553,N_8830,N_8978);
or U14554 (N_14554,N_9422,N_10407);
nor U14555 (N_14555,N_10855,N_11058);
xor U14556 (N_14556,N_10011,N_9160);
nand U14557 (N_14557,N_11934,N_11150);
or U14558 (N_14558,N_10434,N_10105);
or U14559 (N_14559,N_11693,N_8305);
nor U14560 (N_14560,N_11808,N_8956);
and U14561 (N_14561,N_9750,N_9753);
and U14562 (N_14562,N_8645,N_11120);
or U14563 (N_14563,N_10248,N_10701);
nand U14564 (N_14564,N_10203,N_11437);
nand U14565 (N_14565,N_9125,N_8921);
nand U14566 (N_14566,N_9056,N_10878);
and U14567 (N_14567,N_9337,N_8168);
or U14568 (N_14568,N_10062,N_8640);
nor U14569 (N_14569,N_11911,N_10368);
or U14570 (N_14570,N_11664,N_8167);
and U14571 (N_14571,N_10941,N_8471);
or U14572 (N_14572,N_10855,N_8647);
nor U14573 (N_14573,N_11043,N_10124);
nor U14574 (N_14574,N_10719,N_8785);
or U14575 (N_14575,N_10149,N_9331);
nor U14576 (N_14576,N_9908,N_10762);
nor U14577 (N_14577,N_11278,N_10485);
nand U14578 (N_14578,N_9342,N_8456);
and U14579 (N_14579,N_8251,N_10840);
nor U14580 (N_14580,N_8098,N_9673);
or U14581 (N_14581,N_9528,N_11340);
nand U14582 (N_14582,N_10827,N_8735);
and U14583 (N_14583,N_8827,N_9436);
nor U14584 (N_14584,N_10606,N_9057);
nand U14585 (N_14585,N_11425,N_11813);
nor U14586 (N_14586,N_8038,N_8863);
and U14587 (N_14587,N_9998,N_10917);
xnor U14588 (N_14588,N_11658,N_8111);
and U14589 (N_14589,N_11137,N_10089);
and U14590 (N_14590,N_8279,N_11604);
nor U14591 (N_14591,N_11333,N_10789);
nand U14592 (N_14592,N_8549,N_8641);
and U14593 (N_14593,N_8914,N_9915);
or U14594 (N_14594,N_9966,N_10966);
xor U14595 (N_14595,N_11812,N_11469);
nor U14596 (N_14596,N_9844,N_8943);
nor U14597 (N_14597,N_9082,N_10264);
or U14598 (N_14598,N_10998,N_9822);
and U14599 (N_14599,N_11866,N_8717);
nand U14600 (N_14600,N_10922,N_8874);
or U14601 (N_14601,N_11932,N_11217);
nor U14602 (N_14602,N_11610,N_8198);
and U14603 (N_14603,N_10797,N_9454);
and U14604 (N_14604,N_8048,N_8307);
nor U14605 (N_14605,N_11592,N_9288);
or U14606 (N_14606,N_11652,N_11670);
and U14607 (N_14607,N_11959,N_9968);
nor U14608 (N_14608,N_9710,N_8488);
or U14609 (N_14609,N_9315,N_8009);
and U14610 (N_14610,N_11555,N_11795);
nor U14611 (N_14611,N_11680,N_11639);
and U14612 (N_14612,N_11376,N_11041);
and U14613 (N_14613,N_10762,N_11814);
xnor U14614 (N_14614,N_10920,N_8333);
or U14615 (N_14615,N_8495,N_10989);
and U14616 (N_14616,N_11473,N_10389);
nand U14617 (N_14617,N_8767,N_9017);
or U14618 (N_14618,N_10066,N_8865);
or U14619 (N_14619,N_8673,N_11811);
nand U14620 (N_14620,N_10671,N_9642);
xor U14621 (N_14621,N_8001,N_9677);
nand U14622 (N_14622,N_8586,N_10658);
nand U14623 (N_14623,N_10354,N_10435);
and U14624 (N_14624,N_9270,N_11820);
nand U14625 (N_14625,N_10894,N_9812);
or U14626 (N_14626,N_10259,N_9779);
nor U14627 (N_14627,N_9734,N_11995);
and U14628 (N_14628,N_8642,N_10729);
nor U14629 (N_14629,N_11443,N_9980);
nand U14630 (N_14630,N_11978,N_8667);
xor U14631 (N_14631,N_10438,N_9066);
nor U14632 (N_14632,N_8365,N_9772);
nand U14633 (N_14633,N_9308,N_11171);
and U14634 (N_14634,N_9150,N_10292);
nand U14635 (N_14635,N_9190,N_8244);
xnor U14636 (N_14636,N_10668,N_8706);
or U14637 (N_14637,N_9413,N_8961);
or U14638 (N_14638,N_8882,N_9936);
nand U14639 (N_14639,N_10612,N_11591);
or U14640 (N_14640,N_9483,N_10668);
nor U14641 (N_14641,N_8507,N_11516);
nand U14642 (N_14642,N_10848,N_10136);
and U14643 (N_14643,N_9572,N_8244);
xor U14644 (N_14644,N_10973,N_10150);
nor U14645 (N_14645,N_11917,N_8031);
nor U14646 (N_14646,N_10176,N_9411);
and U14647 (N_14647,N_11903,N_11070);
xnor U14648 (N_14648,N_11486,N_8815);
nand U14649 (N_14649,N_9472,N_9109);
or U14650 (N_14650,N_10938,N_10930);
nand U14651 (N_14651,N_9085,N_10652);
or U14652 (N_14652,N_8271,N_11166);
nor U14653 (N_14653,N_8085,N_10589);
nand U14654 (N_14654,N_11828,N_9521);
nand U14655 (N_14655,N_8004,N_11391);
nand U14656 (N_14656,N_10024,N_9069);
and U14657 (N_14657,N_9788,N_9804);
nand U14658 (N_14658,N_9011,N_11369);
and U14659 (N_14659,N_9168,N_10801);
nand U14660 (N_14660,N_8051,N_9958);
or U14661 (N_14661,N_8036,N_10682);
nor U14662 (N_14662,N_11698,N_10945);
or U14663 (N_14663,N_10835,N_11291);
nand U14664 (N_14664,N_8928,N_9732);
or U14665 (N_14665,N_11812,N_10249);
nand U14666 (N_14666,N_8645,N_9399);
nor U14667 (N_14667,N_8949,N_8258);
nand U14668 (N_14668,N_11183,N_11157);
nand U14669 (N_14669,N_9475,N_11291);
or U14670 (N_14670,N_11913,N_11757);
or U14671 (N_14671,N_8058,N_11690);
and U14672 (N_14672,N_8518,N_10876);
and U14673 (N_14673,N_9305,N_10799);
or U14674 (N_14674,N_10219,N_11369);
nand U14675 (N_14675,N_11467,N_10399);
or U14676 (N_14676,N_9818,N_8330);
nand U14677 (N_14677,N_9935,N_10237);
or U14678 (N_14678,N_8065,N_8528);
nand U14679 (N_14679,N_8059,N_9177);
or U14680 (N_14680,N_11532,N_8428);
and U14681 (N_14681,N_10241,N_8908);
and U14682 (N_14682,N_9878,N_10691);
or U14683 (N_14683,N_10918,N_11163);
nand U14684 (N_14684,N_8948,N_8384);
and U14685 (N_14685,N_8182,N_11804);
nor U14686 (N_14686,N_9724,N_11572);
xnor U14687 (N_14687,N_10065,N_11644);
nor U14688 (N_14688,N_9791,N_8913);
or U14689 (N_14689,N_11097,N_8492);
nor U14690 (N_14690,N_10998,N_10541);
and U14691 (N_14691,N_8428,N_8487);
nand U14692 (N_14692,N_11604,N_10680);
or U14693 (N_14693,N_11046,N_8645);
or U14694 (N_14694,N_10655,N_10680);
and U14695 (N_14695,N_11099,N_10176);
and U14696 (N_14696,N_8764,N_9150);
nand U14697 (N_14697,N_11536,N_11666);
nand U14698 (N_14698,N_8035,N_11790);
and U14699 (N_14699,N_9476,N_9843);
and U14700 (N_14700,N_10355,N_11386);
or U14701 (N_14701,N_9026,N_9200);
nor U14702 (N_14702,N_9609,N_9556);
nand U14703 (N_14703,N_11611,N_8863);
nand U14704 (N_14704,N_10804,N_11072);
xnor U14705 (N_14705,N_9101,N_11332);
xnor U14706 (N_14706,N_9300,N_8521);
nor U14707 (N_14707,N_9522,N_10984);
nand U14708 (N_14708,N_11942,N_9011);
nand U14709 (N_14709,N_9037,N_11235);
and U14710 (N_14710,N_8798,N_9207);
or U14711 (N_14711,N_10145,N_10218);
and U14712 (N_14712,N_10486,N_9097);
nand U14713 (N_14713,N_8935,N_11632);
and U14714 (N_14714,N_10726,N_10465);
and U14715 (N_14715,N_9756,N_10694);
xnor U14716 (N_14716,N_11512,N_10592);
and U14717 (N_14717,N_11464,N_8614);
nor U14718 (N_14718,N_9568,N_11039);
nand U14719 (N_14719,N_9844,N_10218);
nor U14720 (N_14720,N_11867,N_11524);
nor U14721 (N_14721,N_8544,N_11438);
nand U14722 (N_14722,N_10852,N_9667);
nor U14723 (N_14723,N_8974,N_11452);
or U14724 (N_14724,N_11585,N_9716);
or U14725 (N_14725,N_8105,N_11467);
nand U14726 (N_14726,N_8760,N_10799);
or U14727 (N_14727,N_8297,N_11264);
or U14728 (N_14728,N_8854,N_11730);
and U14729 (N_14729,N_8044,N_8818);
nand U14730 (N_14730,N_9485,N_8995);
nand U14731 (N_14731,N_9360,N_8584);
or U14732 (N_14732,N_8131,N_8616);
or U14733 (N_14733,N_10215,N_8354);
and U14734 (N_14734,N_9265,N_9805);
or U14735 (N_14735,N_10678,N_8784);
nand U14736 (N_14736,N_11289,N_10188);
and U14737 (N_14737,N_8579,N_9741);
nor U14738 (N_14738,N_8384,N_9038);
nor U14739 (N_14739,N_10431,N_10219);
and U14740 (N_14740,N_9941,N_11585);
and U14741 (N_14741,N_10384,N_9701);
nor U14742 (N_14742,N_8909,N_10497);
nand U14743 (N_14743,N_10586,N_11488);
nand U14744 (N_14744,N_11006,N_10085);
or U14745 (N_14745,N_10938,N_11213);
and U14746 (N_14746,N_11204,N_10985);
nor U14747 (N_14747,N_11191,N_9105);
or U14748 (N_14748,N_11639,N_8542);
nor U14749 (N_14749,N_8719,N_11915);
and U14750 (N_14750,N_11683,N_9872);
xor U14751 (N_14751,N_11120,N_9495);
and U14752 (N_14752,N_10525,N_11864);
and U14753 (N_14753,N_10003,N_8038);
nor U14754 (N_14754,N_8124,N_11483);
xnor U14755 (N_14755,N_11552,N_10635);
and U14756 (N_14756,N_10559,N_10041);
nor U14757 (N_14757,N_8343,N_9153);
or U14758 (N_14758,N_10987,N_10842);
or U14759 (N_14759,N_8553,N_9614);
or U14760 (N_14760,N_10759,N_11821);
nor U14761 (N_14761,N_9639,N_10791);
or U14762 (N_14762,N_8874,N_9647);
nand U14763 (N_14763,N_9160,N_8132);
nor U14764 (N_14764,N_9233,N_11453);
nor U14765 (N_14765,N_9563,N_10032);
or U14766 (N_14766,N_11234,N_11370);
and U14767 (N_14767,N_10895,N_8347);
nand U14768 (N_14768,N_10831,N_9501);
and U14769 (N_14769,N_9860,N_10539);
or U14770 (N_14770,N_9842,N_10415);
or U14771 (N_14771,N_11942,N_10946);
or U14772 (N_14772,N_11304,N_11919);
nor U14773 (N_14773,N_10385,N_9920);
and U14774 (N_14774,N_9893,N_9326);
and U14775 (N_14775,N_8024,N_10350);
nand U14776 (N_14776,N_8846,N_9250);
xor U14777 (N_14777,N_11012,N_11523);
nand U14778 (N_14778,N_10938,N_10907);
nand U14779 (N_14779,N_8451,N_11236);
or U14780 (N_14780,N_8175,N_10108);
nor U14781 (N_14781,N_8717,N_8412);
and U14782 (N_14782,N_11916,N_8567);
or U14783 (N_14783,N_9419,N_10948);
nand U14784 (N_14784,N_8141,N_8733);
nand U14785 (N_14785,N_10911,N_11098);
and U14786 (N_14786,N_9361,N_8292);
and U14787 (N_14787,N_8493,N_11990);
or U14788 (N_14788,N_11329,N_11593);
or U14789 (N_14789,N_9082,N_11285);
nand U14790 (N_14790,N_11346,N_8421);
or U14791 (N_14791,N_11336,N_11230);
and U14792 (N_14792,N_11059,N_10606);
and U14793 (N_14793,N_8184,N_10068);
nand U14794 (N_14794,N_8572,N_11259);
or U14795 (N_14795,N_8620,N_8551);
and U14796 (N_14796,N_10707,N_8627);
xnor U14797 (N_14797,N_10955,N_9946);
nor U14798 (N_14798,N_10518,N_8402);
xor U14799 (N_14799,N_9885,N_8264);
nor U14800 (N_14800,N_9950,N_11042);
xor U14801 (N_14801,N_11041,N_11691);
xor U14802 (N_14802,N_10385,N_11230);
and U14803 (N_14803,N_10185,N_10985);
and U14804 (N_14804,N_9687,N_10746);
xor U14805 (N_14805,N_9376,N_8481);
xnor U14806 (N_14806,N_9622,N_8652);
nand U14807 (N_14807,N_10523,N_10980);
nor U14808 (N_14808,N_10094,N_9351);
nor U14809 (N_14809,N_9985,N_10284);
nand U14810 (N_14810,N_9413,N_8688);
nand U14811 (N_14811,N_10493,N_8708);
and U14812 (N_14812,N_8327,N_8824);
and U14813 (N_14813,N_9258,N_10911);
xor U14814 (N_14814,N_10909,N_10656);
xnor U14815 (N_14815,N_8178,N_11192);
and U14816 (N_14816,N_9502,N_10547);
or U14817 (N_14817,N_8174,N_8760);
nand U14818 (N_14818,N_10041,N_8168);
or U14819 (N_14819,N_9413,N_10607);
or U14820 (N_14820,N_10636,N_10087);
nor U14821 (N_14821,N_8145,N_10596);
or U14822 (N_14822,N_11668,N_8549);
and U14823 (N_14823,N_10273,N_8751);
nand U14824 (N_14824,N_11295,N_11031);
nand U14825 (N_14825,N_9499,N_10800);
nand U14826 (N_14826,N_10360,N_11321);
nor U14827 (N_14827,N_10271,N_8729);
or U14828 (N_14828,N_10694,N_9579);
or U14829 (N_14829,N_9166,N_8008);
and U14830 (N_14830,N_8015,N_8711);
nand U14831 (N_14831,N_8587,N_9590);
nand U14832 (N_14832,N_8320,N_9147);
or U14833 (N_14833,N_10370,N_11757);
or U14834 (N_14834,N_10384,N_10853);
and U14835 (N_14835,N_11925,N_8363);
and U14836 (N_14836,N_8189,N_9721);
or U14837 (N_14837,N_10787,N_11940);
and U14838 (N_14838,N_10021,N_8516);
nand U14839 (N_14839,N_10865,N_11693);
nor U14840 (N_14840,N_8336,N_8410);
nand U14841 (N_14841,N_9641,N_8840);
and U14842 (N_14842,N_10226,N_10287);
nor U14843 (N_14843,N_8700,N_11553);
nor U14844 (N_14844,N_11547,N_11261);
xnor U14845 (N_14845,N_10823,N_10374);
or U14846 (N_14846,N_10367,N_10477);
nand U14847 (N_14847,N_8189,N_8615);
nor U14848 (N_14848,N_10713,N_9652);
or U14849 (N_14849,N_11959,N_11953);
nand U14850 (N_14850,N_11091,N_11173);
or U14851 (N_14851,N_8000,N_11684);
nor U14852 (N_14852,N_11698,N_8264);
nor U14853 (N_14853,N_11604,N_8291);
and U14854 (N_14854,N_9701,N_9217);
nand U14855 (N_14855,N_10840,N_10699);
or U14856 (N_14856,N_10574,N_10007);
or U14857 (N_14857,N_10581,N_8111);
nand U14858 (N_14858,N_9246,N_10834);
nand U14859 (N_14859,N_9013,N_11709);
nor U14860 (N_14860,N_10040,N_10650);
nand U14861 (N_14861,N_8409,N_11425);
or U14862 (N_14862,N_10534,N_9861);
xnor U14863 (N_14863,N_10643,N_9191);
xor U14864 (N_14864,N_8676,N_8174);
nor U14865 (N_14865,N_8623,N_8704);
nand U14866 (N_14866,N_11829,N_11646);
nand U14867 (N_14867,N_9533,N_11705);
nand U14868 (N_14868,N_9714,N_9480);
xnor U14869 (N_14869,N_11358,N_9440);
xnor U14870 (N_14870,N_8153,N_10917);
xnor U14871 (N_14871,N_11795,N_9332);
xor U14872 (N_14872,N_10996,N_10003);
and U14873 (N_14873,N_11902,N_8045);
or U14874 (N_14874,N_10408,N_10785);
or U14875 (N_14875,N_10639,N_8891);
xor U14876 (N_14876,N_11750,N_10046);
or U14877 (N_14877,N_10922,N_8189);
or U14878 (N_14878,N_9586,N_8250);
nand U14879 (N_14879,N_10327,N_10765);
nand U14880 (N_14880,N_8588,N_10687);
nand U14881 (N_14881,N_9159,N_11117);
and U14882 (N_14882,N_9269,N_9631);
xor U14883 (N_14883,N_11785,N_9804);
and U14884 (N_14884,N_8378,N_8046);
nor U14885 (N_14885,N_10474,N_10669);
or U14886 (N_14886,N_11543,N_8821);
and U14887 (N_14887,N_10457,N_8131);
and U14888 (N_14888,N_8017,N_8679);
nand U14889 (N_14889,N_11148,N_11234);
and U14890 (N_14890,N_10612,N_10674);
nand U14891 (N_14891,N_9777,N_11492);
nand U14892 (N_14892,N_8811,N_9553);
nand U14893 (N_14893,N_9051,N_9654);
nand U14894 (N_14894,N_11096,N_9660);
or U14895 (N_14895,N_9042,N_10618);
and U14896 (N_14896,N_8659,N_11939);
nand U14897 (N_14897,N_10997,N_8963);
or U14898 (N_14898,N_8566,N_10885);
nor U14899 (N_14899,N_9768,N_10962);
nand U14900 (N_14900,N_10678,N_8126);
and U14901 (N_14901,N_11343,N_8883);
nand U14902 (N_14902,N_8204,N_10665);
nor U14903 (N_14903,N_8858,N_10871);
and U14904 (N_14904,N_8296,N_9465);
xor U14905 (N_14905,N_9613,N_8256);
and U14906 (N_14906,N_11981,N_9391);
nand U14907 (N_14907,N_9040,N_8962);
nand U14908 (N_14908,N_9595,N_10037);
xor U14909 (N_14909,N_8720,N_11665);
nand U14910 (N_14910,N_11306,N_10206);
nor U14911 (N_14911,N_9224,N_10653);
nand U14912 (N_14912,N_11483,N_10480);
nor U14913 (N_14913,N_11179,N_11632);
and U14914 (N_14914,N_9662,N_9387);
nor U14915 (N_14915,N_8643,N_8228);
or U14916 (N_14916,N_8582,N_11796);
nand U14917 (N_14917,N_11251,N_8461);
nor U14918 (N_14918,N_8198,N_10854);
and U14919 (N_14919,N_10967,N_10671);
xor U14920 (N_14920,N_9824,N_10751);
and U14921 (N_14921,N_10777,N_11811);
xnor U14922 (N_14922,N_11051,N_10581);
nor U14923 (N_14923,N_9616,N_9179);
and U14924 (N_14924,N_9861,N_9953);
nor U14925 (N_14925,N_11951,N_8700);
nand U14926 (N_14926,N_10219,N_11245);
or U14927 (N_14927,N_11488,N_8617);
nand U14928 (N_14928,N_8327,N_10034);
or U14929 (N_14929,N_8044,N_11477);
or U14930 (N_14930,N_10322,N_11214);
nand U14931 (N_14931,N_9120,N_9063);
or U14932 (N_14932,N_11182,N_10673);
xnor U14933 (N_14933,N_9472,N_9378);
nor U14934 (N_14934,N_9840,N_10088);
nand U14935 (N_14935,N_8559,N_9618);
nand U14936 (N_14936,N_10155,N_10147);
and U14937 (N_14937,N_8447,N_11000);
xor U14938 (N_14938,N_11389,N_11501);
nor U14939 (N_14939,N_10956,N_10431);
or U14940 (N_14940,N_11693,N_8129);
and U14941 (N_14941,N_9733,N_8781);
nor U14942 (N_14942,N_10999,N_10651);
nand U14943 (N_14943,N_11371,N_11996);
and U14944 (N_14944,N_11996,N_8140);
nor U14945 (N_14945,N_10699,N_9252);
nand U14946 (N_14946,N_8943,N_11664);
nand U14947 (N_14947,N_8765,N_11320);
and U14948 (N_14948,N_9048,N_8100);
nor U14949 (N_14949,N_11375,N_10373);
nor U14950 (N_14950,N_8697,N_11322);
nor U14951 (N_14951,N_11297,N_11098);
nand U14952 (N_14952,N_11662,N_10757);
nand U14953 (N_14953,N_10564,N_8545);
and U14954 (N_14954,N_10013,N_8335);
nand U14955 (N_14955,N_11594,N_10605);
or U14956 (N_14956,N_10021,N_8205);
nand U14957 (N_14957,N_8793,N_9043);
nand U14958 (N_14958,N_11040,N_9639);
or U14959 (N_14959,N_10953,N_8944);
and U14960 (N_14960,N_8487,N_10931);
or U14961 (N_14961,N_11431,N_11054);
and U14962 (N_14962,N_8394,N_8905);
or U14963 (N_14963,N_11909,N_10613);
nand U14964 (N_14964,N_9307,N_8989);
nand U14965 (N_14965,N_8185,N_9072);
or U14966 (N_14966,N_9643,N_11506);
nand U14967 (N_14967,N_8310,N_11122);
xnor U14968 (N_14968,N_9831,N_8797);
and U14969 (N_14969,N_9459,N_9667);
and U14970 (N_14970,N_11053,N_8184);
and U14971 (N_14971,N_9471,N_11568);
nand U14972 (N_14972,N_11193,N_8076);
or U14973 (N_14973,N_9216,N_9815);
or U14974 (N_14974,N_11175,N_11297);
or U14975 (N_14975,N_10892,N_8920);
and U14976 (N_14976,N_8500,N_8901);
nor U14977 (N_14977,N_9365,N_9354);
nor U14978 (N_14978,N_11737,N_9827);
xnor U14979 (N_14979,N_10805,N_9329);
xor U14980 (N_14980,N_11382,N_9875);
nor U14981 (N_14981,N_8992,N_9740);
xor U14982 (N_14982,N_11370,N_10796);
xnor U14983 (N_14983,N_8411,N_11890);
nor U14984 (N_14984,N_11624,N_9981);
nor U14985 (N_14985,N_11684,N_11467);
and U14986 (N_14986,N_9637,N_10020);
nand U14987 (N_14987,N_9750,N_9430);
xor U14988 (N_14988,N_10538,N_9198);
or U14989 (N_14989,N_8617,N_8768);
nor U14990 (N_14990,N_9019,N_10996);
nand U14991 (N_14991,N_10958,N_10389);
xor U14992 (N_14992,N_10834,N_10360);
or U14993 (N_14993,N_9099,N_8825);
nor U14994 (N_14994,N_10582,N_10622);
nor U14995 (N_14995,N_9557,N_11687);
and U14996 (N_14996,N_10182,N_10143);
nor U14997 (N_14997,N_8491,N_11417);
nor U14998 (N_14998,N_8438,N_9758);
and U14999 (N_14999,N_8215,N_8727);
nand U15000 (N_15000,N_9111,N_11345);
xnor U15001 (N_15001,N_10729,N_11103);
nor U15002 (N_15002,N_8635,N_8010);
xor U15003 (N_15003,N_11865,N_9938);
xnor U15004 (N_15004,N_8964,N_9735);
nand U15005 (N_15005,N_9869,N_10130);
nand U15006 (N_15006,N_8278,N_8784);
and U15007 (N_15007,N_11381,N_8227);
or U15008 (N_15008,N_8634,N_11995);
or U15009 (N_15009,N_9441,N_9315);
and U15010 (N_15010,N_9161,N_9945);
nor U15011 (N_15011,N_10163,N_8218);
or U15012 (N_15012,N_10772,N_11297);
or U15013 (N_15013,N_9344,N_11592);
nand U15014 (N_15014,N_9260,N_9002);
nor U15015 (N_15015,N_10388,N_10994);
nor U15016 (N_15016,N_8423,N_9474);
and U15017 (N_15017,N_10877,N_8103);
nor U15018 (N_15018,N_9989,N_8807);
nor U15019 (N_15019,N_11754,N_8336);
nor U15020 (N_15020,N_8053,N_10492);
nand U15021 (N_15021,N_10031,N_8603);
and U15022 (N_15022,N_9038,N_11456);
and U15023 (N_15023,N_8777,N_11104);
or U15024 (N_15024,N_8307,N_8523);
or U15025 (N_15025,N_10138,N_11669);
xor U15026 (N_15026,N_11600,N_9116);
and U15027 (N_15027,N_10725,N_11567);
or U15028 (N_15028,N_11149,N_11302);
or U15029 (N_15029,N_9508,N_10924);
nor U15030 (N_15030,N_10807,N_9008);
nand U15031 (N_15031,N_11546,N_8643);
nor U15032 (N_15032,N_9901,N_11800);
and U15033 (N_15033,N_9518,N_8807);
nor U15034 (N_15034,N_8361,N_8471);
nor U15035 (N_15035,N_10548,N_8690);
nor U15036 (N_15036,N_8941,N_10379);
nand U15037 (N_15037,N_11382,N_10709);
nor U15038 (N_15038,N_8545,N_9998);
and U15039 (N_15039,N_10621,N_9674);
or U15040 (N_15040,N_9124,N_10422);
nor U15041 (N_15041,N_10618,N_11684);
xnor U15042 (N_15042,N_8888,N_11927);
and U15043 (N_15043,N_9639,N_11251);
xnor U15044 (N_15044,N_9211,N_10057);
nor U15045 (N_15045,N_10406,N_8080);
or U15046 (N_15046,N_9858,N_11316);
or U15047 (N_15047,N_11558,N_11475);
nor U15048 (N_15048,N_8256,N_8981);
nand U15049 (N_15049,N_11034,N_9693);
nand U15050 (N_15050,N_9684,N_11622);
nand U15051 (N_15051,N_11767,N_10275);
xor U15052 (N_15052,N_10385,N_10888);
or U15053 (N_15053,N_10913,N_9949);
or U15054 (N_15054,N_9182,N_8958);
or U15055 (N_15055,N_9873,N_8468);
and U15056 (N_15056,N_9851,N_11642);
nor U15057 (N_15057,N_10147,N_11204);
and U15058 (N_15058,N_11334,N_10083);
nor U15059 (N_15059,N_8584,N_10280);
and U15060 (N_15060,N_8657,N_11536);
nor U15061 (N_15061,N_11360,N_8462);
and U15062 (N_15062,N_11752,N_9952);
and U15063 (N_15063,N_11427,N_10889);
or U15064 (N_15064,N_8415,N_9298);
nor U15065 (N_15065,N_11024,N_9269);
and U15066 (N_15066,N_8036,N_11652);
nor U15067 (N_15067,N_10523,N_9797);
xor U15068 (N_15068,N_9087,N_9905);
nand U15069 (N_15069,N_8658,N_10414);
xnor U15070 (N_15070,N_10309,N_8408);
or U15071 (N_15071,N_9209,N_10600);
and U15072 (N_15072,N_9040,N_8797);
nor U15073 (N_15073,N_11935,N_10711);
xor U15074 (N_15074,N_9462,N_11580);
or U15075 (N_15075,N_11391,N_9089);
nand U15076 (N_15076,N_8980,N_11885);
and U15077 (N_15077,N_8962,N_8845);
and U15078 (N_15078,N_8861,N_11507);
nor U15079 (N_15079,N_11781,N_8937);
nor U15080 (N_15080,N_9060,N_10814);
nand U15081 (N_15081,N_11073,N_8257);
nor U15082 (N_15082,N_11291,N_8747);
and U15083 (N_15083,N_8625,N_9759);
nand U15084 (N_15084,N_9320,N_8259);
and U15085 (N_15085,N_9239,N_9876);
nand U15086 (N_15086,N_9666,N_11521);
nor U15087 (N_15087,N_11046,N_9961);
nor U15088 (N_15088,N_9396,N_10008);
nor U15089 (N_15089,N_11177,N_11370);
and U15090 (N_15090,N_9033,N_11610);
nand U15091 (N_15091,N_8078,N_11506);
or U15092 (N_15092,N_11030,N_8423);
nand U15093 (N_15093,N_9095,N_8741);
and U15094 (N_15094,N_11078,N_9612);
or U15095 (N_15095,N_10997,N_8534);
and U15096 (N_15096,N_8230,N_8724);
nand U15097 (N_15097,N_8951,N_11042);
and U15098 (N_15098,N_9530,N_11827);
nand U15099 (N_15099,N_10615,N_10723);
nand U15100 (N_15100,N_11185,N_11752);
nand U15101 (N_15101,N_10517,N_9118);
nor U15102 (N_15102,N_8842,N_10058);
or U15103 (N_15103,N_10183,N_9012);
nand U15104 (N_15104,N_8741,N_10708);
or U15105 (N_15105,N_9325,N_9681);
or U15106 (N_15106,N_11819,N_11658);
nor U15107 (N_15107,N_11695,N_10270);
nand U15108 (N_15108,N_9972,N_8176);
nand U15109 (N_15109,N_11159,N_8567);
nor U15110 (N_15110,N_8417,N_8586);
nand U15111 (N_15111,N_8334,N_9858);
and U15112 (N_15112,N_8624,N_8861);
nand U15113 (N_15113,N_10162,N_10310);
or U15114 (N_15114,N_10885,N_9754);
xnor U15115 (N_15115,N_11486,N_11654);
xor U15116 (N_15116,N_11555,N_10820);
nand U15117 (N_15117,N_10044,N_8596);
or U15118 (N_15118,N_10800,N_10152);
or U15119 (N_15119,N_10633,N_8115);
xor U15120 (N_15120,N_8143,N_10264);
or U15121 (N_15121,N_8079,N_10013);
nor U15122 (N_15122,N_9712,N_9608);
nor U15123 (N_15123,N_9866,N_8722);
nor U15124 (N_15124,N_11994,N_8558);
and U15125 (N_15125,N_10266,N_8184);
or U15126 (N_15126,N_9471,N_9268);
nand U15127 (N_15127,N_8460,N_10493);
nand U15128 (N_15128,N_9288,N_11080);
and U15129 (N_15129,N_8220,N_10885);
nor U15130 (N_15130,N_9540,N_11121);
xor U15131 (N_15131,N_9436,N_11110);
nor U15132 (N_15132,N_11096,N_9433);
nor U15133 (N_15133,N_11778,N_9633);
or U15134 (N_15134,N_8332,N_10481);
and U15135 (N_15135,N_11754,N_9782);
and U15136 (N_15136,N_11783,N_9592);
nand U15137 (N_15137,N_11936,N_10946);
nand U15138 (N_15138,N_11166,N_9493);
or U15139 (N_15139,N_11906,N_9209);
nand U15140 (N_15140,N_11371,N_10709);
and U15141 (N_15141,N_9646,N_8946);
nor U15142 (N_15142,N_9867,N_11209);
nand U15143 (N_15143,N_9925,N_10970);
xnor U15144 (N_15144,N_8318,N_8233);
and U15145 (N_15145,N_10886,N_8777);
nand U15146 (N_15146,N_8089,N_8563);
nor U15147 (N_15147,N_8185,N_8828);
nor U15148 (N_15148,N_9671,N_11878);
nor U15149 (N_15149,N_10511,N_8742);
nor U15150 (N_15150,N_9560,N_9158);
nor U15151 (N_15151,N_11925,N_10834);
or U15152 (N_15152,N_9193,N_10575);
or U15153 (N_15153,N_8597,N_8847);
nor U15154 (N_15154,N_8577,N_10103);
or U15155 (N_15155,N_8910,N_11740);
nand U15156 (N_15156,N_8588,N_9977);
nor U15157 (N_15157,N_10826,N_10718);
or U15158 (N_15158,N_11601,N_8721);
nand U15159 (N_15159,N_8897,N_11917);
nand U15160 (N_15160,N_8738,N_9275);
or U15161 (N_15161,N_11785,N_9529);
nor U15162 (N_15162,N_10122,N_9590);
or U15163 (N_15163,N_9551,N_11989);
nor U15164 (N_15164,N_10441,N_9501);
and U15165 (N_15165,N_9799,N_8660);
nor U15166 (N_15166,N_11688,N_9230);
and U15167 (N_15167,N_9342,N_11605);
nand U15168 (N_15168,N_8847,N_11158);
or U15169 (N_15169,N_11111,N_11596);
or U15170 (N_15170,N_9948,N_11180);
nor U15171 (N_15171,N_10251,N_8718);
nor U15172 (N_15172,N_10353,N_9457);
nand U15173 (N_15173,N_11387,N_11825);
nand U15174 (N_15174,N_11231,N_8335);
nor U15175 (N_15175,N_11010,N_11652);
nor U15176 (N_15176,N_11127,N_9280);
xor U15177 (N_15177,N_10888,N_9455);
and U15178 (N_15178,N_8738,N_10009);
and U15179 (N_15179,N_9438,N_11706);
and U15180 (N_15180,N_8916,N_9860);
nand U15181 (N_15181,N_11317,N_9866);
nor U15182 (N_15182,N_10651,N_10962);
and U15183 (N_15183,N_8604,N_9447);
xnor U15184 (N_15184,N_11784,N_9795);
nor U15185 (N_15185,N_10202,N_10220);
or U15186 (N_15186,N_10583,N_9525);
and U15187 (N_15187,N_8883,N_9811);
or U15188 (N_15188,N_10161,N_9294);
nor U15189 (N_15189,N_8031,N_8476);
or U15190 (N_15190,N_11727,N_10233);
or U15191 (N_15191,N_9146,N_10188);
and U15192 (N_15192,N_10353,N_8239);
nor U15193 (N_15193,N_10409,N_10341);
nor U15194 (N_15194,N_10787,N_10398);
and U15195 (N_15195,N_9697,N_11842);
nor U15196 (N_15196,N_10024,N_10258);
and U15197 (N_15197,N_11384,N_9620);
or U15198 (N_15198,N_9297,N_8923);
and U15199 (N_15199,N_10832,N_11957);
or U15200 (N_15200,N_8901,N_8529);
xnor U15201 (N_15201,N_11105,N_8196);
xor U15202 (N_15202,N_11959,N_8503);
nor U15203 (N_15203,N_10961,N_8310);
or U15204 (N_15204,N_9581,N_11192);
nor U15205 (N_15205,N_8901,N_11095);
xnor U15206 (N_15206,N_9907,N_10017);
nand U15207 (N_15207,N_11729,N_9065);
nand U15208 (N_15208,N_8528,N_9771);
xor U15209 (N_15209,N_10466,N_11691);
or U15210 (N_15210,N_9437,N_10739);
nor U15211 (N_15211,N_9114,N_8392);
and U15212 (N_15212,N_10874,N_8237);
or U15213 (N_15213,N_10928,N_8719);
and U15214 (N_15214,N_9118,N_9019);
and U15215 (N_15215,N_9605,N_9566);
or U15216 (N_15216,N_9359,N_8886);
and U15217 (N_15217,N_11812,N_11850);
nand U15218 (N_15218,N_9767,N_10963);
xnor U15219 (N_15219,N_9630,N_9121);
nor U15220 (N_15220,N_8133,N_10736);
or U15221 (N_15221,N_8487,N_11743);
or U15222 (N_15222,N_10343,N_10244);
xor U15223 (N_15223,N_8422,N_9516);
nor U15224 (N_15224,N_11435,N_10198);
or U15225 (N_15225,N_10847,N_11756);
xor U15226 (N_15226,N_8904,N_8101);
nand U15227 (N_15227,N_9929,N_10725);
nor U15228 (N_15228,N_10841,N_11260);
or U15229 (N_15229,N_10870,N_10639);
or U15230 (N_15230,N_10593,N_9454);
or U15231 (N_15231,N_8898,N_10499);
nor U15232 (N_15232,N_10725,N_8939);
nand U15233 (N_15233,N_8067,N_10056);
or U15234 (N_15234,N_8525,N_11394);
xnor U15235 (N_15235,N_10854,N_10268);
or U15236 (N_15236,N_8123,N_9126);
or U15237 (N_15237,N_10845,N_9505);
xor U15238 (N_15238,N_9894,N_8653);
and U15239 (N_15239,N_9496,N_9230);
or U15240 (N_15240,N_11027,N_11626);
xnor U15241 (N_15241,N_10657,N_10396);
nand U15242 (N_15242,N_9787,N_8130);
or U15243 (N_15243,N_9200,N_10260);
nand U15244 (N_15244,N_11149,N_10762);
or U15245 (N_15245,N_8233,N_11933);
and U15246 (N_15246,N_8087,N_8008);
nor U15247 (N_15247,N_9665,N_9586);
or U15248 (N_15248,N_8250,N_9067);
nand U15249 (N_15249,N_11624,N_8364);
xnor U15250 (N_15250,N_11544,N_8728);
and U15251 (N_15251,N_9477,N_11814);
or U15252 (N_15252,N_8478,N_10044);
nor U15253 (N_15253,N_9519,N_9383);
nor U15254 (N_15254,N_10972,N_11472);
xor U15255 (N_15255,N_8333,N_11266);
nor U15256 (N_15256,N_11316,N_11375);
and U15257 (N_15257,N_11593,N_9520);
and U15258 (N_15258,N_9665,N_10610);
or U15259 (N_15259,N_9673,N_11711);
and U15260 (N_15260,N_8796,N_11147);
nor U15261 (N_15261,N_11667,N_10054);
nor U15262 (N_15262,N_8993,N_8658);
nor U15263 (N_15263,N_11094,N_11183);
and U15264 (N_15264,N_9582,N_8085);
or U15265 (N_15265,N_10807,N_9215);
nor U15266 (N_15266,N_10064,N_10015);
and U15267 (N_15267,N_9987,N_9048);
and U15268 (N_15268,N_10745,N_8589);
or U15269 (N_15269,N_10223,N_8939);
nand U15270 (N_15270,N_8753,N_10165);
nor U15271 (N_15271,N_11758,N_11027);
or U15272 (N_15272,N_8280,N_10928);
and U15273 (N_15273,N_11863,N_9228);
or U15274 (N_15274,N_11096,N_11208);
and U15275 (N_15275,N_11947,N_8631);
nand U15276 (N_15276,N_10771,N_11201);
nor U15277 (N_15277,N_9350,N_8872);
and U15278 (N_15278,N_11420,N_10008);
nand U15279 (N_15279,N_9233,N_8377);
or U15280 (N_15280,N_11407,N_11064);
xor U15281 (N_15281,N_11316,N_10146);
nand U15282 (N_15282,N_11073,N_10347);
nor U15283 (N_15283,N_9787,N_9714);
or U15284 (N_15284,N_8813,N_8725);
and U15285 (N_15285,N_11978,N_9816);
or U15286 (N_15286,N_10193,N_11376);
xnor U15287 (N_15287,N_11752,N_10081);
nand U15288 (N_15288,N_10047,N_9815);
xnor U15289 (N_15289,N_10478,N_11840);
and U15290 (N_15290,N_11082,N_8069);
and U15291 (N_15291,N_11567,N_9612);
and U15292 (N_15292,N_11669,N_10178);
and U15293 (N_15293,N_10636,N_8011);
and U15294 (N_15294,N_11568,N_11814);
nand U15295 (N_15295,N_9818,N_9442);
nor U15296 (N_15296,N_10237,N_10941);
and U15297 (N_15297,N_9101,N_10639);
and U15298 (N_15298,N_8018,N_11406);
nand U15299 (N_15299,N_10290,N_8471);
nor U15300 (N_15300,N_10830,N_9858);
xnor U15301 (N_15301,N_11710,N_10543);
nor U15302 (N_15302,N_9826,N_10249);
or U15303 (N_15303,N_11481,N_10477);
nor U15304 (N_15304,N_11188,N_8951);
and U15305 (N_15305,N_11710,N_9292);
nor U15306 (N_15306,N_9041,N_11406);
or U15307 (N_15307,N_10096,N_9977);
and U15308 (N_15308,N_8160,N_9740);
and U15309 (N_15309,N_10153,N_10245);
nand U15310 (N_15310,N_11966,N_11793);
or U15311 (N_15311,N_11378,N_10029);
or U15312 (N_15312,N_9373,N_11536);
nor U15313 (N_15313,N_10030,N_8722);
and U15314 (N_15314,N_11743,N_8758);
or U15315 (N_15315,N_9204,N_9677);
nand U15316 (N_15316,N_11591,N_9647);
nand U15317 (N_15317,N_8966,N_8342);
or U15318 (N_15318,N_10381,N_10085);
nor U15319 (N_15319,N_8209,N_8339);
nand U15320 (N_15320,N_10378,N_9213);
and U15321 (N_15321,N_8058,N_10506);
nand U15322 (N_15322,N_9799,N_11525);
nor U15323 (N_15323,N_11991,N_11430);
nand U15324 (N_15324,N_11041,N_11019);
xnor U15325 (N_15325,N_10785,N_8959);
nand U15326 (N_15326,N_10836,N_8040);
or U15327 (N_15327,N_8841,N_11856);
nor U15328 (N_15328,N_11327,N_10209);
nand U15329 (N_15329,N_8413,N_9588);
or U15330 (N_15330,N_9931,N_10556);
or U15331 (N_15331,N_9520,N_11626);
nor U15332 (N_15332,N_8813,N_9535);
and U15333 (N_15333,N_11481,N_11621);
xnor U15334 (N_15334,N_10478,N_11446);
xor U15335 (N_15335,N_9066,N_8748);
and U15336 (N_15336,N_8695,N_8672);
nand U15337 (N_15337,N_10266,N_9430);
or U15338 (N_15338,N_9337,N_10516);
nand U15339 (N_15339,N_11320,N_11837);
xor U15340 (N_15340,N_8271,N_10282);
nand U15341 (N_15341,N_10040,N_9610);
nor U15342 (N_15342,N_11345,N_8474);
nor U15343 (N_15343,N_8771,N_10865);
nand U15344 (N_15344,N_8207,N_9945);
and U15345 (N_15345,N_10191,N_11381);
xor U15346 (N_15346,N_10266,N_10713);
and U15347 (N_15347,N_8563,N_9071);
xnor U15348 (N_15348,N_8976,N_9483);
or U15349 (N_15349,N_11808,N_10788);
or U15350 (N_15350,N_10571,N_11985);
and U15351 (N_15351,N_8320,N_10832);
or U15352 (N_15352,N_9878,N_8435);
xor U15353 (N_15353,N_9380,N_11658);
nor U15354 (N_15354,N_9205,N_10389);
nor U15355 (N_15355,N_11837,N_10316);
nor U15356 (N_15356,N_10056,N_9691);
nand U15357 (N_15357,N_10792,N_9232);
nand U15358 (N_15358,N_8489,N_11645);
or U15359 (N_15359,N_11284,N_9248);
xor U15360 (N_15360,N_9638,N_11344);
nand U15361 (N_15361,N_8666,N_11441);
nand U15362 (N_15362,N_8815,N_8000);
nor U15363 (N_15363,N_10848,N_11087);
nand U15364 (N_15364,N_10563,N_9159);
and U15365 (N_15365,N_8058,N_10059);
nor U15366 (N_15366,N_9170,N_8735);
nand U15367 (N_15367,N_10683,N_9375);
nor U15368 (N_15368,N_10879,N_11590);
or U15369 (N_15369,N_10685,N_10465);
xor U15370 (N_15370,N_11976,N_9568);
and U15371 (N_15371,N_9276,N_11199);
nor U15372 (N_15372,N_10779,N_9566);
nand U15373 (N_15373,N_8150,N_11134);
or U15374 (N_15374,N_10373,N_11390);
or U15375 (N_15375,N_10250,N_9456);
nand U15376 (N_15376,N_8539,N_9982);
and U15377 (N_15377,N_11744,N_11328);
nand U15378 (N_15378,N_11218,N_10126);
nor U15379 (N_15379,N_10274,N_10046);
or U15380 (N_15380,N_8470,N_10900);
nor U15381 (N_15381,N_10542,N_9200);
xor U15382 (N_15382,N_11587,N_9615);
or U15383 (N_15383,N_11978,N_10833);
nand U15384 (N_15384,N_9556,N_9252);
and U15385 (N_15385,N_11013,N_11545);
or U15386 (N_15386,N_10098,N_8421);
nand U15387 (N_15387,N_11779,N_9117);
nor U15388 (N_15388,N_10403,N_8287);
nor U15389 (N_15389,N_8189,N_9796);
nand U15390 (N_15390,N_11040,N_10967);
and U15391 (N_15391,N_8931,N_8458);
or U15392 (N_15392,N_11875,N_8158);
xnor U15393 (N_15393,N_8546,N_11314);
nand U15394 (N_15394,N_9064,N_10647);
or U15395 (N_15395,N_11653,N_11051);
nand U15396 (N_15396,N_8208,N_8775);
nand U15397 (N_15397,N_8664,N_9631);
or U15398 (N_15398,N_8454,N_10684);
nor U15399 (N_15399,N_9635,N_11717);
or U15400 (N_15400,N_11905,N_9934);
and U15401 (N_15401,N_9491,N_11612);
and U15402 (N_15402,N_9953,N_11463);
xnor U15403 (N_15403,N_11928,N_11204);
nand U15404 (N_15404,N_9715,N_8067);
and U15405 (N_15405,N_10692,N_8890);
xor U15406 (N_15406,N_11705,N_9779);
or U15407 (N_15407,N_10380,N_9558);
xor U15408 (N_15408,N_11622,N_11511);
or U15409 (N_15409,N_8667,N_11639);
xor U15410 (N_15410,N_11605,N_11518);
or U15411 (N_15411,N_10331,N_8192);
and U15412 (N_15412,N_9759,N_8752);
nor U15413 (N_15413,N_11773,N_11428);
xor U15414 (N_15414,N_11686,N_11245);
xnor U15415 (N_15415,N_10976,N_8292);
or U15416 (N_15416,N_10800,N_8123);
nor U15417 (N_15417,N_11951,N_10934);
nand U15418 (N_15418,N_10403,N_10054);
xnor U15419 (N_15419,N_8026,N_9192);
or U15420 (N_15420,N_8200,N_9714);
nand U15421 (N_15421,N_11981,N_9692);
or U15422 (N_15422,N_9564,N_8787);
or U15423 (N_15423,N_9653,N_11060);
xnor U15424 (N_15424,N_8145,N_8419);
nor U15425 (N_15425,N_10996,N_9854);
nor U15426 (N_15426,N_10895,N_8589);
nor U15427 (N_15427,N_8255,N_8227);
or U15428 (N_15428,N_9980,N_8801);
and U15429 (N_15429,N_8668,N_8085);
or U15430 (N_15430,N_9902,N_8731);
and U15431 (N_15431,N_8561,N_10238);
and U15432 (N_15432,N_10930,N_8735);
and U15433 (N_15433,N_9382,N_10433);
and U15434 (N_15434,N_10286,N_8493);
and U15435 (N_15435,N_9390,N_10654);
nor U15436 (N_15436,N_9115,N_10792);
nand U15437 (N_15437,N_8387,N_9844);
or U15438 (N_15438,N_10443,N_8363);
nand U15439 (N_15439,N_10868,N_8793);
nand U15440 (N_15440,N_10413,N_10887);
or U15441 (N_15441,N_9395,N_9765);
nand U15442 (N_15442,N_10139,N_9188);
or U15443 (N_15443,N_10619,N_11628);
nor U15444 (N_15444,N_11137,N_8731);
nand U15445 (N_15445,N_8076,N_8453);
nand U15446 (N_15446,N_9515,N_10747);
nor U15447 (N_15447,N_11271,N_10289);
or U15448 (N_15448,N_8805,N_10075);
nor U15449 (N_15449,N_8797,N_9126);
nor U15450 (N_15450,N_9261,N_10661);
nor U15451 (N_15451,N_8113,N_9336);
or U15452 (N_15452,N_10264,N_9915);
or U15453 (N_15453,N_9949,N_8103);
xor U15454 (N_15454,N_10988,N_11391);
or U15455 (N_15455,N_10034,N_11128);
nand U15456 (N_15456,N_10404,N_8966);
xor U15457 (N_15457,N_9395,N_11422);
nor U15458 (N_15458,N_10326,N_11881);
and U15459 (N_15459,N_11282,N_9698);
nor U15460 (N_15460,N_8409,N_8914);
or U15461 (N_15461,N_8508,N_11203);
nand U15462 (N_15462,N_10624,N_8104);
nor U15463 (N_15463,N_11615,N_8977);
xnor U15464 (N_15464,N_9402,N_11852);
or U15465 (N_15465,N_11633,N_8390);
or U15466 (N_15466,N_8871,N_10924);
nor U15467 (N_15467,N_9651,N_10012);
and U15468 (N_15468,N_8368,N_10956);
and U15469 (N_15469,N_11364,N_10805);
and U15470 (N_15470,N_9399,N_11610);
nor U15471 (N_15471,N_9441,N_9428);
or U15472 (N_15472,N_9008,N_9598);
nand U15473 (N_15473,N_8777,N_9244);
xnor U15474 (N_15474,N_10267,N_9861);
or U15475 (N_15475,N_9183,N_10322);
and U15476 (N_15476,N_9828,N_9792);
and U15477 (N_15477,N_11439,N_10297);
nand U15478 (N_15478,N_10959,N_9211);
or U15479 (N_15479,N_9127,N_9067);
or U15480 (N_15480,N_11802,N_8507);
and U15481 (N_15481,N_9850,N_9887);
nor U15482 (N_15482,N_11136,N_10410);
nor U15483 (N_15483,N_10090,N_8443);
nor U15484 (N_15484,N_10109,N_11484);
and U15485 (N_15485,N_9438,N_10204);
nor U15486 (N_15486,N_8229,N_8960);
and U15487 (N_15487,N_9962,N_10793);
nand U15488 (N_15488,N_11004,N_11751);
and U15489 (N_15489,N_10497,N_10180);
nor U15490 (N_15490,N_10499,N_10879);
or U15491 (N_15491,N_9491,N_11430);
and U15492 (N_15492,N_9705,N_11834);
xor U15493 (N_15493,N_11518,N_9029);
nand U15494 (N_15494,N_10449,N_8758);
nor U15495 (N_15495,N_9376,N_8940);
nor U15496 (N_15496,N_9557,N_8388);
or U15497 (N_15497,N_10355,N_8010);
nand U15498 (N_15498,N_11983,N_9011);
nor U15499 (N_15499,N_10276,N_11865);
and U15500 (N_15500,N_8070,N_9753);
nand U15501 (N_15501,N_11479,N_10339);
and U15502 (N_15502,N_11200,N_10322);
and U15503 (N_15503,N_10541,N_11179);
xor U15504 (N_15504,N_9439,N_11805);
xnor U15505 (N_15505,N_11113,N_9661);
and U15506 (N_15506,N_9996,N_10960);
and U15507 (N_15507,N_9735,N_8507);
and U15508 (N_15508,N_9541,N_9046);
and U15509 (N_15509,N_8962,N_11309);
nand U15510 (N_15510,N_11207,N_10504);
and U15511 (N_15511,N_9624,N_11361);
and U15512 (N_15512,N_10674,N_10827);
nor U15513 (N_15513,N_10077,N_8557);
or U15514 (N_15514,N_8003,N_9048);
and U15515 (N_15515,N_10766,N_10068);
and U15516 (N_15516,N_8558,N_8297);
nor U15517 (N_15517,N_10646,N_9781);
or U15518 (N_15518,N_9944,N_9654);
or U15519 (N_15519,N_9436,N_10505);
nor U15520 (N_15520,N_11990,N_8499);
xor U15521 (N_15521,N_9780,N_9914);
nand U15522 (N_15522,N_9686,N_11602);
or U15523 (N_15523,N_10027,N_8086);
or U15524 (N_15524,N_9336,N_10718);
nor U15525 (N_15525,N_8721,N_9206);
and U15526 (N_15526,N_11787,N_10772);
nor U15527 (N_15527,N_8877,N_10811);
xor U15528 (N_15528,N_10622,N_8374);
or U15529 (N_15529,N_8771,N_11598);
xor U15530 (N_15530,N_11442,N_9427);
and U15531 (N_15531,N_9186,N_9247);
xnor U15532 (N_15532,N_8997,N_10368);
and U15533 (N_15533,N_10841,N_8475);
nor U15534 (N_15534,N_9892,N_11239);
and U15535 (N_15535,N_11427,N_8111);
and U15536 (N_15536,N_8035,N_9731);
nand U15537 (N_15537,N_10008,N_11341);
nand U15538 (N_15538,N_9588,N_9916);
and U15539 (N_15539,N_9602,N_9005);
nor U15540 (N_15540,N_9971,N_10453);
and U15541 (N_15541,N_8398,N_11740);
or U15542 (N_15542,N_8280,N_8689);
nor U15543 (N_15543,N_11656,N_10888);
nand U15544 (N_15544,N_10389,N_9600);
and U15545 (N_15545,N_11194,N_10820);
nor U15546 (N_15546,N_9173,N_11862);
xnor U15547 (N_15547,N_10632,N_9895);
and U15548 (N_15548,N_9200,N_8893);
or U15549 (N_15549,N_8506,N_8651);
nand U15550 (N_15550,N_10781,N_8422);
nor U15551 (N_15551,N_9769,N_11186);
nor U15552 (N_15552,N_11924,N_8553);
nand U15553 (N_15553,N_11297,N_8001);
xnor U15554 (N_15554,N_9011,N_9830);
or U15555 (N_15555,N_8698,N_9302);
nor U15556 (N_15556,N_8314,N_9380);
nor U15557 (N_15557,N_11498,N_10172);
and U15558 (N_15558,N_8146,N_11482);
or U15559 (N_15559,N_9651,N_11708);
or U15560 (N_15560,N_9537,N_11408);
nor U15561 (N_15561,N_9849,N_8888);
or U15562 (N_15562,N_10210,N_9876);
or U15563 (N_15563,N_11268,N_9563);
and U15564 (N_15564,N_8704,N_8180);
or U15565 (N_15565,N_8477,N_10540);
xnor U15566 (N_15566,N_8245,N_8968);
or U15567 (N_15567,N_8999,N_11437);
and U15568 (N_15568,N_8863,N_10956);
or U15569 (N_15569,N_8337,N_10219);
or U15570 (N_15570,N_10282,N_10082);
and U15571 (N_15571,N_11500,N_10080);
or U15572 (N_15572,N_9366,N_9269);
and U15573 (N_15573,N_8351,N_9814);
xnor U15574 (N_15574,N_8861,N_10882);
nor U15575 (N_15575,N_9408,N_10241);
or U15576 (N_15576,N_10437,N_8931);
nand U15577 (N_15577,N_8916,N_9333);
nor U15578 (N_15578,N_11844,N_11953);
nand U15579 (N_15579,N_11070,N_8813);
or U15580 (N_15580,N_10479,N_11691);
nand U15581 (N_15581,N_9629,N_11101);
or U15582 (N_15582,N_11210,N_9636);
nor U15583 (N_15583,N_8197,N_10001);
or U15584 (N_15584,N_10105,N_9692);
or U15585 (N_15585,N_10856,N_9843);
or U15586 (N_15586,N_8572,N_8933);
nor U15587 (N_15587,N_8782,N_9739);
and U15588 (N_15588,N_8340,N_11355);
xor U15589 (N_15589,N_9062,N_9491);
and U15590 (N_15590,N_11803,N_8231);
nor U15591 (N_15591,N_11692,N_11734);
and U15592 (N_15592,N_8739,N_11917);
or U15593 (N_15593,N_11371,N_8591);
nand U15594 (N_15594,N_8614,N_9647);
xor U15595 (N_15595,N_11447,N_8208);
nand U15596 (N_15596,N_11854,N_9075);
and U15597 (N_15597,N_9857,N_8765);
nand U15598 (N_15598,N_8439,N_10949);
or U15599 (N_15599,N_9123,N_9882);
nor U15600 (N_15600,N_10200,N_8074);
and U15601 (N_15601,N_9759,N_9314);
and U15602 (N_15602,N_10656,N_8114);
or U15603 (N_15603,N_9075,N_8064);
nand U15604 (N_15604,N_8339,N_8301);
or U15605 (N_15605,N_11577,N_9201);
and U15606 (N_15606,N_10752,N_11666);
or U15607 (N_15607,N_11395,N_9435);
and U15608 (N_15608,N_10771,N_8958);
nor U15609 (N_15609,N_8062,N_10991);
or U15610 (N_15610,N_9467,N_8538);
and U15611 (N_15611,N_11679,N_8819);
or U15612 (N_15612,N_11318,N_10836);
nand U15613 (N_15613,N_11831,N_8179);
xor U15614 (N_15614,N_11775,N_8074);
and U15615 (N_15615,N_9126,N_9181);
nand U15616 (N_15616,N_8794,N_9985);
or U15617 (N_15617,N_10266,N_9697);
nand U15618 (N_15618,N_11071,N_9824);
xor U15619 (N_15619,N_8831,N_8400);
or U15620 (N_15620,N_9611,N_11386);
nor U15621 (N_15621,N_10678,N_11110);
and U15622 (N_15622,N_11198,N_11058);
or U15623 (N_15623,N_8966,N_8304);
or U15624 (N_15624,N_8133,N_8319);
nand U15625 (N_15625,N_8828,N_9625);
nand U15626 (N_15626,N_9698,N_8093);
xor U15627 (N_15627,N_9482,N_8833);
or U15628 (N_15628,N_11352,N_9406);
nor U15629 (N_15629,N_10126,N_8085);
xnor U15630 (N_15630,N_10446,N_11010);
nor U15631 (N_15631,N_8107,N_9364);
or U15632 (N_15632,N_11406,N_11801);
and U15633 (N_15633,N_9728,N_11869);
nand U15634 (N_15634,N_9802,N_8371);
xor U15635 (N_15635,N_8360,N_11474);
and U15636 (N_15636,N_8628,N_8701);
nor U15637 (N_15637,N_9700,N_9788);
nor U15638 (N_15638,N_10756,N_11474);
nor U15639 (N_15639,N_8276,N_11578);
and U15640 (N_15640,N_11272,N_8021);
nand U15641 (N_15641,N_11157,N_9612);
and U15642 (N_15642,N_9704,N_9761);
nor U15643 (N_15643,N_10778,N_9809);
nand U15644 (N_15644,N_11822,N_10288);
nand U15645 (N_15645,N_10605,N_10512);
nor U15646 (N_15646,N_10156,N_9019);
or U15647 (N_15647,N_8929,N_9189);
nand U15648 (N_15648,N_9268,N_11250);
nand U15649 (N_15649,N_10817,N_9401);
nand U15650 (N_15650,N_8867,N_9663);
or U15651 (N_15651,N_11869,N_10004);
nor U15652 (N_15652,N_8327,N_10510);
and U15653 (N_15653,N_11815,N_11017);
nand U15654 (N_15654,N_9090,N_9550);
nand U15655 (N_15655,N_9294,N_10778);
and U15656 (N_15656,N_11542,N_10400);
nor U15657 (N_15657,N_10719,N_8552);
nor U15658 (N_15658,N_9348,N_10912);
and U15659 (N_15659,N_10754,N_10611);
and U15660 (N_15660,N_10402,N_8750);
nor U15661 (N_15661,N_10371,N_8892);
nor U15662 (N_15662,N_11008,N_8978);
and U15663 (N_15663,N_9110,N_10209);
nor U15664 (N_15664,N_11702,N_9500);
or U15665 (N_15665,N_10595,N_9116);
xor U15666 (N_15666,N_11396,N_10910);
and U15667 (N_15667,N_10949,N_11612);
and U15668 (N_15668,N_10158,N_8731);
nand U15669 (N_15669,N_9230,N_8727);
nand U15670 (N_15670,N_11733,N_10788);
nor U15671 (N_15671,N_8910,N_8439);
and U15672 (N_15672,N_11521,N_8906);
or U15673 (N_15673,N_10594,N_10682);
xnor U15674 (N_15674,N_11856,N_8027);
and U15675 (N_15675,N_10161,N_8403);
xnor U15676 (N_15676,N_9637,N_11938);
nor U15677 (N_15677,N_10755,N_9609);
nand U15678 (N_15678,N_10037,N_11627);
xor U15679 (N_15679,N_9516,N_9843);
nand U15680 (N_15680,N_11317,N_8581);
nor U15681 (N_15681,N_8914,N_9078);
or U15682 (N_15682,N_8228,N_11722);
nand U15683 (N_15683,N_10195,N_8191);
nand U15684 (N_15684,N_8806,N_8010);
or U15685 (N_15685,N_8052,N_8902);
nand U15686 (N_15686,N_9927,N_11285);
nor U15687 (N_15687,N_10059,N_9806);
or U15688 (N_15688,N_8830,N_8722);
and U15689 (N_15689,N_8983,N_10171);
nor U15690 (N_15690,N_11418,N_11660);
nand U15691 (N_15691,N_11113,N_11054);
nand U15692 (N_15692,N_10967,N_9819);
nor U15693 (N_15693,N_10645,N_11358);
or U15694 (N_15694,N_8498,N_11873);
or U15695 (N_15695,N_8196,N_11903);
and U15696 (N_15696,N_10088,N_9687);
nor U15697 (N_15697,N_10927,N_10811);
nand U15698 (N_15698,N_11985,N_8660);
nand U15699 (N_15699,N_11842,N_10761);
or U15700 (N_15700,N_11420,N_11100);
and U15701 (N_15701,N_9194,N_11157);
xor U15702 (N_15702,N_10951,N_9253);
nand U15703 (N_15703,N_10107,N_9283);
nor U15704 (N_15704,N_11559,N_9110);
and U15705 (N_15705,N_10865,N_10026);
or U15706 (N_15706,N_9885,N_11386);
nand U15707 (N_15707,N_8023,N_9097);
nand U15708 (N_15708,N_11448,N_9158);
nand U15709 (N_15709,N_10988,N_10735);
nor U15710 (N_15710,N_9842,N_8780);
nor U15711 (N_15711,N_8138,N_9043);
nor U15712 (N_15712,N_9438,N_10771);
and U15713 (N_15713,N_8010,N_8589);
or U15714 (N_15714,N_11005,N_11098);
xnor U15715 (N_15715,N_10915,N_10008);
xor U15716 (N_15716,N_10238,N_10047);
xor U15717 (N_15717,N_9328,N_9384);
nor U15718 (N_15718,N_8372,N_8007);
or U15719 (N_15719,N_8972,N_11226);
or U15720 (N_15720,N_10919,N_10264);
and U15721 (N_15721,N_10081,N_10495);
or U15722 (N_15722,N_9078,N_9081);
nand U15723 (N_15723,N_11617,N_10324);
nand U15724 (N_15724,N_8621,N_8107);
or U15725 (N_15725,N_8781,N_9734);
nand U15726 (N_15726,N_11202,N_8636);
nand U15727 (N_15727,N_10567,N_9576);
nand U15728 (N_15728,N_9878,N_9505);
xnor U15729 (N_15729,N_8349,N_10154);
and U15730 (N_15730,N_11996,N_9302);
nor U15731 (N_15731,N_8814,N_9694);
xnor U15732 (N_15732,N_9843,N_8198);
xor U15733 (N_15733,N_9873,N_11013);
and U15734 (N_15734,N_8412,N_9357);
or U15735 (N_15735,N_9988,N_10652);
nor U15736 (N_15736,N_9541,N_10374);
or U15737 (N_15737,N_10799,N_8055);
nor U15738 (N_15738,N_11611,N_8777);
xor U15739 (N_15739,N_9561,N_11978);
or U15740 (N_15740,N_11316,N_9588);
nand U15741 (N_15741,N_10805,N_11764);
and U15742 (N_15742,N_9293,N_8505);
nor U15743 (N_15743,N_9825,N_8982);
nand U15744 (N_15744,N_10526,N_8551);
and U15745 (N_15745,N_8674,N_10707);
and U15746 (N_15746,N_8689,N_9279);
or U15747 (N_15747,N_8049,N_8349);
nand U15748 (N_15748,N_8040,N_8573);
or U15749 (N_15749,N_11055,N_9309);
nand U15750 (N_15750,N_8605,N_10140);
nor U15751 (N_15751,N_9543,N_8220);
nor U15752 (N_15752,N_11050,N_10628);
nor U15753 (N_15753,N_11959,N_10932);
xor U15754 (N_15754,N_10378,N_9030);
nor U15755 (N_15755,N_11422,N_10029);
and U15756 (N_15756,N_9588,N_9730);
nand U15757 (N_15757,N_8039,N_10747);
xor U15758 (N_15758,N_9258,N_8093);
nand U15759 (N_15759,N_10964,N_8865);
nand U15760 (N_15760,N_11185,N_10280);
nand U15761 (N_15761,N_10879,N_10305);
nor U15762 (N_15762,N_11478,N_9956);
or U15763 (N_15763,N_10323,N_8711);
and U15764 (N_15764,N_8622,N_8827);
xor U15765 (N_15765,N_10245,N_10787);
and U15766 (N_15766,N_9264,N_9021);
nor U15767 (N_15767,N_10881,N_8592);
or U15768 (N_15768,N_9143,N_11486);
nor U15769 (N_15769,N_9348,N_9095);
nor U15770 (N_15770,N_11851,N_9815);
or U15771 (N_15771,N_9851,N_8036);
xor U15772 (N_15772,N_10268,N_10705);
nor U15773 (N_15773,N_8400,N_9052);
nor U15774 (N_15774,N_10399,N_10733);
xnor U15775 (N_15775,N_11015,N_11258);
or U15776 (N_15776,N_10658,N_11822);
and U15777 (N_15777,N_11821,N_10340);
nor U15778 (N_15778,N_11682,N_10389);
and U15779 (N_15779,N_9076,N_11216);
nor U15780 (N_15780,N_8901,N_11059);
or U15781 (N_15781,N_11061,N_8772);
nor U15782 (N_15782,N_11464,N_11906);
nor U15783 (N_15783,N_10073,N_8581);
nand U15784 (N_15784,N_11596,N_10562);
nand U15785 (N_15785,N_8107,N_9226);
nor U15786 (N_15786,N_9527,N_11521);
and U15787 (N_15787,N_8190,N_11808);
nor U15788 (N_15788,N_11923,N_10341);
and U15789 (N_15789,N_9051,N_8526);
nor U15790 (N_15790,N_11436,N_9536);
nor U15791 (N_15791,N_8186,N_11438);
nor U15792 (N_15792,N_11610,N_11944);
or U15793 (N_15793,N_11255,N_9360);
nor U15794 (N_15794,N_9075,N_10521);
or U15795 (N_15795,N_8122,N_8711);
nor U15796 (N_15796,N_11576,N_8501);
nand U15797 (N_15797,N_8954,N_10129);
and U15798 (N_15798,N_9690,N_10497);
or U15799 (N_15799,N_11995,N_9126);
and U15800 (N_15800,N_8349,N_11315);
and U15801 (N_15801,N_10644,N_9754);
or U15802 (N_15802,N_11928,N_9480);
xor U15803 (N_15803,N_9780,N_11734);
nor U15804 (N_15804,N_8086,N_11324);
xnor U15805 (N_15805,N_9934,N_11418);
xnor U15806 (N_15806,N_8138,N_9446);
nor U15807 (N_15807,N_10690,N_10928);
and U15808 (N_15808,N_9265,N_9954);
and U15809 (N_15809,N_10695,N_9445);
and U15810 (N_15810,N_10965,N_8635);
or U15811 (N_15811,N_8064,N_9602);
nor U15812 (N_15812,N_9244,N_10002);
nand U15813 (N_15813,N_9866,N_10590);
xor U15814 (N_15814,N_11547,N_10386);
or U15815 (N_15815,N_9849,N_9009);
and U15816 (N_15816,N_8033,N_8118);
or U15817 (N_15817,N_10197,N_10048);
or U15818 (N_15818,N_10586,N_8632);
nand U15819 (N_15819,N_10720,N_8748);
nor U15820 (N_15820,N_10412,N_11236);
or U15821 (N_15821,N_9402,N_11178);
or U15822 (N_15822,N_8213,N_8644);
nor U15823 (N_15823,N_10882,N_9418);
xor U15824 (N_15824,N_10519,N_9879);
xor U15825 (N_15825,N_8267,N_8134);
and U15826 (N_15826,N_9980,N_9799);
or U15827 (N_15827,N_8073,N_11698);
or U15828 (N_15828,N_8041,N_11779);
and U15829 (N_15829,N_10455,N_9076);
and U15830 (N_15830,N_11724,N_11466);
nand U15831 (N_15831,N_11798,N_10582);
xnor U15832 (N_15832,N_8190,N_10971);
or U15833 (N_15833,N_9790,N_10816);
nor U15834 (N_15834,N_9522,N_11443);
and U15835 (N_15835,N_10689,N_10371);
and U15836 (N_15836,N_8175,N_8367);
nor U15837 (N_15837,N_10397,N_9930);
xnor U15838 (N_15838,N_8838,N_10765);
nand U15839 (N_15839,N_10349,N_11544);
nor U15840 (N_15840,N_11146,N_10580);
nand U15841 (N_15841,N_9505,N_10309);
and U15842 (N_15842,N_8645,N_11720);
or U15843 (N_15843,N_11193,N_11440);
nand U15844 (N_15844,N_8351,N_8681);
nand U15845 (N_15845,N_8247,N_9121);
nand U15846 (N_15846,N_8876,N_11743);
nor U15847 (N_15847,N_9196,N_10076);
or U15848 (N_15848,N_11155,N_9611);
xnor U15849 (N_15849,N_9050,N_9563);
or U15850 (N_15850,N_9734,N_10129);
nor U15851 (N_15851,N_8334,N_11215);
xor U15852 (N_15852,N_11516,N_9303);
and U15853 (N_15853,N_9237,N_8827);
nor U15854 (N_15854,N_9153,N_9455);
or U15855 (N_15855,N_10763,N_10684);
and U15856 (N_15856,N_9956,N_9314);
xor U15857 (N_15857,N_10033,N_8864);
xnor U15858 (N_15858,N_9327,N_10249);
nor U15859 (N_15859,N_11586,N_10565);
and U15860 (N_15860,N_11423,N_8190);
or U15861 (N_15861,N_9289,N_9632);
nor U15862 (N_15862,N_11190,N_11434);
nor U15863 (N_15863,N_8805,N_9553);
nand U15864 (N_15864,N_8569,N_9828);
xor U15865 (N_15865,N_10966,N_11738);
and U15866 (N_15866,N_8417,N_10997);
nor U15867 (N_15867,N_11784,N_10029);
nand U15868 (N_15868,N_10046,N_9900);
nor U15869 (N_15869,N_8834,N_8023);
or U15870 (N_15870,N_8812,N_10524);
nand U15871 (N_15871,N_10639,N_11284);
or U15872 (N_15872,N_10229,N_10931);
and U15873 (N_15873,N_9949,N_8641);
or U15874 (N_15874,N_8719,N_8237);
nor U15875 (N_15875,N_11433,N_9888);
or U15876 (N_15876,N_9779,N_8513);
nand U15877 (N_15877,N_11297,N_8772);
nand U15878 (N_15878,N_9670,N_10055);
or U15879 (N_15879,N_10712,N_10432);
xor U15880 (N_15880,N_9146,N_9634);
and U15881 (N_15881,N_8055,N_9519);
or U15882 (N_15882,N_8362,N_11920);
nor U15883 (N_15883,N_11443,N_10315);
or U15884 (N_15884,N_9885,N_9862);
nand U15885 (N_15885,N_8013,N_11371);
nand U15886 (N_15886,N_11895,N_10070);
xor U15887 (N_15887,N_9466,N_9220);
or U15888 (N_15888,N_8406,N_10201);
or U15889 (N_15889,N_10786,N_9732);
xor U15890 (N_15890,N_9655,N_9620);
and U15891 (N_15891,N_9910,N_9542);
and U15892 (N_15892,N_10467,N_9371);
and U15893 (N_15893,N_11454,N_11363);
nor U15894 (N_15894,N_9809,N_11000);
nand U15895 (N_15895,N_10129,N_11553);
nor U15896 (N_15896,N_9206,N_9458);
or U15897 (N_15897,N_10214,N_9558);
nor U15898 (N_15898,N_10823,N_10504);
and U15899 (N_15899,N_11759,N_9752);
nor U15900 (N_15900,N_8917,N_9670);
and U15901 (N_15901,N_11714,N_10152);
nor U15902 (N_15902,N_10028,N_9297);
nand U15903 (N_15903,N_8750,N_10121);
nor U15904 (N_15904,N_10382,N_9617);
or U15905 (N_15905,N_11736,N_9621);
or U15906 (N_15906,N_10416,N_9444);
and U15907 (N_15907,N_11949,N_9804);
nor U15908 (N_15908,N_8536,N_9094);
or U15909 (N_15909,N_11287,N_9613);
xnor U15910 (N_15910,N_11128,N_8802);
and U15911 (N_15911,N_10993,N_10472);
nor U15912 (N_15912,N_10568,N_8977);
or U15913 (N_15913,N_10000,N_10684);
and U15914 (N_15914,N_11534,N_10800);
nand U15915 (N_15915,N_10206,N_10660);
or U15916 (N_15916,N_8367,N_11237);
nor U15917 (N_15917,N_10468,N_8705);
nand U15918 (N_15918,N_8440,N_11662);
and U15919 (N_15919,N_9110,N_11761);
nor U15920 (N_15920,N_9995,N_9462);
nor U15921 (N_15921,N_9690,N_10206);
or U15922 (N_15922,N_11842,N_9871);
nor U15923 (N_15923,N_9271,N_8356);
and U15924 (N_15924,N_9996,N_10292);
and U15925 (N_15925,N_9238,N_8569);
or U15926 (N_15926,N_8972,N_10113);
xnor U15927 (N_15927,N_9164,N_8111);
and U15928 (N_15928,N_8766,N_10171);
or U15929 (N_15929,N_9136,N_10165);
nor U15930 (N_15930,N_10547,N_10673);
and U15931 (N_15931,N_9392,N_11627);
nor U15932 (N_15932,N_10779,N_9625);
xnor U15933 (N_15933,N_8689,N_10278);
or U15934 (N_15934,N_11824,N_10876);
and U15935 (N_15935,N_10123,N_9807);
nand U15936 (N_15936,N_10887,N_11300);
or U15937 (N_15937,N_9314,N_11011);
nor U15938 (N_15938,N_10550,N_10238);
nor U15939 (N_15939,N_8498,N_11922);
and U15940 (N_15940,N_11336,N_9375);
nand U15941 (N_15941,N_10436,N_8558);
or U15942 (N_15942,N_9970,N_9703);
nand U15943 (N_15943,N_8742,N_11968);
nand U15944 (N_15944,N_10545,N_11882);
or U15945 (N_15945,N_11290,N_10580);
and U15946 (N_15946,N_9247,N_11613);
nand U15947 (N_15947,N_11879,N_11184);
nand U15948 (N_15948,N_11283,N_11782);
xnor U15949 (N_15949,N_11832,N_10227);
nand U15950 (N_15950,N_9957,N_8435);
and U15951 (N_15951,N_10877,N_10816);
and U15952 (N_15952,N_11955,N_9376);
or U15953 (N_15953,N_11991,N_9244);
and U15954 (N_15954,N_8478,N_8813);
nand U15955 (N_15955,N_8689,N_9931);
and U15956 (N_15956,N_11122,N_8869);
nand U15957 (N_15957,N_8802,N_9825);
nand U15958 (N_15958,N_9439,N_9260);
and U15959 (N_15959,N_11696,N_8493);
and U15960 (N_15960,N_10258,N_11461);
nor U15961 (N_15961,N_10252,N_11353);
nand U15962 (N_15962,N_8363,N_10436);
and U15963 (N_15963,N_10476,N_10646);
and U15964 (N_15964,N_8123,N_8331);
nand U15965 (N_15965,N_11506,N_8519);
nor U15966 (N_15966,N_8726,N_8433);
or U15967 (N_15967,N_8986,N_10006);
nand U15968 (N_15968,N_10883,N_11409);
or U15969 (N_15969,N_10498,N_11045);
or U15970 (N_15970,N_10186,N_10172);
and U15971 (N_15971,N_11063,N_10366);
nor U15972 (N_15972,N_9398,N_9429);
and U15973 (N_15973,N_9610,N_9939);
and U15974 (N_15974,N_10634,N_8489);
or U15975 (N_15975,N_10768,N_11433);
xor U15976 (N_15976,N_11363,N_10546);
xnor U15977 (N_15977,N_8545,N_10477);
nor U15978 (N_15978,N_11105,N_11054);
nand U15979 (N_15979,N_11136,N_8882);
and U15980 (N_15980,N_11569,N_8731);
nand U15981 (N_15981,N_8940,N_8475);
or U15982 (N_15982,N_8500,N_9296);
nor U15983 (N_15983,N_11669,N_9212);
and U15984 (N_15984,N_9781,N_10204);
nand U15985 (N_15985,N_10322,N_10850);
nor U15986 (N_15986,N_10678,N_10360);
nor U15987 (N_15987,N_8143,N_9488);
nand U15988 (N_15988,N_8977,N_10702);
and U15989 (N_15989,N_11193,N_10260);
nor U15990 (N_15990,N_8372,N_9520);
xor U15991 (N_15991,N_11495,N_11771);
and U15992 (N_15992,N_11303,N_10703);
or U15993 (N_15993,N_8036,N_9195);
nand U15994 (N_15994,N_11132,N_10690);
or U15995 (N_15995,N_9758,N_10489);
or U15996 (N_15996,N_9774,N_10423);
nor U15997 (N_15997,N_8482,N_10659);
or U15998 (N_15998,N_10001,N_8332);
nor U15999 (N_15999,N_8501,N_10780);
nand U16000 (N_16000,N_12657,N_12570);
or U16001 (N_16001,N_15901,N_15667);
nand U16002 (N_16002,N_14736,N_13121);
nor U16003 (N_16003,N_15652,N_12887);
nand U16004 (N_16004,N_12847,N_14197);
or U16005 (N_16005,N_14720,N_14980);
nand U16006 (N_16006,N_13554,N_15714);
nor U16007 (N_16007,N_12926,N_12295);
or U16008 (N_16008,N_15273,N_15532);
and U16009 (N_16009,N_13021,N_12262);
and U16010 (N_16010,N_14245,N_14686);
nand U16011 (N_16011,N_12667,N_15298);
or U16012 (N_16012,N_12160,N_14178);
xnor U16013 (N_16013,N_14063,N_13447);
and U16014 (N_16014,N_12937,N_15982);
nor U16015 (N_16015,N_12624,N_14750);
nand U16016 (N_16016,N_12360,N_12168);
nand U16017 (N_16017,N_12930,N_12336);
nor U16018 (N_16018,N_15324,N_15183);
or U16019 (N_16019,N_13813,N_12817);
and U16020 (N_16020,N_13287,N_14957);
and U16021 (N_16021,N_13436,N_13179);
or U16022 (N_16022,N_14210,N_14311);
and U16023 (N_16023,N_13797,N_12804);
nor U16024 (N_16024,N_15097,N_14606);
nor U16025 (N_16025,N_13407,N_13917);
or U16026 (N_16026,N_15830,N_15777);
nor U16027 (N_16027,N_12653,N_13138);
nand U16028 (N_16028,N_12454,N_14159);
xnor U16029 (N_16029,N_14240,N_14101);
nor U16030 (N_16030,N_12080,N_14433);
and U16031 (N_16031,N_15340,N_15150);
and U16032 (N_16032,N_12618,N_12430);
or U16033 (N_16033,N_13546,N_14046);
nor U16034 (N_16034,N_14804,N_14819);
nor U16035 (N_16035,N_14473,N_14648);
or U16036 (N_16036,N_13064,N_15804);
nand U16037 (N_16037,N_14891,N_15552);
xnor U16038 (N_16038,N_12464,N_13865);
and U16039 (N_16039,N_15625,N_15424);
nand U16040 (N_16040,N_15789,N_12678);
nand U16041 (N_16041,N_13717,N_12146);
and U16042 (N_16042,N_12461,N_14278);
and U16043 (N_16043,N_14563,N_13847);
nand U16044 (N_16044,N_13539,N_12941);
or U16045 (N_16045,N_13943,N_12712);
xnor U16046 (N_16046,N_13861,N_13697);
nand U16047 (N_16047,N_14286,N_15690);
and U16048 (N_16048,N_14712,N_14139);
or U16049 (N_16049,N_12250,N_13532);
and U16050 (N_16050,N_12518,N_13578);
nor U16051 (N_16051,N_13915,N_12206);
or U16052 (N_16052,N_12153,N_15094);
and U16053 (N_16053,N_14727,N_14077);
or U16054 (N_16054,N_15743,N_15579);
nand U16055 (N_16055,N_14462,N_14468);
or U16056 (N_16056,N_14070,N_12501);
and U16057 (N_16057,N_15359,N_13784);
and U16058 (N_16058,N_13907,N_12021);
nand U16059 (N_16059,N_14066,N_13333);
nand U16060 (N_16060,N_15072,N_15208);
and U16061 (N_16061,N_15343,N_12274);
and U16062 (N_16062,N_14233,N_12876);
and U16063 (N_16063,N_15052,N_15856);
or U16064 (N_16064,N_13780,N_12787);
and U16065 (N_16065,N_12848,N_15556);
and U16066 (N_16066,N_15245,N_13715);
xnor U16067 (N_16067,N_15486,N_14050);
and U16068 (N_16068,N_14342,N_14598);
nand U16069 (N_16069,N_15931,N_13547);
and U16070 (N_16070,N_13485,N_14545);
xnor U16071 (N_16071,N_15685,N_12312);
and U16072 (N_16072,N_13599,N_14882);
xnor U16073 (N_16073,N_14190,N_15733);
or U16074 (N_16074,N_13916,N_14870);
nand U16075 (N_16075,N_14880,N_12695);
or U16076 (N_16076,N_14146,N_15598);
nand U16077 (N_16077,N_13875,N_14605);
nand U16078 (N_16078,N_14835,N_13348);
nand U16079 (N_16079,N_15291,N_12151);
xnor U16080 (N_16080,N_12949,N_13000);
and U16081 (N_16081,N_12414,N_13786);
and U16082 (N_16082,N_12526,N_13020);
and U16083 (N_16083,N_14639,N_14918);
and U16084 (N_16084,N_14215,N_13209);
and U16085 (N_16085,N_12382,N_13375);
nand U16086 (N_16086,N_15588,N_13435);
and U16087 (N_16087,N_13311,N_12664);
nand U16088 (N_16088,N_12942,N_14025);
or U16089 (N_16089,N_14080,N_13391);
nand U16090 (N_16090,N_14948,N_12010);
nand U16091 (N_16091,N_13268,N_14315);
xnor U16092 (N_16092,N_12474,N_14944);
xnor U16093 (N_16093,N_12300,N_14128);
or U16094 (N_16094,N_15122,N_12301);
and U16095 (N_16095,N_14725,N_15670);
or U16096 (N_16096,N_15417,N_15565);
or U16097 (N_16097,N_14372,N_14848);
xnor U16098 (N_16098,N_14138,N_15933);
nor U16099 (N_16099,N_12101,N_12736);
and U16100 (N_16100,N_12686,N_12573);
nor U16101 (N_16101,N_13884,N_14808);
nand U16102 (N_16102,N_12632,N_14553);
and U16103 (N_16103,N_15584,N_12794);
nand U16104 (N_16104,N_13041,N_15649);
nand U16105 (N_16105,N_13291,N_15900);
or U16106 (N_16106,N_15659,N_14551);
and U16107 (N_16107,N_12222,N_15555);
and U16108 (N_16108,N_13814,N_12985);
xnor U16109 (N_16109,N_14478,N_13241);
nor U16110 (N_16110,N_13558,N_15083);
nand U16111 (N_16111,N_12118,N_14923);
xnor U16112 (N_16112,N_13112,N_12568);
nand U16113 (N_16113,N_15802,N_15446);
nor U16114 (N_16114,N_15334,N_13449);
nor U16115 (N_16115,N_12698,N_15215);
nand U16116 (N_16116,N_12096,N_15076);
and U16117 (N_16117,N_12157,N_15525);
nand U16118 (N_16118,N_13973,N_15722);
nand U16119 (N_16119,N_12873,N_14257);
nor U16120 (N_16120,N_12419,N_12557);
nand U16121 (N_16121,N_13626,N_12018);
and U16122 (N_16122,N_15547,N_13747);
or U16123 (N_16123,N_14638,N_14224);
nor U16124 (N_16124,N_13197,N_13308);
nand U16125 (N_16125,N_12633,N_12842);
nand U16126 (N_16126,N_14464,N_12402);
and U16127 (N_16127,N_14792,N_14115);
nor U16128 (N_16128,N_14056,N_13432);
and U16129 (N_16129,N_15026,N_14065);
nand U16130 (N_16130,N_14079,N_14933);
or U16131 (N_16131,N_15842,N_15628);
xnor U16132 (N_16132,N_13018,N_14626);
and U16133 (N_16133,N_14749,N_12676);
nor U16134 (N_16134,N_12838,N_12379);
nand U16135 (N_16135,N_14893,N_14930);
and U16136 (N_16136,N_15730,N_15336);
nand U16137 (N_16137,N_12421,N_13065);
nor U16138 (N_16138,N_13662,N_13836);
or U16139 (N_16139,N_15571,N_15814);
or U16140 (N_16140,N_12580,N_15850);
nand U16141 (N_16141,N_12401,N_13981);
or U16142 (N_16142,N_13500,N_13200);
or U16143 (N_16143,N_15899,N_14603);
and U16144 (N_16144,N_15236,N_13649);
nor U16145 (N_16145,N_12017,N_14807);
or U16146 (N_16146,N_15347,N_13024);
nor U16147 (N_16147,N_13186,N_13322);
nor U16148 (N_16148,N_13983,N_12713);
or U16149 (N_16149,N_13605,N_14150);
nor U16150 (N_16150,N_13923,N_13094);
and U16151 (N_16151,N_15012,N_14732);
and U16152 (N_16152,N_14814,N_12437);
nand U16153 (N_16153,N_14423,N_13853);
and U16154 (N_16154,N_15744,N_13764);
and U16155 (N_16155,N_13690,N_15650);
and U16156 (N_16156,N_12861,N_13515);
nand U16157 (N_16157,N_15606,N_12384);
nand U16158 (N_16158,N_14557,N_12377);
or U16159 (N_16159,N_12614,N_12611);
or U16160 (N_16160,N_14041,N_15767);
and U16161 (N_16161,N_13001,N_15452);
nor U16162 (N_16162,N_12721,N_13410);
nand U16163 (N_16163,N_14986,N_12201);
or U16164 (N_16164,N_12114,N_12183);
xor U16165 (N_16165,N_14533,N_14729);
or U16166 (N_16166,N_12405,N_13686);
nand U16167 (N_16167,N_15871,N_15503);
and U16168 (N_16168,N_15411,N_15855);
xnor U16169 (N_16169,N_14656,N_15320);
or U16170 (N_16170,N_14955,N_12276);
nand U16171 (N_16171,N_14627,N_14906);
nand U16172 (N_16172,N_15870,N_13471);
or U16173 (N_16173,N_12293,N_14359);
and U16174 (N_16174,N_15618,N_13838);
nor U16175 (N_16175,N_12162,N_14486);
nor U16176 (N_16176,N_14477,N_14045);
nand U16177 (N_16177,N_14218,N_13905);
and U16178 (N_16178,N_12703,N_12111);
xor U16179 (N_16179,N_15294,N_13660);
nand U16180 (N_16180,N_13252,N_12292);
or U16181 (N_16181,N_15813,N_13644);
and U16182 (N_16182,N_12576,N_14476);
and U16183 (N_16183,N_15247,N_12148);
nand U16184 (N_16184,N_14508,N_15930);
nand U16185 (N_16185,N_13766,N_14873);
nand U16186 (N_16186,N_14206,N_14043);
nand U16187 (N_16187,N_12383,N_15891);
nand U16188 (N_16188,N_12751,N_15240);
or U16189 (N_16189,N_15926,N_15459);
and U16190 (N_16190,N_13123,N_13188);
nand U16191 (N_16191,N_12762,N_13376);
and U16192 (N_16192,N_12415,N_15084);
xor U16193 (N_16193,N_13840,N_12357);
nor U16194 (N_16194,N_15970,N_12832);
nor U16195 (N_16195,N_12207,N_12475);
nand U16196 (N_16196,N_13210,N_14756);
nor U16197 (N_16197,N_14172,N_15599);
nor U16198 (N_16198,N_15059,N_15011);
or U16199 (N_16199,N_12855,N_14740);
or U16200 (N_16200,N_12287,N_12772);
nand U16201 (N_16201,N_12102,N_14829);
or U16202 (N_16202,N_15302,N_15752);
nor U16203 (N_16203,N_14674,N_12273);
and U16204 (N_16204,N_12359,N_12354);
and U16205 (N_16205,N_13325,N_12725);
and U16206 (N_16206,N_14979,N_12652);
or U16207 (N_16207,N_15818,N_12947);
nand U16208 (N_16208,N_13800,N_12733);
nand U16209 (N_16209,N_14492,N_12124);
nor U16210 (N_16210,N_15402,N_12844);
or U16211 (N_16211,N_14442,N_13839);
nor U16212 (N_16212,N_15536,N_13505);
nand U16213 (N_16213,N_15338,N_15553);
nand U16214 (N_16214,N_12815,N_12409);
and U16215 (N_16215,N_14503,N_13672);
and U16216 (N_16216,N_14386,N_13159);
or U16217 (N_16217,N_15350,N_12885);
and U16218 (N_16218,N_13202,N_14722);
nand U16219 (N_16219,N_13652,N_14459);
and U16220 (N_16220,N_14576,N_15443);
nand U16221 (N_16221,N_13243,N_13193);
nand U16222 (N_16222,N_15176,N_12831);
nor U16223 (N_16223,N_13738,N_13349);
or U16224 (N_16224,N_12058,N_13297);
nand U16225 (N_16225,N_13835,N_14571);
or U16226 (N_16226,N_15389,N_12740);
nor U16227 (N_16227,N_15943,N_15160);
nand U16228 (N_16228,N_15998,N_14723);
nor U16229 (N_16229,N_13882,N_13961);
nor U16230 (N_16230,N_14033,N_13957);
or U16231 (N_16231,N_14775,N_13658);
or U16232 (N_16232,N_12988,N_15626);
nor U16233 (N_16233,N_14482,N_13567);
nand U16234 (N_16234,N_15576,N_13606);
and U16235 (N_16235,N_13426,N_15234);
xor U16236 (N_16236,N_13102,N_12784);
nand U16237 (N_16237,N_13185,N_13063);
nor U16238 (N_16238,N_12412,N_14897);
nand U16239 (N_16239,N_14177,N_12112);
and U16240 (N_16240,N_13373,N_12435);
nor U16241 (N_16241,N_12479,N_15121);
nand U16242 (N_16242,N_12198,N_12285);
or U16243 (N_16243,N_15762,N_12753);
nor U16244 (N_16244,N_14394,N_12852);
or U16245 (N_16245,N_12864,N_14213);
or U16246 (N_16246,N_15647,N_13344);
and U16247 (N_16247,N_13026,N_14573);
nand U16248 (N_16248,N_13509,N_12311);
and U16249 (N_16249,N_13269,N_14840);
xor U16250 (N_16250,N_13396,N_15913);
xor U16251 (N_16251,N_14498,N_13238);
or U16252 (N_16252,N_13248,N_15157);
nand U16253 (N_16253,N_13560,N_15037);
nand U16254 (N_16254,N_13737,N_13191);
and U16255 (N_16255,N_12001,N_12332);
and U16256 (N_16256,N_15041,N_13795);
nand U16257 (N_16257,N_14558,N_13262);
nand U16258 (N_16258,N_15622,N_15677);
xnor U16259 (N_16259,N_12981,N_13691);
or U16260 (N_16260,N_14708,N_13419);
nor U16261 (N_16261,N_13926,N_13870);
or U16262 (N_16262,N_14517,N_14337);
nand U16263 (N_16263,N_15297,N_13592);
or U16264 (N_16264,N_13888,N_12819);
nor U16265 (N_16265,N_14823,N_15429);
and U16266 (N_16266,N_13057,N_14937);
nor U16267 (N_16267,N_12647,N_12398);
or U16268 (N_16268,N_12532,N_13615);
xor U16269 (N_16269,N_13463,N_15885);
nand U16270 (N_16270,N_13139,N_15229);
nand U16271 (N_16271,N_14306,N_14984);
and U16272 (N_16272,N_12980,N_14281);
and U16273 (N_16273,N_12469,N_12404);
or U16274 (N_16274,N_15682,N_15066);
nor U16275 (N_16275,N_15522,N_15688);
nand U16276 (N_16276,N_15373,N_14003);
nor U16277 (N_16277,N_13351,N_15023);
xnor U16278 (N_16278,N_13734,N_14596);
nand U16279 (N_16279,N_12015,N_12498);
nor U16280 (N_16280,N_13997,N_12072);
nor U16281 (N_16281,N_12989,N_15371);
or U16282 (N_16282,N_13183,N_13437);
nor U16283 (N_16283,N_14682,N_15529);
or U16284 (N_16284,N_12269,N_13053);
nor U16285 (N_16285,N_15768,N_13037);
or U16286 (N_16286,N_15868,N_14564);
or U16287 (N_16287,N_13229,N_14529);
xnor U16288 (N_16288,N_12722,N_15039);
xnor U16289 (N_16289,N_12658,N_12438);
and U16290 (N_16290,N_12306,N_12688);
nor U16291 (N_16291,N_15491,N_12105);
nand U16292 (N_16292,N_12602,N_15713);
and U16293 (N_16293,N_15692,N_12245);
and U16294 (N_16294,N_15766,N_14650);
nor U16295 (N_16295,N_12954,N_14554);
nor U16296 (N_16296,N_13707,N_14812);
nand U16297 (N_16297,N_14152,N_15079);
nand U16298 (N_16298,N_14093,N_15672);
or U16299 (N_16299,N_12127,N_15268);
nand U16300 (N_16300,N_12597,N_12541);
nand U16301 (N_16301,N_14832,N_14964);
nand U16302 (N_16302,N_12425,N_15275);
nor U16303 (N_16303,N_15019,N_14616);
or U16304 (N_16304,N_15838,N_12824);
nor U16305 (N_16305,N_12506,N_15852);
nand U16306 (N_16306,N_15957,N_12716);
and U16307 (N_16307,N_12232,N_15138);
or U16308 (N_16308,N_12634,N_13281);
nand U16309 (N_16309,N_14321,N_13453);
nand U16310 (N_16310,N_13153,N_12033);
or U16311 (N_16311,N_13220,N_13806);
nor U16312 (N_16312,N_13774,N_13035);
or U16313 (N_16313,N_13036,N_15004);
nor U16314 (N_16314,N_15758,N_14110);
nand U16315 (N_16315,N_12559,N_14105);
or U16316 (N_16316,N_13616,N_14693);
nand U16317 (N_16317,N_13395,N_12869);
xnor U16318 (N_16318,N_13673,N_15535);
xor U16319 (N_16319,N_13904,N_13052);
and U16320 (N_16320,N_14989,N_15400);
nand U16321 (N_16321,N_13909,N_14324);
nor U16322 (N_16322,N_12279,N_15954);
nor U16323 (N_16323,N_14249,N_15825);
or U16324 (N_16324,N_13594,N_15663);
nand U16325 (N_16325,N_13450,N_12940);
xnor U16326 (N_16326,N_12390,N_14834);
nor U16327 (N_16327,N_15395,N_13060);
nand U16328 (N_16328,N_13571,N_15573);
nand U16329 (N_16329,N_15388,N_13821);
nor U16330 (N_16330,N_14026,N_12860);
or U16331 (N_16331,N_13479,N_13996);
nand U16332 (N_16332,N_13591,N_13557);
and U16333 (N_16333,N_14106,N_15712);
and U16334 (N_16334,N_13086,N_13767);
nor U16335 (N_16335,N_14223,N_12061);
nand U16336 (N_16336,N_15551,N_13131);
and U16337 (N_16337,N_14474,N_15252);
nand U16338 (N_16338,N_13337,N_13951);
and U16339 (N_16339,N_12671,N_15948);
or U16340 (N_16340,N_14828,N_14922);
and U16341 (N_16341,N_12005,N_14861);
nand U16342 (N_16342,N_12076,N_12055);
xnor U16343 (N_16343,N_12303,N_15641);
xor U16344 (N_16344,N_13089,N_13639);
nand U16345 (N_16345,N_14787,N_14597);
nand U16346 (N_16346,N_14670,N_15449);
nand U16347 (N_16347,N_12447,N_12897);
and U16348 (N_16348,N_12830,N_12732);
nand U16349 (N_16349,N_12696,N_14319);
or U16350 (N_16350,N_13440,N_12494);
nand U16351 (N_16351,N_13461,N_14988);
xor U16352 (N_16352,N_14769,N_14538);
and U16353 (N_16353,N_13543,N_14928);
nor U16354 (N_16354,N_14865,N_13489);
or U16355 (N_16355,N_15495,N_12685);
xnor U16356 (N_16356,N_12259,N_12208);
or U16357 (N_16357,N_13666,N_12103);
nor U16358 (N_16358,N_15178,N_14560);
and U16359 (N_16359,N_13977,N_12745);
or U16360 (N_16360,N_12243,N_12452);
or U16361 (N_16361,N_14345,N_15829);
or U16362 (N_16362,N_12814,N_14879);
and U16363 (N_16363,N_13226,N_12534);
nor U16364 (N_16364,N_14577,N_15960);
xnor U16365 (N_16365,N_13796,N_15863);
or U16366 (N_16366,N_15872,N_12434);
nand U16367 (N_16367,N_15005,N_12582);
and U16368 (N_16368,N_15706,N_14440);
nand U16369 (N_16369,N_12145,N_13775);
nor U16370 (N_16370,N_12710,N_15664);
and U16371 (N_16371,N_14509,N_15456);
nand U16372 (N_16372,N_12648,N_12239);
and U16373 (N_16373,N_12347,N_15642);
and U16374 (N_16374,N_14518,N_15008);
or U16375 (N_16375,N_12737,N_12872);
nand U16376 (N_16376,N_15977,N_15660);
and U16377 (N_16377,N_13743,N_13809);
nor U16378 (N_16378,N_13128,N_12829);
nand U16379 (N_16379,N_14241,N_13992);
and U16380 (N_16380,N_14112,N_14734);
nor U16381 (N_16381,N_15082,N_13274);
or U16382 (N_16382,N_14743,N_14731);
or U16383 (N_16383,N_13043,N_14878);
nand U16384 (N_16384,N_15971,N_14718);
nor U16385 (N_16385,N_14364,N_14332);
and U16386 (N_16386,N_13880,N_15187);
nor U16387 (N_16387,N_14211,N_12397);
nor U16388 (N_16388,N_12659,N_14992);
nand U16389 (N_16389,N_12305,N_15624);
nand U16390 (N_16390,N_14636,N_13196);
nand U16391 (N_16391,N_13386,N_13103);
or U16392 (N_16392,N_14131,N_13482);
nand U16393 (N_16393,N_12428,N_13849);
nand U16394 (N_16394,N_15186,N_13326);
and U16395 (N_16395,N_15009,N_14073);
and U16396 (N_16396,N_15638,N_12350);
nor U16397 (N_16397,N_15918,N_13411);
xnor U16398 (N_16398,N_15505,N_12368);
or U16399 (N_16399,N_13045,N_13687);
nor U16400 (N_16400,N_15474,N_14830);
nand U16401 (N_16401,N_15549,N_14011);
nand U16402 (N_16402,N_13228,N_14429);
xor U16403 (N_16403,N_12036,N_12951);
nand U16404 (N_16404,N_12014,N_14029);
nor U16405 (N_16405,N_15678,N_14000);
nor U16406 (N_16406,N_14480,N_12226);
nand U16407 (N_16407,N_12781,N_15578);
xor U16408 (N_16408,N_14569,N_14356);
nand U16409 (N_16409,N_13807,N_15177);
nand U16410 (N_16410,N_12782,N_13712);
or U16411 (N_16411,N_13679,N_15546);
and U16412 (N_16412,N_13412,N_13015);
and U16413 (N_16413,N_14293,N_15194);
xnor U16414 (N_16414,N_12133,N_13858);
nand U16415 (N_16415,N_15086,N_13214);
or U16416 (N_16416,N_14303,N_12436);
nand U16417 (N_16417,N_15633,N_12251);
xor U16418 (N_16418,N_15007,N_14688);
nand U16419 (N_16419,N_13106,N_13418);
nor U16420 (N_16420,N_14212,N_14995);
and U16421 (N_16421,N_15296,N_12349);
nor U16422 (N_16422,N_15407,N_15329);
and U16423 (N_16423,N_13995,N_13250);
or U16424 (N_16424,N_14994,N_14646);
nor U16425 (N_16425,N_14901,N_15498);
and U16426 (N_16426,N_13745,N_15490);
nor U16427 (N_16427,N_13318,N_15447);
and U16428 (N_16428,N_14284,N_13530);
nor U16429 (N_16429,N_15363,N_14120);
and U16430 (N_16430,N_12862,N_15890);
nand U16431 (N_16431,N_15997,N_12047);
nand U16432 (N_16432,N_12955,N_14887);
or U16433 (N_16433,N_15808,N_15413);
xor U16434 (N_16434,N_14299,N_12697);
nand U16435 (N_16435,N_13730,N_13079);
and U16436 (N_16436,N_14341,N_13177);
or U16437 (N_16437,N_12044,N_13946);
and U16438 (N_16438,N_12040,N_13940);
nand U16439 (N_16439,N_12922,N_13478);
or U16440 (N_16440,N_15457,N_14519);
nor U16441 (N_16441,N_12975,N_13285);
and U16442 (N_16442,N_12711,N_15892);
or U16443 (N_16443,N_14430,N_15708);
nor U16444 (N_16444,N_13488,N_14970);
nor U16445 (N_16445,N_14956,N_14811);
xnor U16446 (N_16446,N_12902,N_12063);
nand U16447 (N_16447,N_13335,N_14107);
and U16448 (N_16448,N_14751,N_14161);
or U16449 (N_16449,N_15103,N_15292);
nand U16450 (N_16450,N_15541,N_12598);
and U16451 (N_16451,N_15455,N_12760);
nor U16452 (N_16452,N_14347,N_13618);
nor U16453 (N_16453,N_12215,N_13161);
xnor U16454 (N_16454,N_14242,N_14963);
or U16455 (N_16455,N_13938,N_14782);
nand U16456 (N_16456,N_13319,N_14921);
nor U16457 (N_16457,N_12630,N_14565);
xnor U16458 (N_16458,N_14130,N_12070);
nand U16459 (N_16459,N_12738,N_15366);
and U16460 (N_16460,N_12317,N_15603);
nand U16461 (N_16461,N_12025,N_12179);
nor U16462 (N_16462,N_14491,N_13289);
nand U16463 (N_16463,N_13655,N_14399);
or U16464 (N_16464,N_12073,N_15875);
xor U16465 (N_16465,N_12533,N_12564);
or U16466 (N_16466,N_14783,N_14925);
nand U16467 (N_16467,N_13187,N_13493);
xnor U16468 (N_16468,N_14618,N_15799);
and U16469 (N_16469,N_15837,N_15787);
and U16470 (N_16470,N_13602,N_13523);
and U16471 (N_16471,N_15147,N_14525);
nor U16472 (N_16472,N_14421,N_15662);
nor U16473 (N_16473,N_13312,N_13081);
or U16474 (N_16474,N_15514,N_14987);
or U16475 (N_16475,N_12366,N_14746);
and U16476 (N_16476,N_15054,N_14393);
nor U16477 (N_16477,N_12704,N_15062);
or U16478 (N_16478,N_15462,N_12190);
and U16479 (N_16479,N_12229,N_12050);
and U16480 (N_16480,N_13075,N_15477);
xnor U16481 (N_16481,N_12779,N_13696);
and U16482 (N_16482,N_13182,N_13919);
nand U16483 (N_16483,N_13459,N_13657);
nor U16484 (N_16484,N_13999,N_12159);
or U16485 (N_16485,N_13154,N_12596);
or U16486 (N_16486,N_14758,N_14903);
nor U16487 (N_16487,N_14232,N_12242);
and U16488 (N_16488,N_15902,N_15387);
and U16489 (N_16489,N_15985,N_13711);
and U16490 (N_16490,N_13044,N_14762);
nand U16491 (N_16491,N_13140,N_13347);
nand U16492 (N_16492,N_14199,N_12482);
xor U16493 (N_16493,N_12726,N_14119);
and U16494 (N_16494,N_12846,N_13027);
nand U16495 (N_16495,N_15508,N_15778);
nor U16496 (N_16496,N_12705,N_12592);
or U16497 (N_16497,N_12174,N_12363);
and U16498 (N_16498,N_12458,N_15595);
nor U16499 (N_16499,N_15727,N_14791);
or U16500 (N_16500,N_12042,N_14967);
and U16501 (N_16501,N_13720,N_14827);
or U16502 (N_16502,N_12075,N_15489);
nand U16503 (N_16503,N_15705,N_14037);
nor U16504 (N_16504,N_15096,N_14087);
nor U16505 (N_16505,N_14204,N_14449);
or U16506 (N_16506,N_12545,N_15248);
nor U16507 (N_16507,N_15745,N_12020);
and U16508 (N_16508,N_12600,N_13190);
nor U16509 (N_16509,N_14135,N_15128);
nand U16510 (N_16510,N_13964,N_12087);
nor U16511 (N_16511,N_14927,N_15300);
xnor U16512 (N_16512,N_15637,N_12318);
and U16513 (N_16513,N_13700,N_13481);
nand U16514 (N_16514,N_13096,N_12643);
nand U16515 (N_16515,N_13483,N_14806);
or U16516 (N_16516,N_15952,N_12391);
and U16517 (N_16517,N_14523,N_13815);
xor U16518 (N_16518,N_15791,N_15759);
or U16519 (N_16519,N_12258,N_13744);
nand U16520 (N_16520,N_13842,N_15843);
nand U16521 (N_16521,N_14678,N_13245);
and U16522 (N_16522,N_12086,N_15999);
and U16523 (N_16523,N_12982,N_12097);
and U16524 (N_16524,N_13944,N_14428);
nor U16525 (N_16525,N_15949,N_15718);
or U16526 (N_16526,N_13846,N_14935);
nand U16527 (N_16527,N_14524,N_14309);
or U16528 (N_16528,N_13253,N_13897);
or U16529 (N_16529,N_13778,N_12520);
and U16530 (N_16530,N_12769,N_13793);
and U16531 (N_16531,N_15040,N_15331);
or U16532 (N_16532,N_14623,N_14051);
nand U16533 (N_16533,N_12607,N_13521);
or U16534 (N_16534,N_15807,N_12267);
and U16535 (N_16535,N_12750,N_12752);
and U16536 (N_16536,N_15734,N_13934);
and U16537 (N_16537,N_12283,N_15380);
or U16538 (N_16538,N_15276,N_13549);
nand U16539 (N_16539,N_12903,N_12466);
xnor U16540 (N_16540,N_12535,N_13912);
xnor U16541 (N_16541,N_12770,N_12636);
xor U16542 (N_16542,N_12766,N_13100);
nor U16543 (N_16543,N_13894,N_14996);
nor U16544 (N_16544,N_14990,N_12549);
and U16545 (N_16545,N_12680,N_12008);
nand U16546 (N_16546,N_12593,N_15434);
or U16547 (N_16547,N_13429,N_13498);
nor U16548 (N_16548,N_12759,N_15544);
nor U16549 (N_16549,N_14247,N_15492);
xnor U16550 (N_16550,N_14238,N_15418);
and U16551 (N_16551,N_14192,N_12866);
or U16552 (N_16552,N_12140,N_15305);
nor U16553 (N_16553,N_15639,N_14755);
and U16554 (N_16554,N_13039,N_14877);
nor U16555 (N_16555,N_13785,N_12645);
nor U16556 (N_16556,N_15093,N_13279);
nor U16557 (N_16557,N_14103,N_13092);
and U16558 (N_16558,N_13752,N_12000);
nand U16559 (N_16559,N_12064,N_15835);
nand U16560 (N_16560,N_12192,N_12209);
nor U16561 (N_16561,N_15155,N_12994);
and U16562 (N_16562,N_12211,N_15510);
nand U16563 (N_16563,N_13088,N_12165);
and U16564 (N_16564,N_12032,N_15607);
and U16565 (N_16565,N_13473,N_14274);
nor U16566 (N_16566,N_13540,N_14719);
and U16567 (N_16567,N_13129,N_12356);
and U16568 (N_16568,N_12834,N_12387);
nand U16569 (N_16569,N_13680,N_13513);
nor U16570 (N_16570,N_12623,N_14296);
and U16571 (N_16571,N_14282,N_15381);
nor U16572 (N_16572,N_14259,N_14036);
or U16573 (N_16573,N_14615,N_15220);
or U16574 (N_16574,N_12761,N_14006);
nand U16575 (N_16575,N_12756,N_15360);
or U16576 (N_16576,N_15239,N_15136);
nand U16577 (N_16577,N_15562,N_15785);
nor U16578 (N_16578,N_12135,N_12984);
nor U16579 (N_16579,N_12193,N_13416);
or U16580 (N_16580,N_14612,N_12799);
nand U16581 (N_16581,N_12386,N_12516);
nand U16582 (N_16582,N_14916,N_12868);
and U16583 (N_16583,N_12875,N_12281);
nand U16584 (N_16584,N_15438,N_12631);
nand U16585 (N_16585,N_14378,N_15849);
nor U16586 (N_16586,N_15884,N_13862);
or U16587 (N_16587,N_14116,N_14689);
nor U16588 (N_16588,N_12604,N_13127);
nand U16589 (N_16589,N_13107,N_15906);
nor U16590 (N_16590,N_13506,N_14448);
xor U16591 (N_16591,N_15728,N_13918);
or U16592 (N_16592,N_12039,N_15460);
nor U16593 (N_16593,N_14329,N_13484);
or U16594 (N_16594,N_12825,N_15761);
nor U16595 (N_16595,N_13357,N_14845);
nand U16596 (N_16596,N_13249,N_13804);
xor U16597 (N_16597,N_15224,N_15107);
nor U16598 (N_16598,N_14495,N_14526);
and U16599 (N_16599,N_15038,N_15858);
nand U16600 (N_16600,N_14535,N_13421);
or U16601 (N_16601,N_15738,N_15002);
nand U16602 (N_16602,N_12818,N_12517);
xnor U16603 (N_16603,N_13763,N_15064);
nand U16604 (N_16604,N_13722,N_14562);
or U16605 (N_16605,N_14941,N_14471);
and U16606 (N_16606,N_12244,N_12544);
or U16607 (N_16607,N_13305,N_12969);
and U16608 (N_16608,N_12441,N_12329);
nand U16609 (N_16609,N_15399,N_12575);
nor U16610 (N_16610,N_13405,N_14797);
nor U16611 (N_16611,N_13716,N_14654);
nand U16612 (N_16612,N_13619,N_13073);
nor U16613 (N_16613,N_13544,N_14888);
or U16614 (N_16614,N_15878,N_13490);
or U16615 (N_16615,N_13794,N_13116);
nand U16616 (N_16616,N_12660,N_15161);
or U16617 (N_16617,N_13520,N_14619);
nor U16618 (N_16618,N_14629,N_14088);
and U16619 (N_16619,N_15558,N_15036);
nand U16620 (N_16620,N_14302,N_13910);
nor U16621 (N_16621,N_15317,N_13577);
and U16622 (N_16622,N_14894,N_15749);
nand U16623 (N_16623,N_15694,N_15521);
and U16624 (N_16624,N_15720,N_15115);
nor U16625 (N_16625,N_12361,N_13848);
xor U16626 (N_16626,N_15506,N_15600);
nor U16627 (N_16627,N_15596,N_14643);
and U16628 (N_16628,N_14153,N_15235);
and U16629 (N_16629,N_14010,N_12399);
xor U16630 (N_16630,N_13047,N_13380);
nand U16631 (N_16631,N_15746,N_12187);
nor U16632 (N_16632,N_12218,N_13545);
nand U16633 (N_16633,N_12558,N_12120);
and U16634 (N_16634,N_12049,N_15679);
nor U16635 (N_16635,N_13630,N_12407);
xnor U16636 (N_16636,N_12327,N_14069);
and U16637 (N_16637,N_13585,N_15567);
and U16638 (N_16638,N_14234,N_15335);
and U16639 (N_16639,N_12476,N_13645);
nor U16640 (N_16640,N_15898,N_12572);
nor U16641 (N_16641,N_15233,N_14134);
nor U16642 (N_16642,N_13114,N_15149);
and U16643 (N_16643,N_13176,N_14714);
and U16644 (N_16644,N_13332,N_13782);
and U16645 (N_16645,N_12983,N_12478);
or U16646 (N_16646,N_12473,N_12735);
and U16647 (N_16647,N_15415,N_13962);
nor U16648 (N_16648,N_12141,N_15938);
or U16649 (N_16649,N_15069,N_14264);
nand U16650 (N_16650,N_14334,N_15472);
nor U16651 (N_16651,N_15794,N_14298);
nor U16652 (N_16652,N_13501,N_12205);
or U16653 (N_16653,N_13553,N_13283);
xor U16654 (N_16654,N_14340,N_15151);
nand U16655 (N_16655,N_15634,N_14113);
and U16656 (N_16656,N_12747,N_13298);
xnor U16657 (N_16657,N_15826,N_13508);
and U16658 (N_16658,N_15349,N_12649);
nor U16659 (N_16659,N_13580,N_14265);
nand U16660 (N_16660,N_13869,N_12371);
nand U16661 (N_16661,N_12186,N_14071);
nand U16662 (N_16662,N_13146,N_13422);
or U16663 (N_16663,N_12024,N_15771);
or U16664 (N_16664,N_15687,N_13566);
nor U16665 (N_16665,N_14383,N_13005);
or U16666 (N_16666,N_15436,N_14588);
xor U16667 (N_16667,N_14022,N_13142);
or U16668 (N_16668,N_13109,N_12918);
xnor U16669 (N_16669,N_14475,N_15962);
nor U16670 (N_16670,N_15152,N_15731);
xnor U16671 (N_16671,N_12655,N_12376);
and U16672 (N_16672,N_14450,N_12791);
xor U16673 (N_16673,N_15202,N_14602);
or U16674 (N_16674,N_14697,N_14905);
or U16675 (N_16675,N_13596,N_12635);
or U16676 (N_16676,N_15674,N_15853);
nor U16677 (N_16677,N_15994,N_15001);
nor U16678 (N_16678,N_14360,N_12471);
or U16679 (N_16679,N_12027,N_13320);
and U16680 (N_16680,N_13165,N_13812);
nand U16681 (N_16681,N_14851,N_13406);
or U16682 (N_16682,N_15665,N_12741);
xor U16683 (N_16683,N_12139,N_14488);
nand U16684 (N_16684,N_14427,N_13709);
nor U16685 (N_16685,N_15286,N_13620);
nor U16686 (N_16686,N_14680,N_15604);
nor U16687 (N_16687,N_13756,N_14086);
nand U16688 (N_16688,N_15632,N_14841);
nand U16689 (N_16689,N_12884,N_15266);
nor U16690 (N_16690,N_15669,N_12933);
or U16691 (N_16691,N_15385,N_14484);
and U16692 (N_16692,N_12927,N_12315);
or U16693 (N_16693,N_12874,N_14978);
nor U16694 (N_16694,N_12065,N_12442);
xnor U16695 (N_16695,N_12424,N_13956);
and U16696 (N_16696,N_15190,N_13388);
or U16697 (N_16697,N_15699,N_13040);
xor U16698 (N_16698,N_13642,N_14952);
and U16699 (N_16699,N_13878,N_14225);
or U16700 (N_16700,N_13234,N_13315);
or U16701 (N_16701,N_15085,N_13914);
or U16702 (N_16702,N_13729,N_12925);
xnor U16703 (N_16703,N_13217,N_15163);
nor U16704 (N_16704,N_13452,N_14396);
and U16705 (N_16705,N_13090,N_15698);
and U16706 (N_16706,N_14203,N_15916);
nor U16707 (N_16707,N_15958,N_13256);
and U16708 (N_16708,N_15601,N_12871);
nand U16709 (N_16709,N_14601,N_15458);
nor U16710 (N_16710,N_12684,N_12675);
nand U16711 (N_16711,N_12615,N_14857);
nor U16712 (N_16712,N_12484,N_15511);
and U16713 (N_16713,N_15995,N_12389);
xnor U16714 (N_16714,N_15815,N_14424);
and U16715 (N_16715,N_15270,N_14358);
and U16716 (N_16716,N_13739,N_15993);
nor U16717 (N_16717,N_15451,N_15857);
nor U16718 (N_16718,N_15193,N_15614);
or U16719 (N_16719,N_15527,N_12013);
nand U16720 (N_16720,N_15534,N_13542);
nor U16721 (N_16721,N_14958,N_13514);
and U16722 (N_16722,N_14363,N_15854);
xor U16723 (N_16723,N_12883,N_12298);
or U16724 (N_16724,N_12028,N_14843);
or U16725 (N_16725,N_13003,N_14084);
xor U16726 (N_16726,N_14300,N_14578);
and U16727 (N_16727,N_12007,N_13384);
nor U16728 (N_16728,N_15393,N_12620);
nor U16729 (N_16729,N_13694,N_13781);
xor U16730 (N_16730,N_14920,N_15022);
and U16731 (N_16731,N_13356,N_15016);
nand U16732 (N_16732,N_15561,N_12497);
nor U16733 (N_16733,N_12504,N_13985);
or U16734 (N_16734,N_14123,N_13583);
xnor U16735 (N_16735,N_13381,N_15704);
and U16736 (N_16736,N_12138,N_14929);
xnor U16737 (N_16737,N_14163,N_14831);
xor U16738 (N_16738,N_13049,N_13232);
nor U16739 (N_16739,N_15441,N_14763);
nand U16740 (N_16740,N_15792,N_12893);
nor U16741 (N_16741,N_15479,N_15048);
or U16742 (N_16742,N_12197,N_15589);
nand U16743 (N_16743,N_12012,N_15216);
nand U16744 (N_16744,N_14291,N_12789);
or U16745 (N_16745,N_14133,N_15619);
xor U16746 (N_16746,N_13430,N_15635);
and U16747 (N_16747,N_12979,N_12960);
and U16748 (N_16748,N_12542,N_14158);
or U16749 (N_16749,N_13495,N_12067);
nor U16750 (N_16750,N_15397,N_13982);
or U16751 (N_16751,N_13952,N_15132);
nor U16752 (N_16752,N_13098,N_15228);
or U16753 (N_16753,N_12233,N_14975);
nor U16754 (N_16754,N_14097,N_13574);
and U16755 (N_16755,N_15783,N_14771);
nor U16756 (N_16756,N_15570,N_15108);
nor U16757 (N_16757,N_15355,N_15199);
nand U16758 (N_16758,N_12282,N_12003);
and U16759 (N_16759,N_15288,N_14940);
and U16760 (N_16760,N_12246,N_14122);
nor U16761 (N_16761,N_14585,N_15816);
xor U16762 (N_16762,N_12916,N_12465);
or U16763 (N_16763,N_12053,N_15365);
and U16764 (N_16764,N_12748,N_14574);
or U16765 (N_16765,N_15031,N_14496);
nor U16766 (N_16766,N_12277,N_13953);
nand U16767 (N_16767,N_15127,N_15605);
or U16768 (N_16768,N_15927,N_13370);
nand U16769 (N_16769,N_15118,N_13466);
nand U16770 (N_16770,N_15440,N_12117);
xor U16771 (N_16771,N_15257,N_14774);
xnor U16772 (N_16772,N_14815,N_14721);
or U16773 (N_16773,N_14622,N_15267);
nor U16774 (N_16774,N_13529,N_12637);
or U16775 (N_16775,N_15033,N_15213);
nor U16776 (N_16776,N_13413,N_13314);
nor U16777 (N_16777,N_14422,N_14132);
xor U16778 (N_16778,N_13705,N_14148);
nand U16779 (N_16779,N_15823,N_15285);
xor U16780 (N_16780,N_13702,N_13776);
nand U16781 (N_16781,N_14001,N_15384);
and U16782 (N_16782,N_15691,N_13674);
or U16783 (N_16783,N_15465,N_14497);
or U16784 (N_16784,N_15356,N_12976);
nand U16785 (N_16785,N_14243,N_14683);
and U16786 (N_16786,N_13218,N_12314);
nor U16787 (N_16787,N_14136,N_14889);
nand U16788 (N_16788,N_13562,N_12663);
and U16789 (N_16789,N_12335,N_12904);
nand U16790 (N_16790,N_13830,N_15866);
xor U16791 (N_16791,N_15590,N_12691);
and U16792 (N_16792,N_12900,N_14668);
and U16793 (N_16793,N_15788,N_15379);
nand U16794 (N_16794,N_13931,N_14058);
and U16795 (N_16795,N_14169,N_15277);
nor U16796 (N_16796,N_14244,N_14776);
nor U16797 (N_16797,N_14285,N_14617);
nand U16798 (N_16798,N_12839,N_15043);
or U16799 (N_16799,N_12749,N_13242);
xnor U16800 (N_16800,N_14279,N_12924);
and U16801 (N_16801,N_12788,N_12144);
or U16802 (N_16802,N_12938,N_15179);
or U16803 (N_16803,N_15800,N_13460);
nand U16804 (N_16804,N_14030,N_15702);
nor U16805 (N_16805,N_14726,N_14527);
or U16806 (N_16806,N_14432,N_13573);
nand U16807 (N_16807,N_12629,N_14145);
or U16808 (N_16808,N_13168,N_13331);
xnor U16809 (N_16809,N_12309,N_14481);
or U16810 (N_16810,N_14261,N_13866);
nor U16811 (N_16811,N_12362,N_14528);
nand U16812 (N_16812,N_13288,N_15577);
xnor U16813 (N_16813,N_12963,N_15484);
and U16814 (N_16814,N_15881,N_14977);
xnor U16815 (N_16815,N_13633,N_13002);
or U16816 (N_16816,N_14494,N_15135);
or U16817 (N_16817,N_14516,N_14388);
nor U16818 (N_16818,N_14625,N_12161);
nor U16819 (N_16819,N_12812,N_14632);
and U16820 (N_16820,N_13570,N_12878);
and U16821 (N_16821,N_15124,N_14685);
nand U16822 (N_16822,N_14246,N_15869);
nor U16823 (N_16823,N_12486,N_14943);
and U16824 (N_16824,N_15651,N_12319);
or U16825 (N_16825,N_13363,N_14483);
or U16826 (N_16826,N_13282,N_14104);
xnor U16827 (N_16827,N_12167,N_13458);
and U16828 (N_16828,N_13913,N_14219);
or U16829 (N_16829,N_14092,N_13890);
or U16830 (N_16830,N_12816,N_14675);
or U16831 (N_16831,N_14262,N_12945);
nor U16832 (N_16832,N_12316,N_14401);
nand U16833 (N_16833,N_15071,N_13270);
and U16834 (N_16834,N_13754,N_14355);
nand U16835 (N_16835,N_13474,N_15467);
nor U16836 (N_16836,N_12253,N_13118);
and U16837 (N_16837,N_13516,N_14904);
nand U16838 (N_16838,N_15210,N_14642);
and U16839 (N_16839,N_13860,N_14323);
nand U16840 (N_16840,N_13307,N_15078);
and U16841 (N_16841,N_12006,N_15463);
or U16842 (N_16842,N_13898,N_12595);
and U16843 (N_16843,N_13299,N_12188);
or U16844 (N_16844,N_13303,N_14375);
nor U16845 (N_16845,N_13936,N_14320);
nor U16846 (N_16846,N_14439,N_12802);
nand U16847 (N_16847,N_13339,N_14443);
and U16848 (N_16848,N_15754,N_15981);
and U16849 (N_16849,N_14913,N_14521);
nor U16850 (N_16850,N_12364,N_13760);
and U16851 (N_16851,N_15394,N_14493);
nor U16852 (N_16852,N_13930,N_13457);
and U16853 (N_16853,N_12185,N_14164);
nand U16854 (N_16854,N_15612,N_12882);
and U16855 (N_16855,N_12894,N_13692);
and U16856 (N_16856,N_14384,N_15836);
and U16857 (N_16857,N_13641,N_13343);
xnor U16858 (N_16858,N_15513,N_12297);
and U16859 (N_16859,N_14700,N_14790);
and U16860 (N_16860,N_14042,N_12339);
nand U16861 (N_16861,N_13390,N_12917);
xor U16862 (N_16862,N_13126,N_14837);
and U16863 (N_16863,N_15497,N_13833);
xor U16864 (N_16864,N_14196,N_15893);
nand U16865 (N_16865,N_14336,N_13117);
or U16866 (N_16866,N_12978,N_14917);
and U16867 (N_16867,N_13492,N_13295);
nor U16868 (N_16868,N_12768,N_13517);
nand U16869 (N_16869,N_15032,N_13246);
and U16870 (N_16870,N_13816,N_14501);
and U16871 (N_16871,N_14266,N_14187);
nand U16872 (N_16872,N_13004,N_12672);
or U16873 (N_16873,N_13550,N_14288);
and U16874 (N_16874,N_13537,N_12594);
nand U16875 (N_16875,N_12641,N_14512);
or U16876 (N_16876,N_15499,N_13975);
nand U16877 (N_16877,N_14954,N_12238);
nor U16878 (N_16878,N_12538,N_13414);
or U16879 (N_16879,N_13030,N_13008);
xnor U16880 (N_16880,N_14149,N_15587);
or U16881 (N_16881,N_13487,N_15453);
nor U16882 (N_16882,N_15264,N_13949);
nor U16883 (N_16883,N_12278,N_14381);
nand U16884 (N_16884,N_14805,N_12642);
nor U16885 (N_16885,N_15991,N_12225);
nand U16886 (N_16886,N_13205,N_14593);
xor U16887 (N_16887,N_15299,N_15339);
nor U16888 (N_16888,N_13783,N_15801);
and U16889 (N_16889,N_12619,N_13130);
or U16890 (N_16890,N_12510,N_14062);
xor U16891 (N_16891,N_14584,N_13710);
xor U16892 (N_16892,N_15055,N_14389);
nor U16893 (N_16893,N_12449,N_14507);
and U16894 (N_16894,N_15827,N_13609);
nor U16895 (N_16895,N_13980,N_14181);
nand U16896 (N_16896,N_15200,N_13818);
nor U16897 (N_16897,N_14581,N_12125);
nor U16898 (N_16898,N_12344,N_12638);
and U16899 (N_16899,N_14660,N_13124);
nor U16900 (N_16900,N_13360,N_14398);
and U16901 (N_16901,N_12805,N_12995);
nand U16902 (N_16902,N_15361,N_12723);
and U16903 (N_16903,N_13826,N_15295);
nand U16904 (N_16904,N_13230,N_13172);
and U16905 (N_16905,N_14028,N_15976);
nor U16906 (N_16906,N_13110,N_15736);
nor U16907 (N_16907,N_15328,N_14515);
and U16908 (N_16908,N_13684,N_14052);
nor U16909 (N_16909,N_15928,N_12656);
nor U16910 (N_16910,N_15740,N_13682);
nor U16911 (N_16911,N_15230,N_12088);
and U16912 (N_16912,N_15496,N_12609);
nand U16913 (N_16913,N_13727,N_15087);
xnor U16914 (N_16914,N_13404,N_14611);
nor U16915 (N_16915,N_12308,N_12962);
nor U16916 (N_16916,N_15967,N_13361);
or U16917 (N_16917,N_14325,N_12038);
nor U16918 (N_16918,N_14655,N_14142);
nor U16919 (N_16919,N_13132,N_13612);
nor U16920 (N_16920,N_12396,N_12547);
nor U16921 (N_16921,N_13994,N_15721);
and U16922 (N_16922,N_13507,N_13903);
nor U16923 (N_16923,N_12775,N_15542);
nor U16924 (N_16924,N_14109,N_12577);
nand U16925 (N_16925,N_15029,N_13222);
nand U16926 (N_16926,N_12569,N_12758);
nor U16927 (N_16927,N_14032,N_13087);
or U16928 (N_16928,N_12921,N_12591);
nor U16929 (N_16929,N_14868,N_13896);
and U16930 (N_16930,N_13824,N_12694);
nor U16931 (N_16931,N_12555,N_13120);
and U16932 (N_16932,N_15370,N_13974);
or U16933 (N_16933,N_15666,N_15476);
nor U16934 (N_16934,N_12662,N_12094);
xnor U16935 (N_16935,N_14859,N_14881);
and U16936 (N_16936,N_14251,N_14555);
xor U16937 (N_16937,N_12392,N_14691);
or U16938 (N_16938,N_15142,N_12863);
nand U16939 (N_16939,N_12228,N_12433);
and U16940 (N_16940,N_14572,N_13134);
nor U16941 (N_16941,N_15131,N_12622);
or U16942 (N_16942,N_14312,N_15045);
or U16943 (N_16943,N_14666,N_15312);
nand U16944 (N_16944,N_15408,N_13864);
or U16945 (N_16945,N_14390,N_15524);
or U16946 (N_16946,N_14339,N_12665);
and U16947 (N_16947,N_15695,N_14820);
nor U16948 (N_16948,N_14467,N_14651);
nor U16949 (N_16949,N_12754,N_12227);
or U16950 (N_16950,N_15111,N_12854);
or U16951 (N_16951,N_12351,N_14407);
xnor U16952 (N_16952,N_15911,N_15656);
or U16953 (N_16953,N_14183,N_14926);
and U16954 (N_16954,N_15888,N_13358);
and U16955 (N_16955,N_15482,N_15167);
nor U16956 (N_16956,N_12806,N_13317);
nor U16957 (N_16957,N_15512,N_14361);
nor U16958 (N_16958,N_13922,N_15580);
xor U16959 (N_16959,N_13099,N_13627);
or U16960 (N_16960,N_14365,N_14176);
nand U16961 (N_16961,N_13902,N_13069);
or U16962 (N_16962,N_12936,N_14019);
nor U16963 (N_16963,N_14053,N_13531);
nand U16964 (N_16964,N_15262,N_15877);
or U16965 (N_16965,N_15790,N_15464);
xor U16966 (N_16966,N_12550,N_15185);
nand U16967 (N_16967,N_15341,N_12780);
or U16968 (N_16968,N_14737,N_13823);
or U16969 (N_16969,N_12865,N_15530);
nand U16970 (N_16970,N_15169,N_15081);
nand U16971 (N_16971,N_15166,N_14434);
nor U16972 (N_16972,N_15942,N_12121);
nand U16973 (N_16973,N_12113,N_14784);
nand U16974 (N_16974,N_15332,N_12628);
xnor U16975 (N_16975,N_15847,N_13525);
and U16976 (N_16976,N_14171,N_15700);
and U16977 (N_16977,N_14231,N_13751);
nor U16978 (N_16978,N_12275,N_12972);
nor U16979 (N_16979,N_12155,N_14874);
nand U16980 (N_16980,N_12110,N_13831);
or U16981 (N_16981,N_13601,N_15621);
nand U16982 (N_16982,N_12521,N_12307);
nand U16983 (N_16983,N_14121,N_15141);
and U16984 (N_16984,N_12890,N_14939);
or U16985 (N_16985,N_14801,N_14353);
or U16986 (N_16986,N_13225,N_12480);
nand U16987 (N_16987,N_14799,N_13428);
or U16988 (N_16988,N_15049,N_14411);
nand U16989 (N_16989,N_12367,N_14307);
and U16990 (N_16990,N_14645,N_14760);
nand U16991 (N_16991,N_15969,N_14013);
nor U16992 (N_16992,N_15739,N_12320);
nor U16993 (N_16993,N_12261,N_12967);
or U16994 (N_16994,N_13354,N_13216);
nor U16995 (N_16995,N_13014,N_15063);
and U16996 (N_16996,N_15475,N_12220);
and U16997 (N_16997,N_15423,N_14900);
nand U16998 (N_16998,N_14437,N_12453);
nor U16999 (N_16999,N_14690,N_12247);
nor U17000 (N_17000,N_15050,N_14007);
nand U17001 (N_17001,N_14095,N_13613);
or U17002 (N_17002,N_15217,N_13689);
and U17003 (N_17003,N_14821,N_12858);
and U17004 (N_17004,N_12385,N_13777);
nor U17005 (N_17005,N_12587,N_13638);
or U17006 (N_17006,N_14237,N_15232);
nor U17007 (N_17007,N_12254,N_12961);
nor U17008 (N_17008,N_14707,N_15805);
nand U17009 (N_17009,N_15272,N_14452);
and U17010 (N_17010,N_12393,N_12328);
nor U17011 (N_17011,N_12031,N_14114);
and U17012 (N_17012,N_15445,N_14853);
or U17013 (N_17013,N_12203,N_12164);
nand U17014 (N_17014,N_15932,N_13260);
nor U17015 (N_17015,N_12718,N_15568);
or U17016 (N_17016,N_15105,N_12880);
nor U17017 (N_17017,N_13555,N_15769);
nand U17018 (N_17018,N_13534,N_15274);
nor U17019 (N_17019,N_14455,N_14768);
or U17020 (N_17020,N_13377,N_12709);
nor U17021 (N_17021,N_12644,N_13240);
or U17022 (N_17022,N_14487,N_14739);
and U17023 (N_17023,N_15784,N_13966);
nor U17024 (N_17024,N_13791,N_14287);
nor U17025 (N_17025,N_13799,N_12919);
nor U17026 (N_17026,N_14552,N_15209);
nand U17027 (N_17027,N_13151,N_15261);
and U17028 (N_17028,N_14765,N_15654);
nand U17029 (N_17029,N_15258,N_13970);
xnor U17030 (N_17030,N_13885,N_12509);
nor U17031 (N_17031,N_12977,N_14659);
nor U17032 (N_17032,N_13292,N_15554);
and U17033 (N_17033,N_13841,N_12299);
xnor U17034 (N_17034,N_12757,N_13464);
xor U17035 (N_17035,N_13011,N_14624);
and U17036 (N_17036,N_15741,N_13455);
or U17037 (N_17037,N_14924,N_15965);
xnor U17038 (N_17038,N_15751,N_12310);
or U17039 (N_17039,N_15617,N_15910);
and U17040 (N_17040,N_12082,N_13244);
or U17041 (N_17041,N_13108,N_14255);
nor U17042 (N_17042,N_14665,N_12870);
or U17043 (N_17043,N_15377,N_15680);
and U17044 (N_17044,N_14936,N_14023);
nor U17045 (N_17045,N_14412,N_14147);
and U17046 (N_17046,N_15833,N_13194);
or U17047 (N_17047,N_15279,N_15834);
nand U17048 (N_17048,N_13769,N_15123);
or U17049 (N_17049,N_15882,N_12744);
and U17050 (N_17050,N_15330,N_13906);
and U17051 (N_17051,N_13353,N_12682);
nand U17052 (N_17052,N_12483,N_15470);
nand U17053 (N_17053,N_12523,N_13207);
xor U17054 (N_17054,N_15304,N_12896);
nor U17055 (N_17055,N_13235,N_14713);
or U17056 (N_17056,N_12257,N_14076);
xor U17057 (N_17057,N_12895,N_14741);
nand U17058 (N_17058,N_13551,N_14968);
nor U17059 (N_17059,N_12915,N_12811);
nand U17060 (N_17060,N_15357,N_13504);
nand U17061 (N_17061,N_13597,N_12338);
nor U17062 (N_17062,N_15348,N_15494);
xor U17063 (N_17063,N_12840,N_15732);
and U17064 (N_17064,N_13443,N_14254);
nand U17065 (N_17065,N_12057,N_14226);
xnor U17066 (N_17066,N_12030,N_14470);
nand U17067 (N_17067,N_13586,N_12477);
nand U17068 (N_17068,N_12395,N_12241);
or U17069 (N_17069,N_15061,N_13819);
or U17070 (N_17070,N_14009,N_12200);
or U17071 (N_17071,N_14186,N_12263);
nand U17072 (N_17072,N_12495,N_12527);
xor U17073 (N_17073,N_12763,N_14742);
xnor U17074 (N_17074,N_13111,N_14973);
and U17075 (N_17075,N_15812,N_13212);
nor U17076 (N_17076,N_13732,N_12348);
or U17077 (N_17077,N_15844,N_12271);
nand U17078 (N_17078,N_13267,N_14664);
or U17079 (N_17079,N_13524,N_15164);
nor U17080 (N_17080,N_15437,N_14350);
or U17081 (N_17081,N_15820,N_15308);
and U17082 (N_17082,N_12909,N_13725);
nor U17083 (N_17083,N_12294,N_15092);
nor U17084 (N_17084,N_13622,N_15426);
nand U17085 (N_17085,N_13368,N_12646);
and U17086 (N_17086,N_13887,N_15616);
nand U17087 (N_17087,N_12798,N_12968);
nand U17088 (N_17088,N_13670,N_13828);
and U17089 (N_17089,N_13296,N_13519);
or U17090 (N_17090,N_13979,N_14912);
xnor U17091 (N_17091,N_15250,N_13263);
or U17092 (N_17092,N_15090,N_15566);
and U17093 (N_17093,N_15316,N_15602);
nor U17094 (N_17094,N_13579,N_13765);
nor U17095 (N_17095,N_12426,N_12173);
nand U17096 (N_17096,N_14127,N_14075);
nand U17097 (N_17097,N_12843,N_12513);
nor U17098 (N_17098,N_13236,N_12661);
and U17099 (N_17099,N_15114,N_14796);
or U17100 (N_17100,N_15198,N_14094);
nor U17101 (N_17101,N_14444,N_12952);
and U17102 (N_17102,N_13444,N_12987);
xnor U17103 (N_17103,N_12054,N_14532);
and U17104 (N_17104,N_15538,N_13789);
nand U17105 (N_17105,N_12143,N_12296);
or U17106 (N_17106,N_14579,N_13628);
and U17107 (N_17107,N_12284,N_12605);
or U17108 (N_17108,N_13306,N_15180);
nand U17109 (N_17109,N_12470,N_14671);
nand U17110 (N_17110,N_12590,N_15346);
xor U17111 (N_17111,N_15241,N_14499);
and U17112 (N_17112,N_13265,N_12746);
nand U17113 (N_17113,N_13115,N_14872);
nand U17114 (N_17114,N_14778,N_15231);
nor U17115 (N_17115,N_12715,N_12522);
and U17116 (N_17116,N_14272,N_14902);
nor U17117 (N_17117,N_14570,N_13502);
xor U17118 (N_17118,N_12131,N_12561);
nor U17119 (N_17119,N_14057,N_14441);
nand U17120 (N_17120,N_13723,N_14591);
and U17121 (N_17121,N_15533,N_15159);
or U17122 (N_17122,N_14608,N_13310);
and U17123 (N_17123,N_14630,N_15502);
nor U17124 (N_17124,N_12492,N_12455);
nand U17125 (N_17125,N_13714,N_14283);
nand U17126 (N_17126,N_15110,N_14438);
nor U17127 (N_17127,N_13056,N_15717);
and U17128 (N_17128,N_12821,N_14461);
nand U17129 (N_17129,N_13364,N_14151);
nor U17130 (N_17130,N_15404,N_15227);
and U17131 (N_17131,N_15314,N_15238);
nand U17132 (N_17132,N_14034,N_13261);
nor U17133 (N_17133,N_14351,N_15212);
xnor U17134 (N_17134,N_12971,N_13203);
or U17135 (N_17135,N_12845,N_15917);
or U17136 (N_17136,N_12199,N_12411);
xor U17137 (N_17137,N_13275,N_13874);
nand U17138 (N_17138,N_15523,N_15144);
or U17139 (N_17139,N_13122,N_15146);
nand U17140 (N_17140,N_14847,N_14413);
nor U17141 (N_17141,N_14711,N_13342);
and U17142 (N_17142,N_15398,N_15775);
and U17143 (N_17143,N_15531,N_13595);
nand U17144 (N_17144,N_12828,N_15493);
or U17145 (N_17145,N_12681,N_15392);
or U17146 (N_17146,N_13762,N_15431);
nand U17147 (N_17147,N_12892,N_12074);
nand U17148 (N_17148,N_15256,N_14514);
nor U17149 (N_17149,N_13034,N_14157);
nor U17150 (N_17150,N_14969,N_12388);
nor U17151 (N_17151,N_14772,N_15563);
nand U17152 (N_17152,N_12002,N_15615);
nor U17153 (N_17153,N_13393,N_15068);
nor U17154 (N_17154,N_15326,N_15676);
nand U17155 (N_17155,N_12290,N_14942);
xor U17156 (N_17156,N_15517,N_13768);
and U17157 (N_17157,N_13647,N_15485);
nand U17158 (N_17158,N_15735,N_13071);
or U17159 (N_17159,N_14426,N_15623);
and U17160 (N_17160,N_12224,N_13382);
nor U17161 (N_17161,N_12585,N_15372);
xnor U17162 (N_17162,N_13856,N_12720);
and U17163 (N_17163,N_14330,N_14595);
nand U17164 (N_17164,N_15575,N_13486);
and U17165 (N_17165,N_12221,N_13653);
or U17166 (N_17166,N_14793,N_12403);
nand U17167 (N_17167,N_13336,N_14849);
or U17168 (N_17168,N_13701,N_12934);
or U17169 (N_17169,N_12268,N_12304);
and U17170 (N_17170,N_13755,N_14653);
nand U17171 (N_17171,N_13150,N_13145);
nor U17172 (N_17172,N_14971,N_14400);
and U17173 (N_17173,N_13563,N_12767);
nand U17174 (N_17174,N_14657,N_12163);
or U17175 (N_17175,N_14344,N_13431);
nor U17176 (N_17176,N_13408,N_14322);
nand U17177 (N_17177,N_15375,N_12108);
nand U17178 (N_17178,N_15362,N_14757);
and U17179 (N_17179,N_13503,N_15980);
or U17180 (N_17180,N_13085,N_13199);
nor U17181 (N_17181,N_15027,N_13171);
nor U17182 (N_17182,N_13698,N_12699);
nand U17183 (N_17183,N_14458,N_14141);
xor U17184 (N_17184,N_14730,N_14368);
nor U17185 (N_17185,N_13147,N_12343);
nand U17186 (N_17186,N_15915,N_14024);
xnor U17187 (N_17187,N_15439,N_13022);
and U17188 (N_17188,N_14370,N_15609);
xor U17189 (N_17189,N_14738,N_15428);
or U17190 (N_17190,N_13423,N_15780);
nor U17191 (N_17191,N_13667,N_13272);
or U17192 (N_17192,N_15696,N_13640);
or U17193 (N_17193,N_14005,N_12583);
nand U17194 (N_17194,N_14761,N_15374);
and U17195 (N_17195,N_12429,N_13935);
and U17196 (N_17196,N_15507,N_12783);
and U17197 (N_17197,N_15501,N_14174);
nor U17198 (N_17198,N_12184,N_14295);
or U17199 (N_17199,N_12991,N_13061);
nand U17200 (N_17200,N_14869,N_12514);
or U17201 (N_17201,N_13671,N_14055);
and U17202 (N_17202,N_15966,N_13802);
and U17203 (N_17203,N_13759,N_12126);
nand U17204 (N_17204,N_12052,N_12958);
nand U17205 (N_17205,N_13719,N_14728);
and U17206 (N_17206,N_12764,N_15168);
and U17207 (N_17207,N_13988,N_13023);
nand U17208 (N_17208,N_14209,N_15469);
nor U17209 (N_17209,N_13077,N_13309);
nand U17210 (N_17210,N_14167,N_13286);
or U17211 (N_17211,N_14328,N_13559);
or U17212 (N_17212,N_13659,N_13790);
nand U17213 (N_17213,N_14717,N_14860);
and U17214 (N_17214,N_13178,N_14367);
nand U17215 (N_17215,N_12440,N_13454);
nand U17216 (N_17216,N_15260,N_14326);
or U17217 (N_17217,N_12152,N_14899);
nand U17218 (N_17218,N_15221,N_14892);
or U17219 (N_17219,N_12626,N_15223);
nor U17220 (N_17220,N_12059,N_12776);
and U17221 (N_17221,N_15955,N_15681);
or U17222 (N_17222,N_13070,N_15478);
and U17223 (N_17223,N_14454,N_12372);
nand U17224 (N_17224,N_15935,N_15222);
nand U17225 (N_17225,N_13213,N_12265);
or U17226 (N_17226,N_14362,N_12177);
nand U17227 (N_17227,N_13614,N_12169);
nand U17228 (N_17228,N_13527,N_15887);
and U17229 (N_17229,N_15075,N_14696);
nor U17230 (N_17230,N_12235,N_12093);
xnor U17231 (N_17231,N_14641,N_15053);
or U17232 (N_17232,N_13290,N_13683);
nor U17233 (N_17233,N_14716,N_13876);
and U17234 (N_17234,N_12166,N_14974);
xor U17235 (N_17235,N_12256,N_13067);
or U17236 (N_17236,N_14018,N_12134);
xnor U17237 (N_17237,N_12625,N_12427);
and U17238 (N_17238,N_15874,N_13341);
nor U17239 (N_17239,N_13254,N_14858);
nand U17240 (N_17240,N_15207,N_14703);
or U17241 (N_17241,N_13750,N_14269);
and U17242 (N_17242,N_12413,N_14822);
xor U17243 (N_17243,N_14173,N_13693);
nor U17244 (N_17244,N_15098,N_14754);
and U17245 (N_17245,N_12130,N_12406);
or U17246 (N_17246,N_13082,N_14216);
nor U17247 (N_17247,N_15364,N_14699);
nand U17248 (N_17248,N_15798,N_12508);
and U17249 (N_17249,N_13899,N_14435);
and U17250 (N_17250,N_13221,N_14539);
nand U17251 (N_17251,N_14035,N_14766);
or U17252 (N_17252,N_12463,N_12677);
or U17253 (N_17253,N_14662,N_14338);
nand U17254 (N_17254,N_12467,N_12586);
and U17255 (N_17255,N_14809,N_15644);
or U17256 (N_17256,N_12048,N_13359);
or U17257 (N_17257,N_13927,N_14875);
nand U17258 (N_17258,N_13726,N_14016);
and U17259 (N_17259,N_14540,N_12149);
nand U17260 (N_17260,N_12493,N_15782);
nor U17261 (N_17261,N_15986,N_12459);
nor U17262 (N_17262,N_15515,N_15675);
nor U17263 (N_17263,N_14724,N_15344);
xor U17264 (N_17264,N_12755,N_12264);
nor U17265 (N_17265,N_12334,N_12956);
and U17266 (N_17266,N_13346,N_15013);
or U17267 (N_17267,N_12369,N_15839);
and U17268 (N_17268,N_12325,N_15175);
or U17269 (N_17269,N_13439,N_15406);
or U17270 (N_17270,N_13998,N_15737);
xnor U17271 (N_17271,N_14932,N_12850);
nand U17272 (N_17272,N_15864,N_12809);
or U17273 (N_17273,N_14277,N_12353);
nand U17274 (N_17274,N_15909,N_14382);
nor U17275 (N_17275,N_14951,N_13324);
and U17276 (N_17276,N_13610,N_14096);
nor U17277 (N_17277,N_14965,N_13676);
or U17278 (N_17278,N_13032,N_15352);
and U17279 (N_17279,N_13434,N_12487);
nor U17280 (N_17280,N_15219,N_14966);
xor U17281 (N_17281,N_13076,N_15726);
and U17282 (N_17282,N_15897,N_14543);
or U17283 (N_17283,N_13646,N_15886);
nand U17284 (N_17284,N_15526,N_14582);
and U17285 (N_17285,N_15889,N_12679);
and U17286 (N_17286,N_15102,N_14144);
nand U17287 (N_17287,N_12439,N_13164);
nor U17288 (N_17288,N_13713,N_12786);
nand U17289 (N_17289,N_12512,N_12939);
nand U17290 (N_17290,N_13845,N_15488);
and U17291 (N_17291,N_14911,N_12931);
nor U17292 (N_17292,N_13433,N_14846);
or U17293 (N_17293,N_12537,N_12889);
nor U17294 (N_17294,N_12137,N_14883);
nand U17295 (N_17295,N_15369,N_14380);
nor U17296 (N_17296,N_12330,N_15077);
or U17297 (N_17297,N_12004,N_14854);
and U17298 (N_17298,N_12905,N_13323);
or U17299 (N_17299,N_15776,N_12795);
and U17300 (N_17300,N_14541,N_14522);
and U17301 (N_17301,N_12898,N_13855);
nor U17302 (N_17302,N_15100,N_14867);
and U17303 (N_17303,N_14681,N_15367);
and U17304 (N_17304,N_15422,N_12906);
nor U17305 (N_17305,N_13277,N_12581);
nor U17306 (N_17306,N_14946,N_13636);
nor U17307 (N_17307,N_14313,N_13937);
xnor U17308 (N_17308,N_13801,N_15973);
nor U17309 (N_17309,N_12996,N_13392);
nor U17310 (N_17310,N_13010,N_15810);
and U17311 (N_17311,N_14798,N_14592);
and U17312 (N_17312,N_13624,N_12946);
or U17313 (N_17313,N_14862,N_13420);
nand U17314 (N_17314,N_14628,N_14836);
or U17315 (N_17315,N_15903,N_13062);
or U17316 (N_17316,N_15824,N_14701);
nor U17317 (N_17317,N_14221,N_12690);
nand U17318 (N_17318,N_12515,N_14402);
nand U17319 (N_17319,N_12539,N_14280);
or U17320 (N_17320,N_12035,N_12589);
nand U17321 (N_17321,N_12019,N_15992);
nand U17322 (N_17322,N_12765,N_13859);
nand U17323 (N_17323,N_13772,N_13499);
or U17324 (N_17324,N_15860,N_15303);
or U17325 (N_17325,N_12326,N_12380);
nor U17326 (N_17326,N_15290,N_13068);
nand U17327 (N_17327,N_13608,N_15017);
and U17328 (N_17328,N_14856,N_14366);
or U17329 (N_17329,N_15319,N_12260);
or U17330 (N_17330,N_12240,N_13895);
nand U17331 (N_17331,N_15188,N_12974);
or U17332 (N_17332,N_12654,N_14934);
nor U17333 (N_17333,N_15821,N_14125);
or U17334 (N_17334,N_14012,N_12077);
and U17335 (N_17335,N_13991,N_13104);
nand U17336 (N_17336,N_14294,N_14547);
xor U17337 (N_17337,N_14357,N_14898);
nand U17338 (N_17338,N_15306,N_14789);
or U17339 (N_17339,N_13029,N_14614);
nand U17340 (N_17340,N_13012,N_14864);
or U17341 (N_17341,N_15630,N_13631);
and U17342 (N_17342,N_15586,N_13740);
xnor U17343 (N_17343,N_12104,N_14008);
nand U17344 (N_17344,N_15640,N_14568);
or U17345 (N_17345,N_15793,N_14465);
xnor U17346 (N_17346,N_15753,N_15795);
nor U17347 (N_17347,N_15435,N_13162);
or U17348 (N_17348,N_15259,N_15841);
xnor U17349 (N_17349,N_15117,N_12701);
nand U17350 (N_17350,N_12796,N_13264);
nand U17351 (N_17351,N_13480,N_12881);
and U17352 (N_17352,N_15559,N_12416);
nand U17353 (N_17353,N_14371,N_13561);
xor U17354 (N_17354,N_12997,N_12132);
nand U17355 (N_17355,N_14915,N_15432);
or U17356 (N_17356,N_14735,N_14405);
or U17357 (N_17357,N_14960,N_13496);
nor U17358 (N_17358,N_14549,N_13582);
nor U17359 (N_17359,N_15597,N_13892);
and U17360 (N_17360,N_13208,N_14542);
xnor U17361 (N_17361,N_13851,N_14706);
xor U17362 (N_17362,N_15165,N_14684);
nand U17363 (N_17363,N_13987,N_15520);
and U17364 (N_17364,N_15796,N_15920);
nor U17365 (N_17365,N_15201,N_14271);
nor U17366 (N_17366,N_13192,N_14118);
xor U17367 (N_17367,N_12252,N_15106);
nand U17368 (N_17368,N_15653,N_14048);
xnor U17369 (N_17369,N_15473,N_15908);
and U17370 (N_17370,N_13251,N_15225);
xor U17371 (N_17371,N_15773,N_13695);
or U17372 (N_17372,N_15764,N_15089);
and U17373 (N_17373,N_15709,N_14673);
nor U17374 (N_17374,N_12079,N_13007);
or U17375 (N_17375,N_13113,N_12519);
nand U17376 (N_17376,N_12970,N_14081);
nor U17377 (N_17377,N_14228,N_14844);
nor U17378 (N_17378,N_15126,N_14331);
and U17379 (N_17379,N_12321,N_12992);
or U17380 (N_17380,N_12195,N_15310);
xnor U17381 (N_17381,N_13803,N_14085);
and U17382 (N_17382,N_15113,N_12673);
or U17383 (N_17383,N_14816,N_13850);
and U17384 (N_17384,N_13383,N_15953);
nor U17385 (N_17385,N_13989,N_14031);
and U17386 (N_17386,N_15545,N_15403);
nor U17387 (N_17387,N_14395,N_13548);
nand U17388 (N_17388,N_13355,N_12352);
nor U17389 (N_17389,N_14504,N_15109);
and U17390 (N_17390,N_12841,N_15088);
or U17391 (N_17391,N_12029,N_14479);
nand U17392 (N_17392,N_14376,N_12078);
or U17393 (N_17393,N_13441,N_12128);
nor U17394 (N_17394,N_13438,N_14377);
nand U17395 (N_17395,N_12313,N_14884);
or U17396 (N_17396,N_14580,N_15342);
nand U17397 (N_17397,N_12115,N_13316);
nor U17398 (N_17398,N_15416,N_13590);
nor U17399 (N_17399,N_14327,N_15327);
nor U17400 (N_17400,N_15946,N_12170);
nor U17401 (N_17401,N_12833,N_15284);
or U17402 (N_17402,N_15070,N_13462);
nand U17403 (N_17403,N_13080,N_13867);
and U17404 (N_17404,N_12669,N_13844);
nand U17405 (N_17405,N_12026,N_13871);
nand U17406 (N_17406,N_14301,N_13091);
nand U17407 (N_17407,N_15480,N_13078);
or U17408 (N_17408,N_14833,N_13006);
nand U17409 (N_17409,N_13526,N_14297);
xor U17410 (N_17410,N_15828,N_13552);
nand U17411 (N_17411,N_13345,N_14408);
nor U17412 (N_17412,N_13271,N_14195);
and U17413 (N_17413,N_12856,N_14694);
and U17414 (N_17414,N_13367,N_15689);
or U17415 (N_17415,N_12456,N_15156);
or U17416 (N_17416,N_14124,N_14207);
nor U17417 (N_17417,N_13528,N_14414);
nand U17418 (N_17418,N_12608,N_15382);
and U17419 (N_17419,N_13389,N_13733);
xnor U17420 (N_17420,N_14268,N_15211);
nor U17421 (N_17421,N_13965,N_12731);
nor U17422 (N_17422,N_15378,N_14235);
nand U17423 (N_17423,N_14089,N_14959);
nor U17424 (N_17424,N_13703,N_14644);
nor U17425 (N_17425,N_12771,N_13046);
xnor U17426 (N_17426,N_13604,N_13066);
nor U17427 (N_17427,N_13472,N_12739);
xnor U17428 (N_17428,N_15173,N_15282);
xnor U17429 (N_17429,N_15254,N_12965);
or U17430 (N_17430,N_13535,N_14702);
or U17431 (N_17431,N_13681,N_14200);
nand U17432 (N_17432,N_15421,N_15581);
nor U17433 (N_17433,N_15278,N_14425);
nor U17434 (N_17434,N_13607,N_14154);
and U17435 (N_17435,N_15968,N_12156);
nand U17436 (N_17436,N_12912,N_15214);
nand U17437 (N_17437,N_15811,N_12910);
and U17438 (N_17438,N_15539,N_15074);
nand U17439 (N_17439,N_14290,N_15044);
or U17440 (N_17440,N_12472,N_14409);
nand U17441 (N_17441,N_15035,N_15354);
or U17442 (N_17442,N_15937,N_15265);
nand U17443 (N_17443,N_12932,N_13611);
or U17444 (N_17444,N_15218,N_15851);
or U17445 (N_17445,N_15627,N_14072);
and U17446 (N_17446,N_15703,N_14871);
nand U17447 (N_17447,N_14253,N_12217);
xor U17448 (N_17448,N_15923,N_14044);
nand U17449 (N_17449,N_13901,N_13273);
nand U17450 (N_17450,N_12460,N_12432);
or U17451 (N_17451,N_13156,N_13266);
nand U17452 (N_17452,N_14745,N_13625);
nand U17453 (N_17453,N_12907,N_14802);
nand U17454 (N_17454,N_13939,N_15293);
nand U17455 (N_17455,N_12266,N_15729);
and U17456 (N_17456,N_12668,N_12062);
or U17457 (N_17457,N_15139,N_14559);
or U17458 (N_17458,N_12616,N_13257);
nand U17459 (N_17459,N_14909,N_12488);
or U17460 (N_17460,N_14637,N_12507);
and U17461 (N_17461,N_14083,N_12574);
and U17462 (N_17462,N_15671,N_14607);
and U17463 (N_17463,N_14613,N_13371);
nand U17464 (N_17464,N_15569,N_14067);
or U17465 (N_17465,N_15057,N_12729);
nor U17466 (N_17466,N_14410,N_15896);
or U17467 (N_17467,N_15430,N_15091);
or U17468 (N_17468,N_14276,N_15028);
nand U17469 (N_17469,N_14586,N_14817);
and U17470 (N_17470,N_15725,N_13925);
and U17471 (N_17471,N_15323,N_15560);
nand U17472 (N_17472,N_15765,N_12457);
xor U17473 (N_17473,N_15358,N_14550);
or U17474 (N_17474,N_13635,N_12565);
nand U17475 (N_17475,N_15748,N_13900);
and U17476 (N_17476,N_14180,N_14227);
nand U17477 (N_17477,N_15876,N_15410);
and U17478 (N_17478,N_12706,N_14140);
and U17479 (N_17479,N_12505,N_12204);
and U17480 (N_17480,N_15716,N_13181);
nor U17481 (N_17481,N_13379,N_12913);
nor U17482 (N_17482,N_15042,N_12835);
nor U17483 (N_17483,N_15433,N_14544);
nand U17484 (N_17484,N_13133,N_12666);
or U17485 (N_17485,N_15822,N_14705);
nor U17486 (N_17486,N_12248,N_14885);
nand U17487 (N_17487,N_14369,N_14126);
and U17488 (N_17488,N_14640,N_15309);
nand U17489 (N_17489,N_12707,N_14387);
nand U17490 (N_17490,N_14777,N_13148);
nand U17491 (N_17491,N_13259,N_14431);
nor U17492 (N_17492,N_14074,N_15191);
or U17493 (N_17493,N_12986,N_15483);
and U17494 (N_17494,N_13832,N_15945);
and U17495 (N_17495,N_12400,N_14785);
nor U17496 (N_17496,N_14910,N_14391);
or U17497 (N_17497,N_15046,N_15301);
or U17498 (N_17498,N_13877,N_13779);
xor U17499 (N_17499,N_14354,N_15668);
or U17500 (N_17500,N_14679,N_15610);
or U17501 (N_17501,N_14886,N_15056);
nand U17502 (N_17502,N_12355,N_13144);
and U17503 (N_17503,N_15396,N_13741);
xnor U17504 (N_17504,N_15192,N_13746);
or U17505 (N_17505,N_14589,N_13048);
and U17506 (N_17506,N_15051,N_15172);
nand U17507 (N_17507,N_15961,N_13280);
nand U17508 (N_17508,N_15951,N_13206);
and U17509 (N_17509,N_15419,N_14520);
nor U17510 (N_17510,N_14004,N_14972);
nor U17511 (N_17511,N_13180,N_13825);
nor U17512 (N_17512,N_14676,N_12374);
nor U17513 (N_17513,N_15919,N_12837);
or U17514 (N_17514,N_13304,N_13967);
and U17515 (N_17515,N_15528,N_12959);
nor U17516 (N_17516,N_14610,N_12683);
nor U17517 (N_17517,N_15325,N_15848);
nor U17518 (N_17518,N_15592,N_13227);
or U17519 (N_17519,N_14175,N_13724);
or U17520 (N_17520,N_12551,N_13211);
or U17521 (N_17521,N_13731,N_14385);
and U17522 (N_17522,N_15921,N_15519);
or U17523 (N_17523,N_12540,N_14594);
and U17524 (N_17524,N_14047,N_12820);
and U17525 (N_17525,N_12886,N_12051);
or U17526 (N_17526,N_15724,N_14229);
or U17527 (N_17527,N_13477,N_13442);
xor U17528 (N_17528,N_14182,N_14609);
nand U17529 (N_17529,N_12443,N_12503);
nor U17530 (N_17530,N_15984,N_14961);
nor U17531 (N_17531,N_15646,N_12171);
and U17532 (N_17532,N_13445,N_15756);
or U17533 (N_17533,N_14098,N_13857);
nand U17534 (N_17534,N_13166,N_14600);
nor U17535 (N_17535,N_12627,N_13155);
or U17536 (N_17536,N_13643,N_12154);
nand U17537 (N_17537,N_14451,N_14852);
nand U17538 (N_17538,N_15537,N_15974);
xnor U17539 (N_17539,N_14931,N_12530);
or U17540 (N_17540,N_13854,N_15487);
nor U17541 (N_17541,N_14335,N_12109);
and U17542 (N_17542,N_15383,N_13278);
or U17543 (N_17543,N_15405,N_12929);
nor U17544 (N_17544,N_13175,N_14813);
or U17545 (N_17545,N_14346,N_12901);
nand U17546 (N_17546,N_15409,N_12182);
xor U17547 (N_17547,N_12851,N_13565);
nor U17548 (N_17548,N_12797,N_12603);
nor U17549 (N_17549,N_13321,N_13728);
nand U17550 (N_17550,N_14667,N_14530);
nand U17551 (N_17551,N_13675,N_12107);
and U17552 (N_17552,N_15655,N_13753);
and U17553 (N_17553,N_12491,N_14252);
nand U17554 (N_17554,N_15988,N_15313);
nand U17555 (N_17555,N_15244,N_14863);
nand U17556 (N_17556,N_15253,N_14463);
xnor U17557 (N_17557,N_14620,N_12719);
or U17558 (N_17558,N_12536,N_15130);
nand U17559 (N_17559,N_15333,N_13184);
nand U17560 (N_17560,N_13491,N_13541);
nand U17561 (N_17561,N_13581,N_13533);
xor U17562 (N_17562,N_13083,N_13648);
nand U17563 (N_17563,N_12375,N_14054);
or U17564 (N_17564,N_12056,N_12490);
nor U17565 (N_17565,N_12468,N_13805);
nand U17566 (N_17566,N_13169,N_15963);
and U17567 (N_17567,N_15170,N_12045);
nor U17568 (N_17568,N_12340,N_14788);
nand U17569 (N_17569,N_13125,N_12068);
nand U17570 (N_17570,N_15929,N_13811);
nor U17571 (N_17571,N_13497,N_15594);
nor U17572 (N_17572,N_13334,N_14333);
nor U17573 (N_17573,N_13365,N_15572);
or U17574 (N_17574,N_13198,N_14184);
and U17575 (N_17575,N_13042,N_14631);
nor U17576 (N_17576,N_14417,N_12237);
nor U17577 (N_17577,N_14404,N_12908);
nor U17578 (N_17578,N_15018,N_12826);
and U17579 (N_17579,N_12270,N_15468);
xor U17580 (N_17580,N_12462,N_13928);
nand U17581 (N_17581,N_14780,N_12849);
nand U17582 (N_17582,N_13685,N_13820);
xor U17583 (N_17583,N_15162,N_15206);
or U17584 (N_17584,N_12973,N_13947);
xor U17585 (N_17585,N_13058,N_15034);
nand U17586 (N_17586,N_14999,N_15543);
nand U17587 (N_17587,N_12651,N_14895);
and U17588 (N_17588,N_13394,N_12743);
nand U17589 (N_17589,N_14534,N_13598);
nor U17590 (N_17590,N_15376,N_13167);
nor U17591 (N_17591,N_15585,N_13510);
nor U17592 (N_17592,N_14137,N_15574);
or U17593 (N_17593,N_14217,N_12444);
nand U17594 (N_17594,N_13284,N_14567);
xor U17595 (N_17595,N_15145,N_13511);
or U17596 (N_17596,N_14672,N_12928);
nand U17597 (N_17597,N_14222,N_13650);
and U17598 (N_17598,N_12230,N_15645);
or U17599 (N_17599,N_15629,N_13669);
nand U17600 (N_17600,N_15119,N_15959);
or U17601 (N_17601,N_12689,N_12728);
and U17602 (N_17602,N_14753,N_15620);
and U17603 (N_17603,N_15770,N_12085);
and U17604 (N_17604,N_14947,N_12613);
and U17605 (N_17605,N_15368,N_14143);
and U17606 (N_17606,N_13665,N_13822);
nand U17607 (N_17607,N_14621,N_13808);
or U17608 (N_17608,N_13258,N_15060);
and U17609 (N_17609,N_15318,N_14002);
or U17610 (N_17610,N_13663,N_12322);
nor U17611 (N_17611,N_15693,N_15701);
nor U17612 (N_17612,N_12408,N_15134);
nor U17613 (N_17613,N_14310,N_13163);
or U17614 (N_17614,N_13742,N_12567);
and U17615 (N_17615,N_14314,N_14759);
or U17616 (N_17616,N_13881,N_12923);
xor U17617 (N_17617,N_15723,N_12272);
and U17618 (N_17618,N_12176,N_13074);
nor U17619 (N_17619,N_13512,N_15947);
nand U17620 (N_17620,N_13576,N_14318);
nor U17621 (N_17621,N_13362,N_13948);
and U17622 (N_17622,N_13761,N_15181);
nand U17623 (N_17623,N_12289,N_15845);
or U17624 (N_17624,N_12911,N_14634);
nand U17625 (N_17625,N_14981,N_12189);
nand U17626 (N_17626,N_12280,N_15710);
nand U17627 (N_17627,N_15500,N_14220);
or U17628 (N_17628,N_15104,N_15003);
nand U17629 (N_17629,N_13224,N_13494);
nor U17630 (N_17630,N_13757,N_14419);
nor U17631 (N_17631,N_15015,N_13059);
nand U17632 (N_17632,N_14165,N_13247);
nor U17633 (N_17633,N_13972,N_14824);
nor U17634 (N_17634,N_12502,N_15781);
or U17635 (N_17635,N_15636,N_15846);
nor U17636 (N_17636,N_14039,N_13810);
nand U17637 (N_17637,N_13941,N_15643);
xor U17638 (N_17638,N_12612,N_12011);
and U17639 (N_17639,N_15125,N_12446);
nand U17640 (N_17640,N_12158,N_15189);
nor U17641 (N_17641,N_15006,N_13137);
xnor U17642 (N_17642,N_13817,N_13141);
xnor U17643 (N_17643,N_14436,N_14800);
and U17644 (N_17644,N_15171,N_12687);
nand U17645 (N_17645,N_15611,N_13637);
and U17646 (N_17646,N_13568,N_14208);
nor U17647 (N_17647,N_13587,N_12291);
nand U17648 (N_17648,N_14061,N_12774);
xor U17649 (N_17649,N_15772,N_13055);
and U17650 (N_17650,N_15583,N_14604);
xor U17651 (N_17651,N_12529,N_13470);
xnor U17652 (N_17652,N_12800,N_15182);
nor U17653 (N_17653,N_14020,N_15711);
or U17654 (N_17654,N_12617,N_14373);
and U17655 (N_17655,N_13019,N_15939);
or U17656 (N_17656,N_15289,N_13748);
or U17657 (N_17657,N_12823,N_13170);
xor U17658 (N_17658,N_12324,N_14260);
nand U17659 (N_17659,N_14027,N_13787);
and U17660 (N_17660,N_14230,N_12777);
and U17661 (N_17661,N_12579,N_13718);
nor U17662 (N_17662,N_12370,N_15420);
and U17663 (N_17663,N_13424,N_13468);
nor U17664 (N_17664,N_15442,N_15148);
nor U17665 (N_17665,N_15661,N_13101);
or U17666 (N_17666,N_12571,N_13097);
nor U17667 (N_17667,N_15914,N_15425);
xor U17668 (N_17668,N_13302,N_13770);
or U17669 (N_17669,N_14406,N_15263);
and U17670 (N_17670,N_15466,N_12822);
and U17671 (N_17671,N_13963,N_12548);
xor U17672 (N_17672,N_15564,N_12877);
or U17673 (N_17673,N_14962,N_13798);
and U17674 (N_17674,N_15116,N_12827);
nand U17675 (N_17675,N_13451,N_13958);
nor U17676 (N_17676,N_15806,N_15140);
nor U17677 (N_17677,N_13978,N_14304);
nand U17678 (N_17678,N_13300,N_15321);
and U17679 (N_17679,N_14850,N_13398);
nor U17680 (N_17680,N_13033,N_14839);
and U17681 (N_17681,N_15817,N_12785);
and U17682 (N_17682,N_14289,N_12172);
nor U17683 (N_17683,N_13399,N_14818);
nor U17684 (N_17684,N_15516,N_12302);
or U17685 (N_17685,N_15944,N_14201);
nor U17686 (N_17686,N_14236,N_15242);
xor U17687 (N_17687,N_13834,N_12191);
nor U17688 (N_17688,N_12034,N_14752);
or U17689 (N_17689,N_15067,N_15307);
or U17690 (N_17690,N_15648,N_15412);
or U17691 (N_17691,N_12792,N_14446);
and U17692 (N_17692,N_12023,N_14587);
or U17693 (N_17693,N_13837,N_13873);
nor U17694 (N_17694,N_15707,N_15673);
nand U17695 (N_17695,N_14583,N_15907);
nand U17696 (N_17696,N_12957,N_15518);
and U17697 (N_17697,N_13600,N_13960);
and U17698 (N_17698,N_13084,N_14091);
nor U17699 (N_17699,N_15686,N_13469);
or U17700 (N_17700,N_15204,N_14908);
nor U17701 (N_17701,N_12485,N_12801);
nand U17702 (N_17702,N_14256,N_13329);
and U17703 (N_17703,N_14349,N_14506);
or U17704 (N_17704,N_13158,N_12948);
or U17705 (N_17705,N_15972,N_12066);
nand U17706 (N_17706,N_14343,N_14983);
nand U17707 (N_17707,N_12724,N_13971);
and U17708 (N_17708,N_15504,N_12793);
nand U17709 (N_17709,N_15471,N_12345);
nand U17710 (N_17710,N_12451,N_12116);
and U17711 (N_17711,N_13569,N_14633);
or U17712 (N_17712,N_15803,N_14082);
xnor U17713 (N_17713,N_13623,N_13219);
nand U17714 (N_17714,N_13239,N_13195);
nand U17715 (N_17715,N_12346,N_13749);
nand U17716 (N_17716,N_15196,N_12119);
or U17717 (N_17717,N_13522,N_13575);
nand U17718 (N_17718,N_12859,N_15287);
or U17719 (N_17719,N_12993,N_14420);
xor U17720 (N_17720,N_13736,N_14695);
or U17721 (N_17721,N_12708,N_13908);
and U17722 (N_17722,N_13891,N_14117);
and U17723 (N_17723,N_14998,N_14415);
nor U17724 (N_17724,N_12216,N_13400);
or U17725 (N_17725,N_15401,N_14403);
nor U17726 (N_17726,N_15030,N_13629);
or U17727 (N_17727,N_14652,N_15996);
nor U17728 (N_17728,N_15448,N_14747);
nor U17729 (N_17729,N_13792,N_13385);
or U17730 (N_17730,N_12194,N_13189);
nor U17731 (N_17731,N_14258,N_14500);
and U17732 (N_17732,N_14456,N_15195);
or U17733 (N_17733,N_12060,N_14193);
nand U17734 (N_17734,N_13593,N_13143);
nand U17735 (N_17735,N_13959,N_14198);
or U17736 (N_17736,N_15174,N_15337);
or U17737 (N_17737,N_15742,N_15950);
xnor U17738 (N_17738,N_14453,N_15879);
nand U17739 (N_17739,N_14687,N_12129);
or U17740 (N_17740,N_14546,N_12810);
or U17741 (N_17741,N_14794,N_13932);
nor U17742 (N_17742,N_15010,N_12944);
nor U17743 (N_17743,N_14914,N_13072);
and U17744 (N_17744,N_15865,N_14786);
or U17745 (N_17745,N_14661,N_15557);
nor U17746 (N_17746,N_15509,N_13149);
nor U17747 (N_17747,N_15322,N_12288);
nand U17748 (N_17748,N_13038,N_15080);
or U17749 (N_17749,N_13538,N_15779);
nand U17750 (N_17750,N_14460,N_15281);
nor U17751 (N_17751,N_12420,N_12150);
and U17752 (N_17752,N_12836,N_12234);
or U17753 (N_17753,N_13293,N_14275);
nor U17754 (N_17754,N_14855,N_13976);
or U17755 (N_17755,N_15613,N_12175);
nor U17756 (N_17756,N_13911,N_12100);
and U17757 (N_17757,N_15763,N_12879);
or U17758 (N_17758,N_15345,N_15205);
or U17759 (N_17759,N_15861,N_12450);
and U17760 (N_17760,N_15058,N_14188);
or U17761 (N_17761,N_14513,N_15154);
nor U17762 (N_17762,N_14392,N_13157);
nand U17763 (N_17763,N_13476,N_13955);
and U17764 (N_17764,N_13617,N_12714);
nor U17765 (N_17765,N_14982,N_15862);
nand U17766 (N_17766,N_14214,N_14049);
nor U17767 (N_17767,N_13564,N_13301);
nand U17768 (N_17768,N_13465,N_15137);
or U17769 (N_17769,N_12702,N_13661);
and U17770 (N_17770,N_12935,N_15311);
xor U17771 (N_17771,N_12650,N_14472);
nor U17772 (N_17772,N_12560,N_13993);
nor U17773 (N_17773,N_15905,N_13009);
or U17774 (N_17774,N_13231,N_13893);
nor U17775 (N_17775,N_12606,N_13448);
xor U17776 (N_17776,N_12106,N_14160);
or U17777 (N_17777,N_14985,N_15883);
nor U17778 (N_17778,N_13403,N_13031);
or U17779 (N_17779,N_12223,N_15047);
nand U17780 (N_17780,N_15684,N_12041);
xor U17781 (N_17781,N_15757,N_14194);
nor U17782 (N_17782,N_13771,N_13387);
or U17783 (N_17783,N_13340,N_12693);
nand U17784 (N_17784,N_13427,N_12920);
nor U17785 (N_17785,N_15390,N_13201);
and U17786 (N_17786,N_13369,N_12212);
and U17787 (N_17787,N_14505,N_13025);
or U17788 (N_17788,N_12214,N_15608);
nand U17789 (N_17789,N_13237,N_12998);
nor U17790 (N_17790,N_12578,N_14976);
or U17791 (N_17791,N_12378,N_14040);
nor U17792 (N_17792,N_13924,N_12181);
or U17793 (N_17793,N_15983,N_14015);
nor U17794 (N_17794,N_14418,N_12016);
nor U17795 (N_17795,N_12123,N_15020);
and U17796 (N_17796,N_15283,N_15197);
and U17797 (N_17797,N_14317,N_15904);
nor U17798 (N_17798,N_15481,N_14305);
nor U17799 (N_17799,N_15548,N_14489);
and U17800 (N_17800,N_13233,N_13409);
and U17801 (N_17801,N_12953,N_14021);
nor U17802 (N_17802,N_13294,N_15025);
and U17803 (N_17803,N_13704,N_13883);
nand U17804 (N_17804,N_14090,N_14795);
or U17805 (N_17805,N_14842,N_14710);
nor U17806 (N_17806,N_14263,N_12083);
nand U17807 (N_17807,N_15697,N_13017);
or U17808 (N_17808,N_14308,N_15251);
nor U17809 (N_17809,N_15386,N_14490);
or U17810 (N_17810,N_13968,N_15797);
nor U17811 (N_17811,N_15133,N_13417);
nand U17812 (N_17812,N_12381,N_14108);
and U17813 (N_17813,N_15631,N_12730);
or U17814 (N_17814,N_12046,N_12090);
nand U17815 (N_17815,N_15658,N_13397);
xor U17816 (N_17816,N_13456,N_15255);
and U17817 (N_17817,N_12095,N_13446);
or U17818 (N_17818,N_13366,N_13708);
or U17819 (N_17819,N_14155,N_12122);
nor U17820 (N_17820,N_13152,N_13093);
nand U17821 (N_17821,N_12563,N_12423);
nor U17822 (N_17822,N_15073,N_14896);
xnor U17823 (N_17823,N_12734,N_12323);
and U17824 (N_17824,N_12249,N_13536);
nor U17825 (N_17825,N_15880,N_15859);
and U17826 (N_17826,N_12448,N_14953);
and U17827 (N_17827,N_15940,N_14416);
and U17828 (N_17828,N_12196,N_15112);
and U17829 (N_17829,N_13843,N_14949);
nor U17830 (N_17830,N_15444,N_14191);
and U17831 (N_17831,N_15956,N_13467);
and U17832 (N_17832,N_13350,N_14537);
nor U17833 (N_17833,N_13758,N_14715);
nand U17834 (N_17834,N_15975,N_13050);
and U17835 (N_17835,N_12588,N_14068);
or U17836 (N_17836,N_15979,N_13584);
nand U17837 (N_17837,N_14162,N_14770);
nor U17838 (N_17838,N_15755,N_14635);
nor U17839 (N_17839,N_15591,N_13706);
nand U17840 (N_17840,N_12692,N_13028);
nor U17841 (N_17841,N_13054,N_13872);
nand U17842 (N_17842,N_13735,N_12337);
or U17843 (N_17843,N_14647,N_12891);
and U17844 (N_17844,N_12943,N_13920);
or U17845 (N_17845,N_12333,N_12210);
or U17846 (N_17846,N_12562,N_12566);
and U17847 (N_17847,N_13632,N_14510);
and U17848 (N_17848,N_15065,N_12022);
xor U17849 (N_17849,N_14919,N_13223);
nand U17850 (N_17850,N_12500,N_12950);
and U17851 (N_17851,N_15450,N_14838);
nor U17852 (N_17852,N_12553,N_14017);
and U17853 (N_17853,N_14767,N_13721);
nor U17854 (N_17854,N_15936,N_15747);
and U17855 (N_17855,N_14156,N_14826);
and U17856 (N_17856,N_15246,N_13868);
xor U17857 (N_17857,N_12966,N_12202);
nand U17858 (N_17858,N_12990,N_12422);
and U17859 (N_17859,N_14698,N_12331);
nand U17860 (N_17860,N_12742,N_14649);
and U17861 (N_17861,N_15414,N_14445);
and U17862 (N_17862,N_13372,N_15989);
and U17863 (N_17863,N_14945,N_14078);
nand U17864 (N_17864,N_14248,N_13518);
and U17865 (N_17865,N_14100,N_13338);
nor U17866 (N_17866,N_15750,N_13204);
nand U17867 (N_17867,N_14189,N_14502);
and U17868 (N_17868,N_13827,N_12803);
and U17869 (N_17869,N_14466,N_14677);
nor U17870 (N_17870,N_15280,N_14531);
or U17871 (N_17871,N_15867,N_14202);
nand U17872 (N_17872,N_12525,N_13276);
or U17873 (N_17873,N_13950,N_12790);
nand U17874 (N_17874,N_15832,N_15000);
or U17875 (N_17875,N_15786,N_12496);
or U17876 (N_17876,N_15095,N_12610);
nand U17877 (N_17877,N_15550,N_15924);
and U17878 (N_17878,N_14205,N_15941);
or U17879 (N_17879,N_15143,N_13174);
and U17880 (N_17880,N_13929,N_13969);
or U17881 (N_17881,N_12552,N_13475);
xnor U17882 (N_17882,N_13603,N_12410);
and U17883 (N_17883,N_12089,N_12554);
nand U17884 (N_17884,N_13588,N_12489);
or U17885 (N_17885,N_13378,N_13105);
or U17886 (N_17886,N_12043,N_14038);
or U17887 (N_17887,N_12219,N_13013);
nor U17888 (N_17888,N_13135,N_12136);
and U17889 (N_17889,N_12009,N_14556);
or U17890 (N_17890,N_15774,N_15831);
or U17891 (N_17891,N_13415,N_14447);
and U17892 (N_17892,N_15203,N_15760);
nand U17893 (N_17893,N_15249,N_15024);
nand U17894 (N_17894,N_12341,N_13016);
nor U17895 (N_17895,N_15454,N_15540);
and U17896 (N_17896,N_12091,N_15351);
nand U17897 (N_17897,N_14561,N_15184);
nor U17898 (N_17898,N_15391,N_15269);
or U17899 (N_17899,N_13945,N_15158);
and U17900 (N_17900,N_13621,N_14485);
and U17901 (N_17901,N_12807,N_14669);
xnor U17902 (N_17902,N_14511,N_14250);
nand U17903 (N_17903,N_15237,N_12099);
nor U17904 (N_17904,N_12546,N_12037);
and U17905 (N_17905,N_14168,N_15840);
nor U17906 (N_17906,N_14866,N_14779);
nand U17907 (N_17907,N_14658,N_12640);
nand U17908 (N_17908,N_15226,N_13327);
or U17909 (N_17909,N_15978,N_14733);
nor U17910 (N_17910,N_15315,N_13051);
nor U17911 (N_17911,N_14663,N_14810);
nand U17912 (N_17912,N_13879,N_13654);
and U17913 (N_17913,N_14352,N_12147);
and U17914 (N_17914,N_13852,N_14566);
nand U17915 (N_17915,N_15925,N_15243);
xor U17916 (N_17916,N_12556,N_12584);
and U17917 (N_17917,N_13954,N_13255);
and U17918 (N_17918,N_14993,N_12394);
nand U17919 (N_17919,N_12531,N_14709);
or U17920 (N_17920,N_14825,N_12670);
xor U17921 (N_17921,N_13402,N_15593);
nand U17922 (N_17922,N_15934,N_14704);
nand U17923 (N_17923,N_14270,N_12621);
xor U17924 (N_17924,N_14185,N_13656);
xnor U17925 (N_17925,N_14773,N_12142);
and U17926 (N_17926,N_14348,N_13886);
or U17927 (N_17927,N_12373,N_12524);
or U17928 (N_17928,N_14239,N_14170);
and U17929 (N_17929,N_14997,N_14064);
and U17930 (N_17930,N_12286,N_15427);
nor U17931 (N_17931,N_14014,N_12773);
or U17932 (N_17932,N_13986,N_14938);
xnor U17933 (N_17933,N_12417,N_14536);
nor U17934 (N_17934,N_14876,N_12445);
or U17935 (N_17935,N_14397,N_12857);
nor U17936 (N_17936,N_12481,N_15894);
and U17937 (N_17937,N_15873,N_13136);
nor U17938 (N_17938,N_12255,N_13313);
nand U17939 (N_17939,N_13589,N_13664);
xnor U17940 (N_17940,N_13374,N_14764);
nand U17941 (N_17941,N_15922,N_13160);
and U17942 (N_17942,N_15461,N_14179);
nand U17943 (N_17943,N_14575,N_15895);
nor U17944 (N_17944,N_14781,N_14292);
nor U17945 (N_17945,N_15101,N_12867);
and U17946 (N_17946,N_15129,N_15014);
or U17947 (N_17947,N_13173,N_15912);
nand U17948 (N_17948,N_12528,N_13215);
and U17949 (N_17949,N_13921,N_12727);
nand U17950 (N_17950,N_12964,N_14692);
or U17951 (N_17951,N_13688,N_12213);
nor U17952 (N_17952,N_14457,N_12358);
nor U17953 (N_17953,N_12888,N_12813);
or U17954 (N_17954,N_13699,N_15719);
and U17955 (N_17955,N_13788,N_14748);
nand U17956 (N_17956,N_13352,N_14129);
and U17957 (N_17957,N_12365,N_13889);
or U17958 (N_17958,N_13773,N_14099);
and U17959 (N_17959,N_15099,N_14599);
nand U17960 (N_17960,N_15657,N_14890);
or U17961 (N_17961,N_13933,N_14803);
and U17962 (N_17962,N_12601,N_12231);
xnor U17963 (N_17963,N_15809,N_14469);
or U17964 (N_17964,N_14060,N_13651);
xnor U17965 (N_17965,N_12431,N_12674);
nand U17966 (N_17966,N_15582,N_13678);
nand U17967 (N_17967,N_13942,N_14590);
xnor U17968 (N_17968,N_14111,N_12418);
nor U17969 (N_17969,N_12853,N_15683);
nand U17970 (N_17970,N_15120,N_15353);
nor U17971 (N_17971,N_13119,N_12808);
xnor U17972 (N_17972,N_13328,N_14102);
and U17973 (N_17973,N_15021,N_12511);
and U17974 (N_17974,N_14273,N_12639);
nor U17975 (N_17975,N_12499,N_13668);
nor U17976 (N_17976,N_12717,N_12178);
nand U17977 (N_17977,N_15153,N_12543);
nand U17978 (N_17978,N_14267,N_13401);
xor U17979 (N_17979,N_13984,N_13095);
nand U17980 (N_17980,N_14548,N_12092);
nand U17981 (N_17981,N_15715,N_14907);
and U17982 (N_17982,N_12914,N_13330);
nor U17983 (N_17983,N_12071,N_14374);
and U17984 (N_17984,N_14316,N_12778);
or U17985 (N_17985,N_15990,N_12069);
and U17986 (N_17986,N_15987,N_15964);
and U17987 (N_17987,N_14950,N_15819);
xnor U17988 (N_17988,N_12899,N_12236);
nor U17989 (N_17989,N_12599,N_12700);
nor U17990 (N_17990,N_12084,N_12999);
nand U17991 (N_17991,N_12098,N_14744);
nand U17992 (N_17992,N_13425,N_12342);
or U17993 (N_17993,N_14166,N_13572);
nor U17994 (N_17994,N_13677,N_13829);
xnor U17995 (N_17995,N_14059,N_13634);
or U17996 (N_17996,N_14991,N_15271);
or U17997 (N_17997,N_13556,N_12081);
and U17998 (N_17998,N_12180,N_13863);
nor U17999 (N_17999,N_14379,N_13990);
xor U18000 (N_18000,N_12740,N_12291);
and U18001 (N_18001,N_12009,N_13316);
and U18002 (N_18002,N_12510,N_12610);
or U18003 (N_18003,N_13082,N_13981);
and U18004 (N_18004,N_15459,N_13127);
and U18005 (N_18005,N_12803,N_15686);
nor U18006 (N_18006,N_15587,N_14646);
and U18007 (N_18007,N_15106,N_12267);
or U18008 (N_18008,N_14043,N_15804);
or U18009 (N_18009,N_14768,N_13376);
xnor U18010 (N_18010,N_15236,N_14745);
or U18011 (N_18011,N_13347,N_13976);
and U18012 (N_18012,N_15432,N_15763);
nand U18013 (N_18013,N_12388,N_13278);
and U18014 (N_18014,N_13720,N_12230);
nand U18015 (N_18015,N_12049,N_12692);
or U18016 (N_18016,N_14984,N_14357);
nand U18017 (N_18017,N_15220,N_13273);
nand U18018 (N_18018,N_15578,N_15204);
and U18019 (N_18019,N_14994,N_12641);
nor U18020 (N_18020,N_15540,N_14693);
nand U18021 (N_18021,N_15583,N_14540);
nor U18022 (N_18022,N_13977,N_14436);
and U18023 (N_18023,N_14107,N_12354);
nor U18024 (N_18024,N_14435,N_15115);
xor U18025 (N_18025,N_13610,N_12829);
and U18026 (N_18026,N_14832,N_13769);
and U18027 (N_18027,N_12441,N_14651);
or U18028 (N_18028,N_12773,N_14571);
nand U18029 (N_18029,N_12816,N_12907);
or U18030 (N_18030,N_14772,N_15673);
or U18031 (N_18031,N_12675,N_13491);
nor U18032 (N_18032,N_12547,N_12111);
or U18033 (N_18033,N_12225,N_14841);
nor U18034 (N_18034,N_13847,N_15868);
nand U18035 (N_18035,N_14843,N_15282);
nand U18036 (N_18036,N_14417,N_15379);
nor U18037 (N_18037,N_15552,N_12764);
nand U18038 (N_18038,N_13436,N_13124);
and U18039 (N_18039,N_12244,N_15891);
nand U18040 (N_18040,N_15305,N_15230);
xor U18041 (N_18041,N_14840,N_12854);
or U18042 (N_18042,N_14092,N_12744);
or U18043 (N_18043,N_15986,N_13013);
nand U18044 (N_18044,N_15331,N_12618);
and U18045 (N_18045,N_15908,N_15030);
xnor U18046 (N_18046,N_12355,N_12334);
nor U18047 (N_18047,N_12207,N_13466);
nor U18048 (N_18048,N_15110,N_14388);
or U18049 (N_18049,N_12487,N_14947);
or U18050 (N_18050,N_15594,N_15932);
nor U18051 (N_18051,N_13858,N_13511);
nand U18052 (N_18052,N_14202,N_13502);
or U18053 (N_18053,N_13234,N_14914);
xnor U18054 (N_18054,N_13634,N_12009);
xnor U18055 (N_18055,N_14674,N_12120);
and U18056 (N_18056,N_14252,N_12446);
and U18057 (N_18057,N_12619,N_14656);
and U18058 (N_18058,N_14010,N_14585);
nand U18059 (N_18059,N_15168,N_12707);
and U18060 (N_18060,N_15592,N_15807);
or U18061 (N_18061,N_13836,N_12585);
and U18062 (N_18062,N_14552,N_12615);
nor U18063 (N_18063,N_14254,N_12132);
and U18064 (N_18064,N_14193,N_12812);
xnor U18065 (N_18065,N_15661,N_13331);
or U18066 (N_18066,N_14795,N_13499);
or U18067 (N_18067,N_12259,N_12615);
or U18068 (N_18068,N_13575,N_14565);
nand U18069 (N_18069,N_15001,N_15982);
xor U18070 (N_18070,N_15954,N_13619);
and U18071 (N_18071,N_12719,N_12723);
or U18072 (N_18072,N_13987,N_12951);
or U18073 (N_18073,N_12647,N_13064);
nand U18074 (N_18074,N_13265,N_14709);
nor U18075 (N_18075,N_12955,N_15858);
nor U18076 (N_18076,N_12309,N_13600);
or U18077 (N_18077,N_14288,N_15379);
nand U18078 (N_18078,N_14195,N_14904);
and U18079 (N_18079,N_15836,N_13142);
nand U18080 (N_18080,N_14469,N_15270);
and U18081 (N_18081,N_14874,N_14916);
or U18082 (N_18082,N_14578,N_15345);
nand U18083 (N_18083,N_15244,N_15835);
nand U18084 (N_18084,N_15770,N_12588);
or U18085 (N_18085,N_15638,N_14583);
or U18086 (N_18086,N_15909,N_12375);
nor U18087 (N_18087,N_15411,N_13409);
nand U18088 (N_18088,N_13255,N_13962);
nor U18089 (N_18089,N_14451,N_14767);
nor U18090 (N_18090,N_13656,N_14789);
nand U18091 (N_18091,N_15368,N_15805);
and U18092 (N_18092,N_12440,N_13595);
or U18093 (N_18093,N_12326,N_14438);
or U18094 (N_18094,N_12385,N_15346);
nor U18095 (N_18095,N_12692,N_15215);
nand U18096 (N_18096,N_13664,N_15947);
nor U18097 (N_18097,N_15391,N_12995);
or U18098 (N_18098,N_15106,N_14952);
nor U18099 (N_18099,N_14139,N_14035);
and U18100 (N_18100,N_13690,N_15368);
and U18101 (N_18101,N_13918,N_15799);
nor U18102 (N_18102,N_14031,N_14998);
nand U18103 (N_18103,N_14698,N_12373);
nor U18104 (N_18104,N_15012,N_12091);
and U18105 (N_18105,N_14820,N_14078);
nand U18106 (N_18106,N_15881,N_14237);
nand U18107 (N_18107,N_15157,N_15193);
nor U18108 (N_18108,N_14094,N_12297);
xor U18109 (N_18109,N_12521,N_13771);
nor U18110 (N_18110,N_13056,N_14864);
nor U18111 (N_18111,N_12627,N_12619);
nor U18112 (N_18112,N_14406,N_14133);
and U18113 (N_18113,N_15368,N_12249);
nor U18114 (N_18114,N_12709,N_14953);
and U18115 (N_18115,N_13949,N_13737);
and U18116 (N_18116,N_14811,N_12558);
nor U18117 (N_18117,N_15560,N_15802);
and U18118 (N_18118,N_12599,N_12907);
nor U18119 (N_18119,N_13976,N_15742);
xor U18120 (N_18120,N_12091,N_12782);
and U18121 (N_18121,N_15464,N_14599);
and U18122 (N_18122,N_15363,N_15139);
and U18123 (N_18123,N_14930,N_15785);
and U18124 (N_18124,N_14972,N_13392);
nand U18125 (N_18125,N_15082,N_13678);
nor U18126 (N_18126,N_15696,N_13238);
and U18127 (N_18127,N_13438,N_14142);
nand U18128 (N_18128,N_12343,N_12915);
nor U18129 (N_18129,N_13162,N_12108);
nor U18130 (N_18130,N_12777,N_14726);
and U18131 (N_18131,N_15899,N_13417);
and U18132 (N_18132,N_15775,N_13837);
or U18133 (N_18133,N_12579,N_15282);
nor U18134 (N_18134,N_15607,N_13403);
or U18135 (N_18135,N_13043,N_15372);
and U18136 (N_18136,N_13307,N_14736);
nand U18137 (N_18137,N_12484,N_15295);
nor U18138 (N_18138,N_14197,N_13031);
nor U18139 (N_18139,N_14800,N_15254);
and U18140 (N_18140,N_15322,N_15805);
xnor U18141 (N_18141,N_15874,N_13140);
nor U18142 (N_18142,N_15004,N_15799);
nor U18143 (N_18143,N_12237,N_15890);
and U18144 (N_18144,N_15123,N_13492);
or U18145 (N_18145,N_14413,N_12233);
or U18146 (N_18146,N_14430,N_14193);
nand U18147 (N_18147,N_12517,N_15236);
nor U18148 (N_18148,N_13947,N_13908);
nand U18149 (N_18149,N_13635,N_14215);
nand U18150 (N_18150,N_13429,N_14273);
nand U18151 (N_18151,N_14418,N_14551);
nand U18152 (N_18152,N_14686,N_15685);
nor U18153 (N_18153,N_13043,N_13007);
and U18154 (N_18154,N_13523,N_14444);
nor U18155 (N_18155,N_13402,N_14749);
and U18156 (N_18156,N_14992,N_14538);
and U18157 (N_18157,N_12976,N_15632);
nand U18158 (N_18158,N_15682,N_13939);
nand U18159 (N_18159,N_12159,N_15329);
xor U18160 (N_18160,N_13110,N_13758);
or U18161 (N_18161,N_15203,N_12849);
and U18162 (N_18162,N_13375,N_12343);
xnor U18163 (N_18163,N_15094,N_15659);
xor U18164 (N_18164,N_15918,N_15802);
or U18165 (N_18165,N_13283,N_14951);
nor U18166 (N_18166,N_15184,N_13905);
nor U18167 (N_18167,N_12212,N_14970);
nor U18168 (N_18168,N_12510,N_14180);
and U18169 (N_18169,N_12677,N_12522);
xnor U18170 (N_18170,N_15222,N_13595);
and U18171 (N_18171,N_12885,N_14457);
nand U18172 (N_18172,N_13061,N_12803);
and U18173 (N_18173,N_12437,N_13062);
xor U18174 (N_18174,N_14909,N_13955);
nor U18175 (N_18175,N_13809,N_13623);
or U18176 (N_18176,N_12393,N_12667);
nand U18177 (N_18177,N_15216,N_13599);
and U18178 (N_18178,N_13680,N_14464);
nor U18179 (N_18179,N_15756,N_14755);
nor U18180 (N_18180,N_13953,N_14064);
nand U18181 (N_18181,N_12075,N_15284);
nand U18182 (N_18182,N_14086,N_15936);
or U18183 (N_18183,N_14269,N_12808);
nor U18184 (N_18184,N_13776,N_15644);
and U18185 (N_18185,N_14116,N_14913);
nor U18186 (N_18186,N_12572,N_12604);
nand U18187 (N_18187,N_15574,N_15471);
or U18188 (N_18188,N_15803,N_15703);
xnor U18189 (N_18189,N_15446,N_15940);
nand U18190 (N_18190,N_14936,N_14704);
or U18191 (N_18191,N_14646,N_13275);
nor U18192 (N_18192,N_14305,N_14520);
xor U18193 (N_18193,N_15196,N_12671);
nand U18194 (N_18194,N_12164,N_14944);
nor U18195 (N_18195,N_15175,N_13856);
nor U18196 (N_18196,N_12859,N_14723);
nor U18197 (N_18197,N_15446,N_12822);
nor U18198 (N_18198,N_12885,N_14583);
nand U18199 (N_18199,N_12092,N_14710);
and U18200 (N_18200,N_14320,N_12220);
or U18201 (N_18201,N_14925,N_14633);
nor U18202 (N_18202,N_13313,N_12789);
nor U18203 (N_18203,N_15726,N_15194);
xnor U18204 (N_18204,N_13734,N_13714);
and U18205 (N_18205,N_12525,N_13593);
or U18206 (N_18206,N_12292,N_14532);
or U18207 (N_18207,N_14875,N_15079);
nor U18208 (N_18208,N_13921,N_14294);
and U18209 (N_18209,N_15421,N_12320);
and U18210 (N_18210,N_15569,N_14243);
nor U18211 (N_18211,N_14261,N_15750);
and U18212 (N_18212,N_13993,N_12931);
or U18213 (N_18213,N_13541,N_14499);
or U18214 (N_18214,N_12277,N_13577);
nor U18215 (N_18215,N_15048,N_14067);
or U18216 (N_18216,N_14317,N_14893);
nor U18217 (N_18217,N_14647,N_14315);
xnor U18218 (N_18218,N_13990,N_15403);
or U18219 (N_18219,N_15644,N_15347);
or U18220 (N_18220,N_15603,N_12394);
or U18221 (N_18221,N_14282,N_13863);
or U18222 (N_18222,N_12758,N_15509);
nand U18223 (N_18223,N_12636,N_15934);
and U18224 (N_18224,N_12542,N_14817);
nor U18225 (N_18225,N_14542,N_12851);
and U18226 (N_18226,N_15436,N_13033);
nor U18227 (N_18227,N_13850,N_15179);
nand U18228 (N_18228,N_14703,N_12247);
nor U18229 (N_18229,N_14833,N_15148);
nor U18230 (N_18230,N_15679,N_15459);
nand U18231 (N_18231,N_12629,N_13523);
or U18232 (N_18232,N_15460,N_14291);
nand U18233 (N_18233,N_15355,N_14619);
and U18234 (N_18234,N_13382,N_14008);
nor U18235 (N_18235,N_12095,N_13757);
nor U18236 (N_18236,N_13388,N_13477);
and U18237 (N_18237,N_13307,N_14412);
nand U18238 (N_18238,N_15912,N_12105);
and U18239 (N_18239,N_13435,N_14540);
nand U18240 (N_18240,N_15557,N_12718);
nand U18241 (N_18241,N_15232,N_13955);
and U18242 (N_18242,N_15919,N_12834);
xor U18243 (N_18243,N_15093,N_13101);
xor U18244 (N_18244,N_12077,N_13914);
nand U18245 (N_18245,N_12491,N_12940);
nor U18246 (N_18246,N_12872,N_15199);
nand U18247 (N_18247,N_14415,N_12497);
nor U18248 (N_18248,N_14205,N_12555);
xnor U18249 (N_18249,N_14990,N_15472);
nand U18250 (N_18250,N_15432,N_15515);
xnor U18251 (N_18251,N_15183,N_12028);
and U18252 (N_18252,N_14945,N_14586);
nor U18253 (N_18253,N_15970,N_14316);
nor U18254 (N_18254,N_15410,N_13219);
nor U18255 (N_18255,N_13191,N_12129);
and U18256 (N_18256,N_12893,N_12624);
nand U18257 (N_18257,N_15069,N_15406);
nor U18258 (N_18258,N_15645,N_12715);
and U18259 (N_18259,N_12664,N_14618);
nor U18260 (N_18260,N_14968,N_15021);
nor U18261 (N_18261,N_15825,N_13088);
or U18262 (N_18262,N_12942,N_13334);
or U18263 (N_18263,N_13429,N_15449);
nor U18264 (N_18264,N_14035,N_12109);
and U18265 (N_18265,N_15504,N_14964);
or U18266 (N_18266,N_15646,N_12217);
or U18267 (N_18267,N_13047,N_15498);
nand U18268 (N_18268,N_12262,N_15522);
nand U18269 (N_18269,N_14974,N_15072);
nor U18270 (N_18270,N_12263,N_13277);
or U18271 (N_18271,N_13903,N_12616);
or U18272 (N_18272,N_13808,N_13522);
nor U18273 (N_18273,N_12996,N_15531);
and U18274 (N_18274,N_12686,N_13388);
xnor U18275 (N_18275,N_13810,N_14533);
or U18276 (N_18276,N_14339,N_13864);
nand U18277 (N_18277,N_15639,N_12742);
and U18278 (N_18278,N_13520,N_14043);
and U18279 (N_18279,N_15071,N_14817);
or U18280 (N_18280,N_15962,N_12185);
nor U18281 (N_18281,N_13069,N_15672);
nor U18282 (N_18282,N_15078,N_12561);
nand U18283 (N_18283,N_14423,N_13562);
and U18284 (N_18284,N_15485,N_12100);
and U18285 (N_18285,N_15937,N_15990);
and U18286 (N_18286,N_15382,N_12621);
xor U18287 (N_18287,N_15694,N_13903);
nor U18288 (N_18288,N_12701,N_14090);
and U18289 (N_18289,N_13760,N_15158);
and U18290 (N_18290,N_15842,N_12727);
nand U18291 (N_18291,N_15805,N_13540);
nor U18292 (N_18292,N_15900,N_15930);
or U18293 (N_18293,N_14252,N_15587);
or U18294 (N_18294,N_14622,N_14992);
or U18295 (N_18295,N_14406,N_15347);
and U18296 (N_18296,N_12743,N_15098);
xnor U18297 (N_18297,N_12840,N_14515);
and U18298 (N_18298,N_13882,N_12419);
nor U18299 (N_18299,N_12389,N_14857);
nor U18300 (N_18300,N_13643,N_15117);
or U18301 (N_18301,N_12345,N_15849);
and U18302 (N_18302,N_15639,N_12843);
nor U18303 (N_18303,N_14572,N_14675);
nand U18304 (N_18304,N_12534,N_15316);
nor U18305 (N_18305,N_13716,N_12006);
nand U18306 (N_18306,N_15551,N_13634);
nand U18307 (N_18307,N_15658,N_13164);
nor U18308 (N_18308,N_13998,N_14189);
and U18309 (N_18309,N_15466,N_13821);
nand U18310 (N_18310,N_15267,N_13215);
nand U18311 (N_18311,N_12058,N_14737);
and U18312 (N_18312,N_13039,N_12183);
or U18313 (N_18313,N_15223,N_15550);
nor U18314 (N_18314,N_15708,N_13940);
nand U18315 (N_18315,N_13108,N_12356);
nor U18316 (N_18316,N_15564,N_13083);
nand U18317 (N_18317,N_13801,N_13184);
and U18318 (N_18318,N_14889,N_13614);
or U18319 (N_18319,N_15424,N_12684);
or U18320 (N_18320,N_13335,N_15659);
nand U18321 (N_18321,N_13495,N_13211);
nand U18322 (N_18322,N_12849,N_14904);
and U18323 (N_18323,N_14640,N_12687);
nor U18324 (N_18324,N_12200,N_13924);
nand U18325 (N_18325,N_12307,N_12001);
or U18326 (N_18326,N_14001,N_12066);
or U18327 (N_18327,N_15220,N_12811);
and U18328 (N_18328,N_14852,N_15050);
and U18329 (N_18329,N_13371,N_15066);
and U18330 (N_18330,N_15979,N_14522);
nand U18331 (N_18331,N_14687,N_14831);
nor U18332 (N_18332,N_14710,N_12489);
nand U18333 (N_18333,N_15994,N_15703);
and U18334 (N_18334,N_12105,N_12129);
xnor U18335 (N_18335,N_15339,N_15124);
nand U18336 (N_18336,N_14591,N_13039);
and U18337 (N_18337,N_12201,N_15895);
and U18338 (N_18338,N_15446,N_15663);
and U18339 (N_18339,N_14263,N_12972);
nand U18340 (N_18340,N_15889,N_15472);
and U18341 (N_18341,N_12492,N_14200);
xor U18342 (N_18342,N_15482,N_14926);
nor U18343 (N_18343,N_15872,N_15323);
nand U18344 (N_18344,N_12798,N_14404);
nor U18345 (N_18345,N_15681,N_12246);
or U18346 (N_18346,N_15903,N_14085);
nand U18347 (N_18347,N_15415,N_15628);
nand U18348 (N_18348,N_15793,N_15271);
nand U18349 (N_18349,N_13796,N_14596);
or U18350 (N_18350,N_15558,N_13265);
or U18351 (N_18351,N_15776,N_15578);
and U18352 (N_18352,N_12905,N_13979);
nand U18353 (N_18353,N_12491,N_14573);
nand U18354 (N_18354,N_15715,N_12037);
and U18355 (N_18355,N_15971,N_12175);
nand U18356 (N_18356,N_12425,N_12440);
nand U18357 (N_18357,N_12684,N_14076);
nand U18358 (N_18358,N_12526,N_12806);
and U18359 (N_18359,N_12310,N_14566);
and U18360 (N_18360,N_14496,N_15206);
nand U18361 (N_18361,N_12977,N_12531);
or U18362 (N_18362,N_13290,N_15799);
and U18363 (N_18363,N_14855,N_13599);
nand U18364 (N_18364,N_15157,N_12252);
nand U18365 (N_18365,N_13899,N_12685);
and U18366 (N_18366,N_13994,N_14957);
nor U18367 (N_18367,N_14251,N_15985);
nor U18368 (N_18368,N_12667,N_13988);
nand U18369 (N_18369,N_14812,N_13503);
xnor U18370 (N_18370,N_14291,N_13690);
or U18371 (N_18371,N_15319,N_12487);
nor U18372 (N_18372,N_14536,N_13365);
and U18373 (N_18373,N_13704,N_15615);
nor U18374 (N_18374,N_12475,N_14886);
and U18375 (N_18375,N_12178,N_15900);
nand U18376 (N_18376,N_15889,N_13563);
nand U18377 (N_18377,N_13642,N_14538);
nor U18378 (N_18378,N_15666,N_14389);
and U18379 (N_18379,N_13230,N_12734);
or U18380 (N_18380,N_12512,N_13753);
or U18381 (N_18381,N_12092,N_15641);
or U18382 (N_18382,N_13745,N_12614);
or U18383 (N_18383,N_13180,N_14700);
or U18384 (N_18384,N_13640,N_15380);
and U18385 (N_18385,N_14167,N_13163);
nand U18386 (N_18386,N_15032,N_13817);
xnor U18387 (N_18387,N_15644,N_12749);
nor U18388 (N_18388,N_13502,N_13678);
and U18389 (N_18389,N_15055,N_15082);
or U18390 (N_18390,N_14688,N_15234);
nor U18391 (N_18391,N_14633,N_14371);
xnor U18392 (N_18392,N_12858,N_15937);
and U18393 (N_18393,N_12766,N_14665);
xnor U18394 (N_18394,N_15082,N_14690);
nand U18395 (N_18395,N_15074,N_13930);
or U18396 (N_18396,N_13565,N_14300);
and U18397 (N_18397,N_13865,N_14596);
xnor U18398 (N_18398,N_14525,N_15535);
nand U18399 (N_18399,N_15400,N_13316);
nand U18400 (N_18400,N_13007,N_14240);
nand U18401 (N_18401,N_15151,N_15843);
nor U18402 (N_18402,N_12622,N_12734);
xor U18403 (N_18403,N_13352,N_14050);
xnor U18404 (N_18404,N_12474,N_15618);
nor U18405 (N_18405,N_12838,N_12797);
nand U18406 (N_18406,N_14094,N_15953);
nand U18407 (N_18407,N_13783,N_14943);
nand U18408 (N_18408,N_12230,N_12920);
or U18409 (N_18409,N_13500,N_14357);
and U18410 (N_18410,N_14421,N_13496);
and U18411 (N_18411,N_15807,N_15830);
and U18412 (N_18412,N_14486,N_13662);
xor U18413 (N_18413,N_14314,N_13011);
xor U18414 (N_18414,N_15427,N_13492);
or U18415 (N_18415,N_12662,N_12174);
or U18416 (N_18416,N_14584,N_12526);
nand U18417 (N_18417,N_13181,N_13559);
nand U18418 (N_18418,N_13988,N_12211);
and U18419 (N_18419,N_13470,N_14988);
and U18420 (N_18420,N_13684,N_14348);
nor U18421 (N_18421,N_12155,N_14491);
or U18422 (N_18422,N_15863,N_14293);
nor U18423 (N_18423,N_14357,N_15167);
or U18424 (N_18424,N_14801,N_15791);
nor U18425 (N_18425,N_13040,N_15211);
or U18426 (N_18426,N_12702,N_15068);
xnor U18427 (N_18427,N_12103,N_15305);
or U18428 (N_18428,N_12004,N_15273);
or U18429 (N_18429,N_14701,N_13932);
nor U18430 (N_18430,N_12928,N_14352);
or U18431 (N_18431,N_13154,N_13414);
nor U18432 (N_18432,N_12063,N_13102);
and U18433 (N_18433,N_15981,N_14732);
or U18434 (N_18434,N_15086,N_14963);
or U18435 (N_18435,N_12174,N_13555);
and U18436 (N_18436,N_13167,N_12146);
xnor U18437 (N_18437,N_15236,N_12803);
nor U18438 (N_18438,N_15392,N_13256);
nand U18439 (N_18439,N_15607,N_13122);
nand U18440 (N_18440,N_12380,N_15683);
nor U18441 (N_18441,N_15497,N_13596);
and U18442 (N_18442,N_12003,N_15457);
nand U18443 (N_18443,N_15946,N_12603);
xnor U18444 (N_18444,N_14886,N_12321);
and U18445 (N_18445,N_12262,N_12054);
or U18446 (N_18446,N_14104,N_12182);
and U18447 (N_18447,N_15462,N_14200);
or U18448 (N_18448,N_14953,N_14784);
xnor U18449 (N_18449,N_13937,N_13985);
xnor U18450 (N_18450,N_14958,N_13633);
xor U18451 (N_18451,N_15332,N_14085);
and U18452 (N_18452,N_15143,N_14269);
and U18453 (N_18453,N_14859,N_14928);
or U18454 (N_18454,N_12470,N_15419);
and U18455 (N_18455,N_13880,N_14221);
nor U18456 (N_18456,N_14426,N_13803);
nor U18457 (N_18457,N_14504,N_13957);
nand U18458 (N_18458,N_12103,N_12966);
or U18459 (N_18459,N_15182,N_13320);
nand U18460 (N_18460,N_12582,N_14750);
nand U18461 (N_18461,N_13232,N_13514);
nand U18462 (N_18462,N_13056,N_12313);
nand U18463 (N_18463,N_14564,N_13213);
nand U18464 (N_18464,N_13569,N_14480);
and U18465 (N_18465,N_12421,N_15417);
and U18466 (N_18466,N_15796,N_14666);
nand U18467 (N_18467,N_15453,N_13813);
nor U18468 (N_18468,N_14779,N_12433);
or U18469 (N_18469,N_13768,N_12244);
xnor U18470 (N_18470,N_13133,N_15319);
and U18471 (N_18471,N_14842,N_14033);
or U18472 (N_18472,N_13859,N_13064);
nor U18473 (N_18473,N_13556,N_15511);
or U18474 (N_18474,N_14561,N_12295);
or U18475 (N_18475,N_15996,N_15381);
or U18476 (N_18476,N_12351,N_12940);
xor U18477 (N_18477,N_12308,N_14845);
nor U18478 (N_18478,N_13083,N_15639);
and U18479 (N_18479,N_12918,N_13099);
nor U18480 (N_18480,N_12086,N_12926);
nand U18481 (N_18481,N_14144,N_13612);
nand U18482 (N_18482,N_12733,N_13190);
or U18483 (N_18483,N_14058,N_15639);
and U18484 (N_18484,N_15245,N_15798);
nand U18485 (N_18485,N_12242,N_13826);
nand U18486 (N_18486,N_15316,N_12959);
nor U18487 (N_18487,N_15916,N_12062);
xor U18488 (N_18488,N_14837,N_12196);
nand U18489 (N_18489,N_13608,N_12385);
or U18490 (N_18490,N_15493,N_12465);
or U18491 (N_18491,N_12907,N_15085);
or U18492 (N_18492,N_13005,N_14490);
nor U18493 (N_18493,N_12925,N_15080);
xnor U18494 (N_18494,N_15991,N_14637);
or U18495 (N_18495,N_13240,N_14396);
nor U18496 (N_18496,N_14306,N_14760);
and U18497 (N_18497,N_14800,N_14870);
or U18498 (N_18498,N_13260,N_15329);
and U18499 (N_18499,N_14475,N_12292);
and U18500 (N_18500,N_13436,N_13018);
xnor U18501 (N_18501,N_12065,N_13197);
nand U18502 (N_18502,N_15221,N_12627);
nor U18503 (N_18503,N_12872,N_15599);
or U18504 (N_18504,N_13082,N_12025);
or U18505 (N_18505,N_14775,N_14488);
and U18506 (N_18506,N_13765,N_15018);
and U18507 (N_18507,N_15971,N_15282);
xnor U18508 (N_18508,N_13449,N_12670);
nand U18509 (N_18509,N_14301,N_15382);
xnor U18510 (N_18510,N_15112,N_15559);
and U18511 (N_18511,N_15197,N_12687);
nor U18512 (N_18512,N_14062,N_15233);
or U18513 (N_18513,N_13534,N_15232);
and U18514 (N_18514,N_15538,N_15933);
nand U18515 (N_18515,N_12628,N_12458);
or U18516 (N_18516,N_14155,N_15787);
and U18517 (N_18517,N_15196,N_12182);
and U18518 (N_18518,N_13641,N_13043);
or U18519 (N_18519,N_13977,N_15300);
and U18520 (N_18520,N_14379,N_13370);
nand U18521 (N_18521,N_15720,N_12884);
nor U18522 (N_18522,N_14857,N_14748);
nand U18523 (N_18523,N_15185,N_14149);
nand U18524 (N_18524,N_14802,N_15260);
nand U18525 (N_18525,N_13557,N_13633);
nor U18526 (N_18526,N_14366,N_15332);
or U18527 (N_18527,N_15271,N_13914);
nand U18528 (N_18528,N_14320,N_14779);
nor U18529 (N_18529,N_15648,N_14632);
and U18530 (N_18530,N_13519,N_14683);
or U18531 (N_18531,N_13235,N_15474);
or U18532 (N_18532,N_12708,N_14864);
or U18533 (N_18533,N_15487,N_15654);
xnor U18534 (N_18534,N_15438,N_14658);
or U18535 (N_18535,N_15627,N_12070);
nand U18536 (N_18536,N_12910,N_15144);
or U18537 (N_18537,N_13856,N_13016);
or U18538 (N_18538,N_13044,N_12855);
nor U18539 (N_18539,N_13314,N_13438);
or U18540 (N_18540,N_13787,N_12738);
or U18541 (N_18541,N_12908,N_12592);
and U18542 (N_18542,N_14020,N_13085);
or U18543 (N_18543,N_12134,N_14679);
xor U18544 (N_18544,N_13398,N_12069);
and U18545 (N_18545,N_14271,N_13834);
xor U18546 (N_18546,N_14362,N_15908);
or U18547 (N_18547,N_12070,N_14517);
or U18548 (N_18548,N_13780,N_15596);
or U18549 (N_18549,N_15069,N_15968);
nand U18550 (N_18550,N_12971,N_13758);
nand U18551 (N_18551,N_12463,N_14102);
nor U18552 (N_18552,N_15859,N_14523);
and U18553 (N_18553,N_12082,N_15983);
nand U18554 (N_18554,N_14245,N_14566);
xor U18555 (N_18555,N_13596,N_14729);
and U18556 (N_18556,N_15505,N_15721);
or U18557 (N_18557,N_12278,N_13324);
or U18558 (N_18558,N_15318,N_15337);
nand U18559 (N_18559,N_13236,N_13406);
or U18560 (N_18560,N_13872,N_15807);
or U18561 (N_18561,N_13494,N_14439);
nor U18562 (N_18562,N_13331,N_13907);
and U18563 (N_18563,N_12461,N_12707);
nor U18564 (N_18564,N_12982,N_12458);
and U18565 (N_18565,N_13627,N_12051);
and U18566 (N_18566,N_14372,N_15139);
or U18567 (N_18567,N_13429,N_15921);
and U18568 (N_18568,N_12433,N_15081);
or U18569 (N_18569,N_15329,N_15123);
and U18570 (N_18570,N_15659,N_13807);
and U18571 (N_18571,N_14904,N_15113);
nand U18572 (N_18572,N_14937,N_13521);
nor U18573 (N_18573,N_14707,N_14390);
and U18574 (N_18574,N_14770,N_12584);
nand U18575 (N_18575,N_13745,N_12470);
or U18576 (N_18576,N_15658,N_14285);
or U18577 (N_18577,N_15299,N_13002);
and U18578 (N_18578,N_12303,N_12101);
nand U18579 (N_18579,N_14405,N_14875);
and U18580 (N_18580,N_15067,N_13057);
nor U18581 (N_18581,N_14318,N_14994);
nand U18582 (N_18582,N_15558,N_14958);
nor U18583 (N_18583,N_14862,N_13389);
and U18584 (N_18584,N_15714,N_13431);
or U18585 (N_18585,N_12136,N_12701);
and U18586 (N_18586,N_13234,N_15649);
nor U18587 (N_18587,N_14389,N_15387);
xnor U18588 (N_18588,N_14331,N_15156);
or U18589 (N_18589,N_12520,N_12955);
nor U18590 (N_18590,N_12340,N_15091);
and U18591 (N_18591,N_13928,N_15317);
nor U18592 (N_18592,N_14890,N_12642);
xor U18593 (N_18593,N_15068,N_15256);
nand U18594 (N_18594,N_13541,N_14687);
nor U18595 (N_18595,N_12608,N_15248);
nand U18596 (N_18596,N_12133,N_13209);
xor U18597 (N_18597,N_14459,N_12614);
nand U18598 (N_18598,N_13724,N_14555);
and U18599 (N_18599,N_13098,N_14794);
nor U18600 (N_18600,N_12546,N_12270);
xor U18601 (N_18601,N_13375,N_13049);
nand U18602 (N_18602,N_15117,N_13291);
xor U18603 (N_18603,N_14206,N_13664);
and U18604 (N_18604,N_15162,N_14644);
nand U18605 (N_18605,N_13053,N_12708);
nor U18606 (N_18606,N_14880,N_12495);
and U18607 (N_18607,N_12144,N_15457);
and U18608 (N_18608,N_15412,N_13706);
or U18609 (N_18609,N_13093,N_15940);
nor U18610 (N_18610,N_13063,N_13569);
and U18611 (N_18611,N_14064,N_12355);
nand U18612 (N_18612,N_14987,N_13438);
nand U18613 (N_18613,N_14047,N_14099);
and U18614 (N_18614,N_13877,N_15844);
xnor U18615 (N_18615,N_12956,N_15706);
or U18616 (N_18616,N_13087,N_14279);
nor U18617 (N_18617,N_14124,N_14355);
or U18618 (N_18618,N_13929,N_14250);
or U18619 (N_18619,N_14817,N_14274);
and U18620 (N_18620,N_13238,N_12416);
nand U18621 (N_18621,N_14620,N_12538);
or U18622 (N_18622,N_13329,N_13378);
or U18623 (N_18623,N_13127,N_14261);
xor U18624 (N_18624,N_12607,N_15076);
xor U18625 (N_18625,N_14878,N_14632);
nand U18626 (N_18626,N_14525,N_12351);
or U18627 (N_18627,N_14470,N_13964);
and U18628 (N_18628,N_13080,N_12186);
nand U18629 (N_18629,N_12478,N_14717);
and U18630 (N_18630,N_15813,N_15573);
and U18631 (N_18631,N_12235,N_12015);
nand U18632 (N_18632,N_14835,N_15264);
nand U18633 (N_18633,N_14810,N_15130);
nor U18634 (N_18634,N_13648,N_12940);
or U18635 (N_18635,N_13324,N_12686);
or U18636 (N_18636,N_14013,N_12779);
nor U18637 (N_18637,N_13564,N_14813);
or U18638 (N_18638,N_12251,N_13818);
nor U18639 (N_18639,N_12269,N_13255);
nor U18640 (N_18640,N_14316,N_14636);
and U18641 (N_18641,N_12366,N_14149);
nor U18642 (N_18642,N_14473,N_14062);
nand U18643 (N_18643,N_14010,N_12802);
and U18644 (N_18644,N_14470,N_12370);
or U18645 (N_18645,N_15186,N_13691);
and U18646 (N_18646,N_15141,N_14695);
and U18647 (N_18647,N_15541,N_15877);
or U18648 (N_18648,N_13719,N_13606);
and U18649 (N_18649,N_13135,N_15255);
nor U18650 (N_18650,N_15363,N_13481);
or U18651 (N_18651,N_12245,N_14807);
or U18652 (N_18652,N_12694,N_13786);
nor U18653 (N_18653,N_15178,N_14202);
nor U18654 (N_18654,N_14606,N_15470);
nand U18655 (N_18655,N_13234,N_15115);
and U18656 (N_18656,N_12070,N_14271);
or U18657 (N_18657,N_12138,N_14768);
or U18658 (N_18658,N_15696,N_12172);
or U18659 (N_18659,N_14716,N_13044);
or U18660 (N_18660,N_13324,N_14137);
nor U18661 (N_18661,N_15208,N_14848);
nand U18662 (N_18662,N_13115,N_12109);
nand U18663 (N_18663,N_14333,N_13901);
xnor U18664 (N_18664,N_12599,N_13803);
nor U18665 (N_18665,N_15857,N_14972);
nor U18666 (N_18666,N_12249,N_14795);
or U18667 (N_18667,N_15296,N_14950);
nand U18668 (N_18668,N_14031,N_14822);
or U18669 (N_18669,N_14517,N_12839);
xor U18670 (N_18670,N_13185,N_12574);
or U18671 (N_18671,N_14478,N_12206);
or U18672 (N_18672,N_15404,N_13373);
or U18673 (N_18673,N_13997,N_14751);
or U18674 (N_18674,N_12896,N_14902);
nand U18675 (N_18675,N_15890,N_14668);
and U18676 (N_18676,N_13009,N_14590);
and U18677 (N_18677,N_13939,N_12663);
nor U18678 (N_18678,N_12979,N_12685);
nor U18679 (N_18679,N_15534,N_12047);
or U18680 (N_18680,N_14718,N_12778);
and U18681 (N_18681,N_12573,N_15521);
nor U18682 (N_18682,N_14259,N_15601);
nand U18683 (N_18683,N_13208,N_12583);
and U18684 (N_18684,N_13006,N_14859);
nor U18685 (N_18685,N_15992,N_14037);
xnor U18686 (N_18686,N_12456,N_12561);
nor U18687 (N_18687,N_15153,N_12839);
nor U18688 (N_18688,N_12569,N_13722);
nor U18689 (N_18689,N_12058,N_15508);
xor U18690 (N_18690,N_15024,N_12094);
and U18691 (N_18691,N_12333,N_12091);
or U18692 (N_18692,N_13501,N_14793);
or U18693 (N_18693,N_13559,N_15858);
or U18694 (N_18694,N_15969,N_12477);
nand U18695 (N_18695,N_14139,N_12595);
or U18696 (N_18696,N_15892,N_14353);
nor U18697 (N_18697,N_12041,N_14492);
or U18698 (N_18698,N_13383,N_12776);
nor U18699 (N_18699,N_15807,N_12326);
or U18700 (N_18700,N_14642,N_15743);
nand U18701 (N_18701,N_12479,N_13844);
xor U18702 (N_18702,N_14922,N_14585);
nor U18703 (N_18703,N_12978,N_12484);
xnor U18704 (N_18704,N_12382,N_12681);
nor U18705 (N_18705,N_12512,N_12678);
nand U18706 (N_18706,N_14027,N_12520);
or U18707 (N_18707,N_12746,N_14604);
nor U18708 (N_18708,N_15450,N_14614);
nor U18709 (N_18709,N_15401,N_14558);
nand U18710 (N_18710,N_12006,N_14524);
nand U18711 (N_18711,N_12776,N_13273);
and U18712 (N_18712,N_14256,N_14624);
xor U18713 (N_18713,N_14026,N_12156);
or U18714 (N_18714,N_12125,N_13526);
and U18715 (N_18715,N_13360,N_14924);
xnor U18716 (N_18716,N_13061,N_15531);
nor U18717 (N_18717,N_15392,N_14369);
xnor U18718 (N_18718,N_15887,N_13833);
and U18719 (N_18719,N_13394,N_14638);
and U18720 (N_18720,N_13877,N_14221);
or U18721 (N_18721,N_12629,N_13610);
and U18722 (N_18722,N_13204,N_12504);
or U18723 (N_18723,N_12407,N_14921);
and U18724 (N_18724,N_12299,N_13456);
nand U18725 (N_18725,N_13891,N_15890);
or U18726 (N_18726,N_15715,N_12899);
or U18727 (N_18727,N_13870,N_14512);
or U18728 (N_18728,N_13908,N_14088);
or U18729 (N_18729,N_14955,N_13452);
or U18730 (N_18730,N_14473,N_13674);
nor U18731 (N_18731,N_14978,N_12769);
nor U18732 (N_18732,N_13867,N_12484);
and U18733 (N_18733,N_15802,N_12041);
and U18734 (N_18734,N_12755,N_13246);
or U18735 (N_18735,N_14116,N_14277);
nand U18736 (N_18736,N_13432,N_14652);
or U18737 (N_18737,N_13925,N_12362);
or U18738 (N_18738,N_12399,N_12630);
nor U18739 (N_18739,N_15899,N_15413);
nor U18740 (N_18740,N_13879,N_15772);
nor U18741 (N_18741,N_14209,N_13124);
or U18742 (N_18742,N_12855,N_13649);
and U18743 (N_18743,N_14282,N_12110);
and U18744 (N_18744,N_13284,N_14549);
and U18745 (N_18745,N_14430,N_14024);
nor U18746 (N_18746,N_14886,N_13563);
and U18747 (N_18747,N_15861,N_13758);
or U18748 (N_18748,N_13983,N_12532);
and U18749 (N_18749,N_14320,N_15029);
and U18750 (N_18750,N_13787,N_13438);
or U18751 (N_18751,N_14286,N_12362);
nor U18752 (N_18752,N_14850,N_14522);
nor U18753 (N_18753,N_15246,N_14814);
nand U18754 (N_18754,N_14636,N_13247);
nand U18755 (N_18755,N_14599,N_12836);
and U18756 (N_18756,N_14308,N_14641);
nand U18757 (N_18757,N_13319,N_12022);
nand U18758 (N_18758,N_12100,N_15621);
nand U18759 (N_18759,N_13535,N_13634);
or U18760 (N_18760,N_12290,N_13492);
and U18761 (N_18761,N_15572,N_15429);
and U18762 (N_18762,N_15970,N_14356);
and U18763 (N_18763,N_14965,N_15058);
nor U18764 (N_18764,N_12462,N_15428);
nand U18765 (N_18765,N_12793,N_13646);
and U18766 (N_18766,N_12697,N_15177);
nor U18767 (N_18767,N_13261,N_13334);
and U18768 (N_18768,N_12849,N_12765);
or U18769 (N_18769,N_13737,N_12528);
or U18770 (N_18770,N_13199,N_15390);
nor U18771 (N_18771,N_13269,N_15158);
nand U18772 (N_18772,N_14039,N_14886);
nand U18773 (N_18773,N_15723,N_12303);
nor U18774 (N_18774,N_12765,N_13437);
and U18775 (N_18775,N_12144,N_13337);
nand U18776 (N_18776,N_12319,N_12311);
or U18777 (N_18777,N_15913,N_15004);
nand U18778 (N_18778,N_15411,N_12039);
nor U18779 (N_18779,N_12071,N_12304);
and U18780 (N_18780,N_15188,N_13602);
nor U18781 (N_18781,N_14440,N_14923);
nor U18782 (N_18782,N_15669,N_13173);
and U18783 (N_18783,N_13914,N_14413);
nand U18784 (N_18784,N_12342,N_13466);
nor U18785 (N_18785,N_14545,N_12706);
nor U18786 (N_18786,N_15791,N_12796);
xnor U18787 (N_18787,N_15877,N_15757);
and U18788 (N_18788,N_12408,N_14686);
nand U18789 (N_18789,N_14614,N_13670);
xor U18790 (N_18790,N_13995,N_12125);
nor U18791 (N_18791,N_12489,N_14978);
and U18792 (N_18792,N_14808,N_12550);
or U18793 (N_18793,N_12908,N_14961);
nor U18794 (N_18794,N_14646,N_12976);
and U18795 (N_18795,N_12218,N_14828);
xor U18796 (N_18796,N_13033,N_15190);
xor U18797 (N_18797,N_12604,N_15954);
or U18798 (N_18798,N_12235,N_14795);
and U18799 (N_18799,N_13774,N_13012);
or U18800 (N_18800,N_15253,N_14732);
xor U18801 (N_18801,N_15784,N_12383);
nor U18802 (N_18802,N_15430,N_13887);
or U18803 (N_18803,N_13421,N_14355);
or U18804 (N_18804,N_15787,N_15766);
nand U18805 (N_18805,N_12693,N_12037);
nand U18806 (N_18806,N_14951,N_15421);
nand U18807 (N_18807,N_14112,N_15986);
nor U18808 (N_18808,N_15984,N_15110);
nor U18809 (N_18809,N_14593,N_13094);
and U18810 (N_18810,N_14026,N_14783);
and U18811 (N_18811,N_12206,N_12056);
and U18812 (N_18812,N_14942,N_14826);
and U18813 (N_18813,N_15789,N_12229);
and U18814 (N_18814,N_13558,N_14917);
nand U18815 (N_18815,N_14691,N_14562);
or U18816 (N_18816,N_14420,N_15916);
nand U18817 (N_18817,N_12444,N_12649);
and U18818 (N_18818,N_15510,N_13371);
nor U18819 (N_18819,N_13868,N_14264);
xnor U18820 (N_18820,N_13489,N_12021);
nor U18821 (N_18821,N_12222,N_14555);
and U18822 (N_18822,N_13982,N_13327);
nand U18823 (N_18823,N_13297,N_12092);
xor U18824 (N_18824,N_15633,N_13685);
or U18825 (N_18825,N_14016,N_12955);
and U18826 (N_18826,N_15263,N_13231);
nor U18827 (N_18827,N_13223,N_15763);
and U18828 (N_18828,N_15554,N_12218);
nor U18829 (N_18829,N_14821,N_14409);
nand U18830 (N_18830,N_15929,N_13530);
nor U18831 (N_18831,N_14716,N_12974);
or U18832 (N_18832,N_14443,N_12764);
and U18833 (N_18833,N_12017,N_13466);
or U18834 (N_18834,N_13639,N_13979);
nor U18835 (N_18835,N_14872,N_15751);
or U18836 (N_18836,N_15210,N_12238);
nor U18837 (N_18837,N_14246,N_15926);
nand U18838 (N_18838,N_13359,N_15102);
and U18839 (N_18839,N_14264,N_12748);
and U18840 (N_18840,N_15237,N_15161);
or U18841 (N_18841,N_15133,N_12732);
or U18842 (N_18842,N_13544,N_13827);
nor U18843 (N_18843,N_13136,N_13455);
and U18844 (N_18844,N_15436,N_15470);
nand U18845 (N_18845,N_14361,N_14619);
and U18846 (N_18846,N_15678,N_12110);
nand U18847 (N_18847,N_14009,N_15646);
and U18848 (N_18848,N_15771,N_14401);
nand U18849 (N_18849,N_14907,N_15209);
and U18850 (N_18850,N_15837,N_13964);
nand U18851 (N_18851,N_15885,N_14319);
xnor U18852 (N_18852,N_12815,N_13540);
nor U18853 (N_18853,N_13425,N_12379);
and U18854 (N_18854,N_12164,N_14457);
xnor U18855 (N_18855,N_12989,N_15736);
nand U18856 (N_18856,N_15091,N_14607);
and U18857 (N_18857,N_12820,N_12773);
nor U18858 (N_18858,N_15223,N_12430);
or U18859 (N_18859,N_14198,N_12470);
nand U18860 (N_18860,N_15844,N_13662);
nand U18861 (N_18861,N_14182,N_13847);
and U18862 (N_18862,N_12250,N_15521);
nor U18863 (N_18863,N_13317,N_13682);
or U18864 (N_18864,N_14301,N_13345);
and U18865 (N_18865,N_14232,N_13420);
nand U18866 (N_18866,N_12432,N_14243);
nand U18867 (N_18867,N_15422,N_12850);
nor U18868 (N_18868,N_13352,N_13672);
xnor U18869 (N_18869,N_12448,N_14361);
or U18870 (N_18870,N_15256,N_14102);
nor U18871 (N_18871,N_15273,N_13829);
or U18872 (N_18872,N_12587,N_14591);
or U18873 (N_18873,N_15795,N_13315);
or U18874 (N_18874,N_13458,N_13171);
and U18875 (N_18875,N_12341,N_12313);
and U18876 (N_18876,N_15903,N_12419);
nand U18877 (N_18877,N_12082,N_13968);
nor U18878 (N_18878,N_14678,N_13202);
nand U18879 (N_18879,N_13107,N_13780);
and U18880 (N_18880,N_12795,N_12324);
and U18881 (N_18881,N_14510,N_12840);
or U18882 (N_18882,N_12437,N_12753);
nor U18883 (N_18883,N_13337,N_15760);
nor U18884 (N_18884,N_14225,N_12094);
or U18885 (N_18885,N_15040,N_13870);
or U18886 (N_18886,N_15564,N_14823);
nor U18887 (N_18887,N_12245,N_15043);
nor U18888 (N_18888,N_13768,N_14487);
xnor U18889 (N_18889,N_14987,N_12096);
nor U18890 (N_18890,N_13451,N_15152);
or U18891 (N_18891,N_12505,N_14263);
nor U18892 (N_18892,N_13639,N_13507);
or U18893 (N_18893,N_12852,N_15940);
or U18894 (N_18894,N_13975,N_13356);
and U18895 (N_18895,N_12571,N_14660);
or U18896 (N_18896,N_15336,N_15219);
nand U18897 (N_18897,N_14191,N_14258);
or U18898 (N_18898,N_12120,N_12496);
xor U18899 (N_18899,N_13967,N_15057);
nor U18900 (N_18900,N_13341,N_15340);
nand U18901 (N_18901,N_12171,N_14562);
and U18902 (N_18902,N_13010,N_13176);
or U18903 (N_18903,N_15844,N_12226);
and U18904 (N_18904,N_14160,N_14392);
nor U18905 (N_18905,N_14150,N_15945);
and U18906 (N_18906,N_13204,N_13952);
or U18907 (N_18907,N_13300,N_14030);
or U18908 (N_18908,N_14166,N_12779);
nor U18909 (N_18909,N_14658,N_13577);
or U18910 (N_18910,N_15748,N_13824);
and U18911 (N_18911,N_15025,N_14899);
xnor U18912 (N_18912,N_12594,N_15371);
xnor U18913 (N_18913,N_13149,N_13905);
and U18914 (N_18914,N_12211,N_15162);
nor U18915 (N_18915,N_14163,N_15540);
nand U18916 (N_18916,N_14668,N_13187);
xnor U18917 (N_18917,N_14240,N_12668);
or U18918 (N_18918,N_14808,N_14267);
nor U18919 (N_18919,N_13638,N_12705);
nor U18920 (N_18920,N_15238,N_15284);
and U18921 (N_18921,N_15393,N_14662);
or U18922 (N_18922,N_12515,N_12069);
and U18923 (N_18923,N_14750,N_14600);
nor U18924 (N_18924,N_12413,N_12338);
or U18925 (N_18925,N_15606,N_13757);
and U18926 (N_18926,N_13914,N_15835);
nand U18927 (N_18927,N_15963,N_15327);
and U18928 (N_18928,N_13245,N_15872);
xor U18929 (N_18929,N_12825,N_14056);
and U18930 (N_18930,N_13614,N_14536);
nor U18931 (N_18931,N_15668,N_15764);
and U18932 (N_18932,N_15514,N_15942);
nand U18933 (N_18933,N_13883,N_12467);
nor U18934 (N_18934,N_14143,N_12263);
nand U18935 (N_18935,N_15118,N_13503);
nand U18936 (N_18936,N_15132,N_12046);
xor U18937 (N_18937,N_12734,N_12592);
and U18938 (N_18938,N_14500,N_13882);
nand U18939 (N_18939,N_12832,N_12859);
or U18940 (N_18940,N_15835,N_12619);
nor U18941 (N_18941,N_12330,N_13065);
nand U18942 (N_18942,N_14996,N_14864);
or U18943 (N_18943,N_12283,N_12469);
and U18944 (N_18944,N_12896,N_14550);
nor U18945 (N_18945,N_12868,N_12628);
nor U18946 (N_18946,N_12048,N_15764);
and U18947 (N_18947,N_12209,N_12653);
nor U18948 (N_18948,N_15849,N_14628);
nand U18949 (N_18949,N_15287,N_15659);
nor U18950 (N_18950,N_15167,N_13477);
and U18951 (N_18951,N_12262,N_15140);
and U18952 (N_18952,N_15915,N_14182);
xor U18953 (N_18953,N_15172,N_12278);
and U18954 (N_18954,N_12479,N_15074);
nand U18955 (N_18955,N_13872,N_12561);
and U18956 (N_18956,N_13348,N_12791);
nand U18957 (N_18957,N_12146,N_14932);
nand U18958 (N_18958,N_15853,N_13631);
or U18959 (N_18959,N_12329,N_14137);
and U18960 (N_18960,N_15518,N_14275);
and U18961 (N_18961,N_14049,N_15047);
and U18962 (N_18962,N_12612,N_13352);
or U18963 (N_18963,N_12117,N_13333);
nand U18964 (N_18964,N_14207,N_12428);
nand U18965 (N_18965,N_12791,N_13741);
nand U18966 (N_18966,N_13573,N_12762);
nor U18967 (N_18967,N_15338,N_15595);
nand U18968 (N_18968,N_12290,N_13408);
xnor U18969 (N_18969,N_15194,N_12802);
nand U18970 (N_18970,N_14149,N_15726);
nand U18971 (N_18971,N_13480,N_15976);
nor U18972 (N_18972,N_12064,N_15363);
and U18973 (N_18973,N_15678,N_15307);
nand U18974 (N_18974,N_15478,N_13399);
or U18975 (N_18975,N_14126,N_14436);
or U18976 (N_18976,N_12915,N_13090);
and U18977 (N_18977,N_13549,N_12082);
or U18978 (N_18978,N_15037,N_13096);
xor U18979 (N_18979,N_12362,N_15416);
and U18980 (N_18980,N_13261,N_13602);
and U18981 (N_18981,N_13346,N_12341);
or U18982 (N_18982,N_14537,N_13672);
or U18983 (N_18983,N_15411,N_15293);
nand U18984 (N_18984,N_13336,N_13760);
or U18985 (N_18985,N_12695,N_13713);
nand U18986 (N_18986,N_14918,N_12651);
nand U18987 (N_18987,N_13279,N_14545);
nand U18988 (N_18988,N_15794,N_14107);
or U18989 (N_18989,N_14109,N_13307);
or U18990 (N_18990,N_12746,N_13587);
nor U18991 (N_18991,N_12469,N_15413);
or U18992 (N_18992,N_13802,N_15570);
or U18993 (N_18993,N_12035,N_14985);
and U18994 (N_18994,N_15926,N_14236);
nor U18995 (N_18995,N_12660,N_12941);
xor U18996 (N_18996,N_13106,N_13632);
xor U18997 (N_18997,N_13175,N_13827);
or U18998 (N_18998,N_15398,N_14769);
and U18999 (N_18999,N_12094,N_13835);
xor U19000 (N_19000,N_15685,N_15281);
and U19001 (N_19001,N_15364,N_15946);
and U19002 (N_19002,N_13596,N_14742);
nor U19003 (N_19003,N_15382,N_15249);
and U19004 (N_19004,N_14697,N_14459);
or U19005 (N_19005,N_13875,N_13629);
nand U19006 (N_19006,N_12625,N_12247);
and U19007 (N_19007,N_14482,N_12483);
or U19008 (N_19008,N_12313,N_12041);
and U19009 (N_19009,N_14589,N_15671);
nor U19010 (N_19010,N_14428,N_14720);
and U19011 (N_19011,N_14844,N_14696);
and U19012 (N_19012,N_13739,N_15603);
nor U19013 (N_19013,N_14042,N_14473);
and U19014 (N_19014,N_15839,N_12788);
nor U19015 (N_19015,N_15841,N_13911);
or U19016 (N_19016,N_14813,N_13916);
and U19017 (N_19017,N_15823,N_14167);
and U19018 (N_19018,N_14263,N_15350);
nor U19019 (N_19019,N_12500,N_14771);
xor U19020 (N_19020,N_15829,N_15868);
nor U19021 (N_19021,N_15698,N_14656);
or U19022 (N_19022,N_15441,N_12188);
nor U19023 (N_19023,N_14143,N_12057);
and U19024 (N_19024,N_14662,N_14210);
and U19025 (N_19025,N_12088,N_15136);
nor U19026 (N_19026,N_15176,N_14344);
nand U19027 (N_19027,N_13797,N_12103);
xnor U19028 (N_19028,N_15359,N_12718);
nand U19029 (N_19029,N_13790,N_13530);
nand U19030 (N_19030,N_13383,N_15319);
and U19031 (N_19031,N_14024,N_15583);
nor U19032 (N_19032,N_15680,N_14763);
and U19033 (N_19033,N_13552,N_12038);
xor U19034 (N_19034,N_15943,N_14582);
and U19035 (N_19035,N_12869,N_12817);
or U19036 (N_19036,N_14997,N_12725);
and U19037 (N_19037,N_13364,N_15257);
nand U19038 (N_19038,N_13027,N_13309);
nand U19039 (N_19039,N_15618,N_14805);
nand U19040 (N_19040,N_12174,N_14708);
and U19041 (N_19041,N_13069,N_12952);
nand U19042 (N_19042,N_15159,N_14855);
xnor U19043 (N_19043,N_14459,N_14142);
nand U19044 (N_19044,N_14018,N_14659);
and U19045 (N_19045,N_12758,N_13146);
or U19046 (N_19046,N_15574,N_14275);
and U19047 (N_19047,N_14267,N_12389);
nor U19048 (N_19048,N_12842,N_14460);
and U19049 (N_19049,N_14405,N_12051);
nand U19050 (N_19050,N_13998,N_13512);
nor U19051 (N_19051,N_14224,N_12077);
nand U19052 (N_19052,N_12364,N_13919);
and U19053 (N_19053,N_12708,N_15328);
nand U19054 (N_19054,N_14811,N_15911);
nand U19055 (N_19055,N_12069,N_12550);
nand U19056 (N_19056,N_15960,N_14342);
and U19057 (N_19057,N_14085,N_13726);
nand U19058 (N_19058,N_13940,N_12126);
nor U19059 (N_19059,N_13061,N_13907);
nor U19060 (N_19060,N_15060,N_13711);
nand U19061 (N_19061,N_15488,N_14593);
or U19062 (N_19062,N_14942,N_12138);
xnor U19063 (N_19063,N_14234,N_13823);
or U19064 (N_19064,N_15529,N_15462);
or U19065 (N_19065,N_15105,N_15636);
and U19066 (N_19066,N_15189,N_12204);
nand U19067 (N_19067,N_13627,N_12568);
nand U19068 (N_19068,N_15626,N_14435);
nor U19069 (N_19069,N_12591,N_12945);
nand U19070 (N_19070,N_15189,N_12945);
nand U19071 (N_19071,N_15896,N_12788);
and U19072 (N_19072,N_13744,N_12359);
or U19073 (N_19073,N_14457,N_12216);
or U19074 (N_19074,N_12395,N_15622);
nor U19075 (N_19075,N_13507,N_13975);
xnor U19076 (N_19076,N_14104,N_15727);
or U19077 (N_19077,N_14380,N_15388);
or U19078 (N_19078,N_14680,N_15983);
nor U19079 (N_19079,N_13912,N_14140);
xor U19080 (N_19080,N_12401,N_13000);
nand U19081 (N_19081,N_13086,N_12862);
and U19082 (N_19082,N_15771,N_13138);
and U19083 (N_19083,N_13453,N_14174);
and U19084 (N_19084,N_13860,N_14521);
or U19085 (N_19085,N_15548,N_14116);
xor U19086 (N_19086,N_14245,N_15893);
nor U19087 (N_19087,N_14675,N_12587);
nor U19088 (N_19088,N_14924,N_14494);
and U19089 (N_19089,N_14980,N_14557);
or U19090 (N_19090,N_12112,N_14132);
nor U19091 (N_19091,N_15905,N_15644);
nand U19092 (N_19092,N_12881,N_12578);
nand U19093 (N_19093,N_13222,N_13553);
nand U19094 (N_19094,N_13351,N_15544);
nor U19095 (N_19095,N_13583,N_15708);
or U19096 (N_19096,N_15072,N_12807);
and U19097 (N_19097,N_14478,N_12482);
nor U19098 (N_19098,N_12986,N_12595);
xnor U19099 (N_19099,N_15140,N_12099);
or U19100 (N_19100,N_13015,N_12615);
and U19101 (N_19101,N_14184,N_15025);
nor U19102 (N_19102,N_14788,N_14458);
or U19103 (N_19103,N_15656,N_14537);
or U19104 (N_19104,N_14962,N_12349);
nor U19105 (N_19105,N_13766,N_14359);
nor U19106 (N_19106,N_14248,N_14055);
or U19107 (N_19107,N_15744,N_15637);
nor U19108 (N_19108,N_13441,N_12178);
nor U19109 (N_19109,N_14744,N_12940);
nor U19110 (N_19110,N_14567,N_12624);
nand U19111 (N_19111,N_14410,N_14362);
or U19112 (N_19112,N_15262,N_13741);
or U19113 (N_19113,N_14335,N_12259);
and U19114 (N_19114,N_14624,N_15162);
or U19115 (N_19115,N_13221,N_15434);
and U19116 (N_19116,N_13632,N_14967);
nand U19117 (N_19117,N_15341,N_15306);
and U19118 (N_19118,N_13778,N_15973);
or U19119 (N_19119,N_14157,N_14956);
nor U19120 (N_19120,N_15892,N_12586);
nand U19121 (N_19121,N_14361,N_14156);
and U19122 (N_19122,N_15998,N_12914);
nor U19123 (N_19123,N_14677,N_14389);
and U19124 (N_19124,N_13830,N_12729);
nand U19125 (N_19125,N_15989,N_15951);
nor U19126 (N_19126,N_14742,N_14204);
or U19127 (N_19127,N_12463,N_13174);
and U19128 (N_19128,N_15019,N_13257);
or U19129 (N_19129,N_14957,N_15120);
or U19130 (N_19130,N_13877,N_14840);
nor U19131 (N_19131,N_15886,N_14257);
and U19132 (N_19132,N_13240,N_15194);
nor U19133 (N_19133,N_14028,N_14892);
xor U19134 (N_19134,N_13143,N_15489);
and U19135 (N_19135,N_15309,N_14504);
and U19136 (N_19136,N_14151,N_14051);
xor U19137 (N_19137,N_13200,N_13701);
nand U19138 (N_19138,N_12881,N_14588);
nand U19139 (N_19139,N_12282,N_13730);
nand U19140 (N_19140,N_13072,N_15544);
nand U19141 (N_19141,N_14495,N_15934);
nor U19142 (N_19142,N_12131,N_14098);
xor U19143 (N_19143,N_13815,N_12010);
xnor U19144 (N_19144,N_12884,N_14758);
nor U19145 (N_19145,N_15180,N_12043);
or U19146 (N_19146,N_14250,N_14152);
and U19147 (N_19147,N_14448,N_15547);
nor U19148 (N_19148,N_14596,N_13488);
nor U19149 (N_19149,N_14904,N_14342);
and U19150 (N_19150,N_15741,N_15618);
or U19151 (N_19151,N_14343,N_14828);
or U19152 (N_19152,N_12564,N_15674);
or U19153 (N_19153,N_14437,N_14451);
nand U19154 (N_19154,N_13821,N_14062);
nor U19155 (N_19155,N_13156,N_13386);
nand U19156 (N_19156,N_15610,N_13492);
nor U19157 (N_19157,N_15730,N_12893);
and U19158 (N_19158,N_12132,N_13411);
and U19159 (N_19159,N_12402,N_15176);
xnor U19160 (N_19160,N_14618,N_14068);
nand U19161 (N_19161,N_14133,N_14974);
nand U19162 (N_19162,N_14343,N_15402);
nand U19163 (N_19163,N_12669,N_12116);
nand U19164 (N_19164,N_12294,N_14521);
and U19165 (N_19165,N_14576,N_15788);
and U19166 (N_19166,N_14945,N_12781);
nor U19167 (N_19167,N_14162,N_13975);
nand U19168 (N_19168,N_14496,N_13857);
nand U19169 (N_19169,N_15224,N_12289);
or U19170 (N_19170,N_15485,N_12114);
or U19171 (N_19171,N_15245,N_14383);
and U19172 (N_19172,N_14058,N_14393);
xor U19173 (N_19173,N_15233,N_14316);
nand U19174 (N_19174,N_15109,N_14376);
and U19175 (N_19175,N_14109,N_15037);
and U19176 (N_19176,N_15262,N_15051);
and U19177 (N_19177,N_13850,N_14643);
and U19178 (N_19178,N_12541,N_13674);
xnor U19179 (N_19179,N_12765,N_14828);
nor U19180 (N_19180,N_14862,N_13308);
nand U19181 (N_19181,N_12262,N_13561);
or U19182 (N_19182,N_14653,N_13668);
and U19183 (N_19183,N_12475,N_12679);
xor U19184 (N_19184,N_12399,N_14161);
or U19185 (N_19185,N_12381,N_12178);
or U19186 (N_19186,N_15653,N_15451);
or U19187 (N_19187,N_12741,N_15910);
nor U19188 (N_19188,N_15924,N_12629);
and U19189 (N_19189,N_14342,N_12596);
nand U19190 (N_19190,N_12077,N_13570);
and U19191 (N_19191,N_12766,N_14365);
and U19192 (N_19192,N_14030,N_14221);
and U19193 (N_19193,N_13070,N_14305);
and U19194 (N_19194,N_13658,N_14947);
or U19195 (N_19195,N_14309,N_15002);
nor U19196 (N_19196,N_14233,N_14314);
and U19197 (N_19197,N_14352,N_13182);
nor U19198 (N_19198,N_13944,N_13162);
nor U19199 (N_19199,N_14639,N_13360);
or U19200 (N_19200,N_14213,N_12013);
nand U19201 (N_19201,N_13334,N_13744);
nand U19202 (N_19202,N_12900,N_12925);
nand U19203 (N_19203,N_15997,N_15626);
xor U19204 (N_19204,N_14961,N_13961);
nor U19205 (N_19205,N_15753,N_14051);
nor U19206 (N_19206,N_12958,N_15311);
nor U19207 (N_19207,N_12102,N_12202);
xnor U19208 (N_19208,N_14377,N_13798);
and U19209 (N_19209,N_14427,N_13915);
nand U19210 (N_19210,N_15701,N_13230);
nand U19211 (N_19211,N_13257,N_15434);
nand U19212 (N_19212,N_12583,N_15728);
xnor U19213 (N_19213,N_12706,N_13756);
xnor U19214 (N_19214,N_12491,N_14293);
and U19215 (N_19215,N_15909,N_15252);
and U19216 (N_19216,N_14256,N_15631);
nor U19217 (N_19217,N_12968,N_14958);
and U19218 (N_19218,N_14050,N_12988);
or U19219 (N_19219,N_12078,N_13358);
and U19220 (N_19220,N_13135,N_15367);
or U19221 (N_19221,N_13661,N_13596);
xor U19222 (N_19222,N_14276,N_15694);
xor U19223 (N_19223,N_12201,N_15231);
and U19224 (N_19224,N_14379,N_13106);
or U19225 (N_19225,N_15626,N_15675);
nand U19226 (N_19226,N_13297,N_12094);
nand U19227 (N_19227,N_15838,N_14716);
nand U19228 (N_19228,N_13298,N_15108);
xnor U19229 (N_19229,N_13514,N_12081);
and U19230 (N_19230,N_13883,N_15984);
xor U19231 (N_19231,N_15076,N_12333);
xor U19232 (N_19232,N_13904,N_12047);
nor U19233 (N_19233,N_13418,N_13698);
nand U19234 (N_19234,N_12753,N_14945);
nor U19235 (N_19235,N_15392,N_12048);
or U19236 (N_19236,N_13733,N_12365);
nand U19237 (N_19237,N_14610,N_13461);
or U19238 (N_19238,N_14732,N_14624);
nand U19239 (N_19239,N_15385,N_15624);
or U19240 (N_19240,N_15261,N_13117);
or U19241 (N_19241,N_14634,N_13792);
nor U19242 (N_19242,N_14358,N_15353);
and U19243 (N_19243,N_13383,N_15541);
nand U19244 (N_19244,N_13825,N_12038);
or U19245 (N_19245,N_12430,N_14066);
nor U19246 (N_19246,N_15830,N_12805);
xor U19247 (N_19247,N_15620,N_14496);
or U19248 (N_19248,N_14342,N_12828);
nand U19249 (N_19249,N_15004,N_14150);
nor U19250 (N_19250,N_15146,N_14228);
xnor U19251 (N_19251,N_13484,N_14025);
nand U19252 (N_19252,N_15515,N_12354);
nor U19253 (N_19253,N_12866,N_14907);
or U19254 (N_19254,N_15493,N_13876);
nor U19255 (N_19255,N_12906,N_14328);
nand U19256 (N_19256,N_13338,N_14579);
and U19257 (N_19257,N_14553,N_12155);
nand U19258 (N_19258,N_12719,N_14095);
or U19259 (N_19259,N_13453,N_13554);
or U19260 (N_19260,N_15283,N_12194);
and U19261 (N_19261,N_12457,N_14817);
or U19262 (N_19262,N_13497,N_14825);
nand U19263 (N_19263,N_14159,N_12576);
nor U19264 (N_19264,N_14356,N_13352);
xor U19265 (N_19265,N_15309,N_14884);
and U19266 (N_19266,N_13917,N_15836);
nand U19267 (N_19267,N_12644,N_13398);
or U19268 (N_19268,N_14993,N_14045);
nand U19269 (N_19269,N_15333,N_13731);
nor U19270 (N_19270,N_12401,N_13110);
nor U19271 (N_19271,N_12612,N_15488);
and U19272 (N_19272,N_13301,N_12521);
or U19273 (N_19273,N_12073,N_13789);
or U19274 (N_19274,N_14737,N_14333);
nor U19275 (N_19275,N_13554,N_14572);
nor U19276 (N_19276,N_15289,N_15038);
nor U19277 (N_19277,N_12183,N_12910);
xor U19278 (N_19278,N_13448,N_15276);
and U19279 (N_19279,N_12500,N_13417);
and U19280 (N_19280,N_13597,N_13159);
nand U19281 (N_19281,N_14791,N_15383);
nor U19282 (N_19282,N_15190,N_12039);
nand U19283 (N_19283,N_13463,N_15935);
and U19284 (N_19284,N_15056,N_15403);
xor U19285 (N_19285,N_14282,N_14098);
and U19286 (N_19286,N_12774,N_13349);
and U19287 (N_19287,N_15004,N_12065);
nand U19288 (N_19288,N_14468,N_13540);
or U19289 (N_19289,N_14858,N_12047);
nor U19290 (N_19290,N_13815,N_15178);
or U19291 (N_19291,N_13984,N_12930);
xnor U19292 (N_19292,N_12811,N_15646);
nand U19293 (N_19293,N_14171,N_12719);
or U19294 (N_19294,N_13890,N_14702);
and U19295 (N_19295,N_13048,N_15433);
nand U19296 (N_19296,N_14373,N_15172);
or U19297 (N_19297,N_13420,N_14473);
and U19298 (N_19298,N_13124,N_12684);
nor U19299 (N_19299,N_15928,N_12184);
nand U19300 (N_19300,N_14697,N_12043);
nand U19301 (N_19301,N_13571,N_15882);
and U19302 (N_19302,N_12074,N_15637);
or U19303 (N_19303,N_12855,N_14514);
xnor U19304 (N_19304,N_14864,N_15975);
nand U19305 (N_19305,N_13874,N_14794);
nor U19306 (N_19306,N_12837,N_13140);
nand U19307 (N_19307,N_14201,N_12852);
or U19308 (N_19308,N_14974,N_13843);
or U19309 (N_19309,N_15057,N_14621);
or U19310 (N_19310,N_14115,N_14828);
and U19311 (N_19311,N_12561,N_13243);
xor U19312 (N_19312,N_12182,N_13297);
nand U19313 (N_19313,N_14514,N_12444);
nand U19314 (N_19314,N_12665,N_15134);
xnor U19315 (N_19315,N_14989,N_12590);
nand U19316 (N_19316,N_12863,N_15449);
nor U19317 (N_19317,N_15769,N_12138);
nand U19318 (N_19318,N_13382,N_13554);
or U19319 (N_19319,N_15897,N_13948);
nand U19320 (N_19320,N_12425,N_15471);
or U19321 (N_19321,N_15399,N_12792);
xor U19322 (N_19322,N_13419,N_15428);
or U19323 (N_19323,N_14503,N_15109);
or U19324 (N_19324,N_14363,N_13207);
or U19325 (N_19325,N_15711,N_14148);
nor U19326 (N_19326,N_13026,N_15412);
and U19327 (N_19327,N_12624,N_13904);
or U19328 (N_19328,N_15855,N_13195);
or U19329 (N_19329,N_13008,N_15878);
and U19330 (N_19330,N_15298,N_14510);
nor U19331 (N_19331,N_14947,N_15004);
and U19332 (N_19332,N_13174,N_12046);
or U19333 (N_19333,N_13519,N_13900);
and U19334 (N_19334,N_15090,N_13912);
and U19335 (N_19335,N_12905,N_13689);
and U19336 (N_19336,N_13900,N_15467);
nor U19337 (N_19337,N_14978,N_12036);
xor U19338 (N_19338,N_15591,N_12893);
nand U19339 (N_19339,N_15750,N_13664);
nand U19340 (N_19340,N_12702,N_13626);
or U19341 (N_19341,N_12416,N_14829);
nor U19342 (N_19342,N_14424,N_14863);
nand U19343 (N_19343,N_15858,N_14230);
nand U19344 (N_19344,N_13678,N_12482);
nand U19345 (N_19345,N_12272,N_15185);
nand U19346 (N_19346,N_14841,N_13259);
xnor U19347 (N_19347,N_12450,N_14364);
and U19348 (N_19348,N_13946,N_14861);
and U19349 (N_19349,N_14914,N_15185);
nand U19350 (N_19350,N_13166,N_12402);
nor U19351 (N_19351,N_14876,N_12669);
nor U19352 (N_19352,N_13649,N_15164);
or U19353 (N_19353,N_15902,N_14213);
nor U19354 (N_19354,N_12258,N_14058);
and U19355 (N_19355,N_13005,N_13088);
nor U19356 (N_19356,N_12233,N_13926);
nor U19357 (N_19357,N_15830,N_12562);
nor U19358 (N_19358,N_15018,N_15928);
and U19359 (N_19359,N_14388,N_12528);
nor U19360 (N_19360,N_13343,N_14535);
nor U19361 (N_19361,N_15810,N_15951);
or U19362 (N_19362,N_12484,N_14075);
or U19363 (N_19363,N_14535,N_13289);
or U19364 (N_19364,N_13830,N_12342);
or U19365 (N_19365,N_15602,N_13287);
and U19366 (N_19366,N_15917,N_12123);
xnor U19367 (N_19367,N_14655,N_12055);
nor U19368 (N_19368,N_13582,N_12024);
xor U19369 (N_19369,N_13874,N_13409);
nand U19370 (N_19370,N_15061,N_13518);
nand U19371 (N_19371,N_15774,N_12595);
nand U19372 (N_19372,N_15321,N_14901);
nand U19373 (N_19373,N_12378,N_13697);
nor U19374 (N_19374,N_14529,N_14696);
xor U19375 (N_19375,N_15215,N_15151);
and U19376 (N_19376,N_15272,N_14739);
nand U19377 (N_19377,N_15125,N_14164);
xor U19378 (N_19378,N_15942,N_15688);
and U19379 (N_19379,N_13391,N_14418);
xnor U19380 (N_19380,N_12979,N_14576);
and U19381 (N_19381,N_12950,N_14123);
or U19382 (N_19382,N_13705,N_12677);
nor U19383 (N_19383,N_15850,N_14284);
nand U19384 (N_19384,N_14329,N_14209);
xor U19385 (N_19385,N_12127,N_15724);
or U19386 (N_19386,N_14631,N_14396);
or U19387 (N_19387,N_15034,N_13763);
nor U19388 (N_19388,N_13549,N_13191);
nand U19389 (N_19389,N_14278,N_14822);
nand U19390 (N_19390,N_14741,N_12856);
nor U19391 (N_19391,N_12192,N_14845);
or U19392 (N_19392,N_14242,N_14424);
nor U19393 (N_19393,N_12108,N_13358);
nand U19394 (N_19394,N_12857,N_15224);
nor U19395 (N_19395,N_15494,N_15037);
nand U19396 (N_19396,N_12808,N_13202);
nand U19397 (N_19397,N_12051,N_13977);
and U19398 (N_19398,N_12978,N_12867);
nand U19399 (N_19399,N_14104,N_15919);
and U19400 (N_19400,N_12319,N_13479);
xnor U19401 (N_19401,N_12249,N_14206);
nor U19402 (N_19402,N_13618,N_12467);
or U19403 (N_19403,N_15195,N_12973);
and U19404 (N_19404,N_13465,N_13684);
or U19405 (N_19405,N_13548,N_13206);
or U19406 (N_19406,N_13352,N_14764);
nand U19407 (N_19407,N_13512,N_14950);
or U19408 (N_19408,N_14924,N_12610);
and U19409 (N_19409,N_15979,N_12691);
nand U19410 (N_19410,N_12421,N_15321);
nor U19411 (N_19411,N_12147,N_15569);
nor U19412 (N_19412,N_15066,N_12549);
and U19413 (N_19413,N_15237,N_12092);
nor U19414 (N_19414,N_14893,N_15301);
nor U19415 (N_19415,N_15261,N_14975);
or U19416 (N_19416,N_13796,N_13346);
nor U19417 (N_19417,N_14321,N_14761);
nand U19418 (N_19418,N_13244,N_14413);
nor U19419 (N_19419,N_15664,N_12318);
nand U19420 (N_19420,N_12119,N_15523);
or U19421 (N_19421,N_13450,N_13886);
or U19422 (N_19422,N_14364,N_14901);
nand U19423 (N_19423,N_14644,N_13764);
or U19424 (N_19424,N_15561,N_14708);
nor U19425 (N_19425,N_15342,N_14572);
and U19426 (N_19426,N_13619,N_13297);
or U19427 (N_19427,N_15431,N_13253);
or U19428 (N_19428,N_15338,N_13079);
or U19429 (N_19429,N_13630,N_15571);
nor U19430 (N_19430,N_12628,N_15396);
and U19431 (N_19431,N_15691,N_13513);
nor U19432 (N_19432,N_12107,N_13153);
nor U19433 (N_19433,N_12029,N_12774);
nor U19434 (N_19434,N_15199,N_12497);
nand U19435 (N_19435,N_14564,N_15101);
nor U19436 (N_19436,N_15927,N_14183);
nor U19437 (N_19437,N_12669,N_14737);
and U19438 (N_19438,N_12843,N_15085);
and U19439 (N_19439,N_14708,N_13475);
nand U19440 (N_19440,N_14118,N_12177);
nor U19441 (N_19441,N_13840,N_15928);
or U19442 (N_19442,N_13260,N_15649);
or U19443 (N_19443,N_12836,N_12050);
or U19444 (N_19444,N_15012,N_14197);
nor U19445 (N_19445,N_13739,N_12732);
or U19446 (N_19446,N_12565,N_12262);
and U19447 (N_19447,N_12293,N_14030);
nand U19448 (N_19448,N_14880,N_13484);
and U19449 (N_19449,N_12598,N_12786);
or U19450 (N_19450,N_12137,N_12439);
or U19451 (N_19451,N_14062,N_14544);
nor U19452 (N_19452,N_13787,N_13349);
xnor U19453 (N_19453,N_15427,N_15390);
or U19454 (N_19454,N_12169,N_15158);
xnor U19455 (N_19455,N_15233,N_15852);
nand U19456 (N_19456,N_13910,N_14128);
or U19457 (N_19457,N_13763,N_13695);
nor U19458 (N_19458,N_15594,N_14321);
nor U19459 (N_19459,N_12731,N_13685);
nor U19460 (N_19460,N_15807,N_12102);
nor U19461 (N_19461,N_13594,N_14108);
xor U19462 (N_19462,N_14697,N_14912);
or U19463 (N_19463,N_12510,N_15077);
xnor U19464 (N_19464,N_15951,N_14737);
nand U19465 (N_19465,N_13500,N_13073);
nand U19466 (N_19466,N_12111,N_14784);
or U19467 (N_19467,N_13922,N_12952);
or U19468 (N_19468,N_12056,N_13429);
or U19469 (N_19469,N_12444,N_14432);
and U19470 (N_19470,N_13637,N_12313);
or U19471 (N_19471,N_13841,N_14821);
nand U19472 (N_19472,N_12038,N_12995);
or U19473 (N_19473,N_15273,N_13180);
or U19474 (N_19474,N_15087,N_14483);
and U19475 (N_19475,N_12402,N_12835);
nor U19476 (N_19476,N_13789,N_14890);
nor U19477 (N_19477,N_15881,N_14141);
nand U19478 (N_19478,N_13966,N_13110);
and U19479 (N_19479,N_15855,N_12343);
and U19480 (N_19480,N_14809,N_12415);
and U19481 (N_19481,N_14048,N_12318);
or U19482 (N_19482,N_14260,N_12614);
and U19483 (N_19483,N_12574,N_13293);
and U19484 (N_19484,N_14628,N_14110);
nand U19485 (N_19485,N_14135,N_14700);
and U19486 (N_19486,N_13803,N_15264);
xnor U19487 (N_19487,N_12920,N_14834);
and U19488 (N_19488,N_14487,N_12378);
xnor U19489 (N_19489,N_13771,N_15911);
xor U19490 (N_19490,N_12312,N_15252);
or U19491 (N_19491,N_12117,N_14346);
xnor U19492 (N_19492,N_12247,N_15790);
or U19493 (N_19493,N_13876,N_15967);
nor U19494 (N_19494,N_15751,N_14227);
nor U19495 (N_19495,N_15359,N_14418);
or U19496 (N_19496,N_14399,N_13906);
xor U19497 (N_19497,N_12794,N_15195);
nand U19498 (N_19498,N_15457,N_14181);
nor U19499 (N_19499,N_15187,N_14438);
or U19500 (N_19500,N_12486,N_13819);
and U19501 (N_19501,N_14367,N_12376);
or U19502 (N_19502,N_13844,N_15405);
or U19503 (N_19503,N_14203,N_15365);
or U19504 (N_19504,N_15959,N_13064);
xnor U19505 (N_19505,N_15071,N_12277);
and U19506 (N_19506,N_14638,N_15347);
or U19507 (N_19507,N_14859,N_14162);
or U19508 (N_19508,N_14164,N_14702);
nand U19509 (N_19509,N_13243,N_13261);
nand U19510 (N_19510,N_14245,N_12837);
or U19511 (N_19511,N_13067,N_14838);
xor U19512 (N_19512,N_14973,N_15000);
or U19513 (N_19513,N_15244,N_14764);
or U19514 (N_19514,N_12464,N_12310);
or U19515 (N_19515,N_14469,N_14855);
nor U19516 (N_19516,N_13335,N_14633);
nand U19517 (N_19517,N_12244,N_12431);
and U19518 (N_19518,N_15598,N_14521);
nor U19519 (N_19519,N_14871,N_14170);
nand U19520 (N_19520,N_14933,N_15818);
nand U19521 (N_19521,N_12536,N_15906);
or U19522 (N_19522,N_15033,N_13051);
or U19523 (N_19523,N_13003,N_14963);
nor U19524 (N_19524,N_12152,N_12632);
and U19525 (N_19525,N_12219,N_15649);
and U19526 (N_19526,N_14137,N_14383);
nor U19527 (N_19527,N_12392,N_13770);
and U19528 (N_19528,N_14629,N_13762);
xnor U19529 (N_19529,N_12605,N_14231);
or U19530 (N_19530,N_12248,N_13758);
or U19531 (N_19531,N_12278,N_14934);
nor U19532 (N_19532,N_12684,N_12413);
nand U19533 (N_19533,N_15486,N_13458);
or U19534 (N_19534,N_13143,N_13781);
nor U19535 (N_19535,N_14474,N_13652);
xor U19536 (N_19536,N_13548,N_13949);
or U19537 (N_19537,N_13881,N_14546);
or U19538 (N_19538,N_12139,N_13117);
nand U19539 (N_19539,N_12145,N_13750);
or U19540 (N_19540,N_13264,N_12382);
nand U19541 (N_19541,N_14395,N_12117);
nand U19542 (N_19542,N_14409,N_15436);
and U19543 (N_19543,N_12821,N_13069);
or U19544 (N_19544,N_13260,N_15018);
nand U19545 (N_19545,N_14648,N_15503);
or U19546 (N_19546,N_13351,N_13746);
or U19547 (N_19547,N_12533,N_13588);
or U19548 (N_19548,N_15966,N_12640);
or U19549 (N_19549,N_15852,N_12647);
nand U19550 (N_19550,N_15520,N_14348);
nand U19551 (N_19551,N_12253,N_12815);
and U19552 (N_19552,N_13590,N_13650);
nand U19553 (N_19553,N_12030,N_15290);
or U19554 (N_19554,N_12663,N_14149);
nor U19555 (N_19555,N_15829,N_15505);
or U19556 (N_19556,N_14629,N_12493);
or U19557 (N_19557,N_12273,N_12920);
and U19558 (N_19558,N_12159,N_15423);
or U19559 (N_19559,N_13407,N_12348);
and U19560 (N_19560,N_13697,N_15065);
xnor U19561 (N_19561,N_13426,N_13690);
or U19562 (N_19562,N_12198,N_13727);
nor U19563 (N_19563,N_15094,N_12851);
nand U19564 (N_19564,N_15683,N_13572);
and U19565 (N_19565,N_15332,N_14336);
and U19566 (N_19566,N_12176,N_15196);
and U19567 (N_19567,N_14425,N_12495);
or U19568 (N_19568,N_13816,N_15068);
and U19569 (N_19569,N_15749,N_13210);
nor U19570 (N_19570,N_14500,N_15371);
or U19571 (N_19571,N_14031,N_14230);
nand U19572 (N_19572,N_15996,N_14891);
nand U19573 (N_19573,N_12631,N_13286);
nor U19574 (N_19574,N_13321,N_13666);
and U19575 (N_19575,N_15886,N_15381);
nor U19576 (N_19576,N_14711,N_13334);
nand U19577 (N_19577,N_14401,N_15792);
and U19578 (N_19578,N_15520,N_15753);
nor U19579 (N_19579,N_14422,N_15453);
xnor U19580 (N_19580,N_14886,N_15618);
or U19581 (N_19581,N_12031,N_14351);
or U19582 (N_19582,N_15192,N_13570);
nand U19583 (N_19583,N_12833,N_14926);
xor U19584 (N_19584,N_12280,N_13493);
and U19585 (N_19585,N_13026,N_14360);
or U19586 (N_19586,N_14795,N_12341);
and U19587 (N_19587,N_14708,N_13550);
nor U19588 (N_19588,N_12962,N_15119);
or U19589 (N_19589,N_15140,N_14762);
nor U19590 (N_19590,N_14666,N_12789);
nand U19591 (N_19591,N_13353,N_13697);
nor U19592 (N_19592,N_13398,N_14015);
or U19593 (N_19593,N_14440,N_13728);
xor U19594 (N_19594,N_15096,N_14565);
nand U19595 (N_19595,N_12557,N_15715);
and U19596 (N_19596,N_15091,N_14399);
and U19597 (N_19597,N_15128,N_12699);
or U19598 (N_19598,N_14045,N_14831);
and U19599 (N_19599,N_14702,N_12525);
and U19600 (N_19600,N_13991,N_12149);
or U19601 (N_19601,N_14608,N_15718);
nand U19602 (N_19602,N_15301,N_12622);
nand U19603 (N_19603,N_13298,N_14303);
nor U19604 (N_19604,N_12943,N_14716);
and U19605 (N_19605,N_12818,N_12886);
nor U19606 (N_19606,N_13148,N_14064);
nand U19607 (N_19607,N_12681,N_15967);
nand U19608 (N_19608,N_13448,N_12089);
and U19609 (N_19609,N_13530,N_12414);
nor U19610 (N_19610,N_14061,N_12169);
xor U19611 (N_19611,N_13140,N_13702);
or U19612 (N_19612,N_13332,N_14216);
nor U19613 (N_19613,N_13558,N_13776);
or U19614 (N_19614,N_14470,N_13329);
nand U19615 (N_19615,N_12682,N_12737);
nor U19616 (N_19616,N_14160,N_13917);
or U19617 (N_19617,N_12296,N_14015);
or U19618 (N_19618,N_12029,N_13935);
nor U19619 (N_19619,N_12197,N_14863);
and U19620 (N_19620,N_13481,N_15405);
xor U19621 (N_19621,N_14444,N_15558);
nor U19622 (N_19622,N_14657,N_12521);
or U19623 (N_19623,N_14911,N_14324);
xor U19624 (N_19624,N_14829,N_12297);
and U19625 (N_19625,N_14586,N_14680);
or U19626 (N_19626,N_13649,N_13869);
and U19627 (N_19627,N_13194,N_15325);
and U19628 (N_19628,N_12900,N_14574);
and U19629 (N_19629,N_13312,N_15647);
or U19630 (N_19630,N_13761,N_14653);
nor U19631 (N_19631,N_14489,N_12728);
nand U19632 (N_19632,N_15518,N_15952);
nand U19633 (N_19633,N_14649,N_12804);
nand U19634 (N_19634,N_14792,N_15024);
xor U19635 (N_19635,N_14408,N_15600);
and U19636 (N_19636,N_12751,N_14491);
nand U19637 (N_19637,N_15983,N_12915);
nor U19638 (N_19638,N_13580,N_12660);
nand U19639 (N_19639,N_14195,N_12957);
nor U19640 (N_19640,N_15132,N_13098);
and U19641 (N_19641,N_13503,N_15342);
nor U19642 (N_19642,N_12542,N_13577);
and U19643 (N_19643,N_14930,N_13674);
and U19644 (N_19644,N_15169,N_13766);
nand U19645 (N_19645,N_13716,N_14899);
or U19646 (N_19646,N_12248,N_14131);
and U19647 (N_19647,N_12819,N_15110);
nand U19648 (N_19648,N_14995,N_15137);
or U19649 (N_19649,N_13800,N_15586);
or U19650 (N_19650,N_12762,N_13394);
and U19651 (N_19651,N_15346,N_14635);
nand U19652 (N_19652,N_15271,N_15380);
xnor U19653 (N_19653,N_14575,N_15055);
and U19654 (N_19654,N_15415,N_15273);
and U19655 (N_19655,N_12920,N_14181);
nand U19656 (N_19656,N_12196,N_15412);
or U19657 (N_19657,N_13257,N_15363);
or U19658 (N_19658,N_13231,N_12366);
and U19659 (N_19659,N_15662,N_14508);
or U19660 (N_19660,N_15664,N_12355);
nor U19661 (N_19661,N_15049,N_14745);
xnor U19662 (N_19662,N_12419,N_13334);
nand U19663 (N_19663,N_14324,N_15572);
or U19664 (N_19664,N_15168,N_15423);
or U19665 (N_19665,N_15124,N_15217);
nand U19666 (N_19666,N_12134,N_13503);
nor U19667 (N_19667,N_15311,N_15857);
or U19668 (N_19668,N_15501,N_15962);
and U19669 (N_19669,N_14456,N_15259);
nand U19670 (N_19670,N_13242,N_15651);
or U19671 (N_19671,N_14275,N_15312);
and U19672 (N_19672,N_15834,N_15318);
and U19673 (N_19673,N_14956,N_12351);
and U19674 (N_19674,N_15475,N_13083);
nand U19675 (N_19675,N_13262,N_13976);
nand U19676 (N_19676,N_12858,N_14070);
nand U19677 (N_19677,N_12648,N_13412);
nor U19678 (N_19678,N_13404,N_12124);
and U19679 (N_19679,N_15138,N_15662);
and U19680 (N_19680,N_12790,N_15412);
nand U19681 (N_19681,N_14749,N_12730);
or U19682 (N_19682,N_13074,N_14681);
and U19683 (N_19683,N_15463,N_15557);
and U19684 (N_19684,N_15600,N_14426);
nand U19685 (N_19685,N_15870,N_13518);
nand U19686 (N_19686,N_12767,N_12375);
or U19687 (N_19687,N_13419,N_12240);
and U19688 (N_19688,N_12725,N_15361);
nand U19689 (N_19689,N_15001,N_13446);
xor U19690 (N_19690,N_14009,N_13509);
nor U19691 (N_19691,N_13953,N_12078);
or U19692 (N_19692,N_14161,N_12022);
and U19693 (N_19693,N_15267,N_14943);
nand U19694 (N_19694,N_14942,N_15900);
nor U19695 (N_19695,N_15753,N_13735);
or U19696 (N_19696,N_15580,N_13048);
and U19697 (N_19697,N_12925,N_12513);
nand U19698 (N_19698,N_14958,N_15005);
nand U19699 (N_19699,N_14654,N_14318);
and U19700 (N_19700,N_13410,N_14256);
nor U19701 (N_19701,N_13852,N_13967);
nand U19702 (N_19702,N_13586,N_14039);
xor U19703 (N_19703,N_15063,N_13414);
nor U19704 (N_19704,N_13693,N_15495);
xnor U19705 (N_19705,N_14715,N_12477);
nand U19706 (N_19706,N_13793,N_12791);
nor U19707 (N_19707,N_15498,N_15894);
nor U19708 (N_19708,N_13548,N_15859);
nor U19709 (N_19709,N_13218,N_15749);
nor U19710 (N_19710,N_14199,N_14946);
nand U19711 (N_19711,N_15034,N_14389);
nor U19712 (N_19712,N_14676,N_14824);
nor U19713 (N_19713,N_12643,N_13722);
or U19714 (N_19714,N_14204,N_12561);
nand U19715 (N_19715,N_15921,N_15774);
xnor U19716 (N_19716,N_14055,N_15637);
or U19717 (N_19717,N_14439,N_14677);
xor U19718 (N_19718,N_12323,N_13064);
xor U19719 (N_19719,N_14092,N_14205);
nand U19720 (N_19720,N_13459,N_12700);
and U19721 (N_19721,N_12366,N_13221);
or U19722 (N_19722,N_12690,N_15277);
nor U19723 (N_19723,N_14494,N_12716);
and U19724 (N_19724,N_12252,N_12665);
and U19725 (N_19725,N_13518,N_15929);
xor U19726 (N_19726,N_15725,N_14263);
nand U19727 (N_19727,N_12659,N_15404);
nand U19728 (N_19728,N_13564,N_14737);
or U19729 (N_19729,N_12855,N_14433);
and U19730 (N_19730,N_15590,N_14917);
and U19731 (N_19731,N_13988,N_13971);
and U19732 (N_19732,N_15582,N_13938);
nor U19733 (N_19733,N_12811,N_12153);
and U19734 (N_19734,N_12404,N_13178);
xor U19735 (N_19735,N_13449,N_14835);
and U19736 (N_19736,N_13714,N_13198);
nand U19737 (N_19737,N_15591,N_14231);
nor U19738 (N_19738,N_13986,N_13910);
xor U19739 (N_19739,N_13225,N_12750);
nor U19740 (N_19740,N_13576,N_12181);
or U19741 (N_19741,N_13612,N_13752);
or U19742 (N_19742,N_14576,N_14174);
nand U19743 (N_19743,N_15462,N_15552);
and U19744 (N_19744,N_12964,N_12064);
and U19745 (N_19745,N_14006,N_13509);
xnor U19746 (N_19746,N_14777,N_12560);
nand U19747 (N_19747,N_14452,N_12788);
nor U19748 (N_19748,N_14710,N_14103);
or U19749 (N_19749,N_13597,N_15150);
xnor U19750 (N_19750,N_13272,N_15557);
or U19751 (N_19751,N_13907,N_15247);
nand U19752 (N_19752,N_13410,N_14476);
or U19753 (N_19753,N_12626,N_15318);
xnor U19754 (N_19754,N_15139,N_15693);
and U19755 (N_19755,N_14402,N_12133);
nor U19756 (N_19756,N_13641,N_15279);
nand U19757 (N_19757,N_14952,N_15780);
xnor U19758 (N_19758,N_12325,N_13889);
and U19759 (N_19759,N_12718,N_15696);
nand U19760 (N_19760,N_14040,N_15865);
or U19761 (N_19761,N_12281,N_12735);
or U19762 (N_19762,N_12115,N_12609);
and U19763 (N_19763,N_15848,N_14346);
xor U19764 (N_19764,N_14867,N_12212);
and U19765 (N_19765,N_14767,N_12708);
or U19766 (N_19766,N_14513,N_15439);
xor U19767 (N_19767,N_12375,N_14904);
nand U19768 (N_19768,N_12270,N_13403);
nand U19769 (N_19769,N_14383,N_12083);
nand U19770 (N_19770,N_15931,N_15954);
nor U19771 (N_19771,N_12866,N_15309);
nor U19772 (N_19772,N_13276,N_12492);
nor U19773 (N_19773,N_15675,N_14419);
and U19774 (N_19774,N_12762,N_14899);
and U19775 (N_19775,N_15261,N_13463);
and U19776 (N_19776,N_15272,N_15244);
or U19777 (N_19777,N_15915,N_14115);
nor U19778 (N_19778,N_15572,N_15143);
nand U19779 (N_19779,N_12671,N_14903);
nor U19780 (N_19780,N_13085,N_14316);
or U19781 (N_19781,N_12196,N_14653);
nor U19782 (N_19782,N_12913,N_14664);
or U19783 (N_19783,N_15062,N_15674);
nor U19784 (N_19784,N_15202,N_13567);
xor U19785 (N_19785,N_13741,N_12411);
and U19786 (N_19786,N_15060,N_14314);
xor U19787 (N_19787,N_15636,N_14899);
xor U19788 (N_19788,N_13292,N_12401);
nor U19789 (N_19789,N_13546,N_12497);
or U19790 (N_19790,N_12747,N_12094);
xnor U19791 (N_19791,N_15125,N_13588);
xor U19792 (N_19792,N_13010,N_15497);
nand U19793 (N_19793,N_15094,N_14889);
and U19794 (N_19794,N_15880,N_12570);
and U19795 (N_19795,N_12079,N_13340);
nand U19796 (N_19796,N_12794,N_14858);
or U19797 (N_19797,N_12399,N_12921);
xnor U19798 (N_19798,N_12794,N_14302);
and U19799 (N_19799,N_14751,N_14526);
nand U19800 (N_19800,N_12998,N_13345);
and U19801 (N_19801,N_13358,N_14563);
or U19802 (N_19802,N_15070,N_15606);
or U19803 (N_19803,N_15268,N_14553);
and U19804 (N_19804,N_15324,N_12818);
or U19805 (N_19805,N_12925,N_12269);
nor U19806 (N_19806,N_12543,N_12863);
xor U19807 (N_19807,N_14738,N_14473);
nor U19808 (N_19808,N_12030,N_15630);
nor U19809 (N_19809,N_13684,N_12846);
xnor U19810 (N_19810,N_13897,N_13620);
and U19811 (N_19811,N_12525,N_15655);
xor U19812 (N_19812,N_14740,N_13286);
nand U19813 (N_19813,N_12538,N_14777);
nand U19814 (N_19814,N_12344,N_15520);
nor U19815 (N_19815,N_13590,N_13612);
nor U19816 (N_19816,N_15387,N_15240);
nand U19817 (N_19817,N_15680,N_14234);
xnor U19818 (N_19818,N_15372,N_12478);
and U19819 (N_19819,N_15354,N_12134);
nand U19820 (N_19820,N_14512,N_12412);
or U19821 (N_19821,N_14100,N_13518);
nand U19822 (N_19822,N_14502,N_14419);
nor U19823 (N_19823,N_13622,N_14126);
and U19824 (N_19824,N_15250,N_12428);
or U19825 (N_19825,N_15252,N_13517);
nor U19826 (N_19826,N_14777,N_13244);
xnor U19827 (N_19827,N_14598,N_13390);
and U19828 (N_19828,N_13718,N_12860);
nand U19829 (N_19829,N_12157,N_13507);
nor U19830 (N_19830,N_12717,N_14656);
nor U19831 (N_19831,N_12800,N_13263);
or U19832 (N_19832,N_13989,N_12477);
nand U19833 (N_19833,N_15905,N_15431);
nand U19834 (N_19834,N_14606,N_13489);
or U19835 (N_19835,N_14971,N_15979);
xor U19836 (N_19836,N_12663,N_14835);
nor U19837 (N_19837,N_12884,N_15129);
nand U19838 (N_19838,N_12167,N_13784);
or U19839 (N_19839,N_13723,N_13707);
nor U19840 (N_19840,N_14729,N_12127);
nor U19841 (N_19841,N_12709,N_13556);
or U19842 (N_19842,N_12368,N_12502);
nand U19843 (N_19843,N_15747,N_14036);
nor U19844 (N_19844,N_14876,N_14562);
nor U19845 (N_19845,N_14929,N_15043);
and U19846 (N_19846,N_12165,N_15966);
nor U19847 (N_19847,N_13620,N_14867);
nand U19848 (N_19848,N_12805,N_15417);
nand U19849 (N_19849,N_14613,N_12523);
nor U19850 (N_19850,N_13801,N_13934);
xor U19851 (N_19851,N_13866,N_13541);
or U19852 (N_19852,N_14080,N_13540);
nor U19853 (N_19853,N_12718,N_13934);
nand U19854 (N_19854,N_13517,N_14523);
and U19855 (N_19855,N_12630,N_14580);
nor U19856 (N_19856,N_15486,N_14949);
nand U19857 (N_19857,N_12861,N_14867);
nand U19858 (N_19858,N_13902,N_13867);
and U19859 (N_19859,N_12277,N_12081);
and U19860 (N_19860,N_14183,N_13922);
nor U19861 (N_19861,N_14642,N_15127);
and U19862 (N_19862,N_14160,N_15451);
and U19863 (N_19863,N_14771,N_14740);
nand U19864 (N_19864,N_15643,N_15258);
nand U19865 (N_19865,N_13151,N_15946);
and U19866 (N_19866,N_13836,N_12630);
and U19867 (N_19867,N_15751,N_13359);
nand U19868 (N_19868,N_15323,N_14135);
and U19869 (N_19869,N_12338,N_15274);
and U19870 (N_19870,N_15264,N_12934);
nor U19871 (N_19871,N_13257,N_12185);
nor U19872 (N_19872,N_15008,N_12981);
or U19873 (N_19873,N_15300,N_13211);
and U19874 (N_19874,N_12540,N_12440);
and U19875 (N_19875,N_15984,N_14887);
nand U19876 (N_19876,N_15283,N_15079);
or U19877 (N_19877,N_13131,N_13107);
nand U19878 (N_19878,N_14615,N_15095);
or U19879 (N_19879,N_13056,N_15353);
nand U19880 (N_19880,N_15608,N_13017);
and U19881 (N_19881,N_15359,N_15188);
nand U19882 (N_19882,N_13543,N_12039);
or U19883 (N_19883,N_14326,N_15384);
nand U19884 (N_19884,N_14730,N_14340);
nor U19885 (N_19885,N_15449,N_13833);
and U19886 (N_19886,N_13032,N_15488);
xor U19887 (N_19887,N_14454,N_15810);
or U19888 (N_19888,N_15244,N_12409);
nand U19889 (N_19889,N_14041,N_14854);
nor U19890 (N_19890,N_14966,N_14081);
xnor U19891 (N_19891,N_13920,N_14652);
nand U19892 (N_19892,N_15951,N_13135);
nor U19893 (N_19893,N_12134,N_12480);
nor U19894 (N_19894,N_14456,N_14972);
nand U19895 (N_19895,N_12546,N_13789);
nor U19896 (N_19896,N_12071,N_12535);
nor U19897 (N_19897,N_12011,N_12887);
xnor U19898 (N_19898,N_12277,N_12323);
and U19899 (N_19899,N_15511,N_12086);
xor U19900 (N_19900,N_15323,N_12345);
and U19901 (N_19901,N_14842,N_12819);
and U19902 (N_19902,N_14756,N_12696);
nand U19903 (N_19903,N_13617,N_12399);
or U19904 (N_19904,N_14682,N_15635);
and U19905 (N_19905,N_12095,N_13275);
nand U19906 (N_19906,N_14072,N_14911);
nor U19907 (N_19907,N_15381,N_15979);
nor U19908 (N_19908,N_13509,N_12908);
and U19909 (N_19909,N_13128,N_15841);
and U19910 (N_19910,N_14531,N_14511);
nor U19911 (N_19911,N_12541,N_12088);
or U19912 (N_19912,N_15800,N_13725);
nand U19913 (N_19913,N_15633,N_13237);
nand U19914 (N_19914,N_14724,N_13292);
nand U19915 (N_19915,N_13066,N_12914);
nor U19916 (N_19916,N_12417,N_13958);
nand U19917 (N_19917,N_13252,N_14694);
or U19918 (N_19918,N_14774,N_14571);
or U19919 (N_19919,N_14396,N_13491);
nor U19920 (N_19920,N_14252,N_15922);
xor U19921 (N_19921,N_13227,N_13615);
nor U19922 (N_19922,N_12396,N_12200);
and U19923 (N_19923,N_13672,N_15449);
xnor U19924 (N_19924,N_15736,N_14652);
nand U19925 (N_19925,N_13664,N_13314);
xor U19926 (N_19926,N_14048,N_14943);
or U19927 (N_19927,N_15346,N_15879);
nand U19928 (N_19928,N_13575,N_14892);
and U19929 (N_19929,N_15303,N_15049);
xor U19930 (N_19930,N_12491,N_14027);
xnor U19931 (N_19931,N_13520,N_13841);
nor U19932 (N_19932,N_14021,N_12037);
and U19933 (N_19933,N_15720,N_15229);
nor U19934 (N_19934,N_14654,N_13755);
or U19935 (N_19935,N_15899,N_15243);
or U19936 (N_19936,N_15692,N_15898);
xor U19937 (N_19937,N_14897,N_13486);
or U19938 (N_19938,N_13610,N_12156);
or U19939 (N_19939,N_14516,N_12553);
nor U19940 (N_19940,N_14912,N_15074);
or U19941 (N_19941,N_12541,N_15747);
nand U19942 (N_19942,N_14993,N_15574);
or U19943 (N_19943,N_14586,N_13340);
nor U19944 (N_19944,N_15479,N_14509);
and U19945 (N_19945,N_14152,N_14328);
nand U19946 (N_19946,N_14296,N_12205);
nand U19947 (N_19947,N_15655,N_12954);
xor U19948 (N_19948,N_13514,N_12615);
and U19949 (N_19949,N_13240,N_14181);
xnor U19950 (N_19950,N_15051,N_14859);
nor U19951 (N_19951,N_14700,N_15768);
xor U19952 (N_19952,N_13809,N_13441);
or U19953 (N_19953,N_14054,N_12119);
and U19954 (N_19954,N_12636,N_13476);
or U19955 (N_19955,N_14951,N_13185);
nor U19956 (N_19956,N_15043,N_14175);
and U19957 (N_19957,N_12268,N_13040);
xnor U19958 (N_19958,N_14857,N_15865);
nand U19959 (N_19959,N_12498,N_12280);
and U19960 (N_19960,N_12769,N_13216);
or U19961 (N_19961,N_15303,N_15557);
or U19962 (N_19962,N_14015,N_12752);
and U19963 (N_19963,N_12811,N_13355);
xnor U19964 (N_19964,N_15488,N_12194);
and U19965 (N_19965,N_15133,N_15699);
nand U19966 (N_19966,N_14440,N_15434);
or U19967 (N_19967,N_14133,N_13163);
nand U19968 (N_19968,N_13778,N_15364);
nand U19969 (N_19969,N_15563,N_13814);
nor U19970 (N_19970,N_14229,N_13539);
nand U19971 (N_19971,N_15645,N_14584);
and U19972 (N_19972,N_13570,N_12594);
or U19973 (N_19973,N_13387,N_13918);
or U19974 (N_19974,N_14526,N_12614);
nand U19975 (N_19975,N_13591,N_13133);
and U19976 (N_19976,N_13894,N_13981);
nor U19977 (N_19977,N_12959,N_13801);
or U19978 (N_19978,N_13433,N_13230);
nor U19979 (N_19979,N_13913,N_15453);
nand U19980 (N_19980,N_13667,N_12504);
nand U19981 (N_19981,N_15049,N_13297);
nand U19982 (N_19982,N_12428,N_13238);
nand U19983 (N_19983,N_13688,N_12119);
nand U19984 (N_19984,N_12697,N_15063);
and U19985 (N_19985,N_14320,N_13317);
nor U19986 (N_19986,N_13844,N_14741);
or U19987 (N_19987,N_13482,N_12274);
nand U19988 (N_19988,N_15017,N_12735);
nand U19989 (N_19989,N_12365,N_13595);
and U19990 (N_19990,N_13895,N_15567);
or U19991 (N_19991,N_15961,N_12581);
or U19992 (N_19992,N_12796,N_15284);
and U19993 (N_19993,N_15732,N_14978);
nor U19994 (N_19994,N_13727,N_14703);
nand U19995 (N_19995,N_15204,N_15462);
nor U19996 (N_19996,N_15221,N_14245);
nor U19997 (N_19997,N_14858,N_14035);
or U19998 (N_19998,N_15168,N_12104);
and U19999 (N_19999,N_12164,N_12259);
or UO_0 (O_0,N_19712,N_18116);
and UO_1 (O_1,N_17535,N_17895);
and UO_2 (O_2,N_16202,N_16286);
and UO_3 (O_3,N_17705,N_18405);
or UO_4 (O_4,N_16462,N_17515);
or UO_5 (O_5,N_16718,N_18721);
nor UO_6 (O_6,N_16349,N_17943);
xor UO_7 (O_7,N_17749,N_18449);
nand UO_8 (O_8,N_19993,N_17393);
nor UO_9 (O_9,N_16482,N_19222);
or UO_10 (O_10,N_17485,N_16691);
nand UO_11 (O_11,N_19081,N_18626);
or UO_12 (O_12,N_17824,N_16635);
nor UO_13 (O_13,N_18538,N_16016);
nor UO_14 (O_14,N_19412,N_19158);
and UO_15 (O_15,N_16786,N_18041);
or UO_16 (O_16,N_16353,N_16325);
or UO_17 (O_17,N_19469,N_17622);
or UO_18 (O_18,N_18432,N_18563);
nor UO_19 (O_19,N_18586,N_16201);
and UO_20 (O_20,N_16378,N_17383);
nand UO_21 (O_21,N_19762,N_17037);
and UO_22 (O_22,N_19023,N_19849);
or UO_23 (O_23,N_16308,N_17302);
nor UO_24 (O_24,N_18680,N_18751);
nor UO_25 (O_25,N_17073,N_16847);
nor UO_26 (O_26,N_16200,N_18720);
nand UO_27 (O_27,N_18959,N_17980);
nor UO_28 (O_28,N_18649,N_16788);
xor UO_29 (O_29,N_19384,N_18302);
xnor UO_30 (O_30,N_19866,N_16487);
nor UO_31 (O_31,N_17333,N_17153);
xnor UO_32 (O_32,N_16185,N_18105);
and UO_33 (O_33,N_16221,N_17735);
or UO_34 (O_34,N_17084,N_16442);
and UO_35 (O_35,N_16828,N_18241);
nand UO_36 (O_36,N_16524,N_17412);
and UO_37 (O_37,N_17507,N_18977);
nand UO_38 (O_38,N_18776,N_16696);
and UO_39 (O_39,N_16947,N_18320);
nor UO_40 (O_40,N_17774,N_16671);
or UO_41 (O_41,N_19183,N_17669);
or UO_42 (O_42,N_19970,N_17240);
nand UO_43 (O_43,N_18203,N_17626);
nand UO_44 (O_44,N_17413,N_19487);
nand UO_45 (O_45,N_18306,N_19287);
or UO_46 (O_46,N_16994,N_17827);
xor UO_47 (O_47,N_17139,N_19278);
and UO_48 (O_48,N_17221,N_17104);
xor UO_49 (O_49,N_18814,N_16931);
and UO_50 (O_50,N_18469,N_17094);
and UO_51 (O_51,N_19978,N_16575);
nand UO_52 (O_52,N_18522,N_16273);
nor UO_53 (O_53,N_17658,N_19696);
nor UO_54 (O_54,N_19284,N_17055);
or UO_55 (O_55,N_16305,N_16035);
nor UO_56 (O_56,N_18610,N_16337);
or UO_57 (O_57,N_19215,N_17367);
nand UO_58 (O_58,N_19262,N_17384);
or UO_59 (O_59,N_19524,N_17899);
and UO_60 (O_60,N_19920,N_18612);
nand UO_61 (O_61,N_17711,N_16050);
nand UO_62 (O_62,N_16204,N_18699);
nor UO_63 (O_63,N_16107,N_19156);
nor UO_64 (O_64,N_19893,N_19693);
nor UO_65 (O_65,N_18953,N_19488);
or UO_66 (O_66,N_18892,N_18485);
or UO_67 (O_67,N_18236,N_17461);
nand UO_68 (O_68,N_16448,N_18781);
nor UO_69 (O_69,N_19100,N_19432);
nand UO_70 (O_70,N_17432,N_18848);
nor UO_71 (O_71,N_16407,N_18755);
nor UO_72 (O_72,N_16972,N_18537);
nand UO_73 (O_73,N_19144,N_18006);
or UO_74 (O_74,N_17045,N_16344);
nand UO_75 (O_75,N_19324,N_18792);
nor UO_76 (O_76,N_19787,N_17152);
and UO_77 (O_77,N_16490,N_17307);
and UO_78 (O_78,N_16164,N_17066);
nand UO_79 (O_79,N_19083,N_18211);
nor UO_80 (O_80,N_16052,N_19502);
and UO_81 (O_81,N_19011,N_18961);
and UO_82 (O_82,N_18322,N_17419);
and UO_83 (O_83,N_17575,N_17835);
or UO_84 (O_84,N_19881,N_16705);
and UO_85 (O_85,N_19180,N_18616);
xnor UO_86 (O_86,N_19937,N_19179);
or UO_87 (O_87,N_18825,N_17613);
and UO_88 (O_88,N_19120,N_16198);
nor UO_89 (O_89,N_17662,N_19140);
nand UO_90 (O_90,N_16795,N_18341);
nand UO_91 (O_91,N_17378,N_18713);
nor UO_92 (O_92,N_19961,N_19602);
nor UO_93 (O_93,N_16034,N_18507);
or UO_94 (O_94,N_17633,N_16592);
nand UO_95 (O_95,N_19211,N_17530);
or UO_96 (O_96,N_17491,N_19754);
nand UO_97 (O_97,N_18017,N_18905);
nor UO_98 (O_98,N_16215,N_16626);
and UO_99 (O_99,N_17523,N_17617);
nand UO_100 (O_100,N_19705,N_17060);
nor UO_101 (O_101,N_17075,N_17916);
or UO_102 (O_102,N_19472,N_18960);
or UO_103 (O_103,N_19767,N_19938);
nand UO_104 (O_104,N_17505,N_18127);
or UO_105 (O_105,N_16382,N_19649);
or UO_106 (O_106,N_18256,N_18108);
nor UO_107 (O_107,N_17609,N_19036);
nand UO_108 (O_108,N_17100,N_19005);
nand UO_109 (O_109,N_19723,N_16372);
nand UO_110 (O_110,N_16561,N_19288);
nand UO_111 (O_111,N_16359,N_18172);
and UO_112 (O_112,N_17193,N_17851);
xnor UO_113 (O_113,N_19348,N_18804);
nor UO_114 (O_114,N_18424,N_18873);
xor UO_115 (O_115,N_19667,N_19437);
or UO_116 (O_116,N_17959,N_19119);
xnor UO_117 (O_117,N_16942,N_17165);
xnor UO_118 (O_118,N_17767,N_17479);
and UO_119 (O_119,N_17667,N_18901);
xor UO_120 (O_120,N_17181,N_19743);
and UO_121 (O_121,N_18069,N_16319);
or UO_122 (O_122,N_16083,N_16664);
xnor UO_123 (O_123,N_18859,N_19742);
or UO_124 (O_124,N_18487,N_19124);
xor UO_125 (O_125,N_16429,N_18922);
nor UO_126 (O_126,N_18219,N_18559);
nor UO_127 (O_127,N_17727,N_19740);
nor UO_128 (O_128,N_18893,N_17733);
xor UO_129 (O_129,N_17738,N_16357);
or UO_130 (O_130,N_19720,N_19417);
nor UO_131 (O_131,N_19890,N_17740);
and UO_132 (O_132,N_18524,N_18508);
xnor UO_133 (O_133,N_18654,N_18237);
nand UO_134 (O_134,N_16342,N_16264);
nand UO_135 (O_135,N_19968,N_16982);
nor UO_136 (O_136,N_17166,N_19515);
and UO_137 (O_137,N_16038,N_17162);
or UO_138 (O_138,N_17114,N_17587);
nand UO_139 (O_139,N_17698,N_18160);
nor UO_140 (O_140,N_17846,N_18433);
nor UO_141 (O_141,N_16595,N_19589);
nor UO_142 (O_142,N_16499,N_19208);
nand UO_143 (O_143,N_16347,N_17951);
nand UO_144 (O_144,N_17024,N_18476);
or UO_145 (O_145,N_17143,N_17049);
or UO_146 (O_146,N_19292,N_16167);
nand UO_147 (O_147,N_19805,N_19072);
or UO_148 (O_148,N_17929,N_16617);
nand UO_149 (O_149,N_18448,N_18951);
and UO_150 (O_150,N_16329,N_16436);
nand UO_151 (O_151,N_16842,N_18214);
xnor UO_152 (O_152,N_16126,N_16205);
nand UO_153 (O_153,N_17005,N_19984);
and UO_154 (O_154,N_19695,N_19854);
or UO_155 (O_155,N_16686,N_17945);
or UO_156 (O_156,N_18638,N_19707);
and UO_157 (O_157,N_19570,N_19503);
nor UO_158 (O_158,N_19798,N_16778);
xnor UO_159 (O_159,N_16328,N_16518);
and UO_160 (O_160,N_16489,N_19664);
and UO_161 (O_161,N_16775,N_17919);
nor UO_162 (O_162,N_16973,N_17340);
or UO_163 (O_163,N_17909,N_16491);
nor UO_164 (O_164,N_18503,N_17370);
and UO_165 (O_165,N_19572,N_16365);
or UO_166 (O_166,N_19044,N_18074);
or UO_167 (O_167,N_19370,N_16820);
nand UO_168 (O_168,N_19520,N_19789);
or UO_169 (O_169,N_17216,N_19852);
nand UO_170 (O_170,N_19191,N_17910);
nor UO_171 (O_171,N_16822,N_16764);
and UO_172 (O_172,N_16173,N_17962);
nand UO_173 (O_173,N_16494,N_18714);
or UO_174 (O_174,N_16709,N_19241);
nor UO_175 (O_175,N_19851,N_16024);
and UO_176 (O_176,N_16739,N_17852);
or UO_177 (O_177,N_16109,N_19657);
or UO_178 (O_178,N_19733,N_19212);
or UO_179 (O_179,N_17879,N_18881);
and UO_180 (O_180,N_16249,N_19500);
xnor UO_181 (O_181,N_17288,N_19547);
xor UO_182 (O_182,N_19091,N_16145);
nand UO_183 (O_183,N_16320,N_16356);
and UO_184 (O_184,N_18351,N_19910);
nand UO_185 (O_185,N_16299,N_16488);
or UO_186 (O_186,N_16928,N_17939);
or UO_187 (O_187,N_19346,N_18981);
xor UO_188 (O_188,N_16158,N_18246);
or UO_189 (O_189,N_18934,N_18132);
or UO_190 (O_190,N_16608,N_17512);
nand UO_191 (O_191,N_19041,N_17047);
or UO_192 (O_192,N_18597,N_19795);
nor UO_193 (O_193,N_19297,N_17022);
and UO_194 (O_194,N_16611,N_16551);
nand UO_195 (O_195,N_17361,N_18223);
xor UO_196 (O_196,N_19645,N_18962);
or UO_197 (O_197,N_16999,N_18190);
or UO_198 (O_198,N_17121,N_16332);
nor UO_199 (O_199,N_19224,N_18590);
nor UO_200 (O_200,N_19616,N_19489);
nor UO_201 (O_201,N_17746,N_17376);
nand UO_202 (O_202,N_16986,N_19505);
xor UO_203 (O_203,N_17913,N_17858);
nand UO_204 (O_204,N_16437,N_18533);
xnor UO_205 (O_205,N_16929,N_18001);
nand UO_206 (O_206,N_18300,N_16333);
nand UO_207 (O_207,N_17242,N_16208);
nand UO_208 (O_208,N_18785,N_18312);
nand UO_209 (O_209,N_18845,N_18491);
and UO_210 (O_210,N_16250,N_19397);
and UO_211 (O_211,N_17815,N_16948);
and UO_212 (O_212,N_17516,N_16965);
nor UO_213 (O_213,N_19186,N_17406);
and UO_214 (O_214,N_16995,N_17141);
or UO_215 (O_215,N_18393,N_17580);
nor UO_216 (O_216,N_16717,N_18583);
nor UO_217 (O_217,N_16312,N_16501);
or UO_218 (O_218,N_16259,N_18502);
and UO_219 (O_219,N_17117,N_18196);
and UO_220 (O_220,N_18715,N_16878);
nand UO_221 (O_221,N_18414,N_17392);
nand UO_222 (O_222,N_16427,N_18677);
nor UO_223 (O_223,N_18044,N_19408);
or UO_224 (O_224,N_17606,N_18920);
and UO_225 (O_225,N_19359,N_19187);
nand UO_226 (O_226,N_16559,N_17071);
and UO_227 (O_227,N_19646,N_16841);
and UO_228 (O_228,N_19722,N_19601);
nand UO_229 (O_229,N_19115,N_18411);
nand UO_230 (O_230,N_17217,N_18602);
nor UO_231 (O_231,N_19928,N_19133);
nor UO_232 (O_232,N_17784,N_16096);
nand UO_233 (O_233,N_17093,N_16257);
or UO_234 (O_234,N_16036,N_19266);
nor UO_235 (O_235,N_18059,N_16529);
nand UO_236 (O_236,N_18192,N_16882);
and UO_237 (O_237,N_19612,N_19776);
nand UO_238 (O_238,N_17985,N_16628);
xnor UO_239 (O_239,N_16370,N_17002);
and UO_240 (O_240,N_16891,N_19609);
and UO_241 (O_241,N_18226,N_19847);
or UO_242 (O_242,N_19495,N_19433);
nor UO_243 (O_243,N_17446,N_17509);
and UO_244 (O_244,N_16420,N_18511);
nor UO_245 (O_245,N_19032,N_19989);
nor UO_246 (O_246,N_19353,N_17965);
nor UO_247 (O_247,N_17739,N_16552);
or UO_248 (O_248,N_16458,N_18420);
nand UO_249 (O_249,N_19319,N_17826);
or UO_250 (O_250,N_19167,N_18852);
and UO_251 (O_251,N_19730,N_16178);
or UO_252 (O_252,N_16859,N_17898);
and UO_253 (O_253,N_16459,N_17487);
nand UO_254 (O_254,N_17700,N_19986);
nand UO_255 (O_255,N_16738,N_16974);
nor UO_256 (O_256,N_16057,N_17381);
and UO_257 (O_257,N_16888,N_18161);
and UO_258 (O_258,N_17940,N_16291);
or UO_259 (O_259,N_16441,N_18983);
and UO_260 (O_260,N_16886,N_16470);
nor UO_261 (O_261,N_19242,N_19685);
nor UO_262 (O_262,N_18095,N_16450);
and UO_263 (O_263,N_18000,N_16930);
or UO_264 (O_264,N_17565,N_18745);
and UO_265 (O_265,N_17081,N_18191);
xnor UO_266 (O_266,N_16687,N_16189);
xnor UO_267 (O_267,N_16751,N_16246);
or UO_268 (O_268,N_17668,N_16180);
or UO_269 (O_269,N_16695,N_18767);
or UO_270 (O_270,N_19007,N_18676);
nor UO_271 (O_271,N_18276,N_19234);
nor UO_272 (O_272,N_16182,N_17044);
nand UO_273 (O_273,N_16354,N_19148);
nor UO_274 (O_274,N_17229,N_19010);
and UO_275 (O_275,N_18762,N_16066);
nand UO_276 (O_276,N_18443,N_19871);
and UO_277 (O_277,N_16946,N_19111);
xor UO_278 (O_278,N_16360,N_17619);
nor UO_279 (O_279,N_16379,N_17737);
nand UO_280 (O_280,N_17797,N_17593);
and UO_281 (O_281,N_18376,N_16702);
and UO_282 (O_282,N_18188,N_19629);
or UO_283 (O_283,N_16725,N_17409);
or UO_284 (O_284,N_16019,N_17365);
or UO_285 (O_285,N_17471,N_17431);
or UO_286 (O_286,N_19981,N_17731);
or UO_287 (O_287,N_17486,N_18952);
xor UO_288 (O_288,N_19448,N_17390);
nor UO_289 (O_289,N_18679,N_18628);
and UO_290 (O_290,N_16772,N_18747);
nor UO_291 (O_291,N_18897,N_18769);
nand UO_292 (O_292,N_17110,N_16027);
nand UO_293 (O_293,N_17291,N_16440);
or UO_294 (O_294,N_16316,N_19037);
nand UO_295 (O_295,N_18247,N_18771);
and UO_296 (O_296,N_17138,N_17878);
and UO_297 (O_297,N_19216,N_19603);
nand UO_298 (O_298,N_18644,N_17837);
or UO_299 (O_299,N_19425,N_19845);
and UO_300 (O_300,N_18130,N_17896);
and UO_301 (O_301,N_16884,N_18282);
or UO_302 (O_302,N_19253,N_18674);
nor UO_303 (O_303,N_16517,N_18637);
xor UO_304 (O_304,N_16514,N_16322);
nand UO_305 (O_305,N_19352,N_16817);
or UO_306 (O_306,N_19046,N_19074);
nand UO_307 (O_307,N_16646,N_16823);
or UO_308 (O_308,N_19966,N_17567);
or UO_309 (O_309,N_18774,N_17219);
nor UO_310 (O_310,N_18890,N_19940);
nor UO_311 (O_311,N_16300,N_17258);
xnor UO_312 (O_312,N_17761,N_18931);
and UO_313 (O_313,N_16438,N_19135);
and UO_314 (O_314,N_17556,N_16402);
nor UO_315 (O_315,N_19302,N_19314);
nor UO_316 (O_316,N_19271,N_18576);
nand UO_317 (O_317,N_18947,N_16054);
nor UO_318 (O_318,N_18513,N_16502);
nor UO_319 (O_319,N_19518,N_16421);
nor UO_320 (O_320,N_19658,N_18259);
and UO_321 (O_321,N_18182,N_16274);
nand UO_322 (O_322,N_17867,N_18023);
nand UO_323 (O_323,N_18800,N_16439);
and UO_324 (O_324,N_19451,N_19022);
and UO_325 (O_325,N_16449,N_19899);
nor UO_326 (O_326,N_16051,N_16576);
and UO_327 (O_327,N_18332,N_18627);
nand UO_328 (O_328,N_19643,N_16265);
nand UO_329 (O_329,N_18055,N_16025);
or UO_330 (O_330,N_18565,N_19939);
nor UO_331 (O_331,N_16335,N_19277);
or UO_332 (O_332,N_17877,N_18170);
nand UO_333 (O_333,N_16682,N_17988);
nand UO_334 (O_334,N_19865,N_19574);
and UO_335 (O_335,N_17177,N_18561);
or UO_336 (O_336,N_17801,N_16782);
xnor UO_337 (O_337,N_17467,N_17142);
xor UO_338 (O_338,N_19249,N_16883);
or UO_339 (O_339,N_16234,N_18415);
nor UO_340 (O_340,N_18743,N_17574);
or UO_341 (O_341,N_17666,N_19107);
or UO_342 (O_342,N_17953,N_18969);
nor UO_343 (O_343,N_19625,N_17414);
and UO_344 (O_344,N_19808,N_19872);
nor UO_345 (O_345,N_18400,N_18594);
or UO_346 (O_346,N_18435,N_16610);
or UO_347 (O_347,N_18361,N_17079);
or UO_348 (O_348,N_17007,N_18461);
nand UO_349 (O_349,N_17764,N_18648);
xnor UO_350 (O_350,N_16901,N_16028);
xnor UO_351 (O_351,N_19699,N_18615);
nand UO_352 (O_352,N_17663,N_17129);
nand UO_353 (O_353,N_16479,N_16138);
and UO_354 (O_354,N_17758,N_19141);
or UO_355 (O_355,N_16485,N_16471);
or UO_356 (O_356,N_17279,N_19057);
nand UO_357 (O_357,N_19824,N_19713);
nor UO_358 (O_358,N_17744,N_19626);
xnor UO_359 (O_359,N_18145,N_19479);
nor UO_360 (O_360,N_17434,N_18821);
or UO_361 (O_361,N_18801,N_16845);
nand UO_362 (O_362,N_19496,N_19145);
nor UO_363 (O_363,N_19517,N_17199);
nand UO_364 (O_364,N_16769,N_17402);
nand UO_365 (O_365,N_16937,N_17277);
nor UO_366 (O_366,N_19098,N_18984);
nand UO_367 (O_367,N_18996,N_19185);
and UO_368 (O_368,N_18497,N_19221);
and UO_369 (O_369,N_17424,N_19876);
nand UO_370 (O_370,N_18484,N_17148);
xnor UO_371 (O_371,N_19741,N_18081);
or UO_372 (O_372,N_17892,N_18046);
and UO_373 (O_373,N_18352,N_16454);
nand UO_374 (O_374,N_17092,N_17912);
nor UO_375 (O_375,N_19554,N_18163);
nand UO_376 (O_376,N_18248,N_17548);
or UO_377 (O_377,N_16396,N_18661);
nor UO_378 (O_378,N_16615,N_19861);
nand UO_379 (O_379,N_16645,N_19672);
and UO_380 (O_380,N_17544,N_19510);
nor UO_381 (O_381,N_18668,N_18782);
and UO_382 (O_382,N_19552,N_17429);
nand UO_383 (O_383,N_16818,N_19560);
nor UO_384 (O_384,N_18707,N_16248);
nor UO_385 (O_385,N_18562,N_19407);
and UO_386 (O_386,N_16129,N_16311);
and UO_387 (O_387,N_16416,N_18718);
nand UO_388 (O_388,N_17861,N_17379);
nor UO_389 (O_389,N_16880,N_18991);
nand UO_390 (O_390,N_18275,N_17589);
and UO_391 (O_391,N_16679,N_16814);
xor UO_392 (O_392,N_19809,N_17303);
or UO_393 (O_393,N_16476,N_19586);
nor UO_394 (O_394,N_17154,N_16266);
nand UO_395 (O_395,N_18141,N_16860);
nand UO_396 (O_396,N_19209,N_17451);
or UO_397 (O_397,N_17335,N_19239);
or UO_398 (O_398,N_16724,N_18967);
nand UO_399 (O_399,N_17396,N_19551);
and UO_400 (O_400,N_19474,N_19739);
nor UO_401 (O_401,N_18311,N_19295);
and UO_402 (O_402,N_19024,N_16582);
nor UO_403 (O_403,N_19411,N_16916);
nor UO_404 (O_404,N_17888,N_16924);
nor UO_405 (O_405,N_19677,N_16546);
xor UO_406 (O_406,N_16506,N_17660);
or UO_407 (O_407,N_16081,N_18082);
nand UO_408 (O_408,N_17082,N_16708);
nand UO_409 (O_409,N_18641,N_18742);
nand UO_410 (O_410,N_18906,N_19285);
nor UO_411 (O_411,N_17292,N_17052);
nor UO_412 (O_412,N_18406,N_16543);
nor UO_413 (O_413,N_19656,N_18383);
nand UO_414 (O_414,N_19323,N_18837);
nand UO_415 (O_415,N_18752,N_18222);
nor UO_416 (O_416,N_19903,N_17720);
or UO_417 (O_417,N_19527,N_16681);
and UO_418 (O_418,N_17294,N_17834);
and UO_419 (O_419,N_17811,N_16445);
or UO_420 (O_420,N_18392,N_16780);
nand UO_421 (O_421,N_16009,N_19429);
nor UO_422 (O_422,N_19283,N_18595);
xor UO_423 (O_423,N_18536,N_19594);
nand UO_424 (O_424,N_18086,N_16759);
and UO_425 (O_425,N_16560,N_16136);
nand UO_426 (O_426,N_19567,N_17651);
nand UO_427 (O_427,N_17533,N_17604);
nor UO_428 (O_428,N_16956,N_19084);
and UO_429 (O_429,N_16836,N_18992);
or UO_430 (O_430,N_19190,N_16275);
nand UO_431 (O_431,N_17194,N_19790);
and UO_432 (O_432,N_19329,N_18280);
and UO_433 (O_433,N_16125,N_17135);
nor UO_434 (O_434,N_16252,N_16134);
or UO_435 (O_435,N_19675,N_19485);
nand UO_436 (O_436,N_19347,N_17699);
and UO_437 (O_437,N_17195,N_19843);
and UO_438 (O_438,N_17197,N_16157);
nand UO_439 (O_439,N_17284,N_18685);
or UO_440 (O_440,N_18314,N_17914);
nor UO_441 (O_441,N_16032,N_17665);
nor UO_442 (O_442,N_19233,N_17492);
or UO_443 (O_443,N_18467,N_16675);
nand UO_444 (O_444,N_19836,N_18370);
or UO_445 (O_445,N_17348,N_18474);
nor UO_446 (O_446,N_18805,N_19152);
and UO_447 (O_447,N_17000,N_18272);
nor UO_448 (O_448,N_19877,N_19834);
nor UO_449 (O_449,N_18657,N_17691);
xor UO_450 (O_450,N_18466,N_16075);
nor UO_451 (O_451,N_17400,N_17713);
or UO_452 (O_452,N_17853,N_16169);
or UO_453 (O_453,N_19138,N_19727);
nor UO_454 (O_454,N_19704,N_18639);
nor UO_455 (O_455,N_17180,N_16371);
or UO_456 (O_456,N_16390,N_18812);
xor UO_457 (O_457,N_19470,N_16699);
nor UO_458 (O_458,N_18052,N_19653);
nand UO_459 (O_459,N_17831,N_18647);
nand UO_460 (O_460,N_16810,N_19692);
nand UO_461 (O_461,N_18740,N_17098);
and UO_462 (O_462,N_19134,N_19207);
nand UO_463 (O_463,N_19611,N_18486);
or UO_464 (O_464,N_18770,N_18764);
nor UO_465 (O_465,N_18501,N_18238);
nor UO_466 (O_466,N_17207,N_17090);
and UO_467 (O_467,N_16230,N_17457);
nor UO_468 (O_468,N_17190,N_18345);
xnor UO_469 (O_469,N_19306,N_19565);
or UO_470 (O_470,N_17564,N_16062);
xnor UO_471 (O_471,N_18340,N_19194);
or UO_472 (O_472,N_17987,N_16103);
nand UO_473 (O_473,N_16563,N_19436);
and UO_474 (O_474,N_19172,N_17272);
and UO_475 (O_475,N_18463,N_17124);
and UO_476 (O_476,N_17977,N_19325);
nor UO_477 (O_477,N_19842,N_18941);
xor UO_478 (O_478,N_19462,N_18360);
or UO_479 (O_479,N_18450,N_19584);
xor UO_480 (O_480,N_19568,N_18481);
xor UO_481 (O_481,N_17173,N_18019);
and UO_482 (O_482,N_17301,N_19912);
or UO_483 (O_483,N_18839,N_19456);
and UO_484 (O_484,N_18877,N_19673);
nand UO_485 (O_485,N_16355,N_19259);
nand UO_486 (O_486,N_17653,N_18206);
or UO_487 (O_487,N_17146,N_18077);
and UO_488 (O_488,N_18784,N_17783);
nor UO_489 (O_489,N_17941,N_19682);
or UO_490 (O_490,N_18636,N_17032);
or UO_491 (O_491,N_19227,N_19576);
and UO_492 (O_492,N_17541,N_17261);
and UO_493 (O_493,N_19240,N_17765);
or UO_494 (O_494,N_18540,N_16621);
nor UO_495 (O_495,N_17779,N_17127);
or UO_496 (O_496,N_19827,N_19291);
or UO_497 (O_497,N_16294,N_17246);
or UO_498 (O_498,N_17862,N_16412);
nand UO_499 (O_499,N_19763,N_16911);
nand UO_500 (O_500,N_19773,N_16241);
or UO_501 (O_501,N_18696,N_17820);
or UO_502 (O_502,N_18047,N_16642);
and UO_503 (O_503,N_18035,N_18840);
nor UO_504 (O_504,N_16376,N_16978);
nand UO_505 (O_505,N_16415,N_16540);
and UO_506 (O_506,N_19832,N_16128);
or UO_507 (O_507,N_16877,N_19823);
and UO_508 (O_508,N_18719,N_19651);
and UO_509 (O_509,N_16826,N_16478);
or UO_510 (O_510,N_17116,N_18724);
xnor UO_511 (O_511,N_19361,N_16622);
xor UO_512 (O_512,N_19894,N_19086);
nor UO_513 (O_513,N_16115,N_17891);
nand UO_514 (O_514,N_19588,N_17027);
and UO_515 (O_515,N_18043,N_17125);
nor UO_516 (O_516,N_17841,N_16007);
or UO_517 (O_517,N_19587,N_17796);
and UO_518 (O_518,N_16116,N_18976);
or UO_519 (O_519,N_16525,N_17174);
and UO_520 (O_520,N_17313,N_18966);
and UO_521 (O_521,N_16614,N_17785);
and UO_522 (O_522,N_18338,N_17042);
nand UO_523 (O_523,N_17747,N_16897);
nand UO_524 (O_524,N_19963,N_18235);
and UO_525 (O_525,N_17577,N_17675);
nand UO_526 (O_526,N_16481,N_19058);
nor UO_527 (O_527,N_17183,N_17592);
nor UO_528 (O_528,N_18554,N_19440);
or UO_529 (O_529,N_16447,N_17102);
or UO_530 (O_530,N_17426,N_16846);
nor UO_531 (O_531,N_19294,N_16612);
nand UO_532 (O_532,N_17113,N_16701);
nor UO_533 (O_533,N_16925,N_16292);
or UO_534 (O_534,N_17865,N_16692);
xnor UO_535 (O_535,N_18150,N_18927);
nor UO_536 (O_536,N_18887,N_19630);
nand UO_537 (O_537,N_18874,N_16594);
nor UO_538 (O_538,N_17268,N_18847);
or UO_539 (O_539,N_17976,N_17478);
and UO_540 (O_540,N_18032,N_18321);
nor UO_541 (O_541,N_16072,N_18545);
and UO_542 (O_542,N_19009,N_19930);
nand UO_543 (O_543,N_19315,N_18293);
nand UO_544 (O_544,N_18571,N_18057);
nor UO_545 (O_545,N_19096,N_17836);
or UO_546 (O_546,N_18104,N_18475);
and UO_547 (O_547,N_18207,N_16314);
or UO_548 (O_548,N_17029,N_17549);
and UO_549 (O_549,N_18122,N_19373);
nor UO_550 (O_550,N_16315,N_18935);
nand UO_551 (O_551,N_16636,N_18357);
and UO_552 (O_552,N_16118,N_18273);
nor UO_553 (O_553,N_17009,N_19883);
nor UO_554 (O_554,N_19755,N_16222);
and UO_555 (O_555,N_18665,N_16766);
or UO_556 (O_556,N_18264,N_17115);
or UO_557 (O_557,N_17799,N_16338);
nor UO_558 (O_558,N_16669,N_19117);
nor UO_559 (O_559,N_16711,N_19724);
or UO_560 (O_560,N_17692,N_18441);
nand UO_561 (O_561,N_18896,N_17339);
and UO_562 (O_562,N_19927,N_18317);
or UO_563 (O_563,N_16907,N_16730);
nor UO_564 (O_564,N_19494,N_18727);
nor UO_565 (O_565,N_19702,N_19243);
xnor UO_566 (O_566,N_16497,N_16176);
or UO_567 (O_567,N_19464,N_19817);
or UO_568 (O_568,N_16987,N_19105);
nor UO_569 (O_569,N_16528,N_17062);
xnor UO_570 (O_570,N_16511,N_17828);
and UO_571 (O_571,N_16923,N_17465);
nor UO_572 (O_572,N_19250,N_19480);
or UO_573 (O_573,N_18144,N_17464);
nand UO_574 (O_574,N_17149,N_17198);
or UO_575 (O_575,N_17998,N_16604);
nor UO_576 (O_576,N_18539,N_18579);
or UO_577 (O_577,N_19228,N_17063);
nand UO_578 (O_578,N_19200,N_16397);
xnor UO_579 (O_579,N_16092,N_16288);
nor UO_580 (O_580,N_18787,N_19623);
and UO_581 (O_581,N_18642,N_18629);
or UO_582 (O_582,N_17300,N_18518);
nor UO_583 (O_583,N_16743,N_19504);
or UO_584 (O_584,N_19441,N_19729);
nand UO_585 (O_585,N_17961,N_18999);
and UO_586 (O_586,N_16271,N_18523);
nor UO_587 (O_587,N_17703,N_16253);
and UO_588 (O_588,N_18166,N_17059);
nand UO_589 (O_589,N_19582,N_19175);
and UO_590 (O_590,N_18058,N_16808);
or UO_591 (O_591,N_19457,N_17839);
xor UO_592 (O_592,N_17050,N_16532);
and UO_593 (O_593,N_18613,N_19631);
or UO_594 (O_594,N_19443,N_19015);
or UO_595 (O_595,N_17819,N_17097);
or UO_596 (O_596,N_18667,N_17926);
nand UO_597 (O_597,N_19758,N_17028);
nor UO_598 (O_598,N_16309,N_16553);
nor UO_599 (O_599,N_17437,N_16833);
xor UO_600 (O_600,N_16465,N_17894);
or UO_601 (O_601,N_19593,N_16678);
nand UO_602 (O_602,N_17130,N_16295);
and UO_603 (O_603,N_16154,N_18088);
nor UO_604 (O_604,N_17215,N_16168);
nand UO_605 (O_605,N_18224,N_16231);
nor UO_606 (O_606,N_19698,N_19863);
nor UO_607 (O_607,N_17949,N_18717);
nand UO_608 (O_608,N_17741,N_16261);
and UO_609 (O_609,N_19301,N_19996);
nor UO_610 (O_610,N_19694,N_16734);
and UO_611 (O_611,N_16564,N_19087);
or UO_612 (O_612,N_18936,N_16398);
or UO_613 (O_613,N_19785,N_19744);
xor UO_614 (O_614,N_16939,N_19676);
and UO_615 (O_615,N_16117,N_19027);
or UO_616 (O_616,N_17218,N_18103);
xnor UO_617 (O_617,N_16813,N_17902);
or UO_618 (O_618,N_17245,N_16601);
nand UO_619 (O_619,N_16393,N_16346);
nor UO_620 (O_620,N_17186,N_18564);
and UO_621 (O_621,N_17825,N_17095);
xor UO_622 (O_622,N_18168,N_19363);
or UO_623 (O_623,N_18438,N_17353);
and UO_624 (O_624,N_18490,N_19461);
and UO_625 (O_625,N_16464,N_19830);
nor UO_626 (O_626,N_17520,N_17710);
nor UO_627 (O_627,N_16161,N_19199);
nor UO_628 (O_628,N_19042,N_17872);
nor UO_629 (O_629,N_19613,N_17595);
nor UO_630 (O_630,N_19248,N_16013);
and UO_631 (O_631,N_16959,N_18945);
or UO_632 (O_632,N_19177,N_17096);
xor UO_633 (O_633,N_16729,N_17224);
and UO_634 (O_634,N_18640,N_18009);
and UO_635 (O_635,N_17267,N_19463);
xnor UO_636 (O_636,N_17517,N_16981);
nand UO_637 (O_637,N_17754,N_16565);
nor UO_638 (O_638,N_18492,N_19331);
nor UO_639 (O_639,N_19178,N_18795);
nand UO_640 (O_640,N_17455,N_16568);
nand UO_641 (O_641,N_18888,N_18878);
xor UO_642 (O_642,N_17800,N_16750);
nand UO_643 (O_643,N_16133,N_17439);
and UO_644 (O_644,N_18147,N_16850);
nor UO_645 (O_645,N_17238,N_17583);
or UO_646 (O_646,N_19607,N_19226);
and UO_647 (O_647,N_18730,N_18835);
nor UO_648 (O_648,N_16263,N_19082);
nand UO_649 (O_649,N_19304,N_16387);
and UO_650 (O_650,N_17880,N_17388);
xor UO_651 (O_651,N_19635,N_16426);
nand UO_652 (O_652,N_16555,N_16589);
or UO_653 (O_653,N_18712,N_16651);
nor UO_654 (O_654,N_18865,N_18817);
or UO_655 (O_655,N_19109,N_18971);
nor UO_656 (O_656,N_16801,N_17856);
and UO_657 (O_657,N_18735,N_16262);
and UO_658 (O_658,N_19513,N_17854);
nor UO_659 (O_659,N_19404,N_18318);
nor UO_660 (O_660,N_19137,N_19674);
nor UO_661 (O_661,N_19136,N_18532);
and UO_662 (O_662,N_18919,N_16124);
nand UO_663 (O_663,N_19390,N_18510);
nor UO_664 (O_664,N_17420,N_18218);
nor UO_665 (O_665,N_18851,N_18281);
nor UO_666 (O_666,N_17771,N_17859);
nand UO_667 (O_667,N_16326,N_18410);
nand UO_668 (O_668,N_18367,N_19534);
nor UO_669 (O_669,N_17161,N_16741);
nand UO_670 (O_670,N_19516,N_18291);
nor UO_671 (O_671,N_18635,N_19703);
or UO_672 (O_672,N_18687,N_16391);
or UO_673 (O_673,N_18296,N_17723);
and UO_674 (O_674,N_18625,N_18783);
and UO_675 (O_675,N_17472,N_17118);
xor UO_676 (O_676,N_19219,N_17967);
nand UO_677 (O_677,N_16430,N_16659);
nand UO_678 (O_678,N_17493,N_16170);
nand UO_679 (O_679,N_17968,N_18886);
xnor UO_680 (O_680,N_19737,N_18725);
nand UO_681 (O_681,N_16704,N_19947);
nor UO_682 (O_682,N_19049,N_17614);
nor UO_683 (O_683,N_19701,N_17586);
nand UO_684 (O_684,N_16648,N_19258);
and UO_685 (O_685,N_19622,N_16712);
and UO_686 (O_686,N_16345,N_18773);
and UO_687 (O_687,N_19279,N_16079);
and UO_688 (O_688,N_16673,N_16369);
nand UO_689 (O_689,N_16544,N_17539);
and UO_690 (O_690,N_18778,N_19995);
nand UO_691 (O_691,N_18506,N_19129);
nand UO_692 (O_692,N_19318,N_19615);
or UO_693 (O_693,N_19056,N_17947);
nand UO_694 (O_694,N_18429,N_19142);
nor UO_695 (O_695,N_19542,N_19308);
xor UO_696 (O_696,N_16541,N_16643);
or UO_697 (O_697,N_16306,N_18633);
nor UO_698 (O_698,N_17568,N_16493);
nand UO_699 (O_699,N_17974,N_18292);
xor UO_700 (O_700,N_18864,N_19711);
nand UO_701 (O_701,N_16707,N_18089);
and UO_702 (O_702,N_16395,N_16434);
or UO_703 (O_703,N_16155,N_17722);
or UO_704 (O_704,N_17308,N_16219);
nor UO_705 (O_705,N_18164,N_17441);
and UO_706 (O_706,N_18465,N_19697);
and UO_707 (O_707,N_16943,N_19272);
nand UO_708 (O_708,N_17873,N_19925);
nand UO_709 (O_709,N_19008,N_17585);
nand UO_710 (O_710,N_18954,N_16794);
xor UO_711 (O_711,N_19659,N_19732);
or UO_712 (O_712,N_18528,N_19336);
nor UO_713 (O_713,N_19777,N_18021);
nor UO_714 (O_714,N_18843,N_18209);
or UO_715 (O_715,N_19237,N_18593);
xor UO_716 (O_716,N_17123,N_17391);
nor UO_717 (O_717,N_16419,N_16777);
or UO_718 (O_718,N_16689,N_16466);
and UO_719 (O_719,N_18478,N_16131);
nor UO_720 (O_720,N_17488,N_19097);
nor UO_721 (O_721,N_17674,N_18330);
nor UO_722 (O_722,N_17086,N_17103);
nand UO_723 (O_723,N_19062,N_18663);
xnor UO_724 (O_724,N_18997,N_16985);
or UO_725 (O_725,N_16195,N_17282);
nor UO_726 (O_726,N_18195,N_19377);
or UO_727 (O_727,N_19439,N_18250);
or UO_728 (O_728,N_18498,N_16915);
nand UO_729 (O_729,N_17232,N_16021);
nand UO_730 (O_730,N_18809,N_18356);
and UO_731 (O_731,N_18558,N_18867);
or UO_732 (O_732,N_16630,N_19452);
and UO_733 (O_733,N_16074,N_17717);
nand UO_734 (O_734,N_17745,N_16535);
or UO_735 (O_735,N_19261,N_18600);
nand UO_736 (O_736,N_16593,N_18184);
xnor UO_737 (O_737,N_17030,N_16570);
nor UO_738 (O_738,N_16556,N_17158);
nor UO_739 (O_739,N_18002,N_18695);
or UO_740 (O_740,N_18208,N_18353);
nand UO_741 (O_741,N_17842,N_17270);
nor UO_742 (O_742,N_19624,N_19003);
or UO_743 (O_743,N_18903,N_18950);
nand UO_744 (O_744,N_18434,N_18117);
and UO_745 (O_745,N_18451,N_17725);
xor UO_746 (O_746,N_19640,N_17371);
or UO_747 (O_747,N_19918,N_18011);
nor UO_748 (O_748,N_16647,N_16918);
nand UO_749 (O_749,N_19077,N_19281);
and UO_750 (O_750,N_16736,N_17552);
and UO_751 (O_751,N_19303,N_17048);
nor UO_752 (O_752,N_17654,N_17421);
nor UO_753 (O_753,N_19196,N_16015);
and UO_754 (O_754,N_19340,N_16197);
or UO_755 (O_755,N_16287,N_16358);
and UO_756 (O_756,N_19367,N_19873);
nor UO_757 (O_757,N_16098,N_17829);
nand UO_758 (O_758,N_17743,N_17337);
and UO_759 (O_759,N_17994,N_16658);
nor UO_760 (O_760,N_16586,N_17077);
or UO_761 (O_761,N_17787,N_18899);
and UO_762 (O_762,N_18157,N_17715);
nand UO_763 (O_763,N_19637,N_18181);
nor UO_764 (O_764,N_18051,N_18326);
and UO_765 (O_765,N_18705,N_18832);
or UO_766 (O_766,N_17518,N_16703);
and UO_767 (O_767,N_19438,N_16410);
xor UO_768 (O_768,N_16858,N_17706);
nor UO_769 (O_769,N_19573,N_17628);
or UO_770 (O_770,N_16500,N_19955);
or UO_771 (O_771,N_18263,N_19231);
nor UO_772 (O_772,N_19065,N_17209);
nor UO_773 (O_773,N_16228,N_16600);
and UO_774 (O_774,N_19931,N_19636);
nor UO_775 (O_775,N_18162,N_19770);
nand UO_776 (O_776,N_16199,N_19811);
or UO_777 (O_777,N_18358,N_19717);
nand UO_778 (O_778,N_19174,N_16606);
and UO_779 (O_779,N_19379,N_18350);
nand UO_780 (O_780,N_18323,N_17600);
xor UO_781 (O_781,N_19033,N_17510);
or UO_782 (O_782,N_19418,N_17925);
xnor UO_783 (O_783,N_17954,N_19016);
nand UO_784 (O_784,N_16244,N_19421);
or UO_785 (O_785,N_19521,N_17356);
nor UO_786 (O_786,N_19714,N_17844);
xnor UO_787 (O_787,N_18940,N_16014);
and UO_788 (O_788,N_18142,N_18020);
nor UO_789 (O_789,N_19427,N_19247);
xor UO_790 (O_790,N_19164,N_16000);
nand UO_791 (O_791,N_19310,N_18728);
nand UO_792 (O_792,N_19532,N_18123);
and UO_793 (O_793,N_17588,N_18099);
or UO_794 (O_794,N_17524,N_16577);
xor UO_795 (O_795,N_19073,N_17649);
and UO_796 (O_796,N_19671,N_16844);
nand UO_797 (O_797,N_19113,N_18242);
and UO_798 (O_798,N_18087,N_18025);
or UO_799 (O_799,N_17946,N_17775);
nor UO_800 (O_800,N_18869,N_18090);
and UO_801 (O_801,N_17990,N_19747);
nand UO_802 (O_802,N_16112,N_18101);
and UO_803 (O_803,N_17869,N_18741);
and UO_804 (O_804,N_18584,N_17080);
and UO_805 (O_805,N_17610,N_18608);
nand UO_806 (O_806,N_17690,N_19424);
nor UO_807 (O_807,N_18870,N_17026);
or UO_808 (O_808,N_19540,N_16706);
nor UO_809 (O_809,N_19909,N_19431);
or UO_810 (O_810,N_16655,N_16251);
nand UO_811 (O_811,N_18283,N_16830);
or UO_812 (O_812,N_16033,N_18343);
nor UO_813 (O_813,N_18325,N_19193);
and UO_814 (O_814,N_19621,N_19826);
xor UO_815 (O_815,N_18255,N_17832);
nor UO_816 (O_816,N_17536,N_17160);
nor UO_817 (O_817,N_16721,N_18710);
and UO_818 (O_818,N_17213,N_18174);
or UO_819 (O_819,N_16313,N_19992);
and UO_820 (O_820,N_17368,N_18592);
nand UO_821 (O_821,N_16723,N_19924);
nand UO_822 (O_822,N_19498,N_18980);
nor UO_823 (O_823,N_19322,N_19684);
xnor UO_824 (O_824,N_16953,N_19332);
nor UO_825 (O_825,N_18137,N_18309);
nor UO_826 (O_826,N_17061,N_16106);
nor UO_827 (O_827,N_17168,N_16049);
and UO_828 (O_828,N_16181,N_18830);
and UO_829 (O_829,N_16148,N_19202);
and UO_830 (O_830,N_19997,N_18653);
and UO_831 (O_831,N_16728,N_17830);
nand UO_832 (O_832,N_18267,N_18898);
nor UO_833 (O_833,N_17855,N_16233);
nor UO_834 (O_834,N_19647,N_19490);
xnor UO_835 (O_835,N_17417,N_19901);
or UO_836 (O_836,N_16095,N_18124);
nor UO_837 (O_837,N_19691,N_19343);
xor UO_838 (O_838,N_18091,N_18862);
nor UO_839 (O_839,N_16627,N_19954);
or UO_840 (O_840,N_16977,N_18912);
xor UO_841 (O_841,N_19217,N_18514);
nor UO_842 (O_842,N_19812,N_17405);
xnor UO_843 (O_843,N_19539,N_18133);
nand UO_844 (O_844,N_16424,N_17297);
and UO_845 (O_845,N_16910,N_18975);
nand UO_846 (O_846,N_19837,N_17602);
xor UO_847 (O_847,N_19875,N_18307);
and UO_848 (O_848,N_17311,N_19149);
and UO_849 (O_849,N_17656,N_18261);
xnor UO_850 (O_850,N_18289,N_19907);
nor UO_851 (O_851,N_19416,N_19169);
nor UO_852 (O_852,N_18786,N_17336);
or UO_853 (O_853,N_16892,N_16871);
and UO_854 (O_854,N_19189,N_17377);
or UO_855 (O_855,N_19544,N_18505);
nand UO_856 (O_856,N_17714,N_17025);
xnor UO_857 (O_857,N_19163,N_17997);
or UO_858 (O_858,N_16688,N_19764);
or UO_859 (O_859,N_16745,N_17164);
nor UO_860 (O_860,N_16889,N_17304);
xnor UO_861 (O_861,N_16752,N_16957);
nand UO_862 (O_862,N_16143,N_17056);
or UO_863 (O_863,N_17921,N_18397);
and UO_864 (O_864,N_18093,N_17572);
nor UO_865 (O_865,N_18570,N_18389);
nor UO_866 (O_866,N_17952,N_18085);
and UO_867 (O_867,N_16101,N_19563);
nand UO_868 (O_868,N_18152,N_16584);
nand UO_869 (O_869,N_17864,N_19556);
xnor UO_870 (O_870,N_18048,N_17623);
or UO_871 (O_871,N_19326,N_19959);
or UO_872 (O_872,N_19759,N_18297);
nor UO_873 (O_873,N_18071,N_18468);
nor UO_874 (O_874,N_17814,N_19751);
nand UO_875 (O_875,N_19342,N_19274);
or UO_876 (O_876,N_18569,N_16574);
xnor UO_877 (O_877,N_18304,N_18489);
nor UO_878 (O_878,N_16077,N_16289);
and UO_879 (O_879,N_18107,N_16225);
nand UO_880 (O_880,N_16807,N_17108);
nor UO_881 (O_881,N_19976,N_17670);
xor UO_882 (O_882,N_18173,N_16868);
nor UO_883 (O_883,N_19031,N_16091);
and UO_884 (O_884,N_19392,N_18342);
or UO_885 (O_885,N_19887,N_19998);
nor UO_886 (O_886,N_17680,N_16088);
nand UO_887 (O_887,N_17222,N_18128);
nand UO_888 (O_888,N_19792,N_16756);
and UO_889 (O_889,N_16389,N_17559);
nand UO_890 (O_890,N_19820,N_16151);
and UO_891 (O_891,N_17849,N_16805);
nand UO_892 (O_892,N_19333,N_19680);
nor UO_893 (O_893,N_17014,N_17427);
nor UO_894 (O_894,N_18114,N_18989);
and UO_895 (O_895,N_18948,N_19922);
nand UO_896 (O_896,N_18440,N_16697);
and UO_897 (O_897,N_16123,N_16475);
nor UO_898 (O_898,N_19364,N_17263);
nand UO_899 (O_899,N_18185,N_18858);
and UO_900 (O_900,N_16362,N_17971);
and UO_901 (O_901,N_18972,N_19591);
nor UO_902 (O_902,N_16041,N_19710);
nor UO_903 (O_903,N_16991,N_17635);
xnor UO_904 (O_904,N_16663,N_19974);
nand UO_905 (O_905,N_17375,N_17352);
or UO_906 (O_906,N_16971,N_18234);
nor UO_907 (O_907,N_18165,N_18894);
nor UO_908 (O_908,N_16791,N_16336);
and UO_909 (O_909,N_16146,N_17070);
nand UO_910 (O_910,N_16276,N_18791);
nor UO_911 (O_911,N_19372,N_18460);
and UO_912 (O_912,N_19882,N_17231);
nand UO_913 (O_913,N_16992,N_19964);
or UO_914 (O_914,N_18136,N_18257);
nor UO_915 (O_915,N_19473,N_17021);
nor UO_916 (O_916,N_16159,N_18883);
nand UO_917 (O_917,N_18131,N_17561);
nor UO_918 (O_918,N_19898,N_16229);
nor UO_919 (O_919,N_16340,N_19977);
nand UO_920 (O_920,N_18249,N_18956);
nand UO_921 (O_921,N_18802,N_19388);
and UO_922 (O_922,N_16536,N_16023);
or UO_923 (O_923,N_18907,N_18842);
nor UO_924 (O_924,N_17930,N_17345);
nand UO_925 (O_925,N_19409,N_18904);
nor UO_926 (O_926,N_19184,N_16526);
or UO_927 (O_927,N_19289,N_19089);
nor UO_928 (O_928,N_18880,N_17645);
and UO_929 (O_929,N_17342,N_19375);
nand UO_930 (O_930,N_18946,N_17893);
nor UO_931 (O_931,N_17470,N_17305);
or UO_932 (O_932,N_17637,N_16324);
nand UO_933 (O_933,N_19121,N_16043);
or UO_934 (O_934,N_18096,N_18990);
xnor UO_935 (O_935,N_17995,N_19254);
nand UO_936 (O_936,N_16094,N_17058);
or UO_937 (O_937,N_19543,N_19130);
or UO_938 (O_938,N_17897,N_16105);
xnor UO_939 (O_939,N_18768,N_16662);
or UO_940 (O_940,N_18678,N_16837);
nand UO_941 (O_941,N_16067,N_19300);
nor UO_942 (O_942,N_19848,N_17235);
or UO_943 (O_943,N_16504,N_19466);
nand UO_944 (O_944,N_18422,N_19523);
and UO_945 (O_945,N_16350,N_18146);
nor UO_946 (O_946,N_18175,N_17611);
nor UO_947 (O_947,N_16666,N_19160);
nor UO_948 (O_948,N_18495,N_18706);
nor UO_949 (O_949,N_18373,N_17701);
and UO_950 (O_950,N_18807,N_17252);
or UO_951 (O_951,N_19358,N_16144);
nor UO_952 (O_952,N_18158,N_17543);
xnor UO_953 (O_953,N_16099,N_19391);
nor UO_954 (O_954,N_19561,N_16761);
xnor UO_955 (O_955,N_18974,N_18265);
and UO_956 (O_956,N_18754,N_19071);
or UO_957 (O_957,N_19396,N_16549);
nand UO_958 (O_958,N_19230,N_16076);
and UO_959 (O_959,N_19368,N_16900);
nor UO_960 (O_960,N_17359,N_17763);
or UO_961 (O_961,N_17769,N_16238);
nor UO_962 (O_962,N_16039,N_18251);
nand UO_963 (O_963,N_19991,N_19050);
and UO_964 (O_964,N_19273,N_17210);
or UO_965 (O_965,N_16187,N_19929);
nand UO_966 (O_966,N_18385,N_19596);
and UO_967 (O_967,N_16451,N_17795);
and UO_968 (O_968,N_17496,N_18408);
nor UO_969 (O_969,N_17169,N_19155);
or UO_970 (O_970,N_18750,N_16086);
or UO_971 (O_971,N_19118,N_18315);
xor UO_972 (O_972,N_18402,N_16163);
or UO_973 (O_973,N_16885,N_16865);
and UO_974 (O_974,N_19879,N_16310);
xnor UO_975 (O_975,N_19067,N_16301);
nor UO_976 (O_976,N_16684,N_19590);
and UO_977 (O_977,N_17448,N_19350);
or UO_978 (O_978,N_17957,N_18910);
xnor UO_979 (O_979,N_19905,N_16588);
xor UO_980 (O_980,N_16207,N_16242);
and UO_981 (O_981,N_16733,N_19028);
or UO_982 (O_982,N_18456,N_17927);
nand UO_983 (O_983,N_18993,N_17085);
or UO_984 (O_984,N_19632,N_17212);
and UO_985 (O_985,N_19362,N_19530);
and UO_986 (O_986,N_17243,N_19054);
or UO_987 (O_987,N_18871,N_16455);
or UO_988 (O_988,N_18688,N_16270);
xor UO_989 (O_989,N_16411,N_19257);
nand UO_990 (O_990,N_17239,N_17459);
nor UO_991 (O_991,N_18274,N_16983);
nor UO_992 (O_992,N_17495,N_17147);
nor UO_993 (O_993,N_18018,N_17806);
nor UO_994 (O_994,N_19605,N_17285);
nor UO_995 (O_995,N_19816,N_17034);
and UO_996 (O_996,N_16962,N_17481);
and UO_997 (O_997,N_19814,N_16873);
xor UO_998 (O_998,N_16631,N_19614);
and UO_999 (O_999,N_16003,N_17155);
and UO_1000 (O_1000,N_17970,N_18271);
or UO_1001 (O_1001,N_17860,N_18229);
or UO_1002 (O_1002,N_17355,N_16331);
and UO_1003 (O_1003,N_19103,N_17780);
nand UO_1004 (O_1004,N_19205,N_18582);
and UO_1005 (O_1005,N_19381,N_19578);
nand UO_1006 (O_1006,N_18398,N_18759);
nor UO_1007 (O_1007,N_17760,N_18591);
nor UO_1008 (O_1008,N_16694,N_19020);
nand UO_1009 (O_1009,N_18227,N_19445);
nor UO_1010 (O_1010,N_19665,N_19948);
nand UO_1011 (O_1011,N_18987,N_17823);
and UO_1012 (O_1012,N_18381,N_19943);
nand UO_1013 (O_1013,N_19831,N_19825);
or UO_1014 (O_1014,N_17629,N_19157);
nand UO_1015 (O_1015,N_18793,N_16632);
xnor UO_1016 (O_1016,N_19892,N_18454);
xnor UO_1017 (O_1017,N_17283,N_18978);
nand UO_1018 (O_1018,N_16849,N_19176);
or UO_1019 (O_1019,N_16516,N_17944);
nand UO_1020 (O_1020,N_16758,N_16996);
and UO_1021 (O_1021,N_17363,N_19296);
xnor UO_1022 (O_1022,N_19004,N_17254);
xnor UO_1023 (O_1023,N_18632,N_18177);
nor UO_1024 (O_1024,N_16368,N_16330);
xnor UO_1025 (O_1025,N_18915,N_17237);
nor UO_1026 (O_1026,N_17499,N_17200);
nand UO_1027 (O_1027,N_16469,N_19146);
and UO_1028 (O_1028,N_16890,N_18694);
xnor UO_1029 (O_1029,N_19639,N_17416);
nor UO_1030 (O_1030,N_16418,N_17001);
or UO_1031 (O_1031,N_17707,N_17719);
nor UO_1032 (O_1032,N_16732,N_19765);
xnor UO_1033 (O_1033,N_16089,N_17870);
nand UO_1034 (O_1034,N_16984,N_18149);
and UO_1035 (O_1035,N_18850,N_18689);
nor UO_1036 (O_1036,N_19030,N_16864);
xnor UO_1037 (O_1037,N_18210,N_19538);
nand UO_1038 (O_1038,N_17937,N_16677);
or UO_1039 (O_1039,N_19110,N_18827);
nor UO_1040 (O_1040,N_17244,N_16171);
nor UO_1041 (O_1041,N_19541,N_18884);
or UO_1042 (O_1042,N_16190,N_17338);
or UO_1043 (O_1043,N_17091,N_18703);
xor UO_1044 (O_1044,N_17876,N_19492);
xor UO_1045 (O_1045,N_18630,N_18140);
nor UO_1046 (O_1046,N_19889,N_16279);
or UO_1047 (O_1047,N_18917,N_16811);
and UO_1048 (O_1048,N_19499,N_17176);
and UO_1049 (O_1049,N_16142,N_17956);
nand UO_1050 (O_1050,N_17545,N_17394);
xor UO_1051 (O_1051,N_16361,N_17528);
nand UO_1052 (O_1052,N_17850,N_17640);
nand UO_1053 (O_1053,N_18496,N_18777);
or UO_1054 (O_1054,N_17398,N_18567);
xor UO_1055 (O_1055,N_16521,N_19280);
nor UO_1056 (O_1056,N_19857,N_18620);
nand UO_1057 (O_1057,N_17310,N_16373);
and UO_1058 (O_1058,N_19245,N_17247);
or UO_1059 (O_1059,N_16523,N_16824);
nand UO_1060 (O_1060,N_19360,N_19979);
xnor UO_1061 (O_1061,N_16004,N_19188);
or UO_1062 (O_1062,N_16386,N_18364);
nor UO_1063 (O_1063,N_16394,N_17621);
nor UO_1064 (O_1064,N_16065,N_17506);
and UO_1065 (O_1065,N_19555,N_19061);
and UO_1066 (O_1066,N_18921,N_17225);
nand UO_1067 (O_1067,N_18125,N_16486);
nor UO_1068 (O_1068,N_16919,N_18943);
and UO_1069 (O_1069,N_18631,N_19168);
and UO_1070 (O_1070,N_19150,N_18369);
and UO_1071 (O_1071,N_18651,N_16572);
nor UO_1072 (O_1072,N_17752,N_18348);
nor UO_1073 (O_1073,N_17256,N_17742);
and UO_1074 (O_1074,N_18815,N_19597);
or UO_1075 (O_1075,N_18228,N_17253);
and UO_1076 (O_1076,N_18494,N_17016);
nand UO_1077 (O_1077,N_16967,N_19330);
and UO_1078 (O_1078,N_18765,N_18875);
nor UO_1079 (O_1079,N_18581,N_16623);
xor UO_1080 (O_1080,N_19519,N_19458);
nand UO_1081 (O_1081,N_17547,N_18799);
xnor UO_1082 (O_1082,N_16838,N_19655);
or UO_1083 (O_1083,N_17596,N_16232);
nand UO_1084 (O_1084,N_16819,N_17134);
or UO_1085 (O_1085,N_17612,N_17020);
and UO_1086 (O_1086,N_19471,N_19719);
nor UO_1087 (O_1087,N_17766,N_18916);
nor UO_1088 (O_1088,N_17319,N_17782);
or UO_1089 (O_1089,N_18404,N_19559);
nor UO_1090 (O_1090,N_17196,N_18605);
or UO_1091 (O_1091,N_16912,N_19286);
or UO_1092 (O_1092,N_17555,N_17172);
nand UO_1093 (O_1093,N_17885,N_18808);
xnor UO_1094 (O_1094,N_17099,N_16179);
or UO_1095 (O_1095,N_16784,N_17278);
or UO_1096 (O_1096,N_19366,N_16763);
nor UO_1097 (O_1097,N_18779,N_19104);
and UO_1098 (O_1098,N_17150,N_17068);
nor UO_1099 (O_1099,N_17248,N_17106);
nand UO_1100 (O_1100,N_17329,N_18186);
or UO_1101 (O_1101,N_19446,N_17107);
nand UO_1102 (O_1102,N_19935,N_16998);
or UO_1103 (O_1103,N_16254,N_19916);
nor UO_1104 (O_1104,N_19687,N_17227);
nor UO_1105 (O_1105,N_19039,N_17903);
and UO_1106 (O_1106,N_19750,N_18578);
nor UO_1107 (O_1107,N_18260,N_19617);
or UO_1108 (O_1108,N_19618,N_18305);
or UO_1109 (O_1109,N_18126,N_17145);
nand UO_1110 (O_1110,N_17498,N_19093);
xor UO_1111 (O_1111,N_16399,N_19275);
xnor UO_1112 (O_1112,N_18621,N_19967);
and UO_1113 (O_1113,N_19819,N_17863);
or UO_1114 (O_1114,N_16017,N_19255);
or UO_1115 (O_1115,N_19896,N_19734);
nor UO_1116 (O_1116,N_17309,N_18939);
and UO_1117 (O_1117,N_19365,N_19085);
or UO_1118 (O_1118,N_16881,N_16637);
or UO_1119 (O_1119,N_17033,N_16284);
and UO_1120 (O_1120,N_18349,N_17018);
xor UO_1121 (O_1121,N_16070,N_19159);
nand UO_1122 (O_1122,N_17265,N_19807);
or UO_1123 (O_1123,N_16917,N_18618);
or UO_1124 (O_1124,N_19236,N_17299);
nor UO_1125 (O_1125,N_16639,N_18416);
nor UO_1126 (O_1126,N_16829,N_17724);
xor UO_1127 (O_1127,N_16520,N_17721);
and UO_1128 (O_1128,N_16767,N_17704);
nor UO_1129 (O_1129,N_19395,N_16031);
nand UO_1130 (O_1130,N_19410,N_17230);
xnor UO_1131 (O_1131,N_16656,N_16388);
or UO_1132 (O_1132,N_19577,N_18387);
or UO_1133 (O_1133,N_16921,N_17755);
nor UO_1134 (O_1134,N_18477,N_16653);
and UO_1135 (O_1135,N_16800,N_18143);
or UO_1136 (O_1136,N_18816,N_16063);
nor UO_1137 (O_1137,N_16423,N_17241);
or UO_1138 (O_1138,N_19579,N_18362);
and UO_1139 (O_1139,N_16713,N_19804);
and UO_1140 (O_1140,N_19945,N_19678);
or UO_1141 (O_1141,N_16403,N_18599);
or UO_1142 (O_1142,N_16260,N_17644);
nand UO_1143 (O_1143,N_17041,N_19092);
or UO_1144 (O_1144,N_16044,N_16573);
nand UO_1145 (O_1145,N_18918,N_17228);
or UO_1146 (O_1146,N_19801,N_16719);
nand UO_1147 (O_1147,N_18709,N_16720);
nor UO_1148 (O_1148,N_17793,N_17551);
and UO_1149 (O_1149,N_17332,N_19756);
nand UO_1150 (O_1150,N_17920,N_16011);
nor UO_1151 (O_1151,N_16194,N_19999);
or UO_1152 (O_1152,N_19850,N_16010);
or UO_1153 (O_1153,N_19839,N_17380);
and UO_1154 (O_1154,N_16665,N_17452);
and UO_1155 (O_1155,N_17702,N_19969);
or UO_1156 (O_1156,N_18377,N_19002);
nand UO_1157 (O_1157,N_19413,N_16156);
or UO_1158 (O_1158,N_18798,N_18671);
or UO_1159 (O_1159,N_19511,N_16875);
and UO_1160 (O_1160,N_16803,N_17264);
nor UO_1161 (O_1161,N_17482,N_16870);
or UO_1162 (O_1162,N_16936,N_19213);
and UO_1163 (O_1163,N_19988,N_17682);
nand UO_1164 (O_1164,N_17650,N_16509);
nand UO_1165 (O_1165,N_16209,N_19270);
nand UO_1166 (O_1166,N_17011,N_16147);
xnor UO_1167 (O_1167,N_16700,N_18995);
and UO_1168 (O_1168,N_18831,N_19497);
nand UO_1169 (O_1169,N_16863,N_19884);
nor UO_1170 (O_1170,N_18516,N_18482);
nand UO_1171 (O_1171,N_16443,N_16184);
nor UO_1172 (O_1172,N_16165,N_18344);
and UO_1173 (O_1173,N_16933,N_18180);
and UO_1174 (O_1174,N_16510,N_17500);
or UO_1175 (O_1175,N_19749,N_17907);
or UO_1176 (O_1176,N_18673,N_17318);
and UO_1177 (O_1177,N_17989,N_17314);
and UO_1178 (O_1178,N_19921,N_18587);
or UO_1179 (O_1179,N_16297,N_17986);
and UO_1180 (O_1180,N_19349,N_17950);
nor UO_1181 (O_1181,N_16816,N_18003);
nor UO_1182 (O_1182,N_17280,N_16055);
and UO_1183 (O_1183,N_18167,N_17657);
and UO_1184 (O_1184,N_16210,N_17573);
or UO_1185 (O_1185,N_18458,N_17581);
and UO_1186 (O_1186,N_19768,N_18588);
and UO_1187 (O_1187,N_19244,N_16383);
nand UO_1188 (O_1188,N_17993,N_17772);
xnor UO_1189 (O_1189,N_16714,N_16237);
or UO_1190 (O_1190,N_16020,N_19533);
and UO_1191 (O_1191,N_16603,N_19900);
or UO_1192 (O_1192,N_16934,N_18270);
nand UO_1193 (O_1193,N_17347,N_16256);
xor UO_1194 (O_1194,N_19311,N_19143);
nand UO_1195 (O_1195,N_17905,N_17430);
or UO_1196 (O_1196,N_17908,N_16160);
or UO_1197 (O_1197,N_16245,N_18462);
and UO_1198 (O_1198,N_19599,N_16854);
or UO_1199 (O_1199,N_18262,N_19856);
nor UO_1200 (O_1200,N_18189,N_19566);
nand UO_1201 (O_1201,N_19965,N_19950);
and UO_1202 (O_1202,N_17132,N_17601);
and UO_1203 (O_1203,N_17736,N_18520);
or UO_1204 (O_1204,N_18436,N_17206);
nand UO_1205 (O_1205,N_16318,N_16001);
nand UO_1206 (O_1206,N_16905,N_16896);
nor UO_1207 (O_1207,N_17973,N_17984);
nand UO_1208 (O_1208,N_17942,N_17726);
or UO_1209 (O_1209,N_19971,N_18205);
and UO_1210 (O_1210,N_17679,N_17632);
or UO_1211 (O_1211,N_17374,N_16258);
nor UO_1212 (O_1212,N_18836,N_16255);
or UO_1213 (O_1213,N_16137,N_17789);
and UO_1214 (O_1214,N_19718,N_19080);
nand UO_1215 (O_1215,N_19806,N_19214);
nand UO_1216 (O_1216,N_19246,N_16484);
or UO_1217 (O_1217,N_17179,N_18775);
and UO_1218 (O_1218,N_18923,N_18589);
and UO_1219 (O_1219,N_16683,N_19162);
nor UO_1220 (O_1220,N_17295,N_16650);
nor UO_1221 (O_1221,N_18118,N_16492);
nor UO_1222 (O_1222,N_18193,N_19357);
or UO_1223 (O_1223,N_18225,N_16296);
or UO_1224 (O_1224,N_17399,N_16380);
nand UO_1225 (O_1225,N_19980,N_18119);
or UO_1226 (O_1226,N_19780,N_18655);
or UO_1227 (O_1227,N_18601,N_17931);
nor UO_1228 (O_1228,N_19838,N_16191);
or UO_1229 (O_1229,N_18650,N_19840);
or UO_1230 (O_1230,N_16140,N_18050);
or UO_1231 (O_1231,N_18746,N_16667);
and UO_1232 (O_1232,N_17550,N_16961);
nor UO_1233 (O_1233,N_17202,N_16042);
or UO_1234 (O_1234,N_18604,N_16220);
or UO_1235 (O_1235,N_16771,N_16381);
nor UO_1236 (O_1236,N_19666,N_17566);
and UO_1237 (O_1237,N_19256,N_19752);
or UO_1238 (O_1238,N_19951,N_17716);
and UO_1239 (O_1239,N_17211,N_19276);
nor UO_1240 (O_1240,N_19700,N_18459);
or UO_1241 (O_1241,N_16071,N_16085);
xnor UO_1242 (O_1242,N_17395,N_18030);
and UO_1243 (O_1243,N_19619,N_19052);
or UO_1244 (O_1244,N_17251,N_17462);
nand UO_1245 (O_1245,N_16211,N_18753);
nor UO_1246 (O_1246,N_17693,N_18068);
and UO_1247 (O_1247,N_18329,N_16609);
nor UO_1248 (O_1248,N_19116,N_19779);
or UO_1249 (O_1249,N_18652,N_17590);
nor UO_1250 (O_1250,N_16483,N_19268);
and UO_1251 (O_1251,N_16668,N_19914);
nand UO_1252 (O_1252,N_17322,N_17661);
or UO_1253 (O_1253,N_18425,N_16218);
xnor UO_1254 (O_1254,N_18958,N_19307);
nand UO_1255 (O_1255,N_19267,N_17019);
or UO_1256 (O_1256,N_16090,N_19783);
nor UO_1257 (O_1257,N_19895,N_17677);
nand UO_1258 (O_1258,N_19201,N_18803);
or UO_1259 (O_1259,N_18221,N_16174);
or UO_1260 (O_1260,N_19405,N_18788);
nand UO_1261 (O_1261,N_18098,N_16433);
nor UO_1262 (O_1262,N_19415,N_18022);
and UO_1263 (O_1263,N_19114,N_19069);
xnor UO_1264 (O_1264,N_18027,N_17349);
or UO_1265 (O_1265,N_19161,N_17605);
nor UO_1266 (O_1266,N_19309,N_18233);
nor UO_1267 (O_1267,N_18378,N_19982);
nand UO_1268 (O_1268,N_18854,N_18614);
nand UO_1269 (O_1269,N_19772,N_19317);
nor UO_1270 (O_1270,N_17404,N_16940);
xor UO_1271 (O_1271,N_17271,N_17015);
xor UO_1272 (O_1272,N_18169,N_17494);
nor UO_1273 (O_1273,N_17350,N_19949);
or UO_1274 (O_1274,N_19447,N_18038);
nor UO_1275 (O_1275,N_19334,N_17540);
nor UO_1276 (O_1276,N_18841,N_16385);
or UO_1277 (O_1277,N_19444,N_16087);
nand UO_1278 (O_1278,N_18337,N_18634);
and UO_1279 (O_1279,N_18037,N_16152);
nand UO_1280 (O_1280,N_18547,N_16935);
and UO_1281 (O_1281,N_17659,N_16384);
nor UO_1282 (O_1282,N_16135,N_17109);
nor UO_1283 (O_1283,N_17732,N_17882);
xnor UO_1284 (O_1284,N_17694,N_18418);
xor UO_1285 (O_1285,N_17475,N_17067);
and UO_1286 (O_1286,N_16018,N_19771);
xor UO_1287 (O_1287,N_19385,N_18824);
nor UO_1288 (O_1288,N_16557,N_16080);
and UO_1289 (O_1289,N_18924,N_17389);
nand UO_1290 (O_1290,N_18409,N_19878);
nand UO_1291 (O_1291,N_16366,N_18431);
or UO_1292 (O_1292,N_18198,N_17330);
or UO_1293 (O_1293,N_17928,N_17233);
or UO_1294 (O_1294,N_17249,N_18925);
or UO_1295 (O_1295,N_16113,N_16303);
and UO_1296 (O_1296,N_18833,N_17344);
nand UO_1297 (O_1297,N_18550,N_18748);
and UO_1298 (O_1298,N_16792,N_18876);
or UO_1299 (O_1299,N_16848,N_19064);
nand UO_1300 (O_1300,N_17324,N_17445);
or UO_1301 (O_1301,N_17120,N_17144);
xnor UO_1302 (O_1302,N_19125,N_19913);
xnor UO_1303 (O_1303,N_18277,N_16809);
nand UO_1304 (O_1304,N_16422,N_17364);
and UO_1305 (O_1305,N_18955,N_18354);
or UO_1306 (O_1306,N_18937,N_17289);
or UO_1307 (O_1307,N_17273,N_19374);
or UO_1308 (O_1308,N_19627,N_16468);
and UO_1309 (O_1309,N_16446,N_19282);
nand UO_1310 (O_1310,N_17435,N_17443);
and UO_1311 (O_1311,N_18698,N_17089);
nor UO_1312 (O_1312,N_18151,N_18541);
nand UO_1313 (O_1313,N_18187,N_16539);
nand UO_1314 (O_1314,N_18914,N_18573);
nor UO_1315 (O_1315,N_19654,N_17357);
nor UO_1316 (O_1316,N_18509,N_17576);
or UO_1317 (O_1317,N_18930,N_19728);
or UO_1318 (O_1318,N_17433,N_18846);
nand UO_1319 (O_1319,N_18220,N_16474);
nor UO_1320 (O_1320,N_16920,N_18070);
or UO_1321 (O_1321,N_18199,N_17881);
nand UO_1322 (O_1322,N_17615,N_19394);
or UO_1323 (O_1323,N_17346,N_19220);
nor UO_1324 (O_1324,N_18965,N_16649);
nand UO_1325 (O_1325,N_19864,N_19508);
nor UO_1326 (O_1326,N_19781,N_19491);
nor UO_1327 (O_1327,N_16432,N_16405);
nand UO_1328 (O_1328,N_18766,N_18772);
nor UO_1329 (O_1329,N_18985,N_18856);
xor UO_1330 (O_1330,N_18860,N_19581);
or UO_1331 (O_1331,N_18659,N_16843);
or UO_1332 (O_1332,N_16545,N_17525);
nor UO_1333 (O_1333,N_17316,N_16941);
and UO_1334 (O_1334,N_16059,N_17208);
and UO_1335 (O_1335,N_19012,N_16569);
nand UO_1336 (O_1336,N_17794,N_16364);
nand UO_1337 (O_1337,N_17936,N_18928);
nor UO_1338 (O_1338,N_16339,N_18446);
or UO_1339 (O_1339,N_17410,N_16213);
nor UO_1340 (O_1340,N_17810,N_16581);
nand UO_1341 (O_1341,N_16121,N_19106);
nor UO_1342 (O_1342,N_18757,N_16227);
nor UO_1343 (O_1343,N_16904,N_17924);
and UO_1344 (O_1344,N_16976,N_16797);
nor UO_1345 (O_1345,N_17817,N_19210);
or UO_1346 (O_1346,N_18258,N_19960);
and UO_1347 (O_1347,N_18012,N_18572);
nor UO_1348 (O_1348,N_19060,N_16212);
or UO_1349 (O_1349,N_19420,N_17537);
nand UO_1350 (O_1350,N_16855,N_17504);
nor UO_1351 (O_1351,N_17554,N_19419);
nand UO_1352 (O_1352,N_19260,N_17900);
and UO_1353 (O_1353,N_18932,N_17140);
and UO_1354 (O_1354,N_17734,N_17579);
nor UO_1355 (O_1355,N_16272,N_17643);
or UO_1356 (O_1356,N_19844,N_16672);
and UO_1357 (O_1357,N_19197,N_19536);
nor UO_1358 (O_1358,N_16591,N_18327);
or UO_1359 (O_1359,N_16744,N_16130);
nor UO_1360 (O_1360,N_18857,N_19853);
and UO_1361 (O_1361,N_16866,N_16566);
or UO_1362 (O_1362,N_18623,N_16579);
nand UO_1363 (O_1363,N_19251,N_17366);
and UO_1364 (O_1364,N_18029,N_17128);
nand UO_1365 (O_1365,N_16644,N_16068);
nor UO_1366 (O_1366,N_19218,N_19670);
and UO_1367 (O_1367,N_19766,N_17562);
nor UO_1368 (O_1368,N_18112,N_18739);
and UO_1369 (O_1369,N_17320,N_17035);
and UO_1370 (O_1370,N_17636,N_19537);
nor UO_1371 (O_1371,N_19128,N_17642);
and UO_1372 (O_1372,N_17932,N_18853);
nand UO_1373 (O_1373,N_16922,N_18202);
nand UO_1374 (O_1374,N_17327,N_19788);
and UO_1375 (O_1375,N_18316,N_17808);
or UO_1376 (O_1376,N_16832,N_19459);
and UO_1377 (O_1377,N_19634,N_18957);
and UO_1378 (O_1378,N_17136,N_18729);
nor UO_1379 (O_1379,N_19662,N_17423);
and UO_1380 (O_1380,N_16993,N_17236);
and UO_1381 (O_1381,N_19355,N_18413);
or UO_1382 (O_1382,N_18013,N_19558);
nand UO_1383 (O_1383,N_17039,N_17157);
or UO_1384 (O_1384,N_16352,N_18521);
nand UO_1385 (O_1385,N_16341,N_19858);
nand UO_1386 (O_1386,N_19526,N_18500);
nand UO_1387 (O_1387,N_19716,N_18111);
nor UO_1388 (O_1388,N_18575,N_17748);
nor UO_1389 (O_1389,N_16110,N_17137);
xor UO_1390 (O_1390,N_18008,N_18731);
xor UO_1391 (O_1391,N_17689,N_17991);
or UO_1392 (O_1392,N_16400,N_17546);
and UO_1393 (O_1393,N_19813,N_16367);
or UO_1394 (O_1394,N_18154,N_17053);
nor UO_1395 (O_1395,N_19919,N_19774);
nand UO_1396 (O_1396,N_19681,N_19465);
xor UO_1397 (O_1397,N_17269,N_18139);
and UO_1398 (O_1398,N_16002,N_17960);
xnor UO_1399 (O_1399,N_16990,N_19477);
or UO_1400 (O_1400,N_19828,N_18526);
and UO_1401 (O_1401,N_19936,N_18566);
or UO_1402 (O_1402,N_17678,N_16958);
or UO_1403 (O_1403,N_16674,N_16053);
nor UO_1404 (O_1404,N_17447,N_17341);
nor UO_1405 (O_1405,N_18384,N_19428);
and UO_1406 (O_1406,N_19725,N_18546);
or UO_1407 (O_1407,N_16282,N_16406);
nor UO_1408 (O_1408,N_19040,N_17051);
nor UO_1409 (O_1409,N_18763,N_18176);
and UO_1410 (O_1410,N_18266,N_18796);
and UO_1411 (O_1411,N_18780,N_17382);
nand UO_1412 (O_1412,N_18553,N_19575);
nor UO_1413 (O_1413,N_16547,N_16583);
nor UO_1414 (O_1414,N_16435,N_19166);
nor UO_1415 (O_1415,N_19501,N_19869);
and UO_1416 (O_1416,N_19478,N_18902);
nand UO_1417 (O_1417,N_16030,N_17584);
and UO_1418 (O_1418,N_17006,N_16153);
xnor UO_1419 (O_1419,N_19822,N_18609);
xnor UO_1420 (O_1420,N_17317,N_18075);
or UO_1421 (O_1421,N_18968,N_17904);
nand UO_1422 (O_1422,N_17838,N_19112);
xor UO_1423 (O_1423,N_16542,N_16654);
and UO_1424 (O_1424,N_19514,N_16515);
nand UO_1425 (O_1425,N_16192,N_18049);
nor UO_1426 (O_1426,N_16676,N_16796);
nor UO_1427 (O_1427,N_17458,N_19131);
xor UO_1428 (O_1428,N_17428,N_17276);
nor UO_1429 (O_1429,N_17234,N_16802);
nand UO_1430 (O_1430,N_19799,N_16727);
and UO_1431 (O_1431,N_18031,N_16776);
nand UO_1432 (O_1432,N_17768,N_17119);
or UO_1433 (O_1433,N_16787,N_18386);
xor UO_1434 (O_1434,N_17023,N_16267);
xnor UO_1435 (O_1435,N_19525,N_17886);
and UO_1436 (O_1436,N_18861,N_17983);
nand UO_1437 (O_1437,N_16753,N_19610);
or UO_1438 (O_1438,N_18294,N_19430);
or UO_1439 (O_1439,N_18823,N_17201);
nand UO_1440 (O_1440,N_18844,N_16006);
and UO_1441 (O_1441,N_19264,N_18015);
and UO_1442 (O_1442,N_17298,N_17529);
xnor UO_1443 (O_1443,N_18179,N_18834);
nand UO_1444 (O_1444,N_18097,N_19633);
xor UO_1445 (O_1445,N_19944,N_17630);
nand UO_1446 (O_1446,N_18109,N_16530);
and UO_1447 (O_1447,N_16952,N_16634);
or UO_1448 (O_1448,N_19341,N_19708);
nor UO_1449 (O_1449,N_18439,N_17112);
nand UO_1450 (O_1450,N_17975,N_17054);
or UO_1451 (O_1451,N_17250,N_16278);
nand UO_1452 (O_1452,N_16348,N_19585);
and UO_1453 (O_1453,N_16827,N_17557);
and UO_1454 (O_1454,N_19102,N_17321);
and UO_1455 (O_1455,N_17057,N_17010);
or UO_1456 (O_1456,N_18535,N_17185);
or UO_1457 (O_1457,N_18239,N_17444);
and UO_1458 (O_1458,N_19638,N_19859);
nor UO_1459 (O_1459,N_17972,N_16548);
xor UO_1460 (O_1460,N_19063,N_16177);
xnor UO_1461 (O_1461,N_18135,N_17178);
nor UO_1462 (O_1462,N_16872,N_17915);
or UO_1463 (O_1463,N_16102,N_17275);
nor UO_1464 (O_1464,N_18217,N_18664);
or UO_1465 (O_1465,N_16765,N_16735);
nor UO_1466 (O_1466,N_17553,N_19860);
or UO_1467 (O_1467,N_18368,N_19669);
nor UO_1468 (O_1468,N_19108,N_18039);
nor UO_1469 (O_1469,N_19170,N_19351);
or UO_1470 (O_1470,N_19055,N_17101);
nor UO_1471 (O_1471,N_17728,N_16108);
xor UO_1472 (O_1472,N_16236,N_19339);
and UO_1473 (O_1473,N_17522,N_17351);
nor UO_1474 (O_1474,N_16084,N_17750);
or UO_1475 (O_1475,N_19802,N_18704);
or UO_1476 (O_1476,N_16812,N_16283);
or UO_1477 (O_1477,N_16186,N_17822);
nand UO_1478 (O_1478,N_17489,N_18005);
and UO_1479 (O_1479,N_16048,N_18670);
nor UO_1480 (O_1480,N_16821,N_18515);
and UO_1481 (O_1481,N_16097,N_17538);
or UO_1482 (O_1482,N_16428,N_16127);
nand UO_1483 (O_1483,N_16856,N_19426);
nand UO_1484 (O_1484,N_17759,N_16064);
or UO_1485 (O_1485,N_16715,N_17501);
nand UO_1486 (O_1486,N_18702,N_18908);
nor UO_1487 (O_1487,N_16964,N_16298);
or UO_1488 (O_1488,N_17671,N_18662);
nand UO_1489 (O_1489,N_16005,N_18347);
nand UO_1490 (O_1490,N_18693,N_17440);
nor UO_1491 (O_1491,N_18138,N_16122);
or UO_1492 (O_1492,N_19688,N_19934);
and UO_1493 (O_1493,N_16119,N_18938);
nand UO_1494 (O_1494,N_17620,N_18480);
nor UO_1495 (O_1495,N_18004,N_17918);
nand UO_1496 (O_1496,N_18585,N_17105);
nand UO_1497 (O_1497,N_16413,N_18447);
nand UO_1498 (O_1498,N_17683,N_16363);
nand UO_1499 (O_1499,N_18313,N_18072);
and UO_1500 (O_1500,N_17334,N_16452);
nand UO_1501 (O_1501,N_18056,N_16580);
nor UO_1502 (O_1502,N_17845,N_16781);
or UO_1503 (O_1503,N_16304,N_19548);
and UO_1504 (O_1504,N_17641,N_18555);
nand UO_1505 (O_1505,N_18683,N_17133);
or UO_1506 (O_1506,N_19721,N_16522);
nor UO_1507 (O_1507,N_18216,N_16773);
xor UO_1508 (O_1508,N_16141,N_17813);
or UO_1509 (O_1509,N_17182,N_16806);
nand UO_1510 (O_1510,N_18430,N_16562);
or UO_1511 (O_1511,N_16554,N_18308);
and UO_1512 (O_1512,N_16505,N_18076);
and UO_1513 (O_1513,N_18493,N_19099);
nand UO_1514 (O_1514,N_17331,N_18063);
nor UO_1515 (O_1515,N_19648,N_17624);
and UO_1516 (O_1516,N_17483,N_19423);
nand UO_1517 (O_1517,N_18444,N_16926);
nor UO_1518 (O_1518,N_18499,N_16722);
or UO_1519 (O_1519,N_19021,N_16307);
or UO_1520 (O_1520,N_19679,N_16913);
xnor UO_1521 (O_1521,N_19026,N_17188);
xnor UO_1522 (O_1522,N_16618,N_16768);
nor UO_1523 (O_1523,N_17408,N_16747);
xnor UO_1524 (O_1524,N_17223,N_18473);
and UO_1525 (O_1525,N_18083,N_19053);
xnor UO_1526 (O_1526,N_18442,N_16226);
nand UO_1527 (O_1527,N_19460,N_18129);
or UO_1528 (O_1528,N_18790,N_17184);
xor UO_1529 (O_1529,N_19549,N_19204);
and UO_1530 (O_1530,N_17685,N_17205);
nand UO_1531 (O_1531,N_17031,N_19915);
xor UO_1532 (O_1532,N_19235,N_19546);
nor UO_1533 (O_1533,N_17730,N_18504);
and UO_1534 (O_1534,N_17171,N_19414);
nand UO_1535 (O_1535,N_19628,N_17214);
nor UO_1536 (O_1536,N_19946,N_18574);
nor UO_1537 (O_1537,N_18423,N_18115);
nor UO_1538 (O_1538,N_18619,N_17220);
nor UO_1539 (O_1539,N_19870,N_19512);
nand UO_1540 (O_1540,N_17695,N_18826);
or UO_1541 (O_1541,N_17527,N_17790);
or UO_1542 (O_1542,N_16472,N_16799);
nand UO_1543 (O_1543,N_18253,N_16214);
xor UO_1544 (O_1544,N_18328,N_19223);
nand UO_1545 (O_1545,N_19604,N_17189);
nand UO_1546 (O_1546,N_18736,N_19090);
nand UO_1547 (O_1547,N_16613,N_19468);
nand UO_1548 (O_1548,N_19580,N_18412);
nor UO_1549 (O_1549,N_19035,N_19962);
nand UO_1550 (O_1550,N_17040,N_19815);
and UO_1551 (O_1551,N_18457,N_18624);
nand UO_1552 (O_1552,N_17287,N_16533);
or UO_1553 (O_1553,N_17639,N_19369);
nor UO_1554 (O_1554,N_17385,N_19642);
and UO_1555 (O_1555,N_16793,N_18606);
nand UO_1556 (O_1556,N_16624,N_18045);
nor UO_1557 (O_1557,N_19775,N_19380);
nor UO_1558 (O_1558,N_18611,N_18806);
nor UO_1559 (O_1559,N_19761,N_16597);
nand UO_1560 (O_1560,N_19550,N_18737);
and UO_1561 (O_1561,N_16737,N_16456);
nor UO_1562 (O_1562,N_17126,N_18374);
nand UO_1563 (O_1563,N_17474,N_19335);
and UO_1564 (O_1564,N_17038,N_17751);
xnor UO_1565 (O_1565,N_16779,N_19731);
nand UO_1566 (O_1566,N_16392,N_18690);
or UO_1567 (O_1567,N_19389,N_16473);
xor UO_1568 (O_1568,N_18660,N_18453);
nand UO_1569 (O_1569,N_17513,N_18178);
nand UO_1570 (O_1570,N_19075,N_17999);
or UO_1571 (O_1571,N_17681,N_18286);
xor UO_1572 (O_1572,N_17718,N_18053);
nor UO_1573 (O_1573,N_19088,N_16804);
xor UO_1574 (O_1574,N_16840,N_18534);
nand UO_1575 (O_1575,N_16012,N_16149);
xor UO_1576 (O_1576,N_16790,N_18672);
nor UO_1577 (O_1577,N_19506,N_18279);
or UO_1578 (O_1578,N_17982,N_17616);
and UO_1579 (O_1579,N_19475,N_16979);
nand UO_1580 (O_1580,N_18929,N_18544);
and UO_1581 (O_1581,N_19265,N_17978);
nand UO_1582 (O_1582,N_17786,N_16040);
or UO_1583 (O_1583,N_18394,N_19641);
nor UO_1584 (O_1584,N_18531,N_16578);
and UO_1585 (O_1585,N_19668,N_16496);
nor UO_1586 (O_1586,N_19592,N_19017);
nor UO_1587 (O_1587,N_18872,N_17069);
and UO_1588 (O_1588,N_18646,N_17923);
nand UO_1589 (O_1589,N_16693,N_16534);
nor UO_1590 (O_1590,N_19661,N_16037);
nand UO_1591 (O_1591,N_19001,N_19476);
or UO_1592 (O_1592,N_19398,N_19045);
nand UO_1593 (O_1593,N_17418,N_17407);
nand UO_1594 (O_1594,N_17607,N_18197);
nor UO_1595 (O_1595,N_16290,N_19051);
and UO_1596 (O_1596,N_17170,N_17648);
or UO_1597 (O_1597,N_19400,N_18065);
nand UO_1598 (O_1598,N_17111,N_16908);
nand UO_1599 (O_1599,N_19886,N_16874);
nor UO_1600 (O_1600,N_17204,N_19182);
xor UO_1601 (O_1601,N_16602,N_19171);
nor UO_1602 (O_1602,N_17560,N_16078);
and UO_1603 (O_1603,N_16377,N_17078);
and UO_1604 (O_1604,N_19800,N_19689);
nand UO_1605 (O_1605,N_17664,N_18194);
or UO_1606 (O_1606,N_18243,N_19070);
nand UO_1607 (O_1607,N_17514,N_19263);
and UO_1608 (O_1608,N_19094,N_16480);
nor UO_1609 (O_1609,N_16660,N_17631);
nor UO_1610 (O_1610,N_19987,N_17686);
nand UO_1611 (O_1611,N_16216,N_19422);
or UO_1612 (O_1612,N_16815,N_16268);
or UO_1613 (O_1613,N_17362,N_19715);
and UO_1614 (O_1614,N_19029,N_18042);
nand UO_1615 (O_1615,N_18722,N_18040);
nor UO_1616 (O_1616,N_18761,N_16100);
xor UO_1617 (O_1617,N_18697,N_18855);
and UO_1618 (O_1618,N_18359,N_18598);
nor UO_1619 (O_1619,N_17712,N_19312);
xnor UO_1620 (O_1620,N_17757,N_17469);
nand UO_1621 (O_1621,N_17122,N_16056);
nand UO_1622 (O_1622,N_19290,N_18278);
or UO_1623 (O_1623,N_16966,N_18519);
and UO_1624 (O_1624,N_16641,N_18033);
nor UO_1625 (O_1625,N_18675,N_16302);
nor UO_1626 (O_1626,N_18822,N_18708);
and UO_1627 (O_1627,N_19203,N_16620);
xor UO_1628 (O_1628,N_19529,N_19835);
nor UO_1629 (O_1629,N_19006,N_19371);
nand UO_1630 (O_1630,N_16698,N_18551);
nand UO_1631 (O_1631,N_18372,N_19994);
xnor UO_1632 (O_1632,N_18159,N_19195);
and UO_1633 (O_1633,N_18036,N_16334);
nor UO_1634 (O_1634,N_18963,N_17687);
and UO_1635 (O_1635,N_19173,N_18113);
or UO_1636 (O_1636,N_16680,N_19595);
nand UO_1637 (O_1637,N_19402,N_17480);
or UO_1638 (O_1638,N_17151,N_19127);
or UO_1639 (O_1639,N_17449,N_18303);
or UO_1640 (O_1640,N_18365,N_16243);
or UO_1641 (O_1641,N_16327,N_17709);
xor UO_1642 (O_1642,N_17373,N_19313);
xnor UO_1643 (O_1643,N_17159,N_16742);
nand UO_1644 (O_1644,N_16321,N_17935);
and UO_1645 (O_1645,N_17843,N_16599);
or UO_1646 (O_1646,N_18682,N_18231);
and UO_1647 (O_1647,N_16746,N_19917);
xnor UO_1648 (O_1648,N_16690,N_18346);
nand UO_1649 (O_1649,N_17511,N_18701);
and UO_1650 (O_1650,N_17792,N_17889);
nor UO_1651 (O_1651,N_19562,N_18339);
nor UO_1652 (O_1652,N_16247,N_16825);
or UO_1653 (O_1653,N_17260,N_18658);
or UO_1654 (O_1654,N_16625,N_19983);
xor UO_1655 (O_1655,N_16235,N_17438);
and UO_1656 (O_1656,N_18153,N_16914);
xnor UO_1657 (O_1657,N_18716,N_17992);
or UO_1658 (O_1658,N_19769,N_16754);
nand UO_1659 (O_1659,N_16046,N_17569);
and UO_1660 (O_1660,N_16457,N_17652);
nor UO_1661 (O_1661,N_16927,N_16616);
and UO_1662 (O_1662,N_19818,N_18891);
and UO_1663 (O_1663,N_16047,N_19608);
nor UO_1664 (O_1664,N_18895,N_19778);
nand UO_1665 (O_1665,N_17922,N_16104);
or UO_1666 (O_1666,N_17955,N_18666);
nand UO_1667 (O_1667,N_19198,N_16710);
xor UO_1668 (O_1668,N_16774,N_19598);
nand UO_1669 (O_1669,N_17156,N_18335);
nor UO_1670 (O_1670,N_16239,N_19153);
or UO_1671 (O_1671,N_19043,N_18986);
or UO_1672 (O_1672,N_19132,N_16968);
nand UO_1673 (O_1673,N_18964,N_16839);
xnor UO_1674 (O_1674,N_16351,N_16975);
nand UO_1675 (O_1675,N_19293,N_18464);
or UO_1676 (O_1676,N_19952,N_17286);
or UO_1677 (O_1677,N_16444,N_17369);
nor UO_1678 (O_1678,N_19683,N_18472);
or UO_1679 (O_1679,N_19139,N_17948);
nor UO_1680 (O_1680,N_18982,N_19450);
nor UO_1681 (O_1681,N_16950,N_18933);
or UO_1682 (O_1682,N_19165,N_16851);
nand UO_1683 (O_1683,N_19571,N_16893);
nand UO_1684 (O_1684,N_18744,N_18252);
and UO_1685 (O_1685,N_16431,N_17884);
or UO_1686 (O_1686,N_18333,N_16938);
or UO_1687 (O_1687,N_16280,N_19735);
nor UO_1688 (O_1688,N_18838,N_16898);
and UO_1689 (O_1689,N_16638,N_19382);
nand UO_1690 (O_1690,N_19973,N_19321);
xor UO_1691 (O_1691,N_17468,N_17979);
nor UO_1692 (O_1692,N_17688,N_19269);
or UO_1693 (O_1693,N_16495,N_17756);
and UO_1694 (O_1694,N_18230,N_19535);
and UO_1695 (O_1695,N_17226,N_18155);
nor UO_1696 (O_1696,N_19784,N_17401);
or UO_1697 (O_1697,N_17672,N_16114);
or UO_1698 (O_1698,N_18024,N_18470);
nand UO_1699 (O_1699,N_16740,N_17323);
and UO_1700 (O_1700,N_17874,N_16887);
nor UO_1701 (O_1701,N_19434,N_17386);
nor UO_1702 (O_1702,N_19047,N_18692);
nor UO_1703 (O_1703,N_18726,N_18007);
nand UO_1704 (O_1704,N_19902,N_18607);
or UO_1705 (O_1705,N_18483,N_19868);
and UO_1706 (O_1706,N_16073,N_17526);
nor UO_1707 (O_1707,N_16507,N_17599);
nand UO_1708 (O_1708,N_19399,N_18552);
xnor UO_1709 (O_1709,N_19454,N_17013);
xnor UO_1710 (O_1710,N_19327,N_16132);
or UO_1711 (O_1711,N_16852,N_18686);
and UO_1712 (O_1712,N_19442,N_16906);
and UO_1713 (O_1713,N_19782,N_19690);
nand UO_1714 (O_1714,N_19650,N_16861);
or UO_1715 (O_1715,N_18026,N_17087);
xor UO_1716 (O_1716,N_19181,N_16862);
or UO_1717 (O_1717,N_17848,N_18548);
nand UO_1718 (O_1718,N_16685,N_18201);
nor UO_1719 (O_1719,N_18866,N_16293);
nand UO_1720 (O_1720,N_18577,N_16857);
and UO_1721 (O_1721,N_19013,N_19620);
and UO_1722 (O_1722,N_16120,N_17397);
and UO_1723 (O_1723,N_17043,N_17798);
xnor UO_1724 (O_1724,N_19038,N_16512);
and UO_1725 (O_1725,N_16531,N_16558);
nor UO_1726 (O_1726,N_19305,N_17436);
or UO_1727 (O_1727,N_17088,N_17773);
or UO_1728 (O_1728,N_18388,N_19320);
nand UO_1729 (O_1729,N_18034,N_16217);
xnor UO_1730 (O_1730,N_18882,N_18016);
and UO_1731 (O_1731,N_17598,N_17274);
nand UO_1732 (O_1732,N_19101,N_19829);
and UO_1733 (O_1733,N_19345,N_17532);
nor UO_1734 (O_1734,N_18691,N_18066);
nand UO_1735 (O_1735,N_18760,N_17422);
nor UO_1736 (O_1736,N_16223,N_18711);
and UO_1737 (O_1737,N_17076,N_19600);
and UO_1738 (O_1738,N_18944,N_18380);
nand UO_1739 (O_1739,N_17804,N_18094);
nand UO_1740 (O_1740,N_17933,N_17647);
and UO_1741 (O_1741,N_16770,N_18656);
nor UO_1742 (O_1742,N_19957,N_19386);
and UO_1743 (O_1743,N_16932,N_17868);
and UO_1744 (O_1744,N_16895,N_17503);
and UO_1745 (O_1745,N_18911,N_19975);
and UO_1746 (O_1746,N_18813,N_18213);
nand UO_1747 (O_1747,N_19401,N_16945);
nand UO_1748 (O_1748,N_18994,N_17816);
and UO_1749 (O_1749,N_16587,N_17777);
and UO_1750 (O_1750,N_16903,N_19034);
nand UO_1751 (O_1751,N_19095,N_18215);
and UO_1752 (O_1752,N_18403,N_19483);
nand UO_1753 (O_1753,N_18527,N_18723);
xor UO_1754 (O_1754,N_19206,N_16757);
nand UO_1755 (O_1755,N_16997,N_16748);
and UO_1756 (O_1756,N_18355,N_18421);
nor UO_1757 (O_1757,N_18900,N_18596);
nor UO_1758 (O_1758,N_17463,N_19833);
nor UO_1759 (O_1759,N_19748,N_19467);
nor UO_1760 (O_1760,N_17167,N_17017);
nor UO_1761 (O_1761,N_16567,N_17625);
nor UO_1762 (O_1762,N_17563,N_17996);
nor UO_1763 (O_1763,N_16409,N_18054);
xnor UO_1764 (O_1764,N_19122,N_18366);
or UO_1765 (O_1765,N_19736,N_18336);
xnor UO_1766 (O_1766,N_19803,N_16954);
nor UO_1767 (O_1767,N_17508,N_17911);
and UO_1768 (O_1768,N_17866,N_18067);
xnor UO_1769 (O_1769,N_17403,N_16026);
nor UO_1770 (O_1770,N_16093,N_16414);
nand UO_1771 (O_1771,N_17964,N_17476);
nand UO_1772 (O_1772,N_17770,N_19528);
nor UO_1773 (O_1773,N_17594,N_17696);
nor UO_1774 (O_1774,N_17387,N_17812);
and UO_1775 (O_1775,N_19126,N_18299);
nand UO_1776 (O_1776,N_16980,N_16538);
nand UO_1777 (O_1777,N_18391,N_16277);
and UO_1778 (O_1778,N_18471,N_16834);
nor UO_1779 (O_1779,N_16281,N_19000);
nand UO_1780 (O_1780,N_18183,N_17266);
nor UO_1781 (O_1781,N_16183,N_19956);
nor UO_1782 (O_1782,N_17012,N_17306);
or UO_1783 (O_1783,N_19252,N_17571);
and UO_1784 (O_1784,N_19796,N_17934);
nand UO_1785 (O_1785,N_19486,N_16188);
and UO_1786 (O_1786,N_17818,N_19923);
or UO_1787 (O_1787,N_16716,N_18560);
nand UO_1788 (O_1788,N_16951,N_18645);
nor UO_1789 (O_1789,N_17328,N_19481);
and UO_1790 (O_1790,N_18390,N_19482);
nor UO_1791 (O_1791,N_19862,N_18684);
and UO_1792 (O_1792,N_18542,N_16970);
xnor UO_1793 (O_1793,N_19557,N_17442);
nor UO_1794 (O_1794,N_18382,N_16193);
nor UO_1795 (O_1795,N_18028,N_16835);
and UO_1796 (O_1796,N_17697,N_17290);
nand UO_1797 (O_1797,N_17519,N_16605);
or UO_1798 (O_1798,N_17753,N_16876);
nand UO_1799 (O_1799,N_19885,N_19793);
nand UO_1800 (O_1800,N_17776,N_17781);
nand UO_1801 (O_1801,N_19151,N_19926);
or UO_1802 (O_1802,N_17966,N_16853);
and UO_1803 (O_1803,N_18073,N_16045);
nor UO_1804 (O_1804,N_19794,N_17875);
and UO_1805 (O_1805,N_18445,N_16944);
or UO_1806 (O_1806,N_19958,N_16058);
and UO_1807 (O_1807,N_17578,N_17473);
or UO_1808 (O_1808,N_17192,N_19564);
nor UO_1809 (O_1809,N_19874,N_17634);
and UO_1810 (O_1810,N_18092,N_19435);
and UO_1811 (O_1811,N_16537,N_18120);
or UO_1812 (O_1812,N_16960,N_16785);
nand UO_1813 (O_1813,N_18643,N_17570);
and UO_1814 (O_1814,N_18455,N_17901);
nor UO_1815 (O_1815,N_19972,N_17490);
or UO_1816 (O_1816,N_19846,N_19880);
nand UO_1817 (O_1817,N_16869,N_17802);
or UO_1818 (O_1818,N_17655,N_19531);
nand UO_1819 (O_1819,N_17542,N_17360);
or UO_1820 (O_1820,N_16224,N_17906);
or UO_1821 (O_1821,N_17072,N_18401);
nand UO_1822 (O_1822,N_17358,N_18078);
nand UO_1823 (O_1823,N_16657,N_18363);
nand UO_1824 (O_1824,N_17046,N_18417);
nand UO_1825 (O_1825,N_18530,N_16894);
nor UO_1826 (O_1826,N_18818,N_17453);
xor UO_1827 (O_1827,N_16652,N_19147);
xor UO_1828 (O_1828,N_18794,N_19791);
nand UO_1829 (O_1829,N_19932,N_17497);
nand UO_1830 (O_1830,N_16317,N_17958);
nand UO_1831 (O_1831,N_19356,N_17521);
nand UO_1832 (O_1832,N_19059,N_17460);
or UO_1833 (O_1833,N_17603,N_18061);
and UO_1834 (O_1834,N_18949,N_18749);
nor UO_1835 (O_1835,N_16401,N_17257);
or UO_1836 (O_1836,N_19484,N_16069);
nor UO_1837 (O_1837,N_18889,N_19154);
and UO_1838 (O_1838,N_18828,N_17673);
nor UO_1839 (O_1839,N_17074,N_19229);
or UO_1840 (O_1840,N_17203,N_19298);
nor UO_1841 (O_1841,N_19238,N_19545);
or UO_1842 (O_1842,N_18810,N_16082);
and UO_1843 (O_1843,N_18603,N_17608);
or UO_1844 (O_1844,N_16969,N_17326);
or UO_1845 (O_1845,N_17847,N_19953);
or UO_1846 (O_1846,N_19908,N_16343);
and UO_1847 (O_1847,N_18014,N_18811);
nand UO_1848 (O_1848,N_16670,N_19123);
nand UO_1849 (O_1849,N_19663,N_19328);
or UO_1850 (O_1850,N_16726,N_18254);
xor UO_1851 (O_1851,N_18557,N_19453);
xor UO_1852 (O_1852,N_18549,N_17871);
nor UO_1853 (O_1853,N_19786,N_17890);
nor UO_1854 (O_1854,N_18200,N_19867);
nand UO_1855 (O_1855,N_17293,N_17312);
nand UO_1856 (O_1856,N_16203,N_17262);
or UO_1857 (O_1857,N_18079,N_18334);
xor UO_1858 (O_1858,N_19079,N_18284);
or UO_1859 (O_1859,N_17466,N_17676);
nand UO_1860 (O_1860,N_18732,N_16111);
xnor UO_1861 (O_1861,N_16029,N_17646);
nor UO_1862 (O_1862,N_18084,N_18290);
nand UO_1863 (O_1863,N_16323,N_17415);
nor UO_1864 (O_1864,N_18909,N_18913);
nand UO_1865 (O_1865,N_18452,N_18556);
nand UO_1866 (O_1866,N_17502,N_16640);
or UO_1867 (O_1867,N_19393,N_19583);
or UO_1868 (O_1868,N_18681,N_19757);
nand UO_1869 (O_1869,N_17065,N_18395);
and UO_1870 (O_1870,N_16902,N_19338);
xor UO_1871 (O_1871,N_17372,N_17187);
nand UO_1872 (O_1872,N_19760,N_16596);
nor UO_1873 (O_1873,N_16503,N_17582);
and UO_1874 (O_1874,N_16417,N_17969);
or UO_1875 (O_1875,N_19068,N_19888);
nor UO_1876 (O_1876,N_16783,N_16519);
nand UO_1877 (O_1877,N_16060,N_18988);
or UO_1878 (O_1878,N_17425,N_17788);
and UO_1879 (O_1879,N_17805,N_18437);
xnor UO_1880 (O_1880,N_17809,N_18110);
or UO_1881 (O_1881,N_19553,N_17004);
and UO_1882 (O_1882,N_18819,N_16909);
nand UO_1883 (O_1883,N_16453,N_18789);
nor UO_1884 (O_1884,N_16571,N_19841);
nor UO_1885 (O_1885,N_19018,N_18756);
nand UO_1886 (O_1886,N_16513,N_18512);
nand UO_1887 (O_1887,N_19316,N_17684);
and UO_1888 (O_1888,N_16550,N_19745);
nor UO_1889 (O_1889,N_16467,N_16789);
or UO_1890 (O_1890,N_19906,N_18268);
or UO_1891 (O_1891,N_18820,N_17354);
nand UO_1892 (O_1892,N_17191,N_19821);
and UO_1893 (O_1893,N_19738,N_18734);
and UO_1894 (O_1894,N_18064,N_18010);
or UO_1895 (O_1895,N_18529,N_18758);
and UO_1896 (O_1896,N_19076,N_18148);
nor UO_1897 (O_1897,N_18970,N_18371);
nor UO_1898 (O_1898,N_17833,N_17255);
or UO_1899 (O_1899,N_18979,N_16899);
nand UO_1900 (O_1900,N_19078,N_17917);
nor UO_1901 (O_1901,N_17477,N_18926);
xnor UO_1902 (O_1902,N_19709,N_18288);
or UO_1903 (O_1903,N_16175,N_19726);
and UO_1904 (O_1904,N_19606,N_17778);
nand UO_1905 (O_1905,N_18868,N_16463);
and UO_1906 (O_1906,N_18738,N_16629);
or UO_1907 (O_1907,N_18407,N_17821);
and UO_1908 (O_1908,N_17296,N_18580);
xnor UO_1909 (O_1909,N_18700,N_18331);
nand UO_1910 (O_1910,N_16955,N_18998);
nand UO_1911 (O_1911,N_19855,N_18204);
and UO_1912 (O_1912,N_17259,N_19387);
or UO_1913 (O_1913,N_18121,N_16166);
and UO_1914 (O_1914,N_18319,N_17558);
or UO_1915 (O_1915,N_18419,N_18285);
and UO_1916 (O_1916,N_19376,N_16755);
nor UO_1917 (O_1917,N_19019,N_17531);
or UO_1918 (O_1918,N_16607,N_18525);
nor UO_1919 (O_1919,N_16831,N_18301);
xnor UO_1920 (O_1920,N_17008,N_19507);
and UO_1921 (O_1921,N_18849,N_16498);
nor UO_1922 (O_1922,N_19810,N_17411);
or UO_1923 (O_1923,N_18942,N_18295);
and UO_1924 (O_1924,N_19569,N_19383);
or UO_1925 (O_1925,N_19192,N_18427);
nor UO_1926 (O_1926,N_19797,N_17597);
nand UO_1927 (O_1927,N_19493,N_18102);
or UO_1928 (O_1928,N_17315,N_16375);
nand UO_1929 (O_1929,N_19225,N_17840);
or UO_1930 (O_1930,N_16408,N_18543);
nor UO_1931 (O_1931,N_18244,N_16461);
and UO_1932 (O_1932,N_17938,N_18426);
and UO_1933 (O_1933,N_17791,N_18885);
or UO_1934 (O_1934,N_19753,N_16172);
and UO_1935 (O_1935,N_19014,N_18973);
or UO_1936 (O_1936,N_18568,N_16162);
or UO_1937 (O_1937,N_17484,N_17343);
xor UO_1938 (O_1938,N_18240,N_17454);
nand UO_1939 (O_1939,N_16150,N_19660);
xor UO_1940 (O_1940,N_18156,N_18245);
xnor UO_1941 (O_1941,N_16460,N_18060);
or UO_1942 (O_1942,N_18134,N_16619);
nand UO_1943 (O_1943,N_19891,N_17131);
nor UO_1944 (O_1944,N_17857,N_18379);
nor UO_1945 (O_1945,N_19904,N_17534);
nor UO_1946 (O_1946,N_16988,N_16633);
or UO_1947 (O_1947,N_16760,N_16425);
xnor UO_1948 (O_1948,N_16590,N_19990);
xor UO_1949 (O_1949,N_17163,N_19344);
nand UO_1950 (O_1950,N_19509,N_18479);
or UO_1951 (O_1951,N_18622,N_19406);
and UO_1952 (O_1952,N_19337,N_19048);
or UO_1953 (O_1953,N_19746,N_16008);
and UO_1954 (O_1954,N_19941,N_19933);
or UO_1955 (O_1955,N_17762,N_18375);
and UO_1956 (O_1956,N_16867,N_18062);
or UO_1957 (O_1957,N_19522,N_16598);
and UO_1958 (O_1958,N_17981,N_17708);
or UO_1959 (O_1959,N_17325,N_19897);
and UO_1960 (O_1960,N_18100,N_19449);
and UO_1961 (O_1961,N_18617,N_16731);
or UO_1962 (O_1962,N_18310,N_19911);
and UO_1963 (O_1963,N_16879,N_18399);
and UO_1964 (O_1964,N_17003,N_19378);
nor UO_1965 (O_1965,N_16798,N_18733);
and UO_1966 (O_1966,N_18396,N_17963);
and UO_1967 (O_1967,N_19942,N_17456);
nand UO_1968 (O_1968,N_19985,N_19652);
nand UO_1969 (O_1969,N_19066,N_18488);
nor UO_1970 (O_1970,N_17883,N_16374);
or UO_1971 (O_1971,N_19686,N_16963);
nand UO_1972 (O_1972,N_18669,N_19232);
nand UO_1973 (O_1973,N_18324,N_17887);
nor UO_1974 (O_1974,N_16240,N_17807);
nand UO_1975 (O_1975,N_17618,N_17064);
nand UO_1976 (O_1976,N_18879,N_17627);
or UO_1977 (O_1977,N_16949,N_18863);
xnor UO_1978 (O_1978,N_16285,N_19455);
nand UO_1979 (O_1979,N_16989,N_17638);
nand UO_1980 (O_1980,N_16661,N_16762);
or UO_1981 (O_1981,N_17450,N_17083);
xnor UO_1982 (O_1982,N_18212,N_17281);
xor UO_1983 (O_1983,N_18232,N_18269);
and UO_1984 (O_1984,N_18080,N_16749);
or UO_1985 (O_1985,N_16404,N_17175);
and UO_1986 (O_1986,N_17803,N_18106);
nand UO_1987 (O_1987,N_16585,N_18829);
xor UO_1988 (O_1988,N_16022,N_19299);
nor UO_1989 (O_1989,N_19644,N_16527);
nand UO_1990 (O_1990,N_16477,N_16269);
xnor UO_1991 (O_1991,N_18171,N_17729);
xor UO_1992 (O_1992,N_16508,N_19354);
and UO_1993 (O_1993,N_18287,N_18517);
nand UO_1994 (O_1994,N_16061,N_19025);
nor UO_1995 (O_1995,N_19706,N_16206);
or UO_1996 (O_1996,N_17591,N_17036);
or UO_1997 (O_1997,N_18298,N_18428);
nand UO_1998 (O_1998,N_16139,N_16196);
and UO_1999 (O_1999,N_19403,N_18797);
and UO_2000 (O_2000,N_16796,N_17303);
nand UO_2001 (O_2001,N_19618,N_17384);
nand UO_2002 (O_2002,N_19205,N_17249);
nand UO_2003 (O_2003,N_19265,N_19906);
or UO_2004 (O_2004,N_19894,N_19202);
nor UO_2005 (O_2005,N_18676,N_18041);
and UO_2006 (O_2006,N_18510,N_16312);
nand UO_2007 (O_2007,N_19841,N_19827);
or UO_2008 (O_2008,N_19813,N_17450);
nor UO_2009 (O_2009,N_16941,N_16299);
nand UO_2010 (O_2010,N_17390,N_16644);
nand UO_2011 (O_2011,N_16382,N_19509);
xor UO_2012 (O_2012,N_18045,N_16826);
xor UO_2013 (O_2013,N_18437,N_19670);
nand UO_2014 (O_2014,N_18386,N_18443);
and UO_2015 (O_2015,N_17870,N_18523);
and UO_2016 (O_2016,N_17028,N_19650);
xor UO_2017 (O_2017,N_18983,N_17248);
and UO_2018 (O_2018,N_17963,N_17713);
or UO_2019 (O_2019,N_17533,N_19443);
xnor UO_2020 (O_2020,N_16565,N_19350);
nor UO_2021 (O_2021,N_19293,N_19221);
and UO_2022 (O_2022,N_17591,N_17861);
and UO_2023 (O_2023,N_18254,N_18966);
nand UO_2024 (O_2024,N_17669,N_17040);
and UO_2025 (O_2025,N_17321,N_19973);
nand UO_2026 (O_2026,N_18012,N_18161);
nor UO_2027 (O_2027,N_19077,N_17966);
xnor UO_2028 (O_2028,N_16213,N_18943);
and UO_2029 (O_2029,N_16743,N_16403);
and UO_2030 (O_2030,N_19912,N_18661);
nand UO_2031 (O_2031,N_17691,N_18038);
nand UO_2032 (O_2032,N_16668,N_19706);
or UO_2033 (O_2033,N_18751,N_19481);
nor UO_2034 (O_2034,N_16206,N_18947);
and UO_2035 (O_2035,N_16827,N_19273);
nand UO_2036 (O_2036,N_18256,N_18751);
nand UO_2037 (O_2037,N_18503,N_18472);
nand UO_2038 (O_2038,N_16407,N_16380);
nor UO_2039 (O_2039,N_19851,N_18428);
or UO_2040 (O_2040,N_19903,N_16841);
nand UO_2041 (O_2041,N_17744,N_17600);
nor UO_2042 (O_2042,N_18091,N_19167);
nor UO_2043 (O_2043,N_17050,N_17807);
nand UO_2044 (O_2044,N_18296,N_18756);
nor UO_2045 (O_2045,N_18594,N_16149);
or UO_2046 (O_2046,N_19162,N_18473);
or UO_2047 (O_2047,N_19710,N_16528);
and UO_2048 (O_2048,N_17991,N_17881);
nand UO_2049 (O_2049,N_16655,N_19007);
nand UO_2050 (O_2050,N_19841,N_16954);
nand UO_2051 (O_2051,N_16804,N_19259);
or UO_2052 (O_2052,N_19864,N_18859);
or UO_2053 (O_2053,N_18136,N_19772);
nand UO_2054 (O_2054,N_16874,N_18408);
nor UO_2055 (O_2055,N_18170,N_16062);
nor UO_2056 (O_2056,N_19917,N_16206);
nor UO_2057 (O_2057,N_16315,N_16394);
nand UO_2058 (O_2058,N_18044,N_18861);
and UO_2059 (O_2059,N_17442,N_19027);
and UO_2060 (O_2060,N_19726,N_18066);
nand UO_2061 (O_2061,N_16205,N_16160);
nand UO_2062 (O_2062,N_16225,N_19303);
xor UO_2063 (O_2063,N_19639,N_16509);
or UO_2064 (O_2064,N_17674,N_19329);
or UO_2065 (O_2065,N_19209,N_16454);
or UO_2066 (O_2066,N_17107,N_17206);
nand UO_2067 (O_2067,N_19546,N_18689);
nand UO_2068 (O_2068,N_17393,N_19779);
nor UO_2069 (O_2069,N_17890,N_17078);
nor UO_2070 (O_2070,N_18419,N_16123);
nand UO_2071 (O_2071,N_17194,N_18237);
and UO_2072 (O_2072,N_19565,N_18061);
nand UO_2073 (O_2073,N_16947,N_17609);
nand UO_2074 (O_2074,N_18236,N_17931);
and UO_2075 (O_2075,N_16951,N_19312);
nor UO_2076 (O_2076,N_19199,N_16564);
or UO_2077 (O_2077,N_18676,N_19076);
nor UO_2078 (O_2078,N_17097,N_19651);
xnor UO_2079 (O_2079,N_19704,N_19932);
and UO_2080 (O_2080,N_16627,N_18319);
nor UO_2081 (O_2081,N_16558,N_16173);
nor UO_2082 (O_2082,N_16096,N_17268);
nor UO_2083 (O_2083,N_17400,N_17035);
or UO_2084 (O_2084,N_17053,N_17576);
nand UO_2085 (O_2085,N_16505,N_18061);
nor UO_2086 (O_2086,N_18598,N_18978);
or UO_2087 (O_2087,N_19745,N_16693);
nor UO_2088 (O_2088,N_16169,N_18241);
nand UO_2089 (O_2089,N_19496,N_18867);
nand UO_2090 (O_2090,N_17316,N_16319);
and UO_2091 (O_2091,N_17528,N_17010);
and UO_2092 (O_2092,N_17351,N_19423);
and UO_2093 (O_2093,N_17866,N_18823);
nand UO_2094 (O_2094,N_16974,N_18069);
nand UO_2095 (O_2095,N_19549,N_16264);
nor UO_2096 (O_2096,N_17502,N_17324);
nor UO_2097 (O_2097,N_19021,N_19849);
nand UO_2098 (O_2098,N_18046,N_18446);
or UO_2099 (O_2099,N_16640,N_19698);
nand UO_2100 (O_2100,N_19241,N_18419);
and UO_2101 (O_2101,N_19678,N_18508);
nand UO_2102 (O_2102,N_18065,N_16857);
or UO_2103 (O_2103,N_17320,N_17703);
or UO_2104 (O_2104,N_18348,N_16661);
nor UO_2105 (O_2105,N_17700,N_17204);
nand UO_2106 (O_2106,N_18633,N_18097);
and UO_2107 (O_2107,N_19893,N_16474);
nand UO_2108 (O_2108,N_18808,N_16470);
and UO_2109 (O_2109,N_17450,N_16743);
xnor UO_2110 (O_2110,N_16792,N_16176);
or UO_2111 (O_2111,N_18958,N_19538);
or UO_2112 (O_2112,N_16277,N_18348);
or UO_2113 (O_2113,N_17327,N_16444);
or UO_2114 (O_2114,N_18300,N_18890);
nand UO_2115 (O_2115,N_19030,N_17802);
and UO_2116 (O_2116,N_18493,N_17960);
or UO_2117 (O_2117,N_17019,N_19769);
nor UO_2118 (O_2118,N_17054,N_18152);
nor UO_2119 (O_2119,N_16465,N_17589);
nand UO_2120 (O_2120,N_17574,N_17600);
or UO_2121 (O_2121,N_18750,N_17537);
nand UO_2122 (O_2122,N_19211,N_16594);
and UO_2123 (O_2123,N_19592,N_17245);
or UO_2124 (O_2124,N_18186,N_18283);
xnor UO_2125 (O_2125,N_19711,N_18695);
or UO_2126 (O_2126,N_19318,N_18483);
or UO_2127 (O_2127,N_18211,N_18659);
nor UO_2128 (O_2128,N_17840,N_18788);
xor UO_2129 (O_2129,N_19871,N_19951);
nor UO_2130 (O_2130,N_17279,N_18938);
or UO_2131 (O_2131,N_19109,N_17780);
nor UO_2132 (O_2132,N_16995,N_18328);
nand UO_2133 (O_2133,N_19278,N_19005);
and UO_2134 (O_2134,N_19767,N_18416);
nand UO_2135 (O_2135,N_19178,N_19824);
xor UO_2136 (O_2136,N_17857,N_18401);
nor UO_2137 (O_2137,N_16836,N_19129);
nor UO_2138 (O_2138,N_17754,N_16271);
xor UO_2139 (O_2139,N_19894,N_17212);
nor UO_2140 (O_2140,N_16085,N_19175);
or UO_2141 (O_2141,N_17676,N_18957);
nand UO_2142 (O_2142,N_16100,N_17578);
xor UO_2143 (O_2143,N_17771,N_17430);
and UO_2144 (O_2144,N_18405,N_17916);
nor UO_2145 (O_2145,N_17168,N_19480);
nand UO_2146 (O_2146,N_18092,N_17997);
nand UO_2147 (O_2147,N_16748,N_16471);
and UO_2148 (O_2148,N_17348,N_18469);
and UO_2149 (O_2149,N_17670,N_16083);
xor UO_2150 (O_2150,N_16849,N_17178);
xnor UO_2151 (O_2151,N_16334,N_16423);
and UO_2152 (O_2152,N_18939,N_19067);
and UO_2153 (O_2153,N_18288,N_17089);
nand UO_2154 (O_2154,N_16243,N_19535);
and UO_2155 (O_2155,N_17152,N_19010);
nand UO_2156 (O_2156,N_19719,N_19253);
and UO_2157 (O_2157,N_17471,N_19893);
nor UO_2158 (O_2158,N_17501,N_16321);
and UO_2159 (O_2159,N_18353,N_16454);
and UO_2160 (O_2160,N_19595,N_18207);
nor UO_2161 (O_2161,N_19159,N_18793);
nor UO_2162 (O_2162,N_17468,N_17750);
or UO_2163 (O_2163,N_16186,N_19788);
nand UO_2164 (O_2164,N_18053,N_19997);
or UO_2165 (O_2165,N_17697,N_17111);
nand UO_2166 (O_2166,N_16960,N_19740);
nor UO_2167 (O_2167,N_17665,N_17781);
nand UO_2168 (O_2168,N_19723,N_17205);
nor UO_2169 (O_2169,N_19147,N_18359);
and UO_2170 (O_2170,N_17757,N_19330);
xor UO_2171 (O_2171,N_19255,N_19534);
xnor UO_2172 (O_2172,N_19202,N_17365);
or UO_2173 (O_2173,N_19650,N_17124);
xnor UO_2174 (O_2174,N_19037,N_19642);
or UO_2175 (O_2175,N_18080,N_16442);
xnor UO_2176 (O_2176,N_17074,N_16728);
nand UO_2177 (O_2177,N_16111,N_17372);
nand UO_2178 (O_2178,N_18510,N_19909);
or UO_2179 (O_2179,N_17718,N_16672);
xor UO_2180 (O_2180,N_18963,N_18967);
or UO_2181 (O_2181,N_18511,N_18002);
or UO_2182 (O_2182,N_16484,N_18404);
nor UO_2183 (O_2183,N_16964,N_18513);
or UO_2184 (O_2184,N_19365,N_17460);
xor UO_2185 (O_2185,N_16259,N_18267);
nor UO_2186 (O_2186,N_17295,N_19086);
nand UO_2187 (O_2187,N_17525,N_19961);
nand UO_2188 (O_2188,N_16316,N_18208);
or UO_2189 (O_2189,N_19067,N_18049);
and UO_2190 (O_2190,N_18768,N_17531);
nand UO_2191 (O_2191,N_16249,N_16324);
nand UO_2192 (O_2192,N_19371,N_17675);
nand UO_2193 (O_2193,N_19788,N_18774);
nor UO_2194 (O_2194,N_16114,N_16956);
and UO_2195 (O_2195,N_19799,N_17805);
nor UO_2196 (O_2196,N_19098,N_18039);
nor UO_2197 (O_2197,N_16846,N_19474);
and UO_2198 (O_2198,N_18917,N_16902);
nand UO_2199 (O_2199,N_18658,N_17277);
nand UO_2200 (O_2200,N_19526,N_16408);
xnor UO_2201 (O_2201,N_19770,N_16669);
or UO_2202 (O_2202,N_16550,N_18531);
nand UO_2203 (O_2203,N_17796,N_18145);
nand UO_2204 (O_2204,N_19454,N_17205);
nor UO_2205 (O_2205,N_16373,N_16260);
and UO_2206 (O_2206,N_17069,N_18770);
and UO_2207 (O_2207,N_19072,N_18558);
nand UO_2208 (O_2208,N_19640,N_19375);
nand UO_2209 (O_2209,N_16759,N_19353);
nand UO_2210 (O_2210,N_17326,N_16683);
or UO_2211 (O_2211,N_19772,N_17069);
nor UO_2212 (O_2212,N_19621,N_18800);
and UO_2213 (O_2213,N_16949,N_17058);
nand UO_2214 (O_2214,N_18138,N_17722);
and UO_2215 (O_2215,N_16445,N_19933);
nor UO_2216 (O_2216,N_17004,N_18247);
or UO_2217 (O_2217,N_18408,N_17535);
and UO_2218 (O_2218,N_18914,N_19281);
and UO_2219 (O_2219,N_17387,N_16771);
and UO_2220 (O_2220,N_17616,N_16731);
or UO_2221 (O_2221,N_16542,N_17923);
nand UO_2222 (O_2222,N_16402,N_19027);
nor UO_2223 (O_2223,N_17670,N_18991);
and UO_2224 (O_2224,N_18757,N_18608);
and UO_2225 (O_2225,N_19222,N_18894);
nand UO_2226 (O_2226,N_18864,N_19118);
nor UO_2227 (O_2227,N_16494,N_18484);
or UO_2228 (O_2228,N_17446,N_19125);
or UO_2229 (O_2229,N_16678,N_16823);
xnor UO_2230 (O_2230,N_19175,N_19670);
nor UO_2231 (O_2231,N_18752,N_19827);
nor UO_2232 (O_2232,N_18933,N_18902);
nor UO_2233 (O_2233,N_18489,N_18832);
and UO_2234 (O_2234,N_18209,N_18418);
nand UO_2235 (O_2235,N_16200,N_16445);
nand UO_2236 (O_2236,N_17957,N_17432);
nor UO_2237 (O_2237,N_19278,N_16398);
nor UO_2238 (O_2238,N_17142,N_18709);
nand UO_2239 (O_2239,N_19567,N_19857);
xor UO_2240 (O_2240,N_17597,N_16118);
and UO_2241 (O_2241,N_16246,N_17455);
nor UO_2242 (O_2242,N_18871,N_18165);
and UO_2243 (O_2243,N_19636,N_16019);
xnor UO_2244 (O_2244,N_16744,N_18702);
and UO_2245 (O_2245,N_18915,N_17002);
or UO_2246 (O_2246,N_17828,N_18038);
nor UO_2247 (O_2247,N_16799,N_18373);
nand UO_2248 (O_2248,N_18297,N_18972);
nand UO_2249 (O_2249,N_17747,N_17150);
and UO_2250 (O_2250,N_18711,N_16733);
nand UO_2251 (O_2251,N_18069,N_17658);
and UO_2252 (O_2252,N_16376,N_18037);
nor UO_2253 (O_2253,N_16056,N_17465);
and UO_2254 (O_2254,N_19543,N_19751);
or UO_2255 (O_2255,N_17620,N_17649);
nand UO_2256 (O_2256,N_19462,N_17171);
nand UO_2257 (O_2257,N_19738,N_19355);
or UO_2258 (O_2258,N_18407,N_19635);
nand UO_2259 (O_2259,N_16986,N_19582);
nand UO_2260 (O_2260,N_19063,N_17895);
nand UO_2261 (O_2261,N_16510,N_17915);
and UO_2262 (O_2262,N_19725,N_19890);
or UO_2263 (O_2263,N_18262,N_18785);
nand UO_2264 (O_2264,N_17659,N_16096);
or UO_2265 (O_2265,N_18023,N_17139);
or UO_2266 (O_2266,N_17265,N_19777);
nand UO_2267 (O_2267,N_19157,N_19450);
or UO_2268 (O_2268,N_19667,N_19488);
nor UO_2269 (O_2269,N_18799,N_19312);
nand UO_2270 (O_2270,N_18304,N_17784);
and UO_2271 (O_2271,N_17621,N_19221);
xnor UO_2272 (O_2272,N_19333,N_17540);
or UO_2273 (O_2273,N_16962,N_18082);
xor UO_2274 (O_2274,N_17539,N_18076);
nand UO_2275 (O_2275,N_18500,N_17162);
and UO_2276 (O_2276,N_17120,N_16023);
or UO_2277 (O_2277,N_19393,N_19237);
nand UO_2278 (O_2278,N_16278,N_19570);
and UO_2279 (O_2279,N_19953,N_19661);
or UO_2280 (O_2280,N_19561,N_19913);
and UO_2281 (O_2281,N_16340,N_16130);
nand UO_2282 (O_2282,N_17164,N_16673);
nor UO_2283 (O_2283,N_19296,N_17161);
or UO_2284 (O_2284,N_19160,N_19961);
or UO_2285 (O_2285,N_18173,N_17165);
and UO_2286 (O_2286,N_18803,N_18087);
xor UO_2287 (O_2287,N_18003,N_17405);
or UO_2288 (O_2288,N_18412,N_18820);
nand UO_2289 (O_2289,N_17111,N_18916);
nor UO_2290 (O_2290,N_17703,N_19228);
and UO_2291 (O_2291,N_17032,N_17454);
and UO_2292 (O_2292,N_16662,N_16882);
nand UO_2293 (O_2293,N_18327,N_16129);
and UO_2294 (O_2294,N_19157,N_18303);
xnor UO_2295 (O_2295,N_18935,N_17888);
or UO_2296 (O_2296,N_16444,N_19850);
nand UO_2297 (O_2297,N_18347,N_19930);
nor UO_2298 (O_2298,N_19478,N_16752);
and UO_2299 (O_2299,N_17837,N_16366);
and UO_2300 (O_2300,N_16249,N_16532);
or UO_2301 (O_2301,N_17700,N_18423);
and UO_2302 (O_2302,N_18360,N_18216);
xor UO_2303 (O_2303,N_19591,N_16852);
or UO_2304 (O_2304,N_16512,N_19128);
nor UO_2305 (O_2305,N_19876,N_19723);
nand UO_2306 (O_2306,N_16519,N_17974);
nor UO_2307 (O_2307,N_16487,N_16254);
nand UO_2308 (O_2308,N_17715,N_18714);
nand UO_2309 (O_2309,N_17080,N_19705);
xor UO_2310 (O_2310,N_17339,N_18656);
or UO_2311 (O_2311,N_19610,N_17920);
nor UO_2312 (O_2312,N_19286,N_17504);
and UO_2313 (O_2313,N_16255,N_19166);
nand UO_2314 (O_2314,N_19601,N_18669);
or UO_2315 (O_2315,N_19343,N_18329);
xnor UO_2316 (O_2316,N_16460,N_18115);
and UO_2317 (O_2317,N_16552,N_18753);
nand UO_2318 (O_2318,N_17593,N_17262);
nand UO_2319 (O_2319,N_17460,N_19393);
nand UO_2320 (O_2320,N_17736,N_19217);
nand UO_2321 (O_2321,N_18370,N_19785);
or UO_2322 (O_2322,N_17990,N_18103);
and UO_2323 (O_2323,N_19783,N_19499);
and UO_2324 (O_2324,N_17591,N_17994);
and UO_2325 (O_2325,N_19534,N_19972);
nor UO_2326 (O_2326,N_18729,N_18453);
and UO_2327 (O_2327,N_17998,N_16135);
or UO_2328 (O_2328,N_16746,N_17265);
or UO_2329 (O_2329,N_19705,N_18809);
or UO_2330 (O_2330,N_18879,N_18558);
xnor UO_2331 (O_2331,N_18047,N_18942);
nand UO_2332 (O_2332,N_17531,N_19130);
nor UO_2333 (O_2333,N_17999,N_19266);
nor UO_2334 (O_2334,N_19540,N_18738);
or UO_2335 (O_2335,N_16356,N_19431);
nor UO_2336 (O_2336,N_19264,N_16422);
or UO_2337 (O_2337,N_18468,N_19821);
or UO_2338 (O_2338,N_17164,N_18504);
and UO_2339 (O_2339,N_18809,N_18636);
and UO_2340 (O_2340,N_17176,N_16739);
or UO_2341 (O_2341,N_19120,N_17257);
and UO_2342 (O_2342,N_16867,N_18822);
nand UO_2343 (O_2343,N_16750,N_18577);
nand UO_2344 (O_2344,N_19817,N_16158);
xnor UO_2345 (O_2345,N_17007,N_18271);
nor UO_2346 (O_2346,N_16988,N_18125);
and UO_2347 (O_2347,N_18685,N_19168);
nand UO_2348 (O_2348,N_19094,N_17304);
xnor UO_2349 (O_2349,N_18055,N_17103);
xnor UO_2350 (O_2350,N_17101,N_16189);
and UO_2351 (O_2351,N_16432,N_16109);
or UO_2352 (O_2352,N_17009,N_18185);
or UO_2353 (O_2353,N_17473,N_19766);
xor UO_2354 (O_2354,N_17101,N_19730);
nand UO_2355 (O_2355,N_18508,N_17911);
nor UO_2356 (O_2356,N_18255,N_18360);
nand UO_2357 (O_2357,N_16815,N_16589);
nor UO_2358 (O_2358,N_17358,N_18992);
nor UO_2359 (O_2359,N_17185,N_16526);
or UO_2360 (O_2360,N_16113,N_17313);
nor UO_2361 (O_2361,N_17491,N_17852);
or UO_2362 (O_2362,N_18663,N_19197);
and UO_2363 (O_2363,N_17927,N_18739);
and UO_2364 (O_2364,N_19681,N_18568);
or UO_2365 (O_2365,N_16954,N_16400);
nand UO_2366 (O_2366,N_18791,N_18350);
nor UO_2367 (O_2367,N_16385,N_18524);
nand UO_2368 (O_2368,N_17818,N_16965);
or UO_2369 (O_2369,N_16061,N_18502);
nand UO_2370 (O_2370,N_16806,N_17013);
or UO_2371 (O_2371,N_18143,N_17012);
or UO_2372 (O_2372,N_18924,N_17012);
nor UO_2373 (O_2373,N_17807,N_17953);
nor UO_2374 (O_2374,N_16319,N_17570);
nor UO_2375 (O_2375,N_17514,N_16541);
or UO_2376 (O_2376,N_16457,N_16028);
and UO_2377 (O_2377,N_18470,N_17225);
and UO_2378 (O_2378,N_19584,N_17784);
xor UO_2379 (O_2379,N_18227,N_19059);
and UO_2380 (O_2380,N_19402,N_18259);
xnor UO_2381 (O_2381,N_19892,N_17574);
nand UO_2382 (O_2382,N_17852,N_17893);
and UO_2383 (O_2383,N_18123,N_18161);
or UO_2384 (O_2384,N_16316,N_16097);
nand UO_2385 (O_2385,N_19403,N_16051);
and UO_2386 (O_2386,N_19365,N_17825);
nor UO_2387 (O_2387,N_18434,N_16434);
nor UO_2388 (O_2388,N_16395,N_17625);
nand UO_2389 (O_2389,N_19507,N_18388);
nand UO_2390 (O_2390,N_18958,N_17396);
or UO_2391 (O_2391,N_17932,N_16890);
nor UO_2392 (O_2392,N_17832,N_16487);
and UO_2393 (O_2393,N_17474,N_18291);
or UO_2394 (O_2394,N_17787,N_19411);
nand UO_2395 (O_2395,N_17073,N_18935);
and UO_2396 (O_2396,N_18433,N_18456);
nand UO_2397 (O_2397,N_17633,N_19393);
and UO_2398 (O_2398,N_16750,N_16148);
nor UO_2399 (O_2399,N_17231,N_19590);
or UO_2400 (O_2400,N_19853,N_19275);
or UO_2401 (O_2401,N_16792,N_16668);
and UO_2402 (O_2402,N_18600,N_18437);
and UO_2403 (O_2403,N_18676,N_16009);
nor UO_2404 (O_2404,N_19927,N_19443);
or UO_2405 (O_2405,N_19485,N_17077);
nand UO_2406 (O_2406,N_19295,N_17989);
or UO_2407 (O_2407,N_16081,N_18507);
or UO_2408 (O_2408,N_17376,N_19747);
xor UO_2409 (O_2409,N_19286,N_16823);
nand UO_2410 (O_2410,N_17312,N_17212);
and UO_2411 (O_2411,N_19691,N_19270);
or UO_2412 (O_2412,N_17157,N_18771);
or UO_2413 (O_2413,N_19811,N_18108);
or UO_2414 (O_2414,N_17726,N_18203);
xor UO_2415 (O_2415,N_17894,N_17502);
nor UO_2416 (O_2416,N_17755,N_17692);
nor UO_2417 (O_2417,N_16029,N_19042);
nor UO_2418 (O_2418,N_16968,N_19707);
and UO_2419 (O_2419,N_16548,N_18761);
nand UO_2420 (O_2420,N_16379,N_16355);
or UO_2421 (O_2421,N_17616,N_19446);
or UO_2422 (O_2422,N_16765,N_19156);
nand UO_2423 (O_2423,N_19029,N_18788);
nor UO_2424 (O_2424,N_18432,N_19868);
or UO_2425 (O_2425,N_18351,N_19109);
nand UO_2426 (O_2426,N_19189,N_18391);
nand UO_2427 (O_2427,N_19217,N_16895);
nand UO_2428 (O_2428,N_17588,N_17426);
xor UO_2429 (O_2429,N_18912,N_17623);
or UO_2430 (O_2430,N_17309,N_16748);
nor UO_2431 (O_2431,N_16663,N_16466);
nor UO_2432 (O_2432,N_18797,N_16881);
nor UO_2433 (O_2433,N_19574,N_17729);
and UO_2434 (O_2434,N_17152,N_17180);
and UO_2435 (O_2435,N_16868,N_19886);
nor UO_2436 (O_2436,N_17887,N_19562);
nand UO_2437 (O_2437,N_16716,N_17054);
xnor UO_2438 (O_2438,N_17777,N_18118);
nand UO_2439 (O_2439,N_18040,N_16378);
and UO_2440 (O_2440,N_16830,N_18840);
and UO_2441 (O_2441,N_16139,N_17862);
or UO_2442 (O_2442,N_18464,N_18652);
xnor UO_2443 (O_2443,N_18844,N_16221);
nand UO_2444 (O_2444,N_19377,N_16673);
nand UO_2445 (O_2445,N_17309,N_19715);
xnor UO_2446 (O_2446,N_18148,N_18152);
and UO_2447 (O_2447,N_17353,N_16334);
nor UO_2448 (O_2448,N_18513,N_19653);
nor UO_2449 (O_2449,N_18865,N_17132);
nand UO_2450 (O_2450,N_18796,N_17115);
nor UO_2451 (O_2451,N_17228,N_18327);
and UO_2452 (O_2452,N_16036,N_18212);
nand UO_2453 (O_2453,N_18545,N_16058);
or UO_2454 (O_2454,N_18436,N_19999);
or UO_2455 (O_2455,N_19244,N_19628);
and UO_2456 (O_2456,N_16847,N_19195);
and UO_2457 (O_2457,N_17876,N_17321);
nand UO_2458 (O_2458,N_18442,N_18621);
and UO_2459 (O_2459,N_16542,N_19396);
and UO_2460 (O_2460,N_17480,N_16939);
nor UO_2461 (O_2461,N_17777,N_16639);
or UO_2462 (O_2462,N_19337,N_19743);
nor UO_2463 (O_2463,N_16081,N_16167);
nor UO_2464 (O_2464,N_19279,N_17440);
nor UO_2465 (O_2465,N_16540,N_17619);
nand UO_2466 (O_2466,N_18618,N_19509);
nor UO_2467 (O_2467,N_18602,N_16848);
nor UO_2468 (O_2468,N_19896,N_18340);
or UO_2469 (O_2469,N_19412,N_19181);
nand UO_2470 (O_2470,N_18217,N_16695);
nand UO_2471 (O_2471,N_16398,N_18793);
nand UO_2472 (O_2472,N_18110,N_17354);
and UO_2473 (O_2473,N_16868,N_16245);
nor UO_2474 (O_2474,N_17086,N_19511);
xnor UO_2475 (O_2475,N_17989,N_18964);
or UO_2476 (O_2476,N_16146,N_16659);
nand UO_2477 (O_2477,N_18784,N_16349);
and UO_2478 (O_2478,N_16971,N_19538);
xor UO_2479 (O_2479,N_16295,N_18847);
and UO_2480 (O_2480,N_17540,N_16827);
xor UO_2481 (O_2481,N_16719,N_18318);
or UO_2482 (O_2482,N_18321,N_16076);
nand UO_2483 (O_2483,N_19782,N_16423);
nand UO_2484 (O_2484,N_17895,N_19164);
or UO_2485 (O_2485,N_16038,N_17648);
nor UO_2486 (O_2486,N_17854,N_16276);
and UO_2487 (O_2487,N_16269,N_19031);
and UO_2488 (O_2488,N_18327,N_16774);
and UO_2489 (O_2489,N_16972,N_19928);
nor UO_2490 (O_2490,N_17855,N_18561);
and UO_2491 (O_2491,N_16410,N_16963);
xor UO_2492 (O_2492,N_18019,N_19091);
or UO_2493 (O_2493,N_18381,N_17411);
or UO_2494 (O_2494,N_17247,N_18472);
and UO_2495 (O_2495,N_19129,N_19514);
nor UO_2496 (O_2496,N_17425,N_19400);
nor UO_2497 (O_2497,N_19389,N_17573);
nor UO_2498 (O_2498,N_17988,N_19896);
and UO_2499 (O_2499,N_17663,N_16838);
endmodule