module basic_5000_50000_5000_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_2147,In_299);
or U1 (N_1,In_1268,In_450);
xnor U2 (N_2,In_3495,In_2777);
nor U3 (N_3,In_4458,In_2918);
or U4 (N_4,In_2518,In_2114);
and U5 (N_5,In_4111,In_876);
and U6 (N_6,In_686,In_1652);
nor U7 (N_7,In_2190,In_4141);
nand U8 (N_8,In_1358,In_4201);
nor U9 (N_9,In_3986,In_1735);
and U10 (N_10,In_3172,In_600);
nand U11 (N_11,In_1991,In_3686);
or U12 (N_12,In_3559,In_2782);
xnor U13 (N_13,In_29,In_1870);
nor U14 (N_14,In_37,In_992);
nand U15 (N_15,In_4855,In_4103);
or U16 (N_16,In_4820,In_1861);
nor U17 (N_17,In_566,In_3410);
xnor U18 (N_18,In_3133,In_2880);
nand U19 (N_19,In_954,In_4396);
nor U20 (N_20,In_2286,In_1212);
and U21 (N_21,In_731,In_3781);
xor U22 (N_22,In_724,In_2496);
or U23 (N_23,In_732,In_1131);
or U24 (N_24,In_4900,In_52);
xor U25 (N_25,In_2311,In_3914);
nor U26 (N_26,In_4957,In_26);
nand U27 (N_27,In_401,In_369);
nand U28 (N_28,In_4156,In_3078);
and U29 (N_29,In_1666,In_3115);
nor U30 (N_30,In_1320,In_2099);
xor U31 (N_31,In_4801,In_4427);
and U32 (N_32,In_2781,In_766);
and U33 (N_33,In_2040,In_1468);
or U34 (N_34,In_2422,In_4);
xnor U35 (N_35,In_3585,In_2107);
nand U36 (N_36,In_3232,In_4868);
or U37 (N_37,In_843,In_171);
xnor U38 (N_38,In_4232,In_1348);
nand U39 (N_39,In_3441,In_1981);
xor U40 (N_40,In_4846,In_4492);
xnor U41 (N_41,In_2624,In_2587);
nor U42 (N_42,In_3198,In_877);
nand U43 (N_43,In_4324,In_3875);
xnor U44 (N_44,In_3493,In_3009);
nor U45 (N_45,In_95,In_4649);
xor U46 (N_46,In_183,In_2870);
nor U47 (N_47,In_2800,In_2690);
nand U48 (N_48,In_4574,In_2710);
xnor U49 (N_49,In_4524,In_1311);
nand U50 (N_50,In_2684,In_3934);
nand U51 (N_51,In_474,In_1332);
xnor U52 (N_52,In_1768,In_442);
or U53 (N_53,In_1473,In_2689);
nor U54 (N_54,In_2441,In_2192);
or U55 (N_55,In_2671,In_2277);
nand U56 (N_56,In_4695,In_1542);
nor U57 (N_57,In_2351,In_3558);
and U58 (N_58,In_4843,In_1974);
nor U59 (N_59,In_2626,In_4025);
nand U60 (N_60,In_3208,In_2036);
nor U61 (N_61,In_727,In_886);
nand U62 (N_62,In_2084,In_2322);
and U63 (N_63,In_3784,In_759);
or U64 (N_64,In_1241,In_697);
nand U65 (N_65,In_1979,In_3600);
nor U66 (N_66,In_1699,In_792);
xnor U67 (N_67,In_1580,In_788);
nor U68 (N_68,In_2071,In_2905);
nand U69 (N_69,In_162,In_1539);
xor U70 (N_70,In_3615,In_468);
nor U71 (N_71,In_3161,In_1236);
nor U72 (N_72,In_2180,In_1294);
xor U73 (N_73,In_3909,In_1327);
nand U74 (N_74,In_1692,In_1915);
and U75 (N_75,In_2733,In_247);
xor U76 (N_76,In_2120,In_2765);
nor U77 (N_77,In_201,In_2605);
nand U78 (N_78,In_167,In_4892);
xor U79 (N_79,In_2279,In_4350);
or U80 (N_80,In_3206,In_3478);
nand U81 (N_81,In_3840,In_4496);
nand U82 (N_82,In_4858,In_3060);
and U83 (N_83,In_3173,In_2961);
or U84 (N_84,In_4887,In_1078);
and U85 (N_85,In_885,In_2149);
and U86 (N_86,In_3066,In_1695);
or U87 (N_87,In_879,In_4857);
and U88 (N_88,In_4126,In_2810);
and U89 (N_89,In_3494,In_4880);
or U90 (N_90,In_1086,In_1193);
nor U91 (N_91,In_24,In_3728);
xor U92 (N_92,In_113,In_2720);
and U93 (N_93,In_4726,In_2478);
xnor U94 (N_94,In_1724,In_3873);
nor U95 (N_95,In_748,In_605);
and U96 (N_96,In_1855,In_3705);
xnor U97 (N_97,In_1544,In_4230);
or U98 (N_98,In_4135,In_2318);
or U99 (N_99,In_4040,In_812);
nand U100 (N_100,In_4883,In_1484);
xnor U101 (N_101,In_1481,In_3136);
xnor U102 (N_102,In_826,In_1156);
xnor U103 (N_103,In_2725,In_875);
nand U104 (N_104,In_1992,In_4722);
xor U105 (N_105,In_152,In_1373);
and U106 (N_106,In_578,In_439);
xor U107 (N_107,In_2230,In_2039);
or U108 (N_108,In_4631,In_915);
and U109 (N_109,In_3313,In_2968);
nand U110 (N_110,In_1231,In_88);
xnor U111 (N_111,In_4203,In_1017);
and U112 (N_112,In_1164,In_185);
or U113 (N_113,In_1772,In_4371);
xor U114 (N_114,In_4504,In_583);
xnor U115 (N_115,In_3716,In_3997);
or U116 (N_116,In_3552,In_1764);
xor U117 (N_117,In_4788,In_3393);
nor U118 (N_118,In_3423,In_391);
or U119 (N_119,In_2633,In_1219);
nor U120 (N_120,In_548,In_4740);
nand U121 (N_121,In_1020,In_4784);
and U122 (N_122,In_3646,In_778);
nor U123 (N_123,In_3571,In_1505);
nand U124 (N_124,In_4196,In_3853);
xnor U125 (N_125,In_4330,In_1963);
or U126 (N_126,In_2111,In_2297);
or U127 (N_127,In_2571,In_2257);
xor U128 (N_128,In_136,In_2704);
or U129 (N_129,In_1530,In_4790);
xnor U130 (N_130,In_1006,In_2523);
or U131 (N_131,In_4665,In_3012);
and U132 (N_132,In_4739,In_4598);
nand U133 (N_133,In_4848,In_2421);
nand U134 (N_134,In_404,In_3209);
and U135 (N_135,In_3202,In_4377);
nor U136 (N_136,In_2520,In_1947);
or U137 (N_137,In_2525,In_77);
nor U138 (N_138,In_4394,In_2156);
and U139 (N_139,In_2592,In_4837);
nor U140 (N_140,In_365,In_4208);
nor U141 (N_141,In_1988,In_713);
and U142 (N_142,In_3946,In_4529);
nor U143 (N_143,In_1689,In_4656);
xnor U144 (N_144,In_485,In_475);
or U145 (N_145,In_2160,In_3471);
nor U146 (N_146,In_232,In_4193);
and U147 (N_147,In_4482,In_830);
nor U148 (N_148,In_2555,In_2137);
nand U149 (N_149,In_2695,In_2657);
xnor U150 (N_150,In_4319,In_1548);
nor U151 (N_151,In_619,In_2983);
xnor U152 (N_152,In_208,In_603);
xor U153 (N_153,In_3735,In_1985);
xnor U154 (N_154,In_899,In_3910);
nor U155 (N_155,In_1182,In_747);
and U156 (N_156,In_3469,In_2197);
or U157 (N_157,In_3847,In_2390);
or U158 (N_158,In_3556,In_2463);
xor U159 (N_159,In_402,In_3650);
xnor U160 (N_160,In_3015,In_4229);
xnor U161 (N_161,In_4045,In_416);
nor U162 (N_162,In_4415,In_4092);
nor U163 (N_163,In_3708,In_1595);
and U164 (N_164,In_4516,In_9);
nor U165 (N_165,In_2090,In_317);
or U166 (N_166,In_2429,In_3971);
nor U167 (N_167,In_3288,In_470);
xnor U168 (N_168,In_4931,In_2260);
nor U169 (N_169,In_4617,In_3320);
xor U170 (N_170,In_4948,In_4460);
nand U171 (N_171,In_126,In_4834);
nand U172 (N_172,In_1611,In_4452);
nand U173 (N_173,In_2258,In_3635);
nor U174 (N_174,In_1584,In_1977);
xnor U175 (N_175,In_3321,In_1546);
nand U176 (N_176,In_139,In_2508);
or U177 (N_177,In_488,In_2759);
xor U178 (N_178,In_3129,In_4685);
nor U179 (N_179,In_4313,In_370);
xnor U180 (N_180,In_3003,In_698);
or U181 (N_181,In_3700,In_1079);
xnor U182 (N_182,In_4218,In_4076);
xor U183 (N_183,In_1346,In_3151);
nand U184 (N_184,In_4199,In_170);
nand U185 (N_185,In_1383,In_1970);
xor U186 (N_186,In_949,In_4128);
xnor U187 (N_187,In_3818,In_522);
xor U188 (N_188,In_498,In_829);
nand U189 (N_189,In_4778,In_1005);
xnor U190 (N_190,In_2977,In_1293);
xor U191 (N_191,In_2616,In_3597);
xnor U192 (N_192,In_1479,In_3276);
nor U193 (N_193,In_4873,In_3497);
and U194 (N_194,In_2025,In_1978);
nor U195 (N_195,In_3359,In_3079);
and U196 (N_196,In_48,In_2970);
nand U197 (N_197,In_2467,In_1269);
and U198 (N_198,In_1625,In_2221);
nor U199 (N_199,In_2858,In_2900);
xnor U200 (N_200,In_4049,In_358);
or U201 (N_201,In_1547,In_4202);
and U202 (N_202,In_1066,In_258);
nor U203 (N_203,In_2802,In_4992);
or U204 (N_204,In_814,In_371);
nand U205 (N_205,In_3724,In_245);
and U206 (N_206,In_460,In_852);
nand U207 (N_207,In_2327,In_1853);
or U208 (N_208,In_3395,In_1845);
or U209 (N_209,In_880,In_959);
and U210 (N_210,In_284,In_702);
nor U211 (N_211,In_1921,In_2052);
xor U212 (N_212,In_4105,In_133);
or U213 (N_213,In_4023,In_3461);
xor U214 (N_214,In_3622,In_1372);
nand U215 (N_215,In_4961,In_325);
xor U216 (N_216,In_4949,In_1141);
nor U217 (N_217,In_2404,In_3425);
or U218 (N_218,In_525,In_2722);
and U219 (N_219,In_4247,In_776);
nand U220 (N_220,In_2285,In_2771);
or U221 (N_221,In_4558,In_3987);
nor U222 (N_222,In_492,In_3500);
nor U223 (N_223,In_2335,In_1564);
nor U224 (N_224,In_907,In_2964);
xor U225 (N_225,In_586,In_3007);
and U226 (N_226,In_2339,In_173);
nand U227 (N_227,In_4954,In_1211);
nand U228 (N_228,In_1379,In_1550);
nand U229 (N_229,In_3286,In_1744);
xor U230 (N_230,In_4173,In_4764);
and U231 (N_231,In_2187,In_582);
nor U232 (N_232,In_2979,In_970);
nor U233 (N_233,In_769,In_4802);
xor U234 (N_234,In_3326,In_952);
nor U235 (N_235,In_4502,In_408);
and U236 (N_236,In_1682,In_2564);
or U237 (N_237,In_4355,In_782);
xor U238 (N_238,In_4841,In_2613);
nor U239 (N_239,In_914,In_2691);
and U240 (N_240,In_432,In_39);
nor U241 (N_241,In_4024,In_335);
and U242 (N_242,In_656,In_3357);
or U243 (N_243,In_226,In_2313);
xnor U244 (N_244,In_3034,In_1901);
and U245 (N_245,In_3611,In_2216);
nor U246 (N_246,In_2888,In_1387);
and U247 (N_247,In_3898,In_524);
or U248 (N_248,In_2239,In_2790);
or U249 (N_249,In_93,In_3316);
nor U250 (N_250,In_1408,In_1265);
nand U251 (N_251,In_602,In_2761);
nor U252 (N_252,In_4192,In_3435);
or U253 (N_253,In_4941,In_3373);
xnor U254 (N_254,In_1810,In_2031);
nand U255 (N_255,In_2213,In_84);
xor U256 (N_256,In_1030,In_2336);
nor U257 (N_257,In_3107,In_2032);
xnor U258 (N_258,In_833,In_4937);
and U259 (N_259,In_339,In_1951);
nand U260 (N_260,In_3103,In_1579);
nor U261 (N_261,In_699,In_4683);
and U262 (N_262,In_4181,In_2576);
nor U263 (N_263,In_3630,In_4386);
xor U264 (N_264,In_2927,In_2836);
and U265 (N_265,In_2075,In_3117);
xor U266 (N_266,In_2848,In_2009);
nand U267 (N_267,In_2632,In_683);
nor U268 (N_268,In_2565,In_206);
nand U269 (N_269,In_3950,In_517);
or U270 (N_270,In_212,In_1752);
or U271 (N_271,In_4719,In_4073);
xor U272 (N_272,In_3381,In_3959);
nand U273 (N_273,In_1899,In_3045);
xnor U274 (N_274,In_4870,In_2225);
or U275 (N_275,In_4256,In_3838);
and U276 (N_276,In_387,In_4531);
nand U277 (N_277,In_3119,In_2340);
or U278 (N_278,In_1248,In_3280);
nor U279 (N_279,In_3805,In_1421);
nor U280 (N_280,In_2492,In_967);
xor U281 (N_281,In_446,In_2003);
or U282 (N_282,In_3140,In_2358);
nand U283 (N_283,In_4109,In_240);
and U284 (N_284,In_2083,In_4430);
and U285 (N_285,In_4162,In_1243);
xor U286 (N_286,In_3148,In_3989);
xor U287 (N_287,In_3378,In_4535);
xor U288 (N_288,In_72,In_4602);
nor U289 (N_289,In_4331,In_2312);
and U290 (N_290,In_3601,In_2785);
and U291 (N_291,In_503,In_1249);
or U292 (N_292,In_2569,In_803);
or U293 (N_293,In_3549,In_1043);
xor U294 (N_294,In_3037,In_754);
nand U295 (N_295,In_3331,In_2686);
nand U296 (N_296,In_4470,In_4865);
or U297 (N_297,In_250,In_112);
xor U298 (N_298,In_4952,In_2857);
or U299 (N_299,In_41,In_3257);
nand U300 (N_300,In_1700,In_943);
nand U301 (N_301,In_308,In_2756);
or U302 (N_302,In_4048,In_2195);
nand U303 (N_303,In_922,In_1759);
nand U304 (N_304,In_1185,In_558);
xnor U305 (N_305,In_944,In_584);
or U306 (N_306,In_2899,In_4812);
nand U307 (N_307,In_1897,In_4494);
or U308 (N_308,In_4225,In_4720);
nor U309 (N_309,In_4673,In_4353);
or U310 (N_310,In_3044,In_1707);
nor U311 (N_311,In_3083,In_2519);
xnor U312 (N_312,In_806,In_4786);
and U313 (N_313,In_4484,In_1391);
nand U314 (N_314,In_3504,In_4804);
nor U315 (N_315,In_489,In_2367);
and U316 (N_316,In_3391,In_1696);
nor U317 (N_317,In_4099,In_1366);
nor U318 (N_318,In_4934,In_2374);
nand U319 (N_319,In_4258,In_1889);
xnor U320 (N_320,In_83,In_4140);
or U321 (N_321,In_2353,In_3598);
nand U322 (N_322,In_1990,In_3297);
or U323 (N_323,In_2643,In_1177);
nor U324 (N_324,In_4606,In_2490);
or U325 (N_325,In_2506,In_1057);
nand U326 (N_326,In_2646,In_1957);
nor U327 (N_327,In_1198,In_4479);
xor U328 (N_328,In_1021,In_1515);
xor U329 (N_329,In_3932,In_4416);
nand U330 (N_330,In_60,In_4002);
nand U331 (N_331,In_2469,In_2864);
xor U332 (N_332,In_1954,In_2893);
xor U333 (N_333,In_2935,In_4457);
or U334 (N_334,In_3019,In_599);
nor U335 (N_335,In_628,In_4972);
xnor U336 (N_336,In_2826,In_4495);
xnor U337 (N_337,In_2162,In_3918);
xnor U338 (N_338,In_1636,In_4565);
or U339 (N_339,In_2892,In_1235);
and U340 (N_340,In_2247,In_3564);
or U341 (N_341,In_2678,In_1702);
nand U342 (N_342,In_3962,In_3570);
nor U343 (N_343,In_1731,In_3548);
nor U344 (N_344,In_497,In_1723);
nand U345 (N_345,In_2282,In_4985);
nor U346 (N_346,In_2827,In_4071);
and U347 (N_347,In_3056,In_2941);
nor U348 (N_348,In_2499,In_4263);
nor U349 (N_349,In_405,In_1382);
or U350 (N_350,In_62,In_815);
xor U351 (N_351,In_3820,In_2098);
or U352 (N_352,In_4155,In_3372);
or U353 (N_353,In_4669,In_3744);
xnor U354 (N_354,In_2673,In_3569);
nor U355 (N_355,In_2168,In_714);
xnor U356 (N_356,In_3546,In_3167);
nand U357 (N_357,In_641,In_1423);
and U358 (N_358,In_1307,In_1342);
xor U359 (N_359,In_2152,In_1047);
nor U360 (N_360,In_1393,In_3138);
or U361 (N_361,In_3530,In_2418);
nand U362 (N_362,In_1830,In_1628);
or U363 (N_363,In_2489,In_1354);
nand U364 (N_364,In_2922,In_4754);
nand U365 (N_365,In_3089,In_2253);
xnor U366 (N_366,In_2459,In_3018);
and U367 (N_367,In_3480,In_3868);
or U368 (N_368,In_636,In_1167);
and U369 (N_369,In_42,In_244);
or U370 (N_370,In_4036,In_75);
xor U371 (N_371,In_1704,In_4997);
xnor U372 (N_372,In_3978,In_3751);
and U373 (N_373,In_1869,In_608);
nor U374 (N_374,In_1642,In_2682);
xnor U375 (N_375,In_1326,In_398);
and U376 (N_376,In_4026,In_1074);
or U377 (N_377,In_2602,In_2159);
or U378 (N_378,In_4051,In_1728);
nor U379 (N_379,In_2234,In_700);
and U380 (N_380,In_3839,In_809);
nand U381 (N_381,In_4833,In_2360);
nor U382 (N_382,In_4815,In_298);
and U383 (N_383,In_2661,In_4775);
nand U384 (N_384,In_1431,In_860);
xnor U385 (N_385,In_2373,In_672);
nand U386 (N_386,In_4907,In_891);
nor U387 (N_387,In_4269,In_651);
nor U388 (N_388,In_1280,In_4862);
xnor U389 (N_389,In_4487,In_2537);
and U390 (N_390,In_3205,In_2536);
and U391 (N_391,In_2488,In_2882);
and U392 (N_392,In_1753,In_1446);
or U393 (N_393,In_4559,In_3656);
and U394 (N_394,In_2862,In_3464);
nand U395 (N_395,In_4534,In_1649);
xnor U396 (N_396,In_1173,In_2116);
and U397 (N_397,In_307,In_1794);
or U398 (N_398,In_2744,In_4762);
and U399 (N_399,In_1864,In_4178);
and U400 (N_400,In_4747,In_1333);
nand U401 (N_401,In_4399,In_2881);
nand U402 (N_402,In_3879,In_3443);
nand U403 (N_403,In_2685,In_3057);
nor U404 (N_404,In_3929,In_33);
nor U405 (N_405,In_81,In_3524);
nor U406 (N_406,In_3479,In_690);
xor U407 (N_407,In_3455,In_4185);
nand U408 (N_408,In_4551,In_4710);
nand U409 (N_409,In_3251,In_3557);
and U410 (N_410,In_3177,In_4736);
and U411 (N_411,In_2971,In_2144);
and U412 (N_412,In_65,In_1925);
and U413 (N_413,In_606,In_69);
and U414 (N_414,In_3030,In_1129);
xor U415 (N_415,In_4237,In_2424);
or U416 (N_416,In_594,In_4876);
or U417 (N_417,In_4299,In_1594);
nand U418 (N_418,In_2430,In_4822);
and U419 (N_419,In_2076,In_1306);
nand U420 (N_420,In_1982,In_1045);
nand U421 (N_421,In_310,In_4465);
nand U422 (N_422,In_1619,In_1205);
or U423 (N_423,In_3289,In_3399);
and U424 (N_424,In_1412,In_3587);
or U425 (N_425,In_3884,In_900);
or U426 (N_426,In_2997,In_3295);
nor U427 (N_427,In_4334,In_3786);
xor U428 (N_428,In_2333,In_4031);
or U429 (N_429,In_3091,In_462);
nor U430 (N_430,In_729,In_4339);
nand U431 (N_431,In_314,In_4962);
nor U432 (N_432,In_137,In_4806);
xnor U433 (N_433,In_1487,In_2635);
nor U434 (N_434,In_4279,In_287);
xnor U435 (N_435,In_1471,In_740);
and U436 (N_436,In_768,In_1827);
xor U437 (N_437,In_3024,In_242);
nand U438 (N_438,In_246,In_2805);
and U439 (N_439,In_3709,In_3125);
and U440 (N_440,In_2603,In_3970);
nand U441 (N_441,In_3921,In_1763);
nand U442 (N_442,In_3219,In_1941);
nor U443 (N_443,In_591,In_2474);
or U444 (N_444,In_4012,In_1821);
and U445 (N_445,In_741,In_4356);
nor U446 (N_446,In_1739,In_1210);
or U447 (N_447,In_3513,In_4976);
and U448 (N_448,In_1305,In_1665);
nand U449 (N_449,In_2804,In_3649);
nor U450 (N_450,In_2020,In_3156);
xnor U451 (N_451,In_3106,In_2687);
nand U452 (N_452,In_3163,In_1409);
and U453 (N_453,In_3896,In_2109);
or U454 (N_454,In_3434,In_1557);
xnor U455 (N_455,In_4715,In_1968);
nor U456 (N_456,In_3269,In_3991);
or U457 (N_457,In_4898,In_4829);
nor U458 (N_458,In_3722,In_3127);
xor U459 (N_459,In_1247,In_1742);
nand U460 (N_460,In_4944,In_388);
xnor U461 (N_461,In_2302,In_571);
and U462 (N_462,In_67,In_1002);
xor U463 (N_463,In_3666,In_2991);
and U464 (N_464,In_3928,In_2341);
nor U465 (N_465,In_3942,In_3827);
or U466 (N_466,In_4498,In_3953);
nor U467 (N_467,In_3406,In_1110);
xnor U468 (N_468,In_2960,In_4159);
or U469 (N_469,In_2165,In_527);
and U470 (N_470,In_8,In_4338);
and U471 (N_471,In_4364,In_502);
nand U472 (N_472,In_3327,In_3301);
nand U473 (N_473,In_4995,In_3528);
and U474 (N_474,In_4176,In_3706);
nor U475 (N_475,In_3927,In_887);
nand U476 (N_476,In_273,In_3804);
or U477 (N_477,In_3926,In_3794);
nand U478 (N_478,In_961,In_1256);
nand U479 (N_479,In_4453,In_2011);
or U480 (N_480,In_4821,In_2493);
xnor U481 (N_481,In_919,In_2219);
nor U482 (N_482,In_3508,In_718);
nand U483 (N_483,In_2609,In_1840);
xor U484 (N_484,In_3193,In_4861);
nand U485 (N_485,In_1132,In_3977);
or U486 (N_486,In_147,In_169);
nor U487 (N_487,In_3312,In_615);
nand U488 (N_488,In_4456,In_3484);
xor U489 (N_489,In_1761,In_3711);
or U490 (N_490,In_3618,In_1832);
xnor U491 (N_491,In_3667,In_719);
xor U492 (N_492,In_4958,In_1819);
or U493 (N_493,In_4678,In_665);
nand U494 (N_494,In_2588,In_1658);
or U495 (N_495,In_1520,In_1806);
or U496 (N_496,In_4904,In_1715);
nand U497 (N_497,In_4780,In_260);
nand U498 (N_498,In_4632,In_4426);
and U499 (N_499,In_3768,In_4630);
and U500 (N_500,In_2223,In_1113);
or U501 (N_501,In_4368,In_1778);
nand U502 (N_502,In_323,In_3956);
and U503 (N_503,In_3064,In_4517);
and U504 (N_504,In_4046,In_2698);
nor U505 (N_505,In_2731,In_901);
xnor U506 (N_506,In_312,In_2191);
and U507 (N_507,In_4971,In_4127);
nor U508 (N_508,In_2411,In_2167);
nand U509 (N_509,In_3499,In_2739);
and U510 (N_510,In_3973,In_4610);
nor U511 (N_511,In_3438,In_2129);
and U512 (N_512,In_3885,In_596);
or U513 (N_513,In_3645,In_111);
xor U514 (N_514,In_3099,In_2679);
or U515 (N_515,In_1524,In_4627);
xnor U516 (N_516,In_4578,In_2141);
nor U517 (N_517,In_4645,In_397);
and U518 (N_518,In_1894,In_4851);
or U519 (N_519,In_3290,In_706);
xor U520 (N_520,In_351,In_908);
or U521 (N_521,In_2064,In_3258);
or U522 (N_522,In_3603,In_1614);
nand U523 (N_523,In_2701,In_487);
and U524 (N_524,In_4360,In_1470);
and U525 (N_525,In_4303,In_3743);
xor U526 (N_526,In_3002,In_196);
or U527 (N_527,In_438,In_3848);
nand U528 (N_528,In_1621,In_1558);
nand U529 (N_529,In_2153,In_2504);
and U530 (N_530,In_491,In_4807);
xnor U531 (N_531,In_4342,In_1790);
nor U532 (N_532,In_4867,In_1023);
or U533 (N_533,In_4800,In_2948);
nor U534 (N_534,In_4318,In_4891);
xnor U535 (N_535,In_3979,In_3476);
or U536 (N_536,In_775,In_4007);
xnor U537 (N_537,In_345,In_4871);
and U538 (N_538,In_1106,In_3566);
nand U539 (N_539,In_2926,In_3067);
or U540 (N_540,In_2178,In_2772);
nor U541 (N_541,In_4792,In_4357);
or U542 (N_542,In_3878,In_966);
nand U543 (N_543,In_3980,In_2329);
and U544 (N_544,In_3159,In_629);
nand U545 (N_545,In_3539,In_2887);
and U546 (N_546,In_1807,In_4566);
xor U547 (N_547,In_3574,In_4511);
xnor U548 (N_548,In_4349,In_361);
and U549 (N_549,In_1049,In_4284);
or U550 (N_550,In_1678,In_4179);
xor U551 (N_551,In_984,In_4696);
and U552 (N_552,In_3561,In_1202);
and U553 (N_553,In_403,In_1290);
nor U554 (N_554,In_4276,In_3006);
nor U555 (N_555,In_2362,In_4096);
nor U556 (N_556,In_215,In_2319);
nand U557 (N_557,In_2974,In_1606);
xor U558 (N_558,In_1802,In_3033);
xor U559 (N_559,In_4682,In_4010);
and U560 (N_560,In_3254,In_50);
and U561 (N_561,In_449,In_296);
and U562 (N_562,In_471,In_534);
nand U563 (N_563,In_2818,In_3826);
nand U564 (N_564,In_2204,In_2133);
nor U565 (N_565,In_1615,In_2610);
nor U566 (N_566,In_2397,In_4358);
nor U567 (N_567,In_4908,In_2017);
nor U568 (N_568,In_749,In_4047);
and U569 (N_569,In_3800,In_35);
and U570 (N_570,In_516,In_1805);
or U571 (N_571,In_2950,In_873);
nor U572 (N_572,In_4850,In_2929);
nand U573 (N_573,In_597,In_4896);
or U574 (N_574,In_1116,In_3329);
nor U575 (N_575,In_4413,In_3139);
or U576 (N_576,In_4760,In_1643);
and U577 (N_577,In_367,In_3305);
nor U578 (N_578,In_3184,In_3769);
or U579 (N_579,In_642,In_2649);
or U580 (N_580,In_211,In_12);
or U581 (N_581,In_300,In_3682);
or U582 (N_582,In_227,In_3562);
or U583 (N_583,In_1851,In_1750);
and U584 (N_584,In_3352,In_4414);
or U585 (N_585,In_236,In_4583);
nand U586 (N_586,In_2956,In_1267);
or U587 (N_587,In_1053,In_1622);
nor U588 (N_588,In_4171,In_329);
nor U589 (N_589,In_1835,In_705);
xnor U590 (N_590,In_3851,In_2269);
nor U591 (N_591,In_3542,In_181);
or U592 (N_592,In_3354,In_3368);
nor U593 (N_593,In_4499,In_1814);
or U594 (N_594,In_722,In_3203);
xor U595 (N_595,In_3846,In_1285);
and U596 (N_596,In_2057,In_1822);
xnor U597 (N_597,In_3068,In_4875);
nand U598 (N_598,In_2189,In_3102);
nor U599 (N_599,In_565,In_2224);
and U600 (N_600,In_1148,In_575);
or U601 (N_601,In_4869,In_3902);
or U602 (N_602,In_2295,In_3748);
and U603 (N_603,In_2259,In_2041);
nor U604 (N_604,In_3070,In_1910);
and U605 (N_605,In_2112,In_1708);
nand U606 (N_606,In_1850,In_892);
nand U607 (N_607,In_4455,In_3467);
nand U608 (N_608,In_2483,In_3685);
nand U609 (N_609,In_4477,In_2018);
xor U610 (N_610,In_3581,In_1025);
nor U611 (N_611,In_1599,In_840);
and U612 (N_612,In_1999,In_3533);
nand U613 (N_613,In_2254,In_1858);
xor U614 (N_614,In_3105,In_2395);
and U615 (N_615,In_3224,In_3988);
or U616 (N_616,In_2370,In_3841);
or U617 (N_617,In_935,In_3338);
nand U618 (N_618,In_1261,In_1007);
nand U619 (N_619,In_3101,In_4068);
and U620 (N_620,In_2629,In_623);
nor U621 (N_621,In_4252,In_1157);
xnor U622 (N_622,In_2650,In_607);
or U623 (N_623,In_2473,In_3418);
nor U624 (N_624,In_950,In_904);
or U625 (N_625,In_654,In_1533);
or U626 (N_626,In_556,In_1693);
xnor U627 (N_627,In_121,In_384);
nand U628 (N_628,In_1300,In_2348);
nor U629 (N_629,In_2487,In_2108);
nand U630 (N_630,In_2540,In_1062);
or U631 (N_631,In_1959,In_2222);
xor U632 (N_632,In_3594,In_3080);
and U633 (N_633,In_2066,In_1318);
nand U634 (N_634,In_677,In_853);
xnor U635 (N_635,In_521,In_2524);
nor U636 (N_636,In_2821,In_3732);
xnor U637 (N_637,In_1077,In_494);
nor U638 (N_638,In_59,In_1691);
and U639 (N_639,In_4637,In_1811);
and U640 (N_640,In_3725,In_1415);
nand U641 (N_641,In_4735,In_1140);
xnor U642 (N_642,In_4309,In_3757);
nor U643 (N_643,In_3755,In_4044);
xnor U644 (N_644,In_3050,In_878);
nand U645 (N_645,In_3882,In_1426);
or U646 (N_646,In_3216,In_1093);
xor U647 (N_647,In_3382,In_1698);
or U648 (N_648,In_4038,In_2659);
xor U649 (N_649,In_3488,In_3249);
nand U650 (N_650,In_4652,In_2732);
and U651 (N_651,In_1996,In_3220);
nor U652 (N_652,In_3937,In_1168);
and U653 (N_653,In_4432,In_4991);
nand U654 (N_654,In_1741,In_3659);
nor U655 (N_655,In_4582,In_2012);
nor U656 (N_656,In_3259,In_2859);
or U657 (N_657,In_2442,In_1390);
nor U658 (N_658,In_3131,In_1879);
nor U659 (N_659,In_3903,In_1197);
nand U660 (N_660,In_153,In_1499);
xor U661 (N_661,In_140,In_3069);
xnor U662 (N_662,In_3958,In_376);
and U663 (N_663,In_3128,In_2644);
and U664 (N_664,In_2202,In_2349);
xor U665 (N_665,In_4996,In_3141);
and U666 (N_666,In_4332,In_3752);
or U667 (N_667,In_248,In_4708);
nand U668 (N_668,In_2126,In_3941);
nand U669 (N_669,In_4088,In_4072);
nand U670 (N_670,In_862,In_507);
or U671 (N_671,In_3766,In_1514);
nor U672 (N_672,In_311,In_3309);
and U673 (N_673,In_817,In_1801);
xnor U674 (N_674,In_3887,In_4226);
or U675 (N_675,In_2501,In_1588);
nand U676 (N_676,In_4227,In_4737);
or U677 (N_677,In_294,In_1122);
xor U678 (N_678,In_4429,In_4572);
nand U679 (N_679,In_1195,In_73);
nor U680 (N_680,In_1798,In_1559);
nor U681 (N_681,In_3639,In_477);
and U682 (N_682,In_1142,In_1532);
and U683 (N_683,In_4605,In_4940);
and U684 (N_684,In_4508,In_723);
nand U685 (N_685,In_4005,In_129);
xnor U686 (N_686,In_3404,In_3351);
xnor U687 (N_687,In_3417,In_3680);
or U688 (N_688,In_3591,In_4098);
or U689 (N_689,In_479,In_306);
or U690 (N_690,In_4294,In_51);
xnor U691 (N_691,In_1048,In_2766);
and U692 (N_692,In_2078,In_657);
or U693 (N_693,In_1402,In_1826);
or U694 (N_694,In_1161,In_1174);
and U695 (N_695,In_78,In_4419);
nor U696 (N_696,In_1089,In_1638);
nor U697 (N_697,In_3093,In_3165);
or U698 (N_698,In_3714,In_2205);
nor U699 (N_699,In_4174,In_3111);
xnor U700 (N_700,In_363,In_2023);
xor U701 (N_701,In_4717,In_1799);
xnor U702 (N_702,In_2871,In_906);
nand U703 (N_703,In_4700,In_531);
xor U704 (N_704,In_1808,In_2444);
nand U705 (N_705,In_1782,In_218);
nand U706 (N_706,In_2396,In_664);
xnor U707 (N_707,In_4160,In_1872);
or U708 (N_708,In_1685,In_4505);
and U709 (N_709,In_186,In_3814);
nand U710 (N_710,In_155,In_1867);
or U711 (N_711,In_3745,In_4439);
and U712 (N_712,In_3923,In_3341);
nor U713 (N_713,In_457,In_4009);
nor U714 (N_714,In_913,In_415);
xor U715 (N_715,In_832,In_1068);
nand U716 (N_716,In_4235,In_2070);
or U717 (N_717,In_1151,In_36);
or U718 (N_718,In_4543,In_4286);
nand U719 (N_719,In_2642,In_574);
nand U720 (N_720,In_1166,In_1458);
or U721 (N_721,In_1895,In_3054);
nand U722 (N_722,In_277,In_822);
or U723 (N_723,In_58,In_496);
and U724 (N_724,In_1476,In_1730);
xor U725 (N_725,In_3737,In_3966);
nor U726 (N_726,In_2238,In_4372);
xor U727 (N_727,In_4351,In_356);
and U728 (N_728,In_3081,In_1883);
and U729 (N_729,In_3323,In_4446);
and U730 (N_730,In_4897,In_4878);
or U731 (N_731,In_559,In_637);
or U732 (N_732,In_4134,In_1440);
or U733 (N_733,In_1629,In_64);
nor U734 (N_734,In_1781,In_1163);
and U735 (N_735,In_4677,In_426);
nor U736 (N_736,In_4395,In_2303);
nand U737 (N_737,In_813,In_704);
nand U738 (N_738,In_1430,In_2828);
and U739 (N_739,In_3631,In_1466);
nand U740 (N_740,In_845,In_2952);
or U741 (N_741,In_4734,In_392);
nor U742 (N_742,In_2102,In_4233);
and U743 (N_743,In_235,In_1125);
nand U744 (N_744,In_3892,In_4293);
nand U745 (N_745,In_604,In_2403);
xor U746 (N_746,In_2751,In_2740);
nor U747 (N_747,In_1509,In_1083);
and U748 (N_748,In_381,In_3654);
nor U749 (N_749,In_3416,In_1726);
and U750 (N_750,In_220,In_4785);
nor U751 (N_751,In_3629,In_625);
nand U752 (N_752,In_989,In_4404);
xor U753 (N_753,In_4307,In_2807);
nor U754 (N_754,In_2125,In_243);
or U755 (N_755,In_1462,In_4621);
xnor U756 (N_756,In_2516,In_4753);
or U757 (N_757,In_400,In_3097);
or U758 (N_758,In_541,In_645);
and U759 (N_759,In_2,In_3616);
and U760 (N_760,In_2528,In_4794);
and U761 (N_761,In_4362,In_1881);
or U762 (N_762,In_2572,In_2969);
xor U763 (N_763,In_580,In_2631);
nor U764 (N_764,In_1111,In_156);
xor U765 (N_765,In_546,In_4333);
or U766 (N_766,In_1414,In_1134);
nand U767 (N_767,In_1108,In_2154);
nor U768 (N_768,In_3974,In_302);
nor U769 (N_769,In_1329,In_4367);
nor U770 (N_770,In_1732,In_781);
or U771 (N_771,In_1605,In_962);
nand U772 (N_772,In_2611,In_4927);
nor U773 (N_773,In_2276,In_4003);
xnor U774 (N_774,In_4058,In_3211);
or U775 (N_775,In_2658,In_4266);
xnor U776 (N_776,In_1276,In_1287);
nand U777 (N_777,In_4301,In_266);
xnor U778 (N_778,In_2580,In_4261);
nor U779 (N_779,In_2907,In_4172);
nor U780 (N_780,In_4709,In_1031);
xnor U781 (N_781,In_480,In_4315);
nor U782 (N_782,In_2829,In_4189);
nand U783 (N_783,In_1427,In_469);
or U784 (N_784,In_2868,In_2115);
or U785 (N_785,In_1158,In_1203);
nand U786 (N_786,In_4664,In_1404);
xnor U787 (N_787,In_4112,In_676);
or U788 (N_788,In_923,In_418);
xnor U789 (N_789,In_1461,In_2215);
and U790 (N_790,In_4589,In_1733);
xnor U791 (N_791,In_2482,In_2174);
and U792 (N_792,In_199,In_2408);
or U793 (N_793,In_1304,In_4809);
nand U794 (N_794,In_3271,In_2415);
or U795 (N_795,In_1124,In_4013);
xor U796 (N_796,In_3279,In_3049);
nand U797 (N_797,In_1135,In_3662);
and U798 (N_798,In_4445,In_2290);
nor U799 (N_799,In_14,In_2817);
xor U800 (N_800,In_3292,In_1289);
nor U801 (N_801,In_2177,In_3199);
nand U802 (N_802,In_2006,In_4744);
nand U803 (N_803,In_1491,In_2916);
and U804 (N_804,In_4808,In_1362);
nand U805 (N_805,In_2793,In_406);
nor U806 (N_806,In_4066,In_1075);
xnor U807 (N_807,In_3463,In_4206);
nand U808 (N_808,In_3931,In_11);
xor U809 (N_809,In_659,In_1922);
xnor U810 (N_810,In_3252,In_4724);
xnor U811 (N_811,In_3891,In_4831);
or U812 (N_812,In_3731,In_2914);
nand U813 (N_813,In_3537,In_4981);
xnor U814 (N_814,In_3789,In_932);
and U815 (N_815,In_557,In_3608);
nor U816 (N_816,In_4278,In_1312);
or U817 (N_817,In_3032,In_1647);
and U818 (N_818,In_627,In_303);
and U819 (N_819,In_4601,In_4953);
xnor U820 (N_820,In_4273,In_2591);
or U821 (N_821,In_4305,In_2433);
nor U822 (N_822,In_2080,In_1213);
xnor U823 (N_823,In_2988,In_3697);
nor U824 (N_824,In_1296,In_2620);
nor U825 (N_825,In_3756,In_1567);
nand U826 (N_826,In_1264,In_1187);
nor U827 (N_827,In_289,In_1224);
and U828 (N_828,In_1688,In_2990);
xnor U829 (N_829,In_4200,In_1989);
nor U830 (N_830,In_2059,In_4636);
nor U831 (N_831,In_1586,In_4894);
and U832 (N_832,In_2709,In_1225);
xnor U833 (N_833,In_3108,In_2513);
xnor U834 (N_834,In_4078,In_4905);
and U835 (N_835,In_1012,In_3710);
or U836 (N_836,In_2432,In_3375);
nor U837 (N_837,In_2884,In_2809);
and U838 (N_838,In_1186,In_2896);
and U839 (N_839,In_2885,In_1920);
or U840 (N_840,In_145,In_3554);
and U841 (N_841,In_4923,In_281);
nand U842 (N_842,In_3643,In_4343);
xnor U843 (N_843,In_2000,In_4466);
or U844 (N_844,In_4341,In_883);
xnor U845 (N_845,In_773,In_3046);
nand U846 (N_846,In_3636,In_2248);
or U847 (N_847,In_1380,In_4557);
nand U848 (N_848,In_3339,In_2250);
and U849 (N_849,In_3330,In_1714);
nor U850 (N_850,In_3187,In_3501);
nor U851 (N_851,In_2551,In_630);
nand U852 (N_852,In_2235,In_780);
or U853 (N_853,In_4547,In_2300);
nor U854 (N_854,In_1036,In_164);
nor U855 (N_855,In_573,In_1448);
and U856 (N_856,In_1035,In_1604);
and U857 (N_857,In_53,In_1659);
nor U858 (N_858,In_2825,In_4629);
xnor U859 (N_859,In_1145,In_4978);
nor U860 (N_860,In_1657,In_3540);
or U861 (N_861,In_2578,In_529);
nor U862 (N_862,In_4312,In_2532);
or U863 (N_863,In_4522,In_2727);
nand U864 (N_864,In_3483,In_3761);
xor U865 (N_865,In_2450,In_2618);
xnor U866 (N_866,In_3632,In_1597);
xor U867 (N_867,In_777,In_1956);
or U868 (N_868,In_2412,In_666);
or U869 (N_869,In_1712,In_4503);
nor U870 (N_870,In_3833,In_1748);
nand U871 (N_871,In_570,In_1422);
nor U872 (N_872,In_4835,In_3021);
xor U873 (N_873,In_3010,In_721);
or U874 (N_874,In_1841,In_2863);
or U875 (N_875,In_2366,In_2806);
and U876 (N_876,In_3189,In_1893);
nand U877 (N_877,In_3401,In_1252);
nor U878 (N_878,In_3039,In_3328);
nand U879 (N_879,In_1650,In_609);
and U880 (N_880,In_1206,In_1686);
nor U881 (N_881,In_3073,In_4836);
xnor U882 (N_882,In_894,In_3055);
or U883 (N_883,In_1627,In_1812);
nand U884 (N_884,In_1478,In_1653);
and U885 (N_885,In_6,In_3486);
and U886 (N_886,In_1934,In_2672);
xnor U887 (N_887,In_3578,In_4519);
xor U888 (N_888,In_1620,In_2867);
or U889 (N_889,In_1441,In_3344);
xor U890 (N_890,In_1818,In_61);
nand U891 (N_891,In_3451,In_551);
or U892 (N_892,In_1442,In_4169);
and U893 (N_893,In_466,In_2101);
or U894 (N_894,In_771,In_2494);
or U895 (N_895,In_930,In_4210);
or U896 (N_896,In_295,In_1705);
nor U897 (N_897,In_1208,In_4177);
or U898 (N_898,In_1144,In_643);
or U899 (N_899,In_3704,In_1189);
xor U900 (N_900,In_4947,In_4507);
or U901 (N_901,In_4545,In_4964);
xnor U902 (N_902,In_669,In_4770);
xor U903 (N_903,In_3759,In_549);
nor U904 (N_904,In_2791,In_241);
nand U905 (N_905,In_2559,In_1377);
or U906 (N_906,In_2556,In_1517);
or U907 (N_907,In_4746,In_1971);
and U908 (N_908,In_2797,In_4646);
xnor U909 (N_909,In_2324,In_455);
or U910 (N_910,In_1278,In_3110);
or U911 (N_911,In_4306,In_229);
xor U912 (N_912,In_1871,In_2094);
nor U913 (N_913,In_658,In_805);
nand U914 (N_914,In_1833,In_1022);
xor U915 (N_915,In_844,In_4936);
xor U916 (N_916,In_982,In_2716);
xor U917 (N_917,In_553,In_4776);
nand U918 (N_918,In_175,In_4655);
or U919 (N_919,In_3132,In_1411);
nand U920 (N_920,In_2535,In_3703);
nor U921 (N_921,In_4373,In_1923);
and U922 (N_922,In_790,In_758);
nor U923 (N_923,In_1935,In_1194);
or U924 (N_924,In_784,In_920);
xor U925 (N_925,In_2767,In_890);
nand U926 (N_926,In_188,In_4542);
and U927 (N_927,In_617,In_804);
or U928 (N_928,In_3626,In_4793);
nand U929 (N_929,In_601,In_3907);
xor U930 (N_930,In_1527,In_3095);
nand U931 (N_931,In_2392,In_4077);
xnor U932 (N_932,In_871,In_2304);
and U933 (N_933,In_3674,In_3553);
xor U934 (N_934,In_1403,In_429);
and U935 (N_935,In_87,In_4114);
nor U936 (N_936,In_3171,In_2049);
nor U937 (N_937,In_1469,In_2873);
nand U938 (N_938,In_2575,In_646);
or U939 (N_939,In_3773,In_2595);
and U940 (N_940,In_760,In_4768);
xnor U941 (N_941,In_4560,In_3595);
and U942 (N_942,In_4741,In_1507);
and U943 (N_943,In_2001,In_166);
and U944 (N_944,In_1349,In_101);
and U945 (N_945,In_1084,In_4436);
nand U946 (N_946,In_3236,In_3881);
and U947 (N_947,In_2428,In_4145);
and U948 (N_948,In_2999,In_261);
nor U949 (N_949,In_4634,In_4661);
nand U950 (N_950,In_4346,In_1302);
nand U951 (N_951,In_2021,In_3149);
nand U952 (N_952,In_3961,In_3377);
or U953 (N_953,In_3816,In_4592);
or U954 (N_954,In_968,In_688);
and U955 (N_955,In_3449,In_801);
and U956 (N_956,In_110,In_1316);
xor U957 (N_957,In_422,In_964);
and U958 (N_958,In_1368,In_182);
nor U959 (N_959,In_726,In_4593);
nor U960 (N_960,In_2628,In_3255);
xor U961 (N_961,In_2742,In_2376);
or U962 (N_962,In_4567,In_3);
xor U963 (N_963,In_955,In_1590);
nor U964 (N_964,In_378,In_4242);
and U965 (N_965,In_4352,In_3623);
nand U966 (N_966,In_1034,In_4761);
xor U967 (N_967,In_3925,In_1361);
xnor U968 (N_968,In_4859,In_4093);
or U969 (N_969,In_811,In_2323);
nand U970 (N_970,In_1165,In_257);
and U971 (N_971,In_2437,In_934);
and U972 (N_972,In_3376,In_2110);
nand U973 (N_973,In_146,In_589);
nand U974 (N_974,In_3719,In_120);
nor U975 (N_975,In_4287,In_854);
nand U976 (N_976,In_1785,In_3681);
nor U977 (N_977,In_1796,In_1898);
nor U978 (N_978,In_1109,In_1218);
xor U979 (N_979,In_2604,In_1085);
nand U980 (N_980,In_2465,In_1722);
nor U981 (N_981,In_2703,In_734);
or U982 (N_982,In_1453,In_3607);
xor U983 (N_983,In_1529,In_2135);
or U984 (N_984,In_4594,In_4379);
nor U985 (N_985,In_4745,In_2393);
xnor U986 (N_986,In_3013,In_428);
and U987 (N_987,In_4310,In_3758);
or U988 (N_988,In_3233,In_3573);
nand U989 (N_989,In_2521,In_772);
nor U990 (N_990,In_2236,In_2476);
xnor U991 (N_991,In_1245,In_3869);
nand U992 (N_992,In_55,In_4670);
nand U993 (N_993,In_2240,In_678);
nor U994 (N_994,In_916,In_4701);
xnor U995 (N_995,In_4123,In_3300);
nor U996 (N_996,In_798,In_3519);
or U997 (N_997,In_427,In_2700);
xnor U998 (N_998,In_290,In_1518);
nor U999 (N_999,In_4929,In_960);
or U1000 (N_1000,In_1800,In_3121);
nand U1001 (N_1001,In_4915,In_1829);
nor U1002 (N_1002,In_3746,In_4097);
xor U1003 (N_1003,In_2486,In_1424);
nor U1004 (N_1004,In_2773,In_5);
or U1005 (N_1005,In_4340,In_3020);
nand U1006 (N_1006,In_3261,In_2816);
or U1007 (N_1007,In_2315,In_3408);
nand U1008 (N_1008,In_4255,In_3701);
nor U1009 (N_1009,In_3308,In_1737);
nor U1010 (N_1010,In_2780,In_4376);
nor U1011 (N_1011,In_1758,In_3318);
and U1012 (N_1012,In_3828,In_4554);
nand U1013 (N_1013,In_3342,In_3837);
and U1014 (N_1014,In_3061,In_4983);
xor U1015 (N_1015,In_1651,In_4087);
nor U1016 (N_1016,In_4039,In_4819);
nand U1017 (N_1017,In_3076,In_2923);
or U1018 (N_1018,In_4845,In_4298);
xnor U1019 (N_1019,In_4437,In_4712);
nand U1020 (N_1020,In_2485,In_3852);
or U1021 (N_1021,In_2119,In_143);
nor U1022 (N_1022,In_555,In_3358);
nor U1023 (N_1023,In_4471,In_2386);
and U1024 (N_1024,In_3426,In_3063);
nand U1025 (N_1025,In_3669,In_2675);
and U1026 (N_1026,In_268,In_1475);
xor U1027 (N_1027,In_614,In_2981);
xnor U1028 (N_1028,In_1780,In_435);
nand U1029 (N_1029,In_685,In_1919);
xor U1030 (N_1030,In_4348,In_3332);
nor U1031 (N_1031,In_2140,In_1936);
or U1032 (N_1032,In_998,In_2166);
nand U1033 (N_1033,In_1143,In_2930);
nand U1034 (N_1034,In_3400,In_2998);
xor U1035 (N_1035,In_103,In_3665);
xor U1036 (N_1036,In_4119,In_2719);
nor U1037 (N_1037,In_4718,In_253);
xor U1038 (N_1038,In_1958,In_4813);
nor U1039 (N_1039,In_1997,In_2924);
nand U1040 (N_1040,In_693,In_2855);
xnor U1041 (N_1041,In_4796,In_1438);
xor U1042 (N_1042,In_4587,In_3796);
and U1043 (N_1043,In_165,In_1051);
nand U1044 (N_1044,In_4021,In_3547);
or U1045 (N_1045,In_3849,In_2869);
or U1046 (N_1046,In_2662,In_2007);
xor U1047 (N_1047,In_3981,In_2752);
nand U1048 (N_1048,In_533,In_942);
nor U1049 (N_1049,In_189,In_2309);
or U1050 (N_1050,In_2898,In_3911);
or U1051 (N_1051,In_2452,In_2934);
nand U1052 (N_1052,In_4642,In_4914);
nor U1053 (N_1053,In_2173,In_4314);
and U1054 (N_1054,In_445,In_4779);
nand U1055 (N_1055,In_2056,In_1891);
and U1056 (N_1056,In_4165,In_1169);
nand U1057 (N_1057,In_670,In_4546);
nand U1058 (N_1058,In_969,In_3606);
and U1059 (N_1059,In_452,In_2266);
xor U1060 (N_1060,In_3661,In_905);
nor U1061 (N_1061,In_2231,In_4061);
xnor U1062 (N_1062,In_4069,In_2909);
or U1063 (N_1063,In_1907,In_3084);
nand U1064 (N_1064,In_1784,In_3821);
nor U1065 (N_1065,In_3468,In_4990);
or U1066 (N_1066,In_831,In_3798);
and U1067 (N_1067,In_4168,In_2526);
and U1068 (N_1068,In_4433,In_1216);
and U1069 (N_1069,In_3153,In_4955);
nor U1070 (N_1070,In_3644,In_1640);
nor U1071 (N_1071,In_1953,In_1233);
or U1072 (N_1072,In_1445,In_3023);
nand U1073 (N_1073,In_1376,In_2242);
xnor U1074 (N_1074,In_327,In_3496);
and U1075 (N_1075,In_988,In_2028);
nand U1076 (N_1076,In_461,In_1234);
nor U1077 (N_1077,In_3917,In_720);
or U1078 (N_1078,In_4475,In_757);
or U1079 (N_1079,In_2280,In_4704);
or U1080 (N_1080,In_3964,In_2919);
xor U1081 (N_1081,In_1172,In_1877);
xnor U1082 (N_1082,In_2653,In_1952);
nor U1083 (N_1083,In_2345,In_4316);
nor U1084 (N_1084,In_1938,In_135);
nand U1085 (N_1085,In_2045,In_993);
xnor U1086 (N_1086,In_1966,In_4956);
or U1087 (N_1087,In_4231,In_1288);
or U1088 (N_1088,In_482,In_1560);
nand U1089 (N_1089,In_4390,In_1905);
nor U1090 (N_1090,In_3657,In_1965);
nand U1091 (N_1091,In_2715,In_2246);
or U1092 (N_1092,In_3813,In_4549);
xor U1093 (N_1093,In_2065,In_675);
xor U1094 (N_1094,In_3204,In_3190);
or U1095 (N_1095,In_2077,In_626);
xnor U1096 (N_1096,In_1587,In_1964);
nand U1097 (N_1097,In_2364,In_4311);
nor U1098 (N_1098,In_1449,In_1955);
nor U1099 (N_1099,In_2786,In_3545);
and U1100 (N_1100,In_765,In_3637);
and U1101 (N_1101,In_671,In_2146);
nor U1102 (N_1102,In_2705,In_1054);
and U1103 (N_1103,In_598,In_2298);
and U1104 (N_1104,In_4690,In_3456);
nor U1105 (N_1105,In_3311,In_4150);
nand U1106 (N_1106,In_2562,In_1270);
and U1107 (N_1107,In_3446,In_512);
xnor U1108 (N_1108,In_2275,In_996);
and U1109 (N_1109,In_4158,In_2784);
and U1110 (N_1110,In_1634,In_1200);
xor U1111 (N_1111,In_1170,In_4412);
or U1112 (N_1112,In_343,In_3322);
xor U1113 (N_1113,In_1986,In_3137);
and U1114 (N_1114,In_4175,In_4101);
xor U1115 (N_1115,In_1713,In_3000);
nand U1116 (N_1116,In_285,In_4777);
nor U1117 (N_1117,In_1866,In_4260);
or U1118 (N_1118,In_3770,In_2843);
nand U1119 (N_1119,In_1972,In_122);
or U1120 (N_1120,In_3579,In_379);
or U1121 (N_1121,In_3938,In_1095);
xnor U1122 (N_1122,In_4692,In_3831);
and U1123 (N_1123,In_4195,In_3957);
and U1124 (N_1124,In_3531,In_4493);
and U1125 (N_1125,In_1498,In_4699);
xnor U1126 (N_1126,In_1338,In_262);
nand U1127 (N_1127,In_3505,In_2557);
and U1128 (N_1128,In_4403,In_859);
or U1129 (N_1129,In_4275,In_1983);
and U1130 (N_1130,In_179,In_4902);
nor U1131 (N_1131,In_3031,In_4217);
nand U1132 (N_1132,In_3437,In_304);
nor U1133 (N_1133,In_3325,In_4555);
nor U1134 (N_1134,In_3952,In_2420);
and U1135 (N_1135,In_3265,In_2130);
xor U1136 (N_1136,In_1147,In_4089);
nand U1137 (N_1137,In_3477,In_2837);
nand U1138 (N_1138,In_4619,In_3447);
xor U1139 (N_1139,In_4094,In_150);
xor U1140 (N_1140,In_4138,In_1502);
nor U1141 (N_1141,In_1112,In_1323);
or U1142 (N_1142,In_2992,In_535);
nand U1143 (N_1143,In_3900,In_368);
or U1144 (N_1144,In_1823,In_1837);
nand U1145 (N_1145,In_4183,In_1711);
or U1146 (N_1146,In_2737,In_4707);
nand U1147 (N_1147,In_279,In_3374);
and U1148 (N_1148,In_733,In_1561);
nand U1149 (N_1149,In_2198,In_2713);
and U1150 (N_1150,In_794,In_2947);
nor U1151 (N_1151,In_1976,In_2013);
and U1152 (N_1152,In_2798,In_3799);
or U1153 (N_1153,In_3908,In_3192);
nand U1154 (N_1154,In_2819,In_4228);
nor U1155 (N_1155,In_1363,In_4803);
or U1156 (N_1156,In_2890,In_331);
xor U1157 (N_1157,In_3041,In_1668);
or U1158 (N_1158,In_1314,In_544);
xor U1159 (N_1159,In_2172,In_3253);
xor U1160 (N_1160,In_3919,In_1137);
and U1161 (N_1161,In_1646,In_3651);
xnor U1162 (N_1162,In_1260,In_92);
nor U1163 (N_1163,In_4728,In_3527);
nand U1164 (N_1164,In_2966,In_2439);
nor U1165 (N_1165,In_4810,In_3897);
xnor U1166 (N_1166,In_4214,In_16);
and U1167 (N_1167,In_3776,In_2347);
nor U1168 (N_1168,In_2155,In_3231);
nand U1169 (N_1169,In_436,In_4946);
nor U1170 (N_1170,In_2558,In_4576);
or U1171 (N_1171,In_4124,In_3421);
nor U1172 (N_1172,In_4781,In_2127);
and U1173 (N_1173,In_1369,In_115);
xor U1174 (N_1174,In_4591,In_1082);
and U1175 (N_1175,In_1146,In_3843);
or U1176 (N_1176,In_157,In_3475);
xnor U1177 (N_1177,In_486,In_1846);
or U1178 (N_1178,In_4828,In_4019);
xnor U1179 (N_1179,In_4015,In_4122);
xor U1180 (N_1180,In_2497,In_1960);
nand U1181 (N_1181,In_3001,In_3683);
nor U1182 (N_1182,In_3906,In_233);
or U1183 (N_1183,In_4691,In_4186);
nor U1184 (N_1184,In_2566,In_2911);
or U1185 (N_1185,In_1756,In_1246);
and U1186 (N_1186,In_423,In_3762);
nor U1187 (N_1187,In_25,In_2570);
or U1188 (N_1188,In_653,In_198);
and U1189 (N_1189,In_123,In_2457);
xnor U1190 (N_1190,In_85,In_3998);
xnor U1191 (N_1191,In_2762,In_2320);
xor U1192 (N_1192,In_1439,In_2832);
nor U1193 (N_1193,In_763,In_1612);
nor U1194 (N_1194,In_2456,In_1117);
or U1195 (N_1195,In_46,In_3777);
or U1196 (N_1196,In_3535,In_1456);
and U1197 (N_1197,In_3118,In_1418);
nor U1198 (N_1198,In_951,In_1395);
xnor U1199 (N_1199,In_4030,In_3238);
xnor U1200 (N_1200,In_3324,In_2917);
nand U1201 (N_1201,In_3454,In_4603);
nor U1202 (N_1202,In_2449,In_3765);
nand U1203 (N_1203,In_3345,In_2033);
nor U1204 (N_1204,In_4249,In_3888);
nor U1205 (N_1205,In_413,In_4791);
or U1206 (N_1206,In_234,In_484);
nand U1207 (N_1207,In_1880,In_481);
xor U1208 (N_1208,In_3729,In_2783);
and U1209 (N_1209,In_3836,In_1281);
or U1210 (N_1210,In_2694,In_7);
and U1211 (N_1211,In_2104,In_1504);
and U1212 (N_1212,In_4730,In_3285);
and U1213 (N_1213,In_3431,In_3915);
nand U1214 (N_1214,In_739,In_288);
and U1215 (N_1215,In_2458,In_3444);
nor U1216 (N_1216,In_2426,In_320);
or U1217 (N_1217,In_2959,In_4336);
nor U1218 (N_1218,In_272,In_3523);
xor U1219 (N_1219,In_4550,In_639);
nand U1220 (N_1220,In_1258,In_2024);
nand U1221 (N_1221,In_4856,In_4697);
xor U1222 (N_1222,In_708,In_1239);
xor U1223 (N_1223,In_1751,In_3842);
or U1224 (N_1224,In_124,In_2398);
xor U1225 (N_1225,In_2669,In_4644);
and U1226 (N_1226,In_4108,In_538);
and U1227 (N_1227,In_4879,In_1540);
xor U1228 (N_1228,In_701,In_2615);
nor U1229 (N_1229,In_2724,In_269);
nand U1230 (N_1230,In_707,In_895);
and U1231 (N_1231,In_2060,In_2651);
and U1232 (N_1232,In_1121,In_3196);
nor U1233 (N_1233,In_4895,In_1360);
nor U1234 (N_1234,In_4532,In_2978);
nand U1235 (N_1235,In_2748,In_2047);
or U1236 (N_1236,In_216,In_228);
xnor U1237 (N_1237,In_4823,In_3699);
and U1238 (N_1238,In_1617,In_2531);
nor U1239 (N_1239,In_4966,In_4635);
xor U1240 (N_1240,In_4965,In_1191);
or U1241 (N_1241,In_1654,In_4623);
or U1242 (N_1242,In_3960,In_1884);
nor U1243 (N_1243,In_936,In_2015);
and U1244 (N_1244,In_1865,In_3284);
and U1245 (N_1245,In_4640,In_2831);
and U1246 (N_1246,In_4633,In_4713);
nand U1247 (N_1247,In_730,In_184);
and U1248 (N_1248,In_3788,In_1754);
or U1249 (N_1249,In_4191,In_3648);
and U1250 (N_1250,In_618,In_1779);
nor U1251 (N_1251,In_4763,In_3337);
nor U1252 (N_1252,In_2193,In_981);
nor U1253 (N_1253,In_1573,In_4187);
and U1254 (N_1254,In_561,In_1480);
nand U1255 (N_1255,In_4090,In_3503);
nand U1256 (N_1256,In_4363,In_4488);
nor U1257 (N_1257,In_4799,In_357);
nor U1258 (N_1258,In_3899,In_4107);
xor U1259 (N_1259,In_2957,In_2391);
or U1260 (N_1260,In_2903,In_3951);
or U1261 (N_1261,In_1184,In_4451);
or U1262 (N_1262,In_821,In_4520);
and U1263 (N_1263,In_1024,In_409);
xnor U1264 (N_1264,In_319,In_520);
and U1265 (N_1265,In_3247,In_1324);
nor U1266 (N_1266,In_3520,In_3583);
xor U1267 (N_1267,In_1486,In_4209);
nor U1268 (N_1268,In_3319,In_1838);
and U1269 (N_1269,In_1254,In_3155);
nand U1270 (N_1270,In_4028,In_2938);
nor U1271 (N_1271,In_3538,In_2645);
nand U1272 (N_1272,In_2976,In_4345);
xor U1273 (N_1273,In_3775,In_2093);
and U1274 (N_1274,In_2734,In_3450);
nand U1275 (N_1275,In_4431,In_2278);
or U1276 (N_1276,In_649,In_3584);
nand U1277 (N_1277,In_4443,In_1940);
nand U1278 (N_1278,In_1221,In_3385);
and U1279 (N_1279,In_839,In_2164);
and U1280 (N_1280,In_4752,In_1455);
and U1281 (N_1281,In_4616,In_4274);
nor U1282 (N_1282,In_3610,In_802);
and U1283 (N_1283,In_4525,In_4877);
or U1284 (N_1284,In_313,In_1046);
or U1285 (N_1285,In_2895,In_2527);
or U1286 (N_1286,In_163,In_1637);
nor U1287 (N_1287,In_2511,In_545);
xnor U1288 (N_1288,In_735,In_148);
nand U1289 (N_1289,In_3146,In_1398);
or U1290 (N_1290,In_1183,In_673);
xnor U1291 (N_1291,In_3109,In_1885);
and U1292 (N_1292,In_1762,In_353);
nand U1293 (N_1293,In_2702,In_3638);
nand U1294 (N_1294,In_3609,In_3602);
and U1295 (N_1295,In_1738,In_2117);
xor U1296 (N_1296,In_2005,In_2228);
and U1297 (N_1297,In_3605,In_82);
and U1298 (N_1298,In_1171,In_340);
and U1299 (N_1299,In_2106,In_4359);
or U1300 (N_1300,In_4553,In_2388);
nand U1301 (N_1301,In_465,In_3760);
or U1302 (N_1302,In_3343,In_2943);
nor U1303 (N_1303,In_1575,In_2529);
nand U1304 (N_1304,In_3158,In_3855);
nand U1305 (N_1305,In_1222,In_717);
nand U1306 (N_1306,In_3890,In_142);
xnor U1307 (N_1307,In_851,In_3336);
nor U1308 (N_1308,In_2951,In_4653);
xor U1309 (N_1309,In_13,In_1950);
nor U1310 (N_1310,In_2962,In_3143);
nor U1311 (N_1311,In_1204,In_2207);
xnor U1312 (N_1312,In_3734,In_4556);
or U1313 (N_1313,In_3740,In_2002);
xor U1314 (N_1314,In_3747,In_344);
nor U1315 (N_1315,In_3660,In_3916);
or U1316 (N_1316,In_4065,In_4688);
nor U1317 (N_1317,In_1788,In_4916);
nor U1318 (N_1318,In_4935,In_161);
xnor U1319 (N_1319,In_3428,In_1795);
xnor U1320 (N_1320,In_3947,In_3306);
or U1321 (N_1321,In_816,In_3310);
and U1322 (N_1322,In_3871,In_1459);
nor U1323 (N_1323,In_1613,In_3802);
nor U1324 (N_1324,In_2545,In_4787);
or U1325 (N_1325,In_1703,In_276);
or U1326 (N_1326,In_1511,In_1767);
and U1327 (N_1327,In_3780,In_2410);
or U1328 (N_1328,In_2623,In_2550);
and U1329 (N_1329,In_4672,In_4987);
xor U1330 (N_1330,In_1257,In_4121);
nor U1331 (N_1331,In_4920,In_2753);
nand U1332 (N_1332,In_3774,In_1633);
xnor U1333 (N_1333,In_3228,In_1100);
nor U1334 (N_1334,In_1791,In_3048);
nand U1335 (N_1335,In_501,In_4422);
xor U1336 (N_1336,In_443,In_3370);
nor U1337 (N_1337,In_622,In_270);
xnor U1338 (N_1338,In_149,In_4283);
xnor U1339 (N_1339,In_197,In_267);
nand U1340 (N_1340,In_3094,In_2058);
nor U1341 (N_1341,In_2925,In_1230);
nand U1342 (N_1342,In_3874,In_1196);
nor U1343 (N_1343,In_1598,In_4840);
nor U1344 (N_1344,In_2637,In_774);
or U1345 (N_1345,In_2380,In_1008);
and U1346 (N_1346,In_3474,In_4042);
nor U1347 (N_1347,In_4074,In_2477);
nand U1348 (N_1348,In_4989,In_1138);
xnor U1349 (N_1349,In_209,In_4890);
nand U1350 (N_1350,In_4643,In_447);
xor U1351 (N_1351,In_725,In_560);
nand U1352 (N_1352,In_917,In_4759);
xnor U1353 (N_1353,In_350,In_2105);
xnor U1354 (N_1354,In_4666,In_3051);
and U1355 (N_1355,In_3053,In_820);
and U1356 (N_1356,In_328,In_4849);
or U1357 (N_1357,In_898,In_4982);
nand U1358 (N_1358,In_1572,In_4689);
and U1359 (N_1359,In_1740,In_1495);
or U1360 (N_1360,In_4651,In_2296);
nand U1361 (N_1361,In_3245,In_1190);
nor U1362 (N_1362,In_76,In_2226);
or U1363 (N_1363,In_4943,In_709);
nand U1364 (N_1364,In_1107,In_1725);
xor U1365 (N_1365,In_858,In_828);
and U1366 (N_1366,In_751,In_1064);
xor U1367 (N_1367,In_4618,In_3694);
and U1368 (N_1368,In_2436,In_4271);
or U1369 (N_1369,In_2897,In_864);
and U1370 (N_1370,In_4538,In_660);
nor U1371 (N_1371,In_3116,In_239);
nor U1372 (N_1372,In_3809,In_168);
xnor U1373 (N_1373,In_946,In_3278);
nor U1374 (N_1374,In_4671,In_4924);
and U1375 (N_1375,In_2283,In_3867);
xor U1376 (N_1376,In_3655,In_2760);
xnor U1377 (N_1377,In_1032,In_2471);
nand U1378 (N_1378,In_1454,In_738);
and U1379 (N_1379,In_1727,In_519);
xnor U1380 (N_1380,In_1820,In_1255);
nand U1381 (N_1381,In_3100,In_3364);
nand U1382 (N_1382,In_2150,In_4864);
nand U1383 (N_1383,In_1328,In_4686);
or U1384 (N_1384,In_3518,In_4157);
nand U1385 (N_1385,In_4872,In_3170);
or U1386 (N_1386,In_1609,In_3592);
or U1387 (N_1387,In_940,In_2203);
or U1388 (N_1388,In_3522,In_4017);
and U1389 (N_1389,In_4663,In_4378);
xnor U1390 (N_1390,In_2697,In_1766);
or U1391 (N_1391,In_1942,In_440);
and U1392 (N_1392,In_3712,In_4380);
nor U1393 (N_1393,In_918,In_1792);
or U1394 (N_1394,In_4344,In_4257);
nand U1395 (N_1395,In_3676,In_1059);
or U1396 (N_1396,In_297,In_4243);
nand U1397 (N_1397,In_3096,In_3624);
and U1398 (N_1398,In_4548,In_1743);
nor U1399 (N_1399,In_1279,In_2357);
nand U1400 (N_1400,In_997,In_4597);
and U1401 (N_1401,In_4246,In_681);
and U1402 (N_1402,In_1570,In_1489);
or U1403 (N_1403,In_3062,In_4485);
xnor U1404 (N_1404,In_2920,In_3515);
nand U1405 (N_1405,In_3185,In_2886);
nand U1406 (N_1406,In_3652,In_3225);
nand U1407 (N_1407,In_454,In_1684);
xnor U1408 (N_1408,In_679,In_3575);
xor U1409 (N_1409,In_3965,In_1251);
xnor U1410 (N_1410,In_3058,In_2414);
and U1411 (N_1411,In_1706,In_4295);
xnor U1412 (N_1412,In_3383,In_3673);
nand U1413 (N_1413,In_412,In_4585);
xnor U1414 (N_1414,In_1888,In_1917);
or U1415 (N_1415,In_1099,In_1828);
nand U1416 (N_1416,In_2967,In_4590);
or U1417 (N_1417,In_322,In_127);
xnor U1418 (N_1418,In_4693,In_4474);
nand U1419 (N_1419,In_2337,In_346);
nor U1420 (N_1420,In_464,In_2249);
nor U1421 (N_1421,In_2757,In_114);
nand U1422 (N_1422,In_3614,In_1310);
nand U1423 (N_1423,In_2755,In_4481);
or U1424 (N_1424,In_2500,In_1096);
xor U1425 (N_1425,In_4180,In_1528);
or U1426 (N_1426,In_1521,In_1914);
and U1427 (N_1427,In_2196,In_2460);
xor U1428 (N_1428,In_687,In_1932);
nor U1429 (N_1429,In_2594,In_2233);
xor U1430 (N_1430,In_347,In_532);
nand U1431 (N_1431,In_2480,In_3640);
xor U1432 (N_1432,In_818,In_2830);
or U1433 (N_1433,In_973,In_1626);
nand U1434 (N_1434,In_2932,In_976);
or U1435 (N_1435,In_98,In_3992);
nand U1436 (N_1436,In_3433,In_3670);
nand U1437 (N_1437,In_4561,In_4473);
and U1438 (N_1438,In_2597,In_1817);
nor U1439 (N_1439,In_4420,In_4681);
nand U1440 (N_1440,In_3550,In_4899);
or U1441 (N_1441,In_2589,In_2123);
and U1442 (N_1442,In_2401,In_2461);
nand U1443 (N_1443,In_3427,In_4769);
and U1444 (N_1444,In_4847,In_3830);
and U1445 (N_1445,In_3059,In_21);
and U1446 (N_1446,In_668,In_1709);
and U1447 (N_1447,In_4207,In_2029);
or U1448 (N_1448,In_4680,In_4154);
or U1449 (N_1449,In_4280,In_4612);
and U1450 (N_1450,In_3178,In_4423);
nand U1451 (N_1451,In_770,In_957);
nor U1452 (N_1452,In_592,In_1444);
nand U1453 (N_1453,In_202,In_2365);
xor U1454 (N_1454,In_4288,In_2668);
nor U1455 (N_1455,In_3543,In_728);
nand U1456 (N_1456,In_1882,In_3207);
xnor U1457 (N_1457,In_4055,In_4080);
nand U1458 (N_1458,In_3999,In_2865);
and U1459 (N_1459,In_4714,In_4539);
xor U1460 (N_1460,In_1217,In_3590);
xor U1461 (N_1461,In_1676,In_1660);
or U1462 (N_1462,In_855,In_787);
nor U1463 (N_1463,In_4224,In_2852);
xor U1464 (N_1464,In_1944,In_1397);
nand U1465 (N_1465,In_903,In_4909);
xnor U1466 (N_1466,In_2876,In_2142);
nor U1467 (N_1467,In_2067,In_3634);
nand U1468 (N_1468,In_1101,In_106);
and U1469 (N_1469,In_1400,In_3576);
nor U1470 (N_1470,In_334,In_2853);
or U1471 (N_1471,In_1508,In_4116);
xor U1472 (N_1472,In_796,In_3077);
nand U1473 (N_1473,In_3334,In_3448);
nand U1474 (N_1474,In_540,In_1913);
xor U1475 (N_1475,In_3944,In_1667);
nor U1476 (N_1476,In_2186,In_4515);
and U1477 (N_1477,In_4050,In_4239);
nand U1478 (N_1478,In_1435,In_63);
nor U1479 (N_1479,In_2438,In_2940);
nor U1480 (N_1480,In_4968,In_2958);
nor U1481 (N_1481,In_252,In_2534);
and U1482 (N_1482,In_1906,In_4100);
xor U1483 (N_1483,In_716,In_1018);
nand U1484 (N_1484,In_1392,In_1105);
or U1485 (N_1485,In_1,In_1467);
xnor U1486 (N_1486,In_2910,In_4838);
nand U1487 (N_1487,In_4758,In_4043);
and U1488 (N_1488,In_3940,In_1139);
and U1489 (N_1489,In_4628,In_3440);
and U1490 (N_1490,In_2599,In_737);
or U1491 (N_1491,In_4638,In_2883);
nor U1492 (N_1492,In_1496,In_3340);
xnor U1493 (N_1493,In_3985,In_3812);
nand U1494 (N_1494,In_1875,In_2660);
xor U1495 (N_1495,In_493,In_4705);
and U1496 (N_1496,In_947,In_3299);
nor U1497 (N_1497,In_2522,In_3525);
nand U1498 (N_1498,In_490,In_3490);
xnor U1499 (N_1499,In_3181,In_1133);
xor U1500 (N_1500,In_4596,In_1207);
or U1501 (N_1501,In_4139,In_1130);
xnor U1502 (N_1502,In_572,In_995);
and U1503 (N_1503,In_985,In_2044);
nor U1504 (N_1504,In_4926,In_3815);
nor U1505 (N_1505,In_2284,In_4881);
nor U1506 (N_1506,In_909,In_2546);
nor U1507 (N_1507,In_2530,In_4082);
nand U1508 (N_1508,In_2872,In_3367);
or U1509 (N_1509,In_2600,In_463);
or U1510 (N_1510,In_1175,In_444);
or U1511 (N_1511,In_3870,In_999);
and U1512 (N_1512,In_4308,In_3817);
xnor U1513 (N_1513,In_3577,In_3210);
xor U1514 (N_1514,In_176,In_4222);
nand U1515 (N_1515,In_89,In_661);
xor U1516 (N_1516,In_1153,In_1450);
nor U1517 (N_1517,In_710,In_4062);
xnor U1518 (N_1518,In_3234,In_4528);
and U1519 (N_1519,In_1180,In_2158);
or U1520 (N_1520,In_4147,In_1980);
nor U1521 (N_1521,In_3883,In_2996);
and U1522 (N_1522,In_1201,In_1863);
or U1523 (N_1523,In_3790,In_650);
nor U1524 (N_1524,In_2850,In_2143);
nand U1525 (N_1525,In_1250,In_1019);
or U1526 (N_1526,In_3572,In_1571);
nand U1527 (N_1527,In_2281,In_3771);
and U1528 (N_1528,In_4385,In_2936);
nand U1529 (N_1529,In_1209,In_3555);
xor U1530 (N_1530,In_536,In_4190);
or U1531 (N_1531,In_958,In_2484);
nand U1532 (N_1532,In_3641,In_282);
nand U1533 (N_1533,In_1975,In_1516);
nand U1534 (N_1534,In_2987,In_3333);
or U1535 (N_1535,In_4674,In_132);
or U1536 (N_1536,In_1226,In_1967);
and U1537 (N_1537,In_1344,In_3174);
nand U1538 (N_1538,In_4472,In_1506);
xnor U1539 (N_1539,In_2229,In_3186);
or U1540 (N_1540,In_2063,In_3470);
xor U1541 (N_1541,In_1664,In_2583);
or U1542 (N_1542,In_2241,In_514);
nor U1543 (N_1543,In_3281,In_2394);
nand U1544 (N_1544,In_4277,In_3541);
or U1545 (N_1545,In_1081,In_4625);
nor U1546 (N_1546,In_3835,In_1087);
and U1547 (N_1547,In_3993,In_3949);
or U1548 (N_1548,In_3384,In_1321);
or U1549 (N_1549,In_4370,In_2648);
xor U1550 (N_1550,In_2342,In_3420);
xnor U1551 (N_1551,In_2455,In_1355);
nor U1552 (N_1552,In_933,In_1503);
nand U1553 (N_1553,In_1238,In_1721);
nor U1554 (N_1554,In_1061,In_4783);
nand U1555 (N_1555,In_3787,In_848);
nand U1556 (N_1556,In_278,In_3857);
nand U1557 (N_1557,In_117,In_4216);
and U1558 (N_1558,In_0,In_928);
or U1559 (N_1559,In_2984,In_4756);
nand U1560 (N_1560,In_3147,In_2768);
or U1561 (N_1561,In_941,In_2081);
xor U1562 (N_1562,In_2004,In_4771);
or U1563 (N_1563,In_2182,In_2210);
xnor U1564 (N_1564,In_834,In_2749);
xor U1565 (N_1565,In_3726,In_1734);
or U1566 (N_1566,In_18,In_2584);
nand U1567 (N_1567,In_3169,In_1661);
and U1568 (N_1568,In_2262,In_3052);
and U1569 (N_1569,In_3120,In_3653);
or U1570 (N_1570,In_4711,In_585);
nand U1571 (N_1571,In_4374,In_2138);
xor U1572 (N_1572,In_1308,In_2854);
and U1573 (N_1573,In_3239,In_836);
nand U1574 (N_1574,In_3713,In_1317);
nand U1575 (N_1575,In_3485,In_4497);
xor U1576 (N_1576,In_2188,In_4918);
xnor U1577 (N_1577,In_2163,In_79);
nand U1578 (N_1578,In_4967,In_523);
xor U1579 (N_1579,In_4153,In_118);
or U1580 (N_1580,In_1834,In_870);
nand U1581 (N_1581,In_1460,In_3948);
xor U1582 (N_1582,In_2019,In_194);
xor U1583 (N_1583,In_3414,In_3702);
or U1584 (N_1584,In_1825,In_3819);
xnor U1585 (N_1585,In_3424,In_1663);
or U1586 (N_1586,In_4325,In_2577);
or U1587 (N_1587,In_867,In_4259);
nand U1588 (N_1588,In_2718,In_66);
nor U1589 (N_1589,In_3945,In_3355);
and U1590 (N_1590,In_2372,In_1581);
and U1591 (N_1591,In_2596,In_3894);
nand U1592 (N_1592,In_539,In_956);
or U1593 (N_1593,In_692,In_2567);
and U1594 (N_1594,In_3806,In_2801);
and U1595 (N_1595,In_1876,In_1608);
and U1596 (N_1596,In_1399,In_554);
nand U1597 (N_1597,In_4537,In_3675);
nand U1598 (N_1598,In_213,In_360);
and U1599 (N_1599,In_130,In_2794);
nand U1600 (N_1600,In_393,In_4928);
or U1601 (N_1601,In_4459,In_1319);
nand U1602 (N_1602,In_3534,In_2841);
or U1603 (N_1603,In_1492,In_562);
nand U1604 (N_1604,In_2688,In_4041);
nand U1605 (N_1605,In_3642,In_2079);
xnor U1606 (N_1606,In_3668,In_1852);
nand U1607 (N_1607,In_2706,In_810);
xnor U1608 (N_1608,In_3246,In_2273);
xor U1609 (N_1609,In_1776,In_141);
and U1610 (N_1610,In_846,In_1001);
nand U1611 (N_1611,In_1690,In_2711);
and U1612 (N_1612,In_4004,In_2614);
nand U1613 (N_1613,In_1286,In_3394);
nor U1614 (N_1614,In_4852,In_563);
xor U1615 (N_1615,In_3753,In_3088);
and U1616 (N_1616,In_2252,In_1000);
xor U1617 (N_1617,In_2851,In_963);
xor U1618 (N_1618,In_902,In_3688);
or U1619 (N_1619,In_2148,In_2636);
and U1620 (N_1620,In_1351,In_4611);
or U1621 (N_1621,In_22,In_1681);
nor U1622 (N_1622,In_4236,In_2607);
or U1623 (N_1623,In_210,In_663);
or U1624 (N_1624,In_508,In_2692);
nor U1625 (N_1625,In_823,In_1214);
nor U1626 (N_1626,In_2840,In_483);
or U1627 (N_1627,In_158,In_119);
or U1628 (N_1628,In_4086,In_4120);
or U1629 (N_1629,In_3277,In_528);
or U1630 (N_1630,In_71,In_3124);
or U1631 (N_1631,In_1384,In_263);
and U1632 (N_1632,In_3298,In_4789);
xor U1633 (N_1633,In_4573,In_1394);
or U1634 (N_1634,In_3457,In_1013);
nand U1635 (N_1635,In_1428,In_4814);
nand U1636 (N_1636,In_3179,In_2548);
nor U1637 (N_1637,In_2363,In_1472);
nor U1638 (N_1638,In_2776,In_2743);
and U1639 (N_1639,In_1223,In_3620);
nor U1640 (N_1640,In_1995,In_223);
nor U1641 (N_1641,In_3829,In_4911);
nand U1642 (N_1642,In_1694,In_3983);
nor U1643 (N_1643,In_4620,In_291);
xor U1644 (N_1644,In_4827,In_4016);
xnor U1645 (N_1645,In_1038,In_1240);
or U1646 (N_1646,In_2086,In_4921);
nor U1647 (N_1647,In_2381,In_980);
nor U1648 (N_1648,In_2812,In_2560);
nand U1649 (N_1649,In_3664,In_3388);
nor U1650 (N_1650,In_2667,In_1451);
xor U1651 (N_1651,In_2835,In_4888);
nand U1652 (N_1652,In_2128,In_2332);
nand U1653 (N_1653,In_4409,In_433);
and U1654 (N_1654,In_581,In_4930);
nor U1655 (N_1655,In_3984,In_2680);
xor U1656 (N_1656,In_1512,In_3803);
nor U1657 (N_1657,In_800,In_2157);
nand U1658 (N_1658,In_2634,In_3677);
and U1659 (N_1659,In_4447,In_3996);
and U1660 (N_1660,In_4113,In_4675);
or U1661 (N_1661,In_1149,In_2973);
xor U1662 (N_1662,In_1482,In_3419);
and U1663 (N_1663,In_2617,In_3223);
nand U1664 (N_1664,In_3920,In_3293);
xnor U1665 (N_1665,In_4388,In_332);
xnor U1666 (N_1666,In_4115,In_975);
or U1667 (N_1667,In_4442,In_2533);
and U1668 (N_1668,In_4491,In_4659);
nand U1669 (N_1669,In_4544,In_2723);
xor U1670 (N_1670,In_662,In_2183);
xnor U1671 (N_1671,In_4533,In_2779);
nor U1672 (N_1672,In_2328,In_4424);
or U1673 (N_1673,In_4461,In_1860);
and U1674 (N_1674,In_3593,In_2014);
nor U1675 (N_1675,In_4091,In_2199);
nand U1676 (N_1676,In_2385,In_1371);
and U1677 (N_1677,In_1687,In_3130);
or U1678 (N_1678,In_1538,In_4757);
or U1679 (N_1679,In_1073,In_3386);
or U1680 (N_1680,In_138,In_684);
nor U1681 (N_1681,In_3347,In_2169);
nand U1682 (N_1682,In_4647,In_3832);
or U1683 (N_1683,In_2206,In_694);
nor U1684 (N_1684,In_476,In_808);
or U1685 (N_1685,In_4240,In_3240);
or U1686 (N_1686,In_511,In_1670);
and U1687 (N_1687,In_509,In_4027);
nand U1688 (N_1688,In_1386,In_3429);
and U1689 (N_1689,In_3692,In_4067);
xnor U1690 (N_1690,In_2549,In_3647);
nor U1691 (N_1691,In_3047,In_633);
and U1692 (N_1692,In_1593,In_3011);
and U1693 (N_1693,In_1429,In_4449);
nor U1694 (N_1694,In_3218,In_3741);
xor U1695 (N_1695,In_1563,In_4932);
or U1696 (N_1696,In_1437,In_2400);
or U1697 (N_1697,In_1192,In_576);
and U1698 (N_1698,In_4290,In_2813);
xor U1699 (N_1699,In_3580,In_425);
xor U1700 (N_1700,In_2131,In_1273);
xor U1701 (N_1701,In_4727,In_1199);
and U1702 (N_1702,In_2856,In_2792);
nand U1703 (N_1703,In_4136,In_4448);
and U1704 (N_1704,In_4959,In_2237);
xor U1705 (N_1705,In_564,In_1849);
xnor U1706 (N_1706,In_2574,In_1102);
xor U1707 (N_1707,In_4577,In_2443);
nor U1708 (N_1708,In_1039,In_2445);
nor U1709 (N_1709,In_978,In_595);
xnor U1710 (N_1710,In_2683,In_1016);
and U1711 (N_1711,In_4624,In_1313);
and U1712 (N_1712,In_2699,In_2046);
nor U1713 (N_1713,In_1746,In_4884);
nor U1714 (N_1714,In_30,In_326);
or U1715 (N_1715,In_4129,In_1452);
nor U1716 (N_1716,In_807,In_1070);
or U1717 (N_1717,In_4817,In_4570);
xnor U1718 (N_1718,In_4251,In_1315);
nand U1719 (N_1719,In_3176,In_4563);
xnor U1720 (N_1720,In_2475,In_696);
nor U1721 (N_1721,In_2405,In_4398);
nand U1722 (N_1722,In_1909,In_125);
nand U1723 (N_1723,In_3145,In_4070);
nor U1724 (N_1724,In_4441,In_4408);
nand U1725 (N_1725,In_2451,In_4428);
nand U1726 (N_1726,In_652,In_3886);
nor U1727 (N_1727,In_3291,In_4595);
or U1728 (N_1728,In_1029,In_2256);
or U1729 (N_1729,In_1350,In_635);
nor U1730 (N_1730,In_884,In_1356);
or U1731 (N_1731,In_2139,In_1477);
or U1732 (N_1732,In_352,In_2581);
nand U1733 (N_1733,In_193,In_3565);
nor U1734 (N_1734,In_2666,In_1501);
nor U1735 (N_1735,In_2089,In_2912);
xnor U1736 (N_1736,In_2220,In_1232);
or U1737 (N_1737,In_274,In_2568);
and U1738 (N_1738,In_4988,In_2944);
and U1739 (N_1739,In_1259,In_237);
and U1740 (N_1740,In_3707,In_1097);
xnor U1741 (N_1741,In_1645,In_1385);
xor U1742 (N_1742,In_1631,In_1842);
xor U1743 (N_1743,In_4893,In_2541);
nand U1744 (N_1744,In_2879,In_3779);
xnor U1745 (N_1745,In_1777,In_3510);
nor U1746 (N_1746,In_3349,In_1337);
xor U1747 (N_1747,In_2416,In_2553);
or U1748 (N_1748,In_2795,In_4198);
xnor U1749 (N_1749,In_4400,In_1543);
xnor U1750 (N_1750,In_2227,In_4738);
and U1751 (N_1751,In_2325,In_2382);
nor U1752 (N_1752,In_1994,In_866);
and U1753 (N_1753,In_4425,In_2043);
nor U1754 (N_1754,In_3969,In_4748);
or U1755 (N_1755,In_4478,In_912);
or U1756 (N_1756,In_791,In_4588);
and U1757 (N_1757,In_1601,In_3287);
nand U1758 (N_1758,In_4022,In_1760);
nand U1759 (N_1759,In_3248,In_762);
nor U1760 (N_1760,In_1930,In_4056);
xnor U1761 (N_1761,In_1525,In_2670);
and U1762 (N_1762,In_1301,In_4974);
and U1763 (N_1763,In_3797,In_49);
nand U1764 (N_1764,In_4392,In_2217);
nand U1765 (N_1765,In_2263,In_10);
xnor U1766 (N_1766,In_4721,In_2035);
nand U1767 (N_1767,In_3025,In_1591);
or U1768 (N_1768,In_3599,In_2975);
or U1769 (N_1769,In_1330,In_4518);
nor U1770 (N_1770,In_4476,In_1291);
nor U1771 (N_1771,In_1500,In_3718);
nand U1772 (N_1772,In_315,In_3407);
nand U1773 (N_1773,In_2088,In_1092);
nand U1774 (N_1774,In_4607,In_4854);
or U1775 (N_1775,In_214,In_4241);
nand U1776 (N_1776,In_542,In_3036);
and U1777 (N_1777,In_2307,In_2707);
or U1778 (N_1778,In_28,In_1644);
xnor U1779 (N_1779,In_4387,In_3164);
nor U1780 (N_1780,In_1824,In_3684);
or U1781 (N_1781,In_4702,In_4963);
and U1782 (N_1782,In_2310,In_1574);
nand U1783 (N_1783,In_190,In_3465);
xor U1784 (N_1784,In_419,In_896);
xor U1785 (N_1785,In_2849,In_4679);
xnor U1786 (N_1786,In_3679,In_1701);
nand U1787 (N_1787,In_2218,In_420);
xnor U1788 (N_1788,In_1874,In_3150);
xnor U1789 (N_1789,In_4798,In_3134);
or U1790 (N_1790,In_2844,In_478);
or U1791 (N_1791,In_3733,In_2764);
and U1792 (N_1792,In_407,In_3715);
xor U1793 (N_1793,In_2008,In_2306);
or U1794 (N_1794,In_2622,In_4925);
nor U1795 (N_1795,In_4979,In_1228);
and U1796 (N_1796,In_2510,In_910);
or U1797 (N_1797,In_1098,In_34);
nand U1798 (N_1798,In_743,In_354);
or U1799 (N_1799,In_2425,In_1253);
xnor U1800 (N_1800,In_1857,In_3972);
xnor U1801 (N_1801,In_131,In_1928);
xnor U1802 (N_1802,In_3195,In_2022);
xor U1803 (N_1803,In_3346,In_611);
xnor U1804 (N_1804,In_4575,In_1275);
nand U1805 (N_1805,In_2598,In_4490);
nor U1806 (N_1806,In_1568,In_3754);
or U1807 (N_1807,In_283,In_4933);
nor U1808 (N_1808,In_2891,In_1603);
and U1809 (N_1809,In_385,In_1375);
and U1810 (N_1810,In_105,In_4599);
xor U1811 (N_1811,In_2495,In_2606);
xor U1812 (N_1812,In_1566,In_1718);
or U1813 (N_1813,In_1793,In_4018);
nand U1814 (N_1814,In_612,In_2061);
nand U1815 (N_1815,In_2054,In_3390);
xnor U1816 (N_1816,In_4402,In_1065);
nand U1817 (N_1817,In_1357,In_510);
nor U1818 (N_1818,In_4438,In_364);
or U1819 (N_1819,In_377,In_569);
xnor U1820 (N_1820,In_2769,In_868);
nor U1821 (N_1821,In_1420,In_3380);
or U1822 (N_1822,In_4188,In_3191);
and U1823 (N_1823,In_178,In_3122);
nand U1824 (N_1824,In_3617,In_2789);
xor U1825 (N_1825,In_3263,In_587);
nand U1826 (N_1826,In_2889,In_3994);
nand U1827 (N_1827,In_3516,In_2787);
nand U1828 (N_1828,In_2050,In_3498);
nor U1829 (N_1829,In_2554,In_2741);
nor U1830 (N_1830,In_4085,In_3396);
nor U1831 (N_1831,In_410,In_4037);
nand U1832 (N_1832,In_255,In_3215);
nand U1833 (N_1833,In_2453,In_3071);
nand U1834 (N_1834,In_1298,In_1088);
and U1835 (N_1835,In_2440,In_983);
and U1836 (N_1836,In_3182,In_23);
nand U1837 (N_1837,In_4143,In_4267);
or U1838 (N_1838,In_38,In_2593);
and U1839 (N_1839,In_1962,In_1425);
xor U1840 (N_1840,In_4742,In_96);
nand U1841 (N_1841,In_4335,In_1771);
or U1842 (N_1842,In_2184,In_2087);
and U1843 (N_1843,In_4523,In_1924);
or U1844 (N_1844,In_4110,In_4417);
nor U1845 (N_1845,In_4075,In_1669);
and U1846 (N_1846,In_715,In_2954);
xnor U1847 (N_1847,In_1067,In_1610);
or U1848 (N_1848,In_2338,In_655);
or U1849 (N_1849,In_789,In_2435);
and U1850 (N_1850,In_2371,In_2842);
xnor U1851 (N_1851,In_4755,In_3026);
and U1852 (N_1852,In_2446,In_3266);
or U1853 (N_1853,In_1274,In_926);
xnor U1854 (N_1854,In_324,In_2517);
nand U1855 (N_1855,In_2132,In_2582);
and U1856 (N_1856,In_2775,In_472);
xor U1857 (N_1857,In_513,In_4063);
nor U1858 (N_1858,In_1510,In_3845);
or U1859 (N_1859,In_4238,In_4986);
and U1860 (N_1860,In_2251,In_3397);
xor U1861 (N_1861,In_974,In_2097);
xnor U1862 (N_1862,In_1809,In_3356);
nor U1863 (N_1863,In_3412,In_1998);
nand U1864 (N_1864,In_3738,In_1984);
or U1865 (N_1865,In_134,In_2209);
and U1866 (N_1866,In_2314,In_621);
nor U1867 (N_1867,In_3834,In_3460);
xnor U1868 (N_1868,In_4613,In_3922);
and U1869 (N_1869,In_195,In_1745);
or U1870 (N_1870,In_3551,In_1770);
or U1871 (N_1871,In_2989,In_3489);
xor U1872 (N_1872,In_824,In_4650);
nand U1873 (N_1873,In_2272,In_1519);
nor U1874 (N_1874,In_2994,In_4506);
nor U1875 (N_1875,In_1641,In_3183);
nand U1876 (N_1876,In_3627,In_2655);
or U1877 (N_1877,In_631,In_3213);
and U1878 (N_1878,In_1179,In_2538);
nor U1879 (N_1879,In_4951,In_3935);
and U1880 (N_1880,In_4805,In_850);
or U1881 (N_1881,In_2383,In_1749);
or U1882 (N_1882,In_3086,In_4818);
or U1883 (N_1883,In_1583,In_1407);
or U1884 (N_1884,In_1128,In_4569);
xor U1885 (N_1885,In_4489,In_4182);
xor U1886 (N_1886,In_2945,In_3462);
or U1887 (N_1887,In_2171,In_336);
or U1888 (N_1888,In_2933,In_2985);
nand U1889 (N_1889,In_616,In_841);
xnor U1890 (N_1890,In_1041,In_2963);
nor U1891 (N_1891,In_779,In_2027);
nor U1892 (N_1892,In_4292,In_4125);
xnor U1893 (N_1893,In_3521,In_750);
or U1894 (N_1894,In_4170,In_1993);
and U1895 (N_1895,In_249,In_1367);
xor U1896 (N_1896,In_682,In_4950);
and U1897 (N_1897,In_1816,In_4703);
and U1898 (N_1898,In_4468,In_2417);
and U1899 (N_1899,In_2479,In_1272);
and U1900 (N_1900,In_1042,In_191);
nor U1901 (N_1901,In_3188,In_4262);
and U1902 (N_1902,In_3260,In_421);
and U1903 (N_1903,In_4406,In_275);
nor U1904 (N_1904,In_972,In_2161);
nor U1905 (N_1905,In_2407,In_4029);
or U1906 (N_1906,In_4407,In_1720);
xor U1907 (N_1907,In_3612,In_4151);
xnor U1908 (N_1908,In_4513,In_4960);
nand U1909 (N_1909,In_863,In_1071);
nand U1910 (N_1910,In_568,In_1961);
nand U1911 (N_1911,In_2939,In_3482);
nand U1912 (N_1912,In_937,In_1973);
and U1913 (N_1913,In_4253,In_3767);
and U1914 (N_1914,In_1607,In_3275);
xor U1915 (N_1915,In_1903,In_333);
xor U1916 (N_1916,In_4268,In_4604);
nor U1917 (N_1917,In_225,In_921);
xnor U1918 (N_1918,In_2601,In_2811);
nor U1919 (N_1919,In_3824,In_3361);
and U1920 (N_1920,In_526,In_1127);
nand U1921 (N_1921,In_2770,In_395);
xor U1922 (N_1922,In_2822,In_4782);
xnor U1923 (N_1923,In_1464,In_874);
nand U1924 (N_1924,In_1490,In_4265);
xor U1925 (N_1925,In_174,In_4369);
nor U1926 (N_1926,In_4600,In_1003);
nor U1927 (N_1927,In_2051,In_3582);
xnor U1928 (N_1928,In_3168,In_3175);
xnor U1929 (N_1929,In_825,In_4676);
and U1930 (N_1930,In_994,In_3135);
or U1931 (N_1931,In_827,In_3256);
nor U1932 (N_1932,In_2721,In_4579);
xnor U1933 (N_1933,In_4975,In_4919);
nand U1934 (N_1934,In_3967,In_1126);
xor U1935 (N_1935,In_4270,In_3029);
or U1936 (N_1936,In_1044,In_349);
or U1937 (N_1937,In_104,In_613);
xnor U1938 (N_1938,In_90,In_2573);
nand U1939 (N_1939,In_40,In_128);
nand U1940 (N_1940,In_1623,In_203);
xor U1941 (N_1941,In_3866,In_1908);
xnor U1942 (N_1942,In_3028,In_1159);
or U1943 (N_1943,In_3387,In_3235);
nand U1944 (N_1944,In_752,In_1679);
nor U1945 (N_1945,In_495,In_3876);
and U1946 (N_1946,In_2317,In_2211);
and U1947 (N_1947,In_4213,In_4969);
nor U1948 (N_1948,In_2264,In_1343);
nand U1949 (N_1949,In_2505,In_256);
and U1950 (N_1950,In_1413,In_2955);
xor U1951 (N_1951,In_3877,In_1555);
xor U1952 (N_1952,In_4866,In_94);
or U1953 (N_1953,In_3939,In_4300);
or U1954 (N_1954,In_2507,In_2747);
nand U1955 (N_1955,In_3563,In_238);
nand U1956 (N_1956,In_1220,In_3244);
xnor U1957 (N_1957,In_1674,In_1675);
and U1958 (N_1958,In_667,In_348);
nor U1959 (N_1959,In_2103,In_2113);
xnor U1960 (N_1960,In_953,In_857);
or U1961 (N_1961,In_927,In_437);
nand U1962 (N_1962,In_3995,In_3114);
xor U1963 (N_1963,In_3085,In_3663);
nor U1964 (N_1964,In_68,In_3693);
nand U1965 (N_1965,In_2750,In_4375);
nand U1966 (N_1966,In_4945,In_3823);
xnor U1967 (N_1967,In_4562,In_500);
xnor U1968 (N_1968,In_3314,In_4272);
and U1969 (N_1969,In_1616,In_2316);
nand U1970 (N_1970,In_2095,In_2299);
nand U1971 (N_1971,In_430,In_4059);
and U1972 (N_1972,In_1578,In_2402);
or U1973 (N_1973,In_991,In_2758);
and U1974 (N_1974,In_1887,In_3807);
xor U1975 (N_1975,In_1378,In_1299);
xor U1976 (N_1976,In_2729,In_3227);
or U1977 (N_1977,In_4084,In_56);
nand U1978 (N_1978,In_2839,In_2908);
nor U1979 (N_1979,In_4797,In_1292);
xnor U1980 (N_1980,In_543,In_4773);
and U1981 (N_1981,In_3303,In_4571);
nand U1982 (N_1982,In_2389,In_3098);
and U1983 (N_1983,In_2509,In_689);
nor U1984 (N_1984,In_4751,In_2270);
or U1985 (N_1985,In_4215,In_1033);
nand U1986 (N_1986,In_3723,In_2608);
xor U1987 (N_1987,In_837,In_3491);
nor U1988 (N_1988,In_1162,In_1094);
nand U1989 (N_1989,In_4435,In_3865);
or U1990 (N_1990,In_4401,In_3589);
xnor U1991 (N_1991,In_1747,In_2384);
nand U1992 (N_1992,In_4906,In_44);
or U1993 (N_1993,In_4391,In_4527);
or U1994 (N_1994,In_1577,In_4998);
nand U1995 (N_1995,In_3112,In_2301);
or U1996 (N_1996,In_990,In_2708);
and U1997 (N_1997,In_286,In_4220);
xor U1998 (N_1998,In_4221,In_3283);
and U1999 (N_1999,In_2937,In_986);
and U2000 (N_2000,In_1136,In_3409);
or U2001 (N_2001,In_54,In_3250);
xnor U2002 (N_2002,In_4184,In_2746);
or U2003 (N_2003,In_3628,In_2074);
nand U2004 (N_2004,In_1493,In_3445);
nor U2005 (N_2005,In_4826,In_2330);
xor U2006 (N_2006,In_3633,In_2136);
nor U2007 (N_2007,In_1948,In_3315);
or U2008 (N_2008,In_3307,In_2409);
or U2009 (N_2009,In_2427,In_1775);
nor U2010 (N_2010,In_4901,In_2942);
nand U2011 (N_2011,In_552,In_459);
nand U2012 (N_2012,In_4001,In_2055);
nand U2013 (N_2013,In_3092,In_3507);
and U2014 (N_2014,In_2294,In_1277);
nand U2015 (N_2015,In_1585,In_205);
xor U2016 (N_2016,In_280,In_3371);
nand U2017 (N_2017,In_3526,In_362);
nor U2018 (N_2018,In_3506,In_2170);
or U2019 (N_2019,In_1284,In_2735);
nand U2020 (N_2020,In_1602,In_1483);
nand U2021 (N_2021,In_4977,In_2586);
and U2022 (N_2022,In_1340,In_711);
xnor U2023 (N_2023,In_4454,In_869);
nand U2024 (N_2024,In_499,In_3154);
nand U2025 (N_2025,In_4142,In_4381);
nand U2026 (N_2026,In_204,In_1417);
xnor U2027 (N_2027,In_97,In_2292);
xnor U2028 (N_2028,In_3613,In_835);
nor U2029 (N_2029,In_703,In_431);
and U2030 (N_2030,In_1531,In_2334);
xnor U2031 (N_2031,In_3720,In_3982);
xnor U2032 (N_2032,In_2092,In_1494);
xor U2033 (N_2033,In_3317,In_399);
xor U2034 (N_2034,In_1671,In_383);
nor U2035 (N_2035,In_3212,In_3360);
nand U2036 (N_2036,In_4942,In_265);
xor U2037 (N_2037,In_3042,In_4161);
xor U2038 (N_2038,In_4337,In_4514);
or U2039 (N_2039,In_3568,In_3294);
and U2040 (N_2040,In_1946,In_1600);
nor U2041 (N_2041,In_2326,In_3889);
and U2042 (N_2042,In_856,In_4248);
nor U2043 (N_2043,In_1353,In_1322);
nand U2044 (N_2044,In_99,In_4211);
nand U2045 (N_2045,In_3736,In_948);
nor U2046 (N_2046,In_1639,In_4421);
xnor U2047 (N_2047,In_2590,In_3274);
nand U2048 (N_2048,In_4434,In_4816);
nand U2049 (N_2049,In_2356,In_1937);
or U2050 (N_2050,In_4615,In_785);
xnor U2051 (N_2051,In_620,In_925);
or U2052 (N_2052,In_4766,In_4970);
and U2053 (N_2053,In_1786,In_1215);
xnor U2054 (N_2054,In_3588,In_394);
or U2055 (N_2055,In_3862,In_2181);
and U2056 (N_2056,In_4980,In_3544);
or U2057 (N_2057,In_3221,In_610);
or U2058 (N_2058,In_1933,In_2640);
and U2059 (N_2059,In_1868,In_4011);
nor U2060 (N_2060,In_2244,In_897);
nand U2061 (N_2061,In_674,In_4205);
xor U2062 (N_2062,In_4667,In_337);
xor U2063 (N_2063,In_795,In_2464);
xnor U2064 (N_2064,In_1389,In_4285);
nor U2065 (N_2065,In_4102,In_3689);
and U2066 (N_2066,In_1364,In_2665);
xor U2067 (N_2067,In_355,In_4889);
and U2068 (N_2068,In_2823,In_3369);
nand U2069 (N_2069,In_1918,In_3430);
or U2070 (N_2070,In_251,In_4289);
nor U2071 (N_2071,In_929,In_3763);
and U2072 (N_2072,In_230,In_4035);
and U2073 (N_2073,In_4323,In_1188);
xnor U2074 (N_2074,In_3913,In_473);
nand U2075 (N_2075,In_2375,In_4000);
nor U2076 (N_2076,In_2696,In_2245);
xnor U2077 (N_2077,In_47,In_70);
and U2078 (N_2078,In_2778,In_1911);
nor U2079 (N_2079,In_389,In_2638);
xor U2080 (N_2080,In_4984,In_2274);
or U2081 (N_2081,In_2042,In_4034);
or U2082 (N_2082,In_4922,In_1150);
or U2083 (N_2083,In_4354,In_2212);
nand U2084 (N_2084,In_3717,In_2255);
xor U2085 (N_2085,In_3004,In_3005);
nor U2086 (N_2086,In_4512,In_1789);
or U2087 (N_2087,In_2754,In_3453);
nor U2088 (N_2088,In_318,In_2514);
nor U2089 (N_2089,In_634,In_1943);
nor U2090 (N_2090,In_2845,In_57);
or U2091 (N_2091,In_2714,In_4552);
xor U2092 (N_2092,In_1465,In_2652);
and U2093 (N_2093,In_3586,In_1118);
nand U2094 (N_2094,In_316,In_647);
nor U2095 (N_2095,In_4118,In_1370);
and U2096 (N_2096,In_3162,In_293);
nor U2097 (N_2097,In_4317,In_2563);
nand U2098 (N_2098,In_547,In_3864);
or U2099 (N_2099,In_1890,In_4509);
and U2100 (N_2100,In_1050,In_1352);
or U2101 (N_2101,In_3014,In_3403);
nand U2102 (N_2102,In_2287,In_3214);
nand U2103 (N_2103,In_27,In_2368);
xor U2104 (N_2104,In_2208,In_3936);
nor U2105 (N_2105,In_2612,In_4095);
or U2106 (N_2106,In_4993,In_2346);
nor U2107 (N_2107,In_1052,In_4131);
nand U2108 (N_2108,In_939,In_3268);
and U2109 (N_2109,In_3492,In_4568);
xnor U2110 (N_2110,In_2579,In_4393);
and U2111 (N_2111,In_4825,In_1892);
and U2112 (N_2112,In_2377,In_1176);
xnor U2113 (N_2113,In_4526,In_3739);
nor U2114 (N_2114,In_1582,In_4999);
and U2115 (N_2115,In_4521,In_2434);
nand U2116 (N_2116,In_2447,In_2654);
or U2117 (N_2117,In_3825,In_2122);
xor U2118 (N_2118,In_45,In_1522);
xor U2119 (N_2119,In_2808,In_2145);
or U2120 (N_2120,In_4716,In_102);
or U2121 (N_2121,In_2271,In_4444);
or U2122 (N_2122,In_2712,In_2072);
nor U2123 (N_2123,In_4418,In_695);
and U2124 (N_2124,In_2387,In_2656);
nor U2125 (N_2125,In_3458,In_2726);
xor U2126 (N_2126,In_4104,In_2082);
and U2127 (N_2127,In_231,In_847);
nand U2128 (N_2128,In_2561,In_4874);
xor U2129 (N_2129,In_1783,In_4281);
xor U2130 (N_2130,In_3104,In_4694);
or U2131 (N_2131,In_3772,In_3698);
or U2132 (N_2132,In_4321,In_2824);
nor U2133 (N_2133,In_3514,In_32);
or U2134 (N_2134,In_2470,In_1120);
nand U2135 (N_2135,In_3749,In_4706);
and U2136 (N_2136,In_330,In_2763);
nand U2137 (N_2137,In_4973,In_222);
and U2138 (N_2138,In_100,In_3142);
and U2139 (N_2139,In_1672,In_3017);
nand U2140 (N_2140,In_4750,In_411);
xnor U2141 (N_2141,In_4130,In_4839);
nor U2142 (N_2142,In_3432,In_221);
nor U2143 (N_2143,In_1576,In_1004);
xnor U2144 (N_2144,In_144,In_577);
xnor U2145 (N_2145,In_4291,In_3912);
or U2146 (N_2146,In_3065,In_4486);
or U2147 (N_2147,In_1787,In_2268);
and U2148 (N_2148,In_2877,In_4397);
or U2149 (N_2149,In_945,In_3625);
nand U2150 (N_2150,In_4264,In_4795);
or U2151 (N_2151,In_4729,In_4641);
nor U2152 (N_2152,In_1178,In_4698);
nor U2153 (N_2153,In_3043,In_3197);
xor U2154 (N_2154,In_4530,In_1416);
nor U2155 (N_2155,In_3861,In_691);
or U2156 (N_2156,In_4510,In_1119);
or U2157 (N_2157,In_4008,In_3621);
nand U2158 (N_2158,In_1680,In_271);
and U2159 (N_2159,In_453,In_1365);
and U2160 (N_2160,In_1537,In_3487);
and U2161 (N_2161,In_1154,In_2354);
nand U2162 (N_2162,In_1488,In_2728);
xor U2163 (N_2163,In_3764,In_1334);
nor U2164 (N_2164,In_1434,In_3222);
and U2165 (N_2165,In_1069,In_3872);
or U2166 (N_2166,In_3466,In_292);
nor U2167 (N_2167,In_2038,In_2491);
nor U2168 (N_2168,In_187,In_417);
nor U2169 (N_2169,In_372,In_3822);
xor U2170 (N_2170,In_154,In_1848);
nand U2171 (N_2171,In_1433,In_4320);
nor U2172 (N_2172,In_4824,In_2454);
or U2173 (N_2173,In_2291,In_2674);
or U2174 (N_2174,In_414,In_382);
or U2175 (N_2175,In_2378,In_4361);
and U2176 (N_2176,In_1549,In_3241);
nand U2177 (N_2177,In_931,In_2815);
and U2178 (N_2178,In_3856,In_3511);
and U2179 (N_2179,In_342,In_4733);
xnor U2180 (N_2180,In_4297,In_366);
or U2181 (N_2181,In_15,In_744);
nor U2182 (N_2182,In_1710,In_3954);
xnor U2183 (N_2183,In_3090,In_888);
and U2184 (N_2184,In_3273,In_1769);
nand U2185 (N_2185,In_2949,In_1655);
nor U2186 (N_2186,In_1160,In_4006);
xor U2187 (N_2187,In_3509,In_2745);
or U2188 (N_2188,In_3850,In_1309);
and U2189 (N_2189,In_849,In_2542);
nor U2190 (N_2190,In_1896,In_1554);
xnor U2191 (N_2191,In_2904,In_797);
xor U2192 (N_2192,In_4860,In_2946);
xor U2193 (N_2193,In_924,In_1076);
or U2194 (N_2194,In_74,In_842);
and U2195 (N_2195,In_979,In_2664);
nor U2196 (N_2196,In_4723,In_390);
and U2197 (N_2197,In_4913,In_3144);
nor U2198 (N_2198,In_4885,In_889);
nor U2199 (N_2199,In_2068,In_4581);
and U2200 (N_2200,In_259,In_4687);
or U2201 (N_2201,In_4411,In_3027);
nand U2202 (N_2202,In_2466,In_4668);
nand U2203 (N_2203,In_938,In_2352);
nor U2204 (N_2204,In_3901,In_2544);
nor U2205 (N_2205,In_3272,In_3267);
and U2206 (N_2206,In_373,In_3126);
nor U2207 (N_2207,In_4053,In_3811);
nand U2208 (N_2208,In_1103,In_1010);
and U2209 (N_2209,In_593,In_4405);
and U2210 (N_2210,In_456,In_3481);
or U2211 (N_2211,In_2100,In_4501);
nand U2212 (N_2212,In_1014,In_3113);
and U2213 (N_2213,In_1673,In_1886);
nand U2214 (N_2214,In_200,In_380);
nand U2215 (N_2215,In_4832,In_1297);
nand U2216 (N_2216,In_3392,In_515);
or U2217 (N_2217,In_108,In_2982);
nand U2218 (N_2218,In_4057,In_2214);
nor U2219 (N_2219,In_1536,In_1862);
nand U2220 (N_2220,In_1916,In_3473);
nor U2221 (N_2221,In_4564,In_3691);
nor U2222 (N_2222,In_3038,In_2350);
nand U2223 (N_2223,In_1589,In_3695);
xnor U2224 (N_2224,In_4250,In_1904);
nand U2225 (N_2225,In_3858,In_3075);
xnor U2226 (N_2226,In_761,In_3672);
nand U2227 (N_2227,In_644,In_3860);
or U2228 (N_2228,In_3362,In_799);
xnor U2229 (N_2229,In_3413,In_3194);
or U2230 (N_2230,In_1562,In_1436);
nand U2231 (N_2231,In_341,In_160);
nand U2232 (N_2232,In_2833,In_861);
and U2233 (N_2233,In_3270,In_1155);
xor U2234 (N_2234,In_2681,In_2030);
and U2235 (N_2235,In_2730,In_4903);
or U2236 (N_2236,In_2738,In_1080);
nor U2237 (N_2237,In_4322,In_505);
nand U2238 (N_2238,In_2901,In_86);
nand U2239 (N_2239,In_2814,In_3963);
nand U2240 (N_2240,In_3200,In_3924);
or U2241 (N_2241,In_2515,In_1056);
nand U2242 (N_2242,In_4450,In_3229);
nand U2243 (N_2243,In_3335,In_3968);
or U2244 (N_2244,In_1683,In_1931);
or U2245 (N_2245,In_116,In_1648);
nand U2246 (N_2246,In_1374,In_753);
nand U2247 (N_2247,In_1237,In_2265);
and U2248 (N_2248,In_4410,In_1929);
or U2249 (N_2249,In_2134,In_3350);
and U2250 (N_2250,In_4166,In_2293);
nand U2251 (N_2251,In_1443,In_764);
nor U2252 (N_2252,In_2677,In_1526);
nand U2253 (N_2253,In_375,In_177);
nor U2254 (N_2254,In_2972,In_3904);
xnor U2255 (N_2255,In_1553,In_1656);
nor U2256 (N_2256,In_1037,In_1325);
and U2257 (N_2257,In_1815,In_4329);
nor U2258 (N_2258,In_2355,In_624);
or U2259 (N_2259,In_1797,In_3943);
nor U2260 (N_2260,In_4462,In_80);
xor U2261 (N_2261,In_1755,In_3157);
xnor U2262 (N_2262,In_4882,In_4197);
or U2263 (N_2263,In_4536,In_2010);
or U2264 (N_2264,In_3536,In_4731);
or U2265 (N_2265,In_2860,In_2176);
nor U2266 (N_2266,In_3230,In_4244);
and U2267 (N_2267,In_3363,In_2874);
or U2268 (N_2268,In_3082,In_3933);
nand U2269 (N_2269,In_518,In_2625);
nor U2270 (N_2270,In_3955,In_1632);
nand U2271 (N_2271,In_1677,In_2200);
nor U2272 (N_2272,In_1405,In_1551);
or U2273 (N_2273,In_3532,In_3035);
nor U2274 (N_2274,In_1729,In_4767);
xor U2275 (N_2275,In_1060,In_1618);
or U2276 (N_2276,In_2288,In_3237);
nand U2277 (N_2277,In_1719,In_632);
nand U2278 (N_2278,In_4863,In_4743);
and U2279 (N_2279,In_1513,In_1541);
xnor U2280 (N_2280,In_1271,In_2547);
nand U2281 (N_2281,In_3529,In_359);
nand U2282 (N_2282,In_2431,In_3365);
and U2283 (N_2283,In_3619,In_4146);
nor U2284 (N_2284,In_3016,In_1011);
or U2285 (N_2285,In_424,In_3087);
and U2286 (N_2286,In_4654,In_2468);
xnor U2287 (N_2287,In_1063,In_746);
or U2288 (N_2288,In_1844,In_3459);
or U2289 (N_2289,In_3201,In_2543);
xor U2290 (N_2290,In_2875,In_2085);
nand U2291 (N_2291,In_640,In_4204);
or U2292 (N_2292,In_1091,In_4725);
and U2293 (N_2293,In_180,In_712);
nand U2294 (N_2294,In_4609,In_309);
nand U2295 (N_2295,In_1345,In_2413);
or U2296 (N_2296,In_3854,In_4657);
or U2297 (N_2297,In_4302,In_2820);
or U2298 (N_2298,In_1545,In_1803);
xor U2299 (N_2299,In_2462,In_1227);
nor U2300 (N_2300,In_1331,In_3123);
and U2301 (N_2301,In_550,In_971);
nand U2302 (N_2302,In_2902,In_3791);
nor U2303 (N_2303,In_1878,In_1009);
and U2304 (N_2304,In_2331,In_1339);
or U2305 (N_2305,In_1624,In_1926);
nand U2306 (N_2306,In_2062,In_4886);
nor U2307 (N_2307,In_4060,In_224);
and U2308 (N_2308,In_3658,In_159);
and U2309 (N_2309,In_4463,In_1181);
and U2310 (N_2310,In_2121,In_4064);
nand U2311 (N_2311,In_1401,In_2096);
nand U2312 (N_2312,In_4347,In_2861);
nor U2313 (N_2313,In_2619,In_1055);
and U2314 (N_2314,In_4732,In_3152);
nor U2315 (N_2315,In_1015,In_1283);
nand U2316 (N_2316,In_4541,In_4910);
xor U2317 (N_2317,In_2091,In_4148);
and U2318 (N_2318,In_2965,In_1244);
or U2319 (N_2319,In_3810,In_1716);
nor U2320 (N_2320,In_1900,In_338);
nand U2321 (N_2321,In_1104,In_2399);
xnor U2322 (N_2322,In_1457,In_2878);
or U2323 (N_2323,In_4622,In_4684);
nor U2324 (N_2324,In_1939,In_4626);
and U2325 (N_2325,In_3567,In_1027);
and U2326 (N_2326,In_3596,In_386);
nor U2327 (N_2327,In_3517,In_2799);
or U2328 (N_2328,In_3226,In_1295);
xnor U2329 (N_2329,In_305,In_2838);
or U2330 (N_2330,In_4054,In_374);
nor U2331 (N_2331,In_3778,In_4938);
xor U2332 (N_2332,In_3730,In_872);
xnor U2333 (N_2333,In_4133,In_1229);
or U2334 (N_2334,In_4842,In_911);
and U2335 (N_2335,In_4033,In_4469);
xor U2336 (N_2336,In_3792,In_321);
or U2337 (N_2337,In_4296,In_1115);
and U2338 (N_2338,In_1831,In_1736);
or U2339 (N_2339,In_1969,In_2243);
nor U2340 (N_2340,In_448,In_3560);
xnor U2341 (N_2341,In_4440,In_4083);
and U2342 (N_2342,In_3893,In_4152);
or U2343 (N_2343,In_458,In_4540);
and U2344 (N_2344,In_2289,In_1396);
xnor U2345 (N_2345,In_4608,In_3348);
and U2346 (N_2346,In_3690,In_2834);
xnor U2347 (N_2347,In_2846,In_4384);
xnor U2348 (N_2348,In_2026,In_172);
nor U2349 (N_2349,In_3976,In_680);
and U2350 (N_2350,In_2585,In_2717);
xnor U2351 (N_2351,In_3442,In_2343);
and U2352 (N_2352,In_1902,In_2048);
xor U2353 (N_2353,In_965,In_4580);
or U2354 (N_2354,In_2069,In_3905);
xnor U2355 (N_2355,In_4639,In_3366);
or U2356 (N_2356,In_1927,In_2931);
nand U2357 (N_2357,In_3808,In_4326);
nand U2358 (N_2358,In_2913,In_2118);
or U2359 (N_2359,In_2175,In_3405);
nor U2360 (N_2360,In_1336,In_3217);
nor U2361 (N_2361,In_217,In_1847);
xor U2362 (N_2362,In_4500,In_441);
xnor U2363 (N_2363,In_3678,In_1987);
xor U2364 (N_2364,In_783,In_819);
nand U2365 (N_2365,In_2796,In_1381);
nand U2366 (N_2366,In_2736,In_1717);
nand U2367 (N_2367,In_1662,In_1263);
nor U2368 (N_2368,In_1843,In_2928);
nor U2369 (N_2369,In_451,In_2472);
or U2370 (N_2370,In_1839,In_4830);
xnor U2371 (N_2371,In_2344,In_1447);
nor U2372 (N_2372,In_3415,In_1912);
nand U2373 (N_2373,In_2016,In_1090);
nand U2374 (N_2374,In_865,In_2308);
xor U2375 (N_2375,In_588,In_4662);
nand U2376 (N_2376,In_4939,In_1463);
xor U2377 (N_2377,In_1419,In_4614);
or U2378 (N_2378,In_3863,In_3302);
nand U2379 (N_2379,In_3040,In_1242);
nor U2380 (N_2380,In_4660,In_4144);
nor U2381 (N_2381,In_3264,In_3727);
and U2382 (N_2382,In_219,In_1535);
or U2383 (N_2383,In_4032,In_4117);
nor U2384 (N_2384,In_881,In_4774);
xnor U2385 (N_2385,In_3422,In_756);
nor U2386 (N_2386,In_4811,In_3512);
and U2387 (N_2387,In_2194,In_1497);
xor U2388 (N_2388,In_1697,In_1949);
or U2389 (N_2389,In_3990,In_3022);
and U2390 (N_2390,In_506,In_638);
or U2391 (N_2391,In_2552,In_3793);
xor U2392 (N_2392,In_1523,In_1262);
or U2393 (N_2393,In_1765,In_1347);
nand U2394 (N_2394,In_3074,In_2502);
nand U2395 (N_2395,In_4149,In_3687);
xor U2396 (N_2396,In_4464,In_1773);
or U2397 (N_2397,In_786,In_1058);
and U2398 (N_2398,In_1072,In_19);
or U2399 (N_2399,In_2639,In_4327);
nand U2400 (N_2400,In_755,In_4164);
and U2401 (N_2401,In_648,In_4212);
and U2402 (N_2402,In_43,In_301);
nand U2403 (N_2403,In_2185,In_4167);
nor U2404 (N_2404,In_3402,In_2647);
nor U2405 (N_2405,In_3895,In_767);
nor U2406 (N_2406,In_2906,In_3379);
nor U2407 (N_2407,In_2361,In_4137);
or U2408 (N_2408,In_2803,In_2630);
nand U2409 (N_2409,In_2921,In_893);
nand U2410 (N_2410,In_2847,In_3742);
and U2411 (N_2411,In_2448,In_2261);
or U2412 (N_2412,In_1635,In_109);
xnor U2413 (N_2413,In_745,In_4480);
xor U2414 (N_2414,In_3398,In_3975);
and U2415 (N_2415,In_1854,In_3696);
and U2416 (N_2416,In_1266,In_2663);
nand U2417 (N_2417,In_3782,In_2037);
or U2418 (N_2418,In_4163,In_1556);
nand U2419 (N_2419,In_2503,In_4749);
nor U2420 (N_2420,In_2676,In_31);
and U2421 (N_2421,In_3785,In_2201);
nor U2422 (N_2422,In_2693,In_736);
and U2423 (N_2423,In_1774,In_3452);
or U2424 (N_2424,In_1341,In_4382);
or U2425 (N_2425,In_4648,In_882);
xor U2426 (N_2426,In_3353,In_2406);
nand U2427 (N_2427,In_1859,In_1804);
nand U2428 (N_2428,In_4219,In_3721);
or U2429 (N_2429,In_254,In_3180);
or U2430 (N_2430,In_4389,In_4014);
and U2431 (N_2431,In_4106,In_2179);
xnor U2432 (N_2432,In_1565,In_2993);
xor U2433 (N_2433,In_2498,In_1335);
or U2434 (N_2434,In_4304,In_1757);
or U2435 (N_2435,In_4853,In_1569);
or U2436 (N_2436,In_3750,In_396);
or U2437 (N_2437,In_107,In_1028);
and U2438 (N_2438,In_2621,In_1410);
nor U2439 (N_2439,In_4467,In_4254);
xor U2440 (N_2440,In_17,In_2124);
xnor U2441 (N_2441,In_1534,In_3801);
and U2442 (N_2442,In_207,In_3859);
nor U2443 (N_2443,In_2267,In_504);
nand U2444 (N_2444,In_2423,In_4081);
nand U2445 (N_2445,In_1406,In_3160);
nor U2446 (N_2446,In_2369,In_1474);
xor U2447 (N_2447,In_2359,In_2788);
and U2448 (N_2448,In_4912,In_434);
nor U2449 (N_2449,In_3389,In_4765);
and U2450 (N_2450,In_4365,In_151);
xnor U2451 (N_2451,In_1630,In_1856);
or U2452 (N_2452,In_1114,In_537);
xor U2453 (N_2453,In_1596,In_3439);
or U2454 (N_2454,In_2627,In_2305);
xor U2455 (N_2455,In_2866,In_2995);
and U2456 (N_2456,In_1152,In_987);
xor U2457 (N_2457,In_4383,In_579);
or U2458 (N_2458,In_4584,In_2641);
nand U2459 (N_2459,In_530,In_3671);
nor U2460 (N_2460,In_3436,In_4658);
nor U2461 (N_2461,In_1282,In_4079);
nand U2462 (N_2462,In_3880,In_1485);
nor U2463 (N_2463,In_1813,In_793);
nand U2464 (N_2464,In_4586,In_567);
nand U2465 (N_2465,In_4366,In_3282);
or U2466 (N_2466,In_2151,In_3242);
xnor U2467 (N_2467,In_2774,In_2419);
nor U2468 (N_2468,In_20,In_3304);
or U2469 (N_2469,In_1040,In_4132);
and U2470 (N_2470,In_467,In_4020);
and U2471 (N_2471,In_1592,In_3008);
or U2472 (N_2472,In_3844,In_4282);
and U2473 (N_2473,In_2073,In_3072);
nor U2474 (N_2474,In_1388,In_4483);
and U2475 (N_2475,In_4223,In_2232);
nand U2476 (N_2476,In_1552,In_1873);
xor U2477 (N_2477,In_838,In_2915);
nand U2478 (N_2478,In_2980,In_4994);
or U2479 (N_2479,In_1945,In_2034);
and U2480 (N_2480,In_3262,In_590);
nor U2481 (N_2481,In_4234,In_3930);
or U2482 (N_2482,In_192,In_742);
nand U2483 (N_2483,In_91,In_1359);
nand U2484 (N_2484,In_3795,In_1123);
or U2485 (N_2485,In_2321,In_4844);
nand U2486 (N_2486,In_2379,In_3604);
xor U2487 (N_2487,In_264,In_2481);
nor U2488 (N_2488,In_2894,In_4917);
nand U2489 (N_2489,In_2539,In_3472);
nor U2490 (N_2490,In_1303,In_3296);
nand U2491 (N_2491,In_3411,In_3783);
and U2492 (N_2492,In_3502,In_3243);
and U2493 (N_2493,In_1432,In_4772);
or U2494 (N_2494,In_2512,In_4052);
xnor U2495 (N_2495,In_4245,In_1836);
xor U2496 (N_2496,In_2986,In_4194);
or U2497 (N_2497,In_1026,In_2053);
xnor U2498 (N_2498,In_977,In_4328);
and U2499 (N_2499,In_2953,In_3166);
nor U2500 (N_2500,In_868,In_4445);
and U2501 (N_2501,In_3355,In_836);
and U2502 (N_2502,In_1119,In_2866);
or U2503 (N_2503,In_3047,In_3373);
xnor U2504 (N_2504,In_119,In_972);
and U2505 (N_2505,In_4558,In_1034);
and U2506 (N_2506,In_4339,In_1986);
nor U2507 (N_2507,In_1976,In_1069);
or U2508 (N_2508,In_430,In_2337);
and U2509 (N_2509,In_890,In_3296);
nand U2510 (N_2510,In_30,In_2159);
and U2511 (N_2511,In_558,In_3794);
and U2512 (N_2512,In_3744,In_3174);
nor U2513 (N_2513,In_1281,In_1342);
nand U2514 (N_2514,In_4555,In_3687);
and U2515 (N_2515,In_2633,In_4234);
nand U2516 (N_2516,In_4686,In_2673);
and U2517 (N_2517,In_189,In_1495);
or U2518 (N_2518,In_3014,In_232);
nand U2519 (N_2519,In_647,In_922);
nor U2520 (N_2520,In_1210,In_4553);
nor U2521 (N_2521,In_1224,In_181);
and U2522 (N_2522,In_3454,In_4155);
nor U2523 (N_2523,In_1943,In_537);
nand U2524 (N_2524,In_3655,In_264);
or U2525 (N_2525,In_3916,In_3238);
or U2526 (N_2526,In_2589,In_4063);
and U2527 (N_2527,In_2415,In_3338);
or U2528 (N_2528,In_503,In_476);
or U2529 (N_2529,In_1742,In_659);
and U2530 (N_2530,In_2614,In_2837);
or U2531 (N_2531,In_4,In_453);
nand U2532 (N_2532,In_4777,In_2201);
xor U2533 (N_2533,In_1245,In_1171);
and U2534 (N_2534,In_3504,In_282);
and U2535 (N_2535,In_1808,In_4380);
nor U2536 (N_2536,In_185,In_2232);
nor U2537 (N_2537,In_903,In_4588);
nor U2538 (N_2538,In_1671,In_4118);
nor U2539 (N_2539,In_4424,In_1596);
or U2540 (N_2540,In_453,In_1983);
nor U2541 (N_2541,In_3337,In_1949);
or U2542 (N_2542,In_29,In_4629);
nor U2543 (N_2543,In_4617,In_2657);
and U2544 (N_2544,In_1847,In_397);
nor U2545 (N_2545,In_2050,In_1816);
nor U2546 (N_2546,In_3598,In_2674);
xor U2547 (N_2547,In_4785,In_3836);
xor U2548 (N_2548,In_4159,In_4594);
xor U2549 (N_2549,In_1053,In_1532);
or U2550 (N_2550,In_2964,In_3502);
and U2551 (N_2551,In_1727,In_2472);
nand U2552 (N_2552,In_1480,In_4669);
or U2553 (N_2553,In_3546,In_4531);
nor U2554 (N_2554,In_3280,In_1114);
nand U2555 (N_2555,In_1387,In_3612);
or U2556 (N_2556,In_4744,In_3715);
nand U2557 (N_2557,In_4876,In_2412);
nor U2558 (N_2558,In_2086,In_4623);
nand U2559 (N_2559,In_3565,In_934);
and U2560 (N_2560,In_4743,In_3941);
and U2561 (N_2561,In_3947,In_4085);
or U2562 (N_2562,In_4057,In_3862);
and U2563 (N_2563,In_4420,In_3150);
nand U2564 (N_2564,In_2364,In_1989);
or U2565 (N_2565,In_4929,In_4014);
xnor U2566 (N_2566,In_1977,In_3361);
nor U2567 (N_2567,In_1588,In_207);
nor U2568 (N_2568,In_673,In_468);
or U2569 (N_2569,In_1924,In_2018);
and U2570 (N_2570,In_2556,In_1231);
nor U2571 (N_2571,In_3434,In_4994);
xnor U2572 (N_2572,In_350,In_1892);
nand U2573 (N_2573,In_2589,In_399);
and U2574 (N_2574,In_2309,In_2714);
nor U2575 (N_2575,In_3367,In_2901);
or U2576 (N_2576,In_1532,In_3550);
or U2577 (N_2577,In_1329,In_1583);
and U2578 (N_2578,In_4047,In_4854);
or U2579 (N_2579,In_398,In_2768);
nor U2580 (N_2580,In_3992,In_2683);
nand U2581 (N_2581,In_2535,In_1958);
nand U2582 (N_2582,In_2729,In_2004);
and U2583 (N_2583,In_1630,In_4802);
or U2584 (N_2584,In_2169,In_3535);
or U2585 (N_2585,In_3166,In_2369);
xnor U2586 (N_2586,In_126,In_3934);
or U2587 (N_2587,In_2510,In_416);
xnor U2588 (N_2588,In_4914,In_374);
and U2589 (N_2589,In_1157,In_371);
and U2590 (N_2590,In_4294,In_3004);
and U2591 (N_2591,In_3055,In_2395);
or U2592 (N_2592,In_4889,In_1854);
nor U2593 (N_2593,In_255,In_905);
or U2594 (N_2594,In_2928,In_4769);
nor U2595 (N_2595,In_2719,In_3153);
and U2596 (N_2596,In_587,In_4710);
nor U2597 (N_2597,In_2411,In_563);
and U2598 (N_2598,In_2043,In_682);
and U2599 (N_2599,In_65,In_438);
nor U2600 (N_2600,In_1079,In_1424);
xor U2601 (N_2601,In_767,In_4845);
nand U2602 (N_2602,In_2587,In_3909);
nand U2603 (N_2603,In_4037,In_2936);
nor U2604 (N_2604,In_1711,In_2605);
or U2605 (N_2605,In_1116,In_4086);
xnor U2606 (N_2606,In_2027,In_4151);
xor U2607 (N_2607,In_1208,In_2187);
nor U2608 (N_2608,In_2885,In_231);
nor U2609 (N_2609,In_1614,In_1084);
and U2610 (N_2610,In_2413,In_2328);
and U2611 (N_2611,In_2865,In_2090);
or U2612 (N_2612,In_781,In_814);
nand U2613 (N_2613,In_2841,In_3687);
nor U2614 (N_2614,In_2106,In_3872);
xor U2615 (N_2615,In_3020,In_2824);
nor U2616 (N_2616,In_421,In_3);
nand U2617 (N_2617,In_2494,In_2367);
and U2618 (N_2618,In_3747,In_1078);
nand U2619 (N_2619,In_3917,In_3651);
nand U2620 (N_2620,In_4045,In_720);
nand U2621 (N_2621,In_3643,In_3617);
xnor U2622 (N_2622,In_4625,In_1879);
or U2623 (N_2623,In_33,In_3681);
nand U2624 (N_2624,In_261,In_4538);
and U2625 (N_2625,In_3757,In_292);
nor U2626 (N_2626,In_4816,In_1123);
and U2627 (N_2627,In_4605,In_3241);
or U2628 (N_2628,In_4292,In_3672);
nor U2629 (N_2629,In_3103,In_1701);
xnor U2630 (N_2630,In_3210,In_4985);
nor U2631 (N_2631,In_285,In_2636);
xor U2632 (N_2632,In_338,In_3275);
and U2633 (N_2633,In_712,In_935);
nand U2634 (N_2634,In_1328,In_1589);
nand U2635 (N_2635,In_3576,In_4630);
nand U2636 (N_2636,In_4886,In_436);
nor U2637 (N_2637,In_1095,In_3075);
nand U2638 (N_2638,In_3265,In_2407);
nor U2639 (N_2639,In_3731,In_884);
and U2640 (N_2640,In_2033,In_4750);
nor U2641 (N_2641,In_269,In_4221);
xor U2642 (N_2642,In_2472,In_3753);
xor U2643 (N_2643,In_4731,In_2080);
nor U2644 (N_2644,In_910,In_3373);
and U2645 (N_2645,In_3316,In_2306);
and U2646 (N_2646,In_1315,In_3132);
or U2647 (N_2647,In_2756,In_4214);
xnor U2648 (N_2648,In_2881,In_796);
xor U2649 (N_2649,In_244,In_2273);
nand U2650 (N_2650,In_1795,In_42);
xnor U2651 (N_2651,In_3600,In_4254);
nand U2652 (N_2652,In_218,In_2950);
or U2653 (N_2653,In_220,In_562);
and U2654 (N_2654,In_2446,In_2208);
or U2655 (N_2655,In_1513,In_4735);
nor U2656 (N_2656,In_580,In_284);
nor U2657 (N_2657,In_3291,In_4028);
nor U2658 (N_2658,In_4461,In_3071);
xnor U2659 (N_2659,In_4318,In_926);
and U2660 (N_2660,In_2327,In_3114);
nor U2661 (N_2661,In_4374,In_1224);
and U2662 (N_2662,In_872,In_3737);
or U2663 (N_2663,In_4932,In_1194);
and U2664 (N_2664,In_2590,In_2628);
and U2665 (N_2665,In_4720,In_3245);
nand U2666 (N_2666,In_173,In_4962);
xor U2667 (N_2667,In_3861,In_4367);
nand U2668 (N_2668,In_2268,In_21);
xnor U2669 (N_2669,In_960,In_4368);
and U2670 (N_2670,In_2755,In_3545);
and U2671 (N_2671,In_4461,In_939);
and U2672 (N_2672,In_4827,In_4078);
xor U2673 (N_2673,In_608,In_854);
nor U2674 (N_2674,In_774,In_3483);
or U2675 (N_2675,In_599,In_4586);
and U2676 (N_2676,In_940,In_1651);
or U2677 (N_2677,In_3839,In_3000);
or U2678 (N_2678,In_2090,In_2820);
nand U2679 (N_2679,In_1629,In_4804);
nor U2680 (N_2680,In_4182,In_3704);
or U2681 (N_2681,In_2131,In_2764);
nand U2682 (N_2682,In_1438,In_1635);
and U2683 (N_2683,In_1577,In_4940);
nor U2684 (N_2684,In_2808,In_4285);
nor U2685 (N_2685,In_4795,In_3136);
nor U2686 (N_2686,In_4440,In_510);
and U2687 (N_2687,In_4861,In_3561);
or U2688 (N_2688,In_4451,In_2404);
and U2689 (N_2689,In_4207,In_3982);
and U2690 (N_2690,In_1373,In_3871);
xor U2691 (N_2691,In_4001,In_1499);
or U2692 (N_2692,In_2142,In_2455);
and U2693 (N_2693,In_2886,In_1695);
nor U2694 (N_2694,In_542,In_4232);
xor U2695 (N_2695,In_3595,In_590);
and U2696 (N_2696,In_518,In_3904);
xnor U2697 (N_2697,In_2277,In_1348);
xnor U2698 (N_2698,In_3209,In_2386);
or U2699 (N_2699,In_64,In_158);
nor U2700 (N_2700,In_2741,In_2412);
and U2701 (N_2701,In_1366,In_2616);
xor U2702 (N_2702,In_127,In_2582);
or U2703 (N_2703,In_4420,In_1736);
xnor U2704 (N_2704,In_3897,In_1775);
xnor U2705 (N_2705,In_1794,In_1925);
or U2706 (N_2706,In_4553,In_4107);
nor U2707 (N_2707,In_4827,In_2550);
xnor U2708 (N_2708,In_3186,In_379);
nand U2709 (N_2709,In_2741,In_3008);
and U2710 (N_2710,In_4709,In_4954);
nand U2711 (N_2711,In_1791,In_4582);
and U2712 (N_2712,In_4312,In_2696);
nand U2713 (N_2713,In_3358,In_4452);
and U2714 (N_2714,In_2201,In_2711);
nand U2715 (N_2715,In_4372,In_2593);
or U2716 (N_2716,In_3010,In_2541);
nand U2717 (N_2717,In_2786,In_711);
nand U2718 (N_2718,In_148,In_2748);
nand U2719 (N_2719,In_1779,In_3113);
nor U2720 (N_2720,In_1228,In_23);
nor U2721 (N_2721,In_301,In_4568);
xor U2722 (N_2722,In_278,In_2621);
xnor U2723 (N_2723,In_4737,In_3336);
nand U2724 (N_2724,In_4492,In_149);
nor U2725 (N_2725,In_4923,In_2152);
and U2726 (N_2726,In_1503,In_4114);
nand U2727 (N_2727,In_2320,In_182);
or U2728 (N_2728,In_3984,In_3467);
xor U2729 (N_2729,In_4241,In_746);
xor U2730 (N_2730,In_1654,In_4717);
and U2731 (N_2731,In_3167,In_1316);
and U2732 (N_2732,In_4979,In_33);
or U2733 (N_2733,In_1914,In_2503);
xor U2734 (N_2734,In_983,In_2102);
nand U2735 (N_2735,In_1339,In_368);
xnor U2736 (N_2736,In_1246,In_3110);
xor U2737 (N_2737,In_3878,In_1435);
and U2738 (N_2738,In_2757,In_3828);
xnor U2739 (N_2739,In_964,In_4531);
nor U2740 (N_2740,In_2452,In_2459);
or U2741 (N_2741,In_4893,In_852);
nor U2742 (N_2742,In_634,In_2330);
and U2743 (N_2743,In_2057,In_2687);
xor U2744 (N_2744,In_1911,In_1861);
nor U2745 (N_2745,In_4382,In_452);
and U2746 (N_2746,In_2787,In_1480);
nand U2747 (N_2747,In_2250,In_1250);
or U2748 (N_2748,In_1669,In_4179);
nor U2749 (N_2749,In_1166,In_2478);
nand U2750 (N_2750,In_179,In_4745);
nor U2751 (N_2751,In_899,In_2237);
or U2752 (N_2752,In_4632,In_3669);
or U2753 (N_2753,In_4227,In_3463);
and U2754 (N_2754,In_3472,In_2584);
nor U2755 (N_2755,In_4442,In_3279);
and U2756 (N_2756,In_4217,In_568);
nand U2757 (N_2757,In_287,In_3534);
nand U2758 (N_2758,In_3552,In_2175);
nand U2759 (N_2759,In_4141,In_2765);
and U2760 (N_2760,In_1225,In_1215);
xnor U2761 (N_2761,In_2890,In_4548);
nor U2762 (N_2762,In_3550,In_2445);
and U2763 (N_2763,In_161,In_2303);
nor U2764 (N_2764,In_3275,In_3772);
or U2765 (N_2765,In_1524,In_4119);
and U2766 (N_2766,In_476,In_2362);
xor U2767 (N_2767,In_1818,In_4592);
and U2768 (N_2768,In_3535,In_3281);
nand U2769 (N_2769,In_549,In_3392);
xnor U2770 (N_2770,In_3383,In_3052);
or U2771 (N_2771,In_3710,In_1103);
xor U2772 (N_2772,In_1356,In_3553);
xor U2773 (N_2773,In_1255,In_1822);
and U2774 (N_2774,In_2739,In_3403);
nand U2775 (N_2775,In_3631,In_1698);
nand U2776 (N_2776,In_367,In_2436);
nand U2777 (N_2777,In_4249,In_1340);
nor U2778 (N_2778,In_3334,In_4506);
xor U2779 (N_2779,In_4206,In_1426);
and U2780 (N_2780,In_945,In_4498);
nand U2781 (N_2781,In_3299,In_1203);
nand U2782 (N_2782,In_4404,In_4710);
or U2783 (N_2783,In_147,In_3561);
xor U2784 (N_2784,In_4030,In_4454);
and U2785 (N_2785,In_62,In_1484);
and U2786 (N_2786,In_2800,In_1950);
nor U2787 (N_2787,In_2644,In_2293);
nand U2788 (N_2788,In_4283,In_3220);
and U2789 (N_2789,In_428,In_1325);
xnor U2790 (N_2790,In_3036,In_1681);
nor U2791 (N_2791,In_4563,In_1557);
nand U2792 (N_2792,In_4541,In_4438);
nor U2793 (N_2793,In_1633,In_3040);
and U2794 (N_2794,In_4652,In_921);
and U2795 (N_2795,In_478,In_921);
nand U2796 (N_2796,In_2219,In_2370);
and U2797 (N_2797,In_842,In_2772);
and U2798 (N_2798,In_309,In_3896);
xnor U2799 (N_2799,In_3971,In_2945);
nor U2800 (N_2800,In_1083,In_3189);
nand U2801 (N_2801,In_2607,In_1761);
and U2802 (N_2802,In_2023,In_939);
nand U2803 (N_2803,In_1819,In_1522);
nor U2804 (N_2804,In_3735,In_918);
and U2805 (N_2805,In_869,In_3032);
nand U2806 (N_2806,In_4866,In_2009);
xor U2807 (N_2807,In_1598,In_3425);
or U2808 (N_2808,In_2236,In_1630);
xnor U2809 (N_2809,In_2906,In_1878);
nor U2810 (N_2810,In_639,In_1654);
or U2811 (N_2811,In_4449,In_2497);
nor U2812 (N_2812,In_3176,In_3005);
nor U2813 (N_2813,In_3723,In_4874);
or U2814 (N_2814,In_1115,In_3653);
or U2815 (N_2815,In_1399,In_3242);
and U2816 (N_2816,In_1427,In_3935);
and U2817 (N_2817,In_1260,In_2251);
and U2818 (N_2818,In_1597,In_1861);
xnor U2819 (N_2819,In_2514,In_1770);
or U2820 (N_2820,In_3033,In_833);
or U2821 (N_2821,In_1875,In_654);
or U2822 (N_2822,In_1079,In_116);
nand U2823 (N_2823,In_503,In_4066);
nand U2824 (N_2824,In_233,In_2879);
or U2825 (N_2825,In_1408,In_95);
or U2826 (N_2826,In_1055,In_2879);
xnor U2827 (N_2827,In_2638,In_3152);
nand U2828 (N_2828,In_669,In_4098);
and U2829 (N_2829,In_1481,In_3820);
and U2830 (N_2830,In_342,In_2099);
and U2831 (N_2831,In_3960,In_452);
and U2832 (N_2832,In_2386,In_1766);
xor U2833 (N_2833,In_1385,In_325);
or U2834 (N_2834,In_3901,In_4119);
and U2835 (N_2835,In_2931,In_3014);
nand U2836 (N_2836,In_3316,In_2537);
xor U2837 (N_2837,In_4515,In_679);
xnor U2838 (N_2838,In_1818,In_4038);
or U2839 (N_2839,In_3856,In_2433);
xnor U2840 (N_2840,In_3523,In_1350);
nand U2841 (N_2841,In_3940,In_914);
or U2842 (N_2842,In_2232,In_3519);
and U2843 (N_2843,In_4615,In_3966);
or U2844 (N_2844,In_4675,In_1488);
and U2845 (N_2845,In_2501,In_2718);
xnor U2846 (N_2846,In_4546,In_2713);
xnor U2847 (N_2847,In_935,In_460);
and U2848 (N_2848,In_3400,In_4015);
nor U2849 (N_2849,In_884,In_1149);
nand U2850 (N_2850,In_523,In_361);
nor U2851 (N_2851,In_3265,In_243);
or U2852 (N_2852,In_944,In_977);
or U2853 (N_2853,In_263,In_4462);
or U2854 (N_2854,In_3052,In_4835);
and U2855 (N_2855,In_3773,In_2816);
or U2856 (N_2856,In_387,In_1155);
nor U2857 (N_2857,In_725,In_677);
nand U2858 (N_2858,In_4710,In_1083);
xnor U2859 (N_2859,In_687,In_924);
xor U2860 (N_2860,In_150,In_3115);
nor U2861 (N_2861,In_4113,In_3745);
or U2862 (N_2862,In_4264,In_3767);
nand U2863 (N_2863,In_4765,In_4523);
and U2864 (N_2864,In_4938,In_1458);
xor U2865 (N_2865,In_3109,In_2520);
and U2866 (N_2866,In_1054,In_2670);
nor U2867 (N_2867,In_2477,In_166);
and U2868 (N_2868,In_1788,In_4168);
and U2869 (N_2869,In_3664,In_721);
xnor U2870 (N_2870,In_2267,In_2369);
nor U2871 (N_2871,In_4223,In_4324);
and U2872 (N_2872,In_3745,In_2152);
nand U2873 (N_2873,In_478,In_3620);
xnor U2874 (N_2874,In_1833,In_3413);
and U2875 (N_2875,In_3557,In_3188);
or U2876 (N_2876,In_4336,In_2345);
nor U2877 (N_2877,In_996,In_4369);
nand U2878 (N_2878,In_1064,In_2626);
nand U2879 (N_2879,In_1387,In_3110);
nand U2880 (N_2880,In_1380,In_335);
and U2881 (N_2881,In_1158,In_2305);
nand U2882 (N_2882,In_2554,In_184);
xor U2883 (N_2883,In_698,In_854);
or U2884 (N_2884,In_1789,In_2348);
xor U2885 (N_2885,In_4182,In_1680);
or U2886 (N_2886,In_752,In_1989);
nor U2887 (N_2887,In_279,In_1603);
or U2888 (N_2888,In_3332,In_4994);
nor U2889 (N_2889,In_791,In_3866);
or U2890 (N_2890,In_4587,In_4225);
and U2891 (N_2891,In_1687,In_4045);
xor U2892 (N_2892,In_2830,In_2293);
nand U2893 (N_2893,In_3656,In_4555);
nand U2894 (N_2894,In_3380,In_3050);
or U2895 (N_2895,In_334,In_648);
nor U2896 (N_2896,In_1364,In_4243);
xnor U2897 (N_2897,In_4739,In_1478);
nor U2898 (N_2898,In_4852,In_1558);
or U2899 (N_2899,In_3924,In_2451);
or U2900 (N_2900,In_4387,In_2516);
or U2901 (N_2901,In_2713,In_3908);
xor U2902 (N_2902,In_364,In_1671);
nor U2903 (N_2903,In_1007,In_4426);
xnor U2904 (N_2904,In_3835,In_2582);
nand U2905 (N_2905,In_727,In_3766);
xor U2906 (N_2906,In_701,In_3009);
nor U2907 (N_2907,In_4397,In_3272);
or U2908 (N_2908,In_133,In_3451);
xor U2909 (N_2909,In_317,In_2106);
xnor U2910 (N_2910,In_2388,In_3153);
xor U2911 (N_2911,In_105,In_230);
nand U2912 (N_2912,In_4386,In_1526);
xor U2913 (N_2913,In_610,In_4808);
and U2914 (N_2914,In_393,In_1595);
nand U2915 (N_2915,In_2136,In_489);
nand U2916 (N_2916,In_4721,In_1229);
nor U2917 (N_2917,In_1199,In_2108);
or U2918 (N_2918,In_4961,In_4234);
nor U2919 (N_2919,In_2617,In_178);
or U2920 (N_2920,In_271,In_2582);
xor U2921 (N_2921,In_2915,In_3616);
xor U2922 (N_2922,In_3437,In_35);
and U2923 (N_2923,In_14,In_3148);
xnor U2924 (N_2924,In_598,In_453);
or U2925 (N_2925,In_4137,In_3625);
nor U2926 (N_2926,In_3443,In_2788);
nor U2927 (N_2927,In_2187,In_3570);
or U2928 (N_2928,In_3103,In_2891);
or U2929 (N_2929,In_2349,In_3094);
or U2930 (N_2930,In_2492,In_3524);
or U2931 (N_2931,In_2482,In_2142);
and U2932 (N_2932,In_1779,In_3165);
or U2933 (N_2933,In_2472,In_1752);
nand U2934 (N_2934,In_1105,In_3354);
nor U2935 (N_2935,In_3446,In_4305);
xnor U2936 (N_2936,In_795,In_2630);
and U2937 (N_2937,In_944,In_2311);
nand U2938 (N_2938,In_2346,In_4177);
xnor U2939 (N_2939,In_3878,In_439);
or U2940 (N_2940,In_4004,In_3260);
xnor U2941 (N_2941,In_2606,In_4333);
and U2942 (N_2942,In_637,In_1396);
or U2943 (N_2943,In_734,In_3794);
nand U2944 (N_2944,In_658,In_3587);
xor U2945 (N_2945,In_179,In_3120);
nand U2946 (N_2946,In_3217,In_3845);
nor U2947 (N_2947,In_2606,In_2281);
and U2948 (N_2948,In_1150,In_3421);
xnor U2949 (N_2949,In_4803,In_3316);
xor U2950 (N_2950,In_4474,In_1009);
xor U2951 (N_2951,In_2279,In_2129);
and U2952 (N_2952,In_998,In_4160);
or U2953 (N_2953,In_3595,In_4927);
or U2954 (N_2954,In_1214,In_4947);
or U2955 (N_2955,In_2805,In_4450);
or U2956 (N_2956,In_4967,In_2331);
xnor U2957 (N_2957,In_2722,In_694);
or U2958 (N_2958,In_2031,In_3980);
or U2959 (N_2959,In_1812,In_336);
nand U2960 (N_2960,In_3308,In_4797);
or U2961 (N_2961,In_3587,In_211);
xnor U2962 (N_2962,In_2002,In_3346);
and U2963 (N_2963,In_2408,In_4071);
and U2964 (N_2964,In_3767,In_4080);
or U2965 (N_2965,In_437,In_4562);
nor U2966 (N_2966,In_1206,In_2561);
nor U2967 (N_2967,In_2784,In_4226);
nand U2968 (N_2968,In_481,In_1021);
nand U2969 (N_2969,In_2168,In_2802);
nor U2970 (N_2970,In_1083,In_3046);
xnor U2971 (N_2971,In_788,In_257);
and U2972 (N_2972,In_4086,In_4714);
nand U2973 (N_2973,In_3488,In_3412);
or U2974 (N_2974,In_254,In_3672);
nand U2975 (N_2975,In_4227,In_4778);
xor U2976 (N_2976,In_3809,In_4474);
and U2977 (N_2977,In_656,In_1997);
nand U2978 (N_2978,In_2076,In_272);
or U2979 (N_2979,In_2903,In_1541);
nand U2980 (N_2980,In_3441,In_4581);
and U2981 (N_2981,In_1268,In_528);
xnor U2982 (N_2982,In_4021,In_250);
nand U2983 (N_2983,In_289,In_2202);
xnor U2984 (N_2984,In_2032,In_4295);
xor U2985 (N_2985,In_204,In_2947);
and U2986 (N_2986,In_2900,In_1668);
or U2987 (N_2987,In_2585,In_4703);
nand U2988 (N_2988,In_4981,In_2585);
nor U2989 (N_2989,In_4638,In_2569);
and U2990 (N_2990,In_4606,In_1217);
nand U2991 (N_2991,In_4275,In_4641);
nor U2992 (N_2992,In_3564,In_74);
nor U2993 (N_2993,In_11,In_1774);
or U2994 (N_2994,In_2927,In_4388);
nor U2995 (N_2995,In_1475,In_2081);
nor U2996 (N_2996,In_287,In_1099);
xor U2997 (N_2997,In_567,In_965);
xor U2998 (N_2998,In_3974,In_3613);
nand U2999 (N_2999,In_2858,In_3914);
nand U3000 (N_3000,In_2419,In_804);
nor U3001 (N_3001,In_3183,In_935);
nand U3002 (N_3002,In_833,In_3011);
nor U3003 (N_3003,In_390,In_4959);
or U3004 (N_3004,In_4090,In_519);
and U3005 (N_3005,In_3262,In_3304);
and U3006 (N_3006,In_3686,In_3423);
nor U3007 (N_3007,In_4994,In_4051);
nor U3008 (N_3008,In_1737,In_2934);
and U3009 (N_3009,In_4900,In_3883);
or U3010 (N_3010,In_1714,In_886);
or U3011 (N_3011,In_2918,In_1705);
or U3012 (N_3012,In_4967,In_57);
xor U3013 (N_3013,In_868,In_3951);
xnor U3014 (N_3014,In_1207,In_1390);
nor U3015 (N_3015,In_3732,In_979);
or U3016 (N_3016,In_3596,In_1917);
and U3017 (N_3017,In_3732,In_3915);
nand U3018 (N_3018,In_232,In_4320);
nand U3019 (N_3019,In_4430,In_188);
or U3020 (N_3020,In_2527,In_1774);
and U3021 (N_3021,In_2067,In_1589);
nand U3022 (N_3022,In_4744,In_1343);
nor U3023 (N_3023,In_1618,In_1773);
nand U3024 (N_3024,In_4636,In_817);
and U3025 (N_3025,In_3569,In_1072);
nand U3026 (N_3026,In_284,In_3634);
xnor U3027 (N_3027,In_1206,In_4759);
or U3028 (N_3028,In_574,In_1769);
or U3029 (N_3029,In_10,In_2766);
xnor U3030 (N_3030,In_4146,In_3071);
xnor U3031 (N_3031,In_3487,In_640);
nor U3032 (N_3032,In_1554,In_913);
nor U3033 (N_3033,In_391,In_3561);
xnor U3034 (N_3034,In_569,In_365);
nand U3035 (N_3035,In_1110,In_4267);
or U3036 (N_3036,In_3544,In_1056);
xnor U3037 (N_3037,In_760,In_3850);
or U3038 (N_3038,In_579,In_1811);
nand U3039 (N_3039,In_4204,In_751);
xnor U3040 (N_3040,In_804,In_3321);
xnor U3041 (N_3041,In_2675,In_4019);
nand U3042 (N_3042,In_3737,In_3646);
nand U3043 (N_3043,In_1506,In_2100);
and U3044 (N_3044,In_122,In_2162);
or U3045 (N_3045,In_235,In_1354);
or U3046 (N_3046,In_3979,In_4613);
nand U3047 (N_3047,In_1876,In_3832);
nor U3048 (N_3048,In_3666,In_574);
xor U3049 (N_3049,In_1337,In_2813);
or U3050 (N_3050,In_4663,In_376);
or U3051 (N_3051,In_3019,In_3371);
xnor U3052 (N_3052,In_3652,In_4246);
nor U3053 (N_3053,In_4728,In_1068);
and U3054 (N_3054,In_2430,In_4593);
nor U3055 (N_3055,In_2432,In_704);
or U3056 (N_3056,In_1095,In_3258);
or U3057 (N_3057,In_175,In_1118);
or U3058 (N_3058,In_4340,In_1790);
and U3059 (N_3059,In_4396,In_804);
nand U3060 (N_3060,In_3344,In_1850);
xor U3061 (N_3061,In_577,In_3318);
nor U3062 (N_3062,In_1104,In_1135);
nand U3063 (N_3063,In_2545,In_962);
nand U3064 (N_3064,In_939,In_4273);
xnor U3065 (N_3065,In_501,In_89);
nand U3066 (N_3066,In_2968,In_51);
xor U3067 (N_3067,In_2435,In_2231);
nand U3068 (N_3068,In_2957,In_2838);
or U3069 (N_3069,In_3075,In_1566);
or U3070 (N_3070,In_3653,In_94);
xor U3071 (N_3071,In_2676,In_657);
xor U3072 (N_3072,In_2465,In_4546);
nand U3073 (N_3073,In_307,In_2799);
and U3074 (N_3074,In_4133,In_3771);
and U3075 (N_3075,In_4988,In_4818);
xnor U3076 (N_3076,In_1747,In_1317);
and U3077 (N_3077,In_2030,In_4114);
nor U3078 (N_3078,In_4539,In_2719);
or U3079 (N_3079,In_2935,In_415);
nand U3080 (N_3080,In_1627,In_427);
nor U3081 (N_3081,In_584,In_2376);
and U3082 (N_3082,In_1203,In_272);
and U3083 (N_3083,In_3682,In_4828);
and U3084 (N_3084,In_1312,In_450);
xor U3085 (N_3085,In_3986,In_1657);
nand U3086 (N_3086,In_1903,In_834);
nor U3087 (N_3087,In_1205,In_4243);
nor U3088 (N_3088,In_2165,In_4979);
nand U3089 (N_3089,In_789,In_4076);
nor U3090 (N_3090,In_130,In_2286);
and U3091 (N_3091,In_4362,In_2528);
nand U3092 (N_3092,In_3771,In_1009);
or U3093 (N_3093,In_4582,In_1988);
nor U3094 (N_3094,In_3565,In_2986);
nor U3095 (N_3095,In_2132,In_1877);
xor U3096 (N_3096,In_1497,In_982);
or U3097 (N_3097,In_2539,In_4416);
nor U3098 (N_3098,In_3981,In_2702);
and U3099 (N_3099,In_896,In_2979);
and U3100 (N_3100,In_2272,In_2836);
and U3101 (N_3101,In_3096,In_2043);
nand U3102 (N_3102,In_769,In_3344);
nand U3103 (N_3103,In_422,In_395);
or U3104 (N_3104,In_1115,In_1268);
xnor U3105 (N_3105,In_2506,In_4314);
nand U3106 (N_3106,In_3635,In_1558);
nor U3107 (N_3107,In_2439,In_3554);
xnor U3108 (N_3108,In_4983,In_4475);
or U3109 (N_3109,In_3107,In_3840);
and U3110 (N_3110,In_623,In_1426);
nand U3111 (N_3111,In_2498,In_995);
or U3112 (N_3112,In_1675,In_2225);
xnor U3113 (N_3113,In_494,In_1445);
nor U3114 (N_3114,In_1680,In_612);
or U3115 (N_3115,In_3401,In_3708);
and U3116 (N_3116,In_491,In_4388);
and U3117 (N_3117,In_4426,In_1082);
xor U3118 (N_3118,In_3101,In_1195);
nor U3119 (N_3119,In_4704,In_2599);
nor U3120 (N_3120,In_775,In_3472);
nor U3121 (N_3121,In_1932,In_3846);
nor U3122 (N_3122,In_3131,In_4839);
nor U3123 (N_3123,In_520,In_3989);
xor U3124 (N_3124,In_3118,In_4666);
or U3125 (N_3125,In_1577,In_2306);
xor U3126 (N_3126,In_3209,In_2812);
nor U3127 (N_3127,In_4083,In_3593);
and U3128 (N_3128,In_1621,In_4042);
and U3129 (N_3129,In_862,In_2093);
xor U3130 (N_3130,In_2328,In_558);
or U3131 (N_3131,In_2292,In_3931);
nand U3132 (N_3132,In_4983,In_3164);
nand U3133 (N_3133,In_2579,In_3500);
xnor U3134 (N_3134,In_262,In_3802);
nand U3135 (N_3135,In_1280,In_519);
nand U3136 (N_3136,In_4679,In_117);
or U3137 (N_3137,In_2535,In_637);
and U3138 (N_3138,In_3723,In_3152);
nand U3139 (N_3139,In_3057,In_3039);
nand U3140 (N_3140,In_2025,In_2402);
nand U3141 (N_3141,In_2472,In_2538);
nor U3142 (N_3142,In_1331,In_1808);
or U3143 (N_3143,In_4572,In_3960);
or U3144 (N_3144,In_4546,In_2269);
or U3145 (N_3145,In_117,In_2150);
nor U3146 (N_3146,In_1187,In_3735);
and U3147 (N_3147,In_2951,In_4647);
nand U3148 (N_3148,In_1949,In_1245);
or U3149 (N_3149,In_3712,In_1624);
nand U3150 (N_3150,In_1716,In_132);
nor U3151 (N_3151,In_1030,In_507);
or U3152 (N_3152,In_3804,In_4085);
xor U3153 (N_3153,In_4468,In_3369);
nand U3154 (N_3154,In_4685,In_4675);
xor U3155 (N_3155,In_2110,In_2490);
nand U3156 (N_3156,In_1335,In_4001);
xor U3157 (N_3157,In_4333,In_4467);
nand U3158 (N_3158,In_2736,In_3539);
nor U3159 (N_3159,In_210,In_1711);
and U3160 (N_3160,In_4616,In_2223);
xor U3161 (N_3161,In_3262,In_1572);
nor U3162 (N_3162,In_2427,In_268);
xnor U3163 (N_3163,In_1983,In_1193);
xor U3164 (N_3164,In_4188,In_1867);
nor U3165 (N_3165,In_4748,In_149);
nand U3166 (N_3166,In_620,In_4173);
and U3167 (N_3167,In_3702,In_2637);
nand U3168 (N_3168,In_2177,In_2847);
xor U3169 (N_3169,In_1551,In_650);
xor U3170 (N_3170,In_981,In_716);
or U3171 (N_3171,In_3584,In_4950);
xnor U3172 (N_3172,In_4675,In_3795);
xor U3173 (N_3173,In_3210,In_2276);
or U3174 (N_3174,In_393,In_3072);
or U3175 (N_3175,In_1700,In_2777);
nand U3176 (N_3176,In_4388,In_753);
nor U3177 (N_3177,In_614,In_1697);
nor U3178 (N_3178,In_1546,In_4017);
nand U3179 (N_3179,In_1242,In_2749);
xor U3180 (N_3180,In_2729,In_1201);
or U3181 (N_3181,In_1966,In_4102);
or U3182 (N_3182,In_1512,In_2312);
or U3183 (N_3183,In_198,In_3067);
nor U3184 (N_3184,In_1655,In_700);
nor U3185 (N_3185,In_4090,In_101);
and U3186 (N_3186,In_3548,In_4135);
and U3187 (N_3187,In_2294,In_2677);
and U3188 (N_3188,In_619,In_482);
and U3189 (N_3189,In_1870,In_4162);
nand U3190 (N_3190,In_2188,In_4208);
and U3191 (N_3191,In_633,In_2642);
and U3192 (N_3192,In_3908,In_2583);
nand U3193 (N_3193,In_2650,In_1994);
and U3194 (N_3194,In_4815,In_331);
or U3195 (N_3195,In_842,In_4761);
nor U3196 (N_3196,In_4331,In_503);
and U3197 (N_3197,In_1485,In_4951);
nor U3198 (N_3198,In_1997,In_1558);
xor U3199 (N_3199,In_3771,In_2499);
or U3200 (N_3200,In_3118,In_2146);
xor U3201 (N_3201,In_316,In_4932);
xnor U3202 (N_3202,In_4795,In_1468);
xor U3203 (N_3203,In_4386,In_4333);
nor U3204 (N_3204,In_1603,In_4132);
xnor U3205 (N_3205,In_107,In_4254);
xnor U3206 (N_3206,In_2904,In_2388);
and U3207 (N_3207,In_1532,In_3961);
and U3208 (N_3208,In_1979,In_4697);
nand U3209 (N_3209,In_659,In_169);
nand U3210 (N_3210,In_4168,In_3843);
xor U3211 (N_3211,In_1442,In_4647);
or U3212 (N_3212,In_974,In_4435);
nor U3213 (N_3213,In_1856,In_128);
and U3214 (N_3214,In_2115,In_2147);
xor U3215 (N_3215,In_842,In_3919);
xnor U3216 (N_3216,In_3410,In_1774);
xnor U3217 (N_3217,In_429,In_3894);
nand U3218 (N_3218,In_3849,In_4340);
or U3219 (N_3219,In_4172,In_3722);
nor U3220 (N_3220,In_3409,In_4806);
xnor U3221 (N_3221,In_3464,In_4918);
xor U3222 (N_3222,In_1298,In_3472);
or U3223 (N_3223,In_2896,In_4278);
nand U3224 (N_3224,In_1495,In_879);
and U3225 (N_3225,In_4942,In_3274);
nand U3226 (N_3226,In_16,In_3784);
or U3227 (N_3227,In_946,In_215);
and U3228 (N_3228,In_2319,In_1644);
and U3229 (N_3229,In_4351,In_649);
or U3230 (N_3230,In_4533,In_3915);
xnor U3231 (N_3231,In_1980,In_1640);
nor U3232 (N_3232,In_1994,In_2784);
xor U3233 (N_3233,In_27,In_4827);
xnor U3234 (N_3234,In_1097,In_4791);
nor U3235 (N_3235,In_3560,In_4972);
nor U3236 (N_3236,In_3666,In_1573);
xnor U3237 (N_3237,In_4209,In_2132);
nand U3238 (N_3238,In_674,In_1511);
nor U3239 (N_3239,In_703,In_3966);
nand U3240 (N_3240,In_3026,In_3426);
or U3241 (N_3241,In_3621,In_4190);
nand U3242 (N_3242,In_92,In_2150);
nand U3243 (N_3243,In_3806,In_3298);
nor U3244 (N_3244,In_1575,In_3810);
nor U3245 (N_3245,In_4391,In_1774);
xnor U3246 (N_3246,In_2137,In_4682);
nor U3247 (N_3247,In_333,In_3116);
nor U3248 (N_3248,In_4152,In_4707);
xnor U3249 (N_3249,In_1696,In_832);
xnor U3250 (N_3250,In_1798,In_729);
xnor U3251 (N_3251,In_3782,In_2020);
and U3252 (N_3252,In_1889,In_3006);
and U3253 (N_3253,In_3649,In_3909);
or U3254 (N_3254,In_1113,In_1758);
and U3255 (N_3255,In_618,In_3845);
nor U3256 (N_3256,In_2264,In_4685);
and U3257 (N_3257,In_4326,In_1020);
nand U3258 (N_3258,In_2032,In_802);
xor U3259 (N_3259,In_2833,In_1077);
or U3260 (N_3260,In_4680,In_4714);
xor U3261 (N_3261,In_3707,In_2498);
or U3262 (N_3262,In_4013,In_2656);
nand U3263 (N_3263,In_3285,In_592);
xor U3264 (N_3264,In_3558,In_4901);
nor U3265 (N_3265,In_1574,In_355);
nor U3266 (N_3266,In_3801,In_2542);
nand U3267 (N_3267,In_3198,In_1850);
nor U3268 (N_3268,In_1399,In_1679);
nand U3269 (N_3269,In_1168,In_3621);
nor U3270 (N_3270,In_1736,In_3426);
nand U3271 (N_3271,In_685,In_661);
nand U3272 (N_3272,In_4690,In_3538);
xor U3273 (N_3273,In_2336,In_916);
xnor U3274 (N_3274,In_2239,In_3330);
and U3275 (N_3275,In_3422,In_3468);
nor U3276 (N_3276,In_2065,In_2977);
nor U3277 (N_3277,In_2924,In_3821);
and U3278 (N_3278,In_2697,In_2565);
xnor U3279 (N_3279,In_4095,In_2623);
nand U3280 (N_3280,In_1355,In_3820);
nor U3281 (N_3281,In_529,In_4718);
and U3282 (N_3282,In_905,In_4452);
and U3283 (N_3283,In_1623,In_2046);
and U3284 (N_3284,In_3494,In_3596);
xor U3285 (N_3285,In_577,In_3939);
nand U3286 (N_3286,In_4847,In_4741);
xor U3287 (N_3287,In_2125,In_2672);
xor U3288 (N_3288,In_3004,In_3614);
xnor U3289 (N_3289,In_1150,In_2042);
and U3290 (N_3290,In_923,In_4625);
nor U3291 (N_3291,In_4160,In_2912);
nand U3292 (N_3292,In_2561,In_2134);
or U3293 (N_3293,In_2221,In_2403);
or U3294 (N_3294,In_3660,In_308);
or U3295 (N_3295,In_3713,In_2115);
and U3296 (N_3296,In_824,In_4868);
and U3297 (N_3297,In_1257,In_2312);
xor U3298 (N_3298,In_2836,In_2703);
xnor U3299 (N_3299,In_1962,In_552);
nor U3300 (N_3300,In_11,In_1384);
or U3301 (N_3301,In_2685,In_183);
xnor U3302 (N_3302,In_136,In_1836);
xor U3303 (N_3303,In_1958,In_2885);
nand U3304 (N_3304,In_931,In_2561);
nand U3305 (N_3305,In_138,In_851);
and U3306 (N_3306,In_4808,In_3273);
xnor U3307 (N_3307,In_3393,In_1198);
nor U3308 (N_3308,In_4214,In_510);
and U3309 (N_3309,In_3414,In_4796);
and U3310 (N_3310,In_573,In_2311);
nand U3311 (N_3311,In_2854,In_4801);
xor U3312 (N_3312,In_3222,In_4211);
or U3313 (N_3313,In_1342,In_2514);
or U3314 (N_3314,In_2732,In_384);
nor U3315 (N_3315,In_2252,In_3066);
and U3316 (N_3316,In_4556,In_1973);
nor U3317 (N_3317,In_4983,In_1798);
and U3318 (N_3318,In_2625,In_528);
and U3319 (N_3319,In_2517,In_4246);
xor U3320 (N_3320,In_2945,In_517);
or U3321 (N_3321,In_544,In_3856);
xor U3322 (N_3322,In_589,In_358);
nor U3323 (N_3323,In_3063,In_2587);
nor U3324 (N_3324,In_2224,In_3470);
nor U3325 (N_3325,In_1803,In_3601);
or U3326 (N_3326,In_409,In_4913);
nor U3327 (N_3327,In_1062,In_4124);
nor U3328 (N_3328,In_821,In_2876);
nor U3329 (N_3329,In_1149,In_679);
nand U3330 (N_3330,In_143,In_3870);
nor U3331 (N_3331,In_2285,In_3675);
nand U3332 (N_3332,In_1453,In_2572);
xor U3333 (N_3333,In_1600,In_1181);
and U3334 (N_3334,In_4532,In_721);
or U3335 (N_3335,In_4488,In_323);
and U3336 (N_3336,In_3215,In_4551);
nand U3337 (N_3337,In_4474,In_1361);
nand U3338 (N_3338,In_497,In_1479);
xor U3339 (N_3339,In_4219,In_4703);
and U3340 (N_3340,In_4579,In_1811);
nand U3341 (N_3341,In_1059,In_659);
nor U3342 (N_3342,In_1304,In_4024);
or U3343 (N_3343,In_1190,In_105);
nand U3344 (N_3344,In_2358,In_4852);
xor U3345 (N_3345,In_4320,In_2740);
and U3346 (N_3346,In_2831,In_2819);
or U3347 (N_3347,In_1442,In_50);
or U3348 (N_3348,In_2312,In_3056);
or U3349 (N_3349,In_2779,In_3710);
nand U3350 (N_3350,In_958,In_1644);
xor U3351 (N_3351,In_1412,In_3155);
or U3352 (N_3352,In_1520,In_4743);
nand U3353 (N_3353,In_749,In_1214);
or U3354 (N_3354,In_1940,In_2780);
xor U3355 (N_3355,In_1422,In_4600);
and U3356 (N_3356,In_2708,In_1019);
xnor U3357 (N_3357,In_2723,In_2356);
nand U3358 (N_3358,In_359,In_127);
nor U3359 (N_3359,In_4604,In_4542);
nand U3360 (N_3360,In_4582,In_789);
nand U3361 (N_3361,In_1615,In_555);
xnor U3362 (N_3362,In_2941,In_2853);
and U3363 (N_3363,In_1343,In_3);
xor U3364 (N_3364,In_3022,In_3664);
and U3365 (N_3365,In_4539,In_1570);
and U3366 (N_3366,In_93,In_1622);
or U3367 (N_3367,In_2554,In_1432);
nor U3368 (N_3368,In_1632,In_3888);
xor U3369 (N_3369,In_1865,In_2013);
and U3370 (N_3370,In_3791,In_4410);
and U3371 (N_3371,In_1521,In_3003);
nor U3372 (N_3372,In_3154,In_870);
and U3373 (N_3373,In_471,In_2619);
nor U3374 (N_3374,In_3281,In_4537);
xor U3375 (N_3375,In_1507,In_2221);
nor U3376 (N_3376,In_4265,In_3133);
xnor U3377 (N_3377,In_1869,In_979);
nand U3378 (N_3378,In_3067,In_656);
and U3379 (N_3379,In_3622,In_442);
or U3380 (N_3380,In_3378,In_1500);
nand U3381 (N_3381,In_3567,In_4546);
nand U3382 (N_3382,In_4103,In_4434);
nor U3383 (N_3383,In_4960,In_3169);
and U3384 (N_3384,In_4930,In_116);
and U3385 (N_3385,In_1637,In_4220);
nor U3386 (N_3386,In_4042,In_3292);
nand U3387 (N_3387,In_2082,In_1134);
nor U3388 (N_3388,In_4506,In_3861);
and U3389 (N_3389,In_2401,In_4858);
nand U3390 (N_3390,In_1387,In_3684);
or U3391 (N_3391,In_4608,In_2562);
nand U3392 (N_3392,In_2328,In_3673);
or U3393 (N_3393,In_4123,In_3778);
nor U3394 (N_3394,In_3214,In_1884);
xor U3395 (N_3395,In_3164,In_3962);
and U3396 (N_3396,In_2226,In_2371);
nor U3397 (N_3397,In_77,In_4050);
or U3398 (N_3398,In_3325,In_2770);
and U3399 (N_3399,In_4165,In_1534);
and U3400 (N_3400,In_1138,In_1882);
nand U3401 (N_3401,In_4150,In_3826);
nor U3402 (N_3402,In_2985,In_3783);
and U3403 (N_3403,In_4328,In_3745);
and U3404 (N_3404,In_896,In_2700);
nand U3405 (N_3405,In_2038,In_4282);
nor U3406 (N_3406,In_2586,In_2743);
or U3407 (N_3407,In_3567,In_4363);
nor U3408 (N_3408,In_4135,In_1307);
nand U3409 (N_3409,In_1382,In_4161);
nand U3410 (N_3410,In_214,In_3340);
xnor U3411 (N_3411,In_1050,In_3354);
xor U3412 (N_3412,In_556,In_3864);
or U3413 (N_3413,In_2334,In_3511);
nand U3414 (N_3414,In_3328,In_836);
nand U3415 (N_3415,In_4302,In_1456);
or U3416 (N_3416,In_4355,In_170);
or U3417 (N_3417,In_4503,In_235);
xor U3418 (N_3418,In_4230,In_1724);
nor U3419 (N_3419,In_2221,In_4077);
and U3420 (N_3420,In_202,In_2392);
or U3421 (N_3421,In_2760,In_4185);
xor U3422 (N_3422,In_3001,In_3480);
and U3423 (N_3423,In_3242,In_214);
nand U3424 (N_3424,In_1750,In_3511);
nand U3425 (N_3425,In_2969,In_4090);
nor U3426 (N_3426,In_2404,In_1552);
and U3427 (N_3427,In_658,In_4536);
nor U3428 (N_3428,In_366,In_2258);
nand U3429 (N_3429,In_2432,In_1279);
nand U3430 (N_3430,In_2412,In_1513);
or U3431 (N_3431,In_455,In_3118);
xor U3432 (N_3432,In_2172,In_2412);
nor U3433 (N_3433,In_3696,In_1714);
nand U3434 (N_3434,In_640,In_880);
or U3435 (N_3435,In_331,In_3677);
nor U3436 (N_3436,In_4630,In_4657);
nand U3437 (N_3437,In_1544,In_4651);
or U3438 (N_3438,In_3188,In_4841);
nand U3439 (N_3439,In_260,In_121);
xnor U3440 (N_3440,In_2601,In_2564);
nand U3441 (N_3441,In_3333,In_4844);
and U3442 (N_3442,In_3668,In_2124);
nand U3443 (N_3443,In_759,In_1695);
and U3444 (N_3444,In_1300,In_280);
nand U3445 (N_3445,In_4921,In_2045);
or U3446 (N_3446,In_3261,In_4645);
and U3447 (N_3447,In_4791,In_174);
nor U3448 (N_3448,In_3838,In_3217);
nand U3449 (N_3449,In_4932,In_1442);
or U3450 (N_3450,In_3068,In_4088);
or U3451 (N_3451,In_1096,In_973);
nor U3452 (N_3452,In_3206,In_4999);
xor U3453 (N_3453,In_608,In_3900);
xnor U3454 (N_3454,In_3340,In_3056);
nor U3455 (N_3455,In_1041,In_75);
xor U3456 (N_3456,In_1027,In_1770);
nor U3457 (N_3457,In_545,In_748);
xor U3458 (N_3458,In_4592,In_3907);
nand U3459 (N_3459,In_4476,In_3828);
or U3460 (N_3460,In_1689,In_4602);
xor U3461 (N_3461,In_1014,In_3540);
and U3462 (N_3462,In_2082,In_455);
and U3463 (N_3463,In_2295,In_1413);
nor U3464 (N_3464,In_2398,In_3784);
nand U3465 (N_3465,In_1043,In_4615);
nor U3466 (N_3466,In_4166,In_1881);
xnor U3467 (N_3467,In_470,In_3399);
xnor U3468 (N_3468,In_3318,In_4628);
and U3469 (N_3469,In_294,In_801);
xor U3470 (N_3470,In_4831,In_280);
nand U3471 (N_3471,In_828,In_1866);
or U3472 (N_3472,In_2144,In_3018);
or U3473 (N_3473,In_730,In_3731);
and U3474 (N_3474,In_178,In_531);
nand U3475 (N_3475,In_4431,In_2609);
xor U3476 (N_3476,In_1324,In_2104);
nor U3477 (N_3477,In_1361,In_4927);
nand U3478 (N_3478,In_3034,In_987);
nor U3479 (N_3479,In_3814,In_2121);
and U3480 (N_3480,In_3054,In_2465);
nor U3481 (N_3481,In_4460,In_2801);
and U3482 (N_3482,In_553,In_490);
or U3483 (N_3483,In_3569,In_1992);
and U3484 (N_3484,In_4665,In_4839);
nand U3485 (N_3485,In_3341,In_778);
and U3486 (N_3486,In_2695,In_992);
or U3487 (N_3487,In_211,In_872);
and U3488 (N_3488,In_1035,In_4317);
or U3489 (N_3489,In_693,In_3492);
and U3490 (N_3490,In_4156,In_2971);
xnor U3491 (N_3491,In_4411,In_4225);
or U3492 (N_3492,In_767,In_3314);
and U3493 (N_3493,In_4005,In_4063);
and U3494 (N_3494,In_2330,In_3257);
nand U3495 (N_3495,In_4212,In_985);
nor U3496 (N_3496,In_1748,In_4899);
nor U3497 (N_3497,In_893,In_889);
and U3498 (N_3498,In_2774,In_630);
and U3499 (N_3499,In_2011,In_3872);
xnor U3500 (N_3500,In_3621,In_1997);
or U3501 (N_3501,In_553,In_2225);
nor U3502 (N_3502,In_2609,In_2581);
xnor U3503 (N_3503,In_840,In_3324);
xor U3504 (N_3504,In_4396,In_3541);
nor U3505 (N_3505,In_1313,In_797);
nand U3506 (N_3506,In_332,In_2197);
xnor U3507 (N_3507,In_1072,In_471);
and U3508 (N_3508,In_2320,In_1793);
xor U3509 (N_3509,In_3974,In_2477);
nor U3510 (N_3510,In_1757,In_178);
nand U3511 (N_3511,In_4882,In_2632);
or U3512 (N_3512,In_3691,In_3610);
nand U3513 (N_3513,In_2362,In_4372);
or U3514 (N_3514,In_2413,In_4762);
xnor U3515 (N_3515,In_3622,In_4664);
xnor U3516 (N_3516,In_1245,In_1941);
or U3517 (N_3517,In_1868,In_777);
and U3518 (N_3518,In_790,In_1175);
nor U3519 (N_3519,In_1315,In_3445);
or U3520 (N_3520,In_4046,In_3763);
nor U3521 (N_3521,In_4240,In_2384);
nand U3522 (N_3522,In_4763,In_24);
nor U3523 (N_3523,In_2228,In_1304);
nand U3524 (N_3524,In_4223,In_3668);
or U3525 (N_3525,In_4122,In_4979);
nand U3526 (N_3526,In_1668,In_4491);
xnor U3527 (N_3527,In_4863,In_534);
and U3528 (N_3528,In_42,In_198);
nor U3529 (N_3529,In_4502,In_1453);
xnor U3530 (N_3530,In_3315,In_4755);
xor U3531 (N_3531,In_1591,In_1746);
xor U3532 (N_3532,In_1761,In_2150);
xnor U3533 (N_3533,In_1135,In_2678);
and U3534 (N_3534,In_2036,In_2564);
nand U3535 (N_3535,In_3004,In_4215);
nand U3536 (N_3536,In_2929,In_3160);
and U3537 (N_3537,In_1817,In_4557);
xor U3538 (N_3538,In_654,In_4845);
or U3539 (N_3539,In_4300,In_3057);
xor U3540 (N_3540,In_4068,In_4212);
nor U3541 (N_3541,In_1585,In_4208);
and U3542 (N_3542,In_1390,In_1926);
xor U3543 (N_3543,In_679,In_71);
nand U3544 (N_3544,In_1272,In_4225);
and U3545 (N_3545,In_1585,In_1300);
nor U3546 (N_3546,In_2964,In_3747);
nand U3547 (N_3547,In_1254,In_2490);
xor U3548 (N_3548,In_701,In_2729);
xor U3549 (N_3549,In_349,In_2238);
nor U3550 (N_3550,In_2559,In_729);
and U3551 (N_3551,In_3355,In_4416);
nor U3552 (N_3552,In_859,In_4048);
xor U3553 (N_3553,In_4103,In_624);
nand U3554 (N_3554,In_2613,In_428);
xor U3555 (N_3555,In_4181,In_1198);
nor U3556 (N_3556,In_2259,In_3108);
nand U3557 (N_3557,In_645,In_2158);
or U3558 (N_3558,In_3832,In_1579);
or U3559 (N_3559,In_1272,In_1681);
xor U3560 (N_3560,In_2442,In_4256);
or U3561 (N_3561,In_406,In_1911);
nand U3562 (N_3562,In_4893,In_2444);
and U3563 (N_3563,In_2953,In_2582);
nand U3564 (N_3564,In_4462,In_1425);
xnor U3565 (N_3565,In_4656,In_4336);
nor U3566 (N_3566,In_2096,In_1061);
and U3567 (N_3567,In_3664,In_4503);
or U3568 (N_3568,In_1093,In_3467);
xnor U3569 (N_3569,In_2098,In_2577);
xnor U3570 (N_3570,In_4176,In_4449);
and U3571 (N_3571,In_4445,In_20);
and U3572 (N_3572,In_3645,In_3397);
nor U3573 (N_3573,In_2718,In_947);
and U3574 (N_3574,In_3197,In_4967);
and U3575 (N_3575,In_2683,In_199);
or U3576 (N_3576,In_3979,In_912);
nand U3577 (N_3577,In_2698,In_1006);
nand U3578 (N_3578,In_4600,In_4086);
nand U3579 (N_3579,In_922,In_21);
xnor U3580 (N_3580,In_3897,In_453);
nand U3581 (N_3581,In_2287,In_2761);
xnor U3582 (N_3582,In_3313,In_72);
nand U3583 (N_3583,In_400,In_383);
xor U3584 (N_3584,In_4458,In_4301);
and U3585 (N_3585,In_4601,In_4522);
or U3586 (N_3586,In_3169,In_1248);
xor U3587 (N_3587,In_2141,In_1217);
and U3588 (N_3588,In_4543,In_2981);
or U3589 (N_3589,In_4115,In_910);
nand U3590 (N_3590,In_3640,In_4641);
and U3591 (N_3591,In_4651,In_4183);
nand U3592 (N_3592,In_1751,In_41);
nand U3593 (N_3593,In_3781,In_563);
or U3594 (N_3594,In_219,In_990);
nor U3595 (N_3595,In_1834,In_2803);
nor U3596 (N_3596,In_1812,In_4827);
or U3597 (N_3597,In_406,In_670);
xor U3598 (N_3598,In_4541,In_3025);
and U3599 (N_3599,In_2050,In_736);
or U3600 (N_3600,In_200,In_225);
nand U3601 (N_3601,In_3650,In_1811);
and U3602 (N_3602,In_1181,In_1937);
nor U3603 (N_3603,In_385,In_17);
and U3604 (N_3604,In_1257,In_1482);
nand U3605 (N_3605,In_85,In_411);
nor U3606 (N_3606,In_3088,In_650);
or U3607 (N_3607,In_4590,In_204);
and U3608 (N_3608,In_3968,In_433);
nand U3609 (N_3609,In_1924,In_949);
nor U3610 (N_3610,In_3307,In_1824);
xnor U3611 (N_3611,In_4947,In_276);
xor U3612 (N_3612,In_3046,In_3702);
or U3613 (N_3613,In_3790,In_2738);
and U3614 (N_3614,In_848,In_1647);
and U3615 (N_3615,In_1711,In_393);
nand U3616 (N_3616,In_597,In_451);
nand U3617 (N_3617,In_2058,In_3710);
and U3618 (N_3618,In_202,In_2556);
nor U3619 (N_3619,In_2361,In_3157);
nand U3620 (N_3620,In_2834,In_4520);
or U3621 (N_3621,In_1342,In_1743);
or U3622 (N_3622,In_4464,In_4316);
nor U3623 (N_3623,In_4710,In_807);
xnor U3624 (N_3624,In_1293,In_902);
nor U3625 (N_3625,In_1513,In_279);
or U3626 (N_3626,In_2682,In_50);
or U3627 (N_3627,In_2499,In_917);
or U3628 (N_3628,In_199,In_4688);
xnor U3629 (N_3629,In_2182,In_3086);
or U3630 (N_3630,In_1864,In_300);
and U3631 (N_3631,In_4563,In_2261);
or U3632 (N_3632,In_4311,In_1019);
or U3633 (N_3633,In_1724,In_842);
and U3634 (N_3634,In_1783,In_1744);
or U3635 (N_3635,In_1728,In_1507);
nand U3636 (N_3636,In_1046,In_1374);
xnor U3637 (N_3637,In_1266,In_1909);
nand U3638 (N_3638,In_836,In_521);
and U3639 (N_3639,In_1188,In_1605);
xnor U3640 (N_3640,In_1858,In_3503);
and U3641 (N_3641,In_1949,In_4850);
xnor U3642 (N_3642,In_727,In_217);
nor U3643 (N_3643,In_3591,In_4834);
or U3644 (N_3644,In_1585,In_3098);
nor U3645 (N_3645,In_2840,In_4871);
or U3646 (N_3646,In_2538,In_1975);
nand U3647 (N_3647,In_4252,In_4879);
or U3648 (N_3648,In_472,In_2250);
xor U3649 (N_3649,In_963,In_4503);
nor U3650 (N_3650,In_649,In_1206);
or U3651 (N_3651,In_4006,In_436);
xnor U3652 (N_3652,In_3722,In_3041);
nand U3653 (N_3653,In_844,In_1187);
and U3654 (N_3654,In_456,In_2253);
nand U3655 (N_3655,In_1581,In_3124);
nand U3656 (N_3656,In_3129,In_4405);
or U3657 (N_3657,In_2492,In_925);
xnor U3658 (N_3658,In_4581,In_3037);
nor U3659 (N_3659,In_352,In_1252);
nor U3660 (N_3660,In_2480,In_1758);
nor U3661 (N_3661,In_3497,In_3158);
and U3662 (N_3662,In_2688,In_1107);
nand U3663 (N_3663,In_4899,In_4879);
xor U3664 (N_3664,In_4695,In_4812);
nor U3665 (N_3665,In_4485,In_347);
xnor U3666 (N_3666,In_3926,In_1664);
or U3667 (N_3667,In_4256,In_1573);
and U3668 (N_3668,In_2515,In_4868);
and U3669 (N_3669,In_143,In_4336);
nor U3670 (N_3670,In_1019,In_4105);
and U3671 (N_3671,In_3178,In_1980);
nand U3672 (N_3672,In_72,In_3233);
or U3673 (N_3673,In_894,In_1932);
xor U3674 (N_3674,In_2065,In_4581);
and U3675 (N_3675,In_554,In_3953);
nand U3676 (N_3676,In_2002,In_3834);
and U3677 (N_3677,In_3267,In_390);
xor U3678 (N_3678,In_3165,In_4100);
xnor U3679 (N_3679,In_2166,In_4085);
nand U3680 (N_3680,In_1383,In_4855);
or U3681 (N_3681,In_2679,In_2243);
nand U3682 (N_3682,In_355,In_4473);
nor U3683 (N_3683,In_1284,In_2130);
xor U3684 (N_3684,In_432,In_4981);
nand U3685 (N_3685,In_619,In_2310);
or U3686 (N_3686,In_4683,In_195);
nor U3687 (N_3687,In_1402,In_484);
nor U3688 (N_3688,In_2420,In_1264);
nand U3689 (N_3689,In_2064,In_430);
nor U3690 (N_3690,In_1034,In_2884);
or U3691 (N_3691,In_4084,In_4337);
or U3692 (N_3692,In_4488,In_4094);
or U3693 (N_3693,In_3555,In_291);
nor U3694 (N_3694,In_2167,In_4315);
and U3695 (N_3695,In_3664,In_4138);
nand U3696 (N_3696,In_3273,In_385);
or U3697 (N_3697,In_679,In_4620);
nand U3698 (N_3698,In_1841,In_2493);
xnor U3699 (N_3699,In_1989,In_3614);
or U3700 (N_3700,In_3365,In_1277);
xor U3701 (N_3701,In_3539,In_3554);
nand U3702 (N_3702,In_3855,In_1828);
or U3703 (N_3703,In_4838,In_1842);
nor U3704 (N_3704,In_1246,In_736);
nand U3705 (N_3705,In_3604,In_1830);
xnor U3706 (N_3706,In_1574,In_1357);
nand U3707 (N_3707,In_3744,In_3409);
nand U3708 (N_3708,In_3858,In_1883);
nand U3709 (N_3709,In_2635,In_1348);
nand U3710 (N_3710,In_439,In_4402);
nor U3711 (N_3711,In_3680,In_12);
xnor U3712 (N_3712,In_2811,In_4938);
or U3713 (N_3713,In_2907,In_4555);
and U3714 (N_3714,In_2565,In_2437);
nand U3715 (N_3715,In_519,In_4474);
or U3716 (N_3716,In_781,In_3562);
nor U3717 (N_3717,In_2219,In_3051);
nor U3718 (N_3718,In_3859,In_2646);
nor U3719 (N_3719,In_1333,In_537);
nor U3720 (N_3720,In_3209,In_1226);
or U3721 (N_3721,In_3901,In_2039);
nand U3722 (N_3722,In_258,In_3260);
or U3723 (N_3723,In_105,In_4560);
and U3724 (N_3724,In_3268,In_2396);
nor U3725 (N_3725,In_778,In_48);
nand U3726 (N_3726,In_1615,In_577);
xor U3727 (N_3727,In_3048,In_2127);
xnor U3728 (N_3728,In_1051,In_2262);
and U3729 (N_3729,In_2697,In_1074);
xnor U3730 (N_3730,In_4489,In_3779);
nor U3731 (N_3731,In_1533,In_3612);
or U3732 (N_3732,In_1655,In_4057);
nand U3733 (N_3733,In_373,In_2344);
nand U3734 (N_3734,In_351,In_4816);
or U3735 (N_3735,In_65,In_753);
nor U3736 (N_3736,In_765,In_4016);
nand U3737 (N_3737,In_4165,In_4092);
or U3738 (N_3738,In_4982,In_3350);
or U3739 (N_3739,In_1459,In_3084);
xnor U3740 (N_3740,In_3688,In_566);
nor U3741 (N_3741,In_2225,In_2764);
and U3742 (N_3742,In_4704,In_1723);
nor U3743 (N_3743,In_4231,In_2788);
nor U3744 (N_3744,In_4999,In_3441);
xor U3745 (N_3745,In_703,In_3302);
nor U3746 (N_3746,In_4777,In_1488);
xor U3747 (N_3747,In_4392,In_1786);
nor U3748 (N_3748,In_4826,In_1665);
or U3749 (N_3749,In_2505,In_2691);
nor U3750 (N_3750,In_1621,In_4803);
or U3751 (N_3751,In_3624,In_761);
and U3752 (N_3752,In_1165,In_629);
and U3753 (N_3753,In_3742,In_1833);
and U3754 (N_3754,In_4739,In_3892);
or U3755 (N_3755,In_4542,In_3116);
xnor U3756 (N_3756,In_2671,In_1014);
xor U3757 (N_3757,In_375,In_1789);
nor U3758 (N_3758,In_1030,In_2168);
nor U3759 (N_3759,In_376,In_4058);
and U3760 (N_3760,In_786,In_2048);
or U3761 (N_3761,In_332,In_193);
or U3762 (N_3762,In_416,In_1244);
and U3763 (N_3763,In_100,In_3117);
nor U3764 (N_3764,In_4567,In_72);
or U3765 (N_3765,In_2976,In_45);
or U3766 (N_3766,In_3174,In_2602);
and U3767 (N_3767,In_720,In_3031);
or U3768 (N_3768,In_3154,In_4491);
or U3769 (N_3769,In_3539,In_2457);
xnor U3770 (N_3770,In_1348,In_4459);
and U3771 (N_3771,In_4598,In_4732);
nor U3772 (N_3772,In_2400,In_4378);
nor U3773 (N_3773,In_4850,In_2988);
nor U3774 (N_3774,In_4780,In_623);
or U3775 (N_3775,In_4837,In_986);
nand U3776 (N_3776,In_1641,In_3958);
or U3777 (N_3777,In_2899,In_2530);
xor U3778 (N_3778,In_4031,In_3293);
nor U3779 (N_3779,In_1219,In_3750);
nand U3780 (N_3780,In_1752,In_1719);
and U3781 (N_3781,In_2005,In_847);
nor U3782 (N_3782,In_4425,In_3278);
xor U3783 (N_3783,In_4673,In_3710);
nor U3784 (N_3784,In_3345,In_4596);
xnor U3785 (N_3785,In_4145,In_727);
nor U3786 (N_3786,In_4800,In_2957);
and U3787 (N_3787,In_460,In_188);
xnor U3788 (N_3788,In_2428,In_1435);
nand U3789 (N_3789,In_457,In_3562);
xor U3790 (N_3790,In_457,In_493);
xor U3791 (N_3791,In_3044,In_4926);
or U3792 (N_3792,In_4001,In_2857);
or U3793 (N_3793,In_4249,In_2028);
nand U3794 (N_3794,In_0,In_2591);
or U3795 (N_3795,In_1345,In_655);
and U3796 (N_3796,In_1916,In_504);
nand U3797 (N_3797,In_2960,In_3769);
and U3798 (N_3798,In_1992,In_3749);
nand U3799 (N_3799,In_3699,In_1168);
or U3800 (N_3800,In_3521,In_3770);
and U3801 (N_3801,In_4923,In_244);
nor U3802 (N_3802,In_2820,In_4704);
nor U3803 (N_3803,In_905,In_1335);
nor U3804 (N_3804,In_1492,In_4439);
nand U3805 (N_3805,In_3432,In_979);
nor U3806 (N_3806,In_1219,In_4201);
nand U3807 (N_3807,In_76,In_4671);
nor U3808 (N_3808,In_4884,In_3401);
nor U3809 (N_3809,In_1314,In_2568);
and U3810 (N_3810,In_1054,In_2422);
xor U3811 (N_3811,In_969,In_1591);
and U3812 (N_3812,In_1447,In_865);
nor U3813 (N_3813,In_1580,In_1751);
and U3814 (N_3814,In_1013,In_1052);
xnor U3815 (N_3815,In_3296,In_40);
xor U3816 (N_3816,In_3411,In_4653);
nand U3817 (N_3817,In_3435,In_202);
and U3818 (N_3818,In_2739,In_1859);
or U3819 (N_3819,In_3811,In_4855);
xor U3820 (N_3820,In_2082,In_4672);
and U3821 (N_3821,In_1110,In_3142);
and U3822 (N_3822,In_2409,In_654);
nand U3823 (N_3823,In_2292,In_2323);
nand U3824 (N_3824,In_3035,In_982);
nor U3825 (N_3825,In_449,In_1491);
and U3826 (N_3826,In_4536,In_4915);
xnor U3827 (N_3827,In_1218,In_599);
or U3828 (N_3828,In_3405,In_2860);
or U3829 (N_3829,In_760,In_4073);
xnor U3830 (N_3830,In_3684,In_1495);
and U3831 (N_3831,In_1879,In_617);
or U3832 (N_3832,In_3567,In_4996);
and U3833 (N_3833,In_3342,In_2158);
nor U3834 (N_3834,In_518,In_2963);
xor U3835 (N_3835,In_4927,In_472);
and U3836 (N_3836,In_1306,In_4240);
nor U3837 (N_3837,In_3609,In_1133);
nor U3838 (N_3838,In_1705,In_3229);
nand U3839 (N_3839,In_1795,In_230);
xor U3840 (N_3840,In_2288,In_3776);
or U3841 (N_3841,In_4334,In_2239);
nand U3842 (N_3842,In_1373,In_1793);
nor U3843 (N_3843,In_1052,In_1817);
nor U3844 (N_3844,In_2909,In_2855);
xor U3845 (N_3845,In_4641,In_4662);
and U3846 (N_3846,In_2417,In_3186);
nand U3847 (N_3847,In_1732,In_2679);
xor U3848 (N_3848,In_1173,In_2741);
and U3849 (N_3849,In_2665,In_2805);
nor U3850 (N_3850,In_3930,In_2260);
nand U3851 (N_3851,In_2673,In_3548);
or U3852 (N_3852,In_3650,In_3218);
nor U3853 (N_3853,In_3582,In_1204);
or U3854 (N_3854,In_599,In_4148);
and U3855 (N_3855,In_2405,In_1074);
xor U3856 (N_3856,In_3317,In_3725);
xor U3857 (N_3857,In_33,In_1953);
or U3858 (N_3858,In_3699,In_1633);
xor U3859 (N_3859,In_1187,In_2638);
nand U3860 (N_3860,In_2859,In_3538);
nor U3861 (N_3861,In_2565,In_1618);
nor U3862 (N_3862,In_4811,In_2218);
and U3863 (N_3863,In_3178,In_1030);
nand U3864 (N_3864,In_2259,In_1020);
nand U3865 (N_3865,In_1913,In_916);
and U3866 (N_3866,In_4554,In_2227);
nand U3867 (N_3867,In_4936,In_1521);
nand U3868 (N_3868,In_4727,In_4213);
and U3869 (N_3869,In_4604,In_1940);
or U3870 (N_3870,In_3171,In_286);
xnor U3871 (N_3871,In_4926,In_726);
or U3872 (N_3872,In_2214,In_4672);
nand U3873 (N_3873,In_3748,In_937);
or U3874 (N_3874,In_3749,In_4739);
xor U3875 (N_3875,In_367,In_2428);
nor U3876 (N_3876,In_2837,In_3021);
xnor U3877 (N_3877,In_3913,In_1536);
and U3878 (N_3878,In_3398,In_3688);
or U3879 (N_3879,In_4355,In_1497);
xnor U3880 (N_3880,In_2093,In_4934);
nor U3881 (N_3881,In_2994,In_3623);
nor U3882 (N_3882,In_154,In_2728);
nor U3883 (N_3883,In_2724,In_1258);
nor U3884 (N_3884,In_4480,In_2188);
and U3885 (N_3885,In_504,In_3112);
or U3886 (N_3886,In_4925,In_917);
nand U3887 (N_3887,In_4964,In_1167);
and U3888 (N_3888,In_4972,In_1032);
and U3889 (N_3889,In_3449,In_2025);
or U3890 (N_3890,In_2877,In_1224);
nand U3891 (N_3891,In_283,In_663);
nor U3892 (N_3892,In_3329,In_1340);
and U3893 (N_3893,In_1973,In_2754);
xnor U3894 (N_3894,In_4440,In_4747);
and U3895 (N_3895,In_493,In_4735);
nand U3896 (N_3896,In_676,In_2377);
and U3897 (N_3897,In_4638,In_218);
or U3898 (N_3898,In_3059,In_837);
xor U3899 (N_3899,In_2871,In_360);
xor U3900 (N_3900,In_902,In_2626);
and U3901 (N_3901,In_2654,In_2552);
nand U3902 (N_3902,In_670,In_3670);
or U3903 (N_3903,In_3708,In_3958);
xnor U3904 (N_3904,In_3738,In_2475);
xor U3905 (N_3905,In_4987,In_1442);
nand U3906 (N_3906,In_1876,In_4393);
or U3907 (N_3907,In_3601,In_4734);
and U3908 (N_3908,In_2661,In_3889);
or U3909 (N_3909,In_1103,In_1530);
and U3910 (N_3910,In_3511,In_2900);
and U3911 (N_3911,In_3233,In_2964);
and U3912 (N_3912,In_2290,In_3550);
nor U3913 (N_3913,In_337,In_1459);
nor U3914 (N_3914,In_1613,In_3472);
nor U3915 (N_3915,In_3807,In_4729);
nand U3916 (N_3916,In_1572,In_2094);
nand U3917 (N_3917,In_3455,In_3126);
nand U3918 (N_3918,In_3391,In_4607);
and U3919 (N_3919,In_3944,In_1531);
nor U3920 (N_3920,In_1408,In_3435);
nand U3921 (N_3921,In_3086,In_244);
and U3922 (N_3922,In_2144,In_285);
and U3923 (N_3923,In_1526,In_4041);
or U3924 (N_3924,In_4141,In_4733);
nor U3925 (N_3925,In_1964,In_4198);
xnor U3926 (N_3926,In_3238,In_4057);
nor U3927 (N_3927,In_4706,In_197);
nand U3928 (N_3928,In_839,In_3356);
or U3929 (N_3929,In_4135,In_1574);
xnor U3930 (N_3930,In_4868,In_2403);
nand U3931 (N_3931,In_4627,In_3840);
nand U3932 (N_3932,In_2865,In_3351);
or U3933 (N_3933,In_3325,In_595);
xor U3934 (N_3934,In_1606,In_3845);
xor U3935 (N_3935,In_4730,In_3092);
nor U3936 (N_3936,In_3074,In_2940);
xnor U3937 (N_3937,In_119,In_4821);
or U3938 (N_3938,In_1559,In_1504);
or U3939 (N_3939,In_1613,In_1406);
nand U3940 (N_3940,In_3115,In_656);
xor U3941 (N_3941,In_3162,In_1975);
or U3942 (N_3942,In_3553,In_2869);
and U3943 (N_3943,In_279,In_4309);
xor U3944 (N_3944,In_4573,In_317);
xnor U3945 (N_3945,In_2251,In_4839);
nand U3946 (N_3946,In_4162,In_4116);
and U3947 (N_3947,In_4183,In_1377);
xnor U3948 (N_3948,In_3358,In_4937);
nand U3949 (N_3949,In_3308,In_2543);
nand U3950 (N_3950,In_2121,In_4325);
xor U3951 (N_3951,In_2226,In_1656);
xor U3952 (N_3952,In_2429,In_740);
nor U3953 (N_3953,In_4387,In_2710);
and U3954 (N_3954,In_4021,In_3055);
nand U3955 (N_3955,In_4603,In_1267);
and U3956 (N_3956,In_3484,In_1386);
and U3957 (N_3957,In_4744,In_155);
nor U3958 (N_3958,In_4133,In_2771);
xnor U3959 (N_3959,In_3476,In_600);
nor U3960 (N_3960,In_1061,In_4996);
nor U3961 (N_3961,In_3115,In_2803);
xor U3962 (N_3962,In_3252,In_2903);
nor U3963 (N_3963,In_206,In_4632);
nand U3964 (N_3964,In_3840,In_3170);
xor U3965 (N_3965,In_4981,In_2511);
or U3966 (N_3966,In_3458,In_462);
nand U3967 (N_3967,In_1219,In_3779);
nand U3968 (N_3968,In_3455,In_4577);
xnor U3969 (N_3969,In_2472,In_1504);
or U3970 (N_3970,In_973,In_4828);
xnor U3971 (N_3971,In_295,In_1357);
nor U3972 (N_3972,In_3080,In_3939);
nor U3973 (N_3973,In_3247,In_3617);
xnor U3974 (N_3974,In_2030,In_4688);
nand U3975 (N_3975,In_2856,In_2905);
or U3976 (N_3976,In_3508,In_2409);
xnor U3977 (N_3977,In_4066,In_1204);
nand U3978 (N_3978,In_1033,In_1787);
nand U3979 (N_3979,In_1765,In_4946);
nor U3980 (N_3980,In_2720,In_3397);
nor U3981 (N_3981,In_4469,In_2528);
nor U3982 (N_3982,In_588,In_4685);
or U3983 (N_3983,In_4282,In_634);
nor U3984 (N_3984,In_625,In_1896);
nand U3985 (N_3985,In_822,In_809);
nor U3986 (N_3986,In_4675,In_3412);
xor U3987 (N_3987,In_1749,In_1063);
or U3988 (N_3988,In_4799,In_4798);
nand U3989 (N_3989,In_1673,In_2388);
nand U3990 (N_3990,In_1236,In_1661);
or U3991 (N_3991,In_865,In_937);
or U3992 (N_3992,In_4833,In_2935);
nor U3993 (N_3993,In_154,In_4606);
nor U3994 (N_3994,In_301,In_3641);
and U3995 (N_3995,In_2714,In_2010);
or U3996 (N_3996,In_3677,In_1488);
nand U3997 (N_3997,In_4795,In_806);
nand U3998 (N_3998,In_209,In_1817);
nand U3999 (N_3999,In_573,In_4916);
nor U4000 (N_4000,In_88,In_1734);
or U4001 (N_4001,In_3665,In_266);
nor U4002 (N_4002,In_1967,In_4097);
or U4003 (N_4003,In_1996,In_330);
or U4004 (N_4004,In_3237,In_4527);
nand U4005 (N_4005,In_648,In_2041);
xor U4006 (N_4006,In_221,In_2540);
and U4007 (N_4007,In_2968,In_2510);
xnor U4008 (N_4008,In_1456,In_1515);
nor U4009 (N_4009,In_3254,In_3457);
or U4010 (N_4010,In_2717,In_1912);
nand U4011 (N_4011,In_980,In_393);
or U4012 (N_4012,In_3492,In_4464);
or U4013 (N_4013,In_1193,In_4459);
or U4014 (N_4014,In_3301,In_4810);
and U4015 (N_4015,In_2471,In_1878);
and U4016 (N_4016,In_2618,In_1673);
nand U4017 (N_4017,In_3328,In_604);
or U4018 (N_4018,In_3666,In_2349);
nand U4019 (N_4019,In_3575,In_1588);
or U4020 (N_4020,In_1877,In_3313);
xor U4021 (N_4021,In_2589,In_3696);
or U4022 (N_4022,In_2941,In_2569);
and U4023 (N_4023,In_2086,In_4134);
nand U4024 (N_4024,In_3350,In_3549);
nand U4025 (N_4025,In_24,In_2862);
or U4026 (N_4026,In_1608,In_2670);
nand U4027 (N_4027,In_4944,In_3378);
nand U4028 (N_4028,In_2921,In_3683);
nor U4029 (N_4029,In_4758,In_4313);
nand U4030 (N_4030,In_1987,In_2360);
and U4031 (N_4031,In_4983,In_189);
nor U4032 (N_4032,In_1262,In_4252);
or U4033 (N_4033,In_2079,In_742);
nor U4034 (N_4034,In_490,In_4804);
and U4035 (N_4035,In_2310,In_4958);
xnor U4036 (N_4036,In_2343,In_290);
nand U4037 (N_4037,In_1416,In_764);
nor U4038 (N_4038,In_4565,In_3757);
nor U4039 (N_4039,In_3070,In_3697);
or U4040 (N_4040,In_1017,In_2275);
nor U4041 (N_4041,In_3766,In_4624);
nand U4042 (N_4042,In_1720,In_1798);
nor U4043 (N_4043,In_2636,In_4171);
xnor U4044 (N_4044,In_1688,In_1450);
nor U4045 (N_4045,In_377,In_3530);
nor U4046 (N_4046,In_908,In_1006);
nand U4047 (N_4047,In_3985,In_3271);
and U4048 (N_4048,In_3731,In_2821);
nand U4049 (N_4049,In_3969,In_943);
and U4050 (N_4050,In_1162,In_3515);
and U4051 (N_4051,In_4327,In_4491);
nand U4052 (N_4052,In_943,In_4726);
nand U4053 (N_4053,In_2904,In_3031);
xor U4054 (N_4054,In_531,In_4749);
xnor U4055 (N_4055,In_450,In_1571);
xnor U4056 (N_4056,In_2162,In_1419);
or U4057 (N_4057,In_2956,In_3346);
or U4058 (N_4058,In_1000,In_2487);
xnor U4059 (N_4059,In_1162,In_2144);
nor U4060 (N_4060,In_3523,In_3474);
and U4061 (N_4061,In_1161,In_2164);
xnor U4062 (N_4062,In_767,In_3647);
or U4063 (N_4063,In_2930,In_3655);
or U4064 (N_4064,In_2608,In_701);
xnor U4065 (N_4065,In_968,In_2747);
and U4066 (N_4066,In_4734,In_2638);
nand U4067 (N_4067,In_784,In_749);
and U4068 (N_4068,In_1948,In_2490);
or U4069 (N_4069,In_1244,In_302);
or U4070 (N_4070,In_4824,In_2172);
or U4071 (N_4071,In_3059,In_201);
and U4072 (N_4072,In_3395,In_2231);
xnor U4073 (N_4073,In_3258,In_3330);
or U4074 (N_4074,In_4932,In_1635);
xor U4075 (N_4075,In_3204,In_1741);
or U4076 (N_4076,In_368,In_564);
nor U4077 (N_4077,In_2705,In_3296);
or U4078 (N_4078,In_3113,In_110);
or U4079 (N_4079,In_4234,In_3186);
nand U4080 (N_4080,In_4150,In_1610);
xor U4081 (N_4081,In_4848,In_1312);
or U4082 (N_4082,In_2609,In_1068);
nand U4083 (N_4083,In_3739,In_4062);
and U4084 (N_4084,In_2840,In_2088);
or U4085 (N_4085,In_3358,In_1947);
nor U4086 (N_4086,In_706,In_690);
nand U4087 (N_4087,In_1223,In_2597);
nand U4088 (N_4088,In_88,In_1136);
nand U4089 (N_4089,In_2868,In_357);
or U4090 (N_4090,In_3062,In_3525);
nand U4091 (N_4091,In_438,In_3782);
and U4092 (N_4092,In_331,In_4307);
xor U4093 (N_4093,In_1622,In_1362);
nor U4094 (N_4094,In_2723,In_1449);
nand U4095 (N_4095,In_1789,In_3907);
xor U4096 (N_4096,In_4426,In_1557);
xor U4097 (N_4097,In_3661,In_2468);
xor U4098 (N_4098,In_4019,In_1077);
nor U4099 (N_4099,In_2111,In_214);
xnor U4100 (N_4100,In_4052,In_3167);
or U4101 (N_4101,In_3952,In_1559);
nand U4102 (N_4102,In_1527,In_1565);
and U4103 (N_4103,In_262,In_3713);
xor U4104 (N_4104,In_3549,In_3575);
and U4105 (N_4105,In_2275,In_1858);
nand U4106 (N_4106,In_4337,In_2093);
xnor U4107 (N_4107,In_4853,In_1024);
nand U4108 (N_4108,In_2951,In_30);
xor U4109 (N_4109,In_3769,In_3409);
nor U4110 (N_4110,In_830,In_31);
and U4111 (N_4111,In_1178,In_2097);
xor U4112 (N_4112,In_3483,In_2068);
nor U4113 (N_4113,In_318,In_851);
nor U4114 (N_4114,In_1104,In_378);
nor U4115 (N_4115,In_1972,In_783);
nor U4116 (N_4116,In_1917,In_134);
nor U4117 (N_4117,In_3885,In_4290);
xor U4118 (N_4118,In_3205,In_306);
or U4119 (N_4119,In_3656,In_560);
nor U4120 (N_4120,In_4003,In_4181);
xor U4121 (N_4121,In_3484,In_4409);
and U4122 (N_4122,In_460,In_2828);
nor U4123 (N_4123,In_2697,In_4974);
xor U4124 (N_4124,In_2324,In_2562);
xnor U4125 (N_4125,In_4210,In_2008);
and U4126 (N_4126,In_2603,In_3631);
xnor U4127 (N_4127,In_1084,In_3956);
or U4128 (N_4128,In_3710,In_1440);
xnor U4129 (N_4129,In_824,In_3758);
nand U4130 (N_4130,In_4408,In_2737);
or U4131 (N_4131,In_3947,In_2056);
and U4132 (N_4132,In_1914,In_57);
xor U4133 (N_4133,In_1628,In_4138);
xor U4134 (N_4134,In_3193,In_1908);
and U4135 (N_4135,In_2370,In_1957);
nand U4136 (N_4136,In_698,In_892);
and U4137 (N_4137,In_2739,In_2748);
xor U4138 (N_4138,In_1972,In_3802);
nor U4139 (N_4139,In_2281,In_1626);
nor U4140 (N_4140,In_3570,In_897);
and U4141 (N_4141,In_3039,In_2372);
or U4142 (N_4142,In_4300,In_568);
and U4143 (N_4143,In_3902,In_4607);
or U4144 (N_4144,In_336,In_488);
xor U4145 (N_4145,In_1092,In_1882);
or U4146 (N_4146,In_3762,In_2764);
and U4147 (N_4147,In_2672,In_2443);
nor U4148 (N_4148,In_310,In_3952);
xor U4149 (N_4149,In_930,In_610);
xor U4150 (N_4150,In_4169,In_2131);
or U4151 (N_4151,In_3082,In_141);
nor U4152 (N_4152,In_3753,In_2869);
nor U4153 (N_4153,In_252,In_714);
or U4154 (N_4154,In_215,In_3206);
nand U4155 (N_4155,In_235,In_2711);
and U4156 (N_4156,In_2279,In_1624);
or U4157 (N_4157,In_4221,In_831);
nor U4158 (N_4158,In_2644,In_2642);
or U4159 (N_4159,In_1108,In_2012);
and U4160 (N_4160,In_3964,In_4794);
nor U4161 (N_4161,In_4963,In_1343);
and U4162 (N_4162,In_3555,In_447);
nor U4163 (N_4163,In_468,In_3274);
xnor U4164 (N_4164,In_3450,In_4033);
nor U4165 (N_4165,In_4780,In_702);
xnor U4166 (N_4166,In_710,In_1801);
nand U4167 (N_4167,In_4120,In_104);
xor U4168 (N_4168,In_2429,In_4775);
xor U4169 (N_4169,In_3651,In_3189);
nor U4170 (N_4170,In_2615,In_2286);
nand U4171 (N_4171,In_3818,In_1056);
nor U4172 (N_4172,In_2646,In_4427);
nand U4173 (N_4173,In_2826,In_1116);
or U4174 (N_4174,In_1395,In_1075);
xnor U4175 (N_4175,In_2847,In_3834);
nand U4176 (N_4176,In_4016,In_2250);
xnor U4177 (N_4177,In_1112,In_1014);
or U4178 (N_4178,In_4379,In_1222);
or U4179 (N_4179,In_3975,In_1401);
and U4180 (N_4180,In_152,In_167);
and U4181 (N_4181,In_3290,In_2335);
nor U4182 (N_4182,In_4110,In_4883);
xnor U4183 (N_4183,In_4211,In_1670);
or U4184 (N_4184,In_3127,In_3255);
nor U4185 (N_4185,In_1483,In_2858);
nand U4186 (N_4186,In_4259,In_4883);
and U4187 (N_4187,In_214,In_4653);
or U4188 (N_4188,In_2083,In_1760);
or U4189 (N_4189,In_4544,In_3350);
nor U4190 (N_4190,In_63,In_606);
xnor U4191 (N_4191,In_1176,In_54);
nand U4192 (N_4192,In_1025,In_4831);
and U4193 (N_4193,In_328,In_2587);
nor U4194 (N_4194,In_2626,In_2605);
and U4195 (N_4195,In_1630,In_2295);
or U4196 (N_4196,In_4573,In_130);
nand U4197 (N_4197,In_339,In_2889);
or U4198 (N_4198,In_3297,In_1087);
xnor U4199 (N_4199,In_2578,In_2648);
and U4200 (N_4200,In_945,In_2010);
xnor U4201 (N_4201,In_3016,In_4046);
nor U4202 (N_4202,In_4613,In_2450);
and U4203 (N_4203,In_4144,In_3685);
nand U4204 (N_4204,In_1360,In_2458);
or U4205 (N_4205,In_3475,In_3399);
nand U4206 (N_4206,In_4405,In_1867);
and U4207 (N_4207,In_1673,In_943);
nor U4208 (N_4208,In_1300,In_1981);
nand U4209 (N_4209,In_226,In_3691);
or U4210 (N_4210,In_1243,In_3658);
nor U4211 (N_4211,In_798,In_1980);
nor U4212 (N_4212,In_3848,In_2464);
nor U4213 (N_4213,In_4715,In_3212);
xnor U4214 (N_4214,In_4282,In_2817);
nand U4215 (N_4215,In_4911,In_3137);
nor U4216 (N_4216,In_2374,In_3991);
nor U4217 (N_4217,In_4602,In_3910);
and U4218 (N_4218,In_2386,In_4047);
nand U4219 (N_4219,In_3577,In_4105);
or U4220 (N_4220,In_1527,In_794);
nor U4221 (N_4221,In_77,In_572);
or U4222 (N_4222,In_2670,In_1713);
xnor U4223 (N_4223,In_654,In_3140);
nand U4224 (N_4224,In_2637,In_2195);
and U4225 (N_4225,In_268,In_168);
nor U4226 (N_4226,In_1459,In_2490);
nor U4227 (N_4227,In_4287,In_340);
nor U4228 (N_4228,In_316,In_759);
nand U4229 (N_4229,In_3504,In_1455);
xor U4230 (N_4230,In_4294,In_1962);
and U4231 (N_4231,In_4217,In_1192);
or U4232 (N_4232,In_2050,In_2804);
nand U4233 (N_4233,In_1833,In_3175);
nand U4234 (N_4234,In_4833,In_230);
or U4235 (N_4235,In_233,In_25);
nor U4236 (N_4236,In_186,In_237);
and U4237 (N_4237,In_3190,In_1825);
nand U4238 (N_4238,In_4029,In_1049);
xor U4239 (N_4239,In_144,In_446);
nand U4240 (N_4240,In_3850,In_2970);
nand U4241 (N_4241,In_3371,In_486);
and U4242 (N_4242,In_1802,In_2061);
xor U4243 (N_4243,In_3026,In_2277);
or U4244 (N_4244,In_659,In_2122);
or U4245 (N_4245,In_2191,In_812);
or U4246 (N_4246,In_3897,In_4726);
and U4247 (N_4247,In_2955,In_4451);
and U4248 (N_4248,In_516,In_2021);
and U4249 (N_4249,In_861,In_150);
xor U4250 (N_4250,In_1958,In_3276);
nor U4251 (N_4251,In_706,In_2372);
and U4252 (N_4252,In_1620,In_1345);
nor U4253 (N_4253,In_3423,In_3086);
or U4254 (N_4254,In_357,In_2353);
nor U4255 (N_4255,In_39,In_153);
or U4256 (N_4256,In_4508,In_4028);
nor U4257 (N_4257,In_4681,In_1598);
xor U4258 (N_4258,In_514,In_2538);
or U4259 (N_4259,In_2600,In_1649);
and U4260 (N_4260,In_1213,In_3217);
nor U4261 (N_4261,In_3036,In_2332);
nand U4262 (N_4262,In_4865,In_570);
nor U4263 (N_4263,In_946,In_4598);
nor U4264 (N_4264,In_1011,In_1533);
nand U4265 (N_4265,In_1750,In_3899);
or U4266 (N_4266,In_413,In_457);
nor U4267 (N_4267,In_4487,In_3274);
nor U4268 (N_4268,In_2457,In_4492);
xnor U4269 (N_4269,In_2662,In_200);
and U4270 (N_4270,In_1138,In_3527);
xnor U4271 (N_4271,In_3001,In_4172);
or U4272 (N_4272,In_546,In_3091);
xnor U4273 (N_4273,In_4650,In_4186);
and U4274 (N_4274,In_227,In_2294);
xnor U4275 (N_4275,In_4685,In_246);
xnor U4276 (N_4276,In_441,In_1427);
or U4277 (N_4277,In_691,In_3416);
and U4278 (N_4278,In_4328,In_118);
xnor U4279 (N_4279,In_4669,In_37);
and U4280 (N_4280,In_1548,In_4824);
and U4281 (N_4281,In_547,In_1875);
nor U4282 (N_4282,In_886,In_4672);
xnor U4283 (N_4283,In_1770,In_1451);
and U4284 (N_4284,In_2011,In_2676);
nor U4285 (N_4285,In_3959,In_3973);
or U4286 (N_4286,In_946,In_1659);
or U4287 (N_4287,In_3355,In_2854);
nand U4288 (N_4288,In_1282,In_4535);
nor U4289 (N_4289,In_3744,In_2804);
nand U4290 (N_4290,In_1005,In_934);
and U4291 (N_4291,In_3999,In_2923);
or U4292 (N_4292,In_4021,In_2709);
or U4293 (N_4293,In_1264,In_3096);
and U4294 (N_4294,In_3511,In_180);
nor U4295 (N_4295,In_568,In_926);
nor U4296 (N_4296,In_1436,In_4391);
nor U4297 (N_4297,In_1340,In_2940);
or U4298 (N_4298,In_2752,In_4805);
or U4299 (N_4299,In_4707,In_2892);
nand U4300 (N_4300,In_522,In_2728);
nand U4301 (N_4301,In_35,In_3715);
nand U4302 (N_4302,In_1322,In_2987);
nor U4303 (N_4303,In_4037,In_567);
or U4304 (N_4304,In_2008,In_1824);
nor U4305 (N_4305,In_3055,In_2865);
nor U4306 (N_4306,In_4992,In_1783);
or U4307 (N_4307,In_4214,In_1777);
or U4308 (N_4308,In_841,In_4488);
xor U4309 (N_4309,In_3281,In_2827);
or U4310 (N_4310,In_134,In_1123);
nor U4311 (N_4311,In_804,In_3377);
nand U4312 (N_4312,In_916,In_808);
nor U4313 (N_4313,In_4748,In_4740);
and U4314 (N_4314,In_4599,In_1886);
or U4315 (N_4315,In_1830,In_385);
or U4316 (N_4316,In_3829,In_4493);
or U4317 (N_4317,In_3999,In_644);
xnor U4318 (N_4318,In_4056,In_1827);
and U4319 (N_4319,In_1810,In_1821);
nand U4320 (N_4320,In_4174,In_2730);
nand U4321 (N_4321,In_391,In_3938);
xor U4322 (N_4322,In_4455,In_2690);
xor U4323 (N_4323,In_3309,In_4448);
nor U4324 (N_4324,In_3106,In_2789);
and U4325 (N_4325,In_2459,In_3776);
and U4326 (N_4326,In_1881,In_4825);
xor U4327 (N_4327,In_597,In_3227);
nand U4328 (N_4328,In_2656,In_2000);
and U4329 (N_4329,In_559,In_1250);
nor U4330 (N_4330,In_3939,In_3732);
or U4331 (N_4331,In_4962,In_864);
and U4332 (N_4332,In_1504,In_1854);
xor U4333 (N_4333,In_4631,In_3586);
or U4334 (N_4334,In_2026,In_686);
xnor U4335 (N_4335,In_2926,In_2264);
or U4336 (N_4336,In_2888,In_420);
nor U4337 (N_4337,In_1565,In_3899);
and U4338 (N_4338,In_5,In_4276);
nor U4339 (N_4339,In_1105,In_4797);
xnor U4340 (N_4340,In_4105,In_4207);
xor U4341 (N_4341,In_4396,In_2635);
or U4342 (N_4342,In_1746,In_3448);
nand U4343 (N_4343,In_2058,In_2798);
nor U4344 (N_4344,In_4602,In_2460);
or U4345 (N_4345,In_812,In_4494);
nor U4346 (N_4346,In_254,In_1534);
and U4347 (N_4347,In_3626,In_4443);
and U4348 (N_4348,In_1476,In_4351);
and U4349 (N_4349,In_2581,In_3359);
xor U4350 (N_4350,In_3667,In_2788);
xor U4351 (N_4351,In_4779,In_1459);
xnor U4352 (N_4352,In_4108,In_2361);
nor U4353 (N_4353,In_3840,In_3971);
nor U4354 (N_4354,In_4935,In_1692);
nand U4355 (N_4355,In_1487,In_4431);
nor U4356 (N_4356,In_4459,In_4964);
nand U4357 (N_4357,In_4194,In_261);
nor U4358 (N_4358,In_5,In_2730);
and U4359 (N_4359,In_598,In_1133);
and U4360 (N_4360,In_1834,In_1240);
xor U4361 (N_4361,In_254,In_2148);
or U4362 (N_4362,In_3918,In_563);
nor U4363 (N_4363,In_2487,In_3209);
nand U4364 (N_4364,In_1409,In_3595);
or U4365 (N_4365,In_2440,In_1546);
nand U4366 (N_4366,In_3193,In_1989);
xnor U4367 (N_4367,In_1853,In_4198);
xnor U4368 (N_4368,In_1229,In_1997);
nor U4369 (N_4369,In_3513,In_3099);
xor U4370 (N_4370,In_2143,In_862);
and U4371 (N_4371,In_359,In_4460);
nor U4372 (N_4372,In_3903,In_4578);
and U4373 (N_4373,In_4532,In_1519);
xor U4374 (N_4374,In_3390,In_4959);
and U4375 (N_4375,In_2066,In_1307);
nor U4376 (N_4376,In_3549,In_689);
or U4377 (N_4377,In_3625,In_4248);
nand U4378 (N_4378,In_581,In_1074);
and U4379 (N_4379,In_4725,In_68);
nand U4380 (N_4380,In_3047,In_1711);
nand U4381 (N_4381,In_457,In_799);
and U4382 (N_4382,In_1470,In_158);
or U4383 (N_4383,In_2864,In_3892);
and U4384 (N_4384,In_265,In_3518);
nand U4385 (N_4385,In_1026,In_2744);
or U4386 (N_4386,In_3665,In_2819);
nor U4387 (N_4387,In_2388,In_2766);
or U4388 (N_4388,In_3935,In_462);
and U4389 (N_4389,In_2291,In_1297);
or U4390 (N_4390,In_4460,In_3545);
xnor U4391 (N_4391,In_1334,In_3010);
nand U4392 (N_4392,In_3350,In_4529);
nor U4393 (N_4393,In_3006,In_2458);
or U4394 (N_4394,In_887,In_4615);
or U4395 (N_4395,In_413,In_2092);
and U4396 (N_4396,In_3025,In_1370);
and U4397 (N_4397,In_578,In_1091);
or U4398 (N_4398,In_1774,In_1313);
nand U4399 (N_4399,In_3028,In_1305);
nor U4400 (N_4400,In_3782,In_106);
or U4401 (N_4401,In_2088,In_1117);
xor U4402 (N_4402,In_736,In_4175);
xnor U4403 (N_4403,In_1084,In_3965);
and U4404 (N_4404,In_3674,In_1148);
nand U4405 (N_4405,In_1329,In_671);
xnor U4406 (N_4406,In_4119,In_2260);
and U4407 (N_4407,In_2503,In_300);
xnor U4408 (N_4408,In_2692,In_3817);
xnor U4409 (N_4409,In_1012,In_2469);
and U4410 (N_4410,In_745,In_1629);
and U4411 (N_4411,In_793,In_826);
nor U4412 (N_4412,In_26,In_1631);
xnor U4413 (N_4413,In_1309,In_2551);
and U4414 (N_4414,In_1124,In_2600);
and U4415 (N_4415,In_4290,In_4245);
xnor U4416 (N_4416,In_2051,In_1069);
or U4417 (N_4417,In_1433,In_3715);
and U4418 (N_4418,In_3857,In_917);
or U4419 (N_4419,In_4303,In_4049);
nor U4420 (N_4420,In_1952,In_3887);
or U4421 (N_4421,In_2005,In_4958);
nand U4422 (N_4422,In_3082,In_4369);
xnor U4423 (N_4423,In_1863,In_719);
and U4424 (N_4424,In_2798,In_3054);
xor U4425 (N_4425,In_2712,In_2881);
nand U4426 (N_4426,In_323,In_2513);
and U4427 (N_4427,In_1554,In_4796);
nand U4428 (N_4428,In_2609,In_4371);
xnor U4429 (N_4429,In_549,In_4621);
nand U4430 (N_4430,In_1377,In_2711);
xor U4431 (N_4431,In_2753,In_3833);
and U4432 (N_4432,In_4852,In_11);
nand U4433 (N_4433,In_3135,In_817);
nor U4434 (N_4434,In_2381,In_3860);
nor U4435 (N_4435,In_2494,In_146);
nand U4436 (N_4436,In_3522,In_2350);
xnor U4437 (N_4437,In_3353,In_1999);
nand U4438 (N_4438,In_1787,In_1308);
xor U4439 (N_4439,In_1373,In_2652);
and U4440 (N_4440,In_4493,In_4116);
nor U4441 (N_4441,In_2095,In_3441);
nand U4442 (N_4442,In_935,In_4514);
nand U4443 (N_4443,In_1248,In_949);
nor U4444 (N_4444,In_4276,In_408);
nor U4445 (N_4445,In_3059,In_1052);
nand U4446 (N_4446,In_4302,In_2586);
nand U4447 (N_4447,In_1664,In_3957);
nand U4448 (N_4448,In_864,In_140);
or U4449 (N_4449,In_1741,In_2525);
and U4450 (N_4450,In_2512,In_1330);
nor U4451 (N_4451,In_328,In_235);
nand U4452 (N_4452,In_2376,In_2763);
and U4453 (N_4453,In_281,In_2194);
or U4454 (N_4454,In_4497,In_963);
and U4455 (N_4455,In_758,In_2582);
nand U4456 (N_4456,In_2501,In_4342);
or U4457 (N_4457,In_2733,In_1453);
nor U4458 (N_4458,In_4441,In_2583);
nor U4459 (N_4459,In_2238,In_3827);
or U4460 (N_4460,In_2212,In_3263);
nor U4461 (N_4461,In_430,In_969);
and U4462 (N_4462,In_3940,In_1862);
or U4463 (N_4463,In_2875,In_3115);
or U4464 (N_4464,In_2688,In_3664);
and U4465 (N_4465,In_2574,In_657);
nand U4466 (N_4466,In_1365,In_168);
or U4467 (N_4467,In_2574,In_2604);
nand U4468 (N_4468,In_682,In_2048);
nand U4469 (N_4469,In_1624,In_3625);
or U4470 (N_4470,In_2251,In_2414);
and U4471 (N_4471,In_3100,In_524);
xnor U4472 (N_4472,In_3728,In_3676);
or U4473 (N_4473,In_1970,In_3674);
xnor U4474 (N_4474,In_2569,In_2972);
nand U4475 (N_4475,In_4024,In_2055);
nor U4476 (N_4476,In_4545,In_1078);
nand U4477 (N_4477,In_66,In_3770);
nand U4478 (N_4478,In_1634,In_3002);
and U4479 (N_4479,In_308,In_4159);
and U4480 (N_4480,In_2861,In_2039);
or U4481 (N_4481,In_1689,In_4197);
or U4482 (N_4482,In_1192,In_3755);
and U4483 (N_4483,In_3379,In_4175);
or U4484 (N_4484,In_2372,In_1248);
and U4485 (N_4485,In_2704,In_3033);
nand U4486 (N_4486,In_3041,In_4919);
nor U4487 (N_4487,In_3353,In_3410);
xnor U4488 (N_4488,In_4575,In_1444);
and U4489 (N_4489,In_912,In_2970);
and U4490 (N_4490,In_3060,In_716);
and U4491 (N_4491,In_4215,In_7);
and U4492 (N_4492,In_3297,In_3114);
and U4493 (N_4493,In_777,In_1279);
nor U4494 (N_4494,In_1966,In_1353);
nor U4495 (N_4495,In_3449,In_4805);
xnor U4496 (N_4496,In_3403,In_1142);
xor U4497 (N_4497,In_1240,In_1631);
or U4498 (N_4498,In_3107,In_3090);
or U4499 (N_4499,In_3730,In_4121);
nand U4500 (N_4500,In_4658,In_1931);
or U4501 (N_4501,In_1205,In_767);
xor U4502 (N_4502,In_2338,In_2230);
and U4503 (N_4503,In_4060,In_2577);
or U4504 (N_4504,In_1956,In_314);
nor U4505 (N_4505,In_924,In_3372);
or U4506 (N_4506,In_1739,In_1769);
nor U4507 (N_4507,In_853,In_3622);
xor U4508 (N_4508,In_3537,In_2923);
xor U4509 (N_4509,In_4787,In_540);
and U4510 (N_4510,In_4955,In_2548);
nor U4511 (N_4511,In_2701,In_1209);
or U4512 (N_4512,In_4324,In_1223);
and U4513 (N_4513,In_1229,In_4204);
and U4514 (N_4514,In_1078,In_2845);
nor U4515 (N_4515,In_2042,In_1728);
nor U4516 (N_4516,In_4847,In_3416);
xor U4517 (N_4517,In_908,In_1094);
nor U4518 (N_4518,In_3228,In_2298);
and U4519 (N_4519,In_2212,In_791);
nand U4520 (N_4520,In_3362,In_196);
nor U4521 (N_4521,In_3530,In_3879);
nor U4522 (N_4522,In_1375,In_2050);
nand U4523 (N_4523,In_3670,In_1037);
and U4524 (N_4524,In_4262,In_4309);
nor U4525 (N_4525,In_883,In_4692);
nand U4526 (N_4526,In_4585,In_1337);
nor U4527 (N_4527,In_2741,In_4881);
xor U4528 (N_4528,In_2396,In_3719);
or U4529 (N_4529,In_2151,In_3763);
and U4530 (N_4530,In_916,In_4926);
nor U4531 (N_4531,In_891,In_4528);
or U4532 (N_4532,In_1804,In_2626);
xnor U4533 (N_4533,In_2733,In_1312);
nand U4534 (N_4534,In_2947,In_755);
nand U4535 (N_4535,In_3778,In_2553);
nor U4536 (N_4536,In_4154,In_1937);
xor U4537 (N_4537,In_1088,In_3943);
or U4538 (N_4538,In_2457,In_183);
nand U4539 (N_4539,In_3498,In_2262);
xnor U4540 (N_4540,In_74,In_4818);
and U4541 (N_4541,In_2338,In_801);
nor U4542 (N_4542,In_1826,In_1815);
xnor U4543 (N_4543,In_962,In_2394);
nor U4544 (N_4544,In_1967,In_3716);
nor U4545 (N_4545,In_3249,In_4831);
nor U4546 (N_4546,In_903,In_947);
or U4547 (N_4547,In_4466,In_4706);
xnor U4548 (N_4548,In_3227,In_2953);
nor U4549 (N_4549,In_2902,In_1555);
nor U4550 (N_4550,In_3108,In_711);
or U4551 (N_4551,In_3426,In_2305);
xor U4552 (N_4552,In_2857,In_1996);
xor U4553 (N_4553,In_3402,In_1756);
xnor U4554 (N_4554,In_2034,In_2123);
and U4555 (N_4555,In_4488,In_1129);
and U4556 (N_4556,In_3152,In_3885);
nor U4557 (N_4557,In_4681,In_1281);
or U4558 (N_4558,In_495,In_1586);
nand U4559 (N_4559,In_695,In_4156);
and U4560 (N_4560,In_4701,In_2128);
and U4561 (N_4561,In_2531,In_2273);
or U4562 (N_4562,In_2746,In_1295);
nor U4563 (N_4563,In_687,In_2237);
or U4564 (N_4564,In_2936,In_2142);
xnor U4565 (N_4565,In_288,In_1727);
and U4566 (N_4566,In_4137,In_3069);
nor U4567 (N_4567,In_3050,In_66);
nor U4568 (N_4568,In_104,In_4290);
xnor U4569 (N_4569,In_3484,In_2501);
and U4570 (N_4570,In_532,In_4283);
nand U4571 (N_4571,In_753,In_3048);
nand U4572 (N_4572,In_1084,In_50);
nand U4573 (N_4573,In_4523,In_476);
or U4574 (N_4574,In_1698,In_4165);
xnor U4575 (N_4575,In_1442,In_4697);
nor U4576 (N_4576,In_2761,In_2762);
nor U4577 (N_4577,In_3982,In_4190);
nand U4578 (N_4578,In_2361,In_4017);
xor U4579 (N_4579,In_443,In_4342);
nand U4580 (N_4580,In_2138,In_1061);
xnor U4581 (N_4581,In_1539,In_4606);
or U4582 (N_4582,In_4427,In_4050);
or U4583 (N_4583,In_1472,In_4176);
nand U4584 (N_4584,In_1449,In_1178);
nor U4585 (N_4585,In_2698,In_1377);
or U4586 (N_4586,In_3489,In_2689);
xnor U4587 (N_4587,In_4632,In_4897);
nor U4588 (N_4588,In_4331,In_3543);
nor U4589 (N_4589,In_2575,In_2392);
and U4590 (N_4590,In_3755,In_940);
or U4591 (N_4591,In_661,In_2866);
xor U4592 (N_4592,In_2452,In_1858);
nand U4593 (N_4593,In_2360,In_2436);
or U4594 (N_4594,In_1845,In_1798);
or U4595 (N_4595,In_4725,In_1908);
nor U4596 (N_4596,In_2091,In_3564);
or U4597 (N_4597,In_4940,In_850);
xor U4598 (N_4598,In_2867,In_2204);
nand U4599 (N_4599,In_1696,In_3850);
and U4600 (N_4600,In_849,In_3162);
or U4601 (N_4601,In_4292,In_4981);
nand U4602 (N_4602,In_122,In_2013);
nor U4603 (N_4603,In_947,In_2156);
nand U4604 (N_4604,In_4900,In_4241);
or U4605 (N_4605,In_2174,In_396);
nor U4606 (N_4606,In_437,In_2166);
nand U4607 (N_4607,In_254,In_3618);
and U4608 (N_4608,In_2792,In_3024);
nand U4609 (N_4609,In_515,In_1356);
nand U4610 (N_4610,In_4278,In_1615);
and U4611 (N_4611,In_2549,In_4000);
xor U4612 (N_4612,In_690,In_4043);
xor U4613 (N_4613,In_1193,In_2515);
and U4614 (N_4614,In_3796,In_243);
nor U4615 (N_4615,In_2024,In_3721);
xnor U4616 (N_4616,In_4464,In_4616);
or U4617 (N_4617,In_592,In_3327);
or U4618 (N_4618,In_947,In_60);
nand U4619 (N_4619,In_4016,In_2344);
nand U4620 (N_4620,In_3760,In_1621);
or U4621 (N_4621,In_1792,In_635);
and U4622 (N_4622,In_97,In_2644);
nor U4623 (N_4623,In_1461,In_2662);
nand U4624 (N_4624,In_2930,In_1899);
xnor U4625 (N_4625,In_3831,In_872);
and U4626 (N_4626,In_3991,In_2823);
and U4627 (N_4627,In_4776,In_3515);
nor U4628 (N_4628,In_3545,In_3916);
xor U4629 (N_4629,In_1584,In_2027);
and U4630 (N_4630,In_1068,In_43);
xnor U4631 (N_4631,In_4328,In_4044);
nand U4632 (N_4632,In_3041,In_2628);
nand U4633 (N_4633,In_3423,In_3777);
nand U4634 (N_4634,In_4860,In_4138);
nand U4635 (N_4635,In_1849,In_4268);
and U4636 (N_4636,In_4979,In_1250);
nor U4637 (N_4637,In_335,In_952);
xor U4638 (N_4638,In_4543,In_2147);
nor U4639 (N_4639,In_2963,In_4145);
xnor U4640 (N_4640,In_3110,In_1412);
nand U4641 (N_4641,In_3667,In_1076);
or U4642 (N_4642,In_2053,In_2555);
and U4643 (N_4643,In_2699,In_1466);
or U4644 (N_4644,In_1666,In_2794);
xnor U4645 (N_4645,In_186,In_3);
xnor U4646 (N_4646,In_4834,In_1609);
xor U4647 (N_4647,In_3533,In_4080);
nor U4648 (N_4648,In_3354,In_346);
nor U4649 (N_4649,In_4048,In_177);
xnor U4650 (N_4650,In_2362,In_3100);
nand U4651 (N_4651,In_1218,In_2636);
xnor U4652 (N_4652,In_3672,In_4021);
nand U4653 (N_4653,In_2167,In_4102);
or U4654 (N_4654,In_2097,In_4399);
and U4655 (N_4655,In_2726,In_4);
xnor U4656 (N_4656,In_706,In_1011);
xnor U4657 (N_4657,In_839,In_2175);
xor U4658 (N_4658,In_3026,In_2666);
or U4659 (N_4659,In_3939,In_3504);
nand U4660 (N_4660,In_4733,In_4014);
xor U4661 (N_4661,In_3239,In_319);
nand U4662 (N_4662,In_2668,In_1271);
or U4663 (N_4663,In_1091,In_4656);
nor U4664 (N_4664,In_47,In_1204);
or U4665 (N_4665,In_243,In_2016);
xor U4666 (N_4666,In_950,In_3790);
xnor U4667 (N_4667,In_2084,In_1893);
nand U4668 (N_4668,In_3502,In_1095);
or U4669 (N_4669,In_2975,In_2409);
nand U4670 (N_4670,In_650,In_460);
or U4671 (N_4671,In_2266,In_4597);
nand U4672 (N_4672,In_762,In_2201);
xor U4673 (N_4673,In_3479,In_1621);
nand U4674 (N_4674,In_4418,In_4375);
or U4675 (N_4675,In_2757,In_3074);
nand U4676 (N_4676,In_3622,In_344);
and U4677 (N_4677,In_3799,In_1181);
or U4678 (N_4678,In_2585,In_3904);
nand U4679 (N_4679,In_1999,In_3233);
or U4680 (N_4680,In_330,In_787);
or U4681 (N_4681,In_1729,In_3583);
nand U4682 (N_4682,In_2278,In_2840);
nand U4683 (N_4683,In_3648,In_1933);
nor U4684 (N_4684,In_4200,In_4527);
nand U4685 (N_4685,In_3731,In_4624);
or U4686 (N_4686,In_741,In_1091);
or U4687 (N_4687,In_3530,In_4782);
nor U4688 (N_4688,In_452,In_2755);
or U4689 (N_4689,In_1826,In_4495);
nand U4690 (N_4690,In_2061,In_151);
nand U4691 (N_4691,In_17,In_50);
nor U4692 (N_4692,In_2753,In_1744);
nand U4693 (N_4693,In_312,In_1637);
xor U4694 (N_4694,In_707,In_2426);
and U4695 (N_4695,In_153,In_1648);
nand U4696 (N_4696,In_2377,In_4034);
xor U4697 (N_4697,In_2946,In_1440);
nand U4698 (N_4698,In_2615,In_1445);
nand U4699 (N_4699,In_1591,In_1799);
xor U4700 (N_4700,In_449,In_168);
and U4701 (N_4701,In_2274,In_2395);
nor U4702 (N_4702,In_3986,In_3910);
nor U4703 (N_4703,In_3167,In_2738);
nand U4704 (N_4704,In_1624,In_762);
and U4705 (N_4705,In_2071,In_4662);
nand U4706 (N_4706,In_2591,In_4455);
nor U4707 (N_4707,In_206,In_17);
and U4708 (N_4708,In_314,In_4616);
or U4709 (N_4709,In_1096,In_3962);
or U4710 (N_4710,In_1838,In_3937);
nand U4711 (N_4711,In_4617,In_2926);
nor U4712 (N_4712,In_237,In_1471);
nor U4713 (N_4713,In_2377,In_4735);
and U4714 (N_4714,In_834,In_2748);
xor U4715 (N_4715,In_2981,In_3262);
and U4716 (N_4716,In_2082,In_3474);
nand U4717 (N_4717,In_2226,In_4875);
and U4718 (N_4718,In_646,In_3152);
and U4719 (N_4719,In_1016,In_4637);
or U4720 (N_4720,In_3930,In_1747);
nor U4721 (N_4721,In_1689,In_499);
nor U4722 (N_4722,In_3782,In_104);
xor U4723 (N_4723,In_1583,In_4129);
or U4724 (N_4724,In_1560,In_4624);
nor U4725 (N_4725,In_4267,In_3224);
nand U4726 (N_4726,In_2604,In_3712);
xor U4727 (N_4727,In_4097,In_1414);
nor U4728 (N_4728,In_4217,In_2646);
or U4729 (N_4729,In_3048,In_407);
and U4730 (N_4730,In_2569,In_343);
and U4731 (N_4731,In_1272,In_1667);
nor U4732 (N_4732,In_979,In_925);
xnor U4733 (N_4733,In_636,In_1050);
xnor U4734 (N_4734,In_2008,In_3905);
nand U4735 (N_4735,In_4925,In_1721);
nand U4736 (N_4736,In_1968,In_4845);
nor U4737 (N_4737,In_724,In_2497);
and U4738 (N_4738,In_2510,In_966);
or U4739 (N_4739,In_4164,In_4986);
xnor U4740 (N_4740,In_1120,In_4516);
and U4741 (N_4741,In_2090,In_2757);
and U4742 (N_4742,In_1984,In_1742);
or U4743 (N_4743,In_962,In_3204);
and U4744 (N_4744,In_744,In_4951);
nor U4745 (N_4745,In_1110,In_4043);
nor U4746 (N_4746,In_427,In_1147);
nor U4747 (N_4747,In_4588,In_4216);
and U4748 (N_4748,In_1318,In_3300);
nor U4749 (N_4749,In_1847,In_609);
nand U4750 (N_4750,In_3932,In_2560);
or U4751 (N_4751,In_4941,In_3569);
and U4752 (N_4752,In_4907,In_1350);
or U4753 (N_4753,In_2471,In_1415);
nor U4754 (N_4754,In_2565,In_1268);
xor U4755 (N_4755,In_761,In_707);
or U4756 (N_4756,In_4334,In_640);
nor U4757 (N_4757,In_4819,In_4016);
xnor U4758 (N_4758,In_332,In_2109);
xor U4759 (N_4759,In_2692,In_437);
or U4760 (N_4760,In_2036,In_2522);
xor U4761 (N_4761,In_1418,In_3007);
xnor U4762 (N_4762,In_4221,In_3899);
and U4763 (N_4763,In_2345,In_27);
xor U4764 (N_4764,In_4512,In_4306);
or U4765 (N_4765,In_58,In_4286);
xor U4766 (N_4766,In_3401,In_4964);
or U4767 (N_4767,In_1196,In_400);
nor U4768 (N_4768,In_4423,In_1739);
xor U4769 (N_4769,In_506,In_3224);
nand U4770 (N_4770,In_3225,In_2793);
nand U4771 (N_4771,In_4317,In_3617);
nand U4772 (N_4772,In_4805,In_1275);
nand U4773 (N_4773,In_2453,In_3347);
nor U4774 (N_4774,In_2796,In_1138);
xnor U4775 (N_4775,In_820,In_600);
or U4776 (N_4776,In_3196,In_4296);
or U4777 (N_4777,In_1649,In_1540);
or U4778 (N_4778,In_3731,In_3398);
nand U4779 (N_4779,In_3205,In_4539);
and U4780 (N_4780,In_4446,In_1088);
or U4781 (N_4781,In_3922,In_3422);
nor U4782 (N_4782,In_815,In_3669);
or U4783 (N_4783,In_3624,In_132);
and U4784 (N_4784,In_745,In_290);
xor U4785 (N_4785,In_3410,In_2404);
nor U4786 (N_4786,In_3213,In_2015);
nor U4787 (N_4787,In_3050,In_356);
nand U4788 (N_4788,In_3900,In_4560);
and U4789 (N_4789,In_2056,In_4317);
nand U4790 (N_4790,In_470,In_2472);
xor U4791 (N_4791,In_805,In_3103);
or U4792 (N_4792,In_819,In_382);
and U4793 (N_4793,In_449,In_4872);
nand U4794 (N_4794,In_4968,In_3765);
xnor U4795 (N_4795,In_1744,In_1921);
or U4796 (N_4796,In_2045,In_79);
or U4797 (N_4797,In_230,In_2367);
nor U4798 (N_4798,In_2766,In_2201);
nand U4799 (N_4799,In_2378,In_1166);
nor U4800 (N_4800,In_4984,In_2295);
nand U4801 (N_4801,In_2066,In_3391);
nand U4802 (N_4802,In_140,In_3317);
nand U4803 (N_4803,In_422,In_2982);
and U4804 (N_4804,In_1494,In_855);
xnor U4805 (N_4805,In_3943,In_3596);
nor U4806 (N_4806,In_4475,In_2371);
nor U4807 (N_4807,In_219,In_431);
xor U4808 (N_4808,In_4670,In_2728);
nor U4809 (N_4809,In_1457,In_3363);
nor U4810 (N_4810,In_1948,In_503);
xnor U4811 (N_4811,In_1679,In_3844);
or U4812 (N_4812,In_2650,In_769);
xor U4813 (N_4813,In_4814,In_2074);
xnor U4814 (N_4814,In_3782,In_508);
and U4815 (N_4815,In_1665,In_2298);
nand U4816 (N_4816,In_579,In_3414);
or U4817 (N_4817,In_4259,In_429);
or U4818 (N_4818,In_743,In_3984);
xor U4819 (N_4819,In_3677,In_2100);
nor U4820 (N_4820,In_2916,In_2382);
or U4821 (N_4821,In_3011,In_478);
xnor U4822 (N_4822,In_2351,In_2572);
nand U4823 (N_4823,In_515,In_4562);
xnor U4824 (N_4824,In_2375,In_2237);
nor U4825 (N_4825,In_4499,In_2011);
or U4826 (N_4826,In_2146,In_3814);
or U4827 (N_4827,In_3797,In_3937);
nand U4828 (N_4828,In_3874,In_2412);
xor U4829 (N_4829,In_370,In_4290);
or U4830 (N_4830,In_3976,In_3601);
nand U4831 (N_4831,In_1222,In_4083);
nand U4832 (N_4832,In_2110,In_4841);
or U4833 (N_4833,In_4130,In_4077);
and U4834 (N_4834,In_2662,In_1614);
xnor U4835 (N_4835,In_4470,In_1287);
xnor U4836 (N_4836,In_1409,In_1122);
xor U4837 (N_4837,In_2516,In_919);
and U4838 (N_4838,In_4664,In_807);
xor U4839 (N_4839,In_218,In_3326);
xor U4840 (N_4840,In_3301,In_105);
xor U4841 (N_4841,In_1423,In_1297);
and U4842 (N_4842,In_4432,In_621);
nand U4843 (N_4843,In_4946,In_1641);
and U4844 (N_4844,In_1091,In_2952);
xor U4845 (N_4845,In_4428,In_1465);
xor U4846 (N_4846,In_2502,In_1734);
nor U4847 (N_4847,In_2409,In_2865);
and U4848 (N_4848,In_1557,In_4851);
xnor U4849 (N_4849,In_1495,In_4051);
xnor U4850 (N_4850,In_3903,In_1951);
and U4851 (N_4851,In_1814,In_2418);
nor U4852 (N_4852,In_980,In_4624);
nor U4853 (N_4853,In_564,In_4382);
nor U4854 (N_4854,In_1218,In_2341);
and U4855 (N_4855,In_2456,In_2589);
xnor U4856 (N_4856,In_3706,In_345);
nor U4857 (N_4857,In_4256,In_1886);
xnor U4858 (N_4858,In_345,In_2128);
xor U4859 (N_4859,In_4516,In_2537);
nand U4860 (N_4860,In_3192,In_4095);
or U4861 (N_4861,In_3086,In_1490);
and U4862 (N_4862,In_3953,In_691);
and U4863 (N_4863,In_4812,In_3084);
and U4864 (N_4864,In_1826,In_2249);
nand U4865 (N_4865,In_1593,In_4995);
or U4866 (N_4866,In_272,In_3434);
nor U4867 (N_4867,In_2514,In_3614);
and U4868 (N_4868,In_4057,In_3707);
xor U4869 (N_4869,In_1036,In_4541);
nor U4870 (N_4870,In_1850,In_2525);
and U4871 (N_4871,In_3456,In_2052);
or U4872 (N_4872,In_687,In_1611);
or U4873 (N_4873,In_4196,In_1984);
or U4874 (N_4874,In_28,In_4723);
and U4875 (N_4875,In_1991,In_2868);
and U4876 (N_4876,In_3681,In_1365);
and U4877 (N_4877,In_1626,In_802);
xor U4878 (N_4878,In_2902,In_1049);
nand U4879 (N_4879,In_4082,In_823);
nand U4880 (N_4880,In_3554,In_118);
nor U4881 (N_4881,In_2446,In_3441);
nand U4882 (N_4882,In_164,In_3311);
nand U4883 (N_4883,In_739,In_3181);
nand U4884 (N_4884,In_2573,In_2065);
or U4885 (N_4885,In_767,In_689);
xnor U4886 (N_4886,In_797,In_4853);
xnor U4887 (N_4887,In_414,In_38);
nand U4888 (N_4888,In_4670,In_4140);
xnor U4889 (N_4889,In_3870,In_596);
and U4890 (N_4890,In_1499,In_4955);
nor U4891 (N_4891,In_3989,In_4000);
nand U4892 (N_4892,In_305,In_4871);
nand U4893 (N_4893,In_2877,In_4608);
and U4894 (N_4894,In_607,In_3328);
xor U4895 (N_4895,In_3420,In_2208);
and U4896 (N_4896,In_4454,In_4139);
nor U4897 (N_4897,In_1089,In_2014);
xor U4898 (N_4898,In_2211,In_4274);
or U4899 (N_4899,In_3547,In_3393);
nand U4900 (N_4900,In_3135,In_335);
or U4901 (N_4901,In_3225,In_3466);
or U4902 (N_4902,In_1425,In_4575);
xor U4903 (N_4903,In_457,In_2528);
or U4904 (N_4904,In_1580,In_1316);
or U4905 (N_4905,In_3411,In_3503);
or U4906 (N_4906,In_3132,In_2916);
nand U4907 (N_4907,In_4389,In_1278);
nor U4908 (N_4908,In_4798,In_4759);
nor U4909 (N_4909,In_4930,In_998);
and U4910 (N_4910,In_3577,In_4921);
or U4911 (N_4911,In_2757,In_4060);
and U4912 (N_4912,In_148,In_472);
or U4913 (N_4913,In_4064,In_3227);
xnor U4914 (N_4914,In_2316,In_3967);
nand U4915 (N_4915,In_1323,In_552);
or U4916 (N_4916,In_2430,In_2146);
and U4917 (N_4917,In_632,In_4038);
nand U4918 (N_4918,In_4810,In_3715);
nand U4919 (N_4919,In_2688,In_162);
or U4920 (N_4920,In_4543,In_3154);
nor U4921 (N_4921,In_196,In_4084);
xnor U4922 (N_4922,In_417,In_4907);
or U4923 (N_4923,In_4247,In_2965);
xnor U4924 (N_4924,In_4741,In_2105);
and U4925 (N_4925,In_4720,In_9);
nor U4926 (N_4926,In_3738,In_4186);
and U4927 (N_4927,In_4546,In_4867);
nand U4928 (N_4928,In_1950,In_658);
and U4929 (N_4929,In_533,In_3783);
xnor U4930 (N_4930,In_2162,In_1445);
nand U4931 (N_4931,In_3829,In_4735);
and U4932 (N_4932,In_3442,In_1346);
and U4933 (N_4933,In_1905,In_2147);
and U4934 (N_4934,In_2047,In_1486);
or U4935 (N_4935,In_2219,In_3725);
or U4936 (N_4936,In_3631,In_1662);
nand U4937 (N_4937,In_1478,In_914);
or U4938 (N_4938,In_1507,In_4004);
nand U4939 (N_4939,In_443,In_2323);
and U4940 (N_4940,In_3998,In_2537);
nor U4941 (N_4941,In_1232,In_495);
xnor U4942 (N_4942,In_1254,In_1903);
and U4943 (N_4943,In_4583,In_2148);
nor U4944 (N_4944,In_947,In_3912);
and U4945 (N_4945,In_4653,In_4816);
or U4946 (N_4946,In_1289,In_1646);
nand U4947 (N_4947,In_4072,In_3550);
nor U4948 (N_4948,In_4849,In_1520);
nand U4949 (N_4949,In_3977,In_3686);
or U4950 (N_4950,In_235,In_2828);
and U4951 (N_4951,In_2878,In_4311);
and U4952 (N_4952,In_685,In_4905);
xnor U4953 (N_4953,In_2492,In_1238);
xnor U4954 (N_4954,In_4744,In_411);
nor U4955 (N_4955,In_4403,In_3272);
xnor U4956 (N_4956,In_379,In_1464);
or U4957 (N_4957,In_4059,In_1019);
xnor U4958 (N_4958,In_3993,In_2049);
nand U4959 (N_4959,In_3706,In_4397);
and U4960 (N_4960,In_4198,In_3563);
nand U4961 (N_4961,In_943,In_231);
or U4962 (N_4962,In_1381,In_2725);
xor U4963 (N_4963,In_4729,In_1092);
xor U4964 (N_4964,In_4564,In_4061);
and U4965 (N_4965,In_2082,In_3198);
nor U4966 (N_4966,In_3972,In_3390);
xnor U4967 (N_4967,In_1271,In_2360);
or U4968 (N_4968,In_1982,In_3795);
xor U4969 (N_4969,In_3824,In_106);
nor U4970 (N_4970,In_999,In_3958);
nor U4971 (N_4971,In_3423,In_2727);
and U4972 (N_4972,In_2464,In_10);
nor U4973 (N_4973,In_4226,In_3894);
and U4974 (N_4974,In_2652,In_3768);
nor U4975 (N_4975,In_4217,In_3662);
nand U4976 (N_4976,In_4966,In_2973);
or U4977 (N_4977,In_1685,In_4919);
and U4978 (N_4978,In_439,In_371);
nor U4979 (N_4979,In_4601,In_593);
xnor U4980 (N_4980,In_16,In_4965);
or U4981 (N_4981,In_2711,In_2760);
and U4982 (N_4982,In_1140,In_692);
or U4983 (N_4983,In_1624,In_289);
xnor U4984 (N_4984,In_3131,In_4448);
or U4985 (N_4985,In_559,In_4578);
nor U4986 (N_4986,In_875,In_1416);
xor U4987 (N_4987,In_14,In_2670);
nor U4988 (N_4988,In_3925,In_2442);
xor U4989 (N_4989,In_4195,In_283);
and U4990 (N_4990,In_3690,In_3947);
nand U4991 (N_4991,In_3831,In_1439);
or U4992 (N_4992,In_4382,In_1275);
nor U4993 (N_4993,In_3447,In_2534);
nand U4994 (N_4994,In_3430,In_1857);
nand U4995 (N_4995,In_413,In_3264);
nor U4996 (N_4996,In_4067,In_1466);
or U4997 (N_4997,In_1082,In_503);
nand U4998 (N_4998,In_2427,In_947);
nor U4999 (N_4999,In_4205,In_3448);
or U5000 (N_5000,In_1732,In_3845);
and U5001 (N_5001,In_1172,In_350);
nor U5002 (N_5002,In_111,In_3085);
and U5003 (N_5003,In_4221,In_3685);
or U5004 (N_5004,In_2212,In_1420);
nor U5005 (N_5005,In_211,In_476);
and U5006 (N_5006,In_3951,In_3121);
or U5007 (N_5007,In_4677,In_2615);
or U5008 (N_5008,In_400,In_1629);
nand U5009 (N_5009,In_1950,In_2588);
xnor U5010 (N_5010,In_2707,In_3708);
or U5011 (N_5011,In_69,In_4261);
nand U5012 (N_5012,In_4713,In_807);
or U5013 (N_5013,In_3621,In_1046);
nand U5014 (N_5014,In_3691,In_4128);
nand U5015 (N_5015,In_2422,In_3330);
nor U5016 (N_5016,In_1105,In_4822);
and U5017 (N_5017,In_4189,In_1207);
or U5018 (N_5018,In_3967,In_303);
nor U5019 (N_5019,In_4001,In_536);
nor U5020 (N_5020,In_4706,In_4464);
nand U5021 (N_5021,In_1567,In_3993);
or U5022 (N_5022,In_885,In_1264);
xor U5023 (N_5023,In_3608,In_4539);
and U5024 (N_5024,In_508,In_2803);
and U5025 (N_5025,In_2506,In_656);
nand U5026 (N_5026,In_2182,In_1793);
nor U5027 (N_5027,In_3931,In_527);
or U5028 (N_5028,In_4273,In_778);
xnor U5029 (N_5029,In_708,In_2851);
and U5030 (N_5030,In_3939,In_4682);
nand U5031 (N_5031,In_1191,In_2846);
and U5032 (N_5032,In_201,In_2291);
nor U5033 (N_5033,In_2999,In_2583);
xor U5034 (N_5034,In_4170,In_4430);
nor U5035 (N_5035,In_3498,In_1253);
nor U5036 (N_5036,In_929,In_2143);
nor U5037 (N_5037,In_1975,In_4750);
xnor U5038 (N_5038,In_1019,In_4614);
and U5039 (N_5039,In_968,In_4261);
and U5040 (N_5040,In_4203,In_4077);
and U5041 (N_5041,In_2884,In_4874);
nor U5042 (N_5042,In_1838,In_3469);
and U5043 (N_5043,In_4805,In_479);
and U5044 (N_5044,In_3987,In_2989);
nor U5045 (N_5045,In_4351,In_4190);
xor U5046 (N_5046,In_1413,In_4210);
xor U5047 (N_5047,In_4115,In_3945);
xnor U5048 (N_5048,In_491,In_284);
and U5049 (N_5049,In_4380,In_3249);
xor U5050 (N_5050,In_4589,In_4221);
and U5051 (N_5051,In_4649,In_2029);
nand U5052 (N_5052,In_2461,In_3075);
and U5053 (N_5053,In_860,In_557);
xor U5054 (N_5054,In_4716,In_1598);
and U5055 (N_5055,In_4887,In_1469);
nand U5056 (N_5056,In_707,In_2587);
xor U5057 (N_5057,In_1791,In_1179);
nor U5058 (N_5058,In_1216,In_3754);
and U5059 (N_5059,In_1043,In_3235);
or U5060 (N_5060,In_3954,In_2035);
and U5061 (N_5061,In_4168,In_2098);
xnor U5062 (N_5062,In_4016,In_4214);
xnor U5063 (N_5063,In_3278,In_1012);
and U5064 (N_5064,In_3802,In_4896);
nor U5065 (N_5065,In_518,In_1782);
nand U5066 (N_5066,In_1373,In_2591);
xnor U5067 (N_5067,In_4272,In_538);
xor U5068 (N_5068,In_1164,In_2429);
nor U5069 (N_5069,In_168,In_3725);
xnor U5070 (N_5070,In_3277,In_1048);
xor U5071 (N_5071,In_3433,In_2675);
xnor U5072 (N_5072,In_817,In_3415);
nand U5073 (N_5073,In_4217,In_3784);
or U5074 (N_5074,In_1534,In_1567);
and U5075 (N_5075,In_3048,In_2504);
or U5076 (N_5076,In_4203,In_980);
and U5077 (N_5077,In_1119,In_1612);
and U5078 (N_5078,In_345,In_3860);
xor U5079 (N_5079,In_805,In_1989);
xor U5080 (N_5080,In_1268,In_829);
and U5081 (N_5081,In_4994,In_4863);
nor U5082 (N_5082,In_4931,In_1735);
xnor U5083 (N_5083,In_606,In_517);
nor U5084 (N_5084,In_3280,In_2289);
nand U5085 (N_5085,In_3591,In_611);
xor U5086 (N_5086,In_3249,In_704);
xnor U5087 (N_5087,In_3596,In_1612);
xor U5088 (N_5088,In_2006,In_1207);
nor U5089 (N_5089,In_890,In_3028);
and U5090 (N_5090,In_1682,In_787);
or U5091 (N_5091,In_2023,In_237);
xor U5092 (N_5092,In_4060,In_910);
xor U5093 (N_5093,In_1892,In_1161);
nand U5094 (N_5094,In_3663,In_1989);
or U5095 (N_5095,In_1485,In_3964);
or U5096 (N_5096,In_3859,In_832);
xnor U5097 (N_5097,In_281,In_2124);
xnor U5098 (N_5098,In_4262,In_4329);
nor U5099 (N_5099,In_2837,In_966);
and U5100 (N_5100,In_4084,In_4191);
or U5101 (N_5101,In_4291,In_4878);
nand U5102 (N_5102,In_363,In_3182);
nor U5103 (N_5103,In_2914,In_4600);
nand U5104 (N_5104,In_2798,In_4419);
or U5105 (N_5105,In_122,In_853);
nor U5106 (N_5106,In_3,In_4175);
and U5107 (N_5107,In_3964,In_2240);
and U5108 (N_5108,In_3600,In_4732);
nand U5109 (N_5109,In_1784,In_2806);
and U5110 (N_5110,In_1187,In_2859);
or U5111 (N_5111,In_861,In_2425);
and U5112 (N_5112,In_2383,In_4702);
nand U5113 (N_5113,In_2761,In_1141);
and U5114 (N_5114,In_3671,In_4498);
nand U5115 (N_5115,In_1028,In_2996);
or U5116 (N_5116,In_3011,In_2074);
or U5117 (N_5117,In_1124,In_610);
and U5118 (N_5118,In_2526,In_3432);
or U5119 (N_5119,In_3963,In_98);
or U5120 (N_5120,In_2259,In_4720);
and U5121 (N_5121,In_4444,In_4631);
xnor U5122 (N_5122,In_848,In_3485);
nor U5123 (N_5123,In_4000,In_4292);
or U5124 (N_5124,In_2279,In_3781);
xor U5125 (N_5125,In_3558,In_864);
and U5126 (N_5126,In_222,In_1019);
nor U5127 (N_5127,In_3802,In_1656);
nand U5128 (N_5128,In_4701,In_205);
or U5129 (N_5129,In_4221,In_1930);
or U5130 (N_5130,In_4298,In_4978);
nand U5131 (N_5131,In_2905,In_3405);
and U5132 (N_5132,In_2217,In_270);
and U5133 (N_5133,In_461,In_1749);
nand U5134 (N_5134,In_3720,In_2708);
and U5135 (N_5135,In_4396,In_4346);
nand U5136 (N_5136,In_1085,In_3127);
xor U5137 (N_5137,In_3206,In_369);
nor U5138 (N_5138,In_3020,In_4609);
xor U5139 (N_5139,In_3303,In_4166);
and U5140 (N_5140,In_50,In_164);
xor U5141 (N_5141,In_324,In_577);
nor U5142 (N_5142,In_2297,In_3060);
nor U5143 (N_5143,In_3224,In_4570);
or U5144 (N_5144,In_3057,In_3278);
or U5145 (N_5145,In_1299,In_1552);
nor U5146 (N_5146,In_1140,In_1123);
nor U5147 (N_5147,In_3228,In_4480);
nand U5148 (N_5148,In_374,In_621);
nand U5149 (N_5149,In_2024,In_4685);
nand U5150 (N_5150,In_3512,In_2416);
nand U5151 (N_5151,In_4448,In_2419);
or U5152 (N_5152,In_3110,In_943);
xor U5153 (N_5153,In_3807,In_802);
nor U5154 (N_5154,In_2960,In_1521);
xor U5155 (N_5155,In_4783,In_4040);
nand U5156 (N_5156,In_4385,In_291);
xor U5157 (N_5157,In_4900,In_1901);
xor U5158 (N_5158,In_1582,In_2746);
xor U5159 (N_5159,In_2911,In_1979);
xnor U5160 (N_5160,In_4869,In_741);
xnor U5161 (N_5161,In_2237,In_2643);
nand U5162 (N_5162,In_889,In_4870);
and U5163 (N_5163,In_3315,In_3746);
nand U5164 (N_5164,In_2445,In_2858);
nand U5165 (N_5165,In_4907,In_1774);
nand U5166 (N_5166,In_3342,In_4495);
nand U5167 (N_5167,In_3236,In_2893);
and U5168 (N_5168,In_4118,In_804);
xor U5169 (N_5169,In_2373,In_2906);
nor U5170 (N_5170,In_809,In_2901);
xnor U5171 (N_5171,In_3136,In_1621);
xnor U5172 (N_5172,In_756,In_1789);
nand U5173 (N_5173,In_3171,In_2794);
and U5174 (N_5174,In_3498,In_458);
nor U5175 (N_5175,In_3877,In_2858);
xor U5176 (N_5176,In_2946,In_1400);
nor U5177 (N_5177,In_4177,In_2614);
nand U5178 (N_5178,In_94,In_1971);
nor U5179 (N_5179,In_4992,In_2320);
xor U5180 (N_5180,In_4738,In_4590);
xnor U5181 (N_5181,In_4623,In_2796);
xor U5182 (N_5182,In_1288,In_3070);
nand U5183 (N_5183,In_3108,In_2272);
or U5184 (N_5184,In_409,In_2255);
nor U5185 (N_5185,In_1790,In_4699);
and U5186 (N_5186,In_4661,In_594);
or U5187 (N_5187,In_1080,In_715);
nor U5188 (N_5188,In_1892,In_233);
nand U5189 (N_5189,In_1025,In_3098);
xor U5190 (N_5190,In_1725,In_1204);
and U5191 (N_5191,In_2682,In_1411);
or U5192 (N_5192,In_3660,In_1462);
or U5193 (N_5193,In_471,In_3132);
or U5194 (N_5194,In_3398,In_92);
or U5195 (N_5195,In_391,In_4281);
and U5196 (N_5196,In_1948,In_1287);
xor U5197 (N_5197,In_87,In_740);
or U5198 (N_5198,In_1348,In_401);
and U5199 (N_5199,In_862,In_1223);
nand U5200 (N_5200,In_2995,In_492);
nand U5201 (N_5201,In_926,In_4009);
nand U5202 (N_5202,In_890,In_144);
and U5203 (N_5203,In_3453,In_4977);
xor U5204 (N_5204,In_3296,In_3003);
and U5205 (N_5205,In_4535,In_3488);
and U5206 (N_5206,In_3942,In_1027);
and U5207 (N_5207,In_392,In_387);
xnor U5208 (N_5208,In_4730,In_4193);
xor U5209 (N_5209,In_1868,In_2988);
nand U5210 (N_5210,In_4745,In_1764);
or U5211 (N_5211,In_4606,In_956);
nand U5212 (N_5212,In_685,In_1995);
and U5213 (N_5213,In_4318,In_3025);
nor U5214 (N_5214,In_1946,In_4185);
or U5215 (N_5215,In_3399,In_4454);
or U5216 (N_5216,In_4996,In_4039);
and U5217 (N_5217,In_3004,In_3839);
nand U5218 (N_5218,In_1052,In_3812);
nand U5219 (N_5219,In_19,In_4029);
nand U5220 (N_5220,In_1524,In_4358);
xor U5221 (N_5221,In_3415,In_2067);
and U5222 (N_5222,In_1755,In_2936);
nand U5223 (N_5223,In_2338,In_3028);
nand U5224 (N_5224,In_2469,In_2379);
xnor U5225 (N_5225,In_3270,In_4519);
and U5226 (N_5226,In_1350,In_2509);
xnor U5227 (N_5227,In_1675,In_1863);
nand U5228 (N_5228,In_3484,In_1138);
xor U5229 (N_5229,In_4227,In_3978);
and U5230 (N_5230,In_2976,In_2271);
nor U5231 (N_5231,In_2480,In_3940);
or U5232 (N_5232,In_126,In_547);
nand U5233 (N_5233,In_1999,In_2503);
and U5234 (N_5234,In_3032,In_3893);
nand U5235 (N_5235,In_3363,In_4750);
nand U5236 (N_5236,In_4657,In_257);
nor U5237 (N_5237,In_3318,In_1350);
and U5238 (N_5238,In_2313,In_3875);
xnor U5239 (N_5239,In_2598,In_986);
nor U5240 (N_5240,In_3591,In_2825);
and U5241 (N_5241,In_3660,In_4817);
xnor U5242 (N_5242,In_4215,In_2257);
xnor U5243 (N_5243,In_2125,In_3411);
or U5244 (N_5244,In_847,In_861);
and U5245 (N_5245,In_704,In_4811);
or U5246 (N_5246,In_2707,In_3845);
and U5247 (N_5247,In_4026,In_3274);
or U5248 (N_5248,In_3470,In_1090);
nand U5249 (N_5249,In_1552,In_4731);
or U5250 (N_5250,In_1157,In_1606);
xor U5251 (N_5251,In_4081,In_1893);
nor U5252 (N_5252,In_3604,In_4335);
and U5253 (N_5253,In_3553,In_4915);
or U5254 (N_5254,In_1852,In_2471);
nor U5255 (N_5255,In_3123,In_317);
xor U5256 (N_5256,In_1436,In_1374);
and U5257 (N_5257,In_3051,In_784);
nand U5258 (N_5258,In_2309,In_3899);
nor U5259 (N_5259,In_89,In_1442);
and U5260 (N_5260,In_3420,In_3280);
or U5261 (N_5261,In_255,In_1326);
xnor U5262 (N_5262,In_4701,In_452);
xnor U5263 (N_5263,In_397,In_3051);
and U5264 (N_5264,In_2301,In_653);
nand U5265 (N_5265,In_1114,In_4965);
nand U5266 (N_5266,In_3568,In_8);
nand U5267 (N_5267,In_1328,In_850);
and U5268 (N_5268,In_2723,In_972);
and U5269 (N_5269,In_4532,In_1953);
nand U5270 (N_5270,In_1250,In_3383);
or U5271 (N_5271,In_970,In_3680);
nor U5272 (N_5272,In_1728,In_4320);
nor U5273 (N_5273,In_2171,In_1940);
and U5274 (N_5274,In_3856,In_4505);
nand U5275 (N_5275,In_3339,In_3046);
nor U5276 (N_5276,In_3542,In_730);
nand U5277 (N_5277,In_943,In_1946);
and U5278 (N_5278,In_2603,In_3507);
nand U5279 (N_5279,In_1300,In_4918);
and U5280 (N_5280,In_1466,In_288);
and U5281 (N_5281,In_1120,In_1341);
xor U5282 (N_5282,In_3117,In_900);
nand U5283 (N_5283,In_316,In_2154);
xor U5284 (N_5284,In_125,In_392);
and U5285 (N_5285,In_4702,In_2759);
and U5286 (N_5286,In_1971,In_4211);
or U5287 (N_5287,In_839,In_4316);
or U5288 (N_5288,In_1202,In_3051);
xnor U5289 (N_5289,In_652,In_4046);
xnor U5290 (N_5290,In_1159,In_951);
xor U5291 (N_5291,In_2818,In_2185);
xnor U5292 (N_5292,In_1584,In_4823);
nor U5293 (N_5293,In_2026,In_1350);
and U5294 (N_5294,In_367,In_4979);
nor U5295 (N_5295,In_3546,In_3565);
nor U5296 (N_5296,In_2163,In_4154);
nor U5297 (N_5297,In_4124,In_1418);
xor U5298 (N_5298,In_1213,In_837);
nand U5299 (N_5299,In_571,In_32);
and U5300 (N_5300,In_4124,In_73);
xor U5301 (N_5301,In_1529,In_1163);
and U5302 (N_5302,In_4124,In_1639);
or U5303 (N_5303,In_4915,In_2550);
and U5304 (N_5304,In_2444,In_1472);
nor U5305 (N_5305,In_2666,In_2417);
or U5306 (N_5306,In_2015,In_4269);
nor U5307 (N_5307,In_4850,In_1263);
nor U5308 (N_5308,In_1359,In_3706);
and U5309 (N_5309,In_2818,In_4959);
or U5310 (N_5310,In_4593,In_1883);
xor U5311 (N_5311,In_1226,In_499);
xor U5312 (N_5312,In_1493,In_1323);
nand U5313 (N_5313,In_2092,In_2691);
nor U5314 (N_5314,In_3363,In_546);
nand U5315 (N_5315,In_3794,In_126);
or U5316 (N_5316,In_322,In_1832);
and U5317 (N_5317,In_4800,In_1536);
nor U5318 (N_5318,In_4263,In_4661);
nor U5319 (N_5319,In_4946,In_543);
nand U5320 (N_5320,In_4874,In_3879);
or U5321 (N_5321,In_4119,In_481);
nor U5322 (N_5322,In_4722,In_591);
and U5323 (N_5323,In_4710,In_4976);
and U5324 (N_5324,In_2446,In_2043);
nand U5325 (N_5325,In_602,In_2837);
nor U5326 (N_5326,In_3042,In_4701);
or U5327 (N_5327,In_63,In_3556);
and U5328 (N_5328,In_465,In_4445);
nor U5329 (N_5329,In_371,In_3719);
and U5330 (N_5330,In_3339,In_2513);
nor U5331 (N_5331,In_4565,In_4634);
nor U5332 (N_5332,In_3127,In_4022);
or U5333 (N_5333,In_3234,In_2426);
nor U5334 (N_5334,In_4304,In_278);
nor U5335 (N_5335,In_2278,In_3127);
and U5336 (N_5336,In_1366,In_3896);
or U5337 (N_5337,In_1107,In_4886);
nand U5338 (N_5338,In_4461,In_1785);
nor U5339 (N_5339,In_2498,In_4150);
nor U5340 (N_5340,In_4679,In_2240);
and U5341 (N_5341,In_3150,In_1885);
xor U5342 (N_5342,In_3048,In_2212);
xor U5343 (N_5343,In_1444,In_2493);
or U5344 (N_5344,In_523,In_4772);
or U5345 (N_5345,In_2235,In_1258);
and U5346 (N_5346,In_2022,In_593);
and U5347 (N_5347,In_1910,In_3767);
nor U5348 (N_5348,In_1040,In_945);
nand U5349 (N_5349,In_2564,In_736);
or U5350 (N_5350,In_890,In_2736);
or U5351 (N_5351,In_1561,In_4081);
nor U5352 (N_5352,In_2145,In_4295);
or U5353 (N_5353,In_3430,In_842);
xnor U5354 (N_5354,In_4457,In_2205);
xnor U5355 (N_5355,In_4593,In_946);
and U5356 (N_5356,In_2853,In_2799);
nand U5357 (N_5357,In_3863,In_3999);
and U5358 (N_5358,In_800,In_1362);
nor U5359 (N_5359,In_3449,In_4965);
nand U5360 (N_5360,In_1329,In_1069);
nand U5361 (N_5361,In_939,In_1735);
nor U5362 (N_5362,In_599,In_971);
or U5363 (N_5363,In_1658,In_1684);
and U5364 (N_5364,In_1035,In_776);
or U5365 (N_5365,In_1814,In_3605);
nand U5366 (N_5366,In_339,In_369);
nor U5367 (N_5367,In_1291,In_3859);
or U5368 (N_5368,In_4626,In_990);
nand U5369 (N_5369,In_403,In_3910);
nand U5370 (N_5370,In_4660,In_1843);
nor U5371 (N_5371,In_2329,In_2648);
and U5372 (N_5372,In_1438,In_2102);
xor U5373 (N_5373,In_2894,In_4206);
or U5374 (N_5374,In_1031,In_3105);
nand U5375 (N_5375,In_2537,In_373);
nor U5376 (N_5376,In_227,In_382);
nand U5377 (N_5377,In_4785,In_1256);
or U5378 (N_5378,In_416,In_2086);
nor U5379 (N_5379,In_3853,In_368);
xor U5380 (N_5380,In_4222,In_4968);
nand U5381 (N_5381,In_2181,In_241);
or U5382 (N_5382,In_1288,In_4192);
and U5383 (N_5383,In_1730,In_4503);
xnor U5384 (N_5384,In_283,In_233);
and U5385 (N_5385,In_3964,In_2668);
or U5386 (N_5386,In_1559,In_1236);
nand U5387 (N_5387,In_3212,In_516);
xnor U5388 (N_5388,In_1376,In_1342);
or U5389 (N_5389,In_1747,In_2413);
nand U5390 (N_5390,In_1459,In_3006);
xnor U5391 (N_5391,In_4248,In_4957);
xor U5392 (N_5392,In_2062,In_3111);
or U5393 (N_5393,In_2643,In_1037);
xnor U5394 (N_5394,In_566,In_2258);
nand U5395 (N_5395,In_3830,In_409);
nand U5396 (N_5396,In_4211,In_4934);
or U5397 (N_5397,In_3481,In_1781);
or U5398 (N_5398,In_635,In_1618);
nor U5399 (N_5399,In_4952,In_3376);
and U5400 (N_5400,In_4979,In_226);
xnor U5401 (N_5401,In_3932,In_3653);
nor U5402 (N_5402,In_28,In_2708);
and U5403 (N_5403,In_2155,In_2208);
xor U5404 (N_5404,In_1347,In_1164);
nor U5405 (N_5405,In_1945,In_4780);
or U5406 (N_5406,In_753,In_1825);
xor U5407 (N_5407,In_4421,In_1751);
and U5408 (N_5408,In_2269,In_2090);
or U5409 (N_5409,In_205,In_4011);
nand U5410 (N_5410,In_4469,In_3998);
xnor U5411 (N_5411,In_4413,In_526);
or U5412 (N_5412,In_4716,In_3928);
and U5413 (N_5413,In_4629,In_4477);
nand U5414 (N_5414,In_806,In_792);
and U5415 (N_5415,In_185,In_4045);
nor U5416 (N_5416,In_195,In_4865);
or U5417 (N_5417,In_90,In_990);
nand U5418 (N_5418,In_3386,In_3034);
and U5419 (N_5419,In_3806,In_2864);
or U5420 (N_5420,In_3832,In_3760);
nor U5421 (N_5421,In_4696,In_3812);
nand U5422 (N_5422,In_1390,In_2267);
nand U5423 (N_5423,In_2688,In_2837);
or U5424 (N_5424,In_2650,In_3323);
or U5425 (N_5425,In_3010,In_1501);
nand U5426 (N_5426,In_4008,In_71);
and U5427 (N_5427,In_3691,In_1415);
nor U5428 (N_5428,In_346,In_2426);
and U5429 (N_5429,In_4701,In_2246);
nand U5430 (N_5430,In_2867,In_3806);
xnor U5431 (N_5431,In_1039,In_2192);
nand U5432 (N_5432,In_1682,In_3746);
xnor U5433 (N_5433,In_1116,In_4906);
xor U5434 (N_5434,In_357,In_3699);
nand U5435 (N_5435,In_200,In_2336);
xnor U5436 (N_5436,In_58,In_2064);
xnor U5437 (N_5437,In_2819,In_2744);
nor U5438 (N_5438,In_695,In_747);
or U5439 (N_5439,In_3663,In_1379);
and U5440 (N_5440,In_3706,In_3855);
nand U5441 (N_5441,In_4707,In_1109);
nor U5442 (N_5442,In_2972,In_1809);
nor U5443 (N_5443,In_2876,In_1281);
xor U5444 (N_5444,In_2615,In_4591);
xor U5445 (N_5445,In_4565,In_3301);
xnor U5446 (N_5446,In_1077,In_4985);
and U5447 (N_5447,In_4257,In_4697);
nand U5448 (N_5448,In_3380,In_327);
xnor U5449 (N_5449,In_689,In_667);
or U5450 (N_5450,In_635,In_3372);
xor U5451 (N_5451,In_1470,In_757);
xnor U5452 (N_5452,In_203,In_1484);
or U5453 (N_5453,In_1549,In_24);
and U5454 (N_5454,In_2659,In_2355);
or U5455 (N_5455,In_1805,In_629);
nor U5456 (N_5456,In_2165,In_1565);
and U5457 (N_5457,In_131,In_4351);
xnor U5458 (N_5458,In_2108,In_2620);
or U5459 (N_5459,In_4240,In_2640);
or U5460 (N_5460,In_4498,In_2155);
nand U5461 (N_5461,In_4658,In_3);
nand U5462 (N_5462,In_2424,In_2629);
or U5463 (N_5463,In_2467,In_4385);
and U5464 (N_5464,In_2136,In_2733);
nand U5465 (N_5465,In_4795,In_1554);
nand U5466 (N_5466,In_1361,In_479);
and U5467 (N_5467,In_1454,In_839);
nor U5468 (N_5468,In_1374,In_3898);
nand U5469 (N_5469,In_4263,In_2058);
xnor U5470 (N_5470,In_2464,In_3655);
nand U5471 (N_5471,In_3405,In_414);
nand U5472 (N_5472,In_632,In_4675);
and U5473 (N_5473,In_2091,In_4847);
and U5474 (N_5474,In_3534,In_3213);
or U5475 (N_5475,In_2548,In_3225);
nor U5476 (N_5476,In_2693,In_4238);
nand U5477 (N_5477,In_195,In_4408);
or U5478 (N_5478,In_4326,In_3292);
nand U5479 (N_5479,In_3053,In_1229);
or U5480 (N_5480,In_4353,In_2504);
and U5481 (N_5481,In_613,In_3814);
nor U5482 (N_5482,In_1076,In_1797);
xor U5483 (N_5483,In_4022,In_3551);
or U5484 (N_5484,In_1947,In_1002);
xor U5485 (N_5485,In_3994,In_4807);
nor U5486 (N_5486,In_1477,In_2344);
nand U5487 (N_5487,In_2439,In_3293);
or U5488 (N_5488,In_1784,In_2353);
nor U5489 (N_5489,In_2938,In_2120);
or U5490 (N_5490,In_4874,In_3957);
and U5491 (N_5491,In_3205,In_769);
xnor U5492 (N_5492,In_1976,In_968);
or U5493 (N_5493,In_4276,In_479);
nand U5494 (N_5494,In_1056,In_2939);
and U5495 (N_5495,In_384,In_1211);
and U5496 (N_5496,In_4637,In_4298);
nand U5497 (N_5497,In_4262,In_4933);
nand U5498 (N_5498,In_902,In_3630);
or U5499 (N_5499,In_727,In_4542);
nor U5500 (N_5500,In_4953,In_649);
or U5501 (N_5501,In_4905,In_3638);
nor U5502 (N_5502,In_4952,In_2829);
or U5503 (N_5503,In_1725,In_2264);
or U5504 (N_5504,In_1308,In_738);
nor U5505 (N_5505,In_3611,In_4331);
xor U5506 (N_5506,In_4865,In_1245);
or U5507 (N_5507,In_765,In_624);
nor U5508 (N_5508,In_722,In_2859);
xor U5509 (N_5509,In_1989,In_1715);
xnor U5510 (N_5510,In_1360,In_2457);
or U5511 (N_5511,In_3367,In_2992);
or U5512 (N_5512,In_606,In_614);
and U5513 (N_5513,In_1744,In_250);
nand U5514 (N_5514,In_2295,In_4753);
nor U5515 (N_5515,In_2381,In_1040);
xor U5516 (N_5516,In_843,In_3744);
nand U5517 (N_5517,In_3024,In_1151);
and U5518 (N_5518,In_4384,In_3508);
nand U5519 (N_5519,In_2486,In_23);
and U5520 (N_5520,In_3860,In_1274);
nor U5521 (N_5521,In_432,In_783);
or U5522 (N_5522,In_1133,In_1532);
or U5523 (N_5523,In_4352,In_2074);
or U5524 (N_5524,In_4953,In_2086);
or U5525 (N_5525,In_1511,In_1555);
or U5526 (N_5526,In_623,In_2244);
nand U5527 (N_5527,In_3928,In_635);
and U5528 (N_5528,In_1284,In_3176);
nand U5529 (N_5529,In_3367,In_403);
and U5530 (N_5530,In_4986,In_3075);
and U5531 (N_5531,In_4671,In_4105);
nor U5532 (N_5532,In_3338,In_416);
nand U5533 (N_5533,In_845,In_3138);
or U5534 (N_5534,In_4957,In_4985);
nor U5535 (N_5535,In_71,In_1035);
or U5536 (N_5536,In_3897,In_2474);
xnor U5537 (N_5537,In_712,In_923);
and U5538 (N_5538,In_1785,In_2486);
xnor U5539 (N_5539,In_2359,In_1374);
xnor U5540 (N_5540,In_3588,In_2830);
nand U5541 (N_5541,In_4402,In_571);
or U5542 (N_5542,In_1809,In_1859);
or U5543 (N_5543,In_2298,In_3519);
or U5544 (N_5544,In_974,In_304);
xnor U5545 (N_5545,In_568,In_3504);
or U5546 (N_5546,In_1737,In_3920);
xnor U5547 (N_5547,In_1698,In_1563);
nand U5548 (N_5548,In_3179,In_1606);
nand U5549 (N_5549,In_4809,In_3907);
and U5550 (N_5550,In_1832,In_1623);
or U5551 (N_5551,In_4279,In_4774);
nand U5552 (N_5552,In_3102,In_4139);
nand U5553 (N_5553,In_3258,In_3532);
or U5554 (N_5554,In_2364,In_3348);
nor U5555 (N_5555,In_1207,In_1822);
nand U5556 (N_5556,In_4797,In_1356);
xnor U5557 (N_5557,In_1370,In_2841);
nand U5558 (N_5558,In_3176,In_2664);
nand U5559 (N_5559,In_3316,In_997);
nor U5560 (N_5560,In_2346,In_3669);
and U5561 (N_5561,In_3994,In_2165);
or U5562 (N_5562,In_3512,In_3258);
or U5563 (N_5563,In_149,In_2432);
and U5564 (N_5564,In_3858,In_2359);
and U5565 (N_5565,In_4927,In_3992);
xnor U5566 (N_5566,In_161,In_4705);
and U5567 (N_5567,In_3558,In_1872);
nand U5568 (N_5568,In_374,In_1993);
or U5569 (N_5569,In_2043,In_2627);
or U5570 (N_5570,In_2895,In_2373);
nand U5571 (N_5571,In_2462,In_3862);
or U5572 (N_5572,In_3405,In_3958);
nor U5573 (N_5573,In_3930,In_504);
nor U5574 (N_5574,In_1228,In_2417);
nand U5575 (N_5575,In_3539,In_4306);
and U5576 (N_5576,In_4955,In_249);
or U5577 (N_5577,In_4816,In_1697);
nor U5578 (N_5578,In_5,In_17);
nor U5579 (N_5579,In_3643,In_2809);
xor U5580 (N_5580,In_2811,In_2102);
nor U5581 (N_5581,In_756,In_3936);
xnor U5582 (N_5582,In_497,In_884);
or U5583 (N_5583,In_4589,In_4519);
and U5584 (N_5584,In_3603,In_133);
and U5585 (N_5585,In_4204,In_229);
nor U5586 (N_5586,In_1192,In_3444);
nand U5587 (N_5587,In_3053,In_669);
or U5588 (N_5588,In_2691,In_3690);
nor U5589 (N_5589,In_1873,In_1571);
and U5590 (N_5590,In_4337,In_458);
or U5591 (N_5591,In_4640,In_4880);
and U5592 (N_5592,In_3371,In_2405);
nand U5593 (N_5593,In_2263,In_3593);
nand U5594 (N_5594,In_4275,In_1992);
or U5595 (N_5595,In_285,In_1288);
nand U5596 (N_5596,In_3875,In_1032);
xor U5597 (N_5597,In_1925,In_4613);
nor U5598 (N_5598,In_958,In_3639);
xnor U5599 (N_5599,In_2271,In_4672);
nor U5600 (N_5600,In_3841,In_3511);
xnor U5601 (N_5601,In_1466,In_2779);
xor U5602 (N_5602,In_2677,In_3045);
and U5603 (N_5603,In_3976,In_461);
and U5604 (N_5604,In_4684,In_2298);
and U5605 (N_5605,In_1874,In_3905);
or U5606 (N_5606,In_4879,In_4234);
or U5607 (N_5607,In_3545,In_189);
nand U5608 (N_5608,In_1447,In_617);
nor U5609 (N_5609,In_3352,In_4039);
nand U5610 (N_5610,In_2399,In_3327);
xnor U5611 (N_5611,In_3231,In_1445);
or U5612 (N_5612,In_4381,In_111);
and U5613 (N_5613,In_2964,In_275);
nand U5614 (N_5614,In_304,In_3654);
xnor U5615 (N_5615,In_4932,In_2203);
or U5616 (N_5616,In_3937,In_4390);
nand U5617 (N_5617,In_2207,In_2096);
or U5618 (N_5618,In_3946,In_2881);
and U5619 (N_5619,In_3127,In_1253);
or U5620 (N_5620,In_285,In_554);
xor U5621 (N_5621,In_1560,In_3067);
nor U5622 (N_5622,In_1668,In_663);
or U5623 (N_5623,In_886,In_3046);
nor U5624 (N_5624,In_4070,In_2462);
xor U5625 (N_5625,In_4877,In_4317);
or U5626 (N_5626,In_1589,In_2163);
and U5627 (N_5627,In_3112,In_1239);
or U5628 (N_5628,In_4306,In_251);
xnor U5629 (N_5629,In_221,In_3591);
or U5630 (N_5630,In_4297,In_1409);
nor U5631 (N_5631,In_1419,In_4023);
xor U5632 (N_5632,In_4674,In_1710);
nand U5633 (N_5633,In_4381,In_1933);
or U5634 (N_5634,In_2629,In_3590);
and U5635 (N_5635,In_2441,In_1978);
and U5636 (N_5636,In_4484,In_3602);
or U5637 (N_5637,In_4051,In_2323);
or U5638 (N_5638,In_2627,In_3963);
nor U5639 (N_5639,In_2629,In_1270);
or U5640 (N_5640,In_2553,In_3242);
and U5641 (N_5641,In_2149,In_4173);
nor U5642 (N_5642,In_2137,In_525);
nand U5643 (N_5643,In_94,In_3838);
xnor U5644 (N_5644,In_571,In_2052);
or U5645 (N_5645,In_1480,In_288);
nor U5646 (N_5646,In_4210,In_1178);
nor U5647 (N_5647,In_1412,In_3828);
nor U5648 (N_5648,In_1929,In_1386);
xor U5649 (N_5649,In_4449,In_995);
nor U5650 (N_5650,In_1925,In_924);
xnor U5651 (N_5651,In_4993,In_3220);
nor U5652 (N_5652,In_2123,In_3087);
nor U5653 (N_5653,In_171,In_4926);
xnor U5654 (N_5654,In_3906,In_3732);
nor U5655 (N_5655,In_151,In_1766);
nand U5656 (N_5656,In_1981,In_520);
nor U5657 (N_5657,In_4730,In_3531);
or U5658 (N_5658,In_4797,In_4811);
and U5659 (N_5659,In_895,In_1058);
xnor U5660 (N_5660,In_589,In_4666);
and U5661 (N_5661,In_3047,In_2009);
nor U5662 (N_5662,In_3809,In_3173);
nor U5663 (N_5663,In_4492,In_3224);
and U5664 (N_5664,In_3294,In_4245);
xnor U5665 (N_5665,In_4512,In_4430);
and U5666 (N_5666,In_1735,In_3329);
nand U5667 (N_5667,In_2522,In_3597);
nand U5668 (N_5668,In_1776,In_328);
or U5669 (N_5669,In_564,In_2484);
nand U5670 (N_5670,In_3558,In_1669);
xnor U5671 (N_5671,In_2292,In_2847);
nand U5672 (N_5672,In_1289,In_3248);
nor U5673 (N_5673,In_3813,In_3958);
and U5674 (N_5674,In_3566,In_3214);
nand U5675 (N_5675,In_4937,In_2384);
xor U5676 (N_5676,In_4180,In_3865);
xor U5677 (N_5677,In_3240,In_2676);
xor U5678 (N_5678,In_659,In_1048);
or U5679 (N_5679,In_2358,In_2942);
xor U5680 (N_5680,In_1901,In_1216);
nor U5681 (N_5681,In_810,In_4602);
nor U5682 (N_5682,In_4186,In_3525);
nor U5683 (N_5683,In_4567,In_1139);
or U5684 (N_5684,In_3627,In_1874);
or U5685 (N_5685,In_4215,In_1123);
nand U5686 (N_5686,In_4383,In_1655);
nand U5687 (N_5687,In_1588,In_4961);
xor U5688 (N_5688,In_1746,In_2862);
or U5689 (N_5689,In_940,In_2702);
or U5690 (N_5690,In_3651,In_4733);
nor U5691 (N_5691,In_3897,In_691);
xnor U5692 (N_5692,In_4001,In_4287);
and U5693 (N_5693,In_2987,In_752);
and U5694 (N_5694,In_2498,In_4147);
nand U5695 (N_5695,In_3149,In_377);
xor U5696 (N_5696,In_2531,In_3337);
nor U5697 (N_5697,In_2748,In_130);
or U5698 (N_5698,In_3767,In_1925);
or U5699 (N_5699,In_4492,In_4951);
and U5700 (N_5700,In_2520,In_2435);
and U5701 (N_5701,In_2013,In_4694);
nor U5702 (N_5702,In_248,In_716);
xnor U5703 (N_5703,In_1342,In_2297);
nand U5704 (N_5704,In_1039,In_4552);
nor U5705 (N_5705,In_785,In_2297);
and U5706 (N_5706,In_118,In_1458);
and U5707 (N_5707,In_2887,In_2814);
nor U5708 (N_5708,In_3087,In_2170);
and U5709 (N_5709,In_4491,In_4070);
xor U5710 (N_5710,In_2659,In_4288);
xor U5711 (N_5711,In_80,In_2482);
nand U5712 (N_5712,In_2419,In_2578);
or U5713 (N_5713,In_3064,In_3025);
and U5714 (N_5714,In_1914,In_1042);
xnor U5715 (N_5715,In_4281,In_282);
nand U5716 (N_5716,In_4857,In_1731);
or U5717 (N_5717,In_3810,In_4105);
nand U5718 (N_5718,In_2710,In_3245);
nand U5719 (N_5719,In_4550,In_4494);
or U5720 (N_5720,In_2128,In_3746);
or U5721 (N_5721,In_430,In_3977);
xor U5722 (N_5722,In_2311,In_2922);
or U5723 (N_5723,In_1938,In_2455);
or U5724 (N_5724,In_1009,In_4105);
nand U5725 (N_5725,In_3973,In_3045);
or U5726 (N_5726,In_31,In_4504);
xnor U5727 (N_5727,In_3546,In_233);
nor U5728 (N_5728,In_3428,In_4809);
and U5729 (N_5729,In_3924,In_31);
nor U5730 (N_5730,In_2029,In_627);
or U5731 (N_5731,In_1077,In_3873);
nor U5732 (N_5732,In_3840,In_2684);
and U5733 (N_5733,In_1651,In_1357);
nor U5734 (N_5734,In_2033,In_2796);
and U5735 (N_5735,In_3188,In_805);
nand U5736 (N_5736,In_2154,In_288);
or U5737 (N_5737,In_2135,In_4459);
and U5738 (N_5738,In_1956,In_3371);
xor U5739 (N_5739,In_2512,In_1665);
or U5740 (N_5740,In_139,In_1731);
or U5741 (N_5741,In_3788,In_1630);
nor U5742 (N_5742,In_1551,In_2621);
xor U5743 (N_5743,In_1830,In_4685);
nand U5744 (N_5744,In_3749,In_2604);
xnor U5745 (N_5745,In_665,In_4672);
or U5746 (N_5746,In_2923,In_3632);
and U5747 (N_5747,In_3499,In_3239);
and U5748 (N_5748,In_1168,In_181);
nor U5749 (N_5749,In_2889,In_2071);
nand U5750 (N_5750,In_2832,In_4715);
and U5751 (N_5751,In_2148,In_4586);
nand U5752 (N_5752,In_1586,In_2084);
and U5753 (N_5753,In_551,In_4896);
and U5754 (N_5754,In_1838,In_360);
and U5755 (N_5755,In_3133,In_752);
nor U5756 (N_5756,In_2928,In_4227);
and U5757 (N_5757,In_1313,In_1211);
nor U5758 (N_5758,In_2535,In_3741);
nand U5759 (N_5759,In_439,In_4882);
nor U5760 (N_5760,In_1888,In_1179);
nand U5761 (N_5761,In_3512,In_3643);
nand U5762 (N_5762,In_1308,In_3713);
nand U5763 (N_5763,In_2362,In_1803);
nor U5764 (N_5764,In_3927,In_3064);
xnor U5765 (N_5765,In_4385,In_4933);
xnor U5766 (N_5766,In_2451,In_3555);
and U5767 (N_5767,In_1601,In_4999);
and U5768 (N_5768,In_817,In_1573);
nand U5769 (N_5769,In_3365,In_3838);
xor U5770 (N_5770,In_3430,In_1962);
and U5771 (N_5771,In_3328,In_196);
nor U5772 (N_5772,In_2944,In_4869);
nand U5773 (N_5773,In_763,In_2342);
xnor U5774 (N_5774,In_3583,In_86);
or U5775 (N_5775,In_2342,In_1318);
xnor U5776 (N_5776,In_4022,In_4174);
xor U5777 (N_5777,In_3278,In_3158);
or U5778 (N_5778,In_4840,In_4542);
nor U5779 (N_5779,In_3981,In_3380);
or U5780 (N_5780,In_2891,In_2980);
xnor U5781 (N_5781,In_3829,In_3678);
nand U5782 (N_5782,In_4566,In_4077);
and U5783 (N_5783,In_1343,In_962);
nand U5784 (N_5784,In_1749,In_824);
nand U5785 (N_5785,In_3117,In_4285);
or U5786 (N_5786,In_4724,In_2181);
xor U5787 (N_5787,In_2275,In_3468);
nor U5788 (N_5788,In_2732,In_586);
nor U5789 (N_5789,In_1926,In_4444);
or U5790 (N_5790,In_3200,In_2177);
xnor U5791 (N_5791,In_2299,In_1944);
xnor U5792 (N_5792,In_3186,In_1531);
nand U5793 (N_5793,In_2744,In_1927);
nand U5794 (N_5794,In_2919,In_3403);
nor U5795 (N_5795,In_902,In_4841);
or U5796 (N_5796,In_2255,In_3930);
nor U5797 (N_5797,In_4559,In_2606);
and U5798 (N_5798,In_3050,In_4052);
nand U5799 (N_5799,In_861,In_1799);
or U5800 (N_5800,In_500,In_875);
nand U5801 (N_5801,In_1919,In_1041);
and U5802 (N_5802,In_1065,In_4617);
nand U5803 (N_5803,In_594,In_2151);
nand U5804 (N_5804,In_937,In_4855);
nor U5805 (N_5805,In_2435,In_4397);
or U5806 (N_5806,In_4509,In_4738);
xor U5807 (N_5807,In_3812,In_1456);
and U5808 (N_5808,In_2833,In_1565);
nand U5809 (N_5809,In_3190,In_4380);
nand U5810 (N_5810,In_1455,In_1625);
nand U5811 (N_5811,In_4429,In_3643);
and U5812 (N_5812,In_1188,In_1073);
nand U5813 (N_5813,In_1291,In_1227);
nor U5814 (N_5814,In_80,In_3650);
nand U5815 (N_5815,In_1291,In_1035);
or U5816 (N_5816,In_4593,In_1937);
or U5817 (N_5817,In_1993,In_3922);
and U5818 (N_5818,In_658,In_2250);
and U5819 (N_5819,In_1951,In_583);
or U5820 (N_5820,In_39,In_112);
or U5821 (N_5821,In_3311,In_3000);
or U5822 (N_5822,In_1529,In_4970);
xor U5823 (N_5823,In_856,In_2121);
nor U5824 (N_5824,In_2514,In_2475);
xnor U5825 (N_5825,In_350,In_2003);
nor U5826 (N_5826,In_3665,In_2455);
nand U5827 (N_5827,In_3516,In_1241);
or U5828 (N_5828,In_4886,In_3072);
or U5829 (N_5829,In_4221,In_26);
xor U5830 (N_5830,In_393,In_1265);
xnor U5831 (N_5831,In_2773,In_24);
xor U5832 (N_5832,In_2203,In_3615);
or U5833 (N_5833,In_2915,In_4939);
and U5834 (N_5834,In_2857,In_255);
and U5835 (N_5835,In_2465,In_3383);
and U5836 (N_5836,In_2705,In_4359);
or U5837 (N_5837,In_2642,In_4463);
or U5838 (N_5838,In_4434,In_4830);
or U5839 (N_5839,In_3340,In_2756);
nor U5840 (N_5840,In_4064,In_4529);
nor U5841 (N_5841,In_386,In_887);
and U5842 (N_5842,In_3994,In_4057);
nand U5843 (N_5843,In_2850,In_196);
nand U5844 (N_5844,In_4630,In_1330);
xor U5845 (N_5845,In_1067,In_3378);
nor U5846 (N_5846,In_2424,In_2037);
nor U5847 (N_5847,In_1194,In_1818);
and U5848 (N_5848,In_4126,In_4216);
xnor U5849 (N_5849,In_2374,In_2535);
and U5850 (N_5850,In_4897,In_57);
nand U5851 (N_5851,In_4533,In_4534);
and U5852 (N_5852,In_1960,In_4806);
xnor U5853 (N_5853,In_2300,In_4473);
nand U5854 (N_5854,In_2896,In_3135);
nand U5855 (N_5855,In_1244,In_1304);
xor U5856 (N_5856,In_4327,In_585);
and U5857 (N_5857,In_105,In_3734);
xnor U5858 (N_5858,In_4464,In_1765);
nor U5859 (N_5859,In_4914,In_2025);
and U5860 (N_5860,In_1276,In_522);
or U5861 (N_5861,In_2054,In_4255);
nand U5862 (N_5862,In_429,In_2675);
or U5863 (N_5863,In_1937,In_2597);
or U5864 (N_5864,In_1509,In_145);
nand U5865 (N_5865,In_1572,In_2450);
or U5866 (N_5866,In_208,In_321);
or U5867 (N_5867,In_1843,In_3555);
and U5868 (N_5868,In_4034,In_3151);
xnor U5869 (N_5869,In_1837,In_1937);
xor U5870 (N_5870,In_4965,In_1348);
and U5871 (N_5871,In_2595,In_3528);
nor U5872 (N_5872,In_2046,In_3557);
and U5873 (N_5873,In_1698,In_3394);
xor U5874 (N_5874,In_2522,In_3788);
xor U5875 (N_5875,In_4791,In_4109);
and U5876 (N_5876,In_3570,In_1357);
and U5877 (N_5877,In_1272,In_1906);
nor U5878 (N_5878,In_1212,In_3049);
xnor U5879 (N_5879,In_1260,In_35);
or U5880 (N_5880,In_4000,In_2068);
nor U5881 (N_5881,In_4548,In_3607);
xnor U5882 (N_5882,In_2998,In_623);
or U5883 (N_5883,In_1961,In_4574);
and U5884 (N_5884,In_4709,In_2941);
xor U5885 (N_5885,In_2124,In_2567);
nand U5886 (N_5886,In_3779,In_3996);
or U5887 (N_5887,In_317,In_1565);
or U5888 (N_5888,In_661,In_1107);
and U5889 (N_5889,In_1524,In_1807);
nand U5890 (N_5890,In_4445,In_3015);
or U5891 (N_5891,In_2189,In_3628);
nor U5892 (N_5892,In_4478,In_4733);
nor U5893 (N_5893,In_4589,In_3959);
xnor U5894 (N_5894,In_710,In_4452);
or U5895 (N_5895,In_3350,In_3174);
or U5896 (N_5896,In_875,In_2544);
nand U5897 (N_5897,In_3577,In_1253);
nand U5898 (N_5898,In_2059,In_4091);
and U5899 (N_5899,In_1663,In_4264);
xor U5900 (N_5900,In_3648,In_1257);
nand U5901 (N_5901,In_4479,In_4156);
nor U5902 (N_5902,In_1046,In_4510);
nor U5903 (N_5903,In_244,In_3394);
or U5904 (N_5904,In_1616,In_4355);
nor U5905 (N_5905,In_1703,In_1785);
or U5906 (N_5906,In_1769,In_359);
or U5907 (N_5907,In_318,In_795);
nand U5908 (N_5908,In_2692,In_683);
xor U5909 (N_5909,In_2452,In_1619);
xor U5910 (N_5910,In_4130,In_2014);
or U5911 (N_5911,In_3862,In_3670);
or U5912 (N_5912,In_2023,In_3535);
nand U5913 (N_5913,In_885,In_554);
nor U5914 (N_5914,In_322,In_3102);
nand U5915 (N_5915,In_1714,In_4016);
nand U5916 (N_5916,In_1430,In_4073);
nor U5917 (N_5917,In_661,In_3010);
xnor U5918 (N_5918,In_4822,In_4213);
nor U5919 (N_5919,In_4889,In_747);
or U5920 (N_5920,In_3845,In_2794);
nor U5921 (N_5921,In_905,In_467);
nand U5922 (N_5922,In_1873,In_2941);
nor U5923 (N_5923,In_127,In_83);
nor U5924 (N_5924,In_3004,In_1759);
nor U5925 (N_5925,In_4217,In_427);
nand U5926 (N_5926,In_766,In_2456);
or U5927 (N_5927,In_3415,In_2706);
nor U5928 (N_5928,In_3597,In_3061);
nor U5929 (N_5929,In_1043,In_1439);
xor U5930 (N_5930,In_4147,In_1953);
nand U5931 (N_5931,In_1692,In_1862);
nor U5932 (N_5932,In_3281,In_211);
or U5933 (N_5933,In_1061,In_1466);
and U5934 (N_5934,In_2899,In_4896);
xnor U5935 (N_5935,In_2372,In_3379);
or U5936 (N_5936,In_4654,In_4253);
and U5937 (N_5937,In_3148,In_4560);
xnor U5938 (N_5938,In_4441,In_4709);
xor U5939 (N_5939,In_899,In_416);
and U5940 (N_5940,In_482,In_4583);
nand U5941 (N_5941,In_1565,In_3750);
and U5942 (N_5942,In_3747,In_1551);
or U5943 (N_5943,In_341,In_1431);
and U5944 (N_5944,In_4059,In_2007);
or U5945 (N_5945,In_361,In_1736);
xnor U5946 (N_5946,In_3053,In_4903);
or U5947 (N_5947,In_1325,In_3682);
nor U5948 (N_5948,In_4331,In_284);
nand U5949 (N_5949,In_4819,In_3288);
xnor U5950 (N_5950,In_3612,In_437);
or U5951 (N_5951,In_2319,In_3511);
nand U5952 (N_5952,In_213,In_1842);
or U5953 (N_5953,In_4101,In_1190);
nand U5954 (N_5954,In_897,In_1956);
or U5955 (N_5955,In_4839,In_2068);
xnor U5956 (N_5956,In_3169,In_4440);
nor U5957 (N_5957,In_4340,In_4623);
xnor U5958 (N_5958,In_3613,In_1122);
or U5959 (N_5959,In_2370,In_3749);
nand U5960 (N_5960,In_1667,In_204);
and U5961 (N_5961,In_4069,In_3704);
nor U5962 (N_5962,In_690,In_1940);
xnor U5963 (N_5963,In_2526,In_3613);
or U5964 (N_5964,In_4249,In_815);
nand U5965 (N_5965,In_966,In_2493);
and U5966 (N_5966,In_524,In_597);
xnor U5967 (N_5967,In_2930,In_3053);
or U5968 (N_5968,In_3099,In_973);
xor U5969 (N_5969,In_301,In_3211);
xnor U5970 (N_5970,In_1976,In_3306);
or U5971 (N_5971,In_1656,In_4776);
or U5972 (N_5972,In_4190,In_2822);
nand U5973 (N_5973,In_4891,In_1883);
and U5974 (N_5974,In_1515,In_460);
nand U5975 (N_5975,In_4520,In_2118);
nor U5976 (N_5976,In_136,In_1712);
or U5977 (N_5977,In_2627,In_418);
nor U5978 (N_5978,In_419,In_4686);
xor U5979 (N_5979,In_4531,In_444);
nand U5980 (N_5980,In_1866,In_249);
xnor U5981 (N_5981,In_1330,In_1602);
xnor U5982 (N_5982,In_4452,In_3515);
nor U5983 (N_5983,In_2969,In_489);
nor U5984 (N_5984,In_1140,In_1126);
and U5985 (N_5985,In_982,In_4304);
and U5986 (N_5986,In_3969,In_71);
xnor U5987 (N_5987,In_4311,In_667);
or U5988 (N_5988,In_4682,In_574);
xor U5989 (N_5989,In_2962,In_951);
nand U5990 (N_5990,In_1418,In_4912);
or U5991 (N_5991,In_2820,In_3740);
or U5992 (N_5992,In_1532,In_3702);
or U5993 (N_5993,In_272,In_4421);
or U5994 (N_5994,In_4409,In_4905);
nand U5995 (N_5995,In_918,In_3262);
nand U5996 (N_5996,In_2732,In_1660);
or U5997 (N_5997,In_2003,In_1874);
or U5998 (N_5998,In_3263,In_4437);
or U5999 (N_5999,In_3577,In_3184);
nand U6000 (N_6000,In_4606,In_1310);
nand U6001 (N_6001,In_1042,In_4668);
and U6002 (N_6002,In_2828,In_3008);
or U6003 (N_6003,In_4753,In_482);
nor U6004 (N_6004,In_630,In_2165);
and U6005 (N_6005,In_3863,In_1562);
or U6006 (N_6006,In_2931,In_2497);
or U6007 (N_6007,In_1331,In_2554);
xor U6008 (N_6008,In_984,In_1388);
nand U6009 (N_6009,In_4940,In_4812);
or U6010 (N_6010,In_4098,In_2769);
nor U6011 (N_6011,In_3552,In_486);
or U6012 (N_6012,In_3417,In_1398);
xor U6013 (N_6013,In_2299,In_3419);
nor U6014 (N_6014,In_2712,In_3616);
and U6015 (N_6015,In_3341,In_4748);
or U6016 (N_6016,In_4314,In_819);
or U6017 (N_6017,In_969,In_4853);
or U6018 (N_6018,In_235,In_2651);
nand U6019 (N_6019,In_1381,In_1246);
xor U6020 (N_6020,In_618,In_1513);
or U6021 (N_6021,In_871,In_4134);
nor U6022 (N_6022,In_540,In_4651);
nor U6023 (N_6023,In_4130,In_480);
or U6024 (N_6024,In_4771,In_4675);
xnor U6025 (N_6025,In_4514,In_2672);
or U6026 (N_6026,In_3643,In_435);
nor U6027 (N_6027,In_1821,In_1792);
nor U6028 (N_6028,In_2995,In_2952);
or U6029 (N_6029,In_2567,In_1149);
nor U6030 (N_6030,In_3027,In_4240);
xor U6031 (N_6031,In_2302,In_1049);
or U6032 (N_6032,In_659,In_1716);
and U6033 (N_6033,In_1481,In_2388);
nor U6034 (N_6034,In_544,In_2526);
nand U6035 (N_6035,In_3591,In_3964);
and U6036 (N_6036,In_1789,In_507);
nor U6037 (N_6037,In_815,In_2488);
nand U6038 (N_6038,In_4880,In_1269);
xnor U6039 (N_6039,In_1326,In_3397);
nor U6040 (N_6040,In_3217,In_4169);
and U6041 (N_6041,In_2458,In_128);
and U6042 (N_6042,In_904,In_4567);
or U6043 (N_6043,In_2065,In_3454);
nand U6044 (N_6044,In_85,In_1941);
nand U6045 (N_6045,In_4747,In_691);
or U6046 (N_6046,In_1706,In_1059);
nor U6047 (N_6047,In_3435,In_1352);
xnor U6048 (N_6048,In_1042,In_2434);
or U6049 (N_6049,In_2772,In_3917);
nand U6050 (N_6050,In_2414,In_2741);
nand U6051 (N_6051,In_4827,In_3152);
and U6052 (N_6052,In_3939,In_4101);
or U6053 (N_6053,In_4831,In_1503);
xnor U6054 (N_6054,In_4977,In_2801);
and U6055 (N_6055,In_3933,In_1037);
nand U6056 (N_6056,In_3716,In_2939);
xor U6057 (N_6057,In_1213,In_3159);
xor U6058 (N_6058,In_4873,In_2952);
nor U6059 (N_6059,In_543,In_4083);
nor U6060 (N_6060,In_2606,In_2817);
nand U6061 (N_6061,In_1323,In_3265);
nand U6062 (N_6062,In_397,In_1639);
nor U6063 (N_6063,In_472,In_2425);
nor U6064 (N_6064,In_2342,In_4063);
and U6065 (N_6065,In_4460,In_301);
nor U6066 (N_6066,In_2319,In_984);
nand U6067 (N_6067,In_1426,In_3385);
and U6068 (N_6068,In_3565,In_3681);
xnor U6069 (N_6069,In_2494,In_2866);
and U6070 (N_6070,In_3270,In_4117);
and U6071 (N_6071,In_1125,In_4278);
nand U6072 (N_6072,In_4144,In_4659);
xnor U6073 (N_6073,In_3721,In_762);
xnor U6074 (N_6074,In_215,In_3225);
and U6075 (N_6075,In_1230,In_4511);
xor U6076 (N_6076,In_2589,In_2052);
nand U6077 (N_6077,In_4359,In_4684);
nor U6078 (N_6078,In_2961,In_3867);
xnor U6079 (N_6079,In_904,In_4513);
xnor U6080 (N_6080,In_4574,In_4941);
and U6081 (N_6081,In_604,In_1652);
nand U6082 (N_6082,In_3067,In_553);
nand U6083 (N_6083,In_2568,In_4688);
and U6084 (N_6084,In_522,In_590);
and U6085 (N_6085,In_934,In_1602);
and U6086 (N_6086,In_302,In_4946);
nand U6087 (N_6087,In_288,In_3520);
xnor U6088 (N_6088,In_4835,In_1917);
nand U6089 (N_6089,In_3162,In_4282);
xor U6090 (N_6090,In_1775,In_2809);
or U6091 (N_6091,In_3231,In_1390);
nand U6092 (N_6092,In_4065,In_3728);
nand U6093 (N_6093,In_1835,In_3226);
nor U6094 (N_6094,In_2778,In_1225);
nor U6095 (N_6095,In_1578,In_3907);
nor U6096 (N_6096,In_996,In_2535);
and U6097 (N_6097,In_490,In_1656);
or U6098 (N_6098,In_2282,In_4208);
nor U6099 (N_6099,In_1753,In_188);
xnor U6100 (N_6100,In_1798,In_1364);
and U6101 (N_6101,In_4644,In_149);
and U6102 (N_6102,In_3508,In_845);
nand U6103 (N_6103,In_3887,In_1923);
or U6104 (N_6104,In_1216,In_1906);
and U6105 (N_6105,In_936,In_3419);
nand U6106 (N_6106,In_2077,In_1324);
nand U6107 (N_6107,In_3805,In_4644);
nand U6108 (N_6108,In_632,In_2346);
xor U6109 (N_6109,In_1235,In_112);
nor U6110 (N_6110,In_4676,In_1040);
xnor U6111 (N_6111,In_2389,In_821);
or U6112 (N_6112,In_3753,In_1519);
or U6113 (N_6113,In_1916,In_2134);
and U6114 (N_6114,In_892,In_4891);
nor U6115 (N_6115,In_2765,In_4074);
nand U6116 (N_6116,In_4199,In_2968);
nand U6117 (N_6117,In_1985,In_787);
nand U6118 (N_6118,In_4980,In_20);
and U6119 (N_6119,In_750,In_4195);
or U6120 (N_6120,In_4377,In_3842);
or U6121 (N_6121,In_151,In_3762);
xnor U6122 (N_6122,In_3677,In_638);
and U6123 (N_6123,In_3389,In_1038);
or U6124 (N_6124,In_3395,In_4087);
or U6125 (N_6125,In_3474,In_129);
and U6126 (N_6126,In_2899,In_2250);
nand U6127 (N_6127,In_2509,In_4822);
and U6128 (N_6128,In_1869,In_2732);
nor U6129 (N_6129,In_4357,In_1449);
nor U6130 (N_6130,In_651,In_435);
nor U6131 (N_6131,In_45,In_2552);
and U6132 (N_6132,In_1901,In_1820);
and U6133 (N_6133,In_3910,In_4747);
xor U6134 (N_6134,In_3181,In_1249);
nand U6135 (N_6135,In_4149,In_3628);
nor U6136 (N_6136,In_3404,In_159);
xnor U6137 (N_6137,In_3450,In_3502);
or U6138 (N_6138,In_3961,In_3164);
and U6139 (N_6139,In_3543,In_4132);
nor U6140 (N_6140,In_860,In_2659);
nand U6141 (N_6141,In_583,In_1387);
and U6142 (N_6142,In_1643,In_1261);
xnor U6143 (N_6143,In_2716,In_678);
or U6144 (N_6144,In_2653,In_1953);
and U6145 (N_6145,In_2785,In_2069);
xor U6146 (N_6146,In_4911,In_3522);
xnor U6147 (N_6147,In_3436,In_4671);
and U6148 (N_6148,In_2337,In_1474);
nor U6149 (N_6149,In_3563,In_471);
xnor U6150 (N_6150,In_1334,In_898);
or U6151 (N_6151,In_520,In_4685);
and U6152 (N_6152,In_3640,In_1469);
nor U6153 (N_6153,In_8,In_4545);
nand U6154 (N_6154,In_4566,In_1651);
or U6155 (N_6155,In_1514,In_4593);
nand U6156 (N_6156,In_3632,In_2801);
nand U6157 (N_6157,In_2741,In_3537);
nor U6158 (N_6158,In_2056,In_902);
nand U6159 (N_6159,In_350,In_2966);
or U6160 (N_6160,In_3142,In_3750);
and U6161 (N_6161,In_3528,In_3502);
and U6162 (N_6162,In_3084,In_416);
nand U6163 (N_6163,In_2556,In_4948);
nand U6164 (N_6164,In_2569,In_2189);
or U6165 (N_6165,In_2677,In_819);
and U6166 (N_6166,In_1485,In_1183);
nor U6167 (N_6167,In_1057,In_1270);
and U6168 (N_6168,In_703,In_1004);
xnor U6169 (N_6169,In_1590,In_3051);
xor U6170 (N_6170,In_1303,In_4988);
or U6171 (N_6171,In_1327,In_3849);
nor U6172 (N_6172,In_3895,In_1586);
or U6173 (N_6173,In_3055,In_4703);
or U6174 (N_6174,In_3119,In_3056);
or U6175 (N_6175,In_4881,In_1979);
or U6176 (N_6176,In_1255,In_947);
and U6177 (N_6177,In_4318,In_3813);
nor U6178 (N_6178,In_4095,In_4811);
and U6179 (N_6179,In_4464,In_3467);
or U6180 (N_6180,In_4863,In_109);
or U6181 (N_6181,In_958,In_760);
nor U6182 (N_6182,In_4451,In_262);
nand U6183 (N_6183,In_2688,In_291);
and U6184 (N_6184,In_2103,In_2594);
nand U6185 (N_6185,In_2070,In_2768);
xor U6186 (N_6186,In_3770,In_2770);
or U6187 (N_6187,In_3479,In_4999);
xor U6188 (N_6188,In_1488,In_4081);
nand U6189 (N_6189,In_1420,In_1277);
or U6190 (N_6190,In_4431,In_442);
and U6191 (N_6191,In_1929,In_1054);
xor U6192 (N_6192,In_1991,In_1038);
or U6193 (N_6193,In_3572,In_479);
nand U6194 (N_6194,In_4934,In_2041);
xor U6195 (N_6195,In_2937,In_229);
xnor U6196 (N_6196,In_1358,In_3832);
or U6197 (N_6197,In_4365,In_1076);
nor U6198 (N_6198,In_396,In_3339);
nor U6199 (N_6199,In_2363,In_3173);
xnor U6200 (N_6200,In_4260,In_1722);
nor U6201 (N_6201,In_4217,In_3889);
and U6202 (N_6202,In_3196,In_3412);
nor U6203 (N_6203,In_4204,In_475);
xor U6204 (N_6204,In_4748,In_3960);
nand U6205 (N_6205,In_3512,In_2148);
and U6206 (N_6206,In_441,In_288);
and U6207 (N_6207,In_2577,In_1796);
and U6208 (N_6208,In_1927,In_4640);
nor U6209 (N_6209,In_3832,In_449);
nor U6210 (N_6210,In_2823,In_4808);
xor U6211 (N_6211,In_4749,In_425);
or U6212 (N_6212,In_85,In_1547);
xor U6213 (N_6213,In_4987,In_2409);
nand U6214 (N_6214,In_1677,In_1581);
nor U6215 (N_6215,In_973,In_2108);
nor U6216 (N_6216,In_2498,In_1963);
nor U6217 (N_6217,In_879,In_2833);
nand U6218 (N_6218,In_2546,In_3661);
nand U6219 (N_6219,In_2618,In_2716);
nor U6220 (N_6220,In_2038,In_91);
nand U6221 (N_6221,In_2833,In_1860);
or U6222 (N_6222,In_1942,In_3201);
and U6223 (N_6223,In_898,In_4386);
nor U6224 (N_6224,In_4538,In_3066);
nand U6225 (N_6225,In_3674,In_2988);
or U6226 (N_6226,In_2958,In_2337);
xor U6227 (N_6227,In_1605,In_1619);
nand U6228 (N_6228,In_2158,In_1712);
xor U6229 (N_6229,In_327,In_4673);
nor U6230 (N_6230,In_3618,In_2471);
nor U6231 (N_6231,In_3209,In_839);
and U6232 (N_6232,In_2479,In_1957);
xnor U6233 (N_6233,In_3175,In_886);
nor U6234 (N_6234,In_830,In_2508);
nor U6235 (N_6235,In_798,In_4221);
nand U6236 (N_6236,In_923,In_3280);
nor U6237 (N_6237,In_4655,In_2129);
and U6238 (N_6238,In_3497,In_198);
xnor U6239 (N_6239,In_3622,In_3938);
nand U6240 (N_6240,In_82,In_1572);
and U6241 (N_6241,In_1478,In_2278);
xor U6242 (N_6242,In_4952,In_2397);
xor U6243 (N_6243,In_1510,In_4837);
nand U6244 (N_6244,In_2869,In_1380);
and U6245 (N_6245,In_744,In_4482);
nand U6246 (N_6246,In_1285,In_889);
and U6247 (N_6247,In_4422,In_1814);
nor U6248 (N_6248,In_4431,In_1202);
or U6249 (N_6249,In_3732,In_1070);
nand U6250 (N_6250,In_4118,In_3114);
and U6251 (N_6251,In_1261,In_3653);
nor U6252 (N_6252,In_4442,In_3778);
or U6253 (N_6253,In_4473,In_1998);
xor U6254 (N_6254,In_547,In_1159);
xor U6255 (N_6255,In_2947,In_2501);
and U6256 (N_6256,In_2785,In_3459);
xor U6257 (N_6257,In_3146,In_4248);
or U6258 (N_6258,In_4895,In_1071);
and U6259 (N_6259,In_503,In_4667);
xor U6260 (N_6260,In_1477,In_2429);
xnor U6261 (N_6261,In_2553,In_88);
nand U6262 (N_6262,In_2439,In_2298);
and U6263 (N_6263,In_3944,In_31);
nor U6264 (N_6264,In_4284,In_905);
and U6265 (N_6265,In_4717,In_3654);
nand U6266 (N_6266,In_2851,In_4922);
xnor U6267 (N_6267,In_157,In_500);
or U6268 (N_6268,In_4348,In_1923);
and U6269 (N_6269,In_446,In_2274);
and U6270 (N_6270,In_3009,In_2011);
and U6271 (N_6271,In_2438,In_913);
or U6272 (N_6272,In_3547,In_3850);
nor U6273 (N_6273,In_4398,In_717);
xnor U6274 (N_6274,In_2661,In_2857);
xnor U6275 (N_6275,In_1655,In_1844);
nand U6276 (N_6276,In_580,In_4185);
xnor U6277 (N_6277,In_750,In_4024);
xnor U6278 (N_6278,In_257,In_3960);
nand U6279 (N_6279,In_3378,In_3098);
and U6280 (N_6280,In_2454,In_4520);
or U6281 (N_6281,In_1824,In_1248);
and U6282 (N_6282,In_285,In_4527);
xor U6283 (N_6283,In_200,In_170);
and U6284 (N_6284,In_656,In_4610);
xnor U6285 (N_6285,In_2069,In_4698);
or U6286 (N_6286,In_2894,In_3816);
nor U6287 (N_6287,In_3598,In_3312);
xnor U6288 (N_6288,In_3369,In_3654);
or U6289 (N_6289,In_1114,In_4084);
nor U6290 (N_6290,In_2520,In_4269);
xor U6291 (N_6291,In_731,In_209);
nand U6292 (N_6292,In_4373,In_2821);
and U6293 (N_6293,In_2915,In_4899);
and U6294 (N_6294,In_3097,In_4516);
nand U6295 (N_6295,In_675,In_3465);
nand U6296 (N_6296,In_1740,In_563);
xor U6297 (N_6297,In_1763,In_878);
and U6298 (N_6298,In_2819,In_1003);
nor U6299 (N_6299,In_627,In_1603);
xnor U6300 (N_6300,In_2777,In_718);
or U6301 (N_6301,In_2122,In_4283);
nor U6302 (N_6302,In_4989,In_1525);
or U6303 (N_6303,In_4389,In_4916);
nand U6304 (N_6304,In_3983,In_214);
or U6305 (N_6305,In_1052,In_2741);
xor U6306 (N_6306,In_4635,In_4526);
nor U6307 (N_6307,In_3010,In_1637);
nand U6308 (N_6308,In_2608,In_3386);
xor U6309 (N_6309,In_4771,In_729);
xnor U6310 (N_6310,In_2859,In_2210);
xnor U6311 (N_6311,In_4973,In_2882);
and U6312 (N_6312,In_2815,In_4975);
nand U6313 (N_6313,In_4533,In_2084);
nor U6314 (N_6314,In_4246,In_719);
and U6315 (N_6315,In_1874,In_4846);
xnor U6316 (N_6316,In_644,In_4079);
xnor U6317 (N_6317,In_4832,In_3687);
or U6318 (N_6318,In_2777,In_2265);
and U6319 (N_6319,In_4772,In_3822);
nor U6320 (N_6320,In_1374,In_2916);
nand U6321 (N_6321,In_2746,In_3399);
or U6322 (N_6322,In_3242,In_456);
nor U6323 (N_6323,In_1966,In_909);
and U6324 (N_6324,In_2300,In_3781);
nand U6325 (N_6325,In_1235,In_76);
xnor U6326 (N_6326,In_1022,In_2620);
nor U6327 (N_6327,In_4412,In_393);
or U6328 (N_6328,In_3708,In_132);
or U6329 (N_6329,In_2070,In_2666);
nand U6330 (N_6330,In_642,In_653);
or U6331 (N_6331,In_1762,In_2645);
nor U6332 (N_6332,In_866,In_2632);
nor U6333 (N_6333,In_4532,In_3858);
nand U6334 (N_6334,In_3231,In_579);
xor U6335 (N_6335,In_1276,In_989);
nor U6336 (N_6336,In_644,In_4918);
xor U6337 (N_6337,In_872,In_593);
xor U6338 (N_6338,In_3421,In_4882);
and U6339 (N_6339,In_657,In_4183);
xnor U6340 (N_6340,In_3281,In_1261);
xnor U6341 (N_6341,In_793,In_4808);
nand U6342 (N_6342,In_3249,In_4854);
nand U6343 (N_6343,In_2481,In_2928);
xnor U6344 (N_6344,In_3471,In_3707);
nor U6345 (N_6345,In_1225,In_3325);
and U6346 (N_6346,In_2683,In_2250);
and U6347 (N_6347,In_3687,In_4096);
nand U6348 (N_6348,In_2288,In_1596);
and U6349 (N_6349,In_28,In_1169);
and U6350 (N_6350,In_4651,In_355);
or U6351 (N_6351,In_4320,In_356);
nor U6352 (N_6352,In_4203,In_781);
xnor U6353 (N_6353,In_1508,In_3028);
and U6354 (N_6354,In_2456,In_4747);
nor U6355 (N_6355,In_4936,In_245);
nor U6356 (N_6356,In_4697,In_1707);
nor U6357 (N_6357,In_2292,In_3216);
nand U6358 (N_6358,In_3992,In_2839);
nand U6359 (N_6359,In_4536,In_3959);
nor U6360 (N_6360,In_2291,In_2177);
or U6361 (N_6361,In_3660,In_1858);
or U6362 (N_6362,In_3060,In_3563);
or U6363 (N_6363,In_3102,In_927);
and U6364 (N_6364,In_258,In_2966);
nand U6365 (N_6365,In_3757,In_53);
nor U6366 (N_6366,In_4043,In_288);
and U6367 (N_6367,In_2035,In_495);
or U6368 (N_6368,In_4144,In_4250);
nor U6369 (N_6369,In_3005,In_1362);
or U6370 (N_6370,In_3969,In_2950);
or U6371 (N_6371,In_2508,In_2031);
or U6372 (N_6372,In_3817,In_1920);
or U6373 (N_6373,In_1257,In_4460);
nand U6374 (N_6374,In_3527,In_4215);
xor U6375 (N_6375,In_3563,In_4824);
nand U6376 (N_6376,In_644,In_1600);
nand U6377 (N_6377,In_931,In_3356);
and U6378 (N_6378,In_1680,In_1242);
nand U6379 (N_6379,In_4443,In_37);
xor U6380 (N_6380,In_4347,In_4316);
xor U6381 (N_6381,In_1262,In_4422);
or U6382 (N_6382,In_3153,In_46);
nor U6383 (N_6383,In_1295,In_2629);
nor U6384 (N_6384,In_1900,In_566);
xor U6385 (N_6385,In_3873,In_2238);
nor U6386 (N_6386,In_52,In_386);
and U6387 (N_6387,In_2280,In_557);
xnor U6388 (N_6388,In_3633,In_1166);
or U6389 (N_6389,In_2746,In_628);
nand U6390 (N_6390,In_4667,In_516);
nand U6391 (N_6391,In_2969,In_3453);
nand U6392 (N_6392,In_4313,In_3637);
and U6393 (N_6393,In_1007,In_111);
and U6394 (N_6394,In_2689,In_2380);
or U6395 (N_6395,In_2384,In_76);
nand U6396 (N_6396,In_2005,In_1666);
xor U6397 (N_6397,In_3784,In_1358);
xor U6398 (N_6398,In_3416,In_393);
or U6399 (N_6399,In_238,In_2123);
or U6400 (N_6400,In_2835,In_1608);
xnor U6401 (N_6401,In_3678,In_1979);
nand U6402 (N_6402,In_2643,In_4591);
nor U6403 (N_6403,In_2217,In_3386);
and U6404 (N_6404,In_3220,In_765);
or U6405 (N_6405,In_2223,In_2453);
nor U6406 (N_6406,In_3481,In_1082);
or U6407 (N_6407,In_3393,In_872);
nand U6408 (N_6408,In_687,In_4120);
and U6409 (N_6409,In_2572,In_17);
or U6410 (N_6410,In_1229,In_3569);
xor U6411 (N_6411,In_4800,In_178);
or U6412 (N_6412,In_531,In_3123);
xor U6413 (N_6413,In_2776,In_4058);
or U6414 (N_6414,In_4023,In_4006);
and U6415 (N_6415,In_3372,In_4437);
xor U6416 (N_6416,In_3048,In_1599);
xnor U6417 (N_6417,In_1424,In_2726);
xor U6418 (N_6418,In_1638,In_3432);
and U6419 (N_6419,In_825,In_3551);
xnor U6420 (N_6420,In_1720,In_4285);
or U6421 (N_6421,In_666,In_3466);
and U6422 (N_6422,In_187,In_1692);
nand U6423 (N_6423,In_797,In_1331);
nand U6424 (N_6424,In_2761,In_327);
nor U6425 (N_6425,In_4,In_2262);
nand U6426 (N_6426,In_1899,In_3152);
nand U6427 (N_6427,In_3853,In_156);
or U6428 (N_6428,In_2066,In_1659);
nand U6429 (N_6429,In_2312,In_224);
xnor U6430 (N_6430,In_3917,In_4023);
nor U6431 (N_6431,In_649,In_2779);
nand U6432 (N_6432,In_4361,In_3435);
xnor U6433 (N_6433,In_2075,In_1423);
or U6434 (N_6434,In_3507,In_2399);
nand U6435 (N_6435,In_536,In_4543);
xnor U6436 (N_6436,In_4809,In_553);
nor U6437 (N_6437,In_936,In_3067);
or U6438 (N_6438,In_3055,In_2712);
and U6439 (N_6439,In_2690,In_2213);
xor U6440 (N_6440,In_4729,In_2436);
nor U6441 (N_6441,In_4216,In_4218);
or U6442 (N_6442,In_3516,In_4820);
nor U6443 (N_6443,In_1133,In_1342);
and U6444 (N_6444,In_4754,In_2500);
xnor U6445 (N_6445,In_3141,In_3091);
nor U6446 (N_6446,In_2464,In_3779);
nor U6447 (N_6447,In_644,In_2505);
nor U6448 (N_6448,In_4757,In_4387);
nor U6449 (N_6449,In_2860,In_3943);
xor U6450 (N_6450,In_1415,In_4933);
xor U6451 (N_6451,In_2074,In_3191);
and U6452 (N_6452,In_2044,In_2092);
xor U6453 (N_6453,In_1071,In_2023);
nand U6454 (N_6454,In_551,In_4859);
nor U6455 (N_6455,In_4405,In_847);
or U6456 (N_6456,In_1124,In_35);
or U6457 (N_6457,In_1070,In_3166);
nor U6458 (N_6458,In_3583,In_2191);
and U6459 (N_6459,In_4905,In_2411);
nor U6460 (N_6460,In_4104,In_557);
nand U6461 (N_6461,In_3226,In_1102);
and U6462 (N_6462,In_960,In_3666);
and U6463 (N_6463,In_810,In_1483);
nor U6464 (N_6464,In_4635,In_4272);
xnor U6465 (N_6465,In_1557,In_4187);
or U6466 (N_6466,In_2664,In_4789);
nor U6467 (N_6467,In_3406,In_1757);
or U6468 (N_6468,In_4708,In_128);
or U6469 (N_6469,In_1330,In_4958);
xor U6470 (N_6470,In_1737,In_1629);
or U6471 (N_6471,In_3586,In_27);
nand U6472 (N_6472,In_645,In_2122);
or U6473 (N_6473,In_348,In_1011);
or U6474 (N_6474,In_4005,In_682);
nor U6475 (N_6475,In_4831,In_3445);
or U6476 (N_6476,In_3467,In_1878);
and U6477 (N_6477,In_3446,In_3046);
nand U6478 (N_6478,In_19,In_1465);
and U6479 (N_6479,In_996,In_732);
nand U6480 (N_6480,In_2705,In_2558);
and U6481 (N_6481,In_4897,In_983);
and U6482 (N_6482,In_2689,In_203);
or U6483 (N_6483,In_1111,In_4443);
and U6484 (N_6484,In_1057,In_2151);
xnor U6485 (N_6485,In_1193,In_3447);
nand U6486 (N_6486,In_410,In_1253);
xor U6487 (N_6487,In_1004,In_1978);
nor U6488 (N_6488,In_4535,In_4903);
xnor U6489 (N_6489,In_4605,In_1055);
nand U6490 (N_6490,In_467,In_3562);
or U6491 (N_6491,In_3323,In_1942);
xor U6492 (N_6492,In_2719,In_3807);
nand U6493 (N_6493,In_4733,In_2808);
nand U6494 (N_6494,In_2268,In_1219);
nor U6495 (N_6495,In_1919,In_1618);
and U6496 (N_6496,In_4835,In_4259);
nor U6497 (N_6497,In_821,In_3334);
and U6498 (N_6498,In_3370,In_210);
xnor U6499 (N_6499,In_903,In_4846);
or U6500 (N_6500,In_1363,In_1129);
nor U6501 (N_6501,In_4532,In_2510);
and U6502 (N_6502,In_2672,In_491);
and U6503 (N_6503,In_234,In_3430);
nor U6504 (N_6504,In_3117,In_3390);
nand U6505 (N_6505,In_3882,In_1949);
nand U6506 (N_6506,In_303,In_1768);
xnor U6507 (N_6507,In_3330,In_1580);
and U6508 (N_6508,In_3049,In_1339);
or U6509 (N_6509,In_4583,In_1338);
nor U6510 (N_6510,In_4563,In_1952);
or U6511 (N_6511,In_347,In_765);
nor U6512 (N_6512,In_1759,In_2450);
xor U6513 (N_6513,In_4199,In_2978);
and U6514 (N_6514,In_4781,In_3267);
xor U6515 (N_6515,In_2509,In_3742);
or U6516 (N_6516,In_3094,In_1126);
xnor U6517 (N_6517,In_1091,In_4076);
nor U6518 (N_6518,In_1189,In_2850);
nand U6519 (N_6519,In_4395,In_1054);
or U6520 (N_6520,In_131,In_1374);
nor U6521 (N_6521,In_3630,In_2120);
nor U6522 (N_6522,In_3225,In_3833);
nor U6523 (N_6523,In_2092,In_144);
or U6524 (N_6524,In_3926,In_3374);
nor U6525 (N_6525,In_194,In_740);
nand U6526 (N_6526,In_518,In_15);
xnor U6527 (N_6527,In_3614,In_3538);
nand U6528 (N_6528,In_1505,In_3448);
xor U6529 (N_6529,In_532,In_4583);
and U6530 (N_6530,In_2528,In_4715);
xnor U6531 (N_6531,In_2844,In_1113);
or U6532 (N_6532,In_3371,In_4646);
nand U6533 (N_6533,In_2160,In_2638);
nor U6534 (N_6534,In_4316,In_4395);
nor U6535 (N_6535,In_4,In_4240);
xnor U6536 (N_6536,In_4589,In_2821);
or U6537 (N_6537,In_2654,In_464);
xnor U6538 (N_6538,In_200,In_2627);
and U6539 (N_6539,In_3300,In_1522);
or U6540 (N_6540,In_4952,In_3159);
nand U6541 (N_6541,In_510,In_1894);
or U6542 (N_6542,In_1677,In_2572);
nand U6543 (N_6543,In_254,In_242);
xor U6544 (N_6544,In_1525,In_412);
or U6545 (N_6545,In_4744,In_363);
nor U6546 (N_6546,In_1176,In_2172);
and U6547 (N_6547,In_2182,In_2468);
and U6548 (N_6548,In_4531,In_3745);
and U6549 (N_6549,In_3254,In_1269);
nand U6550 (N_6550,In_4586,In_2611);
xnor U6551 (N_6551,In_655,In_2104);
and U6552 (N_6552,In_3180,In_4512);
nor U6553 (N_6553,In_3438,In_3461);
xor U6554 (N_6554,In_3539,In_3865);
nand U6555 (N_6555,In_2779,In_2357);
nand U6556 (N_6556,In_3921,In_1862);
nand U6557 (N_6557,In_2029,In_4034);
nor U6558 (N_6558,In_2490,In_3572);
nor U6559 (N_6559,In_1367,In_3966);
nor U6560 (N_6560,In_3989,In_4872);
nor U6561 (N_6561,In_4578,In_1344);
nor U6562 (N_6562,In_3785,In_3518);
nor U6563 (N_6563,In_614,In_4404);
and U6564 (N_6564,In_3739,In_2701);
and U6565 (N_6565,In_2242,In_926);
and U6566 (N_6566,In_2211,In_4801);
and U6567 (N_6567,In_2043,In_3895);
or U6568 (N_6568,In_964,In_4751);
xnor U6569 (N_6569,In_353,In_2343);
nand U6570 (N_6570,In_2446,In_731);
xor U6571 (N_6571,In_3800,In_663);
nor U6572 (N_6572,In_4467,In_1209);
and U6573 (N_6573,In_800,In_102);
nor U6574 (N_6574,In_2877,In_1529);
or U6575 (N_6575,In_807,In_110);
nor U6576 (N_6576,In_2529,In_3097);
xnor U6577 (N_6577,In_3356,In_1042);
nor U6578 (N_6578,In_698,In_3972);
or U6579 (N_6579,In_2845,In_4302);
xor U6580 (N_6580,In_3841,In_2298);
and U6581 (N_6581,In_3502,In_121);
xnor U6582 (N_6582,In_4901,In_3816);
nor U6583 (N_6583,In_1733,In_2205);
xnor U6584 (N_6584,In_75,In_4293);
nand U6585 (N_6585,In_225,In_3959);
and U6586 (N_6586,In_2438,In_2652);
nand U6587 (N_6587,In_2345,In_2477);
or U6588 (N_6588,In_246,In_3745);
nand U6589 (N_6589,In_4361,In_4930);
nand U6590 (N_6590,In_3722,In_3727);
or U6591 (N_6591,In_4340,In_3169);
and U6592 (N_6592,In_849,In_3986);
nand U6593 (N_6593,In_874,In_4334);
nand U6594 (N_6594,In_3415,In_600);
and U6595 (N_6595,In_2459,In_1386);
nor U6596 (N_6596,In_1107,In_1484);
nor U6597 (N_6597,In_2069,In_2899);
xor U6598 (N_6598,In_2151,In_2193);
nor U6599 (N_6599,In_1974,In_3116);
nand U6600 (N_6600,In_3020,In_2896);
xnor U6601 (N_6601,In_1180,In_1159);
and U6602 (N_6602,In_3748,In_3886);
xnor U6603 (N_6603,In_4679,In_3708);
nand U6604 (N_6604,In_1272,In_3999);
nor U6605 (N_6605,In_401,In_4792);
nand U6606 (N_6606,In_3614,In_2585);
xor U6607 (N_6607,In_3707,In_3211);
and U6608 (N_6608,In_10,In_146);
or U6609 (N_6609,In_1266,In_3228);
and U6610 (N_6610,In_2165,In_1509);
nor U6611 (N_6611,In_4170,In_3836);
or U6612 (N_6612,In_2152,In_4769);
nor U6613 (N_6613,In_257,In_3298);
nor U6614 (N_6614,In_240,In_3232);
or U6615 (N_6615,In_2735,In_2322);
nor U6616 (N_6616,In_394,In_2159);
and U6617 (N_6617,In_2071,In_2204);
xnor U6618 (N_6618,In_1545,In_2285);
nand U6619 (N_6619,In_1516,In_2225);
nand U6620 (N_6620,In_434,In_4463);
nor U6621 (N_6621,In_3328,In_2515);
nand U6622 (N_6622,In_2652,In_4057);
and U6623 (N_6623,In_1712,In_1357);
xnor U6624 (N_6624,In_3364,In_4496);
or U6625 (N_6625,In_430,In_2734);
xor U6626 (N_6626,In_4147,In_4841);
nand U6627 (N_6627,In_2771,In_1143);
nand U6628 (N_6628,In_3846,In_1458);
nand U6629 (N_6629,In_4813,In_1978);
and U6630 (N_6630,In_3910,In_2914);
and U6631 (N_6631,In_2378,In_2870);
and U6632 (N_6632,In_4251,In_1741);
and U6633 (N_6633,In_1429,In_3664);
and U6634 (N_6634,In_4213,In_4532);
nand U6635 (N_6635,In_3896,In_1807);
nand U6636 (N_6636,In_4914,In_1012);
or U6637 (N_6637,In_3205,In_405);
xnor U6638 (N_6638,In_1226,In_755);
nor U6639 (N_6639,In_3097,In_4357);
or U6640 (N_6640,In_2861,In_192);
xor U6641 (N_6641,In_2459,In_2134);
nand U6642 (N_6642,In_2853,In_281);
and U6643 (N_6643,In_3839,In_2261);
and U6644 (N_6644,In_2996,In_2127);
and U6645 (N_6645,In_2373,In_1779);
nor U6646 (N_6646,In_4432,In_3154);
and U6647 (N_6647,In_170,In_4011);
or U6648 (N_6648,In_1042,In_4870);
or U6649 (N_6649,In_1492,In_4185);
and U6650 (N_6650,In_2665,In_1034);
nor U6651 (N_6651,In_441,In_4948);
nand U6652 (N_6652,In_1452,In_4486);
and U6653 (N_6653,In_3618,In_3778);
or U6654 (N_6654,In_613,In_1994);
xnor U6655 (N_6655,In_4065,In_2553);
xnor U6656 (N_6656,In_757,In_4686);
and U6657 (N_6657,In_1463,In_3438);
xnor U6658 (N_6658,In_1502,In_727);
nand U6659 (N_6659,In_4953,In_1495);
and U6660 (N_6660,In_2217,In_312);
nor U6661 (N_6661,In_3928,In_526);
nand U6662 (N_6662,In_3067,In_357);
xor U6663 (N_6663,In_421,In_1430);
nand U6664 (N_6664,In_1587,In_888);
xor U6665 (N_6665,In_3584,In_2167);
and U6666 (N_6666,In_4261,In_3512);
and U6667 (N_6667,In_4532,In_587);
and U6668 (N_6668,In_1343,In_365);
xnor U6669 (N_6669,In_616,In_63);
and U6670 (N_6670,In_4320,In_2848);
nor U6671 (N_6671,In_2065,In_4584);
and U6672 (N_6672,In_4876,In_359);
and U6673 (N_6673,In_3523,In_2178);
or U6674 (N_6674,In_4038,In_3250);
nand U6675 (N_6675,In_81,In_3068);
or U6676 (N_6676,In_1354,In_1414);
or U6677 (N_6677,In_324,In_432);
nand U6678 (N_6678,In_4654,In_2489);
nor U6679 (N_6679,In_2938,In_3961);
nand U6680 (N_6680,In_2933,In_712);
and U6681 (N_6681,In_3168,In_4380);
nand U6682 (N_6682,In_1806,In_2254);
nand U6683 (N_6683,In_1117,In_2516);
xnor U6684 (N_6684,In_3034,In_4941);
nor U6685 (N_6685,In_4318,In_1151);
and U6686 (N_6686,In_4848,In_1967);
nand U6687 (N_6687,In_2377,In_887);
or U6688 (N_6688,In_4619,In_528);
nand U6689 (N_6689,In_2613,In_3267);
nor U6690 (N_6690,In_3735,In_1993);
nand U6691 (N_6691,In_2799,In_1801);
nor U6692 (N_6692,In_4769,In_2884);
xnor U6693 (N_6693,In_4428,In_4520);
or U6694 (N_6694,In_1315,In_1342);
nand U6695 (N_6695,In_1152,In_2754);
nor U6696 (N_6696,In_1375,In_1012);
and U6697 (N_6697,In_2443,In_862);
or U6698 (N_6698,In_3502,In_4126);
and U6699 (N_6699,In_437,In_1388);
or U6700 (N_6700,In_567,In_3993);
and U6701 (N_6701,In_4006,In_2325);
and U6702 (N_6702,In_1,In_4647);
xnor U6703 (N_6703,In_2154,In_1999);
and U6704 (N_6704,In_1952,In_1402);
nand U6705 (N_6705,In_834,In_4264);
and U6706 (N_6706,In_1729,In_145);
nor U6707 (N_6707,In_3638,In_3865);
or U6708 (N_6708,In_942,In_3819);
nor U6709 (N_6709,In_1959,In_2695);
xnor U6710 (N_6710,In_2770,In_3258);
nor U6711 (N_6711,In_2038,In_266);
or U6712 (N_6712,In_3284,In_4640);
and U6713 (N_6713,In_3330,In_2276);
and U6714 (N_6714,In_2468,In_3053);
xor U6715 (N_6715,In_2880,In_745);
nand U6716 (N_6716,In_4385,In_1433);
xnor U6717 (N_6717,In_448,In_3316);
xor U6718 (N_6718,In_4800,In_171);
xnor U6719 (N_6719,In_4860,In_134);
nor U6720 (N_6720,In_3427,In_868);
xor U6721 (N_6721,In_1186,In_3811);
and U6722 (N_6722,In_4826,In_1867);
nor U6723 (N_6723,In_3283,In_2941);
nor U6724 (N_6724,In_4934,In_2634);
nand U6725 (N_6725,In_3551,In_2515);
nand U6726 (N_6726,In_4827,In_1798);
or U6727 (N_6727,In_4970,In_2549);
nand U6728 (N_6728,In_4719,In_3807);
nand U6729 (N_6729,In_3189,In_2199);
nor U6730 (N_6730,In_2519,In_924);
and U6731 (N_6731,In_389,In_2262);
or U6732 (N_6732,In_1441,In_846);
nand U6733 (N_6733,In_226,In_1574);
and U6734 (N_6734,In_2104,In_2992);
nand U6735 (N_6735,In_1281,In_2204);
or U6736 (N_6736,In_868,In_1818);
nand U6737 (N_6737,In_475,In_1733);
or U6738 (N_6738,In_216,In_1666);
and U6739 (N_6739,In_4234,In_3879);
and U6740 (N_6740,In_4212,In_182);
or U6741 (N_6741,In_52,In_1948);
xor U6742 (N_6742,In_3840,In_3755);
and U6743 (N_6743,In_4608,In_1982);
and U6744 (N_6744,In_563,In_4628);
and U6745 (N_6745,In_830,In_93);
or U6746 (N_6746,In_4827,In_4803);
nor U6747 (N_6747,In_3989,In_3442);
nand U6748 (N_6748,In_3116,In_1417);
xor U6749 (N_6749,In_788,In_2436);
xnor U6750 (N_6750,In_3914,In_320);
and U6751 (N_6751,In_2899,In_3988);
or U6752 (N_6752,In_1182,In_1823);
nor U6753 (N_6753,In_2949,In_2884);
nand U6754 (N_6754,In_3266,In_2679);
or U6755 (N_6755,In_4900,In_4397);
nand U6756 (N_6756,In_3903,In_2054);
nor U6757 (N_6757,In_4880,In_3392);
or U6758 (N_6758,In_4263,In_2259);
nor U6759 (N_6759,In_1821,In_2441);
nor U6760 (N_6760,In_2813,In_76);
nor U6761 (N_6761,In_4649,In_2788);
nor U6762 (N_6762,In_4332,In_2288);
nor U6763 (N_6763,In_3649,In_3871);
and U6764 (N_6764,In_633,In_1494);
and U6765 (N_6765,In_3598,In_2777);
nor U6766 (N_6766,In_533,In_3259);
and U6767 (N_6767,In_2350,In_1055);
nand U6768 (N_6768,In_2325,In_2344);
nor U6769 (N_6769,In_3250,In_1080);
nor U6770 (N_6770,In_4437,In_555);
nand U6771 (N_6771,In_1323,In_2458);
nand U6772 (N_6772,In_2403,In_4735);
xnor U6773 (N_6773,In_1406,In_314);
or U6774 (N_6774,In_1654,In_49);
nand U6775 (N_6775,In_859,In_4938);
or U6776 (N_6776,In_3710,In_4073);
xor U6777 (N_6777,In_4908,In_447);
nand U6778 (N_6778,In_4233,In_1953);
and U6779 (N_6779,In_2544,In_2670);
nand U6780 (N_6780,In_3509,In_2991);
and U6781 (N_6781,In_3997,In_1573);
nor U6782 (N_6782,In_965,In_952);
and U6783 (N_6783,In_2910,In_3044);
nand U6784 (N_6784,In_3445,In_1080);
xor U6785 (N_6785,In_4183,In_1499);
nand U6786 (N_6786,In_603,In_3280);
nor U6787 (N_6787,In_3009,In_3710);
xnor U6788 (N_6788,In_3073,In_276);
or U6789 (N_6789,In_1716,In_4752);
and U6790 (N_6790,In_2103,In_3317);
and U6791 (N_6791,In_4320,In_4046);
nor U6792 (N_6792,In_4335,In_4421);
xnor U6793 (N_6793,In_91,In_4046);
or U6794 (N_6794,In_2148,In_4201);
and U6795 (N_6795,In_427,In_1804);
or U6796 (N_6796,In_1833,In_2023);
nand U6797 (N_6797,In_3492,In_3334);
or U6798 (N_6798,In_4252,In_4639);
nand U6799 (N_6799,In_4506,In_3874);
or U6800 (N_6800,In_2852,In_4372);
xor U6801 (N_6801,In_3367,In_2153);
xor U6802 (N_6802,In_10,In_1377);
xor U6803 (N_6803,In_2120,In_3490);
xnor U6804 (N_6804,In_219,In_161);
xor U6805 (N_6805,In_865,In_1181);
nor U6806 (N_6806,In_4141,In_3778);
nor U6807 (N_6807,In_4958,In_1788);
nand U6808 (N_6808,In_235,In_4376);
xnor U6809 (N_6809,In_1182,In_1528);
nand U6810 (N_6810,In_4454,In_616);
nand U6811 (N_6811,In_3530,In_3276);
xnor U6812 (N_6812,In_4619,In_3248);
nand U6813 (N_6813,In_2567,In_4820);
nor U6814 (N_6814,In_4106,In_101);
or U6815 (N_6815,In_1553,In_2188);
or U6816 (N_6816,In_6,In_3330);
nand U6817 (N_6817,In_1806,In_289);
or U6818 (N_6818,In_94,In_3881);
or U6819 (N_6819,In_355,In_1391);
nor U6820 (N_6820,In_2057,In_1648);
nor U6821 (N_6821,In_737,In_1480);
nor U6822 (N_6822,In_992,In_2004);
nand U6823 (N_6823,In_1358,In_1397);
nor U6824 (N_6824,In_1117,In_3786);
nor U6825 (N_6825,In_3328,In_3796);
and U6826 (N_6826,In_3470,In_1219);
nor U6827 (N_6827,In_4886,In_4152);
xor U6828 (N_6828,In_4172,In_3604);
nand U6829 (N_6829,In_221,In_1758);
or U6830 (N_6830,In_4544,In_3750);
and U6831 (N_6831,In_2202,In_1783);
nand U6832 (N_6832,In_4605,In_4417);
or U6833 (N_6833,In_4120,In_4353);
or U6834 (N_6834,In_1348,In_3470);
xor U6835 (N_6835,In_903,In_2313);
nor U6836 (N_6836,In_2183,In_2107);
nand U6837 (N_6837,In_2325,In_3512);
and U6838 (N_6838,In_1847,In_3405);
and U6839 (N_6839,In_3093,In_3806);
nor U6840 (N_6840,In_2941,In_1621);
or U6841 (N_6841,In_1841,In_1670);
nor U6842 (N_6842,In_4599,In_3552);
xnor U6843 (N_6843,In_428,In_2593);
xor U6844 (N_6844,In_3696,In_1746);
or U6845 (N_6845,In_2361,In_1905);
or U6846 (N_6846,In_1679,In_218);
nand U6847 (N_6847,In_3591,In_4427);
nor U6848 (N_6848,In_3846,In_1);
nor U6849 (N_6849,In_174,In_3894);
nand U6850 (N_6850,In_3135,In_2761);
xnor U6851 (N_6851,In_4496,In_2865);
nor U6852 (N_6852,In_2088,In_1137);
or U6853 (N_6853,In_675,In_3813);
nand U6854 (N_6854,In_3354,In_2836);
nand U6855 (N_6855,In_4049,In_4560);
or U6856 (N_6856,In_3799,In_1500);
nand U6857 (N_6857,In_2627,In_1358);
xor U6858 (N_6858,In_2191,In_2374);
nand U6859 (N_6859,In_339,In_240);
nor U6860 (N_6860,In_2250,In_3717);
nor U6861 (N_6861,In_2789,In_3654);
or U6862 (N_6862,In_21,In_4879);
or U6863 (N_6863,In_3593,In_3959);
xnor U6864 (N_6864,In_517,In_4251);
nand U6865 (N_6865,In_2768,In_4506);
nor U6866 (N_6866,In_834,In_3966);
or U6867 (N_6867,In_113,In_2939);
or U6868 (N_6868,In_3236,In_3310);
nor U6869 (N_6869,In_2167,In_335);
or U6870 (N_6870,In_1999,In_841);
nand U6871 (N_6871,In_1716,In_2862);
or U6872 (N_6872,In_4307,In_3320);
xnor U6873 (N_6873,In_1335,In_705);
or U6874 (N_6874,In_1726,In_3746);
xnor U6875 (N_6875,In_1459,In_3927);
xnor U6876 (N_6876,In_2391,In_1169);
and U6877 (N_6877,In_4027,In_3207);
and U6878 (N_6878,In_3843,In_831);
nand U6879 (N_6879,In_4984,In_3176);
or U6880 (N_6880,In_4396,In_2348);
and U6881 (N_6881,In_1354,In_4099);
or U6882 (N_6882,In_1959,In_3918);
xor U6883 (N_6883,In_4029,In_3708);
and U6884 (N_6884,In_3192,In_1375);
nand U6885 (N_6885,In_3377,In_3315);
nand U6886 (N_6886,In_125,In_485);
nor U6887 (N_6887,In_2429,In_4011);
and U6888 (N_6888,In_929,In_941);
nor U6889 (N_6889,In_4929,In_4066);
and U6890 (N_6890,In_4715,In_218);
nand U6891 (N_6891,In_3930,In_1986);
nor U6892 (N_6892,In_649,In_1254);
and U6893 (N_6893,In_3651,In_160);
nor U6894 (N_6894,In_2596,In_153);
nand U6895 (N_6895,In_1896,In_2131);
nand U6896 (N_6896,In_420,In_1134);
nor U6897 (N_6897,In_3740,In_695);
nor U6898 (N_6898,In_1642,In_1183);
or U6899 (N_6899,In_333,In_3812);
nor U6900 (N_6900,In_1798,In_2411);
xnor U6901 (N_6901,In_2134,In_2097);
xnor U6902 (N_6902,In_4220,In_233);
and U6903 (N_6903,In_960,In_4066);
nand U6904 (N_6904,In_1892,In_4247);
nor U6905 (N_6905,In_360,In_446);
nand U6906 (N_6906,In_3209,In_1290);
nor U6907 (N_6907,In_448,In_3424);
nand U6908 (N_6908,In_1864,In_2253);
and U6909 (N_6909,In_4021,In_2464);
or U6910 (N_6910,In_691,In_1184);
and U6911 (N_6911,In_2687,In_4440);
and U6912 (N_6912,In_4332,In_383);
nand U6913 (N_6913,In_3126,In_3003);
nand U6914 (N_6914,In_3197,In_3774);
xnor U6915 (N_6915,In_1585,In_401);
or U6916 (N_6916,In_3928,In_2104);
nor U6917 (N_6917,In_866,In_1807);
nor U6918 (N_6918,In_1199,In_1040);
nand U6919 (N_6919,In_2567,In_247);
nand U6920 (N_6920,In_1308,In_3588);
nand U6921 (N_6921,In_3529,In_3149);
and U6922 (N_6922,In_4994,In_2925);
nand U6923 (N_6923,In_3878,In_1847);
and U6924 (N_6924,In_1370,In_2384);
nor U6925 (N_6925,In_932,In_2814);
nand U6926 (N_6926,In_2760,In_1349);
or U6927 (N_6927,In_2264,In_3870);
and U6928 (N_6928,In_1164,In_3572);
or U6929 (N_6929,In_2389,In_4880);
or U6930 (N_6930,In_1419,In_635);
and U6931 (N_6931,In_3509,In_732);
xnor U6932 (N_6932,In_1117,In_1998);
or U6933 (N_6933,In_2838,In_3857);
nand U6934 (N_6934,In_3954,In_3570);
nor U6935 (N_6935,In_28,In_3375);
nand U6936 (N_6936,In_485,In_2212);
nor U6937 (N_6937,In_1587,In_439);
nor U6938 (N_6938,In_1763,In_3625);
or U6939 (N_6939,In_644,In_557);
nor U6940 (N_6940,In_3701,In_4071);
and U6941 (N_6941,In_3840,In_4326);
xnor U6942 (N_6942,In_250,In_300);
xor U6943 (N_6943,In_1185,In_2075);
or U6944 (N_6944,In_4072,In_3477);
or U6945 (N_6945,In_1584,In_1236);
nor U6946 (N_6946,In_3088,In_2567);
nand U6947 (N_6947,In_651,In_261);
xnor U6948 (N_6948,In_1272,In_4504);
xor U6949 (N_6949,In_3037,In_1900);
nor U6950 (N_6950,In_3472,In_3959);
and U6951 (N_6951,In_1705,In_1653);
and U6952 (N_6952,In_3272,In_3094);
or U6953 (N_6953,In_4701,In_4270);
xnor U6954 (N_6954,In_1518,In_667);
nand U6955 (N_6955,In_4685,In_4377);
or U6956 (N_6956,In_2466,In_2746);
nand U6957 (N_6957,In_2494,In_2009);
or U6958 (N_6958,In_4175,In_1378);
and U6959 (N_6959,In_3381,In_1269);
or U6960 (N_6960,In_887,In_3053);
nor U6961 (N_6961,In_4772,In_1280);
or U6962 (N_6962,In_3066,In_2403);
or U6963 (N_6963,In_479,In_4654);
or U6964 (N_6964,In_3504,In_3475);
nor U6965 (N_6965,In_1434,In_1157);
nand U6966 (N_6966,In_2338,In_4191);
nor U6967 (N_6967,In_464,In_1184);
or U6968 (N_6968,In_4739,In_1217);
nand U6969 (N_6969,In_3265,In_2089);
nor U6970 (N_6970,In_1003,In_3924);
or U6971 (N_6971,In_2262,In_1399);
xor U6972 (N_6972,In_4338,In_4445);
or U6973 (N_6973,In_2516,In_4341);
and U6974 (N_6974,In_730,In_3895);
xnor U6975 (N_6975,In_1506,In_1153);
and U6976 (N_6976,In_2520,In_2281);
nand U6977 (N_6977,In_2843,In_2260);
or U6978 (N_6978,In_3844,In_3429);
xor U6979 (N_6979,In_2366,In_2554);
nand U6980 (N_6980,In_1537,In_4862);
and U6981 (N_6981,In_342,In_453);
and U6982 (N_6982,In_1977,In_2814);
and U6983 (N_6983,In_3743,In_2566);
nand U6984 (N_6984,In_3609,In_1539);
or U6985 (N_6985,In_4908,In_70);
nor U6986 (N_6986,In_4383,In_1501);
nand U6987 (N_6987,In_841,In_4747);
xor U6988 (N_6988,In_1527,In_1481);
and U6989 (N_6989,In_460,In_3623);
nand U6990 (N_6990,In_434,In_4955);
nand U6991 (N_6991,In_3556,In_766);
nand U6992 (N_6992,In_671,In_4321);
nor U6993 (N_6993,In_700,In_3415);
and U6994 (N_6994,In_4905,In_366);
or U6995 (N_6995,In_110,In_4483);
nand U6996 (N_6996,In_2368,In_2171);
nand U6997 (N_6997,In_301,In_4041);
or U6998 (N_6998,In_30,In_2256);
xor U6999 (N_6999,In_849,In_4973);
xnor U7000 (N_7000,In_1232,In_4876);
or U7001 (N_7001,In_4259,In_2584);
nand U7002 (N_7002,In_4748,In_2342);
nor U7003 (N_7003,In_702,In_4036);
nor U7004 (N_7004,In_3314,In_3684);
nand U7005 (N_7005,In_4657,In_2949);
xnor U7006 (N_7006,In_780,In_4418);
nor U7007 (N_7007,In_3360,In_3723);
xnor U7008 (N_7008,In_464,In_701);
and U7009 (N_7009,In_3149,In_1076);
and U7010 (N_7010,In_2383,In_1423);
or U7011 (N_7011,In_1501,In_2538);
xnor U7012 (N_7012,In_2748,In_2532);
nand U7013 (N_7013,In_2967,In_446);
xor U7014 (N_7014,In_4590,In_1688);
xor U7015 (N_7015,In_3213,In_4653);
nand U7016 (N_7016,In_2348,In_3212);
and U7017 (N_7017,In_2742,In_1694);
nand U7018 (N_7018,In_1001,In_1972);
nand U7019 (N_7019,In_2447,In_2454);
or U7020 (N_7020,In_3590,In_2975);
or U7021 (N_7021,In_3314,In_4444);
and U7022 (N_7022,In_3792,In_1619);
nand U7023 (N_7023,In_2422,In_391);
nand U7024 (N_7024,In_1207,In_2424);
nand U7025 (N_7025,In_3649,In_292);
or U7026 (N_7026,In_236,In_1506);
xor U7027 (N_7027,In_2834,In_4514);
nor U7028 (N_7028,In_942,In_134);
nor U7029 (N_7029,In_763,In_321);
or U7030 (N_7030,In_1924,In_1921);
nor U7031 (N_7031,In_3103,In_4415);
and U7032 (N_7032,In_2791,In_3140);
xnor U7033 (N_7033,In_479,In_4092);
xor U7034 (N_7034,In_1923,In_610);
or U7035 (N_7035,In_2125,In_758);
or U7036 (N_7036,In_1242,In_4955);
xnor U7037 (N_7037,In_1761,In_3278);
xnor U7038 (N_7038,In_4500,In_2976);
nor U7039 (N_7039,In_205,In_1460);
and U7040 (N_7040,In_1516,In_1689);
xor U7041 (N_7041,In_830,In_4704);
nor U7042 (N_7042,In_2774,In_1147);
nor U7043 (N_7043,In_154,In_1533);
nor U7044 (N_7044,In_3998,In_752);
nand U7045 (N_7045,In_25,In_3456);
nand U7046 (N_7046,In_4333,In_2614);
nor U7047 (N_7047,In_4137,In_2479);
xnor U7048 (N_7048,In_817,In_4813);
xor U7049 (N_7049,In_2671,In_4497);
nand U7050 (N_7050,In_1169,In_3825);
nand U7051 (N_7051,In_3457,In_613);
xnor U7052 (N_7052,In_3047,In_4058);
nor U7053 (N_7053,In_1120,In_106);
xor U7054 (N_7054,In_1899,In_3966);
nand U7055 (N_7055,In_4097,In_59);
xnor U7056 (N_7056,In_3351,In_728);
xor U7057 (N_7057,In_4211,In_1708);
nor U7058 (N_7058,In_2641,In_3406);
or U7059 (N_7059,In_839,In_2659);
nor U7060 (N_7060,In_2768,In_3487);
xnor U7061 (N_7061,In_241,In_4796);
nand U7062 (N_7062,In_4938,In_4100);
or U7063 (N_7063,In_1633,In_4532);
nand U7064 (N_7064,In_3632,In_3478);
nor U7065 (N_7065,In_4492,In_3383);
nand U7066 (N_7066,In_1709,In_2106);
or U7067 (N_7067,In_854,In_3279);
nand U7068 (N_7068,In_4315,In_3385);
nand U7069 (N_7069,In_2972,In_2885);
or U7070 (N_7070,In_497,In_2084);
nor U7071 (N_7071,In_2870,In_2413);
and U7072 (N_7072,In_3903,In_1381);
nor U7073 (N_7073,In_1478,In_1736);
xor U7074 (N_7074,In_441,In_900);
nor U7075 (N_7075,In_1855,In_4701);
and U7076 (N_7076,In_2490,In_3885);
or U7077 (N_7077,In_223,In_689);
nand U7078 (N_7078,In_3091,In_1119);
nor U7079 (N_7079,In_85,In_3494);
nor U7080 (N_7080,In_3375,In_833);
nor U7081 (N_7081,In_1234,In_3573);
nand U7082 (N_7082,In_2837,In_4730);
nand U7083 (N_7083,In_2643,In_2870);
nor U7084 (N_7084,In_1783,In_2318);
xnor U7085 (N_7085,In_3006,In_1995);
nand U7086 (N_7086,In_3702,In_841);
or U7087 (N_7087,In_2476,In_397);
nand U7088 (N_7088,In_323,In_4254);
nor U7089 (N_7089,In_4429,In_1094);
nor U7090 (N_7090,In_2563,In_3001);
or U7091 (N_7091,In_4145,In_4148);
nor U7092 (N_7092,In_266,In_4430);
and U7093 (N_7093,In_4707,In_4449);
nand U7094 (N_7094,In_2863,In_1412);
nor U7095 (N_7095,In_2134,In_1603);
nor U7096 (N_7096,In_834,In_2843);
or U7097 (N_7097,In_179,In_2740);
nand U7098 (N_7098,In_4495,In_880);
xor U7099 (N_7099,In_2242,In_1569);
and U7100 (N_7100,In_2636,In_1382);
or U7101 (N_7101,In_3748,In_4280);
or U7102 (N_7102,In_1509,In_226);
nand U7103 (N_7103,In_4205,In_2959);
or U7104 (N_7104,In_1419,In_920);
and U7105 (N_7105,In_3124,In_4148);
xnor U7106 (N_7106,In_63,In_2524);
xor U7107 (N_7107,In_2036,In_1507);
nand U7108 (N_7108,In_3212,In_2020);
and U7109 (N_7109,In_3546,In_3613);
nor U7110 (N_7110,In_156,In_345);
nor U7111 (N_7111,In_1484,In_3985);
or U7112 (N_7112,In_4422,In_3372);
nor U7113 (N_7113,In_4465,In_2215);
or U7114 (N_7114,In_2192,In_116);
or U7115 (N_7115,In_1048,In_3157);
xnor U7116 (N_7116,In_4580,In_630);
xor U7117 (N_7117,In_631,In_4543);
nand U7118 (N_7118,In_3704,In_3822);
and U7119 (N_7119,In_4751,In_637);
and U7120 (N_7120,In_4286,In_3488);
xor U7121 (N_7121,In_4602,In_1019);
nor U7122 (N_7122,In_3041,In_3740);
and U7123 (N_7123,In_4653,In_583);
and U7124 (N_7124,In_4239,In_4363);
or U7125 (N_7125,In_880,In_4047);
nand U7126 (N_7126,In_1353,In_3631);
nor U7127 (N_7127,In_1589,In_1959);
xnor U7128 (N_7128,In_2078,In_4020);
or U7129 (N_7129,In_2176,In_2275);
and U7130 (N_7130,In_3134,In_675);
nor U7131 (N_7131,In_4092,In_4883);
and U7132 (N_7132,In_3826,In_418);
nand U7133 (N_7133,In_1445,In_362);
nor U7134 (N_7134,In_3556,In_4240);
nor U7135 (N_7135,In_96,In_4163);
and U7136 (N_7136,In_4456,In_1308);
nand U7137 (N_7137,In_3564,In_3318);
or U7138 (N_7138,In_1476,In_4421);
nand U7139 (N_7139,In_3641,In_2241);
and U7140 (N_7140,In_4598,In_4967);
xor U7141 (N_7141,In_4332,In_157);
nand U7142 (N_7142,In_1845,In_4679);
and U7143 (N_7143,In_375,In_3649);
nor U7144 (N_7144,In_2503,In_975);
nand U7145 (N_7145,In_4867,In_1462);
xnor U7146 (N_7146,In_4238,In_2214);
nand U7147 (N_7147,In_64,In_1447);
nand U7148 (N_7148,In_336,In_4403);
nor U7149 (N_7149,In_9,In_462);
xor U7150 (N_7150,In_583,In_4527);
xnor U7151 (N_7151,In_3310,In_457);
xor U7152 (N_7152,In_760,In_1723);
nor U7153 (N_7153,In_419,In_2207);
xor U7154 (N_7154,In_2120,In_1274);
nor U7155 (N_7155,In_4921,In_3344);
or U7156 (N_7156,In_3757,In_2055);
nand U7157 (N_7157,In_758,In_2490);
and U7158 (N_7158,In_2440,In_2724);
nor U7159 (N_7159,In_2325,In_4353);
nand U7160 (N_7160,In_2103,In_2149);
xnor U7161 (N_7161,In_286,In_145);
xnor U7162 (N_7162,In_3747,In_2345);
xnor U7163 (N_7163,In_3240,In_343);
or U7164 (N_7164,In_1337,In_2342);
and U7165 (N_7165,In_2689,In_4509);
xnor U7166 (N_7166,In_3512,In_154);
nand U7167 (N_7167,In_764,In_1693);
nor U7168 (N_7168,In_3148,In_4044);
or U7169 (N_7169,In_4463,In_3023);
nor U7170 (N_7170,In_2724,In_2533);
and U7171 (N_7171,In_1458,In_2472);
or U7172 (N_7172,In_1781,In_1331);
xor U7173 (N_7173,In_1570,In_1996);
or U7174 (N_7174,In_4646,In_4754);
nor U7175 (N_7175,In_3130,In_3479);
nand U7176 (N_7176,In_483,In_4633);
and U7177 (N_7177,In_1341,In_4937);
and U7178 (N_7178,In_4483,In_3164);
and U7179 (N_7179,In_3534,In_3812);
nand U7180 (N_7180,In_3182,In_1276);
nand U7181 (N_7181,In_2689,In_1802);
xnor U7182 (N_7182,In_356,In_4322);
and U7183 (N_7183,In_3677,In_747);
xnor U7184 (N_7184,In_1994,In_3349);
xor U7185 (N_7185,In_3946,In_1676);
nand U7186 (N_7186,In_4195,In_3557);
or U7187 (N_7187,In_3565,In_142);
or U7188 (N_7188,In_2509,In_4693);
nor U7189 (N_7189,In_4061,In_445);
or U7190 (N_7190,In_4949,In_2734);
nand U7191 (N_7191,In_648,In_4264);
xnor U7192 (N_7192,In_215,In_4194);
and U7193 (N_7193,In_2118,In_1671);
nor U7194 (N_7194,In_4878,In_3046);
xnor U7195 (N_7195,In_551,In_2853);
and U7196 (N_7196,In_146,In_432);
nor U7197 (N_7197,In_2741,In_2935);
or U7198 (N_7198,In_4905,In_2933);
or U7199 (N_7199,In_3489,In_2949);
and U7200 (N_7200,In_1569,In_2168);
nor U7201 (N_7201,In_4290,In_467);
nor U7202 (N_7202,In_4987,In_1179);
and U7203 (N_7203,In_2665,In_4465);
and U7204 (N_7204,In_4009,In_2551);
nand U7205 (N_7205,In_4601,In_1303);
nor U7206 (N_7206,In_3271,In_72);
and U7207 (N_7207,In_4201,In_4133);
nor U7208 (N_7208,In_33,In_4628);
nand U7209 (N_7209,In_883,In_4512);
or U7210 (N_7210,In_255,In_2026);
nand U7211 (N_7211,In_2930,In_4485);
nand U7212 (N_7212,In_440,In_4648);
nand U7213 (N_7213,In_1579,In_816);
nand U7214 (N_7214,In_1852,In_319);
or U7215 (N_7215,In_959,In_2140);
or U7216 (N_7216,In_4495,In_4127);
nand U7217 (N_7217,In_1109,In_4758);
nor U7218 (N_7218,In_41,In_2829);
nand U7219 (N_7219,In_4132,In_3599);
and U7220 (N_7220,In_39,In_4127);
nor U7221 (N_7221,In_635,In_4008);
xnor U7222 (N_7222,In_3985,In_4658);
xor U7223 (N_7223,In_4739,In_490);
nand U7224 (N_7224,In_1606,In_3097);
nand U7225 (N_7225,In_3931,In_687);
nand U7226 (N_7226,In_2851,In_351);
and U7227 (N_7227,In_2503,In_2461);
and U7228 (N_7228,In_957,In_3051);
or U7229 (N_7229,In_2113,In_2389);
and U7230 (N_7230,In_4554,In_3441);
xnor U7231 (N_7231,In_1459,In_1047);
or U7232 (N_7232,In_4621,In_3556);
or U7233 (N_7233,In_3848,In_3573);
nand U7234 (N_7234,In_896,In_4379);
xor U7235 (N_7235,In_1961,In_366);
and U7236 (N_7236,In_4860,In_1856);
xnor U7237 (N_7237,In_3589,In_2590);
nor U7238 (N_7238,In_1261,In_2304);
and U7239 (N_7239,In_4116,In_4743);
xnor U7240 (N_7240,In_1686,In_4722);
and U7241 (N_7241,In_2263,In_1576);
xor U7242 (N_7242,In_488,In_3533);
nor U7243 (N_7243,In_4134,In_3882);
or U7244 (N_7244,In_3430,In_480);
xor U7245 (N_7245,In_2565,In_3991);
and U7246 (N_7246,In_1094,In_2077);
or U7247 (N_7247,In_4807,In_1511);
nand U7248 (N_7248,In_4189,In_4807);
nand U7249 (N_7249,In_2590,In_1900);
nor U7250 (N_7250,In_4472,In_3790);
xnor U7251 (N_7251,In_3701,In_4523);
nor U7252 (N_7252,In_690,In_2881);
nand U7253 (N_7253,In_2716,In_4470);
nand U7254 (N_7254,In_105,In_1431);
and U7255 (N_7255,In_4744,In_4375);
nand U7256 (N_7256,In_1266,In_1993);
or U7257 (N_7257,In_3944,In_398);
nor U7258 (N_7258,In_816,In_431);
and U7259 (N_7259,In_3502,In_3459);
xor U7260 (N_7260,In_2371,In_3185);
or U7261 (N_7261,In_3499,In_2565);
or U7262 (N_7262,In_2729,In_914);
xnor U7263 (N_7263,In_2438,In_2487);
nand U7264 (N_7264,In_3662,In_4557);
nand U7265 (N_7265,In_3872,In_2460);
and U7266 (N_7266,In_1201,In_2465);
xor U7267 (N_7267,In_4166,In_1407);
xor U7268 (N_7268,In_2641,In_3446);
nand U7269 (N_7269,In_3067,In_4994);
xnor U7270 (N_7270,In_1049,In_4136);
xor U7271 (N_7271,In_1699,In_2816);
and U7272 (N_7272,In_4532,In_2974);
or U7273 (N_7273,In_699,In_2130);
and U7274 (N_7274,In_4868,In_4718);
xor U7275 (N_7275,In_1202,In_447);
nand U7276 (N_7276,In_2198,In_4741);
and U7277 (N_7277,In_856,In_4216);
and U7278 (N_7278,In_4348,In_4787);
xor U7279 (N_7279,In_4262,In_1478);
nand U7280 (N_7280,In_1030,In_3310);
or U7281 (N_7281,In_2009,In_318);
nand U7282 (N_7282,In_3824,In_368);
xor U7283 (N_7283,In_3033,In_2077);
nand U7284 (N_7284,In_4732,In_3011);
xnor U7285 (N_7285,In_696,In_796);
and U7286 (N_7286,In_2957,In_1892);
xnor U7287 (N_7287,In_2684,In_4163);
and U7288 (N_7288,In_2293,In_718);
or U7289 (N_7289,In_1187,In_3391);
nor U7290 (N_7290,In_2399,In_3847);
or U7291 (N_7291,In_1110,In_3900);
or U7292 (N_7292,In_3888,In_1971);
xor U7293 (N_7293,In_4801,In_4605);
or U7294 (N_7294,In_670,In_646);
and U7295 (N_7295,In_4060,In_4387);
and U7296 (N_7296,In_2744,In_3954);
nor U7297 (N_7297,In_4986,In_846);
nand U7298 (N_7298,In_3630,In_2647);
nand U7299 (N_7299,In_2507,In_2487);
nand U7300 (N_7300,In_1832,In_126);
nor U7301 (N_7301,In_702,In_1046);
nor U7302 (N_7302,In_4219,In_3222);
and U7303 (N_7303,In_4257,In_4669);
xor U7304 (N_7304,In_152,In_2522);
and U7305 (N_7305,In_4171,In_812);
nor U7306 (N_7306,In_2692,In_4765);
nand U7307 (N_7307,In_2966,In_2056);
nor U7308 (N_7308,In_3333,In_3782);
or U7309 (N_7309,In_1275,In_1164);
or U7310 (N_7310,In_1693,In_3694);
and U7311 (N_7311,In_3439,In_2660);
or U7312 (N_7312,In_1151,In_2566);
and U7313 (N_7313,In_2190,In_4279);
xor U7314 (N_7314,In_863,In_3816);
nor U7315 (N_7315,In_3617,In_4058);
or U7316 (N_7316,In_3919,In_1424);
or U7317 (N_7317,In_3772,In_3243);
nor U7318 (N_7318,In_1160,In_1206);
or U7319 (N_7319,In_2346,In_4068);
nand U7320 (N_7320,In_1343,In_352);
nand U7321 (N_7321,In_3317,In_975);
and U7322 (N_7322,In_3058,In_787);
xor U7323 (N_7323,In_802,In_2842);
and U7324 (N_7324,In_726,In_1201);
or U7325 (N_7325,In_2634,In_2881);
or U7326 (N_7326,In_1126,In_1501);
nor U7327 (N_7327,In_2426,In_2435);
and U7328 (N_7328,In_1611,In_862);
nand U7329 (N_7329,In_861,In_1248);
nand U7330 (N_7330,In_4780,In_966);
xor U7331 (N_7331,In_3362,In_3169);
and U7332 (N_7332,In_1745,In_2224);
nor U7333 (N_7333,In_395,In_187);
nor U7334 (N_7334,In_4285,In_2191);
nor U7335 (N_7335,In_2578,In_1157);
xnor U7336 (N_7336,In_2937,In_3354);
nand U7337 (N_7337,In_3751,In_3119);
nor U7338 (N_7338,In_4022,In_3919);
nor U7339 (N_7339,In_2907,In_1554);
and U7340 (N_7340,In_3136,In_1728);
nor U7341 (N_7341,In_999,In_4331);
and U7342 (N_7342,In_2590,In_4509);
nor U7343 (N_7343,In_3728,In_763);
xnor U7344 (N_7344,In_1235,In_962);
or U7345 (N_7345,In_2766,In_4469);
nor U7346 (N_7346,In_3566,In_1957);
xor U7347 (N_7347,In_1808,In_1960);
or U7348 (N_7348,In_662,In_4079);
nor U7349 (N_7349,In_4283,In_2926);
nand U7350 (N_7350,In_1043,In_2844);
or U7351 (N_7351,In_2576,In_998);
or U7352 (N_7352,In_1092,In_3845);
and U7353 (N_7353,In_1146,In_1138);
xnor U7354 (N_7354,In_1715,In_4264);
xor U7355 (N_7355,In_2338,In_4182);
xnor U7356 (N_7356,In_3947,In_4523);
nor U7357 (N_7357,In_3747,In_3250);
nor U7358 (N_7358,In_2515,In_2491);
nor U7359 (N_7359,In_1790,In_3);
nand U7360 (N_7360,In_1835,In_4053);
xnor U7361 (N_7361,In_48,In_2251);
nand U7362 (N_7362,In_4178,In_1819);
or U7363 (N_7363,In_1466,In_451);
and U7364 (N_7364,In_4473,In_4747);
xor U7365 (N_7365,In_1048,In_4001);
xnor U7366 (N_7366,In_755,In_2745);
xor U7367 (N_7367,In_374,In_4993);
nand U7368 (N_7368,In_4994,In_2972);
and U7369 (N_7369,In_3299,In_596);
nor U7370 (N_7370,In_4027,In_3485);
nor U7371 (N_7371,In_764,In_3888);
and U7372 (N_7372,In_4602,In_3752);
xor U7373 (N_7373,In_374,In_4092);
nor U7374 (N_7374,In_2993,In_239);
nand U7375 (N_7375,In_4144,In_366);
nor U7376 (N_7376,In_4479,In_3524);
nand U7377 (N_7377,In_385,In_428);
or U7378 (N_7378,In_2144,In_2713);
and U7379 (N_7379,In_1041,In_287);
nor U7380 (N_7380,In_2374,In_1654);
or U7381 (N_7381,In_1262,In_2981);
xnor U7382 (N_7382,In_3087,In_3654);
nand U7383 (N_7383,In_2476,In_1598);
xnor U7384 (N_7384,In_2037,In_642);
or U7385 (N_7385,In_4118,In_2995);
or U7386 (N_7386,In_2345,In_569);
or U7387 (N_7387,In_577,In_1854);
nand U7388 (N_7388,In_626,In_4746);
or U7389 (N_7389,In_1164,In_2382);
nand U7390 (N_7390,In_719,In_757);
nor U7391 (N_7391,In_3233,In_2021);
and U7392 (N_7392,In_4923,In_4184);
nor U7393 (N_7393,In_3977,In_1453);
xnor U7394 (N_7394,In_889,In_1997);
and U7395 (N_7395,In_1784,In_1190);
nor U7396 (N_7396,In_4967,In_3020);
nor U7397 (N_7397,In_1885,In_1148);
or U7398 (N_7398,In_1557,In_3788);
nand U7399 (N_7399,In_4061,In_3082);
nand U7400 (N_7400,In_313,In_2490);
nand U7401 (N_7401,In_2121,In_3882);
or U7402 (N_7402,In_885,In_3030);
nand U7403 (N_7403,In_150,In_3394);
nor U7404 (N_7404,In_1360,In_4860);
xnor U7405 (N_7405,In_2143,In_2440);
or U7406 (N_7406,In_4582,In_4697);
nor U7407 (N_7407,In_1720,In_3469);
xor U7408 (N_7408,In_1490,In_457);
or U7409 (N_7409,In_2537,In_3285);
and U7410 (N_7410,In_4184,In_2771);
xor U7411 (N_7411,In_1977,In_702);
or U7412 (N_7412,In_4294,In_2852);
or U7413 (N_7413,In_4286,In_2150);
and U7414 (N_7414,In_2773,In_283);
xnor U7415 (N_7415,In_838,In_1259);
xnor U7416 (N_7416,In_4090,In_974);
or U7417 (N_7417,In_3797,In_2046);
or U7418 (N_7418,In_2246,In_1890);
nor U7419 (N_7419,In_1404,In_1261);
nand U7420 (N_7420,In_4120,In_2875);
xnor U7421 (N_7421,In_1201,In_1108);
or U7422 (N_7422,In_4111,In_3854);
nand U7423 (N_7423,In_1287,In_614);
xor U7424 (N_7424,In_56,In_3712);
and U7425 (N_7425,In_4701,In_3805);
nand U7426 (N_7426,In_3004,In_3594);
nor U7427 (N_7427,In_2456,In_4833);
nand U7428 (N_7428,In_3155,In_2238);
nor U7429 (N_7429,In_4587,In_547);
or U7430 (N_7430,In_4152,In_2931);
nand U7431 (N_7431,In_3468,In_1787);
xnor U7432 (N_7432,In_140,In_364);
or U7433 (N_7433,In_4405,In_2227);
nor U7434 (N_7434,In_2387,In_2533);
xnor U7435 (N_7435,In_4146,In_1191);
and U7436 (N_7436,In_3732,In_2298);
nor U7437 (N_7437,In_4550,In_470);
or U7438 (N_7438,In_4960,In_2254);
xnor U7439 (N_7439,In_286,In_1108);
nand U7440 (N_7440,In_18,In_2731);
nand U7441 (N_7441,In_3378,In_3476);
nor U7442 (N_7442,In_3681,In_1857);
xor U7443 (N_7443,In_1545,In_4512);
or U7444 (N_7444,In_353,In_3718);
nor U7445 (N_7445,In_1616,In_3913);
and U7446 (N_7446,In_2667,In_3920);
nor U7447 (N_7447,In_4052,In_1663);
or U7448 (N_7448,In_4186,In_4048);
xnor U7449 (N_7449,In_1048,In_319);
or U7450 (N_7450,In_856,In_1596);
and U7451 (N_7451,In_1898,In_4818);
or U7452 (N_7452,In_1554,In_2313);
nor U7453 (N_7453,In_3830,In_1010);
xor U7454 (N_7454,In_3978,In_4465);
xor U7455 (N_7455,In_644,In_664);
nor U7456 (N_7456,In_341,In_1850);
and U7457 (N_7457,In_750,In_177);
xor U7458 (N_7458,In_4844,In_4435);
nand U7459 (N_7459,In_4336,In_2514);
nand U7460 (N_7460,In_3452,In_1430);
and U7461 (N_7461,In_1464,In_2404);
xor U7462 (N_7462,In_602,In_3167);
nor U7463 (N_7463,In_2734,In_4410);
xnor U7464 (N_7464,In_2503,In_3607);
nand U7465 (N_7465,In_4364,In_1432);
nand U7466 (N_7466,In_1303,In_4002);
nor U7467 (N_7467,In_3174,In_2788);
and U7468 (N_7468,In_1240,In_4456);
nor U7469 (N_7469,In_1816,In_1660);
nand U7470 (N_7470,In_4331,In_3605);
nand U7471 (N_7471,In_492,In_1341);
or U7472 (N_7472,In_2651,In_4809);
nor U7473 (N_7473,In_3581,In_4966);
nor U7474 (N_7474,In_3981,In_4896);
nand U7475 (N_7475,In_2625,In_1656);
and U7476 (N_7476,In_1845,In_1592);
xor U7477 (N_7477,In_3762,In_639);
and U7478 (N_7478,In_538,In_1692);
or U7479 (N_7479,In_2457,In_4120);
xnor U7480 (N_7480,In_4628,In_2374);
and U7481 (N_7481,In_733,In_713);
and U7482 (N_7482,In_4831,In_149);
and U7483 (N_7483,In_3443,In_1087);
and U7484 (N_7484,In_2331,In_4372);
or U7485 (N_7485,In_1456,In_2998);
xor U7486 (N_7486,In_3333,In_4702);
xor U7487 (N_7487,In_4341,In_2678);
xnor U7488 (N_7488,In_3417,In_988);
nor U7489 (N_7489,In_2006,In_1377);
or U7490 (N_7490,In_1375,In_4470);
and U7491 (N_7491,In_3619,In_4126);
xnor U7492 (N_7492,In_4758,In_3285);
or U7493 (N_7493,In_2066,In_2579);
and U7494 (N_7494,In_387,In_4826);
nor U7495 (N_7495,In_2918,In_862);
xor U7496 (N_7496,In_1282,In_2614);
and U7497 (N_7497,In_3732,In_1527);
nor U7498 (N_7498,In_2953,In_1222);
and U7499 (N_7499,In_1725,In_3184);
nand U7500 (N_7500,In_4158,In_4204);
nor U7501 (N_7501,In_2319,In_4608);
or U7502 (N_7502,In_3448,In_4726);
xor U7503 (N_7503,In_2034,In_1974);
and U7504 (N_7504,In_4424,In_1582);
nor U7505 (N_7505,In_4700,In_2156);
xor U7506 (N_7506,In_2649,In_3593);
or U7507 (N_7507,In_4203,In_2469);
nor U7508 (N_7508,In_3875,In_2147);
xor U7509 (N_7509,In_3230,In_2119);
and U7510 (N_7510,In_1806,In_326);
xnor U7511 (N_7511,In_2243,In_766);
nor U7512 (N_7512,In_703,In_1077);
xor U7513 (N_7513,In_3228,In_392);
or U7514 (N_7514,In_570,In_3920);
and U7515 (N_7515,In_2846,In_4836);
nand U7516 (N_7516,In_2734,In_4167);
xnor U7517 (N_7517,In_1068,In_3820);
and U7518 (N_7518,In_4777,In_1170);
and U7519 (N_7519,In_330,In_3160);
xor U7520 (N_7520,In_2351,In_1228);
nor U7521 (N_7521,In_3802,In_4966);
or U7522 (N_7522,In_1336,In_29);
xor U7523 (N_7523,In_1945,In_4573);
nand U7524 (N_7524,In_4126,In_4973);
nand U7525 (N_7525,In_3579,In_3305);
and U7526 (N_7526,In_2691,In_2800);
nand U7527 (N_7527,In_3544,In_556);
or U7528 (N_7528,In_995,In_1751);
nor U7529 (N_7529,In_415,In_1365);
nand U7530 (N_7530,In_1311,In_1932);
nand U7531 (N_7531,In_0,In_3939);
nor U7532 (N_7532,In_4820,In_4973);
nand U7533 (N_7533,In_788,In_584);
and U7534 (N_7534,In_3235,In_1965);
and U7535 (N_7535,In_421,In_325);
nand U7536 (N_7536,In_2525,In_4355);
or U7537 (N_7537,In_1957,In_3560);
xnor U7538 (N_7538,In_4545,In_3947);
xnor U7539 (N_7539,In_4958,In_3270);
nor U7540 (N_7540,In_3110,In_1018);
or U7541 (N_7541,In_2859,In_2825);
or U7542 (N_7542,In_1057,In_4552);
and U7543 (N_7543,In_1614,In_1796);
or U7544 (N_7544,In_4264,In_4641);
and U7545 (N_7545,In_135,In_2525);
xor U7546 (N_7546,In_2422,In_2678);
or U7547 (N_7547,In_4116,In_4353);
xnor U7548 (N_7548,In_3411,In_4188);
xnor U7549 (N_7549,In_4722,In_313);
and U7550 (N_7550,In_2598,In_335);
or U7551 (N_7551,In_2757,In_1746);
or U7552 (N_7552,In_3881,In_560);
nor U7553 (N_7553,In_831,In_3728);
xor U7554 (N_7554,In_3214,In_1303);
nor U7555 (N_7555,In_4610,In_3301);
nor U7556 (N_7556,In_301,In_2792);
nand U7557 (N_7557,In_4540,In_3587);
or U7558 (N_7558,In_4220,In_1037);
nor U7559 (N_7559,In_4181,In_4267);
nor U7560 (N_7560,In_2166,In_4700);
nand U7561 (N_7561,In_4033,In_88);
xnor U7562 (N_7562,In_1831,In_3769);
or U7563 (N_7563,In_3704,In_3459);
or U7564 (N_7564,In_1095,In_3628);
nor U7565 (N_7565,In_1670,In_200);
or U7566 (N_7566,In_2765,In_1201);
nand U7567 (N_7567,In_385,In_760);
xor U7568 (N_7568,In_1692,In_287);
xor U7569 (N_7569,In_2307,In_1852);
and U7570 (N_7570,In_1852,In_2644);
nand U7571 (N_7571,In_4459,In_3245);
nand U7572 (N_7572,In_2556,In_982);
or U7573 (N_7573,In_2558,In_342);
nand U7574 (N_7574,In_3776,In_1467);
xnor U7575 (N_7575,In_3138,In_818);
or U7576 (N_7576,In_880,In_865);
nor U7577 (N_7577,In_4283,In_4735);
and U7578 (N_7578,In_4243,In_2775);
xnor U7579 (N_7579,In_3813,In_3571);
and U7580 (N_7580,In_1861,In_1255);
and U7581 (N_7581,In_915,In_315);
nor U7582 (N_7582,In_3407,In_4442);
or U7583 (N_7583,In_2339,In_3169);
and U7584 (N_7584,In_4264,In_2083);
or U7585 (N_7585,In_2167,In_2154);
nor U7586 (N_7586,In_1568,In_16);
xor U7587 (N_7587,In_1257,In_2902);
and U7588 (N_7588,In_339,In_520);
xor U7589 (N_7589,In_4911,In_890);
nor U7590 (N_7590,In_1969,In_4649);
nand U7591 (N_7591,In_3926,In_2173);
nand U7592 (N_7592,In_3182,In_3396);
nor U7593 (N_7593,In_298,In_2266);
and U7594 (N_7594,In_2152,In_1571);
nand U7595 (N_7595,In_3888,In_1164);
nor U7596 (N_7596,In_4945,In_2446);
or U7597 (N_7597,In_3841,In_498);
and U7598 (N_7598,In_990,In_2809);
xor U7599 (N_7599,In_993,In_4430);
nor U7600 (N_7600,In_2181,In_3546);
or U7601 (N_7601,In_1739,In_2085);
and U7602 (N_7602,In_938,In_2113);
nand U7603 (N_7603,In_2719,In_3557);
nor U7604 (N_7604,In_915,In_636);
nor U7605 (N_7605,In_2953,In_209);
and U7606 (N_7606,In_2134,In_546);
xor U7607 (N_7607,In_742,In_2858);
xnor U7608 (N_7608,In_3485,In_4135);
xor U7609 (N_7609,In_1252,In_2589);
and U7610 (N_7610,In_1349,In_1184);
nand U7611 (N_7611,In_3628,In_3200);
and U7612 (N_7612,In_2338,In_1419);
nor U7613 (N_7613,In_3781,In_1130);
nor U7614 (N_7614,In_164,In_2604);
and U7615 (N_7615,In_4190,In_2219);
xnor U7616 (N_7616,In_335,In_1568);
nand U7617 (N_7617,In_2435,In_2702);
nor U7618 (N_7618,In_1719,In_2711);
and U7619 (N_7619,In_4707,In_1054);
or U7620 (N_7620,In_4058,In_3713);
nor U7621 (N_7621,In_3008,In_2844);
and U7622 (N_7622,In_4674,In_503);
or U7623 (N_7623,In_1758,In_4436);
xor U7624 (N_7624,In_288,In_2179);
xnor U7625 (N_7625,In_2160,In_2066);
xor U7626 (N_7626,In_2626,In_4443);
or U7627 (N_7627,In_4900,In_1840);
xnor U7628 (N_7628,In_1105,In_729);
nor U7629 (N_7629,In_871,In_2397);
and U7630 (N_7630,In_3239,In_1404);
nor U7631 (N_7631,In_329,In_3988);
nor U7632 (N_7632,In_1014,In_366);
nor U7633 (N_7633,In_2726,In_373);
nand U7634 (N_7634,In_4522,In_1864);
nor U7635 (N_7635,In_3259,In_3861);
and U7636 (N_7636,In_732,In_2754);
nor U7637 (N_7637,In_2252,In_2149);
or U7638 (N_7638,In_2290,In_4235);
or U7639 (N_7639,In_2358,In_1504);
nor U7640 (N_7640,In_4192,In_3794);
or U7641 (N_7641,In_2875,In_346);
nor U7642 (N_7642,In_3711,In_583);
xnor U7643 (N_7643,In_3431,In_2327);
xnor U7644 (N_7644,In_1735,In_1043);
nor U7645 (N_7645,In_86,In_1096);
xnor U7646 (N_7646,In_624,In_822);
nand U7647 (N_7647,In_1769,In_1168);
and U7648 (N_7648,In_798,In_3207);
nand U7649 (N_7649,In_15,In_2018);
nor U7650 (N_7650,In_4783,In_2478);
xor U7651 (N_7651,In_1375,In_4521);
and U7652 (N_7652,In_2504,In_3647);
nor U7653 (N_7653,In_4346,In_237);
or U7654 (N_7654,In_2808,In_2228);
and U7655 (N_7655,In_2013,In_4405);
or U7656 (N_7656,In_2945,In_4014);
xnor U7657 (N_7657,In_727,In_2805);
nand U7658 (N_7658,In_604,In_3703);
nand U7659 (N_7659,In_1055,In_604);
xnor U7660 (N_7660,In_879,In_270);
or U7661 (N_7661,In_1540,In_4296);
xor U7662 (N_7662,In_1071,In_1867);
or U7663 (N_7663,In_1150,In_4253);
xnor U7664 (N_7664,In_3540,In_3920);
nor U7665 (N_7665,In_642,In_4056);
xnor U7666 (N_7666,In_4504,In_3118);
or U7667 (N_7667,In_3234,In_4301);
xnor U7668 (N_7668,In_1589,In_4837);
and U7669 (N_7669,In_600,In_2293);
nor U7670 (N_7670,In_761,In_1515);
xnor U7671 (N_7671,In_3365,In_558);
nand U7672 (N_7672,In_3503,In_4167);
xor U7673 (N_7673,In_4262,In_4580);
and U7674 (N_7674,In_2148,In_2521);
xnor U7675 (N_7675,In_2878,In_882);
and U7676 (N_7676,In_182,In_352);
or U7677 (N_7677,In_3047,In_2948);
xor U7678 (N_7678,In_383,In_1629);
nor U7679 (N_7679,In_338,In_3544);
xnor U7680 (N_7680,In_535,In_901);
nand U7681 (N_7681,In_2167,In_2738);
or U7682 (N_7682,In_1551,In_2337);
xnor U7683 (N_7683,In_4409,In_3958);
and U7684 (N_7684,In_1054,In_3408);
xnor U7685 (N_7685,In_3297,In_213);
nand U7686 (N_7686,In_1973,In_1526);
nor U7687 (N_7687,In_160,In_1518);
nand U7688 (N_7688,In_4557,In_2272);
and U7689 (N_7689,In_1574,In_3247);
nand U7690 (N_7690,In_4078,In_427);
nor U7691 (N_7691,In_168,In_4082);
nor U7692 (N_7692,In_1275,In_325);
nand U7693 (N_7693,In_784,In_4780);
xor U7694 (N_7694,In_2180,In_3028);
nor U7695 (N_7695,In_750,In_4060);
and U7696 (N_7696,In_109,In_3637);
xor U7697 (N_7697,In_908,In_2211);
and U7698 (N_7698,In_3296,In_4984);
nor U7699 (N_7699,In_3347,In_1782);
nand U7700 (N_7700,In_209,In_3737);
and U7701 (N_7701,In_637,In_2764);
or U7702 (N_7702,In_2985,In_1286);
or U7703 (N_7703,In_4696,In_1190);
or U7704 (N_7704,In_4956,In_2526);
nor U7705 (N_7705,In_560,In_917);
xnor U7706 (N_7706,In_4111,In_1421);
nor U7707 (N_7707,In_4546,In_306);
and U7708 (N_7708,In_1504,In_2869);
or U7709 (N_7709,In_3579,In_1580);
nor U7710 (N_7710,In_183,In_4750);
xor U7711 (N_7711,In_786,In_2739);
or U7712 (N_7712,In_3435,In_812);
xor U7713 (N_7713,In_4748,In_2085);
nand U7714 (N_7714,In_4364,In_4547);
or U7715 (N_7715,In_2339,In_3725);
nand U7716 (N_7716,In_2648,In_3570);
nor U7717 (N_7717,In_138,In_1444);
or U7718 (N_7718,In_2032,In_1656);
nor U7719 (N_7719,In_4006,In_4336);
nor U7720 (N_7720,In_4225,In_3041);
nand U7721 (N_7721,In_4603,In_225);
and U7722 (N_7722,In_4762,In_3876);
and U7723 (N_7723,In_3339,In_2869);
nor U7724 (N_7724,In_439,In_2071);
nand U7725 (N_7725,In_0,In_1159);
nand U7726 (N_7726,In_2650,In_4795);
or U7727 (N_7727,In_694,In_2897);
and U7728 (N_7728,In_4870,In_4346);
or U7729 (N_7729,In_4198,In_1152);
nor U7730 (N_7730,In_4365,In_2822);
and U7731 (N_7731,In_3447,In_1361);
and U7732 (N_7732,In_1941,In_4370);
nor U7733 (N_7733,In_355,In_3694);
nor U7734 (N_7734,In_4856,In_4621);
nor U7735 (N_7735,In_957,In_66);
nor U7736 (N_7736,In_548,In_413);
xnor U7737 (N_7737,In_1294,In_1765);
nand U7738 (N_7738,In_2958,In_4386);
nor U7739 (N_7739,In_2669,In_388);
nor U7740 (N_7740,In_4690,In_2989);
nand U7741 (N_7741,In_376,In_2575);
and U7742 (N_7742,In_3178,In_2735);
nor U7743 (N_7743,In_1658,In_1426);
nand U7744 (N_7744,In_841,In_1074);
nor U7745 (N_7745,In_48,In_2476);
xnor U7746 (N_7746,In_1200,In_1675);
nand U7747 (N_7747,In_3145,In_3975);
nor U7748 (N_7748,In_2873,In_301);
nor U7749 (N_7749,In_2752,In_2108);
or U7750 (N_7750,In_2177,In_4179);
nand U7751 (N_7751,In_3509,In_4434);
xor U7752 (N_7752,In_2409,In_3897);
xnor U7753 (N_7753,In_774,In_3565);
xnor U7754 (N_7754,In_1170,In_4922);
xor U7755 (N_7755,In_2833,In_2844);
nand U7756 (N_7756,In_4097,In_345);
nor U7757 (N_7757,In_2455,In_2366);
nor U7758 (N_7758,In_4744,In_3513);
nand U7759 (N_7759,In_4679,In_3321);
or U7760 (N_7760,In_2298,In_3035);
nor U7761 (N_7761,In_849,In_4892);
or U7762 (N_7762,In_1445,In_4254);
and U7763 (N_7763,In_2879,In_2335);
and U7764 (N_7764,In_2540,In_154);
nand U7765 (N_7765,In_4282,In_3628);
nand U7766 (N_7766,In_2350,In_3600);
nor U7767 (N_7767,In_3124,In_518);
or U7768 (N_7768,In_1203,In_1535);
or U7769 (N_7769,In_722,In_3365);
and U7770 (N_7770,In_3120,In_3741);
and U7771 (N_7771,In_4339,In_1814);
nand U7772 (N_7772,In_492,In_4087);
or U7773 (N_7773,In_2671,In_2073);
xnor U7774 (N_7774,In_4355,In_3204);
and U7775 (N_7775,In_1920,In_4573);
xor U7776 (N_7776,In_4279,In_523);
nor U7777 (N_7777,In_1957,In_3307);
nor U7778 (N_7778,In_1754,In_4620);
or U7779 (N_7779,In_2750,In_166);
xnor U7780 (N_7780,In_1729,In_3380);
or U7781 (N_7781,In_4031,In_3776);
nor U7782 (N_7782,In_3328,In_3772);
and U7783 (N_7783,In_1968,In_3301);
and U7784 (N_7784,In_680,In_2427);
and U7785 (N_7785,In_2848,In_4007);
nand U7786 (N_7786,In_4168,In_1245);
xor U7787 (N_7787,In_4127,In_2147);
or U7788 (N_7788,In_2086,In_2266);
nor U7789 (N_7789,In_1583,In_2615);
or U7790 (N_7790,In_2450,In_444);
nand U7791 (N_7791,In_3226,In_2859);
or U7792 (N_7792,In_716,In_459);
nor U7793 (N_7793,In_199,In_1859);
nand U7794 (N_7794,In_4105,In_57);
or U7795 (N_7795,In_4818,In_3269);
nor U7796 (N_7796,In_1391,In_2177);
or U7797 (N_7797,In_1266,In_1541);
nor U7798 (N_7798,In_1422,In_4894);
and U7799 (N_7799,In_322,In_1504);
or U7800 (N_7800,In_2824,In_43);
nand U7801 (N_7801,In_3930,In_4574);
and U7802 (N_7802,In_2152,In_3880);
nor U7803 (N_7803,In_4545,In_910);
nor U7804 (N_7804,In_2078,In_1786);
nand U7805 (N_7805,In_1824,In_843);
nor U7806 (N_7806,In_542,In_1164);
nand U7807 (N_7807,In_3875,In_4849);
nor U7808 (N_7808,In_3926,In_1223);
nand U7809 (N_7809,In_414,In_2543);
nand U7810 (N_7810,In_2658,In_4715);
and U7811 (N_7811,In_4907,In_2020);
or U7812 (N_7812,In_2758,In_3094);
or U7813 (N_7813,In_3302,In_1649);
and U7814 (N_7814,In_2032,In_2316);
xnor U7815 (N_7815,In_2797,In_1157);
nand U7816 (N_7816,In_2611,In_2101);
nand U7817 (N_7817,In_4141,In_997);
xnor U7818 (N_7818,In_1909,In_3146);
nor U7819 (N_7819,In_2936,In_1840);
nor U7820 (N_7820,In_2627,In_283);
xnor U7821 (N_7821,In_2303,In_4133);
nand U7822 (N_7822,In_2009,In_4957);
xnor U7823 (N_7823,In_4155,In_767);
xor U7824 (N_7824,In_4620,In_4605);
xnor U7825 (N_7825,In_2957,In_835);
or U7826 (N_7826,In_1562,In_3659);
or U7827 (N_7827,In_4984,In_2441);
or U7828 (N_7828,In_4302,In_3434);
xnor U7829 (N_7829,In_4201,In_1361);
nand U7830 (N_7830,In_4651,In_955);
and U7831 (N_7831,In_3673,In_3542);
xnor U7832 (N_7832,In_4802,In_3090);
nor U7833 (N_7833,In_1420,In_296);
nor U7834 (N_7834,In_2208,In_1341);
or U7835 (N_7835,In_2733,In_2564);
xnor U7836 (N_7836,In_592,In_1728);
or U7837 (N_7837,In_2154,In_3409);
nand U7838 (N_7838,In_2147,In_320);
and U7839 (N_7839,In_1489,In_4448);
xnor U7840 (N_7840,In_2991,In_294);
nor U7841 (N_7841,In_2753,In_520);
nand U7842 (N_7842,In_4334,In_1113);
or U7843 (N_7843,In_4644,In_3299);
and U7844 (N_7844,In_1411,In_3108);
nor U7845 (N_7845,In_4915,In_4101);
and U7846 (N_7846,In_82,In_217);
and U7847 (N_7847,In_2016,In_1101);
nor U7848 (N_7848,In_1329,In_2173);
xnor U7849 (N_7849,In_4417,In_1228);
or U7850 (N_7850,In_1672,In_373);
and U7851 (N_7851,In_1633,In_3821);
nor U7852 (N_7852,In_4192,In_2902);
and U7853 (N_7853,In_3731,In_708);
or U7854 (N_7854,In_3948,In_3270);
and U7855 (N_7855,In_3384,In_1975);
nand U7856 (N_7856,In_2668,In_2434);
nand U7857 (N_7857,In_2037,In_1003);
nand U7858 (N_7858,In_3006,In_1957);
nor U7859 (N_7859,In_3204,In_3415);
nand U7860 (N_7860,In_4346,In_815);
nor U7861 (N_7861,In_1589,In_431);
nor U7862 (N_7862,In_2396,In_3770);
xnor U7863 (N_7863,In_884,In_1921);
nand U7864 (N_7864,In_683,In_597);
and U7865 (N_7865,In_2945,In_3463);
or U7866 (N_7866,In_2416,In_4814);
or U7867 (N_7867,In_3745,In_1588);
or U7868 (N_7868,In_3802,In_4695);
and U7869 (N_7869,In_2292,In_3867);
xnor U7870 (N_7870,In_2274,In_4265);
xnor U7871 (N_7871,In_2056,In_1592);
nand U7872 (N_7872,In_1730,In_1426);
or U7873 (N_7873,In_813,In_676);
xor U7874 (N_7874,In_911,In_1737);
or U7875 (N_7875,In_1554,In_2497);
or U7876 (N_7876,In_1795,In_3680);
and U7877 (N_7877,In_3530,In_1946);
nand U7878 (N_7878,In_1602,In_3445);
or U7879 (N_7879,In_499,In_3542);
nor U7880 (N_7880,In_307,In_3168);
or U7881 (N_7881,In_3041,In_2974);
or U7882 (N_7882,In_859,In_2838);
xnor U7883 (N_7883,In_2077,In_1938);
nand U7884 (N_7884,In_4808,In_73);
and U7885 (N_7885,In_4000,In_1098);
nand U7886 (N_7886,In_3196,In_3940);
xnor U7887 (N_7887,In_2130,In_3344);
nand U7888 (N_7888,In_2024,In_2068);
nand U7889 (N_7889,In_1822,In_975);
xor U7890 (N_7890,In_4629,In_2721);
or U7891 (N_7891,In_4592,In_1895);
and U7892 (N_7892,In_515,In_3473);
xnor U7893 (N_7893,In_1296,In_3085);
or U7894 (N_7894,In_224,In_2580);
xnor U7895 (N_7895,In_4561,In_681);
nor U7896 (N_7896,In_3693,In_1923);
and U7897 (N_7897,In_2095,In_2470);
nor U7898 (N_7898,In_786,In_1129);
or U7899 (N_7899,In_1962,In_1833);
or U7900 (N_7900,In_291,In_3720);
nand U7901 (N_7901,In_1605,In_4993);
nand U7902 (N_7902,In_2277,In_2346);
or U7903 (N_7903,In_476,In_3074);
nor U7904 (N_7904,In_1039,In_1854);
nor U7905 (N_7905,In_2106,In_2733);
nand U7906 (N_7906,In_1760,In_2915);
or U7907 (N_7907,In_2143,In_1755);
and U7908 (N_7908,In_3622,In_61);
xor U7909 (N_7909,In_3563,In_3695);
xor U7910 (N_7910,In_2942,In_3035);
xnor U7911 (N_7911,In_547,In_1619);
nand U7912 (N_7912,In_19,In_2523);
xnor U7913 (N_7913,In_3511,In_2049);
xor U7914 (N_7914,In_2971,In_2705);
or U7915 (N_7915,In_3788,In_2728);
and U7916 (N_7916,In_3642,In_1503);
or U7917 (N_7917,In_2690,In_859);
nor U7918 (N_7918,In_774,In_4339);
nand U7919 (N_7919,In_3909,In_3592);
xor U7920 (N_7920,In_2966,In_2223);
and U7921 (N_7921,In_1082,In_3757);
nor U7922 (N_7922,In_4003,In_4787);
nor U7923 (N_7923,In_4061,In_3904);
or U7924 (N_7924,In_3205,In_4898);
and U7925 (N_7925,In_2481,In_2005);
or U7926 (N_7926,In_153,In_3428);
and U7927 (N_7927,In_4888,In_4166);
and U7928 (N_7928,In_773,In_1790);
nand U7929 (N_7929,In_93,In_2254);
nand U7930 (N_7930,In_4288,In_875);
and U7931 (N_7931,In_1941,In_2168);
nor U7932 (N_7932,In_4495,In_2717);
or U7933 (N_7933,In_3409,In_1097);
nand U7934 (N_7934,In_228,In_1602);
nand U7935 (N_7935,In_2672,In_1060);
nand U7936 (N_7936,In_4988,In_2654);
xor U7937 (N_7937,In_1085,In_2229);
nand U7938 (N_7938,In_2941,In_2935);
xor U7939 (N_7939,In_844,In_2956);
and U7940 (N_7940,In_3341,In_2867);
or U7941 (N_7941,In_4556,In_4930);
nand U7942 (N_7942,In_4490,In_590);
xnor U7943 (N_7943,In_2634,In_2465);
nor U7944 (N_7944,In_847,In_1870);
or U7945 (N_7945,In_2557,In_2981);
or U7946 (N_7946,In_3858,In_1271);
or U7947 (N_7947,In_540,In_3172);
nor U7948 (N_7948,In_1631,In_781);
xor U7949 (N_7949,In_2480,In_1443);
nand U7950 (N_7950,In_4501,In_2093);
xor U7951 (N_7951,In_271,In_3201);
nor U7952 (N_7952,In_349,In_4651);
xnor U7953 (N_7953,In_3581,In_1917);
xnor U7954 (N_7954,In_4135,In_1389);
or U7955 (N_7955,In_1878,In_754);
xnor U7956 (N_7956,In_4623,In_1728);
nand U7957 (N_7957,In_3130,In_426);
xnor U7958 (N_7958,In_1166,In_3435);
or U7959 (N_7959,In_1000,In_503);
xnor U7960 (N_7960,In_4369,In_948);
nor U7961 (N_7961,In_3920,In_3120);
and U7962 (N_7962,In_3765,In_727);
nor U7963 (N_7963,In_1592,In_3777);
xnor U7964 (N_7964,In_1917,In_3983);
xor U7965 (N_7965,In_3423,In_4673);
or U7966 (N_7966,In_3169,In_4479);
and U7967 (N_7967,In_1670,In_1974);
nand U7968 (N_7968,In_2311,In_1224);
nor U7969 (N_7969,In_1878,In_1609);
xor U7970 (N_7970,In_6,In_1817);
or U7971 (N_7971,In_2875,In_2907);
nor U7972 (N_7972,In_2476,In_1511);
nor U7973 (N_7973,In_874,In_790);
or U7974 (N_7974,In_1337,In_1797);
nand U7975 (N_7975,In_3171,In_234);
and U7976 (N_7976,In_3371,In_1590);
nor U7977 (N_7977,In_3010,In_4342);
xor U7978 (N_7978,In_3792,In_3697);
nor U7979 (N_7979,In_3939,In_1182);
nor U7980 (N_7980,In_1487,In_2750);
or U7981 (N_7981,In_3001,In_842);
or U7982 (N_7982,In_3951,In_385);
and U7983 (N_7983,In_4943,In_2085);
and U7984 (N_7984,In_3894,In_3582);
and U7985 (N_7985,In_4547,In_1439);
xor U7986 (N_7986,In_4567,In_1962);
and U7987 (N_7987,In_701,In_285);
and U7988 (N_7988,In_3278,In_2108);
or U7989 (N_7989,In_3274,In_544);
or U7990 (N_7990,In_1224,In_1305);
xnor U7991 (N_7991,In_4588,In_4445);
nor U7992 (N_7992,In_2197,In_1180);
nor U7993 (N_7993,In_1609,In_2768);
and U7994 (N_7994,In_2466,In_845);
xnor U7995 (N_7995,In_1109,In_1232);
nand U7996 (N_7996,In_3994,In_2612);
nor U7997 (N_7997,In_1935,In_4803);
or U7998 (N_7998,In_1050,In_4520);
and U7999 (N_7999,In_975,In_3115);
and U8000 (N_8000,In_249,In_1023);
and U8001 (N_8001,In_1851,In_1365);
xor U8002 (N_8002,In_96,In_4110);
or U8003 (N_8003,In_2456,In_2489);
and U8004 (N_8004,In_235,In_139);
nand U8005 (N_8005,In_4343,In_3614);
or U8006 (N_8006,In_3699,In_1250);
xnor U8007 (N_8007,In_4713,In_493);
xor U8008 (N_8008,In_1079,In_4948);
nand U8009 (N_8009,In_1728,In_506);
or U8010 (N_8010,In_103,In_3401);
nor U8011 (N_8011,In_2581,In_4997);
or U8012 (N_8012,In_1927,In_1984);
and U8013 (N_8013,In_3749,In_4540);
and U8014 (N_8014,In_2762,In_1781);
or U8015 (N_8015,In_4393,In_3326);
or U8016 (N_8016,In_3457,In_4435);
nor U8017 (N_8017,In_3497,In_3259);
nand U8018 (N_8018,In_131,In_612);
or U8019 (N_8019,In_2172,In_4383);
or U8020 (N_8020,In_1263,In_1963);
xor U8021 (N_8021,In_2498,In_1123);
and U8022 (N_8022,In_2381,In_305);
and U8023 (N_8023,In_3282,In_4391);
and U8024 (N_8024,In_4867,In_264);
nor U8025 (N_8025,In_4666,In_2066);
and U8026 (N_8026,In_1985,In_1475);
nor U8027 (N_8027,In_4718,In_2146);
or U8028 (N_8028,In_2843,In_39);
and U8029 (N_8029,In_4075,In_2527);
or U8030 (N_8030,In_632,In_26);
and U8031 (N_8031,In_2645,In_4598);
nand U8032 (N_8032,In_2149,In_2964);
xnor U8033 (N_8033,In_1034,In_1372);
or U8034 (N_8034,In_1710,In_4269);
and U8035 (N_8035,In_3594,In_3010);
and U8036 (N_8036,In_4847,In_3378);
or U8037 (N_8037,In_3588,In_3098);
or U8038 (N_8038,In_2336,In_4314);
nor U8039 (N_8039,In_349,In_4099);
xor U8040 (N_8040,In_3385,In_3824);
nor U8041 (N_8041,In_4123,In_2057);
nand U8042 (N_8042,In_670,In_3260);
nor U8043 (N_8043,In_3920,In_4142);
and U8044 (N_8044,In_1312,In_2963);
xnor U8045 (N_8045,In_969,In_1735);
xnor U8046 (N_8046,In_603,In_3833);
or U8047 (N_8047,In_4698,In_2082);
nor U8048 (N_8048,In_217,In_2783);
xor U8049 (N_8049,In_3564,In_2611);
or U8050 (N_8050,In_2408,In_4812);
nand U8051 (N_8051,In_1626,In_3474);
or U8052 (N_8052,In_1930,In_383);
xnor U8053 (N_8053,In_4731,In_82);
nand U8054 (N_8054,In_1574,In_2741);
or U8055 (N_8055,In_2701,In_1023);
nand U8056 (N_8056,In_4313,In_2256);
and U8057 (N_8057,In_862,In_2137);
nand U8058 (N_8058,In_4372,In_3677);
nand U8059 (N_8059,In_3549,In_2510);
xnor U8060 (N_8060,In_3501,In_3986);
nand U8061 (N_8061,In_1717,In_4401);
and U8062 (N_8062,In_1025,In_1740);
xor U8063 (N_8063,In_4605,In_233);
and U8064 (N_8064,In_2912,In_1874);
or U8065 (N_8065,In_3893,In_4877);
and U8066 (N_8066,In_1456,In_3821);
and U8067 (N_8067,In_3838,In_2079);
nand U8068 (N_8068,In_50,In_205);
and U8069 (N_8069,In_491,In_2895);
and U8070 (N_8070,In_4502,In_2821);
nand U8071 (N_8071,In_4724,In_4377);
and U8072 (N_8072,In_1125,In_3249);
xnor U8073 (N_8073,In_1233,In_2588);
or U8074 (N_8074,In_3418,In_52);
or U8075 (N_8075,In_632,In_4928);
xnor U8076 (N_8076,In_639,In_4360);
nand U8077 (N_8077,In_2299,In_1480);
nor U8078 (N_8078,In_589,In_592);
or U8079 (N_8079,In_4841,In_1204);
or U8080 (N_8080,In_4959,In_1977);
or U8081 (N_8081,In_2465,In_1762);
nand U8082 (N_8082,In_4634,In_2646);
or U8083 (N_8083,In_1166,In_2988);
nor U8084 (N_8084,In_1506,In_4423);
nand U8085 (N_8085,In_1281,In_2809);
or U8086 (N_8086,In_4780,In_2335);
nand U8087 (N_8087,In_415,In_1142);
nor U8088 (N_8088,In_829,In_4660);
xnor U8089 (N_8089,In_917,In_4261);
nor U8090 (N_8090,In_2701,In_1138);
and U8091 (N_8091,In_3127,In_871);
nor U8092 (N_8092,In_3983,In_1104);
and U8093 (N_8093,In_1329,In_2508);
and U8094 (N_8094,In_92,In_4647);
xnor U8095 (N_8095,In_244,In_2494);
or U8096 (N_8096,In_3286,In_447);
xor U8097 (N_8097,In_2701,In_4201);
nor U8098 (N_8098,In_2292,In_729);
or U8099 (N_8099,In_116,In_1842);
xor U8100 (N_8100,In_604,In_3385);
xor U8101 (N_8101,In_2676,In_4157);
and U8102 (N_8102,In_4204,In_481);
nor U8103 (N_8103,In_4048,In_3630);
and U8104 (N_8104,In_1908,In_1007);
xor U8105 (N_8105,In_4634,In_303);
nand U8106 (N_8106,In_2882,In_3742);
nand U8107 (N_8107,In_3261,In_3807);
or U8108 (N_8108,In_2894,In_3096);
nor U8109 (N_8109,In_1873,In_2817);
nor U8110 (N_8110,In_1114,In_1266);
nand U8111 (N_8111,In_2717,In_3894);
nor U8112 (N_8112,In_4834,In_202);
or U8113 (N_8113,In_1415,In_1709);
or U8114 (N_8114,In_2769,In_866);
nand U8115 (N_8115,In_3816,In_2014);
or U8116 (N_8116,In_2785,In_1749);
xnor U8117 (N_8117,In_3745,In_2814);
and U8118 (N_8118,In_3239,In_3067);
nand U8119 (N_8119,In_4711,In_4706);
nand U8120 (N_8120,In_4574,In_2323);
xor U8121 (N_8121,In_1604,In_3401);
nor U8122 (N_8122,In_2324,In_4611);
and U8123 (N_8123,In_3515,In_1872);
nand U8124 (N_8124,In_3326,In_1690);
nor U8125 (N_8125,In_2601,In_1877);
xor U8126 (N_8126,In_3070,In_49);
or U8127 (N_8127,In_2337,In_4176);
nand U8128 (N_8128,In_1423,In_1757);
nand U8129 (N_8129,In_2557,In_162);
or U8130 (N_8130,In_1008,In_3740);
nor U8131 (N_8131,In_861,In_2826);
nor U8132 (N_8132,In_3417,In_1618);
or U8133 (N_8133,In_4420,In_2573);
xnor U8134 (N_8134,In_2890,In_854);
nor U8135 (N_8135,In_2084,In_2826);
nor U8136 (N_8136,In_4586,In_2417);
and U8137 (N_8137,In_1024,In_2661);
or U8138 (N_8138,In_1267,In_1069);
nand U8139 (N_8139,In_2551,In_1417);
or U8140 (N_8140,In_1543,In_3396);
nand U8141 (N_8141,In_3374,In_2317);
and U8142 (N_8142,In_3241,In_4454);
or U8143 (N_8143,In_2259,In_3118);
xor U8144 (N_8144,In_1776,In_1583);
or U8145 (N_8145,In_4708,In_3495);
nor U8146 (N_8146,In_2637,In_3817);
xor U8147 (N_8147,In_4345,In_4774);
or U8148 (N_8148,In_3673,In_4509);
or U8149 (N_8149,In_928,In_1178);
nor U8150 (N_8150,In_2949,In_4006);
nor U8151 (N_8151,In_3780,In_2389);
nor U8152 (N_8152,In_4499,In_4851);
nand U8153 (N_8153,In_1389,In_3584);
and U8154 (N_8154,In_364,In_4257);
nand U8155 (N_8155,In_1600,In_2548);
and U8156 (N_8156,In_2083,In_4856);
xor U8157 (N_8157,In_1981,In_4530);
and U8158 (N_8158,In_3360,In_591);
xor U8159 (N_8159,In_4845,In_4181);
nor U8160 (N_8160,In_709,In_2761);
or U8161 (N_8161,In_4411,In_4209);
and U8162 (N_8162,In_960,In_4784);
and U8163 (N_8163,In_2235,In_3102);
or U8164 (N_8164,In_767,In_4452);
or U8165 (N_8165,In_4492,In_267);
nand U8166 (N_8166,In_3772,In_3796);
nor U8167 (N_8167,In_1451,In_2011);
nand U8168 (N_8168,In_3852,In_1273);
and U8169 (N_8169,In_2039,In_1534);
nor U8170 (N_8170,In_2191,In_3346);
xor U8171 (N_8171,In_2136,In_2259);
or U8172 (N_8172,In_4296,In_2344);
and U8173 (N_8173,In_4008,In_4770);
or U8174 (N_8174,In_487,In_1377);
xor U8175 (N_8175,In_587,In_1853);
or U8176 (N_8176,In_292,In_1741);
or U8177 (N_8177,In_2332,In_3008);
or U8178 (N_8178,In_185,In_10);
nor U8179 (N_8179,In_4175,In_4096);
or U8180 (N_8180,In_246,In_81);
nand U8181 (N_8181,In_4760,In_3216);
nor U8182 (N_8182,In_3436,In_4737);
and U8183 (N_8183,In_2614,In_2327);
and U8184 (N_8184,In_1475,In_590);
or U8185 (N_8185,In_974,In_1130);
or U8186 (N_8186,In_4026,In_604);
nor U8187 (N_8187,In_3421,In_976);
xor U8188 (N_8188,In_1996,In_3459);
and U8189 (N_8189,In_1409,In_1496);
and U8190 (N_8190,In_32,In_3692);
nand U8191 (N_8191,In_1960,In_4414);
and U8192 (N_8192,In_1126,In_2577);
nor U8193 (N_8193,In_85,In_1204);
and U8194 (N_8194,In_1759,In_4290);
xor U8195 (N_8195,In_2059,In_320);
xor U8196 (N_8196,In_2496,In_628);
xor U8197 (N_8197,In_1493,In_225);
nor U8198 (N_8198,In_4969,In_1588);
or U8199 (N_8199,In_323,In_429);
and U8200 (N_8200,In_3375,In_163);
and U8201 (N_8201,In_4888,In_2366);
or U8202 (N_8202,In_1659,In_2356);
nor U8203 (N_8203,In_1939,In_1280);
xor U8204 (N_8204,In_4475,In_3948);
or U8205 (N_8205,In_809,In_2852);
xor U8206 (N_8206,In_412,In_1722);
nor U8207 (N_8207,In_4550,In_3218);
xnor U8208 (N_8208,In_1995,In_3091);
xor U8209 (N_8209,In_1406,In_3262);
or U8210 (N_8210,In_2791,In_692);
or U8211 (N_8211,In_214,In_4376);
xor U8212 (N_8212,In_1673,In_545);
nand U8213 (N_8213,In_4818,In_3782);
or U8214 (N_8214,In_4765,In_2800);
nor U8215 (N_8215,In_2977,In_4019);
xnor U8216 (N_8216,In_1812,In_4778);
xor U8217 (N_8217,In_1695,In_3745);
or U8218 (N_8218,In_1465,In_2470);
xnor U8219 (N_8219,In_2176,In_555);
nor U8220 (N_8220,In_3833,In_304);
nand U8221 (N_8221,In_1887,In_3806);
or U8222 (N_8222,In_1701,In_1576);
xor U8223 (N_8223,In_2361,In_4078);
nor U8224 (N_8224,In_920,In_4783);
xnor U8225 (N_8225,In_3022,In_2248);
xnor U8226 (N_8226,In_3205,In_1614);
xnor U8227 (N_8227,In_1397,In_4468);
xnor U8228 (N_8228,In_3454,In_1706);
nand U8229 (N_8229,In_1825,In_2951);
and U8230 (N_8230,In_239,In_4888);
nand U8231 (N_8231,In_635,In_1802);
and U8232 (N_8232,In_2722,In_1362);
or U8233 (N_8233,In_4324,In_2258);
nand U8234 (N_8234,In_2088,In_3612);
nand U8235 (N_8235,In_300,In_3460);
nor U8236 (N_8236,In_2181,In_1263);
xnor U8237 (N_8237,In_4386,In_2730);
and U8238 (N_8238,In_2834,In_1565);
nand U8239 (N_8239,In_4306,In_1993);
xnor U8240 (N_8240,In_1840,In_2454);
and U8241 (N_8241,In_4239,In_1622);
or U8242 (N_8242,In_971,In_1866);
and U8243 (N_8243,In_4194,In_2917);
xor U8244 (N_8244,In_3711,In_2488);
nor U8245 (N_8245,In_2844,In_1612);
nand U8246 (N_8246,In_2658,In_21);
or U8247 (N_8247,In_4935,In_994);
nor U8248 (N_8248,In_3347,In_3815);
nand U8249 (N_8249,In_3358,In_521);
and U8250 (N_8250,In_281,In_2706);
nor U8251 (N_8251,In_3015,In_478);
and U8252 (N_8252,In_970,In_1167);
and U8253 (N_8253,In_1964,In_3730);
xor U8254 (N_8254,In_3706,In_4891);
nor U8255 (N_8255,In_1005,In_3504);
and U8256 (N_8256,In_2904,In_2550);
nor U8257 (N_8257,In_685,In_3639);
nor U8258 (N_8258,In_273,In_87);
and U8259 (N_8259,In_490,In_883);
or U8260 (N_8260,In_716,In_3480);
xor U8261 (N_8261,In_1814,In_3415);
nor U8262 (N_8262,In_489,In_1957);
nand U8263 (N_8263,In_1817,In_2873);
xnor U8264 (N_8264,In_3693,In_82);
nor U8265 (N_8265,In_4685,In_1283);
nand U8266 (N_8266,In_723,In_4944);
nor U8267 (N_8267,In_1113,In_1238);
or U8268 (N_8268,In_3112,In_4199);
nor U8269 (N_8269,In_2666,In_3913);
xnor U8270 (N_8270,In_1473,In_32);
and U8271 (N_8271,In_4452,In_2720);
or U8272 (N_8272,In_4643,In_3421);
xnor U8273 (N_8273,In_4356,In_4024);
and U8274 (N_8274,In_1189,In_1133);
xnor U8275 (N_8275,In_3499,In_908);
nand U8276 (N_8276,In_1257,In_1466);
nor U8277 (N_8277,In_3120,In_3150);
nand U8278 (N_8278,In_3772,In_4648);
nand U8279 (N_8279,In_1306,In_4725);
nand U8280 (N_8280,In_3059,In_2727);
nor U8281 (N_8281,In_2294,In_4254);
xor U8282 (N_8282,In_2078,In_1090);
and U8283 (N_8283,In_1894,In_834);
and U8284 (N_8284,In_1161,In_2052);
nand U8285 (N_8285,In_747,In_2140);
nand U8286 (N_8286,In_2263,In_4174);
nor U8287 (N_8287,In_2319,In_1964);
nand U8288 (N_8288,In_3484,In_127);
and U8289 (N_8289,In_1172,In_514);
nand U8290 (N_8290,In_1503,In_399);
nor U8291 (N_8291,In_828,In_3725);
nand U8292 (N_8292,In_2321,In_2225);
xnor U8293 (N_8293,In_3392,In_1492);
and U8294 (N_8294,In_479,In_4554);
xnor U8295 (N_8295,In_1881,In_3466);
nor U8296 (N_8296,In_735,In_3690);
and U8297 (N_8297,In_1725,In_39);
nor U8298 (N_8298,In_1652,In_1436);
and U8299 (N_8299,In_613,In_1611);
nor U8300 (N_8300,In_394,In_4422);
nor U8301 (N_8301,In_3686,In_1454);
nand U8302 (N_8302,In_1052,In_1235);
or U8303 (N_8303,In_1660,In_2114);
xnor U8304 (N_8304,In_4111,In_361);
and U8305 (N_8305,In_609,In_1299);
nor U8306 (N_8306,In_2242,In_3995);
nor U8307 (N_8307,In_2296,In_4703);
and U8308 (N_8308,In_1184,In_360);
xor U8309 (N_8309,In_1701,In_4626);
or U8310 (N_8310,In_3861,In_1138);
and U8311 (N_8311,In_2160,In_3761);
xnor U8312 (N_8312,In_3865,In_3581);
nor U8313 (N_8313,In_4268,In_1309);
nand U8314 (N_8314,In_2348,In_602);
xor U8315 (N_8315,In_2077,In_2116);
nor U8316 (N_8316,In_1862,In_983);
and U8317 (N_8317,In_591,In_3136);
nand U8318 (N_8318,In_1319,In_2034);
and U8319 (N_8319,In_3580,In_3378);
xor U8320 (N_8320,In_2007,In_4124);
nor U8321 (N_8321,In_4749,In_2285);
nor U8322 (N_8322,In_3230,In_2279);
and U8323 (N_8323,In_106,In_2111);
xor U8324 (N_8324,In_1503,In_3989);
xor U8325 (N_8325,In_3676,In_3252);
xor U8326 (N_8326,In_4638,In_1377);
nor U8327 (N_8327,In_2939,In_4695);
xnor U8328 (N_8328,In_2796,In_4463);
nand U8329 (N_8329,In_1422,In_1071);
xor U8330 (N_8330,In_260,In_224);
xnor U8331 (N_8331,In_4375,In_1903);
or U8332 (N_8332,In_515,In_413);
xor U8333 (N_8333,In_150,In_2044);
nand U8334 (N_8334,In_59,In_2843);
or U8335 (N_8335,In_3412,In_1463);
nor U8336 (N_8336,In_3770,In_4161);
or U8337 (N_8337,In_163,In_1420);
nor U8338 (N_8338,In_1220,In_1621);
nor U8339 (N_8339,In_3194,In_137);
and U8340 (N_8340,In_1658,In_393);
xnor U8341 (N_8341,In_3166,In_172);
and U8342 (N_8342,In_948,In_3821);
or U8343 (N_8343,In_1873,In_4640);
or U8344 (N_8344,In_4099,In_4373);
nor U8345 (N_8345,In_4354,In_2619);
xnor U8346 (N_8346,In_2663,In_1621);
xnor U8347 (N_8347,In_4892,In_4966);
nand U8348 (N_8348,In_505,In_1163);
xnor U8349 (N_8349,In_733,In_3260);
nand U8350 (N_8350,In_3971,In_879);
nand U8351 (N_8351,In_567,In_2939);
or U8352 (N_8352,In_585,In_3514);
nand U8353 (N_8353,In_4931,In_4401);
and U8354 (N_8354,In_2876,In_2355);
or U8355 (N_8355,In_215,In_2442);
nand U8356 (N_8356,In_801,In_297);
xor U8357 (N_8357,In_2670,In_4534);
and U8358 (N_8358,In_1039,In_3309);
and U8359 (N_8359,In_25,In_2206);
nand U8360 (N_8360,In_4954,In_3004);
xor U8361 (N_8361,In_37,In_1660);
nor U8362 (N_8362,In_1883,In_952);
or U8363 (N_8363,In_42,In_4507);
and U8364 (N_8364,In_477,In_2094);
or U8365 (N_8365,In_474,In_3729);
or U8366 (N_8366,In_278,In_1613);
and U8367 (N_8367,In_3199,In_2595);
nand U8368 (N_8368,In_972,In_3252);
and U8369 (N_8369,In_3849,In_4861);
or U8370 (N_8370,In_180,In_2392);
or U8371 (N_8371,In_68,In_677);
or U8372 (N_8372,In_3170,In_619);
nand U8373 (N_8373,In_1409,In_2872);
nand U8374 (N_8374,In_772,In_970);
nand U8375 (N_8375,In_4135,In_128);
nand U8376 (N_8376,In_2463,In_2592);
xor U8377 (N_8377,In_4292,In_1089);
and U8378 (N_8378,In_648,In_935);
and U8379 (N_8379,In_3354,In_3264);
and U8380 (N_8380,In_4622,In_4582);
or U8381 (N_8381,In_2887,In_3849);
nand U8382 (N_8382,In_12,In_605);
nand U8383 (N_8383,In_1076,In_1581);
or U8384 (N_8384,In_1315,In_2494);
xor U8385 (N_8385,In_2153,In_4363);
nand U8386 (N_8386,In_730,In_1316);
or U8387 (N_8387,In_132,In_2329);
nor U8388 (N_8388,In_2771,In_275);
or U8389 (N_8389,In_3195,In_4564);
or U8390 (N_8390,In_366,In_3211);
xor U8391 (N_8391,In_4720,In_3628);
or U8392 (N_8392,In_2221,In_143);
nand U8393 (N_8393,In_2846,In_1684);
nor U8394 (N_8394,In_87,In_1752);
nor U8395 (N_8395,In_523,In_1452);
nand U8396 (N_8396,In_1274,In_3627);
nand U8397 (N_8397,In_71,In_2895);
nor U8398 (N_8398,In_89,In_2687);
nor U8399 (N_8399,In_399,In_837);
xnor U8400 (N_8400,In_836,In_2229);
nand U8401 (N_8401,In_1473,In_0);
and U8402 (N_8402,In_375,In_2857);
xor U8403 (N_8403,In_1814,In_1738);
and U8404 (N_8404,In_4257,In_3259);
or U8405 (N_8405,In_3837,In_3548);
nand U8406 (N_8406,In_1883,In_2409);
xnor U8407 (N_8407,In_2852,In_4419);
nand U8408 (N_8408,In_58,In_4910);
nand U8409 (N_8409,In_2073,In_4831);
and U8410 (N_8410,In_4531,In_4955);
nand U8411 (N_8411,In_1375,In_2151);
or U8412 (N_8412,In_361,In_1303);
nor U8413 (N_8413,In_1652,In_372);
nor U8414 (N_8414,In_1202,In_3150);
or U8415 (N_8415,In_911,In_2555);
or U8416 (N_8416,In_3977,In_153);
nor U8417 (N_8417,In_1460,In_2195);
or U8418 (N_8418,In_1800,In_505);
and U8419 (N_8419,In_3235,In_1644);
nand U8420 (N_8420,In_2455,In_4519);
or U8421 (N_8421,In_1907,In_2964);
nand U8422 (N_8422,In_3101,In_1855);
and U8423 (N_8423,In_4975,In_1554);
nand U8424 (N_8424,In_2601,In_1492);
or U8425 (N_8425,In_1555,In_750);
nor U8426 (N_8426,In_948,In_4738);
and U8427 (N_8427,In_2028,In_1072);
xnor U8428 (N_8428,In_462,In_2921);
nor U8429 (N_8429,In_2443,In_4074);
and U8430 (N_8430,In_3377,In_1226);
and U8431 (N_8431,In_2653,In_4194);
xor U8432 (N_8432,In_1749,In_287);
and U8433 (N_8433,In_589,In_1563);
xor U8434 (N_8434,In_920,In_3989);
nor U8435 (N_8435,In_4224,In_4188);
nand U8436 (N_8436,In_1989,In_108);
nand U8437 (N_8437,In_4231,In_4974);
nand U8438 (N_8438,In_4452,In_869);
xor U8439 (N_8439,In_655,In_2534);
or U8440 (N_8440,In_4562,In_2971);
nand U8441 (N_8441,In_2939,In_4006);
or U8442 (N_8442,In_2058,In_2541);
and U8443 (N_8443,In_2279,In_610);
nand U8444 (N_8444,In_3496,In_2574);
or U8445 (N_8445,In_2085,In_2662);
nor U8446 (N_8446,In_128,In_807);
xor U8447 (N_8447,In_296,In_358);
nor U8448 (N_8448,In_4433,In_3916);
and U8449 (N_8449,In_1956,In_946);
or U8450 (N_8450,In_4461,In_4509);
and U8451 (N_8451,In_3157,In_75);
nand U8452 (N_8452,In_3027,In_2854);
nand U8453 (N_8453,In_408,In_2935);
xnor U8454 (N_8454,In_4934,In_732);
and U8455 (N_8455,In_2953,In_3990);
nor U8456 (N_8456,In_325,In_456);
xor U8457 (N_8457,In_1013,In_4648);
or U8458 (N_8458,In_1400,In_3708);
nand U8459 (N_8459,In_2019,In_3166);
nand U8460 (N_8460,In_138,In_3284);
nor U8461 (N_8461,In_3508,In_3391);
xor U8462 (N_8462,In_3019,In_681);
nand U8463 (N_8463,In_3982,In_4378);
or U8464 (N_8464,In_3813,In_1044);
nor U8465 (N_8465,In_1484,In_2815);
and U8466 (N_8466,In_214,In_56);
nand U8467 (N_8467,In_3566,In_3609);
nand U8468 (N_8468,In_4166,In_1767);
and U8469 (N_8469,In_985,In_202);
nand U8470 (N_8470,In_1864,In_2447);
or U8471 (N_8471,In_358,In_1282);
and U8472 (N_8472,In_3256,In_1262);
xnor U8473 (N_8473,In_3309,In_4259);
nand U8474 (N_8474,In_1576,In_4215);
and U8475 (N_8475,In_3910,In_3333);
nand U8476 (N_8476,In_1209,In_3220);
and U8477 (N_8477,In_2685,In_1070);
nand U8478 (N_8478,In_3728,In_557);
and U8479 (N_8479,In_3059,In_1403);
and U8480 (N_8480,In_877,In_4502);
nand U8481 (N_8481,In_4344,In_2242);
xnor U8482 (N_8482,In_968,In_1236);
or U8483 (N_8483,In_2534,In_1209);
and U8484 (N_8484,In_3253,In_3151);
nand U8485 (N_8485,In_2880,In_3342);
nand U8486 (N_8486,In_3934,In_2548);
nor U8487 (N_8487,In_1007,In_4329);
or U8488 (N_8488,In_4311,In_2748);
and U8489 (N_8489,In_1330,In_3154);
nand U8490 (N_8490,In_176,In_2480);
nand U8491 (N_8491,In_1631,In_2866);
nand U8492 (N_8492,In_4668,In_1496);
nor U8493 (N_8493,In_1856,In_1766);
xnor U8494 (N_8494,In_302,In_3643);
nor U8495 (N_8495,In_292,In_790);
nand U8496 (N_8496,In_4790,In_1439);
nand U8497 (N_8497,In_2187,In_3296);
nand U8498 (N_8498,In_3460,In_4042);
nor U8499 (N_8499,In_2428,In_4673);
and U8500 (N_8500,In_419,In_807);
nand U8501 (N_8501,In_2002,In_2943);
or U8502 (N_8502,In_3179,In_878);
nor U8503 (N_8503,In_4804,In_3111);
nor U8504 (N_8504,In_2230,In_3264);
nor U8505 (N_8505,In_3194,In_913);
and U8506 (N_8506,In_828,In_3663);
nand U8507 (N_8507,In_2893,In_1284);
or U8508 (N_8508,In_1470,In_3164);
xor U8509 (N_8509,In_4964,In_4752);
nor U8510 (N_8510,In_3233,In_4365);
nand U8511 (N_8511,In_1751,In_101);
nor U8512 (N_8512,In_3764,In_3356);
xnor U8513 (N_8513,In_3309,In_4742);
and U8514 (N_8514,In_3844,In_3317);
nand U8515 (N_8515,In_4451,In_1272);
and U8516 (N_8516,In_2387,In_2637);
xor U8517 (N_8517,In_4577,In_2161);
nand U8518 (N_8518,In_4984,In_2564);
nor U8519 (N_8519,In_1273,In_942);
nand U8520 (N_8520,In_4797,In_3226);
nor U8521 (N_8521,In_3921,In_3408);
or U8522 (N_8522,In_996,In_4843);
xnor U8523 (N_8523,In_3139,In_584);
and U8524 (N_8524,In_502,In_1211);
or U8525 (N_8525,In_1770,In_3216);
xnor U8526 (N_8526,In_4513,In_4642);
nand U8527 (N_8527,In_1130,In_3659);
nand U8528 (N_8528,In_910,In_4974);
nand U8529 (N_8529,In_25,In_4929);
xnor U8530 (N_8530,In_253,In_2015);
or U8531 (N_8531,In_4857,In_4709);
xnor U8532 (N_8532,In_2095,In_4425);
and U8533 (N_8533,In_1360,In_4262);
nand U8534 (N_8534,In_2619,In_3778);
nand U8535 (N_8535,In_2893,In_2540);
xor U8536 (N_8536,In_3297,In_4000);
nand U8537 (N_8537,In_1479,In_3508);
and U8538 (N_8538,In_608,In_2369);
xor U8539 (N_8539,In_651,In_229);
and U8540 (N_8540,In_3507,In_4066);
or U8541 (N_8541,In_1126,In_1401);
or U8542 (N_8542,In_2038,In_190);
nand U8543 (N_8543,In_3171,In_456);
xnor U8544 (N_8544,In_2325,In_1391);
nor U8545 (N_8545,In_3845,In_3384);
xnor U8546 (N_8546,In_205,In_2242);
nand U8547 (N_8547,In_4383,In_2443);
or U8548 (N_8548,In_4774,In_4846);
and U8549 (N_8549,In_4881,In_852);
nand U8550 (N_8550,In_3348,In_648);
nand U8551 (N_8551,In_2669,In_944);
and U8552 (N_8552,In_4467,In_2735);
nand U8553 (N_8553,In_340,In_2892);
or U8554 (N_8554,In_1487,In_2743);
and U8555 (N_8555,In_485,In_2507);
nand U8556 (N_8556,In_710,In_845);
nand U8557 (N_8557,In_125,In_4708);
and U8558 (N_8558,In_1487,In_3115);
nor U8559 (N_8559,In_3293,In_1884);
nand U8560 (N_8560,In_3437,In_1117);
and U8561 (N_8561,In_2575,In_4296);
nor U8562 (N_8562,In_4031,In_3121);
xnor U8563 (N_8563,In_2616,In_3269);
xnor U8564 (N_8564,In_1522,In_2798);
or U8565 (N_8565,In_395,In_1306);
nor U8566 (N_8566,In_319,In_3176);
nor U8567 (N_8567,In_3818,In_3604);
xnor U8568 (N_8568,In_4752,In_3860);
or U8569 (N_8569,In_2796,In_4858);
xor U8570 (N_8570,In_2163,In_3006);
nor U8571 (N_8571,In_4601,In_1512);
and U8572 (N_8572,In_1875,In_2224);
or U8573 (N_8573,In_860,In_247);
or U8574 (N_8574,In_512,In_394);
and U8575 (N_8575,In_1913,In_3339);
or U8576 (N_8576,In_2188,In_3688);
and U8577 (N_8577,In_413,In_610);
nor U8578 (N_8578,In_3437,In_305);
or U8579 (N_8579,In_3377,In_2007);
xor U8580 (N_8580,In_1628,In_4665);
nand U8581 (N_8581,In_4583,In_2917);
and U8582 (N_8582,In_2905,In_3765);
nor U8583 (N_8583,In_22,In_2567);
xnor U8584 (N_8584,In_1762,In_2443);
xnor U8585 (N_8585,In_4898,In_3119);
xor U8586 (N_8586,In_1678,In_3572);
nor U8587 (N_8587,In_1371,In_3487);
xnor U8588 (N_8588,In_3486,In_3290);
nor U8589 (N_8589,In_3851,In_252);
xnor U8590 (N_8590,In_2383,In_1234);
nand U8591 (N_8591,In_4999,In_3856);
nand U8592 (N_8592,In_999,In_2492);
and U8593 (N_8593,In_1721,In_2401);
and U8594 (N_8594,In_4421,In_3775);
nor U8595 (N_8595,In_499,In_1033);
and U8596 (N_8596,In_1860,In_1686);
nand U8597 (N_8597,In_1155,In_4699);
nand U8598 (N_8598,In_3213,In_1422);
and U8599 (N_8599,In_2682,In_4384);
or U8600 (N_8600,In_2528,In_2600);
and U8601 (N_8601,In_4222,In_1772);
nand U8602 (N_8602,In_3312,In_3796);
or U8603 (N_8603,In_2854,In_3393);
xnor U8604 (N_8604,In_3964,In_855);
nand U8605 (N_8605,In_3618,In_749);
and U8606 (N_8606,In_953,In_3828);
or U8607 (N_8607,In_1056,In_3507);
and U8608 (N_8608,In_83,In_4399);
and U8609 (N_8609,In_3569,In_1640);
xnor U8610 (N_8610,In_1498,In_2874);
nor U8611 (N_8611,In_196,In_3934);
nor U8612 (N_8612,In_870,In_262);
or U8613 (N_8613,In_1414,In_917);
nor U8614 (N_8614,In_2262,In_1085);
or U8615 (N_8615,In_3867,In_875);
xnor U8616 (N_8616,In_3259,In_3547);
and U8617 (N_8617,In_1280,In_2558);
nand U8618 (N_8618,In_335,In_4147);
nand U8619 (N_8619,In_3975,In_2812);
and U8620 (N_8620,In_2984,In_1794);
nor U8621 (N_8621,In_3936,In_462);
xor U8622 (N_8622,In_2591,In_4082);
nor U8623 (N_8623,In_2191,In_2057);
xor U8624 (N_8624,In_4646,In_1286);
nor U8625 (N_8625,In_1244,In_3013);
xnor U8626 (N_8626,In_3927,In_1428);
nand U8627 (N_8627,In_4912,In_961);
nor U8628 (N_8628,In_3916,In_1827);
xor U8629 (N_8629,In_4988,In_2551);
nand U8630 (N_8630,In_569,In_4902);
and U8631 (N_8631,In_4105,In_3266);
and U8632 (N_8632,In_1422,In_3041);
or U8633 (N_8633,In_1356,In_254);
xor U8634 (N_8634,In_1211,In_4818);
or U8635 (N_8635,In_1692,In_1003);
xor U8636 (N_8636,In_2991,In_1662);
and U8637 (N_8637,In_2457,In_702);
or U8638 (N_8638,In_1511,In_1611);
and U8639 (N_8639,In_2947,In_744);
or U8640 (N_8640,In_1822,In_1677);
or U8641 (N_8641,In_4551,In_2718);
nand U8642 (N_8642,In_2580,In_2442);
nand U8643 (N_8643,In_4289,In_4141);
nand U8644 (N_8644,In_639,In_3658);
nor U8645 (N_8645,In_2352,In_1617);
xor U8646 (N_8646,In_1061,In_2323);
nand U8647 (N_8647,In_401,In_2263);
or U8648 (N_8648,In_343,In_3860);
or U8649 (N_8649,In_572,In_3570);
and U8650 (N_8650,In_1806,In_1415);
nor U8651 (N_8651,In_1447,In_2063);
xnor U8652 (N_8652,In_574,In_769);
and U8653 (N_8653,In_623,In_87);
xnor U8654 (N_8654,In_69,In_4690);
xnor U8655 (N_8655,In_2044,In_2731);
nand U8656 (N_8656,In_1973,In_1721);
and U8657 (N_8657,In_3040,In_1928);
nand U8658 (N_8658,In_2152,In_730);
or U8659 (N_8659,In_136,In_16);
nand U8660 (N_8660,In_1161,In_1463);
xor U8661 (N_8661,In_3127,In_663);
and U8662 (N_8662,In_1622,In_2962);
or U8663 (N_8663,In_3874,In_4762);
nor U8664 (N_8664,In_2355,In_1127);
or U8665 (N_8665,In_3247,In_2866);
or U8666 (N_8666,In_4086,In_1373);
and U8667 (N_8667,In_83,In_838);
or U8668 (N_8668,In_4596,In_3578);
nor U8669 (N_8669,In_715,In_4255);
or U8670 (N_8670,In_3615,In_4406);
nand U8671 (N_8671,In_947,In_64);
or U8672 (N_8672,In_2522,In_2145);
nor U8673 (N_8673,In_1843,In_1928);
xnor U8674 (N_8674,In_4992,In_1853);
xor U8675 (N_8675,In_2130,In_2077);
or U8676 (N_8676,In_3911,In_145);
nor U8677 (N_8677,In_2091,In_2948);
or U8678 (N_8678,In_50,In_4371);
nor U8679 (N_8679,In_3499,In_771);
nand U8680 (N_8680,In_4814,In_1524);
or U8681 (N_8681,In_1337,In_4401);
or U8682 (N_8682,In_2471,In_2983);
nor U8683 (N_8683,In_2153,In_2812);
nor U8684 (N_8684,In_4958,In_1345);
nand U8685 (N_8685,In_866,In_4758);
or U8686 (N_8686,In_229,In_4136);
nand U8687 (N_8687,In_3273,In_2170);
or U8688 (N_8688,In_1745,In_4459);
and U8689 (N_8689,In_1566,In_4208);
and U8690 (N_8690,In_1613,In_366);
or U8691 (N_8691,In_3750,In_3714);
xor U8692 (N_8692,In_359,In_1025);
or U8693 (N_8693,In_3265,In_3647);
nor U8694 (N_8694,In_4966,In_580);
or U8695 (N_8695,In_142,In_664);
nand U8696 (N_8696,In_3915,In_4508);
nand U8697 (N_8697,In_2840,In_3694);
nor U8698 (N_8698,In_540,In_2007);
and U8699 (N_8699,In_2911,In_1446);
nand U8700 (N_8700,In_1754,In_824);
or U8701 (N_8701,In_637,In_615);
and U8702 (N_8702,In_4580,In_2553);
nor U8703 (N_8703,In_457,In_2654);
nor U8704 (N_8704,In_2038,In_3022);
nor U8705 (N_8705,In_4311,In_4331);
nand U8706 (N_8706,In_1064,In_997);
or U8707 (N_8707,In_1260,In_3800);
and U8708 (N_8708,In_1780,In_556);
or U8709 (N_8709,In_4483,In_1032);
nand U8710 (N_8710,In_561,In_2674);
and U8711 (N_8711,In_969,In_608);
and U8712 (N_8712,In_43,In_3247);
and U8713 (N_8713,In_763,In_4437);
and U8714 (N_8714,In_732,In_246);
nor U8715 (N_8715,In_247,In_1716);
or U8716 (N_8716,In_2784,In_662);
and U8717 (N_8717,In_3641,In_2483);
nor U8718 (N_8718,In_4896,In_4166);
nand U8719 (N_8719,In_1747,In_2963);
nor U8720 (N_8720,In_1448,In_2229);
and U8721 (N_8721,In_2842,In_155);
xnor U8722 (N_8722,In_4968,In_4719);
nand U8723 (N_8723,In_4849,In_2220);
and U8724 (N_8724,In_2286,In_4312);
nor U8725 (N_8725,In_2601,In_4817);
nor U8726 (N_8726,In_2162,In_4417);
or U8727 (N_8727,In_3287,In_269);
xnor U8728 (N_8728,In_1880,In_4640);
nor U8729 (N_8729,In_3940,In_2254);
nand U8730 (N_8730,In_618,In_3351);
and U8731 (N_8731,In_2996,In_771);
and U8732 (N_8732,In_3145,In_3091);
nor U8733 (N_8733,In_2273,In_4657);
or U8734 (N_8734,In_418,In_1005);
or U8735 (N_8735,In_3699,In_1717);
or U8736 (N_8736,In_1362,In_4331);
or U8737 (N_8737,In_4066,In_437);
and U8738 (N_8738,In_1943,In_1821);
nor U8739 (N_8739,In_1181,In_4850);
nor U8740 (N_8740,In_2573,In_4400);
nor U8741 (N_8741,In_4847,In_3402);
xor U8742 (N_8742,In_2663,In_3797);
or U8743 (N_8743,In_1404,In_2572);
or U8744 (N_8744,In_2427,In_409);
nand U8745 (N_8745,In_677,In_1651);
nor U8746 (N_8746,In_772,In_2796);
xor U8747 (N_8747,In_493,In_3564);
nand U8748 (N_8748,In_1831,In_3078);
nand U8749 (N_8749,In_547,In_2462);
and U8750 (N_8750,In_236,In_1341);
and U8751 (N_8751,In_2301,In_4923);
and U8752 (N_8752,In_4481,In_3115);
xor U8753 (N_8753,In_1703,In_1595);
and U8754 (N_8754,In_224,In_2137);
or U8755 (N_8755,In_4638,In_3056);
xor U8756 (N_8756,In_2810,In_901);
nand U8757 (N_8757,In_2421,In_722);
nor U8758 (N_8758,In_1543,In_1249);
and U8759 (N_8759,In_4816,In_1639);
nor U8760 (N_8760,In_4539,In_2981);
or U8761 (N_8761,In_2843,In_2184);
xor U8762 (N_8762,In_791,In_213);
xnor U8763 (N_8763,In_3898,In_4582);
and U8764 (N_8764,In_2757,In_3862);
xor U8765 (N_8765,In_666,In_3009);
nor U8766 (N_8766,In_1074,In_3638);
or U8767 (N_8767,In_4665,In_3189);
nand U8768 (N_8768,In_1067,In_2396);
nand U8769 (N_8769,In_3266,In_1582);
nand U8770 (N_8770,In_4934,In_2773);
xnor U8771 (N_8771,In_1760,In_2755);
or U8772 (N_8772,In_3495,In_4164);
or U8773 (N_8773,In_3489,In_3968);
or U8774 (N_8774,In_1541,In_977);
xnor U8775 (N_8775,In_1182,In_2157);
nor U8776 (N_8776,In_4392,In_549);
nand U8777 (N_8777,In_2331,In_2997);
or U8778 (N_8778,In_4488,In_3488);
nand U8779 (N_8779,In_3538,In_82);
xnor U8780 (N_8780,In_123,In_2218);
nor U8781 (N_8781,In_12,In_4390);
nand U8782 (N_8782,In_3764,In_4525);
and U8783 (N_8783,In_3411,In_2277);
and U8784 (N_8784,In_1738,In_417);
or U8785 (N_8785,In_152,In_1567);
xor U8786 (N_8786,In_1287,In_1692);
or U8787 (N_8787,In_3450,In_4202);
and U8788 (N_8788,In_1098,In_4755);
or U8789 (N_8789,In_3388,In_3603);
or U8790 (N_8790,In_249,In_4127);
nand U8791 (N_8791,In_2366,In_3267);
nor U8792 (N_8792,In_428,In_3671);
and U8793 (N_8793,In_887,In_4242);
nor U8794 (N_8794,In_159,In_3795);
xor U8795 (N_8795,In_699,In_4654);
nand U8796 (N_8796,In_4228,In_3156);
xor U8797 (N_8797,In_2524,In_4132);
nand U8798 (N_8798,In_309,In_3353);
or U8799 (N_8799,In_387,In_3091);
or U8800 (N_8800,In_4073,In_3348);
nand U8801 (N_8801,In_2704,In_4225);
nor U8802 (N_8802,In_2944,In_2706);
nor U8803 (N_8803,In_3002,In_779);
or U8804 (N_8804,In_2298,In_3932);
and U8805 (N_8805,In_1431,In_576);
nor U8806 (N_8806,In_1804,In_357);
nand U8807 (N_8807,In_3023,In_849);
nor U8808 (N_8808,In_2832,In_3152);
nand U8809 (N_8809,In_2958,In_3458);
nor U8810 (N_8810,In_3115,In_599);
nor U8811 (N_8811,In_3724,In_2671);
nor U8812 (N_8812,In_964,In_3187);
nor U8813 (N_8813,In_788,In_1736);
xor U8814 (N_8814,In_768,In_4736);
and U8815 (N_8815,In_2858,In_1430);
nor U8816 (N_8816,In_4997,In_2531);
xnor U8817 (N_8817,In_4296,In_4464);
xor U8818 (N_8818,In_1443,In_99);
nor U8819 (N_8819,In_55,In_3122);
xnor U8820 (N_8820,In_1246,In_1443);
and U8821 (N_8821,In_2401,In_4044);
xnor U8822 (N_8822,In_987,In_204);
or U8823 (N_8823,In_4580,In_1782);
xnor U8824 (N_8824,In_3705,In_3360);
or U8825 (N_8825,In_3895,In_2645);
xnor U8826 (N_8826,In_3606,In_1230);
xnor U8827 (N_8827,In_1325,In_2976);
nor U8828 (N_8828,In_1610,In_2853);
or U8829 (N_8829,In_2492,In_2738);
and U8830 (N_8830,In_868,In_2685);
nand U8831 (N_8831,In_457,In_111);
and U8832 (N_8832,In_856,In_1701);
nand U8833 (N_8833,In_605,In_4732);
xnor U8834 (N_8834,In_741,In_756);
or U8835 (N_8835,In_4152,In_2120);
xor U8836 (N_8836,In_4326,In_2371);
or U8837 (N_8837,In_1221,In_690);
and U8838 (N_8838,In_3900,In_3856);
nor U8839 (N_8839,In_4076,In_4231);
nor U8840 (N_8840,In_3928,In_722);
nand U8841 (N_8841,In_4617,In_504);
nor U8842 (N_8842,In_2545,In_4017);
and U8843 (N_8843,In_4980,In_3769);
or U8844 (N_8844,In_840,In_2506);
and U8845 (N_8845,In_2196,In_4549);
and U8846 (N_8846,In_143,In_4200);
nor U8847 (N_8847,In_320,In_3655);
or U8848 (N_8848,In_4094,In_768);
nand U8849 (N_8849,In_1779,In_2149);
xor U8850 (N_8850,In_2017,In_4116);
nand U8851 (N_8851,In_1723,In_4677);
nor U8852 (N_8852,In_2252,In_4626);
or U8853 (N_8853,In_3242,In_3018);
xnor U8854 (N_8854,In_4266,In_970);
nand U8855 (N_8855,In_940,In_3184);
xor U8856 (N_8856,In_1254,In_3043);
nor U8857 (N_8857,In_2494,In_2199);
and U8858 (N_8858,In_2004,In_1933);
nand U8859 (N_8859,In_355,In_2909);
nor U8860 (N_8860,In_2484,In_1181);
nor U8861 (N_8861,In_3534,In_1367);
nand U8862 (N_8862,In_2708,In_4418);
or U8863 (N_8863,In_539,In_2616);
and U8864 (N_8864,In_4782,In_4583);
xnor U8865 (N_8865,In_721,In_569);
nor U8866 (N_8866,In_1890,In_4663);
or U8867 (N_8867,In_4099,In_3035);
nand U8868 (N_8868,In_894,In_1559);
and U8869 (N_8869,In_2206,In_3774);
or U8870 (N_8870,In_3985,In_3967);
and U8871 (N_8871,In_3216,In_2903);
or U8872 (N_8872,In_4167,In_1858);
and U8873 (N_8873,In_3579,In_4836);
xnor U8874 (N_8874,In_1034,In_1680);
nor U8875 (N_8875,In_2611,In_2294);
nand U8876 (N_8876,In_3618,In_4270);
or U8877 (N_8877,In_532,In_1520);
and U8878 (N_8878,In_4627,In_2701);
and U8879 (N_8879,In_3008,In_4695);
xnor U8880 (N_8880,In_4934,In_2888);
and U8881 (N_8881,In_752,In_3958);
nor U8882 (N_8882,In_4916,In_2620);
xor U8883 (N_8883,In_4509,In_3787);
nand U8884 (N_8884,In_508,In_144);
nand U8885 (N_8885,In_2813,In_3601);
nand U8886 (N_8886,In_2498,In_2221);
nand U8887 (N_8887,In_3072,In_3507);
nor U8888 (N_8888,In_879,In_2067);
and U8889 (N_8889,In_2824,In_2456);
or U8890 (N_8890,In_3249,In_2995);
nor U8891 (N_8891,In_3061,In_540);
nor U8892 (N_8892,In_4453,In_1518);
nor U8893 (N_8893,In_2316,In_2488);
nor U8894 (N_8894,In_1188,In_3654);
xor U8895 (N_8895,In_1246,In_2622);
and U8896 (N_8896,In_2658,In_2057);
and U8897 (N_8897,In_1614,In_1042);
nor U8898 (N_8898,In_4541,In_4996);
xor U8899 (N_8899,In_3607,In_3748);
nand U8900 (N_8900,In_1411,In_120);
xor U8901 (N_8901,In_4684,In_53);
and U8902 (N_8902,In_3691,In_3018);
or U8903 (N_8903,In_115,In_3547);
nand U8904 (N_8904,In_3110,In_4323);
and U8905 (N_8905,In_1278,In_3509);
nand U8906 (N_8906,In_1931,In_4789);
xor U8907 (N_8907,In_3379,In_355);
xor U8908 (N_8908,In_2662,In_2247);
nor U8909 (N_8909,In_1797,In_2569);
nand U8910 (N_8910,In_3291,In_3161);
nor U8911 (N_8911,In_2322,In_1890);
nand U8912 (N_8912,In_1010,In_2240);
or U8913 (N_8913,In_1342,In_1182);
or U8914 (N_8914,In_2418,In_3433);
xor U8915 (N_8915,In_1703,In_4119);
nand U8916 (N_8916,In_4474,In_1234);
nand U8917 (N_8917,In_1933,In_891);
and U8918 (N_8918,In_3986,In_2434);
nand U8919 (N_8919,In_298,In_4887);
or U8920 (N_8920,In_3552,In_4645);
xnor U8921 (N_8921,In_922,In_2164);
nand U8922 (N_8922,In_4476,In_4920);
nor U8923 (N_8923,In_3129,In_1358);
or U8924 (N_8924,In_1629,In_1326);
nor U8925 (N_8925,In_4505,In_957);
nor U8926 (N_8926,In_4137,In_2993);
nand U8927 (N_8927,In_4510,In_1048);
and U8928 (N_8928,In_1939,In_1850);
or U8929 (N_8929,In_1252,In_3956);
and U8930 (N_8930,In_435,In_3172);
nor U8931 (N_8931,In_2791,In_3153);
nor U8932 (N_8932,In_781,In_1262);
xor U8933 (N_8933,In_2573,In_704);
or U8934 (N_8934,In_1462,In_4118);
and U8935 (N_8935,In_1238,In_3527);
nand U8936 (N_8936,In_1837,In_4758);
nand U8937 (N_8937,In_2519,In_3404);
xnor U8938 (N_8938,In_4080,In_2988);
nor U8939 (N_8939,In_1830,In_3881);
nand U8940 (N_8940,In_4512,In_3240);
xor U8941 (N_8941,In_3778,In_3768);
xnor U8942 (N_8942,In_4451,In_468);
xnor U8943 (N_8943,In_3039,In_1821);
nand U8944 (N_8944,In_3038,In_2425);
or U8945 (N_8945,In_688,In_1185);
nand U8946 (N_8946,In_1371,In_2564);
nor U8947 (N_8947,In_4639,In_3852);
or U8948 (N_8948,In_946,In_776);
nor U8949 (N_8949,In_4960,In_3599);
and U8950 (N_8950,In_4713,In_1179);
or U8951 (N_8951,In_4630,In_4269);
or U8952 (N_8952,In_1514,In_4453);
nor U8953 (N_8953,In_1853,In_1770);
and U8954 (N_8954,In_4273,In_1948);
xor U8955 (N_8955,In_4054,In_2677);
nand U8956 (N_8956,In_3846,In_122);
nand U8957 (N_8957,In_2116,In_4138);
and U8958 (N_8958,In_4385,In_1174);
and U8959 (N_8959,In_3120,In_3195);
nand U8960 (N_8960,In_2852,In_3552);
or U8961 (N_8961,In_4948,In_546);
or U8962 (N_8962,In_904,In_3266);
or U8963 (N_8963,In_1705,In_3130);
and U8964 (N_8964,In_4361,In_202);
or U8965 (N_8965,In_1521,In_3188);
and U8966 (N_8966,In_233,In_1566);
nor U8967 (N_8967,In_4208,In_3389);
nor U8968 (N_8968,In_2089,In_3326);
and U8969 (N_8969,In_2513,In_300);
and U8970 (N_8970,In_4833,In_3770);
nand U8971 (N_8971,In_2000,In_4986);
or U8972 (N_8972,In_4366,In_3205);
nor U8973 (N_8973,In_3058,In_1360);
nor U8974 (N_8974,In_4825,In_1133);
and U8975 (N_8975,In_1603,In_3974);
and U8976 (N_8976,In_3172,In_1210);
xnor U8977 (N_8977,In_2773,In_651);
nor U8978 (N_8978,In_1026,In_2152);
or U8979 (N_8979,In_3279,In_1740);
xnor U8980 (N_8980,In_2457,In_598);
and U8981 (N_8981,In_4794,In_1592);
nor U8982 (N_8982,In_3446,In_2971);
nand U8983 (N_8983,In_4022,In_2976);
nor U8984 (N_8984,In_3742,In_879);
xor U8985 (N_8985,In_4432,In_4399);
nor U8986 (N_8986,In_3448,In_3357);
xnor U8987 (N_8987,In_2911,In_1545);
or U8988 (N_8988,In_468,In_3426);
nor U8989 (N_8989,In_3652,In_4694);
or U8990 (N_8990,In_3972,In_1266);
or U8991 (N_8991,In_2067,In_1203);
nand U8992 (N_8992,In_4706,In_2678);
or U8993 (N_8993,In_3950,In_4906);
nand U8994 (N_8994,In_2940,In_939);
nor U8995 (N_8995,In_1468,In_2151);
or U8996 (N_8996,In_1631,In_215);
or U8997 (N_8997,In_1516,In_888);
nor U8998 (N_8998,In_4519,In_2250);
nand U8999 (N_8999,In_4877,In_2524);
nand U9000 (N_9000,In_484,In_1322);
xnor U9001 (N_9001,In_3301,In_274);
and U9002 (N_9002,In_1669,In_1087);
nor U9003 (N_9003,In_2121,In_3563);
nand U9004 (N_9004,In_2536,In_1067);
xor U9005 (N_9005,In_2616,In_1180);
or U9006 (N_9006,In_4879,In_4554);
or U9007 (N_9007,In_1237,In_1548);
and U9008 (N_9008,In_1613,In_585);
nor U9009 (N_9009,In_2838,In_3095);
nor U9010 (N_9010,In_4009,In_692);
nor U9011 (N_9011,In_4659,In_2144);
and U9012 (N_9012,In_151,In_2443);
or U9013 (N_9013,In_310,In_4815);
or U9014 (N_9014,In_2951,In_4572);
nor U9015 (N_9015,In_4253,In_4324);
xor U9016 (N_9016,In_4611,In_3119);
or U9017 (N_9017,In_179,In_750);
or U9018 (N_9018,In_4339,In_3566);
and U9019 (N_9019,In_2470,In_2610);
nor U9020 (N_9020,In_1817,In_1396);
nand U9021 (N_9021,In_981,In_3434);
xor U9022 (N_9022,In_2892,In_1611);
xnor U9023 (N_9023,In_1649,In_4976);
nand U9024 (N_9024,In_1794,In_4673);
or U9025 (N_9025,In_29,In_4550);
and U9026 (N_9026,In_4779,In_3682);
xnor U9027 (N_9027,In_431,In_1736);
and U9028 (N_9028,In_1543,In_4729);
nand U9029 (N_9029,In_2703,In_3440);
or U9030 (N_9030,In_1887,In_3296);
nand U9031 (N_9031,In_4184,In_728);
or U9032 (N_9032,In_1431,In_3726);
nor U9033 (N_9033,In_4003,In_4359);
or U9034 (N_9034,In_746,In_4733);
nand U9035 (N_9035,In_1066,In_321);
xnor U9036 (N_9036,In_3348,In_2700);
nand U9037 (N_9037,In_2666,In_18);
nand U9038 (N_9038,In_4423,In_3797);
or U9039 (N_9039,In_502,In_1076);
xnor U9040 (N_9040,In_1902,In_3082);
nor U9041 (N_9041,In_1633,In_3624);
xor U9042 (N_9042,In_684,In_3400);
xor U9043 (N_9043,In_4939,In_3777);
or U9044 (N_9044,In_3311,In_619);
nand U9045 (N_9045,In_4744,In_4883);
nor U9046 (N_9046,In_1457,In_4340);
nor U9047 (N_9047,In_4662,In_2070);
nand U9048 (N_9048,In_2546,In_3211);
or U9049 (N_9049,In_2573,In_3836);
xnor U9050 (N_9050,In_270,In_4150);
or U9051 (N_9051,In_493,In_3713);
nor U9052 (N_9052,In_3247,In_318);
nand U9053 (N_9053,In_3016,In_614);
xnor U9054 (N_9054,In_861,In_164);
nand U9055 (N_9055,In_2421,In_4332);
and U9056 (N_9056,In_4196,In_689);
nand U9057 (N_9057,In_2476,In_37);
and U9058 (N_9058,In_980,In_336);
nand U9059 (N_9059,In_526,In_4939);
xor U9060 (N_9060,In_4282,In_347);
or U9061 (N_9061,In_3336,In_771);
nor U9062 (N_9062,In_4930,In_513);
nor U9063 (N_9063,In_3498,In_2529);
nor U9064 (N_9064,In_4899,In_4073);
or U9065 (N_9065,In_4751,In_474);
and U9066 (N_9066,In_210,In_2509);
and U9067 (N_9067,In_1477,In_2722);
nand U9068 (N_9068,In_375,In_2657);
and U9069 (N_9069,In_2204,In_3201);
or U9070 (N_9070,In_4694,In_4232);
nor U9071 (N_9071,In_4132,In_1121);
and U9072 (N_9072,In_3446,In_3793);
xor U9073 (N_9073,In_4916,In_3822);
and U9074 (N_9074,In_206,In_1682);
nand U9075 (N_9075,In_2177,In_1657);
and U9076 (N_9076,In_1654,In_1750);
nand U9077 (N_9077,In_1730,In_3196);
and U9078 (N_9078,In_3677,In_3272);
nand U9079 (N_9079,In_4712,In_2247);
or U9080 (N_9080,In_4111,In_2389);
nand U9081 (N_9081,In_3876,In_2673);
nand U9082 (N_9082,In_1318,In_3260);
and U9083 (N_9083,In_1122,In_3111);
nand U9084 (N_9084,In_761,In_362);
nand U9085 (N_9085,In_3049,In_1023);
nor U9086 (N_9086,In_1692,In_3585);
nor U9087 (N_9087,In_3560,In_3151);
xor U9088 (N_9088,In_4243,In_553);
or U9089 (N_9089,In_3910,In_4518);
or U9090 (N_9090,In_4666,In_1920);
nand U9091 (N_9091,In_465,In_2846);
nand U9092 (N_9092,In_2734,In_3976);
nand U9093 (N_9093,In_4616,In_3666);
and U9094 (N_9094,In_1370,In_915);
and U9095 (N_9095,In_3549,In_2277);
or U9096 (N_9096,In_349,In_4939);
xor U9097 (N_9097,In_2784,In_543);
xnor U9098 (N_9098,In_1378,In_280);
nor U9099 (N_9099,In_819,In_2315);
and U9100 (N_9100,In_3000,In_3251);
xnor U9101 (N_9101,In_1176,In_4578);
nor U9102 (N_9102,In_444,In_885);
or U9103 (N_9103,In_1588,In_823);
xor U9104 (N_9104,In_1379,In_3596);
nand U9105 (N_9105,In_599,In_4789);
or U9106 (N_9106,In_3760,In_2704);
or U9107 (N_9107,In_3315,In_102);
or U9108 (N_9108,In_4798,In_2819);
nor U9109 (N_9109,In_3301,In_2239);
or U9110 (N_9110,In_1067,In_2008);
xnor U9111 (N_9111,In_50,In_1535);
or U9112 (N_9112,In_3612,In_4360);
or U9113 (N_9113,In_4646,In_3951);
and U9114 (N_9114,In_3676,In_3384);
nand U9115 (N_9115,In_32,In_3088);
nand U9116 (N_9116,In_2357,In_1003);
xnor U9117 (N_9117,In_436,In_3836);
nand U9118 (N_9118,In_3125,In_1635);
and U9119 (N_9119,In_1023,In_4407);
or U9120 (N_9120,In_1050,In_1535);
nor U9121 (N_9121,In_1496,In_3241);
xnor U9122 (N_9122,In_2975,In_3882);
or U9123 (N_9123,In_4300,In_1410);
xor U9124 (N_9124,In_1077,In_4785);
nor U9125 (N_9125,In_1170,In_2765);
xnor U9126 (N_9126,In_3926,In_4505);
or U9127 (N_9127,In_3421,In_909);
nand U9128 (N_9128,In_4323,In_2688);
nand U9129 (N_9129,In_2714,In_3723);
xnor U9130 (N_9130,In_2852,In_551);
or U9131 (N_9131,In_2692,In_103);
xor U9132 (N_9132,In_3931,In_1206);
nor U9133 (N_9133,In_4797,In_681);
nor U9134 (N_9134,In_3225,In_901);
xor U9135 (N_9135,In_4584,In_2155);
or U9136 (N_9136,In_1328,In_3691);
nand U9137 (N_9137,In_118,In_2616);
nor U9138 (N_9138,In_4635,In_4614);
xor U9139 (N_9139,In_4392,In_1344);
nand U9140 (N_9140,In_988,In_2436);
and U9141 (N_9141,In_4592,In_2300);
and U9142 (N_9142,In_568,In_3335);
and U9143 (N_9143,In_3484,In_41);
nor U9144 (N_9144,In_2796,In_1923);
xnor U9145 (N_9145,In_1450,In_2280);
nand U9146 (N_9146,In_2706,In_3925);
nand U9147 (N_9147,In_3074,In_2371);
nor U9148 (N_9148,In_4068,In_1105);
or U9149 (N_9149,In_4517,In_99);
or U9150 (N_9150,In_3382,In_2020);
xnor U9151 (N_9151,In_2958,In_2933);
nor U9152 (N_9152,In_1437,In_4617);
or U9153 (N_9153,In_2500,In_2249);
nor U9154 (N_9154,In_788,In_2215);
nand U9155 (N_9155,In_2453,In_4415);
or U9156 (N_9156,In_2905,In_551);
nand U9157 (N_9157,In_4280,In_3975);
nand U9158 (N_9158,In_1944,In_1303);
xnor U9159 (N_9159,In_447,In_1241);
and U9160 (N_9160,In_1675,In_2937);
nand U9161 (N_9161,In_2581,In_4862);
nor U9162 (N_9162,In_1111,In_3098);
xnor U9163 (N_9163,In_2890,In_4277);
and U9164 (N_9164,In_3010,In_1074);
or U9165 (N_9165,In_2005,In_3932);
or U9166 (N_9166,In_2382,In_872);
nand U9167 (N_9167,In_483,In_2784);
nand U9168 (N_9168,In_721,In_296);
and U9169 (N_9169,In_3437,In_607);
nor U9170 (N_9170,In_4336,In_1362);
and U9171 (N_9171,In_260,In_4379);
nand U9172 (N_9172,In_4235,In_709);
or U9173 (N_9173,In_2708,In_2860);
xor U9174 (N_9174,In_1646,In_1587);
xnor U9175 (N_9175,In_4973,In_1623);
or U9176 (N_9176,In_1313,In_4677);
and U9177 (N_9177,In_3809,In_1016);
nor U9178 (N_9178,In_4454,In_4942);
nand U9179 (N_9179,In_2988,In_1057);
and U9180 (N_9180,In_1227,In_1870);
nand U9181 (N_9181,In_451,In_1950);
or U9182 (N_9182,In_2980,In_1188);
and U9183 (N_9183,In_1753,In_3837);
nand U9184 (N_9184,In_3685,In_1433);
nand U9185 (N_9185,In_3370,In_418);
xor U9186 (N_9186,In_75,In_3470);
nand U9187 (N_9187,In_3557,In_1106);
nor U9188 (N_9188,In_578,In_3406);
nand U9189 (N_9189,In_663,In_624);
xnor U9190 (N_9190,In_3651,In_4374);
nand U9191 (N_9191,In_2073,In_3302);
or U9192 (N_9192,In_2453,In_3778);
or U9193 (N_9193,In_4518,In_2516);
nand U9194 (N_9194,In_1925,In_1122);
nand U9195 (N_9195,In_78,In_4781);
nand U9196 (N_9196,In_1937,In_3157);
nand U9197 (N_9197,In_2225,In_2349);
nand U9198 (N_9198,In_2410,In_4481);
and U9199 (N_9199,In_4806,In_908);
nand U9200 (N_9200,In_3850,In_3805);
and U9201 (N_9201,In_2004,In_43);
or U9202 (N_9202,In_4577,In_4550);
or U9203 (N_9203,In_4993,In_4738);
and U9204 (N_9204,In_1695,In_1277);
nand U9205 (N_9205,In_2317,In_4658);
or U9206 (N_9206,In_2656,In_4120);
and U9207 (N_9207,In_4877,In_1706);
nor U9208 (N_9208,In_2865,In_1827);
and U9209 (N_9209,In_609,In_1266);
nor U9210 (N_9210,In_1749,In_1324);
or U9211 (N_9211,In_4590,In_4723);
xnor U9212 (N_9212,In_1837,In_936);
nor U9213 (N_9213,In_1690,In_837);
nand U9214 (N_9214,In_3175,In_878);
nand U9215 (N_9215,In_740,In_2283);
xnor U9216 (N_9216,In_3899,In_3334);
and U9217 (N_9217,In_1062,In_4326);
xnor U9218 (N_9218,In_4505,In_3908);
and U9219 (N_9219,In_4644,In_3797);
and U9220 (N_9220,In_1749,In_3674);
or U9221 (N_9221,In_597,In_1666);
nor U9222 (N_9222,In_1777,In_187);
or U9223 (N_9223,In_1053,In_4411);
or U9224 (N_9224,In_4245,In_338);
xor U9225 (N_9225,In_3926,In_3847);
or U9226 (N_9226,In_4031,In_2772);
nor U9227 (N_9227,In_3016,In_3714);
nand U9228 (N_9228,In_3067,In_36);
and U9229 (N_9229,In_4933,In_4942);
xor U9230 (N_9230,In_921,In_4506);
xnor U9231 (N_9231,In_248,In_1679);
or U9232 (N_9232,In_4265,In_4283);
and U9233 (N_9233,In_1560,In_2676);
or U9234 (N_9234,In_2651,In_1507);
xnor U9235 (N_9235,In_2778,In_3944);
or U9236 (N_9236,In_1190,In_3532);
xor U9237 (N_9237,In_1956,In_1053);
and U9238 (N_9238,In_4168,In_3644);
nand U9239 (N_9239,In_1209,In_4402);
nor U9240 (N_9240,In_2525,In_1188);
nor U9241 (N_9241,In_3788,In_285);
or U9242 (N_9242,In_3850,In_3584);
and U9243 (N_9243,In_471,In_1858);
or U9244 (N_9244,In_3300,In_3682);
or U9245 (N_9245,In_2207,In_2848);
xnor U9246 (N_9246,In_3033,In_4277);
nand U9247 (N_9247,In_3922,In_1618);
and U9248 (N_9248,In_4710,In_416);
nand U9249 (N_9249,In_2495,In_2902);
and U9250 (N_9250,In_3280,In_4498);
and U9251 (N_9251,In_3289,In_2225);
and U9252 (N_9252,In_318,In_694);
xnor U9253 (N_9253,In_1581,In_4347);
nand U9254 (N_9254,In_91,In_2090);
nor U9255 (N_9255,In_1215,In_1656);
xnor U9256 (N_9256,In_250,In_768);
nand U9257 (N_9257,In_1385,In_97);
xnor U9258 (N_9258,In_3071,In_1639);
xnor U9259 (N_9259,In_3122,In_4631);
nand U9260 (N_9260,In_1248,In_2987);
xnor U9261 (N_9261,In_3978,In_2626);
nand U9262 (N_9262,In_4946,In_259);
and U9263 (N_9263,In_138,In_4474);
nand U9264 (N_9264,In_2184,In_2650);
or U9265 (N_9265,In_4282,In_944);
xor U9266 (N_9266,In_487,In_1982);
or U9267 (N_9267,In_3818,In_952);
nand U9268 (N_9268,In_1144,In_3822);
or U9269 (N_9269,In_1461,In_1974);
xnor U9270 (N_9270,In_1996,In_3764);
or U9271 (N_9271,In_2024,In_363);
and U9272 (N_9272,In_4290,In_1691);
nor U9273 (N_9273,In_2179,In_678);
xnor U9274 (N_9274,In_4248,In_2622);
and U9275 (N_9275,In_673,In_4915);
and U9276 (N_9276,In_4816,In_3769);
nor U9277 (N_9277,In_1887,In_498);
and U9278 (N_9278,In_706,In_3577);
and U9279 (N_9279,In_2097,In_1403);
nor U9280 (N_9280,In_3112,In_2267);
or U9281 (N_9281,In_762,In_3127);
nand U9282 (N_9282,In_1820,In_2645);
nor U9283 (N_9283,In_4089,In_1573);
nor U9284 (N_9284,In_557,In_2541);
and U9285 (N_9285,In_3859,In_3055);
xnor U9286 (N_9286,In_3787,In_2973);
nor U9287 (N_9287,In_3165,In_4351);
xnor U9288 (N_9288,In_3536,In_2144);
xnor U9289 (N_9289,In_3078,In_3303);
xor U9290 (N_9290,In_1466,In_3630);
xnor U9291 (N_9291,In_3808,In_3048);
or U9292 (N_9292,In_3837,In_3925);
nand U9293 (N_9293,In_1512,In_4218);
nor U9294 (N_9294,In_4237,In_2171);
and U9295 (N_9295,In_2463,In_4569);
xnor U9296 (N_9296,In_1013,In_1313);
or U9297 (N_9297,In_4407,In_4890);
and U9298 (N_9298,In_490,In_471);
and U9299 (N_9299,In_3290,In_1848);
xnor U9300 (N_9300,In_1836,In_2552);
and U9301 (N_9301,In_3762,In_3787);
or U9302 (N_9302,In_2051,In_971);
nand U9303 (N_9303,In_2784,In_2296);
nor U9304 (N_9304,In_4495,In_2070);
and U9305 (N_9305,In_3273,In_4796);
nor U9306 (N_9306,In_1766,In_3187);
nor U9307 (N_9307,In_2246,In_2634);
or U9308 (N_9308,In_4211,In_901);
xor U9309 (N_9309,In_1512,In_3693);
nand U9310 (N_9310,In_1526,In_185);
nor U9311 (N_9311,In_3992,In_2848);
and U9312 (N_9312,In_3237,In_2293);
nand U9313 (N_9313,In_2176,In_664);
and U9314 (N_9314,In_849,In_704);
nor U9315 (N_9315,In_3369,In_4962);
nor U9316 (N_9316,In_3711,In_1280);
nor U9317 (N_9317,In_3817,In_4470);
xor U9318 (N_9318,In_1930,In_247);
and U9319 (N_9319,In_2472,In_109);
and U9320 (N_9320,In_3884,In_2286);
and U9321 (N_9321,In_1609,In_760);
and U9322 (N_9322,In_4485,In_4723);
xnor U9323 (N_9323,In_4936,In_2600);
nor U9324 (N_9324,In_156,In_3552);
nor U9325 (N_9325,In_994,In_3917);
nand U9326 (N_9326,In_199,In_500);
nand U9327 (N_9327,In_2056,In_1510);
and U9328 (N_9328,In_3951,In_1107);
and U9329 (N_9329,In_4670,In_4708);
xor U9330 (N_9330,In_4260,In_4002);
nor U9331 (N_9331,In_2826,In_2173);
nand U9332 (N_9332,In_685,In_2305);
or U9333 (N_9333,In_1586,In_1230);
nor U9334 (N_9334,In_2452,In_713);
nor U9335 (N_9335,In_1301,In_2812);
xor U9336 (N_9336,In_3512,In_626);
nand U9337 (N_9337,In_708,In_2413);
xnor U9338 (N_9338,In_650,In_3682);
nand U9339 (N_9339,In_176,In_1807);
or U9340 (N_9340,In_1985,In_548);
and U9341 (N_9341,In_4781,In_2993);
or U9342 (N_9342,In_1544,In_3841);
nor U9343 (N_9343,In_164,In_4122);
nor U9344 (N_9344,In_2225,In_285);
nor U9345 (N_9345,In_3640,In_2772);
nand U9346 (N_9346,In_3717,In_4385);
and U9347 (N_9347,In_1271,In_2780);
and U9348 (N_9348,In_1814,In_796);
nor U9349 (N_9349,In_4129,In_551);
nand U9350 (N_9350,In_3606,In_1669);
nor U9351 (N_9351,In_4626,In_4678);
nor U9352 (N_9352,In_1804,In_2865);
and U9353 (N_9353,In_210,In_1292);
or U9354 (N_9354,In_515,In_4669);
and U9355 (N_9355,In_3290,In_4191);
nor U9356 (N_9356,In_2684,In_3771);
and U9357 (N_9357,In_2252,In_2995);
or U9358 (N_9358,In_4984,In_3743);
nor U9359 (N_9359,In_3930,In_1712);
nand U9360 (N_9360,In_4018,In_4143);
or U9361 (N_9361,In_3523,In_3164);
nor U9362 (N_9362,In_81,In_1347);
or U9363 (N_9363,In_1100,In_1011);
nor U9364 (N_9364,In_2311,In_1586);
and U9365 (N_9365,In_4546,In_4542);
and U9366 (N_9366,In_2944,In_101);
and U9367 (N_9367,In_2559,In_927);
xnor U9368 (N_9368,In_4586,In_2320);
nand U9369 (N_9369,In_821,In_1876);
and U9370 (N_9370,In_3738,In_4109);
xor U9371 (N_9371,In_1822,In_1189);
nand U9372 (N_9372,In_3547,In_3742);
xnor U9373 (N_9373,In_3934,In_4003);
xor U9374 (N_9374,In_1120,In_4670);
or U9375 (N_9375,In_1147,In_2815);
nor U9376 (N_9376,In_1848,In_2055);
xor U9377 (N_9377,In_2810,In_1895);
nor U9378 (N_9378,In_3370,In_3389);
nand U9379 (N_9379,In_322,In_819);
nor U9380 (N_9380,In_4286,In_1635);
nand U9381 (N_9381,In_3367,In_3714);
and U9382 (N_9382,In_3510,In_3684);
xnor U9383 (N_9383,In_1044,In_2408);
or U9384 (N_9384,In_4435,In_147);
or U9385 (N_9385,In_809,In_1684);
or U9386 (N_9386,In_2749,In_4685);
nand U9387 (N_9387,In_2609,In_4530);
xor U9388 (N_9388,In_3055,In_4086);
nand U9389 (N_9389,In_1837,In_2137);
and U9390 (N_9390,In_606,In_1027);
nor U9391 (N_9391,In_2256,In_3090);
or U9392 (N_9392,In_1591,In_4988);
xnor U9393 (N_9393,In_4181,In_762);
nand U9394 (N_9394,In_4027,In_4506);
or U9395 (N_9395,In_4847,In_3607);
nand U9396 (N_9396,In_3096,In_346);
xnor U9397 (N_9397,In_4964,In_3665);
nor U9398 (N_9398,In_2075,In_821);
nand U9399 (N_9399,In_4695,In_3016);
nand U9400 (N_9400,In_3684,In_1743);
and U9401 (N_9401,In_4458,In_4308);
and U9402 (N_9402,In_2273,In_1757);
nand U9403 (N_9403,In_380,In_4972);
xnor U9404 (N_9404,In_4866,In_448);
nor U9405 (N_9405,In_2139,In_2317);
xor U9406 (N_9406,In_2617,In_4740);
xor U9407 (N_9407,In_3050,In_2222);
and U9408 (N_9408,In_2372,In_449);
nor U9409 (N_9409,In_2310,In_2897);
and U9410 (N_9410,In_1117,In_4363);
or U9411 (N_9411,In_2283,In_1178);
and U9412 (N_9412,In_2502,In_3945);
nor U9413 (N_9413,In_2777,In_2793);
and U9414 (N_9414,In_1028,In_2028);
and U9415 (N_9415,In_4218,In_4132);
or U9416 (N_9416,In_761,In_949);
xnor U9417 (N_9417,In_1951,In_2780);
nor U9418 (N_9418,In_2793,In_4500);
nand U9419 (N_9419,In_3609,In_2095);
nor U9420 (N_9420,In_2877,In_544);
or U9421 (N_9421,In_564,In_1679);
or U9422 (N_9422,In_1045,In_4961);
xnor U9423 (N_9423,In_4470,In_4770);
and U9424 (N_9424,In_3130,In_1161);
nor U9425 (N_9425,In_4486,In_628);
nor U9426 (N_9426,In_4411,In_4206);
and U9427 (N_9427,In_3980,In_1);
nand U9428 (N_9428,In_747,In_705);
nor U9429 (N_9429,In_691,In_996);
xnor U9430 (N_9430,In_3015,In_1030);
nand U9431 (N_9431,In_1074,In_1125);
nor U9432 (N_9432,In_1402,In_1077);
and U9433 (N_9433,In_1442,In_566);
nand U9434 (N_9434,In_3746,In_2088);
nor U9435 (N_9435,In_3847,In_2671);
nor U9436 (N_9436,In_2482,In_378);
or U9437 (N_9437,In_1493,In_3977);
nor U9438 (N_9438,In_2226,In_2974);
and U9439 (N_9439,In_2237,In_2738);
nor U9440 (N_9440,In_3154,In_678);
and U9441 (N_9441,In_1044,In_3458);
and U9442 (N_9442,In_304,In_4731);
or U9443 (N_9443,In_3043,In_1015);
nand U9444 (N_9444,In_160,In_4674);
nand U9445 (N_9445,In_2260,In_3314);
nand U9446 (N_9446,In_1566,In_4432);
or U9447 (N_9447,In_4582,In_1994);
and U9448 (N_9448,In_4173,In_4935);
nand U9449 (N_9449,In_4077,In_1532);
nor U9450 (N_9450,In_2768,In_3073);
nor U9451 (N_9451,In_455,In_2908);
or U9452 (N_9452,In_4968,In_1013);
and U9453 (N_9453,In_2987,In_3491);
xnor U9454 (N_9454,In_3158,In_3775);
and U9455 (N_9455,In_3738,In_4322);
nand U9456 (N_9456,In_1010,In_3091);
or U9457 (N_9457,In_2556,In_4421);
or U9458 (N_9458,In_3582,In_274);
nor U9459 (N_9459,In_3182,In_1384);
or U9460 (N_9460,In_3040,In_587);
nor U9461 (N_9461,In_3882,In_2707);
nand U9462 (N_9462,In_2497,In_2268);
xor U9463 (N_9463,In_2931,In_3207);
nor U9464 (N_9464,In_2216,In_4575);
xnor U9465 (N_9465,In_4210,In_1886);
xor U9466 (N_9466,In_52,In_4829);
and U9467 (N_9467,In_176,In_1190);
or U9468 (N_9468,In_3419,In_1779);
xnor U9469 (N_9469,In_3780,In_1378);
nor U9470 (N_9470,In_4190,In_248);
nor U9471 (N_9471,In_781,In_1228);
xor U9472 (N_9472,In_3236,In_180);
or U9473 (N_9473,In_4402,In_1712);
nand U9474 (N_9474,In_744,In_1565);
nand U9475 (N_9475,In_2906,In_4761);
and U9476 (N_9476,In_154,In_2705);
xnor U9477 (N_9477,In_79,In_2943);
or U9478 (N_9478,In_3262,In_2139);
nor U9479 (N_9479,In_141,In_1942);
xnor U9480 (N_9480,In_3833,In_739);
xnor U9481 (N_9481,In_2259,In_4112);
nor U9482 (N_9482,In_3619,In_4006);
or U9483 (N_9483,In_3523,In_2887);
xor U9484 (N_9484,In_3830,In_200);
and U9485 (N_9485,In_1982,In_2100);
nor U9486 (N_9486,In_2067,In_4830);
or U9487 (N_9487,In_2397,In_1789);
nor U9488 (N_9488,In_4783,In_2319);
nand U9489 (N_9489,In_455,In_1995);
or U9490 (N_9490,In_4302,In_4090);
and U9491 (N_9491,In_3851,In_1830);
or U9492 (N_9492,In_2098,In_4369);
or U9493 (N_9493,In_341,In_2607);
xnor U9494 (N_9494,In_4187,In_2051);
xor U9495 (N_9495,In_3568,In_4779);
nor U9496 (N_9496,In_3110,In_3136);
and U9497 (N_9497,In_3848,In_4481);
nor U9498 (N_9498,In_3737,In_440);
or U9499 (N_9499,In_3356,In_2575);
xnor U9500 (N_9500,In_2295,In_1522);
nand U9501 (N_9501,In_3207,In_3593);
nor U9502 (N_9502,In_1833,In_3428);
and U9503 (N_9503,In_529,In_4296);
and U9504 (N_9504,In_21,In_429);
or U9505 (N_9505,In_3470,In_1324);
or U9506 (N_9506,In_4698,In_2962);
or U9507 (N_9507,In_3220,In_232);
xor U9508 (N_9508,In_984,In_3248);
nor U9509 (N_9509,In_376,In_3173);
nand U9510 (N_9510,In_2086,In_681);
nor U9511 (N_9511,In_3429,In_4363);
and U9512 (N_9512,In_2669,In_31);
xnor U9513 (N_9513,In_644,In_4626);
and U9514 (N_9514,In_3220,In_1671);
and U9515 (N_9515,In_1349,In_2182);
or U9516 (N_9516,In_172,In_2116);
xor U9517 (N_9517,In_2041,In_1132);
and U9518 (N_9518,In_2235,In_885);
and U9519 (N_9519,In_3211,In_4966);
or U9520 (N_9520,In_3556,In_4524);
nand U9521 (N_9521,In_2462,In_1132);
nor U9522 (N_9522,In_3439,In_4835);
or U9523 (N_9523,In_4328,In_3705);
nand U9524 (N_9524,In_2257,In_1800);
xor U9525 (N_9525,In_3421,In_2099);
and U9526 (N_9526,In_2489,In_810);
and U9527 (N_9527,In_4073,In_2158);
nand U9528 (N_9528,In_4505,In_701);
nor U9529 (N_9529,In_4251,In_4404);
nand U9530 (N_9530,In_1320,In_1398);
nor U9531 (N_9531,In_3312,In_2361);
nor U9532 (N_9532,In_2274,In_3555);
xor U9533 (N_9533,In_2757,In_1339);
nor U9534 (N_9534,In_3332,In_3634);
nand U9535 (N_9535,In_3802,In_2305);
and U9536 (N_9536,In_616,In_1754);
xor U9537 (N_9537,In_701,In_2462);
and U9538 (N_9538,In_3159,In_2021);
nor U9539 (N_9539,In_2027,In_1581);
nand U9540 (N_9540,In_2240,In_796);
or U9541 (N_9541,In_3460,In_1332);
xnor U9542 (N_9542,In_4303,In_4761);
or U9543 (N_9543,In_2113,In_1937);
nand U9544 (N_9544,In_2932,In_1444);
and U9545 (N_9545,In_805,In_2287);
nand U9546 (N_9546,In_3538,In_199);
xnor U9547 (N_9547,In_3832,In_1711);
nand U9548 (N_9548,In_2691,In_1016);
nand U9549 (N_9549,In_4109,In_689);
nand U9550 (N_9550,In_2050,In_3415);
xnor U9551 (N_9551,In_4384,In_2362);
and U9552 (N_9552,In_4230,In_3362);
nand U9553 (N_9553,In_2334,In_4237);
nor U9554 (N_9554,In_3174,In_4224);
xor U9555 (N_9555,In_4040,In_2215);
and U9556 (N_9556,In_450,In_2260);
and U9557 (N_9557,In_2429,In_4574);
nand U9558 (N_9558,In_4548,In_454);
nor U9559 (N_9559,In_2150,In_2835);
nand U9560 (N_9560,In_661,In_303);
nor U9561 (N_9561,In_3141,In_1239);
and U9562 (N_9562,In_1489,In_1052);
or U9563 (N_9563,In_2238,In_1776);
nand U9564 (N_9564,In_1845,In_2594);
xor U9565 (N_9565,In_150,In_4153);
and U9566 (N_9566,In_1927,In_2291);
or U9567 (N_9567,In_536,In_4253);
xor U9568 (N_9568,In_2353,In_1375);
or U9569 (N_9569,In_1675,In_3468);
and U9570 (N_9570,In_4031,In_4444);
nor U9571 (N_9571,In_4576,In_789);
xnor U9572 (N_9572,In_900,In_1749);
nand U9573 (N_9573,In_379,In_991);
nor U9574 (N_9574,In_4325,In_3740);
or U9575 (N_9575,In_41,In_1623);
and U9576 (N_9576,In_2024,In_1335);
or U9577 (N_9577,In_1701,In_2627);
nor U9578 (N_9578,In_243,In_3080);
xor U9579 (N_9579,In_2524,In_1090);
nor U9580 (N_9580,In_2047,In_2488);
or U9581 (N_9581,In_371,In_1170);
and U9582 (N_9582,In_4025,In_2465);
and U9583 (N_9583,In_3073,In_1731);
nand U9584 (N_9584,In_189,In_1674);
nor U9585 (N_9585,In_756,In_4590);
xor U9586 (N_9586,In_214,In_2779);
or U9587 (N_9587,In_2379,In_4427);
nand U9588 (N_9588,In_1692,In_4905);
nand U9589 (N_9589,In_4376,In_4145);
nand U9590 (N_9590,In_2878,In_345);
and U9591 (N_9591,In_2386,In_841);
nor U9592 (N_9592,In_4712,In_3983);
or U9593 (N_9593,In_1936,In_1988);
nor U9594 (N_9594,In_261,In_1997);
nand U9595 (N_9595,In_4217,In_3451);
xnor U9596 (N_9596,In_3203,In_3510);
or U9597 (N_9597,In_1010,In_4762);
or U9598 (N_9598,In_1803,In_2779);
and U9599 (N_9599,In_4197,In_1025);
and U9600 (N_9600,In_1865,In_4950);
and U9601 (N_9601,In_3691,In_3750);
xnor U9602 (N_9602,In_4475,In_1466);
nand U9603 (N_9603,In_1684,In_4526);
nor U9604 (N_9604,In_2979,In_2703);
and U9605 (N_9605,In_1040,In_4949);
nand U9606 (N_9606,In_387,In_1702);
xnor U9607 (N_9607,In_3684,In_3271);
xor U9608 (N_9608,In_303,In_1670);
xor U9609 (N_9609,In_2356,In_3844);
nor U9610 (N_9610,In_2810,In_3330);
nor U9611 (N_9611,In_3032,In_2956);
nand U9612 (N_9612,In_4069,In_410);
or U9613 (N_9613,In_1509,In_3320);
xor U9614 (N_9614,In_189,In_1380);
and U9615 (N_9615,In_2499,In_2259);
nand U9616 (N_9616,In_2276,In_1997);
or U9617 (N_9617,In_1419,In_3327);
or U9618 (N_9618,In_1880,In_203);
and U9619 (N_9619,In_2898,In_3992);
or U9620 (N_9620,In_2702,In_4356);
nand U9621 (N_9621,In_1928,In_140);
nand U9622 (N_9622,In_1172,In_1604);
xor U9623 (N_9623,In_2822,In_3931);
xor U9624 (N_9624,In_4044,In_4703);
nand U9625 (N_9625,In_1857,In_2822);
nor U9626 (N_9626,In_4533,In_1322);
xnor U9627 (N_9627,In_3284,In_1555);
nor U9628 (N_9628,In_2727,In_1093);
nand U9629 (N_9629,In_3818,In_4914);
xor U9630 (N_9630,In_3915,In_2285);
and U9631 (N_9631,In_2240,In_1734);
xnor U9632 (N_9632,In_4072,In_1112);
nor U9633 (N_9633,In_2019,In_2329);
and U9634 (N_9634,In_4440,In_1888);
or U9635 (N_9635,In_792,In_4398);
nor U9636 (N_9636,In_570,In_431);
nor U9637 (N_9637,In_32,In_747);
and U9638 (N_9638,In_2682,In_1105);
and U9639 (N_9639,In_3636,In_174);
xor U9640 (N_9640,In_582,In_673);
xnor U9641 (N_9641,In_3935,In_351);
nand U9642 (N_9642,In_3796,In_4295);
nand U9643 (N_9643,In_40,In_1764);
or U9644 (N_9644,In_2755,In_4921);
xor U9645 (N_9645,In_3082,In_3162);
or U9646 (N_9646,In_4028,In_407);
nor U9647 (N_9647,In_136,In_1649);
and U9648 (N_9648,In_4217,In_3231);
xnor U9649 (N_9649,In_2180,In_1806);
xnor U9650 (N_9650,In_3275,In_2927);
nor U9651 (N_9651,In_287,In_968);
xnor U9652 (N_9652,In_3846,In_573);
and U9653 (N_9653,In_3800,In_1356);
nand U9654 (N_9654,In_4990,In_228);
xor U9655 (N_9655,In_2846,In_4106);
xor U9656 (N_9656,In_3299,In_3483);
and U9657 (N_9657,In_4048,In_1750);
xor U9658 (N_9658,In_1770,In_2787);
nor U9659 (N_9659,In_2786,In_1818);
or U9660 (N_9660,In_3654,In_1952);
and U9661 (N_9661,In_4218,In_1951);
and U9662 (N_9662,In_1041,In_3739);
xor U9663 (N_9663,In_1669,In_2839);
and U9664 (N_9664,In_1800,In_1537);
nor U9665 (N_9665,In_672,In_4163);
nor U9666 (N_9666,In_3550,In_402);
nand U9667 (N_9667,In_1457,In_3277);
and U9668 (N_9668,In_3613,In_3051);
or U9669 (N_9669,In_4297,In_245);
nand U9670 (N_9670,In_1880,In_4106);
nor U9671 (N_9671,In_3102,In_4672);
nand U9672 (N_9672,In_504,In_3836);
and U9673 (N_9673,In_1908,In_2316);
or U9674 (N_9674,In_3960,In_113);
nor U9675 (N_9675,In_1236,In_3949);
nand U9676 (N_9676,In_2751,In_3886);
nand U9677 (N_9677,In_4553,In_149);
and U9678 (N_9678,In_4248,In_4870);
and U9679 (N_9679,In_1405,In_3048);
xnor U9680 (N_9680,In_3322,In_2018);
nand U9681 (N_9681,In_4901,In_2586);
or U9682 (N_9682,In_549,In_3576);
and U9683 (N_9683,In_3521,In_4109);
nor U9684 (N_9684,In_116,In_1855);
and U9685 (N_9685,In_1009,In_2644);
nor U9686 (N_9686,In_4491,In_1204);
xor U9687 (N_9687,In_937,In_2052);
and U9688 (N_9688,In_4760,In_1323);
nor U9689 (N_9689,In_83,In_3273);
nor U9690 (N_9690,In_3407,In_3023);
xnor U9691 (N_9691,In_3580,In_3464);
nor U9692 (N_9692,In_1035,In_3212);
nor U9693 (N_9693,In_3750,In_1837);
nor U9694 (N_9694,In_1410,In_694);
nand U9695 (N_9695,In_2900,In_4456);
nor U9696 (N_9696,In_1331,In_2423);
nand U9697 (N_9697,In_1071,In_887);
and U9698 (N_9698,In_3849,In_2256);
xnor U9699 (N_9699,In_1003,In_916);
nand U9700 (N_9700,In_3636,In_2523);
and U9701 (N_9701,In_4381,In_1889);
nand U9702 (N_9702,In_4089,In_951);
nand U9703 (N_9703,In_2487,In_795);
xor U9704 (N_9704,In_1239,In_1079);
xnor U9705 (N_9705,In_1926,In_4632);
and U9706 (N_9706,In_3478,In_4112);
nand U9707 (N_9707,In_2884,In_3536);
xnor U9708 (N_9708,In_882,In_2223);
or U9709 (N_9709,In_2832,In_2821);
and U9710 (N_9710,In_1041,In_955);
nand U9711 (N_9711,In_455,In_388);
nor U9712 (N_9712,In_412,In_4804);
nor U9713 (N_9713,In_1291,In_3180);
nand U9714 (N_9714,In_1875,In_2802);
xor U9715 (N_9715,In_2403,In_1560);
nor U9716 (N_9716,In_2781,In_687);
nor U9717 (N_9717,In_4372,In_787);
nor U9718 (N_9718,In_3274,In_280);
nand U9719 (N_9719,In_71,In_1798);
and U9720 (N_9720,In_4071,In_3934);
nor U9721 (N_9721,In_2941,In_2789);
nor U9722 (N_9722,In_4361,In_4438);
nand U9723 (N_9723,In_3828,In_876);
or U9724 (N_9724,In_789,In_358);
xnor U9725 (N_9725,In_160,In_1725);
or U9726 (N_9726,In_3170,In_1741);
nand U9727 (N_9727,In_3788,In_1972);
xnor U9728 (N_9728,In_1222,In_2498);
nor U9729 (N_9729,In_1382,In_3373);
nor U9730 (N_9730,In_3034,In_4259);
xnor U9731 (N_9731,In_4473,In_93);
nor U9732 (N_9732,In_1393,In_4901);
nor U9733 (N_9733,In_2775,In_3372);
xnor U9734 (N_9734,In_4802,In_1531);
nand U9735 (N_9735,In_2178,In_2430);
or U9736 (N_9736,In_768,In_2124);
xnor U9737 (N_9737,In_2575,In_2771);
or U9738 (N_9738,In_2429,In_4291);
or U9739 (N_9739,In_1616,In_402);
nand U9740 (N_9740,In_402,In_1183);
or U9741 (N_9741,In_2694,In_2063);
or U9742 (N_9742,In_294,In_3343);
xor U9743 (N_9743,In_716,In_2859);
nand U9744 (N_9744,In_3556,In_2126);
nor U9745 (N_9745,In_3465,In_393);
xnor U9746 (N_9746,In_2297,In_2087);
xnor U9747 (N_9747,In_2200,In_37);
or U9748 (N_9748,In_1263,In_4192);
or U9749 (N_9749,In_2078,In_2606);
and U9750 (N_9750,In_2921,In_1783);
nor U9751 (N_9751,In_233,In_1516);
nor U9752 (N_9752,In_4689,In_9);
nand U9753 (N_9753,In_3893,In_4337);
nand U9754 (N_9754,In_1100,In_773);
xnor U9755 (N_9755,In_2780,In_437);
xor U9756 (N_9756,In_4817,In_4842);
or U9757 (N_9757,In_1731,In_2578);
or U9758 (N_9758,In_77,In_3507);
xor U9759 (N_9759,In_930,In_4918);
and U9760 (N_9760,In_3526,In_707);
or U9761 (N_9761,In_2789,In_1784);
nand U9762 (N_9762,In_3333,In_1925);
or U9763 (N_9763,In_7,In_1833);
nand U9764 (N_9764,In_372,In_1707);
or U9765 (N_9765,In_2984,In_807);
nand U9766 (N_9766,In_4032,In_1813);
or U9767 (N_9767,In_1748,In_1427);
nor U9768 (N_9768,In_4827,In_4418);
xor U9769 (N_9769,In_2785,In_3348);
xnor U9770 (N_9770,In_1225,In_69);
nor U9771 (N_9771,In_4370,In_1822);
or U9772 (N_9772,In_664,In_2177);
xnor U9773 (N_9773,In_2536,In_255);
nor U9774 (N_9774,In_172,In_3606);
xor U9775 (N_9775,In_101,In_3362);
or U9776 (N_9776,In_3252,In_4561);
and U9777 (N_9777,In_3737,In_4406);
and U9778 (N_9778,In_3571,In_4712);
nand U9779 (N_9779,In_653,In_2742);
nor U9780 (N_9780,In_1000,In_3690);
nand U9781 (N_9781,In_4332,In_554);
and U9782 (N_9782,In_1543,In_3345);
or U9783 (N_9783,In_4245,In_3442);
nor U9784 (N_9784,In_2730,In_1795);
and U9785 (N_9785,In_2103,In_2228);
or U9786 (N_9786,In_4585,In_3262);
xor U9787 (N_9787,In_1685,In_3621);
or U9788 (N_9788,In_704,In_2936);
or U9789 (N_9789,In_3314,In_487);
and U9790 (N_9790,In_616,In_3384);
xnor U9791 (N_9791,In_4482,In_998);
nand U9792 (N_9792,In_1364,In_1491);
nand U9793 (N_9793,In_4032,In_2361);
or U9794 (N_9794,In_166,In_845);
or U9795 (N_9795,In_3048,In_4609);
and U9796 (N_9796,In_3097,In_1359);
or U9797 (N_9797,In_2054,In_3634);
xnor U9798 (N_9798,In_979,In_2581);
nand U9799 (N_9799,In_3971,In_3619);
and U9800 (N_9800,In_972,In_761);
xnor U9801 (N_9801,In_2259,In_4287);
and U9802 (N_9802,In_523,In_3811);
nor U9803 (N_9803,In_2518,In_3072);
nand U9804 (N_9804,In_1369,In_2663);
or U9805 (N_9805,In_110,In_4510);
and U9806 (N_9806,In_3929,In_2134);
nand U9807 (N_9807,In_4443,In_1185);
xor U9808 (N_9808,In_2087,In_3750);
nor U9809 (N_9809,In_2244,In_4311);
or U9810 (N_9810,In_4955,In_669);
or U9811 (N_9811,In_36,In_3739);
nand U9812 (N_9812,In_2091,In_4578);
nand U9813 (N_9813,In_355,In_3598);
nor U9814 (N_9814,In_35,In_2621);
and U9815 (N_9815,In_466,In_2855);
and U9816 (N_9816,In_1676,In_4825);
nand U9817 (N_9817,In_3937,In_3583);
xnor U9818 (N_9818,In_2859,In_523);
and U9819 (N_9819,In_1690,In_4274);
or U9820 (N_9820,In_3848,In_4651);
or U9821 (N_9821,In_880,In_4118);
nor U9822 (N_9822,In_3782,In_3754);
or U9823 (N_9823,In_355,In_69);
or U9824 (N_9824,In_3521,In_125);
nand U9825 (N_9825,In_3381,In_3342);
nand U9826 (N_9826,In_2434,In_1610);
nand U9827 (N_9827,In_4077,In_2755);
xnor U9828 (N_9828,In_1212,In_2229);
xor U9829 (N_9829,In_2586,In_1542);
and U9830 (N_9830,In_4992,In_4886);
or U9831 (N_9831,In_4035,In_2102);
or U9832 (N_9832,In_1659,In_1451);
or U9833 (N_9833,In_291,In_1109);
xnor U9834 (N_9834,In_1542,In_2313);
nand U9835 (N_9835,In_2130,In_1981);
or U9836 (N_9836,In_851,In_3570);
xnor U9837 (N_9837,In_628,In_3950);
and U9838 (N_9838,In_2082,In_4411);
nor U9839 (N_9839,In_3430,In_18);
xnor U9840 (N_9840,In_1779,In_4605);
and U9841 (N_9841,In_4633,In_4257);
nand U9842 (N_9842,In_1121,In_4667);
and U9843 (N_9843,In_4876,In_2014);
or U9844 (N_9844,In_1927,In_2486);
and U9845 (N_9845,In_2089,In_3521);
xnor U9846 (N_9846,In_2485,In_2467);
xnor U9847 (N_9847,In_1114,In_3734);
xor U9848 (N_9848,In_4432,In_1373);
nor U9849 (N_9849,In_4391,In_2974);
or U9850 (N_9850,In_4620,In_3836);
nand U9851 (N_9851,In_2909,In_3066);
nand U9852 (N_9852,In_235,In_2721);
or U9853 (N_9853,In_2557,In_3187);
or U9854 (N_9854,In_41,In_2894);
nand U9855 (N_9855,In_1781,In_2302);
xnor U9856 (N_9856,In_4516,In_72);
nand U9857 (N_9857,In_2368,In_438);
xor U9858 (N_9858,In_1768,In_3071);
nand U9859 (N_9859,In_2007,In_593);
nand U9860 (N_9860,In_333,In_2888);
nand U9861 (N_9861,In_256,In_4768);
nor U9862 (N_9862,In_639,In_1144);
or U9863 (N_9863,In_1604,In_4799);
and U9864 (N_9864,In_4520,In_2009);
xor U9865 (N_9865,In_956,In_2649);
and U9866 (N_9866,In_842,In_4487);
xnor U9867 (N_9867,In_318,In_408);
xor U9868 (N_9868,In_3407,In_2493);
and U9869 (N_9869,In_2803,In_79);
nand U9870 (N_9870,In_3254,In_1142);
or U9871 (N_9871,In_4957,In_3976);
or U9872 (N_9872,In_2931,In_2805);
nor U9873 (N_9873,In_2350,In_96);
xnor U9874 (N_9874,In_4377,In_1490);
nand U9875 (N_9875,In_424,In_86);
nand U9876 (N_9876,In_2319,In_4817);
xor U9877 (N_9877,In_848,In_3174);
nand U9878 (N_9878,In_3313,In_1062);
nand U9879 (N_9879,In_2517,In_3258);
and U9880 (N_9880,In_1982,In_4416);
or U9881 (N_9881,In_956,In_263);
xnor U9882 (N_9882,In_2527,In_4312);
and U9883 (N_9883,In_1144,In_1298);
nand U9884 (N_9884,In_4077,In_1708);
and U9885 (N_9885,In_4102,In_280);
nor U9886 (N_9886,In_3279,In_3133);
nand U9887 (N_9887,In_3024,In_4767);
and U9888 (N_9888,In_981,In_4843);
nor U9889 (N_9889,In_4905,In_1287);
and U9890 (N_9890,In_4823,In_2085);
nor U9891 (N_9891,In_2861,In_1457);
and U9892 (N_9892,In_661,In_4164);
and U9893 (N_9893,In_1679,In_4900);
nand U9894 (N_9894,In_2486,In_1940);
xor U9895 (N_9895,In_1064,In_314);
nor U9896 (N_9896,In_2983,In_3893);
or U9897 (N_9897,In_199,In_941);
nor U9898 (N_9898,In_988,In_439);
nor U9899 (N_9899,In_3947,In_232);
and U9900 (N_9900,In_1168,In_3911);
and U9901 (N_9901,In_3133,In_3910);
nor U9902 (N_9902,In_2700,In_1383);
nand U9903 (N_9903,In_428,In_135);
or U9904 (N_9904,In_772,In_1505);
nor U9905 (N_9905,In_3421,In_1131);
nor U9906 (N_9906,In_4985,In_1614);
and U9907 (N_9907,In_561,In_2401);
nor U9908 (N_9908,In_1820,In_4772);
nor U9909 (N_9909,In_1294,In_4855);
or U9910 (N_9910,In_493,In_3241);
xnor U9911 (N_9911,In_1452,In_1316);
and U9912 (N_9912,In_3863,In_1984);
and U9913 (N_9913,In_1525,In_4110);
nand U9914 (N_9914,In_4756,In_4777);
xnor U9915 (N_9915,In_2837,In_4083);
or U9916 (N_9916,In_250,In_3235);
and U9917 (N_9917,In_4097,In_4276);
and U9918 (N_9918,In_2548,In_1026);
nor U9919 (N_9919,In_3410,In_47);
nor U9920 (N_9920,In_3077,In_1383);
xor U9921 (N_9921,In_4335,In_4744);
xor U9922 (N_9922,In_4653,In_1939);
xor U9923 (N_9923,In_3081,In_1485);
and U9924 (N_9924,In_1357,In_3327);
or U9925 (N_9925,In_2713,In_3038);
xnor U9926 (N_9926,In_1518,In_111);
and U9927 (N_9927,In_3075,In_3747);
nor U9928 (N_9928,In_1788,In_3386);
nor U9929 (N_9929,In_4,In_743);
nor U9930 (N_9930,In_2082,In_3600);
xor U9931 (N_9931,In_2772,In_947);
and U9932 (N_9932,In_3713,In_168);
or U9933 (N_9933,In_868,In_246);
or U9934 (N_9934,In_3903,In_3990);
and U9935 (N_9935,In_4091,In_3405);
nor U9936 (N_9936,In_4786,In_3040);
nor U9937 (N_9937,In_4157,In_2934);
xor U9938 (N_9938,In_2566,In_4956);
xor U9939 (N_9939,In_300,In_648);
nor U9940 (N_9940,In_4498,In_2481);
xnor U9941 (N_9941,In_3814,In_1943);
or U9942 (N_9942,In_1211,In_4508);
or U9943 (N_9943,In_1621,In_2685);
and U9944 (N_9944,In_3595,In_4993);
or U9945 (N_9945,In_3813,In_3963);
nand U9946 (N_9946,In_2159,In_3910);
and U9947 (N_9947,In_2098,In_540);
xor U9948 (N_9948,In_1770,In_1578);
and U9949 (N_9949,In_735,In_2500);
nor U9950 (N_9950,In_3127,In_4457);
xor U9951 (N_9951,In_757,In_2610);
xor U9952 (N_9952,In_4743,In_2338);
nand U9953 (N_9953,In_4124,In_3998);
nor U9954 (N_9954,In_247,In_4907);
nand U9955 (N_9955,In_3612,In_944);
nor U9956 (N_9956,In_1434,In_608);
and U9957 (N_9957,In_2221,In_2397);
nand U9958 (N_9958,In_2273,In_2639);
xnor U9959 (N_9959,In_1926,In_879);
nor U9960 (N_9960,In_113,In_96);
nand U9961 (N_9961,In_1666,In_4581);
and U9962 (N_9962,In_1813,In_990);
and U9963 (N_9963,In_2031,In_773);
nor U9964 (N_9964,In_4336,In_1590);
and U9965 (N_9965,In_3600,In_3366);
or U9966 (N_9966,In_3777,In_1405);
xnor U9967 (N_9967,In_3125,In_1099);
nor U9968 (N_9968,In_2859,In_1414);
or U9969 (N_9969,In_2389,In_2617);
xnor U9970 (N_9970,In_1558,In_3381);
xor U9971 (N_9971,In_972,In_3595);
nor U9972 (N_9972,In_315,In_4887);
and U9973 (N_9973,In_1412,In_873);
nor U9974 (N_9974,In_4898,In_493);
nand U9975 (N_9975,In_2045,In_2211);
xor U9976 (N_9976,In_1166,In_4565);
and U9977 (N_9977,In_4452,In_1583);
and U9978 (N_9978,In_456,In_2788);
nor U9979 (N_9979,In_72,In_1958);
nand U9980 (N_9980,In_3345,In_4939);
or U9981 (N_9981,In_692,In_567);
xor U9982 (N_9982,In_2245,In_4081);
nor U9983 (N_9983,In_1539,In_4930);
or U9984 (N_9984,In_2332,In_82);
nand U9985 (N_9985,In_3636,In_2725);
and U9986 (N_9986,In_4,In_3327);
nand U9987 (N_9987,In_561,In_1745);
and U9988 (N_9988,In_4233,In_1720);
xor U9989 (N_9989,In_4261,In_4207);
nand U9990 (N_9990,In_1758,In_170);
xnor U9991 (N_9991,In_4770,In_243);
nor U9992 (N_9992,In_1021,In_2998);
xnor U9993 (N_9993,In_1226,In_2987);
nor U9994 (N_9994,In_253,In_2416);
and U9995 (N_9995,In_2325,In_1348);
xnor U9996 (N_9996,In_1942,In_2774);
xnor U9997 (N_9997,In_4814,In_1877);
and U9998 (N_9998,In_1590,In_2204);
xnor U9999 (N_9999,In_1111,In_2861);
xor U10000 (N_10000,N_8666,N_2824);
xor U10001 (N_10001,N_1472,N_560);
nor U10002 (N_10002,N_4684,N_3347);
nand U10003 (N_10003,N_9838,N_6653);
nor U10004 (N_10004,N_4821,N_5627);
nor U10005 (N_10005,N_8024,N_4789);
nand U10006 (N_10006,N_2041,N_9631);
nor U10007 (N_10007,N_2019,N_6264);
xor U10008 (N_10008,N_22,N_5366);
xnor U10009 (N_10009,N_68,N_1349);
and U10010 (N_10010,N_2459,N_8547);
nor U10011 (N_10011,N_1070,N_5617);
and U10012 (N_10012,N_7444,N_8139);
nand U10013 (N_10013,N_4553,N_925);
or U10014 (N_10014,N_1375,N_1872);
xor U10015 (N_10015,N_1583,N_6925);
or U10016 (N_10016,N_9536,N_6707);
nor U10017 (N_10017,N_7378,N_4763);
or U10018 (N_10018,N_4510,N_5116);
nand U10019 (N_10019,N_7916,N_4425);
and U10020 (N_10020,N_2515,N_4879);
nand U10021 (N_10021,N_4209,N_6050);
nor U10022 (N_10022,N_6260,N_3812);
nand U10023 (N_10023,N_8534,N_1367);
and U10024 (N_10024,N_5289,N_8975);
nor U10025 (N_10025,N_6440,N_4693);
nor U10026 (N_10026,N_1193,N_7415);
xor U10027 (N_10027,N_2032,N_578);
nor U10028 (N_10028,N_1262,N_5471);
nor U10029 (N_10029,N_9343,N_5602);
and U10030 (N_10030,N_7447,N_9914);
nor U10031 (N_10031,N_9622,N_9367);
and U10032 (N_10032,N_533,N_4195);
and U10033 (N_10033,N_1686,N_1157);
nor U10034 (N_10034,N_3071,N_6762);
xor U10035 (N_10035,N_4216,N_3711);
nor U10036 (N_10036,N_6827,N_640);
nand U10037 (N_10037,N_7702,N_2373);
nor U10038 (N_10038,N_8744,N_4492);
and U10039 (N_10039,N_4458,N_2577);
nor U10040 (N_10040,N_8508,N_5914);
nor U10041 (N_10041,N_2859,N_2760);
nand U10042 (N_10042,N_2930,N_9964);
nor U10043 (N_10043,N_9112,N_122);
nor U10044 (N_10044,N_7403,N_4728);
or U10045 (N_10045,N_9886,N_6811);
or U10046 (N_10046,N_1998,N_6730);
and U10047 (N_10047,N_882,N_1425);
or U10048 (N_10048,N_7874,N_7383);
xnor U10049 (N_10049,N_9907,N_6108);
xor U10050 (N_10050,N_7362,N_1544);
and U10051 (N_10051,N_2180,N_4992);
nand U10052 (N_10052,N_4121,N_1230);
or U10053 (N_10053,N_945,N_6324);
nand U10054 (N_10054,N_5944,N_9023);
nand U10055 (N_10055,N_6518,N_9911);
and U10056 (N_10056,N_348,N_6939);
or U10057 (N_10057,N_6763,N_6540);
xnor U10058 (N_10058,N_9065,N_2454);
nand U10059 (N_10059,N_8442,N_6174);
nor U10060 (N_10060,N_5248,N_853);
nand U10061 (N_10061,N_2876,N_3140);
nor U10062 (N_10062,N_2249,N_4165);
nand U10063 (N_10063,N_4945,N_5579);
nand U10064 (N_10064,N_7513,N_6997);
nand U10065 (N_10065,N_6897,N_3519);
or U10066 (N_10066,N_6513,N_2755);
and U10067 (N_10067,N_4241,N_8610);
nor U10068 (N_10068,N_5113,N_105);
xor U10069 (N_10069,N_6726,N_1669);
xor U10070 (N_10070,N_1077,N_10);
nor U10071 (N_10071,N_1996,N_6494);
xor U10072 (N_10072,N_8571,N_2523);
nand U10073 (N_10073,N_1296,N_1018);
or U10074 (N_10074,N_8774,N_7878);
and U10075 (N_10075,N_8363,N_9649);
nor U10076 (N_10076,N_2214,N_2410);
xor U10077 (N_10077,N_4322,N_7186);
and U10078 (N_10078,N_4137,N_6296);
nand U10079 (N_10079,N_4466,N_3075);
nand U10080 (N_10080,N_9916,N_2724);
xor U10081 (N_10081,N_2217,N_7262);
xor U10082 (N_10082,N_4975,N_2204);
xnor U10083 (N_10083,N_7117,N_4974);
nand U10084 (N_10084,N_2420,N_1129);
or U10085 (N_10085,N_553,N_933);
and U10086 (N_10086,N_6477,N_4520);
and U10087 (N_10087,N_417,N_1209);
or U10088 (N_10088,N_7714,N_9475);
xor U10089 (N_10089,N_2589,N_8236);
or U10090 (N_10090,N_5708,N_1338);
nand U10091 (N_10091,N_8423,N_6035);
xor U10092 (N_10092,N_9963,N_9304);
and U10093 (N_10093,N_9761,N_5588);
and U10094 (N_10094,N_5110,N_1920);
nand U10095 (N_10095,N_7073,N_7161);
nand U10096 (N_10096,N_3356,N_3489);
or U10097 (N_10097,N_2132,N_1706);
nor U10098 (N_10098,N_756,N_9194);
or U10099 (N_10099,N_3614,N_5851);
and U10100 (N_10100,N_8295,N_5041);
nand U10101 (N_10101,N_7264,N_4762);
and U10102 (N_10102,N_6369,N_9881);
or U10103 (N_10103,N_644,N_8844);
xor U10104 (N_10104,N_5845,N_9091);
and U10105 (N_10105,N_2475,N_2511);
xor U10106 (N_10106,N_7409,N_5250);
xnor U10107 (N_10107,N_1092,N_4430);
and U10108 (N_10108,N_1903,N_6013);
xor U10109 (N_10109,N_5312,N_3522);
or U10110 (N_10110,N_8581,N_216);
or U10111 (N_10111,N_8014,N_725);
xor U10112 (N_10112,N_3194,N_7826);
xor U10113 (N_10113,N_7341,N_3463);
nor U10114 (N_10114,N_155,N_9311);
nor U10115 (N_10115,N_3192,N_947);
nor U10116 (N_10116,N_8316,N_5799);
nor U10117 (N_10117,N_4387,N_7405);
or U10118 (N_10118,N_9902,N_5216);
or U10119 (N_10119,N_9987,N_1401);
and U10120 (N_10120,N_2654,N_5885);
xor U10121 (N_10121,N_8560,N_7480);
and U10122 (N_10122,N_9181,N_149);
xor U10123 (N_10123,N_2281,N_6219);
nor U10124 (N_10124,N_7519,N_3820);
nor U10125 (N_10125,N_3716,N_8269);
nor U10126 (N_10126,N_8957,N_2178);
nand U10127 (N_10127,N_4905,N_6556);
and U10128 (N_10128,N_845,N_7210);
xor U10129 (N_10129,N_4550,N_9206);
nor U10130 (N_10130,N_3034,N_726);
nor U10131 (N_10131,N_4408,N_613);
nor U10132 (N_10132,N_195,N_8186);
nor U10133 (N_10133,N_5083,N_5576);
xnor U10134 (N_10134,N_4120,N_9732);
and U10135 (N_10135,N_7943,N_6887);
nand U10136 (N_10136,N_557,N_3435);
nand U10137 (N_10137,N_4705,N_3019);
xor U10138 (N_10138,N_113,N_939);
and U10139 (N_10139,N_9388,N_4254);
or U10140 (N_10140,N_6251,N_7274);
and U10141 (N_10141,N_2208,N_5526);
nand U10142 (N_10142,N_7317,N_3022);
and U10143 (N_10143,N_5912,N_2754);
or U10144 (N_10144,N_54,N_7361);
and U10145 (N_10145,N_7438,N_3507);
nor U10146 (N_10146,N_8059,N_318);
and U10147 (N_10147,N_4669,N_6973);
and U10148 (N_10148,N_9210,N_3954);
or U10149 (N_10149,N_5328,N_9609);
and U10150 (N_10150,N_4702,N_5500);
nor U10151 (N_10151,N_8845,N_8340);
and U10152 (N_10152,N_5791,N_4890);
and U10153 (N_10153,N_9734,N_6801);
nor U10154 (N_10154,N_4461,N_2950);
xnor U10155 (N_10155,N_9786,N_9779);
or U10156 (N_10156,N_6528,N_9096);
xnor U10157 (N_10157,N_1139,N_785);
or U10158 (N_10158,N_5468,N_7887);
nor U10159 (N_10159,N_4751,N_2198);
and U10160 (N_10160,N_406,N_234);
and U10161 (N_10161,N_3999,N_2949);
xnor U10162 (N_10162,N_6389,N_4246);
nand U10163 (N_10163,N_3679,N_9917);
nor U10164 (N_10164,N_6685,N_2164);
nor U10165 (N_10165,N_2186,N_2318);
xnor U10166 (N_10166,N_2276,N_6131);
xnor U10167 (N_10167,N_1802,N_2498);
nand U10168 (N_10168,N_8872,N_4987);
nor U10169 (N_10169,N_5833,N_7610);
xnor U10170 (N_10170,N_6866,N_8996);
nor U10171 (N_10171,N_3243,N_1833);
xnor U10172 (N_10172,N_4667,N_2929);
xnor U10173 (N_10173,N_4392,N_3848);
nand U10174 (N_10174,N_5680,N_2645);
nor U10175 (N_10175,N_7573,N_1269);
and U10176 (N_10176,N_2978,N_722);
nor U10177 (N_10177,N_4916,N_1911);
and U10178 (N_10178,N_1803,N_6582);
nand U10179 (N_10179,N_8090,N_683);
and U10180 (N_10180,N_4303,N_7885);
xor U10181 (N_10181,N_2953,N_9281);
nand U10182 (N_10182,N_5266,N_4370);
or U10183 (N_10183,N_5988,N_483);
and U10184 (N_10184,N_3715,N_7538);
nor U10185 (N_10185,N_7678,N_177);
xor U10186 (N_10186,N_1055,N_9748);
or U10187 (N_10187,N_150,N_3048);
xnor U10188 (N_10188,N_3857,N_4131);
or U10189 (N_10189,N_5299,N_9613);
nor U10190 (N_10190,N_5033,N_4270);
xnor U10191 (N_10191,N_7254,N_3426);
xor U10192 (N_10192,N_6509,N_1199);
xor U10193 (N_10193,N_5369,N_2346);
nand U10194 (N_10194,N_8773,N_678);
or U10195 (N_10195,N_3093,N_3753);
or U10196 (N_10196,N_1037,N_9158);
nor U10197 (N_10197,N_607,N_3161);
and U10198 (N_10198,N_4925,N_5970);
nor U10199 (N_10199,N_3494,N_3941);
xor U10200 (N_10200,N_4784,N_8010);
xnor U10201 (N_10201,N_9312,N_6962);
xnor U10202 (N_10202,N_4485,N_4205);
nor U10203 (N_10203,N_3648,N_328);
or U10204 (N_10204,N_1963,N_9105);
and U10205 (N_10205,N_3257,N_6007);
nand U10206 (N_10206,N_6245,N_1529);
xor U10207 (N_10207,N_5212,N_9412);
or U10208 (N_10208,N_6001,N_8523);
and U10209 (N_10209,N_4569,N_4422);
and U10210 (N_10210,N_4943,N_789);
xor U10211 (N_10211,N_1673,N_5812);
and U10212 (N_10212,N_3484,N_1666);
xor U10213 (N_10213,N_8372,N_1723);
xor U10214 (N_10214,N_5207,N_1677);
xor U10215 (N_10215,N_7596,N_362);
nor U10216 (N_10216,N_6226,N_535);
xor U10217 (N_10217,N_7918,N_8748);
and U10218 (N_10218,N_9919,N_4518);
nor U10219 (N_10219,N_3221,N_4039);
or U10220 (N_10220,N_9839,N_190);
nor U10221 (N_10221,N_6676,N_1101);
and U10222 (N_10222,N_3447,N_6617);
xor U10223 (N_10223,N_1302,N_9401);
or U10224 (N_10224,N_145,N_4264);
or U10225 (N_10225,N_4542,N_8675);
nand U10226 (N_10226,N_207,N_4051);
xor U10227 (N_10227,N_2704,N_7029);
xor U10228 (N_10228,N_7934,N_3641);
nand U10229 (N_10229,N_9172,N_4382);
and U10230 (N_10230,N_9676,N_5973);
nor U10231 (N_10231,N_1207,N_3374);
xnor U10232 (N_10232,N_2106,N_3081);
and U10233 (N_10233,N_9151,N_810);
nand U10234 (N_10234,N_6860,N_6207);
and U10235 (N_10235,N_425,N_6285);
or U10236 (N_10236,N_6641,N_241);
nand U10237 (N_10237,N_169,N_3004);
and U10238 (N_10238,N_3297,N_6977);
nor U10239 (N_10239,N_5221,N_5267);
nor U10240 (N_10240,N_4214,N_3681);
nor U10241 (N_10241,N_78,N_1902);
nor U10242 (N_10242,N_1838,N_6067);
xnor U10243 (N_10243,N_9720,N_1484);
and U10244 (N_10244,N_5975,N_9856);
nor U10245 (N_10245,N_4918,N_7996);
or U10246 (N_10246,N_7525,N_8271);
nand U10247 (N_10247,N_6249,N_4219);
or U10248 (N_10248,N_2530,N_8089);
nand U10249 (N_10249,N_1362,N_8398);
nand U10250 (N_10250,N_6668,N_340);
xnor U10251 (N_10251,N_112,N_9217);
nand U10252 (N_10252,N_3881,N_5700);
and U10253 (N_10253,N_6497,N_4380);
and U10254 (N_10254,N_9257,N_6492);
nor U10255 (N_10255,N_9061,N_8541);
xor U10256 (N_10256,N_4796,N_948);
or U10257 (N_10257,N_4083,N_8766);
xor U10258 (N_10258,N_8274,N_2619);
nor U10259 (N_10259,N_567,N_4511);
xor U10260 (N_10260,N_5097,N_796);
and U10261 (N_10261,N_6990,N_8436);
and U10262 (N_10262,N_8317,N_2552);
xor U10263 (N_10263,N_2661,N_1440);
and U10264 (N_10264,N_7789,N_3123);
and U10265 (N_10265,N_9036,N_9527);
nand U10266 (N_10266,N_7666,N_206);
and U10267 (N_10267,N_4428,N_4566);
nand U10268 (N_10268,N_6208,N_2869);
nor U10269 (N_10269,N_7221,N_9468);
nor U10270 (N_10270,N_1474,N_3810);
or U10271 (N_10271,N_4688,N_7511);
nand U10272 (N_10272,N_8535,N_8438);
nor U10273 (N_10273,N_9436,N_8516);
nand U10274 (N_10274,N_5867,N_230);
xnor U10275 (N_10275,N_2177,N_7249);
nand U10276 (N_10276,N_2709,N_7402);
nand U10277 (N_10277,N_7585,N_289);
or U10278 (N_10278,N_8698,N_8205);
nor U10279 (N_10279,N_5692,N_3525);
and U10280 (N_10280,N_4826,N_2768);
nand U10281 (N_10281,N_9123,N_9411);
and U10282 (N_10282,N_9985,N_3380);
nor U10283 (N_10283,N_7856,N_5166);
and U10284 (N_10284,N_9840,N_3249);
nand U10285 (N_10285,N_5333,N_6306);
or U10286 (N_10286,N_3493,N_2226);
nor U10287 (N_10287,N_4801,N_2624);
xnor U10288 (N_10288,N_8652,N_4758);
nor U10289 (N_10289,N_7124,N_2866);
nor U10290 (N_10290,N_7913,N_5219);
and U10291 (N_10291,N_8786,N_8733);
xor U10292 (N_10292,N_7446,N_708);
nor U10293 (N_10293,N_9572,N_6252);
or U10294 (N_10294,N_9244,N_8664);
or U10295 (N_10295,N_7116,N_5928);
or U10296 (N_10296,N_2560,N_6871);
xor U10297 (N_10297,N_1074,N_3814);
xor U10298 (N_10298,N_2550,N_5176);
nand U10299 (N_10299,N_6983,N_44);
xor U10300 (N_10300,N_7459,N_5840);
nand U10301 (N_10301,N_8832,N_3794);
xor U10302 (N_10302,N_5879,N_1189);
or U10303 (N_10303,N_7628,N_226);
or U10304 (N_10304,N_5954,N_7423);
and U10305 (N_10305,N_7851,N_5966);
xnor U10306 (N_10306,N_8716,N_4917);
xnor U10307 (N_10307,N_3864,N_6276);
nor U10308 (N_10308,N_3611,N_8686);
xor U10309 (N_10309,N_3134,N_1355);
or U10310 (N_10310,N_5868,N_2128);
nand U10311 (N_10311,N_4496,N_1825);
or U10312 (N_10312,N_7308,N_6930);
xor U10313 (N_10313,N_2546,N_8580);
or U10314 (N_10314,N_6803,N_4494);
and U10315 (N_10315,N_6737,N_5388);
nand U10316 (N_10316,N_572,N_544);
or U10317 (N_10317,N_9743,N_6642);
or U10318 (N_10318,N_4052,N_4808);
nand U10319 (N_10319,N_543,N_6032);
or U10320 (N_10320,N_6981,N_5479);
nand U10321 (N_10321,N_2853,N_296);
nor U10322 (N_10322,N_9327,N_3311);
nor U10323 (N_10323,N_3241,N_6290);
or U10324 (N_10324,N_2016,N_329);
nand U10325 (N_10325,N_8375,N_9561);
or U10326 (N_10326,N_489,N_1031);
nor U10327 (N_10327,N_6720,N_3181);
and U10328 (N_10328,N_9212,N_6781);
or U10329 (N_10329,N_9554,N_265);
xor U10330 (N_10330,N_278,N_2134);
xnor U10331 (N_10331,N_2377,N_2567);
or U10332 (N_10332,N_781,N_8281);
nor U10333 (N_10333,N_2400,N_8178);
and U10334 (N_10334,N_1514,N_5490);
nor U10335 (N_10335,N_451,N_4994);
and U10336 (N_10336,N_3979,N_8979);
nor U10337 (N_10337,N_5142,N_4746);
nor U10338 (N_10338,N_989,N_1575);
and U10339 (N_10339,N_9021,N_5241);
or U10340 (N_10340,N_2248,N_3084);
xor U10341 (N_10341,N_8154,N_9850);
nand U10342 (N_10342,N_3385,N_5127);
xor U10343 (N_10343,N_6926,N_5887);
or U10344 (N_10344,N_4109,N_9322);
and U10345 (N_10345,N_5288,N_6732);
and U10346 (N_10346,N_6144,N_5018);
nand U10347 (N_10347,N_2957,N_3307);
xor U10348 (N_10348,N_7051,N_1979);
xnor U10349 (N_10349,N_7166,N_6760);
nand U10350 (N_10350,N_8140,N_6381);
xor U10351 (N_10351,N_6865,N_3652);
or U10352 (N_10352,N_3631,N_2118);
nor U10353 (N_10353,N_3919,N_2583);
and U10354 (N_10354,N_6661,N_3174);
and U10355 (N_10355,N_7352,N_370);
xnor U10356 (N_10356,N_630,N_1046);
nor U10357 (N_10357,N_6934,N_8155);
and U10358 (N_10358,N_8417,N_3738);
nor U10359 (N_10359,N_5593,N_9843);
xor U10360 (N_10360,N_1994,N_8548);
or U10361 (N_10361,N_4964,N_465);
nand U10362 (N_10362,N_1347,N_8552);
xor U10363 (N_10363,N_7043,N_6782);
and U10364 (N_10364,N_5681,N_1834);
or U10365 (N_10365,N_8459,N_1991);
or U10366 (N_10366,N_436,N_4913);
or U10367 (N_10367,N_8460,N_3500);
or U10368 (N_10368,N_5819,N_4841);
nor U10369 (N_10369,N_6715,N_9670);
nand U10370 (N_10370,N_1793,N_1959);
nor U10371 (N_10371,N_7129,N_8193);
nand U10372 (N_10372,N_380,N_7690);
or U10373 (N_10373,N_2699,N_9133);
xor U10374 (N_10374,N_5403,N_5828);
and U10375 (N_10375,N_5499,N_9805);
xnor U10376 (N_10376,N_5358,N_5755);
nand U10377 (N_10377,N_235,N_8518);
nor U10378 (N_10378,N_2851,N_186);
nand U10379 (N_10379,N_9699,N_8995);
and U10380 (N_10380,N_9971,N_3399);
nor U10381 (N_10381,N_6132,N_7318);
nor U10382 (N_10382,N_1508,N_2335);
nor U10383 (N_10383,N_5260,N_1191);
nor U10384 (N_10384,N_8859,N_1218);
or U10385 (N_10385,N_666,N_7884);
xor U10386 (N_10386,N_5516,N_6646);
nor U10387 (N_10387,N_2540,N_3609);
or U10388 (N_10388,N_6648,N_4497);
nor U10389 (N_10389,N_959,N_8342);
nor U10390 (N_10390,N_2789,N_4174);
xor U10391 (N_10391,N_5213,N_2967);
nand U10392 (N_10392,N_5880,N_8096);
and U10393 (N_10393,N_127,N_3613);
nor U10394 (N_10394,N_2195,N_5244);
nor U10395 (N_10395,N_5108,N_2192);
xnor U10396 (N_10396,N_336,N_2974);
nand U10397 (N_10397,N_1187,N_5264);
nand U10398 (N_10398,N_1593,N_354);
nand U10399 (N_10399,N_8379,N_7832);
nor U10400 (N_10400,N_2855,N_4168);
or U10401 (N_10401,N_7167,N_7162);
nand U10402 (N_10402,N_9137,N_4465);
xor U10403 (N_10403,N_4468,N_3143);
nor U10404 (N_10404,N_2332,N_277);
and U10405 (N_10405,N_346,N_4376);
or U10406 (N_10406,N_3182,N_5302);
nor U10407 (N_10407,N_6946,N_8282);
or U10408 (N_10408,N_8631,N_7244);
nor U10409 (N_10409,N_6883,N_9107);
nand U10410 (N_10410,N_7529,N_6547);
xnor U10411 (N_10411,N_6688,N_8449);
nor U10412 (N_10412,N_1801,N_3467);
nor U10413 (N_10413,N_453,N_3963);
and U10414 (N_10414,N_8279,N_4170);
xor U10415 (N_10415,N_4523,N_1001);
nand U10416 (N_10416,N_4237,N_5743);
nor U10417 (N_10417,N_9486,N_2895);
xnor U10418 (N_10418,N_337,N_4824);
or U10419 (N_10419,N_5888,N_7138);
nor U10420 (N_10420,N_7998,N_4744);
or U10421 (N_10421,N_2382,N_2296);
and U10422 (N_10422,N_621,N_4527);
xor U10423 (N_10423,N_776,N_8132);
or U10424 (N_10424,N_1357,N_9874);
xor U10425 (N_10425,N_1743,N_1602);
nor U10426 (N_10426,N_7708,N_2328);
nand U10427 (N_10427,N_9371,N_9747);
xor U10428 (N_10428,N_1974,N_2254);
and U10429 (N_10429,N_2057,N_8458);
xor U10430 (N_10430,N_5385,N_5020);
nor U10431 (N_10431,N_4442,N_2607);
or U10432 (N_10432,N_4459,N_3933);
or U10433 (N_10433,N_5744,N_9880);
and U10434 (N_10434,N_2646,N_2660);
nand U10435 (N_10435,N_2937,N_3578);
nand U10436 (N_10436,N_9349,N_6722);
nor U10437 (N_10437,N_6147,N_474);
and U10438 (N_10438,N_7094,N_954);
xor U10439 (N_10439,N_58,N_93);
nand U10440 (N_10440,N_5808,N_1186);
and U10441 (N_10441,N_6745,N_6206);
nor U10442 (N_10442,N_5734,N_4398);
and U10443 (N_10443,N_7236,N_2571);
xor U10444 (N_10444,N_3003,N_4226);
xnor U10445 (N_10445,N_6302,N_9524);
or U10446 (N_10446,N_5177,N_6875);
and U10447 (N_10447,N_7487,N_2877);
xor U10448 (N_10448,N_176,N_4749);
or U10449 (N_10449,N_4594,N_1161);
and U10450 (N_10450,N_3768,N_9605);
and U10451 (N_10451,N_1757,N_675);
nand U10452 (N_10452,N_4780,N_825);
or U10453 (N_10453,N_3981,N_5343);
and U10454 (N_10454,N_911,N_23);
xor U10455 (N_10455,N_6665,N_6767);
nor U10456 (N_10456,N_3410,N_1622);
nand U10457 (N_10457,N_3353,N_4768);
and U10458 (N_10458,N_6605,N_7089);
and U10459 (N_10459,N_131,N_4156);
or U10460 (N_10460,N_642,N_1674);
xnor U10461 (N_10461,N_6281,N_4870);
nor U10462 (N_10462,N_6061,N_286);
nand U10463 (N_10463,N_540,N_1526);
or U10464 (N_10464,N_8118,N_673);
and U10465 (N_10465,N_9289,N_408);
nor U10466 (N_10466,N_9636,N_9272);
nor U10467 (N_10467,N_2474,N_5724);
nand U10468 (N_10468,N_3937,N_2473);
nand U10469 (N_10469,N_3854,N_7570);
xnor U10470 (N_10470,N_2927,N_3189);
or U10471 (N_10471,N_5326,N_9476);
nor U10472 (N_10472,N_7768,N_7135);
nor U10473 (N_10473,N_5414,N_6154);
nor U10474 (N_10474,N_3154,N_3031);
or U10475 (N_10475,N_3600,N_3341);
or U10476 (N_10476,N_254,N_3822);
xor U10477 (N_10477,N_7845,N_9497);
or U10478 (N_10478,N_6846,N_5192);
nand U10479 (N_10479,N_9707,N_9931);
xor U10480 (N_10480,N_950,N_7232);
xnor U10481 (N_10481,N_8724,N_835);
nor U10482 (N_10482,N_2931,N_8620);
nor U10483 (N_10483,N_6921,N_4588);
nand U10484 (N_10484,N_7010,N_9356);
and U10485 (N_10485,N_5433,N_6701);
xnor U10486 (N_10486,N_2203,N_594);
or U10487 (N_10487,N_2986,N_1670);
xor U10488 (N_10488,N_2649,N_7591);
nand U10489 (N_10489,N_8320,N_6307);
nor U10490 (N_10490,N_1713,N_8191);
nor U10491 (N_10491,N_8452,N_3330);
xnor U10492 (N_10492,N_1238,N_3269);
and U10493 (N_10493,N_1935,N_7108);
nand U10494 (N_10494,N_6568,N_7616);
nor U10495 (N_10495,N_3363,N_3667);
or U10496 (N_10496,N_4630,N_2603);
or U10497 (N_10497,N_935,N_3888);
xnor U10498 (N_10498,N_6523,N_6244);
nand U10499 (N_10499,N_1580,N_5498);
xnor U10500 (N_10500,N_3795,N_3351);
xor U10501 (N_10501,N_1100,N_5762);
nor U10502 (N_10502,N_6079,N_3956);
xor U10503 (N_10503,N_9796,N_6438);
nand U10504 (N_10504,N_7827,N_5494);
or U10505 (N_10505,N_741,N_711);
or U10506 (N_10506,N_9704,N_2369);
or U10507 (N_10507,N_2130,N_7521);
xor U10508 (N_10508,N_8762,N_1174);
nor U10509 (N_10509,N_1617,N_2344);
nor U10510 (N_10510,N_5792,N_749);
nor U10511 (N_10511,N_3193,N_9565);
and U10512 (N_10512,N_3655,N_3204);
and U10513 (N_10513,N_7719,N_3044);
xnor U10514 (N_10514,N_2323,N_4998);
xnor U10515 (N_10515,N_2640,N_8804);
or U10516 (N_10516,N_9117,N_8941);
nand U10517 (N_10517,N_48,N_3673);
nand U10518 (N_10518,N_4227,N_1927);
nand U10519 (N_10519,N_393,N_2872);
xor U10520 (N_10520,N_3047,N_8797);
and U10521 (N_10521,N_3553,N_6121);
nor U10522 (N_10522,N_6490,N_5852);
or U10523 (N_10523,N_7384,N_6624);
nand U10524 (N_10524,N_4825,N_3272);
nor U10525 (N_10525,N_5076,N_5847);
or U10526 (N_10526,N_1599,N_9724);
or U10527 (N_10527,N_529,N_1047);
xor U10528 (N_10528,N_5396,N_9160);
or U10529 (N_10529,N_2874,N_1573);
nand U10530 (N_10530,N_561,N_2700);
or U10531 (N_10531,N_8730,N_5061);
or U10532 (N_10532,N_8937,N_5967);
and U10533 (N_10533,N_1787,N_5658);
nor U10534 (N_10534,N_1931,N_6964);
nand U10535 (N_10535,N_9769,N_7860);
xor U10536 (N_10536,N_6670,N_6969);
xor U10537 (N_10537,N_4111,N_1846);
and U10538 (N_10538,N_4915,N_3705);
nand U10539 (N_10539,N_9781,N_7972);
nand U10540 (N_10540,N_5491,N_3465);
nor U10541 (N_10541,N_9228,N_9742);
xnor U10542 (N_10542,N_9694,N_1614);
and U10543 (N_10543,N_914,N_2379);
and U10544 (N_10544,N_5769,N_6343);
xor U10545 (N_10545,N_3037,N_5897);
or U10546 (N_10546,N_1960,N_351);
xor U10547 (N_10547,N_1904,N_8779);
and U10548 (N_10548,N_6751,N_9900);
nand U10549 (N_10549,N_9141,N_5105);
xnor U10550 (N_10550,N_8127,N_6508);
nor U10551 (N_10551,N_7945,N_8050);
xnor U10552 (N_10552,N_9254,N_8917);
nor U10553 (N_10553,N_7631,N_5094);
nand U10554 (N_10554,N_6150,N_3362);
xor U10555 (N_10555,N_4647,N_7615);
or U10556 (N_10556,N_1409,N_3789);
and U10557 (N_10557,N_9788,N_8629);
nand U10558 (N_10558,N_8583,N_4088);
nor U10559 (N_10559,N_1285,N_2191);
or U10560 (N_10560,N_4404,N_1305);
xnor U10561 (N_10561,N_6499,N_3938);
nor U10562 (N_10562,N_5691,N_420);
or U10563 (N_10563,N_2,N_5572);
xnor U10564 (N_10564,N_4555,N_8918);
nor U10565 (N_10565,N_214,N_2314);
or U10566 (N_10566,N_2534,N_9888);
xnor U10567 (N_10567,N_8484,N_8777);
xor U10568 (N_10568,N_4500,N_101);
nor U10569 (N_10569,N_1969,N_6882);
xnor U10570 (N_10570,N_2348,N_3650);
xnor U10571 (N_10571,N_615,N_679);
or U10572 (N_10572,N_3381,N_836);
nand U10573 (N_10573,N_7846,N_4912);
xnor U10574 (N_10574,N_9029,N_6815);
and U10575 (N_10575,N_2482,N_9366);
and U10576 (N_10576,N_6457,N_5263);
xnor U10577 (N_10577,N_9989,N_5410);
or U10578 (N_10578,N_1491,N_4155);
xor U10579 (N_10579,N_2566,N_7240);
and U10580 (N_10580,N_5806,N_3852);
or U10581 (N_10581,N_2313,N_1848);
nor U10582 (N_10582,N_8862,N_2712);
and U10583 (N_10583,N_2888,N_6584);
xnor U10584 (N_10584,N_166,N_7854);
xor U10585 (N_10585,N_4119,N_2936);
nand U10586 (N_10586,N_7344,N_6310);
and U10587 (N_10587,N_9952,N_1344);
and U10588 (N_10588,N_4001,N_4278);
and U10589 (N_10589,N_2520,N_2865);
or U10590 (N_10590,N_7169,N_1500);
or U10591 (N_10591,N_1946,N_3724);
and U10592 (N_10592,N_8453,N_490);
and U10593 (N_10593,N_3620,N_2601);
nor U10594 (N_10594,N_6209,N_470);
nor U10595 (N_10595,N_5505,N_9618);
or U10596 (N_10596,N_3369,N_6452);
xnor U10597 (N_10597,N_6466,N_9296);
nor U10598 (N_10598,N_1481,N_1780);
or U10599 (N_10599,N_9405,N_2113);
xor U10600 (N_10600,N_204,N_3952);
xor U10601 (N_10601,N_6913,N_5741);
nand U10602 (N_10602,N_8468,N_5891);
nor U10603 (N_10603,N_2340,N_8706);
nor U10604 (N_10604,N_477,N_9808);
and U10605 (N_10605,N_2896,N_4973);
nor U10606 (N_10606,N_7099,N_5017);
nand U10607 (N_10607,N_9084,N_2742);
nand U10608 (N_10608,N_7192,N_9922);
xnor U10609 (N_10609,N_5087,N_1581);
nand U10610 (N_10610,N_4456,N_3865);
and U10611 (N_10611,N_5074,N_8812);
nor U10612 (N_10612,N_5090,N_2108);
nand U10613 (N_10613,N_685,N_7778);
and U10614 (N_10614,N_5773,N_2259);
and U10615 (N_10615,N_5103,N_135);
nand U10616 (N_10616,N_634,N_5218);
nand U10617 (N_10617,N_7002,N_9397);
xnor U10618 (N_10618,N_9443,N_2622);
xnor U10619 (N_10619,N_9262,N_302);
or U10620 (N_10620,N_5200,N_4993);
or U10621 (N_10621,N_7790,N_2126);
and U10622 (N_10622,N_9620,N_2136);
nand U10623 (N_10623,N_1806,N_1243);
and U10624 (N_10624,N_2201,N_7040);
and U10625 (N_10625,N_3475,N_7937);
or U10626 (N_10626,N_1831,N_7801);
nand U10627 (N_10627,N_9248,N_8825);
and U10628 (N_10628,N_4927,N_9596);
nor U10629 (N_10629,N_8885,N_5603);
nor U10630 (N_10630,N_2819,N_6691);
nor U10631 (N_10631,N_1064,N_6929);
or U10632 (N_10632,N_9,N_7144);
and U10633 (N_10633,N_2815,N_4650);
and U10634 (N_10634,N_7033,N_8568);
nand U10635 (N_10635,N_8511,N_2677);
or U10636 (N_10636,N_4147,N_2427);
nor U10637 (N_10637,N_6185,N_4659);
xnor U10638 (N_10638,N_7414,N_7389);
xor U10639 (N_10639,N_9030,N_1210);
nor U10640 (N_10640,N_70,N_1875);
xnor U10641 (N_10641,N_1340,N_5437);
nor U10642 (N_10642,N_6374,N_8395);
xnor U10643 (N_10643,N_9718,N_9364);
or U10644 (N_10644,N_5079,N_8319);
or U10645 (N_10645,N_7909,N_6394);
or U10646 (N_10646,N_718,N_2989);
and U10647 (N_10647,N_4926,N_6712);
xnor U10648 (N_10648,N_8800,N_2975);
and U10649 (N_10649,N_1709,N_6056);
xnor U10650 (N_10650,N_9268,N_527);
and U10651 (N_10651,N_8351,N_5298);
nand U10652 (N_10652,N_4770,N_2598);
and U10653 (N_10653,N_188,N_1241);
xor U10654 (N_10654,N_6682,N_5622);
nor U10655 (N_10655,N_5165,N_4935);
nor U10656 (N_10656,N_4384,N_8670);
nand U10657 (N_10657,N_8567,N_252);
or U10658 (N_10658,N_8080,N_9166);
nand U10659 (N_10659,N_2172,N_5637);
and U10660 (N_10660,N_1182,N_3375);
nor U10661 (N_10661,N_5304,N_4363);
or U10662 (N_10662,N_9128,N_9726);
nor U10663 (N_10663,N_620,N_9495);
and U10664 (N_10664,N_2007,N_1304);
and U10665 (N_10665,N_542,N_9652);
nand U10666 (N_10666,N_994,N_4878);
nand U10667 (N_10667,N_1542,N_5911);
nor U10668 (N_10668,N_3400,N_8251);
and U10669 (N_10669,N_4017,N_4192);
or U10670 (N_10670,N_4711,N_5124);
nand U10671 (N_10671,N_9547,N_478);
and U10672 (N_10672,N_4282,N_5549);
or U10673 (N_10673,N_5767,N_9733);
and U10674 (N_10674,N_2060,N_3451);
nand U10675 (N_10675,N_9570,N_390);
xor U10676 (N_10676,N_4769,N_6583);
nand U10677 (N_10677,N_4662,N_988);
and U10678 (N_10678,N_6459,N_9285);
xnor U10679 (N_10679,N_5989,N_6019);
and U10680 (N_10680,N_2903,N_8572);
or U10681 (N_10681,N_4449,N_1134);
xor U10682 (N_10682,N_1980,N_7482);
nand U10683 (N_10683,N_3247,N_7820);
nor U10684 (N_10684,N_9282,N_6723);
nand U10685 (N_10685,N_1025,N_2717);
nor U10686 (N_10686,N_8912,N_3021);
nand U10687 (N_10687,N_6095,N_7655);
xnor U10688 (N_10688,N_4715,N_3121);
nand U10689 (N_10689,N_6672,N_1054);
and U10690 (N_10690,N_7267,N_665);
xnor U10691 (N_10691,N_6211,N_5764);
or U10692 (N_10692,N_2958,N_3207);
and U10693 (N_10693,N_8359,N_72);
xnor U10694 (N_10694,N_5903,N_363);
nand U10695 (N_10695,N_3867,N_3713);
nand U10696 (N_10696,N_3455,N_7821);
nor U10697 (N_10697,N_3365,N_3271);
nand U10698 (N_10698,N_907,N_7983);
nor U10699 (N_10699,N_4366,N_6881);
xnor U10700 (N_10700,N_8704,N_8256);
nand U10701 (N_10701,N_6416,N_6652);
and U10702 (N_10702,N_9705,N_4995);
nand U10703 (N_10703,N_1213,N_9516);
and U10704 (N_10704,N_3967,N_6117);
nand U10705 (N_10705,N_3692,N_9310);
xnor U10706 (N_10706,N_1327,N_9109);
and U10707 (N_10707,N_6300,N_3755);
or U10708 (N_10708,N_3722,N_1127);
nor U10709 (N_10709,N_1148,N_5781);
nor U10710 (N_10710,N_1910,N_1451);
or U10711 (N_10711,N_2720,N_8495);
and U10712 (N_10712,N_1885,N_4886);
or U10713 (N_10713,N_4956,N_6683);
nand U10714 (N_10714,N_8954,N_3498);
and U10715 (N_10715,N_6758,N_2612);
and U10716 (N_10716,N_5287,N_1988);
nand U10717 (N_10717,N_5668,N_423);
or U10718 (N_10718,N_5768,N_2787);
nor U10719 (N_10719,N_872,N_4439);
nor U10720 (N_10720,N_953,N_5240);
nand U10721 (N_10721,N_1841,N_3697);
nand U10722 (N_10722,N_2450,N_1271);
nor U10723 (N_10723,N_5754,N_855);
nand U10724 (N_10724,N_8402,N_7147);
nand U10725 (N_10725,N_5616,N_9883);
nand U10726 (N_10726,N_2669,N_2049);
nor U10727 (N_10727,N_5361,N_3714);
or U10728 (N_10728,N_8091,N_9390);
xnor U10729 (N_10729,N_2630,N_3766);
and U10730 (N_10730,N_6902,N_5909);
xnor U10731 (N_10731,N_4923,N_4427);
nand U10732 (N_10732,N_8942,N_8266);
or U10733 (N_10733,N_9098,N_4986);
nor U10734 (N_10734,N_7209,N_4444);
and U10735 (N_10735,N_5733,N_1360);
and U10736 (N_10736,N_5998,N_6927);
xnor U10737 (N_10737,N_8895,N_9155);
nand U10738 (N_10738,N_3377,N_2467);
and U10739 (N_10739,N_1369,N_4846);
and U10740 (N_10740,N_4725,N_8826);
and U10741 (N_10741,N_1403,N_167);
nand U10742 (N_10742,N_9104,N_8625);
xor U10743 (N_10743,N_9719,N_2090);
and U10744 (N_10744,N_1090,N_325);
and U10745 (N_10745,N_2300,N_6433);
and U10746 (N_10746,N_9479,N_7350);
xnor U10747 (N_10747,N_2221,N_6917);
or U10748 (N_10748,N_3303,N_616);
xor U10749 (N_10749,N_345,N_5546);
or U10750 (N_10750,N_2753,N_3270);
nand U10751 (N_10751,N_8821,N_2470);
or U10752 (N_10752,N_5841,N_5580);
xor U10753 (N_10753,N_9095,N_768);
and U10754 (N_10754,N_6718,N_4967);
or U10755 (N_10755,N_6573,N_4896);
and U10756 (N_10756,N_7340,N_617);
nand U10757 (N_10757,N_3448,N_4761);
and U10758 (N_10758,N_8606,N_4651);
and U10759 (N_10759,N_376,N_6619);
nor U10760 (N_10760,N_5645,N_7707);
or U10761 (N_10761,N_1185,N_8915);
nand U10762 (N_10762,N_8437,N_4615);
or U10763 (N_10763,N_4285,N_6022);
nand U10764 (N_10764,N_4716,N_7425);
and U10765 (N_10765,N_7514,N_2919);
nor U10766 (N_10766,N_9060,N_7145);
nand U10767 (N_10767,N_8300,N_619);
xnor U10768 (N_10768,N_5372,N_1555);
nand U10769 (N_10769,N_1527,N_5028);
xor U10770 (N_10770,N_7156,N_7504);
nor U10771 (N_10771,N_7133,N_793);
or U10772 (N_10772,N_8517,N_499);
or U10773 (N_10773,N_3298,N_9319);
or U10774 (N_10774,N_4513,N_5567);
xor U10775 (N_10775,N_7838,N_707);
and U10776 (N_10776,N_8428,N_1112);
or U10777 (N_10777,N_9571,N_5023);
nand U10778 (N_10778,N_3593,N_4554);
nor U10779 (N_10779,N_3260,N_3658);
nor U10780 (N_10780,N_6246,N_2018);
nand U10781 (N_10781,N_771,N_6644);
nand U10782 (N_10782,N_4534,N_5839);
or U10783 (N_10783,N_5439,N_3013);
and U10784 (N_10784,N_5159,N_2161);
or U10785 (N_10785,N_3560,N_9657);
xnor U10786 (N_10786,N_1021,N_2059);
or U10787 (N_10787,N_1634,N_3007);
and U10788 (N_10788,N_5188,N_217);
or U10789 (N_10789,N_8307,N_3902);
nor U10790 (N_10790,N_9121,N_6023);
xor U10791 (N_10791,N_1760,N_5625);
nor U10792 (N_10792,N_6242,N_4418);
and U10793 (N_10793,N_3458,N_3540);
or U10794 (N_10794,N_9326,N_1006);
nand U10795 (N_10795,N_7803,N_6105);
nand U10796 (N_10796,N_8487,N_1777);
nor U10797 (N_10797,N_8910,N_9949);
xnor U10798 (N_10798,N_5732,N_9247);
xnor U10799 (N_10799,N_7865,N_8827);
nand U10800 (N_10800,N_9871,N_7358);
nor U10801 (N_10801,N_274,N_5881);
nand U10802 (N_10802,N_4884,N_3760);
xnor U10803 (N_10803,N_1888,N_3501);
nor U10804 (N_10804,N_9906,N_2309);
xor U10805 (N_10805,N_2761,N_7258);
xor U10806 (N_10806,N_319,N_8224);
nand U10807 (N_10807,N_8253,N_1525);
nor U10808 (N_10808,N_9428,N_1145);
and U10809 (N_10809,N_9728,N_4085);
nor U10810 (N_10810,N_3858,N_8);
nand U10811 (N_10811,N_7921,N_6664);
and U10812 (N_10812,N_545,N_1232);
nor U10813 (N_10813,N_780,N_8688);
and U10814 (N_10814,N_2905,N_910);
or U10815 (N_10815,N_9939,N_9946);
xnor U10816 (N_10816,N_4665,N_7557);
nor U10817 (N_10817,N_5308,N_3088);
or U10818 (N_10818,N_3787,N_6831);
or U10819 (N_10819,N_9607,N_828);
nor U10820 (N_10820,N_4399,N_4160);
or U10821 (N_10821,N_8640,N_1289);
xnor U10822 (N_10822,N_7148,N_6167);
and U10823 (N_10823,N_7229,N_4256);
nand U10824 (N_10824,N_7576,N_5619);
nand U10825 (N_10825,N_7653,N_1477);
nand U10826 (N_10826,N_4144,N_3211);
and U10827 (N_10827,N_88,N_7782);
nor U10828 (N_10828,N_98,N_3258);
and U10829 (N_10829,N_6044,N_3799);
or U10830 (N_10830,N_2038,N_6198);
nor U10831 (N_10831,N_2750,N_1107);
or U10832 (N_10832,N_2412,N_9854);
nand U10833 (N_10833,N_680,N_9031);
xnor U10834 (N_10834,N_1004,N_7978);
and U10835 (N_10835,N_9928,N_219);
or U10836 (N_10836,N_8968,N_9074);
and U10837 (N_10837,N_2868,N_6693);
xor U10838 (N_10838,N_2349,N_5447);
nor U10839 (N_10839,N_106,N_1696);
nor U10840 (N_10840,N_8532,N_5986);
xnor U10841 (N_10841,N_1752,N_5044);
xnor U10842 (N_10842,N_1160,N_801);
or U10843 (N_10843,N_20,N_1153);
or U10844 (N_10844,N_8283,N_795);
xnor U10845 (N_10845,N_1430,N_7866);
xor U10846 (N_10846,N_8465,N_1828);
xnor U10847 (N_10847,N_1859,N_5683);
xnor U10848 (N_10848,N_256,N_6725);
xor U10849 (N_10849,N_8009,N_7763);
xor U10850 (N_10850,N_5829,N_9591);
or U10851 (N_10851,N_6686,N_5001);
and U10852 (N_10852,N_4820,N_7774);
xnor U10853 (N_10853,N_8149,N_2945);
or U10854 (N_10854,N_4421,N_6063);
nor U10855 (N_10855,N_9722,N_3020);
xor U10856 (N_10856,N_9382,N_4900);
nand U10857 (N_10857,N_6873,N_5663);
nand U10858 (N_10858,N_4686,N_1948);
and U10859 (N_10859,N_9493,N_9597);
and U10860 (N_10860,N_2690,N_1396);
and U10861 (N_10861,N_4386,N_3536);
nor U10862 (N_10862,N_7222,N_3051);
and U10863 (N_10863,N_5539,N_388);
nor U10864 (N_10864,N_8053,N_5307);
xor U10865 (N_10865,N_7474,N_1929);
nand U10866 (N_10866,N_8515,N_9891);
xor U10867 (N_10867,N_1745,N_87);
nor U10868 (N_10868,N_4807,N_8847);
nor U10869 (N_10869,N_3527,N_7042);
and U10870 (N_10870,N_713,N_9291);
or U10871 (N_10871,N_4401,N_4224);
nand U10872 (N_10872,N_2685,N_3539);
or U10873 (N_10873,N_7250,N_1084);
or U10874 (N_10874,N_9972,N_5647);
or U10875 (N_10875,N_6538,N_1088);
xnor U10876 (N_10876,N_3693,N_8993);
nor U10877 (N_10877,N_307,N_5502);
and U10878 (N_10878,N_3130,N_2618);
or U10879 (N_10879,N_2301,N_3551);
nor U10880 (N_10880,N_9634,N_8387);
nand U10881 (N_10881,N_9543,N_9545);
nand U10882 (N_10882,N_9231,N_897);
nor U10883 (N_10883,N_5548,N_9047);
nor U10884 (N_10884,N_3215,N_9526);
nand U10885 (N_10885,N_6429,N_8315);
or U10886 (N_10886,N_259,N_2539);
nor U10887 (N_10887,N_8962,N_1626);
nand U10888 (N_10888,N_3706,N_962);
and U10889 (N_10889,N_7863,N_7022);
xnor U10890 (N_10890,N_5270,N_3384);
nand U10891 (N_10891,N_9127,N_282);
nand U10892 (N_10892,N_2404,N_14);
and U10893 (N_10893,N_3915,N_2326);
and U10894 (N_10894,N_7149,N_4396);
or U10895 (N_10895,N_7437,N_9709);
nor U10896 (N_10896,N_33,N_2247);
nor U10897 (N_10897,N_6432,N_8685);
and U10898 (N_10898,N_8725,N_3368);
or U10899 (N_10899,N_4862,N_7601);
or U10900 (N_10900,N_7449,N_4150);
xnor U10901 (N_10901,N_1683,N_4068);
xor U10902 (N_10902,N_8401,N_9780);
nor U10903 (N_10903,N_3203,N_6891);
nor U10904 (N_10904,N_6439,N_2653);
xor U10905 (N_10905,N_1983,N_2626);
or U10906 (N_10906,N_6543,N_8348);
or U10907 (N_10907,N_2782,N_723);
nor U10908 (N_10908,N_9685,N_4076);
nand U10909 (N_10909,N_9794,N_3376);
or U10910 (N_10910,N_4180,N_9427);
xnor U10911 (N_10911,N_8159,N_3450);
nand U10912 (N_10912,N_8064,N_7932);
or U10913 (N_10913,N_1657,N_8467);
or U10914 (N_10914,N_2381,N_9269);
or U10915 (N_10915,N_5204,N_5849);
nor U10916 (N_10916,N_3544,N_1331);
nand U10917 (N_10917,N_8589,N_8976);
nand U10918 (N_10918,N_4188,N_3216);
or U10919 (N_10919,N_5907,N_6906);
xnor U10920 (N_10920,N_6354,N_9062);
nand U10921 (N_10921,N_2867,N_571);
nand U10922 (N_10922,N_64,N_3280);
nor U10923 (N_10923,N_6818,N_7709);
and U10924 (N_10924,N_5536,N_5961);
nor U10925 (N_10925,N_794,N_6826);
or U10926 (N_10926,N_6761,N_976);
or U10927 (N_10927,N_2516,N_409);
nor U10928 (N_10928,N_7911,N_3036);
or U10929 (N_10929,N_3698,N_32);
nor U10930 (N_10930,N_7539,N_4212);
xnor U10931 (N_10931,N_1775,N_2990);
and U10932 (N_10932,N_1607,N_1458);
and U10933 (N_10933,N_3685,N_8930);
xor U10934 (N_10934,N_705,N_2448);
xor U10935 (N_10935,N_1517,N_5136);
nor U10936 (N_10936,N_9111,N_8994);
xor U10937 (N_10937,N_4549,N_2558);
nor U10938 (N_10938,N_3195,N_7736);
nor U10939 (N_10939,N_9357,N_4617);
or U10940 (N_10940,N_9625,N_6702);
or U10941 (N_10941,N_9557,N_590);
or U10942 (N_10942,N_8439,N_2122);
and U10943 (N_10943,N_5807,N_6177);
xor U10944 (N_10944,N_7510,N_2437);
nand U10945 (N_10945,N_4552,N_8959);
or U10946 (N_10946,N_5556,N_4272);
xnor U10947 (N_10947,N_1377,N_8345);
or U10948 (N_10948,N_1589,N_7575);
nand U10949 (N_10949,N_6423,N_6218);
nor U10950 (N_10950,N_6630,N_3774);
nand U10951 (N_10951,N_232,N_8176);
nand U10952 (N_10952,N_4244,N_4032);
nand U10953 (N_10953,N_2307,N_8177);
or U10954 (N_10954,N_3471,N_7629);
xnor U10955 (N_10955,N_721,N_4633);
or U10956 (N_10956,N_3654,N_3230);
and U10957 (N_10957,N_8124,N_5893);
nand U10958 (N_10958,N_7536,N_8896);
xnor U10959 (N_10959,N_4972,N_2279);
and U10960 (N_10960,N_3418,N_5060);
nor U10961 (N_10961,N_6554,N_8615);
or U10962 (N_10962,N_7445,N_2708);
and U10963 (N_10963,N_2841,N_1402);
nand U10964 (N_10964,N_5397,N_4983);
or U10965 (N_10965,N_229,N_7153);
nor U10966 (N_10966,N_7366,N_2109);
nand U10967 (N_10967,N_4949,N_6173);
nand U10968 (N_10968,N_3396,N_1823);
or U10969 (N_10969,N_3138,N_9352);
and U10970 (N_10970,N_5992,N_201);
or U10971 (N_10971,N_4576,N_3173);
nor U10972 (N_10972,N_1932,N_7816);
nand U10973 (N_10973,N_6954,N_4950);
or U10974 (N_10974,N_1299,N_3895);
and U10975 (N_10975,N_9394,N_5497);
nor U10976 (N_10976,N_2175,N_482);
and U10977 (N_10977,N_9674,N_8498);
xor U10978 (N_10978,N_159,N_6338);
xnor U10979 (N_10979,N_8799,N_2813);
nand U10980 (N_10980,N_4470,N_2494);
xnor U10981 (N_10981,N_5987,N_1579);
and U10982 (N_10982,N_3801,N_468);
or U10983 (N_10983,N_7619,N_114);
or U10984 (N_10984,N_387,N_5836);
or U10985 (N_10985,N_4530,N_3457);
and U10986 (N_10986,N_1098,N_2408);
xnor U10987 (N_10987,N_4351,N_7088);
nor U10988 (N_10988,N_4928,N_668);
xnor U10989 (N_10989,N_6621,N_5581);
xor U10990 (N_10990,N_8781,N_7675);
and U10991 (N_10991,N_2492,N_7791);
nor U10992 (N_10992,N_1094,N_5138);
and U10993 (N_10993,N_7464,N_9132);
nor U10994 (N_10994,N_4567,N_2157);
and U10995 (N_10995,N_8261,N_164);
and U10996 (N_10996,N_2133,N_7930);
and U10997 (N_10997,N_9552,N_3027);
xnor U10998 (N_10998,N_4225,N_8086);
xor U10999 (N_10999,N_8087,N_8947);
or U11000 (N_11000,N_5280,N_1535);
and U11001 (N_11001,N_5699,N_9230);
and U11002 (N_11002,N_279,N_8720);
xor U11003 (N_11003,N_3850,N_1068);
nor U11004 (N_11004,N_3460,N_1057);
or U11005 (N_11005,N_3624,N_8446);
nor U11006 (N_11006,N_50,N_6051);
nor U11007 (N_11007,N_2628,N_3832);
nor U11008 (N_11008,N_3893,N_4799);
and U11009 (N_11009,N_5208,N_877);
or U11010 (N_11010,N_2870,N_9465);
xnor U11011 (N_11011,N_9439,N_389);
or U11012 (N_11012,N_6643,N_7106);
xor U11013 (N_11013,N_6941,N_4850);
and U11014 (N_11014,N_5442,N_3300);
nor U11015 (N_11015,N_5237,N_5621);
and U11016 (N_11016,N_5363,N_8633);
nand U11017 (N_11017,N_4445,N_694);
or U11018 (N_11018,N_42,N_7253);
and U11019 (N_11019,N_444,N_1159);
xor U11020 (N_11020,N_4628,N_9226);
nor U11021 (N_11021,N_2889,N_4940);
or U11022 (N_11022,N_7590,N_8772);
xnor U11023 (N_11023,N_2849,N_1623);
and U11024 (N_11024,N_9182,N_9528);
and U11025 (N_11025,N_6585,N_532);
xnor U11026 (N_11026,N_4601,N_608);
nor U11027 (N_11027,N_9261,N_8380);
xor U11028 (N_11028,N_9211,N_8897);
xnor U11029 (N_11029,N_4991,N_912);
nand U11030 (N_11030,N_6916,N_8657);
xor U11031 (N_11031,N_7829,N_1610);
nand U11032 (N_11032,N_8394,N_9580);
nand U11033 (N_11033,N_8119,N_6511);
xor U11034 (N_11034,N_4295,N_8148);
xnor U11035 (N_11035,N_9877,N_7811);
nand U11036 (N_11036,N_5296,N_8705);
xnor U11037 (N_11037,N_1251,N_4169);
nand U11038 (N_11038,N_202,N_9249);
nand U11039 (N_11039,N_2679,N_1462);
nor U11040 (N_11040,N_7245,N_2535);
xor U11041 (N_11041,N_7045,N_5736);
and U11042 (N_11042,N_5525,N_677);
or U11043 (N_11043,N_7800,N_3993);
xnor U11044 (N_11044,N_3167,N_981);
nor U11045 (N_11045,N_6541,N_5651);
and U11046 (N_11046,N_9462,N_8655);
xor U11047 (N_11047,N_4336,N_1533);
xnor U11048 (N_11048,N_7489,N_9606);
or U11049 (N_11049,N_3045,N_9584);
nand U11050 (N_11050,N_2321,N_9616);
or U11051 (N_11051,N_7671,N_751);
and U11052 (N_11052,N_6153,N_9714);
or U11053 (N_11053,N_1483,N_852);
or U11054 (N_11054,N_2585,N_2555);
nor U11055 (N_11055,N_9455,N_7830);
nor U11056 (N_11056,N_4963,N_6280);
nor U11057 (N_11057,N_982,N_3838);
xnor U11058 (N_11058,N_2858,N_7466);
nand U11059 (N_11059,N_6379,N_3386);
nand U11060 (N_11060,N_5129,N_984);
nand U11061 (N_11061,N_2814,N_2190);
nand U11062 (N_11062,N_2532,N_5429);
or U11063 (N_11063,N_475,N_2702);
or U11064 (N_11064,N_7952,N_2718);
xor U11065 (N_11065,N_3074,N_1504);
or U11066 (N_11066,N_2319,N_9185);
and U11067 (N_11067,N_5077,N_7328);
nor U11068 (N_11068,N_7662,N_5605);
xor U11069 (N_11069,N_1883,N_6700);
and U11070 (N_11070,N_3944,N_5538);
and U11071 (N_11071,N_1445,N_9169);
and U11072 (N_11072,N_8354,N_7097);
nor U11073 (N_11073,N_4043,N_4797);
nor U11074 (N_11074,N_8753,N_538);
nand U11075 (N_11075,N_1867,N_5413);
nand U11076 (N_11076,N_6042,N_9317);
nor U11077 (N_11077,N_334,N_9451);
and U11078 (N_11078,N_517,N_8745);
xor U11079 (N_11079,N_9866,N_365);
and U11080 (N_11080,N_9813,N_5387);
nor U11081 (N_11081,N_3763,N_8873);
nand U11082 (N_11082,N_3939,N_6046);
nand U11083 (N_11083,N_3087,N_4269);
xor U11084 (N_11084,N_9575,N_6660);
xor U11085 (N_11085,N_9354,N_2678);
and U11086 (N_11086,N_2969,N_4318);
nand U11087 (N_11087,N_9429,N_2491);
xnor U11088 (N_11088,N_8020,N_1106);
xor U11089 (N_11089,N_2883,N_1116);
xnor U11090 (N_11090,N_7862,N_424);
nand U11091 (N_11091,N_344,N_130);
xor U11092 (N_11092,N_3372,N_9804);
nand U11093 (N_11093,N_9316,N_6830);
xor U11094 (N_11094,N_1943,N_8058);
nor U11095 (N_11095,N_8988,N_833);
nor U11096 (N_11096,N_9958,N_9256);
nand U11097 (N_11097,N_6963,N_4843);
nand U11098 (N_11098,N_8296,N_4775);
xnor U11099 (N_11099,N_8440,N_8884);
nor U11100 (N_11100,N_5981,N_6857);
nor U11101 (N_11101,N_3214,N_79);
nand U11102 (N_11102,N_7123,N_7796);
nand U11103 (N_11103,N_8758,N_9979);
xnor U11104 (N_11104,N_1290,N_4759);
xor U11105 (N_11105,N_6278,N_709);
and U11106 (N_11106,N_9090,N_3998);
or U11107 (N_11107,N_3325,N_6123);
nand U11108 (N_11108,N_1523,N_3091);
nor U11109 (N_11109,N_1546,N_3175);
and U11110 (N_11110,N_1459,N_3735);
nor U11111 (N_11111,N_7070,N_7286);
and U11112 (N_11112,N_5564,N_3395);
nand U11113 (N_11113,N_7744,N_123);
nor U11114 (N_11114,N_676,N_3238);
or U11115 (N_11115,N_7295,N_2271);
nand U11116 (N_11116,N_1249,N_7087);
or U11117 (N_11117,N_5904,N_1917);
nor U11118 (N_11118,N_6181,N_1655);
xnor U11119 (N_11119,N_4275,N_2105);
nand U11120 (N_11120,N_924,N_3155);
nor U11121 (N_11121,N_3945,N_6919);
or U11122 (N_11122,N_2892,N_5706);
nor U11123 (N_11123,N_7517,N_2176);
or U11124 (N_11124,N_5383,N_5566);
xor U11125 (N_11125,N_2676,N_5664);
or U11126 (N_11126,N_5760,N_9501);
xor U11127 (N_11127,N_9537,N_266);
and U11128 (N_11128,N_3302,N_5426);
or U11129 (N_11129,N_3636,N_7025);
and U11130 (N_11130,N_9025,N_63);
or U11131 (N_11131,N_1328,N_6481);
nor U11132 (N_11132,N_6697,N_9627);
xor U11133 (N_11133,N_6464,N_6163);
and U11134 (N_11134,N_2860,N_4472);
and U11135 (N_11135,N_8163,N_5440);
xor U11136 (N_11136,N_141,N_7773);
nand U11137 (N_11137,N_3185,N_8217);
xor U11138 (N_11138,N_879,N_2125);
and U11139 (N_11139,N_9766,N_786);
nor U11140 (N_11140,N_1625,N_6385);
nand U11141 (N_11141,N_2611,N_8056);
nand U11142 (N_11142,N_2395,N_3577);
and U11143 (N_11143,N_8330,N_7533);
xor U11144 (N_11144,N_2934,N_9086);
and U11145 (N_11145,N_4369,N_6320);
nand U11146 (N_11146,N_3414,N_7520);
or U11147 (N_11147,N_3556,N_1103);
xor U11148 (N_11148,N_7957,N_4362);
xnor U11149 (N_11149,N_3429,N_8488);
and U11150 (N_11150,N_7231,N_5405);
and U11151 (N_11151,N_6948,N_1227);
or U11152 (N_11152,N_547,N_8746);
or U11153 (N_11153,N_3734,N_8479);
nor U11154 (N_11154,N_4013,N_4620);
xnor U11155 (N_11155,N_8519,N_74);
nand U11156 (N_11156,N_8339,N_6986);
and U11157 (N_11157,N_5704,N_7035);
nand U11158 (N_11158,N_9944,N_3388);
xor U11159 (N_11159,N_3703,N_7746);
or U11160 (N_11160,N_7007,N_7541);
or U11161 (N_11161,N_8171,N_2832);
nor U11162 (N_11162,N_8565,N_8735);
and U11163 (N_11163,N_4997,N_4022);
nand U11164 (N_11164,N_2044,N_9020);
nand U11165 (N_11165,N_5929,N_3294);
or U11166 (N_11166,N_3566,N_8926);
nor U11167 (N_11167,N_415,N_8240);
nor U11168 (N_11168,N_9271,N_5871);
or U11169 (N_11169,N_233,N_8494);
nand U11170 (N_11170,N_9912,N_3191);
nand U11171 (N_11171,N_7902,N_942);
xnor U11172 (N_11172,N_6266,N_6824);
or U11173 (N_11173,N_9034,N_5584);
or U11174 (N_11174,N_1860,N_7218);
nor U11175 (N_11175,N_5562,N_1532);
or U11176 (N_11176,N_7030,N_9010);
or U11177 (N_11177,N_4699,N_1915);
or U11178 (N_11178,N_9276,N_1640);
or U11179 (N_11179,N_719,N_782);
or U11180 (N_11180,N_4041,N_7225);
xor U11181 (N_11181,N_9053,N_6176);
or U11182 (N_11182,N_8483,N_3709);
and U11183 (N_11183,N_9336,N_7548);
xnor U11184 (N_11184,N_6924,N_2942);
xnor U11185 (N_11185,N_9103,N_8624);
and U11186 (N_11186,N_1700,N_6000);
or U11187 (N_11187,N_7377,N_9369);
xnor U11188 (N_11188,N_5804,N_8533);
or U11189 (N_11189,N_5949,N_7963);
or U11190 (N_11190,N_844,N_3373);
xnor U11191 (N_11191,N_8215,N_7012);
nand U11192 (N_11192,N_5758,N_8577);
and U11193 (N_11193,N_4696,N_6349);
nor U11194 (N_11194,N_6792,N_6776);
and U11195 (N_11195,N_4582,N_5063);
nor U11196 (N_11196,N_9716,N_9772);
nor U11197 (N_11197,N_9938,N_4695);
nand U11198 (N_11198,N_1562,N_2519);
nand U11199 (N_11199,N_143,N_7990);
nand U11200 (N_11200,N_4839,N_9790);
nor U11201 (N_11201,N_8167,N_6900);
nor U11202 (N_11202,N_4598,N_269);
or U11203 (N_11203,N_9969,N_1730);
nor U11204 (N_11204,N_2011,N_5068);
nand U11205 (N_11205,N_7191,N_9110);
xor U11206 (N_11206,N_3090,N_9578);
xnor U11207 (N_11207,N_9229,N_691);
nor U11208 (N_11208,N_8463,N_2003);
xor U11209 (N_11209,N_8238,N_8450);
nand U11210 (N_11210,N_5757,N_4778);
and U11211 (N_11211,N_8157,N_1335);
nor U11212 (N_11212,N_9189,N_5948);
nand U11213 (N_11213,N_1450,N_5107);
or U11214 (N_11214,N_3267,N_2875);
nand U11215 (N_11215,N_5062,N_1471);
and U11216 (N_11216,N_2014,N_7325);
nor U11217 (N_11217,N_6104,N_3831);
or U11218 (N_11218,N_9688,N_6024);
nand U11219 (N_11219,N_2893,N_1480);
nand U11220 (N_11220,N_8665,N_5120);
nand U11221 (N_11221,N_814,N_7526);
and U11222 (N_11222,N_9267,N_8808);
xor U11223 (N_11223,N_812,N_5826);
xor U11224 (N_11224,N_6258,N_2480);
xnor U11225 (N_11225,N_5091,N_3524);
nand U11226 (N_11226,N_3695,N_7468);
or U11227 (N_11227,N_2580,N_550);
nand U11228 (N_11228,N_1970,N_419);
or U11229 (N_11229,N_5249,N_4783);
nand U11230 (N_11230,N_3702,N_4641);
and U11231 (N_11231,N_8573,N_2792);
xnor U11232 (N_11232,N_9233,N_4007);
nor U11233 (N_11233,N_6903,N_3032);
nor U11234 (N_11234,N_6425,N_6216);
nand U11235 (N_11235,N_2030,N_3903);
xnor U11236 (N_11236,N_9150,N_3606);
and U11237 (N_11237,N_6814,N_172);
nor U11238 (N_11238,N_7323,N_610);
or U11239 (N_11239,N_5258,N_9884);
and U11240 (N_11240,N_7171,N_4431);
xnor U11241 (N_11241,N_8981,N_3358);
nand U11242 (N_11242,N_1192,N_4255);
or U11243 (N_11243,N_5081,N_5745);
xnor U11244 (N_11244,N_7451,N_7008);
and U11245 (N_11245,N_7311,N_9768);
nor U11246 (N_11246,N_7375,N_7270);
nor U11247 (N_11247,N_8505,N_4893);
or U11248 (N_11248,N_8913,N_7143);
or U11249 (N_11249,N_7479,N_891);
or U11250 (N_11250,N_8489,N_2529);
nand U11251 (N_11251,N_38,N_2826);
nor U11252 (N_11252,N_2077,N_7503);
nor U11253 (N_11253,N_7969,N_9472);
or U11254 (N_11254,N_9303,N_1515);
xor U11255 (N_11255,N_9198,N_2274);
and U11256 (N_11256,N_1738,N_3898);
nor U11257 (N_11257,N_8225,N_584);
and U11258 (N_11258,N_4284,N_1386);
xnor U11259 (N_11259,N_558,N_1585);
and U11260 (N_11260,N_8406,N_7818);
and U11261 (N_11261,N_9083,N_4861);
and U11262 (N_11262,N_5555,N_9882);
nor U11263 (N_11263,N_6879,N_7205);
and U11264 (N_11264,N_7917,N_803);
nor U11265 (N_11265,N_4522,N_9463);
or U11266 (N_11266,N_1736,N_8060);
and U11267 (N_11267,N_3042,N_7584);
nor U11268 (N_11268,N_1332,N_9080);
nor U11269 (N_11269,N_1770,N_1109);
or U11270 (N_11270,N_920,N_6616);
nand U11271 (N_11271,N_4354,N_6895);
nand U11272 (N_11272,N_9807,N_5574);
xnor U11273 (N_11273,N_5727,N_2464);
nor U11274 (N_11274,N_4045,N_9723);
xnor U11275 (N_11275,N_5305,N_964);
or U11276 (N_11276,N_1753,N_7101);
nor U11277 (N_11277,N_6901,N_8898);
or U11278 (N_11278,N_1496,N_2752);
or U11279 (N_11279,N_9453,N_1513);
and U11280 (N_11280,N_6721,N_8791);
nand U11281 (N_11281,N_7465,N_7780);
nand U11282 (N_11282,N_2617,N_1383);
nor U11283 (N_11283,N_3287,N_3118);
nor U11284 (N_11284,N_8860,N_5853);
nor U11285 (N_11285,N_3672,N_1179);
or U11286 (N_11286,N_5210,N_6313);
or U11287 (N_11287,N_6411,N_4358);
or U11288 (N_11288,N_6143,N_1422);
and U11289 (N_11289,N_2337,N_9069);
nand U11290 (N_11290,N_3781,N_2644);
or U11291 (N_11291,N_7360,N_5809);
or U11292 (N_11292,N_9740,N_1956);
and U11293 (N_11293,N_3326,N_3268);
and U11294 (N_11294,N_6896,N_7847);
xnor U11295 (N_11295,N_1146,N_1725);
nand U11296 (N_11296,N_570,N_5882);
nor U11297 (N_11297,N_9196,N_1078);
xor U11298 (N_11298,N_4657,N_4675);
nand U11299 (N_11299,N_1488,N_7506);
nand U11300 (N_11300,N_8967,N_956);
nor U11301 (N_11301,N_9384,N_1030);
or U11302 (N_11302,N_6739,N_6711);
or U11303 (N_11303,N_2036,N_7247);
xor U11304 (N_11304,N_5459,N_4021);
or U11305 (N_11305,N_9673,N_7109);
nand U11306 (N_11306,N_5211,N_1022);
xnor U11307 (N_11307,N_3264,N_3732);
nor U11308 (N_11308,N_8426,N_6506);
xnor U11309 (N_11309,N_4683,N_2994);
and U11310 (N_11310,N_7904,N_518);
xor U11311 (N_11311,N_9863,N_5476);
or U11312 (N_11312,N_25,N_2531);
xnor U11313 (N_11313,N_3338,N_7802);
and U11314 (N_11314,N_6436,N_0);
or U11315 (N_11315,N_5449,N_6405);
nand U11316 (N_11316,N_7379,N_7195);
xnor U11317 (N_11317,N_284,N_5501);
or U11318 (N_11318,N_9771,N_6861);
nor U11319 (N_11319,N_5335,N_2028);
and U11320 (N_11320,N_4682,N_3411);
nand U11321 (N_11321,N_396,N_6031);
xnor U11322 (N_11322,N_3314,N_6243);
and U11323 (N_11323,N_5729,N_5626);
or U11324 (N_11324,N_171,N_2333);
nand U11325 (N_11325,N_9066,N_1913);
or U11326 (N_11326,N_6872,N_4410);
and U11327 (N_11327,N_1429,N_1308);
and U11328 (N_11328,N_8081,N_5239);
nand U11329 (N_11329,N_4853,N_7844);
and U11330 (N_11330,N_8645,N_7968);
and U11331 (N_11331,N_6186,N_1804);
nor U11332 (N_11332,N_4329,N_4240);
nand U11333 (N_11333,N_1419,N_2304);
nand U11334 (N_11334,N_5716,N_9921);
xnor U11335 (N_11335,N_1893,N_6335);
xor U11336 (N_11336,N_6836,N_4375);
or U11337 (N_11337,N_3514,N_8242);
or U11338 (N_11338,N_2549,N_9835);
nor U11339 (N_11339,N_3198,N_1682);
and U11340 (N_11340,N_2588,N_5749);
and U11341 (N_11341,N_6043,N_8619);
nand U11342 (N_11342,N_5667,N_6825);
xnor U11343 (N_11343,N_1181,N_3245);
nor U11344 (N_11344,N_1999,N_5730);
and U11345 (N_11345,N_2327,N_4324);
nand U11346 (N_11346,N_2345,N_9700);
or U11347 (N_11347,N_4381,N_5311);
or U11348 (N_11348,N_8005,N_8661);
nor U11349 (N_11349,N_1990,N_435);
or U11350 (N_11350,N_8969,N_2651);
nand U11351 (N_11351,N_8075,N_8699);
xnor U11352 (N_11352,N_6083,N_1810);
or U11353 (N_11353,N_7574,N_3252);
xor U11354 (N_11354,N_1735,N_8358);
nand U11355 (N_11355,N_4198,N_903);
xor U11356 (N_11356,N_1166,N_2272);
nand U11357 (N_11357,N_4875,N_5815);
nand U11358 (N_11358,N_398,N_4424);
nor U11359 (N_11359,N_9621,N_2266);
nor U11360 (N_11360,N_3378,N_9363);
nand U11361 (N_11361,N_889,N_9200);
or U11362 (N_11362,N_716,N_5480);
xor U11363 (N_11363,N_3554,N_9234);
xor U11364 (N_11364,N_745,N_1115);
and U11365 (N_11365,N_6548,N_7933);
nor U11366 (N_11366,N_3949,N_7700);
xor U11367 (N_11367,N_1938,N_2809);
xnor U11368 (N_11368,N_2005,N_215);
nand U11369 (N_11369,N_392,N_5677);
and U11370 (N_11370,N_4112,N_4681);
and U11371 (N_11371,N_4685,N_5234);
and U11372 (N_11372,N_9992,N_6474);
and U11373 (N_11373,N_8741,N_4473);
and U11374 (N_11374,N_9339,N_6418);
xor U11375 (N_11375,N_5157,N_9046);
nand U11376 (N_11376,N_3572,N_4809);
nor U11377 (N_11377,N_8039,N_7298);
xor U11378 (N_11378,N_8461,N_6028);
and U11379 (N_11379,N_2693,N_9459);
xnor U11380 (N_11380,N_5824,N_2545);
nor U11381 (N_11381,N_2864,N_4597);
xor U11382 (N_11382,N_2001,N_4063);
nand U11383 (N_11383,N_8226,N_1705);
and U11384 (N_11384,N_2926,N_8559);
nor U11385 (N_11385,N_3643,N_3892);
or U11386 (N_11386,N_191,N_1089);
xnor U11387 (N_11387,N_581,N_5783);
xor U11388 (N_11388,N_5528,N_3262);
xnor U11389 (N_11389,N_915,N_7454);
nor U11390 (N_11390,N_1541,N_6527);
nand U11391 (N_11391,N_8262,N_1923);
nor U11392 (N_11392,N_6804,N_4251);
or U11393 (N_11393,N_5112,N_9577);
or U11394 (N_11394,N_7115,N_4474);
nand U11395 (N_11395,N_3289,N_8842);
and U11396 (N_11396,N_7857,N_7711);
and U11397 (N_11397,N_7219,N_7031);
nand U11398 (N_11398,N_4828,N_3111);
xor U11399 (N_11399,N_7908,N_1111);
or U11400 (N_11400,N_9659,N_2774);
or U11401 (N_11401,N_40,N_2064);
and U11402 (N_11402,N_7835,N_1858);
nand U11403 (N_11403,N_1234,N_8070);
nand U11404 (N_11404,N_9403,N_7134);
xnor U11405 (N_11405,N_4732,N_3062);
and U11406 (N_11406,N_1023,N_7289);
or U11407 (N_11407,N_3626,N_4462);
or U11408 (N_11408,N_8693,N_9320);
and U11409 (N_11409,N_6933,N_2062);
nor U11410 (N_11410,N_7024,N_9645);
and U11411 (N_11411,N_4299,N_464);
and U11412 (N_11412,N_2088,N_8846);
xnor U11413 (N_11413,N_8408,N_6496);
nor U11414 (N_11414,N_6368,N_7617);
nor U11415 (N_11415,N_3265,N_901);
and U11416 (N_11416,N_8297,N_3101);
or U11417 (N_11417,N_1141,N_1465);
nand U11418 (N_11418,N_7027,N_1774);
or U11419 (N_11419,N_7462,N_2711);
or U11420 (N_11420,N_2596,N_9759);
nand U11421 (N_11421,N_2641,N_1880);
or U11422 (N_11422,N_5448,N_9097);
or U11423 (N_11423,N_4766,N_8546);
or U11424 (N_11424,N_686,N_6911);
or U11425 (N_11425,N_5937,N_6139);
xor U11426 (N_11426,N_4277,N_881);
or U11427 (N_11427,N_7588,N_5649);
nor U11428 (N_11428,N_1194,N_7663);
xor U11429 (N_11429,N_1692,N_1319);
nand U11430 (N_11430,N_4547,N_6127);
xor U11431 (N_11431,N_6570,N_9004);
or U11432 (N_11432,N_7614,N_9129);
nor U11433 (N_11433,N_7745,N_4364);
and U11434 (N_11434,N_9466,N_8017);
or U11435 (N_11435,N_2173,N_6947);
and U11436 (N_11436,N_997,N_7433);
or U11437 (N_11437,N_7960,N_2973);
nand U11438 (N_11438,N_5445,N_4388);
and U11439 (N_11439,N_7261,N_7114);
or U11440 (N_11440,N_1062,N_9122);
nor U11441 (N_11441,N_1764,N_4701);
and U11442 (N_11442,N_5991,N_5942);
nand U11443 (N_11443,N_9703,N_2240);
nand U11444 (N_11444,N_61,N_2746);
and U11445 (N_11445,N_8303,N_2613);
or U11446 (N_11446,N_3321,N_4533);
nor U11447 (N_11447,N_2830,N_7096);
or U11448 (N_11448,N_2786,N_8381);
and U11449 (N_11449,N_999,N_4330);
nand U11450 (N_11450,N_8071,N_6406);
nor U11451 (N_11451,N_1912,N_1528);
nand U11452 (N_11452,N_4231,N_8554);
or U11453 (N_11453,N_1452,N_3542);
and U11454 (N_11454,N_9913,N_4315);
xnor U11455 (N_11455,N_5031,N_352);
nor U11456 (N_11456,N_6265,N_7760);
nand U11457 (N_11457,N_5370,N_1791);
nor U11458 (N_11458,N_440,N_7598);
nand U11459 (N_11459,N_3452,N_9027);
nor U11460 (N_11460,N_6371,N_1954);
nand U11461 (N_11461,N_4632,N_4848);
or U11462 (N_11462,N_5379,N_5969);
nand U11463 (N_11463,N_7882,N_7155);
xor U11464 (N_11464,N_4847,N_8650);
nor U11465 (N_11465,N_899,N_9765);
nor U11466 (N_11466,N_2569,N_3423);
and U11467 (N_11467,N_3630,N_7727);
or U11468 (N_11468,N_4816,N_2899);
nand U11469 (N_11469,N_7733,N_1645);
or U11470 (N_11470,N_1066,N_9175);
or U11471 (N_11471,N_7604,N_520);
nand U11472 (N_11472,N_4726,N_9542);
or U11473 (N_11473,N_8856,N_6066);
or U11474 (N_11474,N_8792,N_8211);
xor U11475 (N_11475,N_9007,N_7556);
or U11476 (N_11476,N_4306,N_5784);
nor U11477 (N_11477,N_6062,N_9576);
and U11478 (N_11478,N_4791,N_9940);
nor U11479 (N_11479,N_2513,N_1768);
nor U11480 (N_11480,N_6191,N_2743);
nor U11481 (N_11481,N_8570,N_8374);
or U11482 (N_11482,N_3950,N_8298);
and U11483 (N_11483,N_1376,N_6059);
nor U11484 (N_11484,N_181,N_646);
and U11485 (N_11485,N_4308,N_7436);
xnor U11486 (N_11486,N_944,N_5095);
or U11487 (N_11487,N_7951,N_7687);
xor U11488 (N_11488,N_2736,N_9220);
nand U11489 (N_11489,N_2938,N_6008);
nand U11490 (N_11490,N_1612,N_2838);
and U11491 (N_11491,N_5648,N_2378);
xnor U11492 (N_11492,N_8607,N_7622);
xnor U11493 (N_11493,N_740,N_1381);
nand U11494 (N_11494,N_4243,N_8062);
and U11495 (N_11495,N_5843,N_4312);
and U11496 (N_11496,N_6446,N_1219);
xnor U11497 (N_11497,N_6678,N_5104);
nand U11498 (N_11498,N_6888,N_6357);
xor U11499 (N_11499,N_8727,N_5789);
or U11500 (N_11500,N_3224,N_8796);
xnor U11501 (N_11501,N_5565,N_222);
or U11502 (N_11502,N_6403,N_6959);
or U11503 (N_11503,N_2155,N_9803);
nor U11504 (N_11504,N_906,N_8235);
and U11505 (N_11505,N_1520,N_729);
or U11506 (N_11506,N_3023,N_8545);
nor U11507 (N_11507,N_6100,N_7342);
xor U11508 (N_11508,N_3094,N_7363);
xor U11509 (N_11509,N_1310,N_2586);
xnor U11510 (N_11510,N_6321,N_4331);
xor U11511 (N_11511,N_5983,N_1026);
nand U11512 (N_11512,N_5265,N_4976);
or U11513 (N_11513,N_116,N_667);
nand U11514 (N_11514,N_1114,N_9865);
nand U11515 (N_11515,N_8798,N_3509);
nand U11516 (N_11516,N_2148,N_7139);
and U11517 (N_11517,N_4952,N_4616);
nor U11518 (N_11518,N_5737,N_2253);
xor U11519 (N_11519,N_9423,N_7562);
xnor U11520 (N_11520,N_5161,N_5662);
and U11521 (N_11521,N_1829,N_5979);
xnor U11522 (N_11522,N_3158,N_7599);
nand U11523 (N_11523,N_7064,N_7532);
nor U11524 (N_11524,N_208,N_5415);
nor U11525 (N_11525,N_913,N_6376);
and U11526 (N_11526,N_2009,N_7630);
and U11527 (N_11527,N_6230,N_635);
nand U11528 (N_11528,N_5675,N_7291);
nor U11529 (N_11529,N_8341,N_6399);
nand U11530 (N_11530,N_5506,N_6904);
nand U11531 (N_11531,N_2418,N_806);
and U11532 (N_11532,N_638,N_3847);
or U11533 (N_11533,N_3821,N_5810);
and U11534 (N_11534,N_983,N_3409);
or U11535 (N_11535,N_8231,N_6708);
nand U11536 (N_11536,N_2620,N_7021);
or U11537 (N_11537,N_6151,N_2297);
xor U11538 (N_11538,N_8882,N_4047);
and U11539 (N_11539,N_5817,N_7664);
nor U11540 (N_11540,N_6360,N_1661);
nor U11541 (N_11541,N_3803,N_7376);
nor U11542 (N_11542,N_3196,N_4229);
or U11543 (N_11543,N_606,N_3179);
xnor U11544 (N_11544,N_6149,N_3914);
nor U11545 (N_11545,N_5310,N_929);
nand U11546 (N_11546,N_2294,N_6110);
or U11547 (N_11547,N_592,N_554);
and U11548 (N_11548,N_7177,N_9077);
and U11549 (N_11549,N_7160,N_2487);
nand U11550 (N_11550,N_6501,N_1438);
and U11551 (N_11551,N_2683,N_1247);
or U11552 (N_11552,N_6288,N_2659);
nand U11553 (N_11553,N_4503,N_1217);
and U11554 (N_11554,N_2024,N_7131);
xnor U11555 (N_11555,N_3468,N_5452);
xor U11556 (N_11556,N_8156,N_3603);
nand U11557 (N_11557,N_1399,N_5406);
or U11558 (N_11558,N_4305,N_322);
and U11559 (N_11559,N_462,N_6833);
or U11560 (N_11560,N_4443,N_6041);
nand U11561 (N_11561,N_9300,N_1636);
nor U11562 (N_11562,N_8476,N_3717);
or U11563 (N_11563,N_3859,N_5259);
nor U11564 (N_11564,N_4830,N_587);
and U11565 (N_11565,N_744,N_5578);
and U11566 (N_11566,N_6334,N_7762);
nand U11567 (N_11567,N_9574,N_3562);
or U11568 (N_11568,N_4416,N_9592);
xnor U11569 (N_11569,N_7689,N_3678);
or U11570 (N_11570,N_1898,N_3645);
nor U11571 (N_11571,N_7683,N_9426);
xor U11572 (N_11572,N_4700,N_4625);
xor U11573 (N_11573,N_1765,N_9331);
or U11574 (N_11574,N_6030,N_3582);
nand U11575 (N_11575,N_656,N_4365);
xor U11576 (N_11576,N_5386,N_1321);
or U11577 (N_11577,N_273,N_9202);
nor U11578 (N_11578,N_6488,N_8871);
or U11579 (N_11579,N_5101,N_7646);
and U11580 (N_11580,N_5713,N_2800);
nand U11581 (N_11581,N_9662,N_3065);
nand U11582 (N_11582,N_1427,N_8932);
xor U11583 (N_11583,N_3137,N_7547);
xnor U11584 (N_11584,N_9345,N_4245);
xor U11585 (N_11585,N_6304,N_1040);
nor U11586 (N_11586,N_7054,N_6742);
nand U11587 (N_11587,N_6431,N_1624);
nand U11588 (N_11588,N_6240,N_6519);
nand U11589 (N_11589,N_9082,N_1693);
nor U11590 (N_11590,N_1135,N_8578);
xnor U11591 (N_11591,N_184,N_2425);
nor U11592 (N_11592,N_6253,N_3908);
nor U11593 (N_11593,N_2721,N_9078);
or U11594 (N_11594,N_8678,N_5118);
and U11595 (N_11595,N_5158,N_783);
and U11596 (N_11596,N_8141,N_3116);
nor U11597 (N_11597,N_8478,N_1852);
xor U11598 (N_11598,N_6807,N_9440);
and U11599 (N_11599,N_476,N_1122);
and U11600 (N_11600,N_1190,N_209);
nor U11601 (N_11601,N_1372,N_6236);
nor U11602 (N_11602,N_5050,N_3840);
and U11603 (N_11603,N_3160,N_2202);
or U11604 (N_11604,N_8562,N_874);
nor U11605 (N_11605,N_9764,N_1267);
or U11606 (N_11606,N_4604,N_3406);
or U11607 (N_11607,N_7788,N_8036);
xor U11608 (N_11608,N_5726,N_412);
xnor U11609 (N_11609,N_865,N_6505);
or U11610 (N_11610,N_1733,N_6282);
or U11611 (N_11611,N_2102,N_19);
nand U11612 (N_11612,N_407,N_8223);
nor U11613 (N_11613,N_7994,N_4777);
xnor U11614 (N_11614,N_9337,N_261);
xor U11615 (N_11615,N_9599,N_9334);
nor U11616 (N_11616,N_4606,N_1680);
or U11617 (N_11617,N_4756,N_7111);
xor U11618 (N_11618,N_1746,N_5513);
nand U11619 (N_11619,N_6344,N_5641);
and U11620 (N_11620,N_1755,N_4333);
xor U11621 (N_11621,N_2757,N_3439);
nor U11622 (N_11622,N_7587,N_2236);
and U11623 (N_11623,N_1882,N_343);
or U11624 (N_11624,N_4954,N_2391);
nand U11625 (N_11625,N_6536,N_6445);
xor U11626 (N_11626,N_8828,N_7864);
nand U11627 (N_11627,N_9962,N_6789);
nand U11628 (N_11628,N_2047,N_6741);
nand U11629 (N_11629,N_7330,N_4593);
xnor U11630 (N_11630,N_8901,N_6112);
nor U11631 (N_11631,N_7920,N_7023);
nor U11632 (N_11632,N_9672,N_5205);
or U11633 (N_11633,N_7084,N_7065);
and U11634 (N_11634,N_5316,N_6160);
xnor U11635 (N_11635,N_9793,N_8850);
or U11636 (N_11636,N_7676,N_9496);
or U11637 (N_11637,N_1945,N_7146);
xnor U11638 (N_11638,N_7284,N_9252);
and U11639 (N_11639,N_7625,N_3349);
nand U11640 (N_11640,N_3758,N_6036);
and U11641 (N_11641,N_3103,N_227);
xor U11642 (N_11642,N_3320,N_7013);
nor U11643 (N_11643,N_4172,N_6936);
and U11644 (N_11644,N_8711,N_4558);
nor U11645 (N_11645,N_9920,N_6223);
and U11646 (N_11646,N_8055,N_9945);
or U11647 (N_11647,N_6689,N_4035);
xor U11648 (N_11648,N_2419,N_3767);
and U11649 (N_11649,N_9445,N_5354);
and U11650 (N_11650,N_7657,N_1150);
xnor U11651 (N_11651,N_6422,N_7701);
nand U11652 (N_11652,N_5517,N_5875);
nand U11653 (N_11653,N_7815,N_1844);
and U11654 (N_11654,N_8868,N_280);
nand U11655 (N_11655,N_7193,N_5146);
xnor U11656 (N_11656,N_305,N_5130);
and U11657 (N_11657,N_2141,N_8837);
nand U11658 (N_11658,N_1558,N_9054);
and U11659 (N_11659,N_1439,N_52);
or U11660 (N_11660,N_3184,N_6233);
nand U11661 (N_11661,N_8471,N_8049);
or U11662 (N_11662,N_5371,N_8414);
nor U11663 (N_11663,N_6315,N_6945);
nand U11664 (N_11664,N_9422,N_1407);
xnor U11665 (N_11665,N_4939,N_8175);
and U11666 (N_11666,N_6448,N_395);
xnor U11667 (N_11667,N_2634,N_2394);
nor U11668 (N_11668,N_3925,N_8787);
and U11669 (N_11669,N_1049,N_9079);
and U11670 (N_11670,N_1165,N_4804);
nand U11671 (N_11671,N_8382,N_8190);
nor U11672 (N_11672,N_955,N_3851);
nor U11673 (N_11673,N_5751,N_8525);
xnor U11674 (N_11674,N_8909,N_7898);
and U11675 (N_11675,N_536,N_1854);
nand U11676 (N_11676,N_2280,N_9393);
and U11677 (N_11677,N_1123,N_8728);
nand U11678 (N_11678,N_7890,N_9915);
and U11679 (N_11679,N_5772,N_3644);
xor U11680 (N_11680,N_6271,N_2065);
xnor U11681 (N_11681,N_3449,N_4036);
nor U11682 (N_11682,N_7976,N_9798);
xor U11683 (N_11683,N_8648,N_2072);
and U11684 (N_11684,N_4056,N_1016);
xnor U11685 (N_11685,N_4080,N_5638);
or U11686 (N_11686,N_4672,N_3646);
xnor U11687 (N_11687,N_7011,N_3420);
and U11688 (N_11688,N_9324,N_1337);
and U11689 (N_11689,N_8454,N_6293);
nand U11690 (N_11690,N_8305,N_7944);
nand U11691 (N_11691,N_8564,N_5132);
nand U11692 (N_11692,N_7450,N_5545);
nor U11693 (N_11693,N_2767,N_9984);
and U11694 (N_11694,N_5990,N_6810);
nor U11695 (N_11695,N_5330,N_9232);
and U11696 (N_11696,N_2250,N_9283);
xnor U11697 (N_11697,N_6533,N_5874);
nand U11698 (N_11698,N_9355,N_8656);
xnor U11699 (N_11699,N_7828,N_7805);
nand U11700 (N_11700,N_4453,N_9737);
nand U11701 (N_11701,N_5896,N_5198);
nand U11702 (N_11702,N_7691,N_7823);
or U11703 (N_11703,N_6816,N_3809);
nand U11704 (N_11704,N_438,N_5376);
or U11705 (N_11705,N_7868,N_7122);
nand U11706 (N_11706,N_5951,N_5390);
or U11707 (N_11707,N_9660,N_5542);
nor U11708 (N_11708,N_8587,N_1769);
nand U11709 (N_11709,N_2092,N_2152);
nor U11710 (N_11710,N_1997,N_5075);
nand U11711 (N_11711,N_2310,N_5905);
xor U11712 (N_11712,N_6130,N_6601);
or U11713 (N_11713,N_2477,N_1379);
or U11714 (N_11714,N_2082,N_3288);
and U11715 (N_11715,N_2362,N_9171);
nand U11716 (N_11716,N_701,N_5589);
nand U11717 (N_11717,N_8147,N_1922);
or U11718 (N_11718,N_3428,N_2234);
nor U11719 (N_11719,N_6080,N_3779);
and U11720 (N_11720,N_8405,N_5171);
nor U11721 (N_11721,N_8550,N_5916);
or U11722 (N_11722,N_2370,N_314);
and U11723 (N_11723,N_2920,N_3328);
nor U11724 (N_11724,N_8304,N_6512);
and U11725 (N_11725,N_3132,N_6806);
nand U11726 (N_11726,N_2801,N_5886);
nand U11727 (N_11727,N_3152,N_6005);
xnor U11728 (N_11728,N_5735,N_1177);
or U11729 (N_11729,N_4040,N_3512);
nor U11730 (N_11730,N_8709,N_3910);
nand U11731 (N_11731,N_126,N_4872);
nand U11732 (N_11732,N_5111,N_9830);
or U11733 (N_11733,N_5543,N_7979);
xor U11734 (N_11734,N_2329,N_2506);
and U11735 (N_11735,N_8970,N_4678);
xor U11736 (N_11736,N_3675,N_9008);
and U11737 (N_11737,N_8931,N_2551);
and U11738 (N_11738,N_231,N_3066);
nor U11739 (N_11739,N_3417,N_5167);
nor U11740 (N_11740,N_5835,N_8097);
and U11741 (N_11741,N_9213,N_3061);
and U11742 (N_11742,N_9435,N_3350);
and U11743 (N_11743,N_4235,N_1000);
and U11744 (N_11744,N_8596,N_2260);
and U11745 (N_11745,N_1167,N_9731);
or U11746 (N_11746,N_7488,N_4631);
and U11747 (N_11747,N_293,N_4595);
nor U11748 (N_11748,N_7000,N_9288);
and U11749 (N_11749,N_8622,N_4015);
nand U11750 (N_11750,N_593,N_5554);
or U11751 (N_11751,N_8023,N_7842);
nor U11752 (N_11752,N_4517,N_8306);
nor U11753 (N_11753,N_6951,N_3335);
or U11754 (N_11754,N_596,N_6791);
xor U11755 (N_11755,N_3228,N_3445);
nor U11756 (N_11756,N_3394,N_4002);
xnor U11757 (N_11757,N_9560,N_1564);
nor U11758 (N_11758,N_7876,N_404);
xor U11759 (N_11759,N_992,N_6675);
xor U11760 (N_11760,N_6114,N_3990);
xnor U11761 (N_11761,N_8485,N_2407);
xor U11762 (N_11762,N_8726,N_6680);
nor U11763 (N_11763,N_1609,N_3601);
nor U11764 (N_11764,N_4966,N_8137);
nand U11765 (N_11765,N_623,N_3664);
nand U11766 (N_11766,N_1571,N_4432);
and U11767 (N_11767,N_8561,N_1093);
xnor U11768 (N_11768,N_4182,N_5340);
nor U11769 (N_11769,N_5238,N_7523);
nand U11770 (N_11770,N_3731,N_8767);
nor U11771 (N_11771,N_6633,N_3590);
or U11772 (N_11772,N_2501,N_4933);
and U11773 (N_11773,N_410,N_5381);
xnor U11774 (N_11774,N_7553,N_9630);
nand U11775 (N_11775,N_5524,N_1203);
xnor U11776 (N_11776,N_7515,N_3431);
xor U11777 (N_11777,N_6392,N_6263);
xnor U11778 (N_11778,N_2104,N_8486);
and U11779 (N_11779,N_7743,N_9936);
or U11780 (N_11780,N_6628,N_3323);
nand U11781 (N_11781,N_958,N_902);
xor U11782 (N_11782,N_3282,N_2183);
nand U11783 (N_11783,N_6631,N_4968);
nor U11784 (N_11784,N_8977,N_182);
nor U11785 (N_11785,N_8085,N_8865);
or U11786 (N_11786,N_2600,N_7761);
nand U11787 (N_11787,N_9598,N_8218);
xor U11788 (N_11788,N_1083,N_1499);
or U11789 (N_11789,N_7004,N_1908);
and U11790 (N_11790,N_3217,N_8614);
xnor U11791 (N_11791,N_5277,N_5045);
nor U11792 (N_11792,N_5000,N_2342);
xnor U11793 (N_11793,N_846,N_7277);
or U11794 (N_11794,N_2843,N_6049);
or U11795 (N_11795,N_1354,N_4279);
xor U11796 (N_11796,N_1464,N_4724);
or U11797 (N_11797,N_8601,N_4738);
or U11798 (N_11798,N_5685,N_2401);
or U11799 (N_11799,N_3871,N_8196);
or U11800 (N_11800,N_4772,N_4055);
nand U11801 (N_11801,N_8911,N_3274);
nand U11802 (N_11802,N_1280,N_8683);
nor U11803 (N_11803,N_6332,N_2794);
and U11804 (N_11804,N_1044,N_6);
or U11805 (N_11805,N_503,N_4343);
nand U11806 (N_11806,N_5321,N_96);
nand U11807 (N_11807,N_9587,N_243);
nand U11808 (N_11808,N_2788,N_8210);
and U11809 (N_11809,N_539,N_9816);
or U11810 (N_11810,N_7419,N_6855);
nand U11811 (N_11811,N_8030,N_6058);
and U11812 (N_11812,N_6388,N_1130);
nand U11813 (N_11813,N_9000,N_9070);
nor U11814 (N_11814,N_8383,N_4451);
nand U11815 (N_11815,N_3492,N_4774);
xor U11816 (N_11816,N_5424,N_5444);
xor U11817 (N_11817,N_3049,N_4562);
xor U11818 (N_11818,N_513,N_5086);
nand U11819 (N_11819,N_9859,N_5125);
or U11820 (N_11820,N_5717,N_1263);
nor U11821 (N_11821,N_5671,N_5257);
nor U11822 (N_11822,N_2070,N_8074);
or U11823 (N_11823,N_6999,N_2156);
and U11824 (N_11824,N_9242,N_839);
xnor U11825 (N_11825,N_8336,N_2982);
or U11826 (N_11826,N_7660,N_5855);
xnor U11827 (N_11827,N_885,N_4924);
nor U11828 (N_11828,N_187,N_3688);
nand U11829 (N_11829,N_4951,N_1311);
nor U11830 (N_11830,N_1180,N_4003);
or U11831 (N_11831,N_9841,N_941);
or U11832 (N_11832,N_7748,N_5469);
nor U11833 (N_11833,N_3344,N_7426);
or U11834 (N_11834,N_3219,N_1300);
and U11835 (N_11835,N_8032,N_7266);
nand U11836 (N_11836,N_9407,N_8126);
nand U11837 (N_11837,N_4203,N_3594);
nor U11838 (N_11838,N_1861,N_7785);
nor U11839 (N_11839,N_7524,N_8416);
xnor U11840 (N_11840,N_8713,N_6397);
or U11841 (N_11841,N_3728,N_8004);
nand U11842 (N_11842,N_7136,N_8802);
nand U11843 (N_11843,N_9653,N_498);
or U11844 (N_11844,N_1832,N_1246);
or U11845 (N_11845,N_7509,N_1261);
xnor U11846 (N_11846,N_5770,N_3434);
nand U11847 (N_11847,N_2575,N_9344);
xor U11848 (N_11848,N_1255,N_35);
or U11849 (N_11849,N_366,N_5492);
and U11850 (N_11850,N_3557,N_8404);
xnor U11851 (N_11851,N_2898,N_3054);
xnor U11852 (N_11852,N_1879,N_2901);
nor U11853 (N_11853,N_5352,N_8203);
and U11854 (N_11854,N_6484,N_6874);
nor U11855 (N_11855,N_290,N_8737);
or U11856 (N_11856,N_4273,N_531);
and U11857 (N_11857,N_9301,N_8384);
and U11858 (N_11858,N_2769,N_6788);
nor U11859 (N_11859,N_4904,N_4490);
and U11860 (N_11860,N_3575,N_1676);
or U11861 (N_11861,N_7105,N_3745);
and U11862 (N_11862,N_6437,N_504);
xor U11863 (N_11863,N_6750,N_2522);
nand U11864 (N_11864,N_4010,N_728);
nor U11865 (N_11865,N_7061,N_9730);
nand U11866 (N_11866,N_1245,N_2797);
nor U11867 (N_11867,N_3741,N_6294);
nor U11868 (N_11868,N_4832,N_6821);
nand U11869 (N_11869,N_7226,N_2354);
or U11870 (N_11870,N_6898,N_8569);
or U11871 (N_11871,N_9420,N_6704);
nand U11872 (N_11872,N_8421,N_6560);
or U11873 (N_11873,N_1731,N_3107);
nor U11874 (N_11874,N_7927,N_5950);
and U11875 (N_11875,N_2962,N_9174);
nor U11876 (N_11876,N_7642,N_3145);
nor U11877 (N_11877,N_5255,N_218);
or U11878 (N_11878,N_6524,N_8841);
xnor U11879 (N_11879,N_8858,N_4840);
nor U11880 (N_11880,N_4218,N_5913);
or U11881 (N_11881,N_7265,N_830);
nand U11882 (N_11882,N_3599,N_3629);
and U11883 (N_11883,N_8732,N_2623);
xnor U11884 (N_11884,N_2971,N_8593);
xnor U11885 (N_11885,N_8455,N_3872);
and U11886 (N_11886,N_1432,N_5297);
nor U11887 (N_11887,N_3285,N_7198);
xor U11888 (N_11888,N_6636,N_5582);
or U11889 (N_11889,N_6279,N_6890);
or U11890 (N_11890,N_4834,N_7398);
xor U11891 (N_11891,N_4764,N_8499);
or U11892 (N_11892,N_5569,N_2267);
nor U11893 (N_11893,N_2504,N_8643);
xor U11894 (N_11894,N_6003,N_8602);
and U11895 (N_11895,N_2471,N_8230);
nand U11896 (N_11896,N_7680,N_3506);
nand U11897 (N_11897,N_7417,N_5036);
nor U11898 (N_11898,N_263,N_2244);
and U11899 (N_11899,N_1158,N_194);
or U11900 (N_11900,N_6220,N_9518);
or U11901 (N_11901,N_7995,N_7435);
xnor U11902 (N_11902,N_8325,N_1473);
nor U11903 (N_11903,N_6834,N_1762);
xor U11904 (N_11904,N_8390,N_7956);
xnor U11905 (N_11905,N_3014,N_534);
nor U11906 (N_11906,N_3638,N_6594);
nand U11907 (N_11907,N_767,N_3986);
or U11908 (N_11908,N_2389,N_1027);
nor U11909 (N_11909,N_3962,N_9532);
xor U11910 (N_11910,N_8172,N_4519);
nor U11911 (N_11911,N_8356,N_3761);
and U11912 (N_11912,N_9216,N_8927);
or U11913 (N_11913,N_8430,N_5963);
and U11914 (N_11914,N_8002,N_3930);
nand U11915 (N_11915,N_6170,N_192);
nor U11916 (N_11916,N_1482,N_5529);
and U11917 (N_11917,N_1740,N_8635);
and U11918 (N_11918,N_3292,N_5320);
nor U11919 (N_11919,N_8166,N_4136);
nand U11920 (N_11920,N_4349,N_3403);
nand U11921 (N_11921,N_9159,N_4574);
xor U11922 (N_11922,N_358,N_8807);
xor U11923 (N_11923,N_8255,N_7184);
nor U11924 (N_11924,N_2197,N_6097);
nand U11925 (N_11925,N_1147,N_5202);
nand U11926 (N_11926,N_8151,N_86);
and U11927 (N_11927,N_4300,N_6535);
and U11928 (N_11928,N_3367,N_5329);
and U11929 (N_11929,N_4377,N_3169);
nor U11930 (N_11930,N_9164,N_8943);
nand U11931 (N_11931,N_4142,N_9754);
and U11932 (N_11932,N_3171,N_7883);
or U11933 (N_11933,N_5696,N_2073);
xor U11934 (N_11934,N_1297,N_4624);
nor U11935 (N_11935,N_6622,N_7309);
nor U11936 (N_11936,N_3253,N_2365);
nand U11937 (N_11937,N_4592,N_5315);
nand U11938 (N_11938,N_3379,N_5945);
and U11939 (N_11939,N_2952,N_3913);
nor U11940 (N_11940,N_8277,N_837);
nand U11941 (N_11941,N_9487,N_9533);
nor U11942 (N_11942,N_6914,N_1225);
or U11943 (N_11943,N_6214,N_712);
xnor U11944 (N_11944,N_1851,N_2894);
nand U11945 (N_11945,N_1710,N_1894);
xnor U11946 (N_11946,N_2710,N_8201);
and U11947 (N_11947,N_3077,N_7185);
xor U11948 (N_11948,N_8676,N_4524);
nand U11949 (N_11949,N_1587,N_2347);
and U11950 (N_11950,N_2573,N_3751);
nand U11951 (N_11951,N_8854,N_8107);
and U11952 (N_11952,N_8492,N_8524);
xnor U11953 (N_11953,N_9315,N_2135);
xor U11954 (N_11954,N_2518,N_1012);
or U11955 (N_11955,N_8623,N_7953);
or U11956 (N_11956,N_1627,N_6503);
and U11957 (N_11957,N_960,N_1767);
xnor U11958 (N_11958,N_9687,N_5927);
or U11959 (N_11959,N_3402,N_7248);
or U11960 (N_11960,N_8712,N_8407);
or U11961 (N_11961,N_8386,N_5514);
nand U11962 (N_11962,N_9924,N_9063);
or U11963 (N_11963,N_7961,N_6734);
xnor U11964 (N_11964,N_7592,N_3747);
xor U11965 (N_11965,N_7408,N_8527);
nor U11966 (N_11966,N_7974,N_9450);
or U11967 (N_11967,N_5793,N_1492);
nand U11968 (N_11968,N_727,N_1631);
or U11969 (N_11969,N_1887,N_9889);
and U11970 (N_11970,N_7452,N_5092);
or U11971 (N_11971,N_1326,N_5364);
nor U11972 (N_11972,N_31,N_6342);
nor U11973 (N_11973,N_3398,N_6203);
and U11974 (N_11974,N_7502,N_7233);
nor U11975 (N_11975,N_1058,N_3771);
or U11976 (N_11976,N_4250,N_1750);
or U11977 (N_11977,N_5043,N_9776);
nor U11978 (N_11978,N_5404,N_5193);
and U11979 (N_11979,N_2215,N_3749);
and U11980 (N_11980,N_3290,N_1373);
and U11981 (N_11981,N_5183,N_7424);
nor U11982 (N_11982,N_739,N_4946);
nor U11983 (N_11983,N_6915,N_9179);
and U11984 (N_11984,N_2050,N_8475);
nor U11985 (N_11985,N_3617,N_7127);
and U11986 (N_11986,N_8742,N_4189);
or U11987 (N_11987,N_1950,N_2124);
nor U11988 (N_11988,N_875,N_4548);
nor U11989 (N_11989,N_2779,N_3584);
nor U11990 (N_11990,N_6993,N_8848);
and U11991 (N_11991,N_5994,N_142);
nor U11992 (N_11992,N_8103,N_6724);
nor U11993 (N_11993,N_3580,N_940);
nand U11994 (N_11994,N_6348,N_4898);
and U11995 (N_11995,N_4596,N_537);
xor U11996 (N_11996,N_2021,N_3309);
or U11997 (N_11997,N_5172,N_3844);
xor U11998 (N_11998,N_2074,N_320);
xnor U11999 (N_11999,N_6892,N_8473);
nor U12000 (N_12000,N_2972,N_5583);
and U12001 (N_12001,N_368,N_823);
nand U12002 (N_12002,N_7770,N_574);
and U12003 (N_12003,N_7654,N_946);
and U12004 (N_12004,N_1878,N_7306);
and U12005 (N_12005,N_6107,N_798);
nor U12006 (N_12006,N_1486,N_8045);
nand U12007 (N_12007,N_2904,N_1590);
or U12008 (N_12008,N_8418,N_5721);
nand U12009 (N_12009,N_8506,N_6077);
nand U12010 (N_12010,N_995,N_7301);
nand U12011 (N_12011,N_8113,N_2584);
nor U12012 (N_12012,N_4694,N_1099);
or U12013 (N_12013,N_6417,N_3135);
or U12014 (N_12014,N_7984,N_3128);
or U12015 (N_12015,N_5917,N_9695);
and U12016 (N_12016,N_585,N_73);
xnor U12017 (N_12017,N_4200,N_7387);
and U12018 (N_12018,N_7392,N_9619);
or U12019 (N_12019,N_472,N_2359);
and U12020 (N_12020,N_8161,N_4208);
nand U12021 (N_12021,N_6330,N_7643);
and U12022 (N_12022,N_5022,N_8216);
xnor U12023 (N_12023,N_7062,N_1749);
nand U12024 (N_12024,N_2350,N_5820);
nor U12025 (N_12025,N_9221,N_6620);
or U12026 (N_12026,N_1805,N_8034);
nand U12027 (N_12027,N_3397,N_4145);
and U12028 (N_12028,N_4881,N_4948);
and U12029 (N_12029,N_8521,N_2909);
and U12030 (N_12030,N_383,N_508);
xnor U12031 (N_12031,N_5416,N_3208);
xor U12032 (N_12032,N_6301,N_7399);
nor U12033 (N_12033,N_860,N_1270);
or U12034 (N_12034,N_5958,N_1398);
xnor U12035 (N_12035,N_1656,N_1412);
nand U12036 (N_12036,N_5278,N_8456);
and U12037 (N_12037,N_99,N_5114);
xnor U12038 (N_12038,N_2103,N_3240);
and U12039 (N_12039,N_2154,N_4194);
or U12040 (N_12040,N_2836,N_8073);
nor U12041 (N_12041,N_3278,N_6182);
and U12042 (N_12042,N_4185,N_5530);
nand U12043 (N_12043,N_311,N_5818);
nor U12044 (N_12044,N_1761,N_4529);
nor U12045 (N_12045,N_8138,N_8955);
xnor U12046 (N_12046,N_4436,N_8805);
and U12047 (N_12047,N_1208,N_1277);
nand U12048 (N_12048,N_7103,N_3046);
xnor U12049 (N_12049,N_8105,N_285);
xor U12050 (N_12050,N_7679,N_6886);
nor U12051 (N_12051,N_4127,N_5782);
or U12052 (N_12052,N_7486,N_6823);
or U12053 (N_12053,N_9581,N_2798);
xnor U12054 (N_12054,N_3783,N_481);
xor U12055 (N_12055,N_3970,N_4623);
nand U12056 (N_12056,N_2582,N_2111);
xor U12057 (N_12057,N_8197,N_7420);
or U12058 (N_12058,N_6703,N_2428);
nand U12059 (N_12059,N_7737,N_978);
xnor U12060 (N_12060,N_1260,N_9995);
and U12061 (N_12061,N_8185,N_1293);
xor U12062 (N_12062,N_7982,N_2966);
or U12063 (N_12063,N_8703,N_671);
nor U12064 (N_12064,N_2386,N_869);
nor U12065 (N_12065,N_3813,N_7731);
xnor U12066 (N_12066,N_9521,N_4906);
nor U12067 (N_12067,N_8780,N_4621);
and U12068 (N_12068,N_4921,N_631);
xor U12069 (N_12069,N_627,N_2461);
xnor U12070 (N_12070,N_1292,N_3477);
nand U12071 (N_12071,N_8966,N_3329);
xor U12072 (N_12072,N_4668,N_8192);
and U12073 (N_12073,N_163,N_479);
and U12074 (N_12074,N_7784,N_6201);
or U12075 (N_12075,N_9795,N_4638);
and U12076 (N_12076,N_4985,N_1886);
or U12077 (N_12077,N_4895,N_1659);
xnor U12078 (N_12078,N_710,N_1387);
nand U12079 (N_12079,N_5178,N_3296);
and U12080 (N_12080,N_6507,N_3720);
or U12081 (N_12081,N_2547,N_5504);
nor U12082 (N_12082,N_6447,N_6493);
and U12083 (N_12083,N_4546,N_7554);
and U12084 (N_12084,N_8734,N_8503);
or U12085 (N_12085,N_427,N_3661);
xor U12086 (N_12086,N_927,N_1621);
and U12087 (N_12087,N_9993,N_5856);
or U12088 (N_12088,N_5327,N_9706);
nand U12089 (N_12089,N_6746,N_6109);
nand U12090 (N_12090,N_7015,N_7852);
and U12091 (N_12091,N_381,N_5084);
and U12092 (N_12092,N_2652,N_3345);
or U12093 (N_12093,N_2503,N_2017);
nand U12094 (N_12094,N_9250,N_3009);
nand U12095 (N_12095,N_3316,N_1476);
xor U12096 (N_12096,N_5763,N_5778);
nand U12097 (N_12097,N_7840,N_7102);
xnor U12098 (N_12098,N_7641,N_736);
nand U12099 (N_12099,N_7949,N_9626);
xnor U12100 (N_12100,N_2834,N_6326);
or U12101 (N_12101,N_6250,N_7910);
xor U12102 (N_12102,N_7501,N_6756);
nor U12103 (N_12103,N_2595,N_8232);
and U12104 (N_12104,N_2544,N_4610);
and U12105 (N_12105,N_6038,N_3334);
xnor U12106 (N_12106,N_6974,N_7950);
nand U12107 (N_12107,N_3225,N_7407);
nand U12108 (N_12108,N_4842,N_9203);
nor U12109 (N_12109,N_8135,N_5844);
nand U12110 (N_12110,N_7936,N_5285);
nand U12111 (N_12111,N_2256,N_6607);
nor U12112 (N_12112,N_8866,N_9826);
nor U12113 (N_12113,N_2637,N_301);
nand U12114 (N_12114,N_1043,N_9611);
xor U12115 (N_12115,N_9447,N_7052);
nor U12116 (N_12116,N_3946,N_5199);
xnor U12117 (N_12117,N_1815,N_6899);
and U12118 (N_12118,N_8415,N_4860);
nor U12119 (N_12119,N_9140,N_6738);
and U12120 (N_12120,N_6006,N_3958);
and U12121 (N_12121,N_5419,N_108);
nand U12122 (N_12122,N_9101,N_1437);
nand U12123 (N_12123,N_7314,N_6200);
and U12124 (N_12124,N_7571,N_9057);
and U12125 (N_12125,N_55,N_4481);
or U12126 (N_12126,N_4589,N_7069);
xor U12127 (N_12127,N_4691,N_5168);
xnor U12128 (N_12128,N_7272,N_6995);
or U12129 (N_12129,N_5890,N_2380);
xor U12130 (N_12130,N_6489,N_2402);
nor U12131 (N_12131,N_6514,N_3205);
xor U12132 (N_12132,N_9876,N_9284);
nand U12133 (N_12133,N_2298,N_583);
or U12134 (N_12134,N_6785,N_1431);
or U12135 (N_12135,N_1239,N_1511);
xnor U12136 (N_12136,N_6359,N_9679);
xnor U12137 (N_12137,N_4280,N_8658);
nor U12138 (N_12138,N_288,N_8309);
nand U12139 (N_12139,N_8367,N_5690);
or U12140 (N_12140,N_103,N_5338);
or U12141 (N_12141,N_2270,N_9867);
and U12142 (N_12142,N_2922,N_5515);
or U12143 (N_12143,N_3089,N_3708);
or U12144 (N_12144,N_5215,N_4328);
or U12145 (N_12145,N_3824,N_3770);
nor U12146 (N_12146,N_9617,N_2616);
xnor U12147 (N_12147,N_7946,N_9359);
xor U12148 (N_12148,N_822,N_4873);
nand U12149 (N_12149,N_3591,N_1307);
and U12150 (N_12150,N_6796,N_1783);
xor U12151 (N_12151,N_9148,N_6564);
nand U12152 (N_12152,N_2823,N_8542);
and U12153 (N_12153,N_5788,N_2206);
and U12154 (N_12154,N_9415,N_8308);
xor U12155 (N_12155,N_8914,N_9116);
nor U12156 (N_12156,N_2006,N_6074);
nand U12157 (N_12157,N_2376,N_1577);
nor U12158 (N_12158,N_6384,N_9147);
or U12159 (N_12159,N_6072,N_8490);
xor U12160 (N_12160,N_6175,N_9512);
and U12161 (N_12161,N_1075,N_8803);
and U12162 (N_12162,N_5014,N_4126);
nand U12163 (N_12163,N_7914,N_7752);
nor U12164 (N_12164,N_2084,N_9071);
and U12165 (N_12165,N_2478,N_4030);
or U12166 (N_12166,N_9456,N_797);
or U12167 (N_12167,N_7492,N_8582);
nor U12168 (N_12168,N_7624,N_857);
nor U12169 (N_12169,N_1786,N_2608);
nand U12170 (N_12170,N_4899,N_1616);
nand U12171 (N_12171,N_6026,N_5924);
nor U12172 (N_12172,N_7896,N_1363);
and U12173 (N_12173,N_3926,N_4677);
and U12174 (N_12174,N_2458,N_5365);
or U12175 (N_12175,N_6396,N_6856);
nand U12176 (N_12176,N_9844,N_6542);
and U12177 (N_12177,N_2984,N_9441);
nand U12178 (N_12178,N_5389,N_2687);
or U12179 (N_12179,N_1015,N_1170);
nor U12180 (N_12180,N_9966,N_447);
nor U12181 (N_12181,N_2775,N_5560);
nand U12182 (N_12182,N_6588,N_5932);
or U12183 (N_12183,N_8180,N_9188);
xnor U12184 (N_12184,N_1313,N_2591);
xnor U12185 (N_12185,N_5231,N_2730);
nand U12186 (N_12186,N_8775,N_4953);
and U12187 (N_12187,N_639,N_1405);
nor U12188 (N_12188,N_6589,N_3712);
xnor U12189 (N_12189,N_1264,N_6372);
xor U12190 (N_12190,N_4079,N_9238);
nor U12191 (N_12191,N_2174,N_4098);
nor U12192 (N_12192,N_6600,N_626);
xor U12193 (N_12193,N_2426,N_1772);
nor U12194 (N_12194,N_6178,N_866);
nand U12195 (N_12195,N_2385,N_1266);
xnor U12196 (N_12196,N_7899,N_9684);
xor U12197 (N_12197,N_7251,N_6254);
nand U12198 (N_12198,N_5345,N_3164);
and U12199 (N_12199,N_1928,N_9093);
nand U12200 (N_12200,N_6404,N_4106);
nand U12201 (N_12201,N_1117,N_4599);
nand U12202 (N_12202,N_1704,N_9492);
nand U12203 (N_12203,N_7841,N_8824);
or U12204 (N_12204,N_4876,N_1242);
nor U12205 (N_12205,N_8667,N_9201);
and U12206 (N_12206,N_2002,N_4084);
nor U12207 (N_12207,N_3635,N_3754);
nand U12208 (N_12208,N_8755,N_2194);
and U12209 (N_12209,N_7989,N_4573);
xnor U12210 (N_12210,N_7076,N_3163);
nand U12211 (N_12211,N_2230,N_4177);
or U12212 (N_12212,N_7551,N_7568);
xnor U12213 (N_12213,N_3012,N_8195);
or U12214 (N_12214,N_9947,N_3971);
nor U12215 (N_12215,N_6295,N_8331);
nand U12216 (N_12216,N_2022,N_1067);
and U12217 (N_12217,N_6256,N_4930);
xor U12218 (N_12218,N_3997,N_6068);
and U12219 (N_12219,N_732,N_3924);
xnor U12220 (N_12220,N_6599,N_3456);
and U12221 (N_12221,N_7287,N_7332);
or U12222 (N_12222,N_5139,N_693);
xor U12223 (N_12223,N_7786,N_1329);
nand U12224 (N_12224,N_1315,N_4400);
or U12225 (N_12225,N_1697,N_1414);
nand U12226 (N_12226,N_6328,N_9910);
nand U12227 (N_12227,N_3982,N_3819);
nand U12228 (N_12228,N_4817,N_6064);
and U12229 (N_12229,N_8902,N_6222);
and U12230 (N_12230,N_1611,N_2991);
and U12231 (N_12231,N_8949,N_3227);
xnor U12232 (N_12232,N_8344,N_1522);
xor U12233 (N_12233,N_8563,N_579);
and U12234 (N_12234,N_3242,N_5650);
or U12235 (N_12235,N_8412,N_6215);
or U12236 (N_12236,N_7234,N_859);
xnor U12237 (N_12237,N_1393,N_6485);
nand U12238 (N_12238,N_805,N_5600);
or U12239 (N_12239,N_1220,N_5594);
nand U12240 (N_12240,N_827,N_7371);
or U12241 (N_12241,N_1087,N_4287);
nand U12242 (N_12242,N_8061,N_4934);
and U12243 (N_12243,N_7335,N_9149);
xnor U12244 (N_12244,N_8007,N_5175);
nand U12245 (N_12245,N_7651,N_6510);
nor U12246 (N_12246,N_7645,N_5920);
or U12247 (N_12247,N_909,N_8663);
xor U12248 (N_12248,N_255,N_8076);
xor U12249 (N_12249,N_7732,N_3736);
xor U12250 (N_12250,N_3953,N_5718);
xnor U12251 (N_12251,N_8574,N_1524);
xnor U12252 (N_12252,N_8887,N_228);
and U12253 (N_12253,N_299,N_5418);
xor U12254 (N_12254,N_8150,N_8311);
nor U12255 (N_12255,N_3829,N_4545);
nand U12256 (N_12256,N_3875,N_2656);
nor U12257 (N_12257,N_4211,N_8123);
and U12258 (N_12258,N_7605,N_7263);
xnor U12259 (N_12259,N_5227,N_3275);
nor U12260 (N_12260,N_861,N_9180);
and U12261 (N_12261,N_1742,N_8422);
nand U12262 (N_12262,N_1050,N_3605);
and U12263 (N_12263,N_1152,N_5720);
xnor U12264 (N_12264,N_7442,N_6629);
and U12265 (N_12265,N_3585,N_3086);
nand U12266 (N_12266,N_9048,N_160);
xnor U12267 (N_12267,N_6575,N_9290);
nor U12268 (N_12268,N_3255,N_7699);
or U12269 (N_12269,N_4334,N_16);
nand U12270 (N_12270,N_7353,N_9421);
nor U12271 (N_12271,N_7413,N_2398);
nor U12272 (N_12272,N_5665,N_1646);
nand U12273 (N_12273,N_7416,N_9163);
xnor U12274 (N_12274,N_2080,N_3112);
nor U12275 (N_12275,N_9639,N_8329);
or U12276 (N_12276,N_5541,N_1444);
and U12277 (N_12277,N_514,N_2489);
and U12278 (N_12278,N_2570,N_8051);
nand U12279 (N_12279,N_4409,N_8538);
or U12280 (N_12280,N_7273,N_4217);
nor U12281 (N_12281,N_7041,N_5348);
nand U12282 (N_12282,N_374,N_9715);
or U12283 (N_12283,N_7669,N_115);
nor U12284 (N_12284,N_5189,N_8057);
or U12285 (N_12285,N_8011,N_9437);
xor U12286 (N_12286,N_6340,N_9192);
nor U12287 (N_12287,N_7712,N_1342);
xor U12288 (N_12288,N_3057,N_2085);
or U12289 (N_12289,N_7656,N_4583);
nand U12290 (N_12290,N_4161,N_9028);
xnor U12291 (N_12291,N_5003,N_8999);
nand U12292 (N_12292,N_4971,N_4697);
nand U12293 (N_12293,N_2780,N_5180);
or U12294 (N_12294,N_8983,N_2013);
and U12295 (N_12295,N_7507,N_7125);
nand U12296 (N_12296,N_7110,N_1773);
xor U12297 (N_12297,N_6650,N_9701);
or U12298 (N_12298,N_5634,N_895);
nand U12299 (N_12299,N_3427,N_591);
nor U12300 (N_12300,N_8820,N_6504);
nand U12301 (N_12301,N_5235,N_1059);
nand U12302 (N_12302,N_5194,N_551);
xnor U12303 (N_12303,N_8206,N_347);
nand U12304 (N_12304,N_815,N_327);
and U12305 (N_12305,N_275,N_4643);
nand U12306 (N_12306,N_4698,N_4580);
or U12307 (N_12307,N_8063,N_7092);
nor U12308 (N_12308,N_4460,N_5402);
or U12309 (N_12309,N_2086,N_4252);
or U12310 (N_12310,N_1615,N_2413);
nand U12311 (N_12311,N_5295,N_7929);
xnor U12312 (N_12312,N_966,N_5901);
or U12313 (N_12313,N_1603,N_6204);
and U12314 (N_12314,N_684,N_2093);
nand U12315 (N_12315,N_763,N_372);
and U12316 (N_12316,N_868,N_746);
and U12317 (N_12317,N_2556,N_5643);
nand U12318 (N_12318,N_5766,N_7216);
nor U12319 (N_12319,N_5026,N_7355);
xor U12320 (N_12320,N_8425,N_6029);
or U12321 (N_12321,N_7157,N_5096);
and U12322 (N_12322,N_505,N_2026);
nand U12323 (N_12323,N_4248,N_7928);
nand U12324 (N_12324,N_5454,N_7739);
and U12325 (N_12325,N_9294,N_8273);
and U12326 (N_12326,N_7650,N_7621);
nand U12327 (N_12327,N_9757,N_6284);
nor U12328 (N_12328,N_102,N_7667);
nand U12329 (N_12329,N_8189,N_456);
and U12330 (N_12330,N_5613,N_8761);
nand U12331 (N_12331,N_245,N_5071);
or U12332 (N_12332,N_3837,N_7132);
nand U12333 (N_12333,N_7180,N_8047);
nor U12334 (N_12334,N_3127,N_9502);
or U12335 (N_12335,N_8462,N_9306);
or U12336 (N_12336,N_5470,N_1987);
nand U12337 (N_12337,N_2765,N_6386);
xnor U12338 (N_12338,N_6905,N_4313);
or U12339 (N_12339,N_5441,N_5780);
nand U12340 (N_12340,N_1876,N_457);
or U12341 (N_12341,N_7705,N_4162);
xor U12342 (N_12342,N_4356,N_1352);
xnor U12343 (N_12343,N_6380,N_223);
nor U12344 (N_12344,N_2658,N_9259);
and U12345 (N_12345,N_2696,N_3992);
nand U12346 (N_12346,N_7583,N_3756);
and U12347 (N_12347,N_4851,N_9977);
or U12348 (N_12348,N_7093,N_9509);
nor U12349 (N_12349,N_18,N_7);
and U12350 (N_12350,N_8973,N_6319);
nand U12351 (N_12351,N_648,N_1973);
nand U12352 (N_12352,N_1566,N_5872);
nor U12353 (N_12353,N_6581,N_2554);
nand U12354 (N_12354,N_9085,N_9089);
xnor U12355 (N_12355,N_7581,N_6333);
and U12356 (N_12356,N_2541,N_6557);
or U12357 (N_12357,N_576,N_1856);
nor U12358 (N_12358,N_9045,N_8144);
nor U12359 (N_12359,N_6076,N_339);
or U12360 (N_12360,N_2330,N_1578);
nand U12361 (N_12361,N_2469,N_9932);
xnor U12362 (N_12362,N_9039,N_8907);
xor U12363 (N_12363,N_8616,N_1924);
and U12364 (N_12364,N_3223,N_4319);
or U12365 (N_12365,N_89,N_1563);
and U12366 (N_12366,N_2916,N_3869);
or U12367 (N_12367,N_6733,N_9338);
and U12368 (N_12368,N_3974,N_5359);
and U12369 (N_12369,N_4183,N_7152);
xnor U12370 (N_12370,N_9380,N_4044);
or U12371 (N_12371,N_6757,N_8377);
nor U12372 (N_12372,N_4092,N_7339);
nand U12373 (N_12373,N_2574,N_1966);
xnor U12374 (N_12374,N_1454,N_5965);
or U12375 (N_12375,N_9858,N_9058);
and U12376 (N_12376,N_9335,N_3016);
nor U12377 (N_12377,N_8194,N_6412);
nand U12378 (N_12378,N_203,N_5624);
xor U12379 (N_12379,N_240,N_496);
and U12380 (N_12380,N_2163,N_4750);
nand U12381 (N_12381,N_4977,N_6336);
nor U12382 (N_12382,N_246,N_773);
nand U12383 (N_12383,N_3920,N_3547);
xnor U12384 (N_12384,N_4988,N_9885);
and U12385 (N_12385,N_3773,N_3942);
xnor U12386 (N_12386,N_6681,N_2353);
and U12387 (N_12387,N_5197,N_1642);
or U12388 (N_12388,N_4332,N_8125);
nand U12389 (N_12389,N_9049,N_3142);
xor U12390 (N_12390,N_3835,N_735);
xor U12391 (N_12391,N_1204,N_1294);
nor U12392 (N_12392,N_7794,N_9664);
nor U12393 (N_12393,N_8584,N_4800);
xor U12394 (N_12394,N_3877,N_8681);
nor U12395 (N_12395,N_8284,N_957);
nand U12396 (N_12396,N_7686,N_8880);
nand U12397 (N_12397,N_7401,N_5246);
or U12398 (N_12398,N_2744,N_9314);
xor U12399 (N_12399,N_2405,N_6705);
nor U12400 (N_12400,N_6387,N_4173);
and U12401 (N_12401,N_2012,N_4581);
and U12402 (N_12402,N_1968,N_4776);
xor U12403 (N_12403,N_8066,N_179);
nand U12404 (N_12404,N_692,N_6221);
and U12405 (N_12405,N_2536,N_9762);
xnor U12406 (N_12406,N_792,N_2415);
nor U12407 (N_12407,N_9809,N_7312);
and U12408 (N_12408,N_6764,N_8543);
nor U12409 (N_12409,N_5153,N_5827);
and U12410 (N_12410,N_8170,N_747);
xor U12411 (N_12411,N_9469,N_8067);
or U12412 (N_12412,N_5279,N_2432);
nor U12413 (N_12413,N_2015,N_7754);
and U12414 (N_12414,N_5190,N_7357);
nand U12415 (N_12415,N_5356,N_9286);
xnor U12416 (N_12416,N_8222,N_5317);
xnor U12417 (N_12417,N_1222,N_3495);
xor U12418 (N_12418,N_9113,N_9130);
xor U12419 (N_12419,N_3100,N_8413);
xnor U12420 (N_12420,N_2325,N_85);
or U12421 (N_12421,N_6118,N_5143);
nor U12422 (N_12422,N_1240,N_2667);
or U12423 (N_12423,N_2763,N_5861);
and U12424 (N_12424,N_9205,N_5612);
nand U12425 (N_12425,N_5805,N_158);
nand U12426 (N_12426,N_6714,N_5351);
xnor U12427 (N_12427,N_6400,N_1727);
and U12428 (N_12428,N_2799,N_300);
nand U12429 (N_12429,N_6780,N_8019);
and U12430 (N_12430,N_2716,N_8131);
nor U12431 (N_12431,N_4869,N_9890);
or U12432 (N_12432,N_1942,N_548);
and U12433 (N_12433,N_7239,N_8613);
and U12434 (N_12434,N_3360,N_8100);
xor U12435 (N_12435,N_7126,N_5010);
or U12436 (N_12436,N_308,N_7516);
or U12437 (N_12437,N_5659,N_3232);
xnor U12438 (N_12438,N_7776,N_3166);
and U12439 (N_12439,N_3497,N_4730);
nor U12440 (N_12440,N_2439,N_1789);
nor U12441 (N_12441,N_3331,N_8861);
xnor U12442 (N_12442,N_9391,N_1436);
xor U12443 (N_12443,N_2466,N_7224);
xor U12444 (N_12444,N_2131,N_9253);
nor U12445 (N_12445,N_437,N_4206);
or U12446 (N_12446,N_2316,N_3068);
or U12447 (N_12447,N_5319,N_5392);
or U12448 (N_12448,N_4629,N_4888);
or U12449 (N_12449,N_1312,N_4102);
or U12450 (N_12450,N_1073,N_1781);
and U12451 (N_12451,N_1390,N_2076);
nand U12452 (N_12452,N_9556,N_4707);
xor U12453 (N_12453,N_7412,N_7326);
nand U12454 (N_12454,N_488,N_9661);
nand U12455 (N_12455,N_6189,N_7958);
and U12456 (N_12456,N_4199,N_4786);
nor U12457 (N_12457,N_5417,N_8204);
nor U12458 (N_12458,N_1163,N_6940);
nand U12459 (N_12459,N_7992,N_7428);
xnor U12460 (N_12460,N_3038,N_92);
nor U12461 (N_12461,N_7912,N_3700);
xor U12462 (N_12462,N_4064,N_411);
or U12463 (N_12463,N_6800,N_5147);
xor U12464 (N_12464,N_7808,N_1449);
or U12465 (N_12465,N_9967,N_3842);
or U12466 (N_12466,N_993,N_8184);
nand U12467 (N_12467,N_7228,N_6194);
or U12468 (N_12468,N_4608,N_4101);
nand U12469 (N_12469,N_6994,N_9689);
nor U12470 (N_12470,N_2636,N_5489);
nand U12471 (N_12471,N_9227,N_1224);
xor U12472 (N_12472,N_9897,N_5282);
nand U12473 (N_12473,N_4437,N_6955);
and U12474 (N_12474,N_9680,N_5425);
or U12475 (N_12475,N_165,N_8752);
and U12476 (N_12476,N_3277,N_5823);
nand U12477 (N_12477,N_8776,N_6169);
and U12478 (N_12478,N_3623,N_7059);
nand U12479 (N_12479,N_3151,N_225);
or U12480 (N_12480,N_951,N_4894);
or U12481 (N_12481,N_1819,N_6812);
xnor U12482 (N_12482,N_1424,N_769);
and U12483 (N_12483,N_2043,N_3546);
and U12484 (N_12484,N_8077,N_9978);
nor U12485 (N_12485,N_1925,N_4342);
nor U12486 (N_12486,N_2738,N_6442);
or U12487 (N_12487,N_2737,N_6289);
xor U12488 (N_12488,N_6698,N_4406);
or U12489 (N_12489,N_9235,N_8327);
nor U12490 (N_12490,N_2331,N_1978);
nand U12491 (N_12491,N_8027,N_4827);
nand U12492 (N_12492,N_6819,N_5346);
xor U12493 (N_12493,N_9506,N_5802);
nor U12494 (N_12494,N_3102,N_1569);
or U12495 (N_12495,N_9812,N_7095);
xnor U12496 (N_12496,N_854,N_8043);
or U12497 (N_12497,N_6421,N_5274);
nand U12498 (N_12498,N_6238,N_5919);
xnor U12499 (N_12499,N_5858,N_125);
or U12500 (N_12500,N_7889,N_9546);
nand U12501 (N_12501,N_5047,N_8611);
xnor U12502 (N_12502,N_9784,N_8950);
xnor U12503 (N_12503,N_7255,N_3256);
nand U12504 (N_12504,N_9525,N_7725);
and U12505 (N_12505,N_4655,N_9274);
nor U12506 (N_12506,N_9744,N_4710);
xor U12507 (N_12507,N_2490,N_2886);
nand U12508 (N_12508,N_9106,N_1718);
nor U12509 (N_12509,N_6052,N_7695);
or U12510 (N_12510,N_3342,N_4868);
nand U12511 (N_12511,N_8696,N_4297);
and U12512 (N_12512,N_7637,N_8986);
nor U12513 (N_12513,N_4411,N_247);
or U12514 (N_12514,N_7418,N_2993);
nand U12515 (N_12515,N_1592,N_699);
or U12516 (N_12516,N_1348,N_9834);
xor U12517 (N_12517,N_9325,N_8397);
xor U12518 (N_12518,N_6775,N_9954);
xnor U12519 (N_12519,N_4213,N_342);
or U12520 (N_12520,N_4433,N_49);
or U12521 (N_12521,N_248,N_1837);
or U12522 (N_12522,N_90,N_5895);
nor U12523 (N_12523,N_1028,N_6257);
nand U12524 (N_12524,N_8886,N_1681);
and U12525 (N_12525,N_9930,N_1324);
and U12526 (N_12526,N_6298,N_9549);
nand U12527 (N_12527,N_7333,N_1126);
xor U12528 (N_12528,N_6269,N_2149);
xnor U12529 (N_12529,N_2997,N_1576);
nor U12530 (N_12530,N_4483,N_2423);
nor U12531 (N_12531,N_8875,N_8536);
or U12532 (N_12532,N_5149,N_2925);
or U12533 (N_12533,N_7692,N_894);
nor U12534 (N_12534,N_3516,N_175);
nor U12535 (N_12535,N_3079,N_9736);
nand U12536 (N_12536,N_788,N_3212);
xnor U12537 (N_12537,N_9483,N_6161);
xnor U12538 (N_12538,N_4158,N_7988);
or U12539 (N_12539,N_5134,N_120);
and U12540 (N_12540,N_6355,N_1584);
or U12541 (N_12541,N_3401,N_9818);
nand U12542 (N_12542,N_7831,N_8992);
and U12543 (N_12543,N_8788,N_5057);
nand U12544 (N_12544,N_1131,N_4845);
nand U12545 (N_12545,N_2008,N_1847);
or U12546 (N_12546,N_8654,N_2825);
or U12547 (N_12547,N_5039,N_6546);
nor U12548 (N_12548,N_8747,N_1620);
xor U12549 (N_12549,N_9458,N_9481);
xor U12550 (N_12550,N_3868,N_3880);
xor U12551 (N_12551,N_8181,N_3793);
or U12552 (N_12552,N_1613,N_9522);
or U12553 (N_12553,N_4822,N_4584);
nor U12554 (N_12554,N_9368,N_5005);
nand U12555 (N_12555,N_4093,N_5342);
and U12556 (N_12556,N_3459,N_4736);
and U12557 (N_12557,N_8026,N_5034);
or U12558 (N_12558,N_3530,N_5229);
nand U12559 (N_12559,N_922,N_4393);
or U12560 (N_12560,N_9991,N_7201);
xnor U12561 (N_12561,N_6449,N_649);
nor U12562 (N_12562,N_3322,N_238);
xnor U12563 (N_12563,N_8243,N_4765);
nand U12564 (N_12564,N_2955,N_373);
and U12565 (N_12565,N_5635,N_2233);
and U12566 (N_12566,N_9827,N_6727);
and U12567 (N_12567,N_4191,N_2219);
xnor U12568 (N_12568,N_4741,N_9448);
nand U12569 (N_12569,N_1694,N_449);
nand U12570 (N_12570,N_8639,N_6179);
nor U12571 (N_12571,N_5066,N_4391);
nand U12572 (N_12572,N_996,N_7199);
xnor U12573 (N_12573,N_1747,N_4429);
nand U12574 (N_12574,N_5186,N_695);
and U12575 (N_12575,N_5999,N_8736);
nand U12576 (N_12576,N_1897,N_4260);
nand U12577 (N_12577,N_153,N_5620);
nand U12578 (N_12578,N_7397,N_8823);
xor U12579 (N_12579,N_1455,N_968);
nand U12580 (N_12580,N_8531,N_1041);
or U12581 (N_12581,N_9799,N_9752);
or U12582 (N_12582,N_3476,N_6909);
nor U12583 (N_12583,N_5597,N_7940);
xnor U12584 (N_12584,N_5630,N_5923);
xnor U12585 (N_12585,N_2862,N_628);
or U12586 (N_12586,N_934,N_4858);
or U12587 (N_12587,N_604,N_1873);
and U12588 (N_12588,N_9241,N_8818);
nand U12589 (N_12589,N_4559,N_7697);
nor U12590 (N_12590,N_9837,N_1944);
or U12591 (N_12591,N_3796,N_7315);
nand U12592 (N_12592,N_4132,N_5746);
and U12593 (N_12593,N_3018,N_2846);
nor U12594 (N_12594,N_9214,N_8893);
nand U12595 (N_12595,N_2882,N_7825);
xor U12596 (N_12596,N_7550,N_2383);
or U12597 (N_12597,N_8919,N_9582);
nand U12598 (N_12598,N_7168,N_6923);
or U12599 (N_12599,N_6122,N_5941);
or U12600 (N_12600,N_7303,N_761);
and U12601 (N_12601,N_1795,N_3777);
nor U12602 (N_12602,N_555,N_502);
nand U12603 (N_12603,N_441,N_5242);
xor U12604 (N_12604,N_9553,N_6098);
or U12605 (N_12605,N_9051,N_4792);
xnor U12606 (N_12606,N_5223,N_1301);
nand U12607 (N_12607,N_2707,N_1421);
nor U12608 (N_12608,N_303,N_1961);
nor U12609 (N_12609,N_9510,N_566);
or U12610 (N_12610,N_9146,N_4810);
xnor U12611 (N_12611,N_9279,N_309);
or U12612 (N_12612,N_2229,N_6719);
xnor U12613 (N_12613,N_2745,N_8689);
nand U12614 (N_12614,N_7347,N_1216);
xor U12615 (N_12615,N_2911,N_898);
xnor U12616 (N_12616,N_7368,N_6604);
and U12617 (N_12617,N_3987,N_6291);
nand U12618 (N_12618,N_2305,N_8514);
and U12619 (N_12619,N_7577,N_4958);
xor U12620 (N_12620,N_7279,N_9087);
and U12621 (N_12621,N_1785,N_4314);
and U12622 (N_12622,N_2117,N_4535);
and U12623 (N_12623,N_4889,N_7612);
and U12624 (N_12624,N_3318,N_6566);
and U12625 (N_12625,N_2406,N_2367);
and U12626 (N_12626,N_9485,N_29);
nand U12627 (N_12627,N_6709,N_1063);
and U12628 (N_12628,N_8991,N_5728);
nand U12629 (N_12629,N_5631,N_4090);
and U12630 (N_12630,N_4309,N_3096);
nor U12631 (N_12631,N_9544,N_9342);
xor U12632 (N_12632,N_8143,N_9224);
and U12633 (N_12633,N_2579,N_6943);
or U12634 (N_12634,N_3660,N_1754);
nor U12635 (N_12635,N_3622,N_414);
and U12636 (N_12636,N_6908,N_3390);
and U12637 (N_12637,N_4,N_2910);
nor U12638 (N_12638,N_5883,N_3254);
xor U12639 (N_12639,N_3124,N_6125);
nand U12640 (N_12640,N_9162,N_2231);
nand U12641 (N_12641,N_3740,N_4674);
or U12642 (N_12642,N_1565,N_6166);
nand U12643 (N_12643,N_2842,N_316);
and U12644 (N_12644,N_432,N_1545);
and U12645 (N_12645,N_8048,N_6443);
xnor U12646 (N_12646,N_8270,N_7496);
nand U12647 (N_12647,N_6468,N_5618);
nand U12648 (N_12648,N_9567,N_8840);
nor U12649 (N_12649,N_2666,N_9698);
nor U12650 (N_12650,N_563,N_2039);
nand U12651 (N_12651,N_8276,N_5456);
or U12652 (N_12652,N_3109,N_136);
or U12653 (N_12653,N_2749,N_4646);
or U12654 (N_12654,N_9417,N_8353);
or U12655 (N_12655,N_317,N_2063);
nor U12656 (N_12656,N_8326,N_147);
and U12657 (N_12657,N_7208,N_6606);
and U12658 (N_12658,N_4941,N_9482);
nand U12659 (N_12659,N_484,N_3466);
nand U12660 (N_12660,N_5599,N_8855);
nor U12661 (N_12661,N_2460,N_6020);
nand U12662 (N_12662,N_8522,N_8934);
or U12663 (N_12663,N_1095,N_1671);
and U12664 (N_12664,N_2946,N_5117);
or U12665 (N_12665,N_5993,N_4027);
and U12666 (N_12666,N_2110,N_2828);
xor U12667 (N_12667,N_1822,N_1007);
and U12668 (N_12668,N_9399,N_6797);
or U12669 (N_12669,N_6184,N_8000);
xor U12670 (N_12670,N_5148,N_3412);
nor U12671 (N_12671,N_8158,N_2075);
and U12672 (N_12672,N_7880,N_2980);
nor U12673 (N_12673,N_3231,N_8116);
nand U12674 (N_12674,N_6795,N_3113);
and U12675 (N_12675,N_3461,N_7107);
or U12676 (N_12676,N_8496,N_8042);
nor U12677 (N_12677,N_3474,N_2890);
xnor U12678 (N_12678,N_9628,N_3306);
nand U12679 (N_12679,N_5813,N_5478);
nor U12680 (N_12680,N_4059,N_1051);
or U12681 (N_12681,N_2284,N_1475);
and U12682 (N_12682,N_4565,N_5889);
nor U12683 (N_12683,N_8628,N_611);
and U12684 (N_12684,N_1919,N_1724);
xnor U12685 (N_12685,N_1257,N_1688);
nand U12686 (N_12686,N_2263,N_2900);
and U12687 (N_12687,N_56,N_1818);
nor U12688 (N_12688,N_3470,N_315);
nand U12689 (N_12689,N_1668,N_144);
or U12690 (N_12690,N_4193,N_9313);
and U12691 (N_12691,N_3029,N_1720);
nor U12692 (N_12692,N_8597,N_7991);
xor U12693 (N_12693,N_6790,N_1643);
xor U12694 (N_12694,N_1635,N_2218);
nor U12695 (N_12695,N_9842,N_3995);
and U12696 (N_12696,N_1782,N_3951);
xor U12697 (N_12697,N_8250,N_7130);
or U12698 (N_12698,N_9153,N_1703);
and U12699 (N_12699,N_6012,N_7497);
nand U12700 (N_12700,N_2258,N_6498);
nor U12701 (N_12701,N_2137,N_8502);
nor U12702 (N_12702,N_1176,N_6190);
and U12703 (N_12703,N_330,N_6783);
or U12704 (N_12704,N_6968,N_270);
and U12705 (N_12705,N_3251,N_4475);
or U12706 (N_12706,N_1457,N_3291);
xnor U12707 (N_12707,N_9073,N_8634);
and U12708 (N_12708,N_3730,N_2286);
or U12709 (N_12709,N_5123,N_5701);
or U12710 (N_12710,N_3615,N_1221);
nand U12711 (N_12711,N_2484,N_9999);
nor U12712 (N_12712,N_1358,N_4359);
and U12713 (N_12713,N_3433,N_9778);
xnor U12714 (N_12714,N_9120,N_4124);
nand U12715 (N_12715,N_2463,N_2713);
or U12716 (N_12716,N_9641,N_7140);
or U12717 (N_12717,N_7327,N_1864);
xor U12718 (N_12718,N_8444,N_1487);
xor U12719 (N_12719,N_733,N_651);
xor U12720 (N_12720,N_6262,N_831);
or U12721 (N_12721,N_1721,N_7726);
or U12722 (N_12722,N_6152,N_5164);
nand U12723 (N_12723,N_2451,N_1490);
or U12724 (N_12724,N_8660,N_6458);
xor U12725 (N_12725,N_9654,N_1660);
nor U12726 (N_12726,N_5474,N_8512);
xnor U12727 (N_12727,N_1967,N_8722);
and U12728 (N_12728,N_1288,N_599);
nand U12729 (N_12729,N_7688,N_6591);
nor U12730 (N_12730,N_9825,N_5608);
nor U12731 (N_12731,N_4122,N_4605);
and U12732 (N_12732,N_3699,N_9050);
nor U12733 (N_12733,N_5065,N_9416);
and U12734 (N_12734,N_9152,N_9717);
or U12735 (N_12735,N_9821,N_9471);
or U12736 (N_12736,N_8838,N_9209);
and U12737 (N_12737,N_197,N_3201);
nor U12738 (N_12738,N_5739,N_3108);
or U12739 (N_12739,N_3043,N_9749);
or U12740 (N_12740,N_5838,N_6645);
xor U12741 (N_12741,N_9297,N_991);
nand U12742 (N_12742,N_8729,N_371);
or U12743 (N_12743,N_2647,N_802);
nor U12744 (N_12744,N_5481,N_9255);
and U12745 (N_12745,N_480,N_168);
and U12746 (N_12746,N_9923,N_3791);
nand U12747 (N_12747,N_6480,N_4352);
xnor U12748 (N_12748,N_1053,N_7658);
nor U12749 (N_12749,N_1416,N_1839);
and U12750 (N_12750,N_2694,N_5256);
nand U12751 (N_12751,N_360,N_3555);
nand U12752 (N_12752,N_6106,N_1559);
nand U12753 (N_12753,N_9026,N_8188);
nor U12754 (N_12754,N_8669,N_9802);
xnor U12755 (N_12755,N_6205,N_8362);
nand U12756 (N_12756,N_8592,N_1633);
xnor U12757 (N_12757,N_4146,N_6748);
nand U12758 (N_12758,N_4139,N_6164);
nand U12759 (N_12759,N_3691,N_759);
and U12760 (N_12760,N_4984,N_6918);
xnor U12761 (N_12761,N_6454,N_2227);
nor U12762 (N_12762,N_7211,N_5225);
xor U12763 (N_12763,N_7718,N_8794);
nor U12764 (N_12764,N_3404,N_6483);
xnor U12765 (N_12765,N_9402,N_2891);
nor U12766 (N_12766,N_220,N_6478);
nor U12767 (N_12767,N_1972,N_5438);
xnor U12768 (N_12768,N_6210,N_1855);
xor U12769 (N_12769,N_4129,N_3634);
xor U12770 (N_12770,N_7563,N_1916);
or U12771 (N_12771,N_9197,N_7338);
nand U12772 (N_12772,N_8012,N_8834);
and U12773 (N_12773,N_3860,N_3587);
nor U12774 (N_12774,N_9511,N_6142);
nor U12775 (N_12775,N_3025,N_4970);
nand U12776 (N_12776,N_7728,N_1684);
or U12777 (N_12777,N_8130,N_3752);
and U12778 (N_12778,N_8553,N_2673);
xnor U12779 (N_12779,N_4859,N_6669);
xnor U12780 (N_12780,N_752,N_9539);
nor U12781 (N_12781,N_8558,N_8202);
and U12782 (N_12782,N_4479,N_5455);
nor U12783 (N_12783,N_8287,N_5598);
or U12784 (N_12784,N_1008,N_5933);
xor U12785 (N_12785,N_2992,N_8749);
or U12786 (N_12786,N_4159,N_8557);
and U12787 (N_12787,N_3921,N_4263);
nor U12788 (N_12788,N_8258,N_4771);
xor U12789 (N_12789,N_6377,N_2147);
nand U12790 (N_12790,N_3162,N_730);
or U12791 (N_12791,N_1664,N_2339);
nand U12792 (N_12792,N_1410,N_1741);
nand U12793 (N_12793,N_8347,N_9831);
xnor U12794 (N_12794,N_9899,N_7494);
nand U12795 (N_12795,N_1516,N_7582);
xor U12796 (N_12796,N_9373,N_3596);
nor U12797 (N_12797,N_2606,N_4577);
nand U12798 (N_12798,N_1550,N_104);
and U12799 (N_12799,N_7246,N_6520);
xnor U12800 (N_12800,N_6239,N_8399);
nand U12801 (N_12801,N_6085,N_5276);
and U12802 (N_12802,N_7879,N_5921);
and U12803 (N_12803,N_2417,N_7200);
or U12804 (N_12804,N_7154,N_1662);
nor U12805 (N_12805,N_5322,N_1343);
xor U12806 (N_12806,N_6373,N_7370);
nor U12807 (N_12807,N_5203,N_9056);
nor U12808 (N_12808,N_7351,N_1707);
nand U12809 (N_12809,N_5976,N_8679);
xnor U12810 (N_12810,N_1065,N_3534);
or U12811 (N_12811,N_1178,N_1717);
and U12812 (N_12812,N_4920,N_5019);
and U12813 (N_12813,N_9519,N_655);
nor U12814 (N_12814,N_9195,N_2288);
or U12815 (N_12815,N_8690,N_6569);
xnor U12816 (N_12816,N_5865,N_9787);
xnor U12817 (N_12817,N_4557,N_4298);
and U12818 (N_12818,N_1982,N_5294);
and U12819 (N_12819,N_486,N_9935);
nor U12820 (N_12820,N_1333,N_742);
xor U12821 (N_12821,N_7939,N_8903);
or U12822 (N_12822,N_5955,N_4140);
and U12823 (N_12823,N_4478,N_9470);
nor U12824 (N_12824,N_4891,N_8101);
and U12825 (N_12825,N_71,N_6268);
nand U12826 (N_12826,N_3765,N_799);
xnor U12827 (N_12827,N_2657,N_6135);
xnor U12828 (N_12828,N_5957,N_1250);
xnor U12829 (N_12829,N_1582,N_9124);
and U12830 (N_12830,N_7283,N_2791);
xnor U12831 (N_12831,N_3932,N_2196);
nor U12832 (N_12832,N_883,N_636);
nor U12833 (N_12833,N_8072,N_418);
nand U12834 (N_12834,N_3782,N_3985);
and U12835 (N_12835,N_6025,N_7659);
and U12836 (N_12836,N_5719,N_7923);
nand U12837 (N_12837,N_3422,N_7715);
and U12838 (N_12838,N_4412,N_8162);
and U12839 (N_12839,N_6613,N_146);
or U12840 (N_12840,N_2533,N_2107);
and U12841 (N_12841,N_335,N_193);
nor U12842 (N_12842,N_3701,N_682);
and U12843 (N_12843,N_8153,N_917);
xnor U12844 (N_12844,N_2881,N_1940);
or U12845 (N_12845,N_9273,N_2827);
xor U12846 (N_12846,N_1339,N_3923);
or U12847 (N_12847,N_9100,N_9165);
or U12848 (N_12848,N_4397,N_9431);
and U12849 (N_12849,N_8411,N_7965);
nor U12850 (N_12850,N_1896,N_6555);
and U12851 (N_12851,N_5284,N_2807);
or U12852 (N_12852,N_2804,N_7485);
xnor U12853 (N_12853,N_267,N_4228);
or U12854 (N_12854,N_1572,N_6193);
nor U12855 (N_12855,N_287,N_3440);
xnor U12856 (N_12856,N_9003,N_5434);
and U12857 (N_12857,N_6325,N_5551);
xnor U12858 (N_12858,N_9295,N_1737);
and U12859 (N_12859,N_3432,N_5341);
nor U12860 (N_12860,N_5252,N_1820);
xor U12861 (N_12861,N_2241,N_4276);
and U12862 (N_12862,N_2964,N_6562);
nand U12863 (N_12863,N_9139,N_3836);
nand U12864 (N_12864,N_8470,N_3078);
xnor U12865 (N_12865,N_8349,N_6574);
nand U12866 (N_12866,N_9052,N_9381);
nor U12867 (N_12867,N_4060,N_2431);
xor U12868 (N_12868,N_7710,N_552);
or U12869 (N_12869,N_3604,N_6212);
and U12870 (N_12870,N_6428,N_1365);
or U12871 (N_12871,N_7966,N_2320);
or U12872 (N_12872,N_5131,N_3984);
and U12873 (N_12873,N_5509,N_9690);
nor U12874 (N_12874,N_8662,N_6965);
xor U12875 (N_12875,N_9341,N_3769);
or U12876 (N_12876,N_9108,N_443);
nor U12877 (N_12877,N_4350,N_9956);
or U12878 (N_12878,N_5586,N_5978);
nand U12879 (N_12879,N_8963,N_3485);
and U12880 (N_12880,N_2497,N_8940);
nand U12881 (N_12881,N_452,N_9755);
nand U12882 (N_12882,N_2269,N_394);
xor U12883 (N_12883,N_6309,N_4794);
or U12884 (N_12884,N_5846,N_8760);
or U12885 (N_12885,N_4476,N_2981);
xnor U12886 (N_12886,N_3657,N_9418);
or U12887 (N_12887,N_4258,N_2703);
nand U12888 (N_12888,N_4885,N_2158);
or U12889 (N_12889,N_9444,N_2885);
nor U12890 (N_12890,N_3538,N_5451);
nor U12891 (N_12891,N_3721,N_2726);
nor U12892 (N_12892,N_5051,N_4654);
and U12893 (N_12893,N_1537,N_932);
xnor U12894 (N_12894,N_9833,N_4719);
or U12895 (N_12895,N_3006,N_8879);
nor U12896 (N_12896,N_6550,N_6482);
and U12897 (N_12897,N_8037,N_3665);
nor U12898 (N_12898,N_6656,N_3828);
xor U12899 (N_12899,N_7886,N_9347);
nand U12900 (N_12900,N_1236,N_784);
xor U12901 (N_12901,N_3718,N_9024);
or U12902 (N_12902,N_4011,N_1011);
xnor U12903 (N_12903,N_2485,N_7044);
nor U12904 (N_12904,N_7721,N_9011);
xor U12905 (N_12905,N_8337,N_1380);
xnor U12906 (N_12906,N_3610,N_3114);
and U12907 (N_12907,N_1728,N_5163);
or U12908 (N_12908,N_5854,N_5873);
nor U12909 (N_12909,N_5013,N_8815);
or U12910 (N_12910,N_9430,N_6980);
and U12911 (N_12911,N_5652,N_1272);
and U12912 (N_12912,N_6534,N_8115);
nand U12913 (N_12913,N_8653,N_3890);
and U12914 (N_12914,N_7850,N_1259);
nand U12915 (N_12915,N_9508,N_704);
nand U12916 (N_12916,N_2505,N_4000);
nor U12917 (N_12917,N_8674,N_4097);
or U12918 (N_12918,N_8065,N_6640);
and U12919 (N_12919,N_3883,N_9092);
and U12920 (N_12920,N_9810,N_1143);
xnor U12921 (N_12921,N_1949,N_1498);
xor U12922 (N_12922,N_7427,N_4283);
nor U12923 (N_12923,N_1608,N_2861);
or U12924 (N_12924,N_6337,N_3878);
and U12925 (N_12925,N_338,N_4855);
nand U12926 (N_12926,N_9156,N_7343);
nor U12927 (N_12927,N_4568,N_9375);
or U12928 (N_12928,N_717,N_6401);
nand U12929 (N_12929,N_919,N_2138);
nand U12930 (N_12930,N_2732,N_5467);
nand U12931 (N_12931,N_3147,N_5368);
or U12932 (N_12932,N_1687,N_4656);
nand U12933 (N_12933,N_2956,N_8839);
nand U12934 (N_12934,N_6522,N_5707);
xnor U12935 (N_12935,N_2784,N_6988);
nor U12936 (N_12936,N_6740,N_7257);
or U12937 (N_12937,N_1843,N_1076);
xor U12938 (N_12938,N_6876,N_1287);
or U12939 (N_12939,N_3125,N_9710);
and U12940 (N_12940,N_5407,N_2199);
nor U12941 (N_12941,N_7346,N_2042);
and U12942 (N_12942,N_2341,N_2046);
nand U12943 (N_12943,N_1665,N_2627);
nor U12944 (N_12944,N_1071,N_1389);
or U12945 (N_12945,N_3746,N_2081);
nand U12946 (N_12946,N_7742,N_3521);
xnor U12947 (N_12947,N_4071,N_8160);
nor U12948 (N_12948,N_6754,N_3957);
nor U12949 (N_12949,N_595,N_974);
xor U12950 (N_12950,N_1201,N_9489);
nor U12951 (N_12951,N_7962,N_8291);
or U12952 (N_12952,N_7834,N_2639);
or U12953 (N_12953,N_5756,N_2944);
xnor U12954 (N_12954,N_2000,N_2324);
and U12955 (N_12955,N_647,N_80);
and U12956 (N_12956,N_2334,N_681);
nor U12957 (N_12957,N_2091,N_6778);
nand U12958 (N_12958,N_4579,N_7527);
xor U12959 (N_12959,N_253,N_6637);
or U12960 (N_12960,N_7703,N_580);
xor U12961 (N_12961,N_6078,N_6531);
or U12962 (N_12962,N_7753,N_3366);
nor U12963 (N_12963,N_8965,N_4544);
or U12964 (N_12964,N_5196,N_3571);
or U12965 (N_12965,N_3052,N_198);
xnor U12966 (N_12966,N_7771,N_3481);
nand U12967 (N_12967,N_1415,N_2121);
nand U12968 (N_12968,N_1540,N_4572);
xnor U12969 (N_12969,N_7499,N_6196);
or U12970 (N_12970,N_281,N_6878);
or U12971 (N_12971,N_6729,N_3055);
xnor U12972 (N_12972,N_7300,N_4221);
nor U12973 (N_12973,N_5709,N_952);
nand U12974 (N_12974,N_6060,N_6799);
and U12975 (N_12975,N_1035,N_4103);
nor U12976 (N_12976,N_170,N_2495);
nor U12977 (N_12977,N_2923,N_3637);
nand U12978 (N_12978,N_3370,N_5367);
xnor U12979 (N_12979,N_4175,N_5980);
xnor U12980 (N_12980,N_2025,N_2854);
nor U12981 (N_12981,N_9980,N_5503);
xor U12982 (N_12982,N_1453,N_4867);
nor U12983 (N_12983,N_8482,N_5040);
and U12984 (N_12984,N_9265,N_7824);
and U12985 (N_12985,N_8403,N_1685);
xor U12986 (N_12986,N_1519,N_847);
nand U12987 (N_12987,N_4556,N_8763);
nor U12988 (N_12988,N_3170,N_1702);
nor U12989 (N_12989,N_4100,N_8288);
xor U12990 (N_12990,N_7388,N_4486);
nand U12991 (N_12991,N_4236,N_1121);
and U12992 (N_12992,N_4480,N_8617);
xor U12993 (N_12993,N_5587,N_298);
and U12994 (N_12994,N_2099,N_6259);
or U12995 (N_12995,N_3846,N_4587);
or U12996 (N_12996,N_1434,N_3092);
xor U12997 (N_12997,N_807,N_6766);
nor U12998 (N_12998,N_2290,N_7292);
nand U12999 (N_12999,N_4645,N_6375);
xor U13000 (N_13000,N_7159,N_132);
or U13001 (N_13001,N_4586,N_8637);
xor U13002 (N_13002,N_3337,N_4281);
nand U13003 (N_13003,N_1933,N_2119);
and U13004 (N_13004,N_4907,N_7176);
or U13005 (N_13005,N_7579,N_7569);
and U13006 (N_13006,N_4811,N_1408);
and U13007 (N_13007,N_3515,N_6822);
or U13008 (N_13008,N_4081,N_7559);
or U13009 (N_13009,N_8604,N_9955);
xnor U13010 (N_13010,N_6710,N_6793);
nand U13011 (N_13011,N_1748,N_1557);
xor U13012 (N_13012,N_5862,N_3916);
nor U13013 (N_13013,N_6120,N_1105);
and U13014 (N_13014,N_492,N_2228);
and U13015 (N_13015,N_9797,N_5997);
or U13016 (N_13016,N_3561,N_6476);
xnor U13017 (N_13017,N_6960,N_1048);
or U13018 (N_13018,N_6092,N_5684);
or U13019 (N_13019,N_349,N_2123);
nor U13020 (N_13020,N_1460,N_331);
xnor U13021 (N_13021,N_9386,N_8951);
or U13022 (N_13022,N_1598,N_2959);
and U13023 (N_13023,N_9490,N_8867);
nand U13024 (N_13024,N_1279,N_6938);
xor U13025 (N_13025,N_4541,N_2684);
nor U13026 (N_13026,N_3097,N_174);
nand U13027 (N_13027,N_9534,N_8285);
or U13028 (N_13028,N_2517,N_2089);
or U13029 (N_13029,N_9887,N_7223);
or U13030 (N_13030,N_7518,N_5935);
xor U13031 (N_13031,N_3934,N_949);
nand U13032 (N_13032,N_2374,N_7894);
nor U13033 (N_13033,N_3550,N_1359);
nor U13034 (N_13034,N_4753,N_4729);
and U13035 (N_13035,N_7293,N_356);
and U13036 (N_13036,N_7280,N_6017);
nand U13037 (N_13037,N_2810,N_4426);
xnor U13038 (N_13038,N_9929,N_5938);
or U13039 (N_13039,N_28,N_4286);
xor U13040 (N_13040,N_1278,N_6666);
xnor U13041 (N_13041,N_7903,N_7319);
or U13042 (N_13042,N_4061,N_6851);
nor U13043 (N_13043,N_2960,N_6283);
and U13044 (N_13044,N_650,N_5533);
and U13045 (N_13045,N_2222,N_1485);
and U13046 (N_13046,N_3737,N_4482);
or U13047 (N_13047,N_5085,N_7543);
or U13048 (N_13048,N_6931,N_7324);
or U13049 (N_13049,N_9610,N_4135);
nor U13050 (N_13050,N_4294,N_8207);
nor U13051 (N_13051,N_1072,N_9823);
nor U13052 (N_13052,N_5373,N_7564);
and U13053 (N_13053,N_7055,N_7120);
nor U13054 (N_13054,N_357,N_7100);
and U13055 (N_13055,N_6187,N_7190);
and U13056 (N_13056,N_4181,N_402);
nand U13057 (N_13057,N_2940,N_653);
nand U13058 (N_13058,N_5640,N_5722);
or U13059 (N_13059,N_2935,N_4077);
xnor U13060 (N_13060,N_890,N_1370);
or U13061 (N_13061,N_1794,N_3392);
and U13062 (N_13062,N_8692,N_2751);
xnor U13063 (N_13063,N_8290,N_3371);
xnor U13064 (N_13064,N_817,N_9022);
and U13065 (N_13065,N_2181,N_6809);
and U13066 (N_13066,N_5482,N_8025);
nor U13067 (N_13067,N_5133,N_8526);
and U13068 (N_13068,N_5088,N_9656);
nor U13069 (N_13069,N_2159,N_6021);
nor U13070 (N_13070,N_7282,N_975);
and U13071 (N_13071,N_4239,N_5374);
xor U13072 (N_13072,N_4065,N_5119);
nor U13073 (N_13073,N_375,N_8809);
nand U13074 (N_13074,N_9918,N_4932);
and U13075 (N_13075,N_6090,N_8945);
and U13076 (N_13076,N_2976,N_7804);
xor U13077 (N_13077,N_2481,N_1096);
and U13078 (N_13078,N_5925,N_4880);
and U13079 (N_13079,N_586,N_9332);
nor U13080 (N_13080,N_7931,N_5610);
xnor U13081 (N_13081,N_3299,N_3528);
and U13082 (N_13082,N_1941,N_6880);
xnor U13083 (N_13083,N_2392,N_9530);
or U13084 (N_13084,N_4722,N_4151);
and U13085 (N_13085,N_8892,N_1256);
nor U13086 (N_13086,N_1798,N_9894);
and U13087 (N_13087,N_5179,N_9933);
nor U13088 (N_13088,N_3424,N_8122);
or U13089 (N_13089,N_7542,N_3480);
xnor U13090 (N_13090,N_8707,N_9075);
and U13091 (N_13091,N_1534,N_4435);
nand U13092 (N_13092,N_7738,N_3446);
nor U13093 (N_13093,N_3834,N_8835);
and U13094 (N_13094,N_8173,N_6577);
or U13095 (N_13095,N_4176,N_5411);
or U13096 (N_13096,N_8208,N_1868);
nand U13097 (N_13097,N_3874,N_2985);
xor U13098 (N_13098,N_2954,N_6838);
nand U13099 (N_13099,N_838,N_3996);
and U13100 (N_13100,N_205,N_4008);
or U13101 (N_13101,N_1428,N_9184);
and U13102 (N_13102,N_5964,N_4417);
nor U13103 (N_13103,N_445,N_602);
nand U13104 (N_13104,N_9579,N_4803);
or U13105 (N_13105,N_3391,N_13);
and U13106 (N_13106,N_921,N_2525);
nand U13107 (N_13107,N_6234,N_463);
nor U13108 (N_13108,N_3095,N_3028);
xor U13109 (N_13109,N_2166,N_1732);
or U13110 (N_13110,N_1561,N_1510);
nand U13111 (N_13111,N_840,N_1939);
and U13112 (N_13112,N_8355,N_295);
xnor U13113 (N_13113,N_3651,N_4291);
and U13114 (N_13114,N_3202,N_5995);
xor U13115 (N_13115,N_4019,N_7173);
nand U13116 (N_13116,N_7704,N_3959);
and U13117 (N_13117,N_4271,N_7558);
xnor U13118 (N_13118,N_4936,N_4955);
nand U13119 (N_13119,N_2670,N_4403);
and U13120 (N_13120,N_4622,N_378);
xnor U13121 (N_13121,N_9898,N_3070);
or U13122 (N_13122,N_9541,N_9517);
nand U13123 (N_13123,N_8671,N_1502);
xnor U13124 (N_13124,N_3315,N_1368);
nand U13125 (N_13125,N_7337,N_5898);
xor U13126 (N_13126,N_9593,N_5457);
and U13127 (N_13127,N_9893,N_5318);
nand U13128 (N_13128,N_2806,N_1596);
or U13129 (N_13129,N_8068,N_7174);
or U13130 (N_13130,N_6172,N_4538);
nand U13131 (N_13131,N_4232,N_5037);
nor U13132 (N_13132,N_2237,N_6849);
xnor U13133 (N_13133,N_8343,N_7508);
nor U13134 (N_13134,N_4551,N_4233);
nand U13135 (N_13135,N_5253,N_9266);
or U13136 (N_13136,N_9246,N_1993);
nor U13137 (N_13137,N_4091,N_4042);
and U13138 (N_13138,N_5884,N_2097);
xor U13139 (N_13139,N_2351,N_8322);
xnor U13140 (N_13140,N_5268,N_8710);
and U13141 (N_13141,N_7795,N_8717);
or U13142 (N_13142,N_133,N_9590);
or U13143 (N_13143,N_943,N_405);
nor U13144 (N_13144,N_5382,N_4942);
and U13145 (N_13145,N_9822,N_7633);
nand U13146 (N_13146,N_8646,N_3235);
nand U13147 (N_13147,N_7421,N_6773);
nand U13148 (N_13148,N_7673,N_2285);
or U13149 (N_13149,N_3686,N_1325);
nand U13150 (N_13150,N_1678,N_1845);
and U13151 (N_13151,N_4721,N_4739);
nand U13152 (N_13152,N_47,N_569);
xnor U13153 (N_13153,N_8811,N_7077);
and U13154 (N_13154,N_3912,N_9114);
or U13155 (N_13155,N_6084,N_7698);
nor U13156 (N_13156,N_4493,N_5486);
nor U13157 (N_13157,N_5254,N_4692);
nor U13158 (N_13158,N_4959,N_7026);
or U13159 (N_13159,N_5011,N_5777);
and U13160 (N_13160,N_1862,N_1039);
nor U13161 (N_13161,N_8694,N_473);
or U13162 (N_13162,N_1604,N_7812);
nor U13163 (N_13163,N_2802,N_8021);
and U13164 (N_13164,N_4498,N_8121);
and U13165 (N_13165,N_6802,N_7213);
nand U13166 (N_13166,N_2668,N_4138);
nor U13167 (N_13167,N_7955,N_1320);
nor U13168 (N_13168,N_6495,N_8246);
nor U13169 (N_13169,N_3855,N_9668);
nor U13170 (N_13170,N_8472,N_3839);
xnor U13171 (N_13171,N_3633,N_6828);
nand U13172 (N_13172,N_3115,N_3918);
nand U13173 (N_13173,N_11,N_2483);
nand U13174 (N_13174,N_4067,N_5695);
xnor U13175 (N_13175,N_7456,N_2112);
and U13176 (N_13176,N_5797,N_6039);
nand U13177 (N_13177,N_7483,N_7268);
and U13178 (N_13178,N_4785,N_6910);
and U13179 (N_13179,N_3473,N_9997);
nand U13180 (N_13180,N_8146,N_7741);
or U13181 (N_13181,N_9696,N_7091);
and U13182 (N_13182,N_6133,N_8474);
or U13183 (N_13183,N_5910,N_7271);
nor U13184 (N_13184,N_3209,N_2390);
or U13185 (N_13185,N_8929,N_1045);
nand U13186 (N_13186,N_871,N_4637);
or U13187 (N_13187,N_9667,N_6845);
nor U13188 (N_13188,N_4901,N_5623);
and U13189 (N_13189,N_5462,N_5049);
and U13190 (N_13190,N_9934,N_5674);
or U13191 (N_13191,N_6461,N_9896);
xor U13192 (N_13192,N_39,N_1003);
and U13193 (N_13193,N_3826,N_6592);
nand U13194 (N_13194,N_605,N_6352);
or U13195 (N_13195,N_156,N_3659);
nor U13196 (N_13196,N_7848,N_4361);
xor U13197 (N_13197,N_5834,N_9016);
and U13198 (N_13198,N_6091,N_4038);
nand U13199 (N_13199,N_6889,N_7053);
xnor U13200 (N_13200,N_4452,N_5878);
nor U13201 (N_13201,N_6985,N_53);
nor U13202 (N_13202,N_4755,N_509);
nand U13203 (N_13203,N_7858,N_9168);
nand U13204 (N_13204,N_4823,N_9408);
xor U13205 (N_13205,N_5408,N_7817);
nor U13206 (N_13206,N_7081,N_4419);
nor U13207 (N_13207,N_7793,N_6840);
nand U13208 (N_13208,N_5170,N_2168);
or U13209 (N_13209,N_1881,N_494);
or U13210 (N_13210,N_9644,N_4752);
or U13211 (N_13211,N_5025,N_3994);
nor U13212 (N_13212,N_6426,N_8108);
or U13213 (N_13213,N_1125,N_3172);
or U13214 (N_13214,N_4619,N_7158);
or U13215 (N_13215,N_2058,N_2918);
xor U13216 (N_13216,N_5427,N_2844);
or U13217 (N_13217,N_4491,N_1019);
or U13218 (N_13218,N_1493,N_1205);
and U13219 (N_13219,N_7822,N_3568);
or U13220 (N_13220,N_2372,N_987);
xor U13221 (N_13221,N_9868,N_9307);
nor U13222 (N_13222,N_5676,N_6089);
xnor U13223 (N_13223,N_9550,N_3598);
or U13224 (N_13224,N_8092,N_9974);
xor U13225 (N_13225,N_9513,N_7696);
nor U13226 (N_13226,N_3969,N_2387);
or U13227 (N_13227,N_4957,N_9925);
or U13228 (N_13228,N_5532,N_3574);
nand U13229 (N_13229,N_3966,N_2409);
nor U13230 (N_13230,N_2363,N_9406);
xnor U13231 (N_13231,N_1813,N_8756);
and U13232 (N_13232,N_97,N_1840);
or U13233 (N_13233,N_2884,N_4337);
nor U13234 (N_13234,N_633,N_3407);
nand U13235 (N_13235,N_5141,N_2368);
and U13236 (N_13236,N_6395,N_9460);
nand U13237 (N_13237,N_9559,N_75);
or U13238 (N_13238,N_2010,N_4757);
xnor U13239 (N_13239,N_8769,N_151);
nand U13240 (N_13240,N_5391,N_4712);
xor U13241 (N_13241,N_1619,N_541);
xor U13242 (N_13242,N_3744,N_5595);
or U13243 (N_13243,N_4664,N_5332);
nor U13244 (N_13244,N_4341,N_5926);
nand U13245 (N_13245,N_9815,N_8883);
and U13246 (N_13246,N_6747,N_9044);
or U13247 (N_13247,N_6835,N_603);
nand U13248 (N_13248,N_748,N_816);
or U13249 (N_13249,N_4979,N_1807);
nor U13250 (N_13250,N_7922,N_1505);
nor U13251 (N_13251,N_8899,N_9432);
nand U13252 (N_13252,N_5521,N_5443);
nand U13253 (N_13253,N_2722,N_9215);
nand U13254 (N_13254,N_6197,N_3244);
or U13255 (N_13255,N_8247,N_8630);
xnor U13256 (N_13256,N_41,N_3917);
and U13257 (N_13257,N_500,N_4402);
or U13258 (N_13258,N_1341,N_1395);
and U13259 (N_13259,N_9125,N_3570);
xnor U13260 (N_13260,N_5245,N_4760);
and U13261 (N_13261,N_589,N_9001);
and U13262 (N_13262,N_2292,N_842);
nor U13263 (N_13263,N_9358,N_3897);
xnor U13264 (N_13264,N_5698,N_8248);
and U13265 (N_13265,N_3663,N_973);
nor U13266 (N_13266,N_3886,N_4731);
and U13267 (N_13267,N_6158,N_59);
or U13268 (N_13268,N_3310,N_3106);
and U13269 (N_13269,N_1164,N_8035);
or U13270 (N_13270,N_3156,N_8088);
or U13271 (N_13271,N_4487,N_3237);
nor U13272 (N_13272,N_1826,N_4658);
xnor U13273 (N_13273,N_8182,N_1884);
or U13274 (N_13274,N_4372,N_8441);
or U13275 (N_13275,N_3904,N_27);
and U13276 (N_13276,N_2650,N_965);
and U13277 (N_13277,N_526,N_4887);
xnor U13278 (N_13278,N_6213,N_6777);
and U13279 (N_13279,N_7819,N_6971);
nor U13280 (N_13280,N_1512,N_7187);
nor U13281 (N_13281,N_262,N_804);
or U13282 (N_13282,N_3178,N_9176);
or U13283 (N_13283,N_888,N_8806);
or U13284 (N_13284,N_5362,N_849);
or U13285 (N_13285,N_1291,N_7170);
and U13286 (N_13286,N_1295,N_3425);
or U13287 (N_13287,N_7316,N_5786);
and U13288 (N_13288,N_670,N_3469);
nand U13289 (N_13289,N_9770,N_7359);
nor U13290 (N_13290,N_1503,N_6626);
or U13291 (N_13291,N_9032,N_1200);
and U13292 (N_13292,N_2831,N_3862);
nor U13293 (N_13293,N_9260,N_654);
or U13294 (N_13294,N_4026,N_4648);
nand U13295 (N_13295,N_2537,N_5012);
xor U13296 (N_13296,N_1446,N_1800);
nand U13297 (N_13297,N_4897,N_6409);
nor U13298 (N_13298,N_1600,N_1276);
nor U13299 (N_13299,N_8923,N_268);
nand U13300 (N_13300,N_1690,N_1417);
and U13301 (N_13301,N_7493,N_1391);
or U13302 (N_13302,N_6912,N_3776);
nor U13303 (N_13303,N_4152,N_887);
xor U13304 (N_13304,N_6953,N_753);
xnor U13305 (N_13305,N_3058,N_6225);
nor U13306 (N_13306,N_2165,N_8328);
or U13307 (N_13307,N_3710,N_3024);
or U13308 (N_13308,N_6859,N_5162);
nand U13309 (N_13309,N_7227,N_4806);
nand U13310 (N_13310,N_5128,N_1712);
xnor U13311 (N_13311,N_7580,N_341);
nor U13312 (N_13312,N_9099,N_5046);
xnor U13313 (N_13313,N_2397,N_3083);
or U13314 (N_13314,N_9378,N_4157);
xnor U13315 (N_13315,N_832,N_8857);
nand U13316 (N_13316,N_4937,N_9464);
and U13317 (N_13317,N_2561,N_2212);
and U13318 (N_13318,N_37,N_6580);
nand U13319 (N_13319,N_364,N_4536);
and U13320 (N_13320,N_3531,N_6323);
xor U13321 (N_13321,N_9362,N_2283);
or U13322 (N_13322,N_1420,N_3479);
or U13323 (N_13323,N_6137,N_6415);
xor U13324 (N_13324,N_3010,N_5027);
or U13325 (N_13325,N_8972,N_2597);
or U13326 (N_13326,N_3222,N_6744);
nand U13327 (N_13327,N_4484,N_7970);
or U13328 (N_13328,N_1223,N_6270);
nand U13329 (N_13329,N_2758,N_562);
nand U13330 (N_13330,N_4222,N_1435);
and U13331 (N_13331,N_2675,N_9309);
and U13332 (N_13332,N_6346,N_3393);
nor U13333 (N_13333,N_4266,N_6684);
xnor U13334 (N_13334,N_3133,N_9442);
nor U13335 (N_13335,N_1905,N_556);
and U13336 (N_13336,N_2697,N_923);
nor U13337 (N_13337,N_6111,N_7067);
xnor U13338 (N_13338,N_487,N_8106);
nor U13339 (N_13339,N_8152,N_2146);
xor U13340 (N_13340,N_1926,N_1418);
nor U13341 (N_13341,N_4509,N_2908);
and U13342 (N_13342,N_1316,N_9777);
or U13343 (N_13343,N_5712,N_6649);
nor U13344 (N_13344,N_413,N_5272);
nand U13345 (N_13345,N_8691,N_829);
or U13346 (N_13346,N_8598,N_7798);
nor U13347 (N_13347,N_7764,N_7471);
nand U13348 (N_13348,N_4590,N_2933);
or U13349 (N_13349,N_8946,N_5495);
xor U13350 (N_13350,N_148,N_6479);
xnor U13351 (N_13351,N_5653,N_609);
nor U13352 (N_13352,N_5697,N_3565);
nand U13353 (N_13353,N_7565,N_4471);
or U13354 (N_13354,N_9943,N_3901);
and U13355 (N_13355,N_2435,N_7839);
and U13356 (N_13356,N_3080,N_7467);
and U13357 (N_13357,N_2592,N_6850);
or U13358 (N_13358,N_1120,N_6322);
nor U13359 (N_13359,N_8765,N_9872);
nor U13360 (N_13360,N_6623,N_2095);
and U13361 (N_13361,N_5550,N_3786);
and U13362 (N_13362,N_4540,N_5007);
nand U13363 (N_13363,N_3060,N_1548);
nand U13364 (N_13364,N_7463,N_7607);
and U13365 (N_13365,N_6329,N_4223);
and U13366 (N_13366,N_663,N_7498);
nor U13367 (N_13367,N_9351,N_4829);
xor U13368 (N_13368,N_8998,N_6611);
or U13369 (N_13369,N_5337,N_5518);
nor U13370 (N_13370,N_9372,N_1252);
nor U13371 (N_13371,N_3569,N_5715);
nand U13372 (N_13372,N_1298,N_1113);
nand U13373 (N_13373,N_7756,N_6674);
and U13374 (N_13374,N_8501,N_2303);
or U13375 (N_13375,N_7038,N_6667);
nor U13376 (N_13376,N_1456,N_7241);
nand U13377 (N_13377,N_9161,N_2521);
nor U13378 (N_13378,N_8971,N_8816);
xnor U13379 (N_13379,N_24,N_9665);
nor U13380 (N_13380,N_2185,N_645);
and U13381 (N_13381,N_9199,N_2465);
and U13382 (N_13382,N_7531,N_2680);
and U13383 (N_13383,N_7048,N_4754);
nand U13384 (N_13384,N_9998,N_6183);
or U13385 (N_13385,N_6339,N_4564);
xnor U13386 (N_13386,N_7172,N_7730);
nor U13387 (N_13387,N_5464,N_5575);
nand U13388 (N_13388,N_2729,N_2839);
and U13389 (N_13389,N_6625,N_8392);
nor U13390 (N_13390,N_2692,N_4210);
xnor U13391 (N_13391,N_4981,N_6011);
nor U13392 (N_13392,N_9223,N_2528);
nor U13393 (N_13393,N_5436,N_283);
xnor U13394 (N_13394,N_893,N_8509);
xnor U13395 (N_13395,N_6844,N_5850);
nor U13396 (N_13396,N_5860,N_715);
and U13397 (N_13397,N_4627,N_8365);
or U13398 (N_13398,N_848,N_662);
nand U13399 (N_13399,N_4818,N_2572);
nand U13400 (N_13400,N_8457,N_2449);
nor U13401 (N_13401,N_9941,N_2924);
nor U13402 (N_13402,N_7382,N_8233);
nand U13403 (N_13403,N_1102,N_1530);
nand U13404 (N_13404,N_2067,N_4164);
nand U13405 (N_13405,N_5678,N_3305);
and U13406 (N_13406,N_6998,N_2235);
or U13407 (N_13407,N_867,N_3387);
and U13408 (N_13408,N_6390,N_6004);
and U13409 (N_13409,N_9186,N_2252);
xnor U13410 (N_13410,N_8599,N_1356);
nor U13411 (N_13411,N_3830,N_9425);
xor U13412 (N_13412,N_8603,N_8003);
or U13413 (N_13413,N_549,N_4204);
or U13414 (N_13414,N_3889,N_7302);
xnor U13415 (N_13415,N_2988,N_4782);
nor U13416 (N_13416,N_3281,N_8718);
nand U13417 (N_13417,N_2695,N_3105);
xnor U13418 (N_13418,N_8982,N_5657);
or U13419 (N_13419,N_4844,N_9507);
or U13420 (N_13420,N_9585,N_2629);
xor U13421 (N_13421,N_7836,N_3104);
and U13422 (N_13422,N_8332,N_8084);
nor U13423 (N_13423,N_1989,N_7891);
and U13424 (N_13424,N_9208,N_6316);
or U13425 (N_13425,N_403,N_1353);
xnor U13426 (N_13426,N_3438,N_5313);
and U13427 (N_13427,N_2220,N_2182);
nor U13428 (N_13428,N_471,N_2614);
nand U13429 (N_13429,N_4477,N_276);
or U13430 (N_13430,N_7861,N_3683);
and U13431 (N_13431,N_4053,N_2096);
and U13432 (N_13432,N_5070,N_2602);
or U13433 (N_13433,N_7060,N_5072);
or U13434 (N_13434,N_6156,N_2587);
xor U13435 (N_13435,N_7003,N_5968);
nor U13436 (N_13436,N_2127,N_2225);
nand U13437 (N_13437,N_4960,N_3293);
nor U13438 (N_13438,N_9183,N_9207);
or U13439 (N_13439,N_1714,N_3355);
nor U13440 (N_13440,N_1531,N_1701);
xor U13441 (N_13441,N_2302,N_6473);
xnor U13442 (N_13442,N_3592,N_421);
and U13443 (N_13443,N_6180,N_3891);
and U13444 (N_13444,N_743,N_7080);
xor U13445 (N_13445,N_3882,N_2213);
nor U13446 (N_13446,N_82,N_8751);
nor U13447 (N_13447,N_6515,N_3668);
xnor U13448 (N_13448,N_5309,N_9333);
nand U13449 (N_13449,N_5,N_8814);
nor U13450 (N_13450,N_21,N_6612);
and U13451 (N_13451,N_4854,N_3552);
or U13452 (N_13452,N_4394,N_3177);
nand U13453 (N_13453,N_6487,N_6057);
nand U13454 (N_13454,N_904,N_8031);
and U13455 (N_13455,N_1667,N_3965);
or U13456 (N_13456,N_3922,N_3273);
xnor U13457 (N_13457,N_4320,N_779);
xor U13458 (N_13458,N_1406,N_4965);
nand U13459 (N_13459,N_2020,N_510);
or U13460 (N_13460,N_3827,N_9982);
nand U13461 (N_13461,N_9976,N_8477);
and U13462 (N_13462,N_154,N_2421);
or U13463 (N_13463,N_8817,N_3619);
and U13464 (N_13464,N_4502,N_430);
nor U13465 (N_13465,N_1317,N_7716);
or U13466 (N_13466,N_688,N_2312);
and U13467 (N_13467,N_8334,N_8431);
nor U13468 (N_13468,N_2211,N_6578);
nand U13469 (N_13469,N_9948,N_3001);
xnor U13470 (N_13470,N_4838,N_6771);
nand U13471 (N_13471,N_5483,N_9981);
nor U13472 (N_13472,N_8672,N_5475);
xnor U13473 (N_13473,N_2150,N_3126);
nand U13474 (N_13474,N_6609,N_6455);
nor U13475 (N_13475,N_5122,N_4242);
xor U13476 (N_13476,N_4057,N_1936);
or U13477 (N_13477,N_3785,N_8361);
or U13478 (N_13478,N_8684,N_9059);
or U13479 (N_13479,N_1384,N_1228);
nor U13480 (N_13480,N_1155,N_3159);
or U13481 (N_13481,N_8933,N_5029);
nor U13482 (N_13482,N_43,N_9551);
or U13483 (N_13483,N_1647,N_310);
or U13484 (N_13484,N_5939,N_3487);
or U13485 (N_13485,N_766,N_8715);
or U13486 (N_13486,N_4413,N_8956);
or U13487 (N_13487,N_2053,N_9647);
or U13488 (N_13488,N_9675,N_3389);
nor U13489 (N_13489,N_6047,N_5794);
nor U13490 (N_13490,N_2907,N_7290);
nand U13491 (N_13491,N_439,N_3748);
and U13492 (N_13492,N_4578,N_5798);
or U13493 (N_13493,N_714,N_2143);
and U13494 (N_13494,N_8790,N_5842);
xnor U13495 (N_13495,N_6713,N_3120);
and U13496 (N_13496,N_8537,N_7980);
or U13497 (N_13497,N_5151,N_2472);
xor U13498 (N_13498,N_3073,N_3775);
nor U13499 (N_13499,N_3327,N_8647);
nor U13500 (N_13500,N_5779,N_6273);
nand U13501 (N_13501,N_3739,N_9240);
nor U13502 (N_13502,N_9081,N_9861);
nand U13503 (N_13503,N_4489,N_8371);
or U13504 (N_13504,N_2486,N_8863);
nor U13505 (N_13505,N_824,N_3472);
nand U13506 (N_13506,N_9811,N_8268);
xnor U13507 (N_13507,N_6345,N_2771);
nand U13508 (N_13508,N_6728,N_5570);
nand U13509 (N_13509,N_7491,N_333);
nand U13510 (N_13510,N_9410,N_416);
or U13511 (N_13511,N_6070,N_7085);
and U13512 (N_13512,N_4390,N_7285);
or U13513 (N_13513,N_12,N_1156);
xnor U13514 (N_13514,N_1538,N_4779);
nand U13515 (N_13515,N_2548,N_9131);
or U13516 (N_13516,N_2393,N_8695);
nand U13517 (N_13517,N_6647,N_5859);
xor U13518 (N_13518,N_775,N_8093);
nand U13519 (N_13519,N_7128,N_8168);
or U13520 (N_13520,N_4197,N_1594);
and U13521 (N_13521,N_6920,N_7374);
or U13522 (N_13522,N_8335,N_6972);
nand U13523 (N_13523,N_4345,N_2299);
and U13524 (N_13524,N_8754,N_4733);
xnor U13525 (N_13525,N_3056,N_9302);
xnor U13526 (N_13526,N_6424,N_9608);
nor U13527 (N_13527,N_8731,N_1140);
or U13528 (N_13528,N_2527,N_4856);
nand U13529 (N_13529,N_2740,N_69);
nand U13530 (N_13530,N_5293,N_7310);
xnor U13531 (N_13531,N_8793,N_7217);
nand U13532 (N_13532,N_6327,N_7603);
nor U13533 (N_13533,N_5952,N_4607);
or U13534 (N_13534,N_8114,N_3975);
or U13535 (N_13535,N_9433,N_6635);
and U13536 (N_13536,N_6893,N_6765);
and U13537 (N_13537,N_9851,N_2139);
or U13538 (N_13538,N_7694,N_7872);
xor U13539 (N_13539,N_2581,N_7634);
nor U13540 (N_13540,N_8228,N_8881);
nor U13541 (N_13541,N_7873,N_8632);
nand U13542 (N_13542,N_8723,N_8078);
xnor U13543 (N_13543,N_6227,N_7947);
xnor U13544 (N_13544,N_459,N_5400);
nand U13545 (N_13545,N_2553,N_2748);
xor U13546 (N_13546,N_8338,N_7005);
and U13547 (N_13547,N_2912,N_1350);
xor U13548 (N_13548,N_446,N_8878);
and U13549 (N_13549,N_5006,N_6277);
nand U13550 (N_13550,N_7685,N_4247);
or U13551 (N_13551,N_313,N_9988);
or U13552 (N_13552,N_9642,N_1654);
nand U13553 (N_13553,N_8822,N_525);
nor U13554 (N_13554,N_1226,N_9414);
or U13555 (N_13555,N_3586,N_2770);
nand U13556 (N_13556,N_2187,N_9305);
nor U13557 (N_13557,N_6984,N_8169);
nor U13558 (N_13558,N_6597,N_2557);
and U13559 (N_13559,N_8833,N_7505);
xor U13560 (N_13560,N_9488,N_3804);
or U13561 (N_13561,N_2848,N_9632);
and U13562 (N_13562,N_9474,N_774);
or U13563 (N_13563,N_6571,N_8429);
or U13564 (N_13564,N_26,N_6303);
nor U13565 (N_13565,N_9568,N_6146);
xor U13566 (N_13566,N_9588,N_9329);
or U13567 (N_13567,N_3259,N_7639);
nand U13568 (N_13568,N_7668,N_7769);
xnor U13569 (N_13569,N_9491,N_5614);
or U13570 (N_13570,N_1934,N_4947);
or U13571 (N_13571,N_6129,N_9832);
nand U13572 (N_13572,N_1618,N_433);
and U13573 (N_13573,N_2741,N_62);
nand U13574 (N_13574,N_8513,N_2655);
nor U13575 (N_13575,N_2306,N_6521);
xor U13576 (N_13576,N_1132,N_8618);
xor U13577 (N_13577,N_3348,N_9767);
or U13578 (N_13578,N_382,N_6128);
or U13579 (N_13579,N_7434,N_8445);
nand U13580 (N_13580,N_5870,N_2445);
nand U13581 (N_13581,N_3666,N_6864);
xnor U13582 (N_13582,N_6148,N_3416);
nor U13583 (N_13583,N_8528,N_4202);
nand U13584 (N_13584,N_4561,N_4990);
nor U13585 (N_13585,N_7855,N_3361);
or U13586 (N_13586,N_8241,N_5568);
and U13587 (N_13587,N_95,N_6867);
nor U13588 (N_13588,N_9857,N_2947);
xor U13589 (N_13589,N_2599,N_5115);
nand U13590 (N_13590,N_7875,N_2293);
nor U13591 (N_13591,N_4153,N_8117);
or U13592 (N_13592,N_564,N_7411);
or U13593 (N_13593,N_7083,N_9800);
xnor U13594 (N_13594,N_2728,N_7781);
nor U13595 (N_13595,N_2273,N_3900);
or U13596 (N_13596,N_6928,N_7713);
nor U13597 (N_13597,N_4317,N_9646);
nor U13598 (N_13598,N_2766,N_5972);
xnor U13599 (N_13599,N_9523,N_8935);
xnor U13600 (N_13600,N_3157,N_5761);
or U13601 (N_13601,N_4795,N_9691);
nand U13602 (N_13602,N_8052,N_3861);
or U13603 (N_13603,N_9994,N_6863);
or U13604 (N_13604,N_4516,N_813);
xor U13605 (N_13605,N_6659,N_2850);
and U13606 (N_13606,N_3674,N_9873);
nor U13607 (N_13607,N_1404,N_1779);
nor U13608 (N_13608,N_1017,N_4105);
nand U13609 (N_13609,N_3940,N_2996);
xnor U13610 (N_13610,N_3978,N_4996);
and U13611 (N_13611,N_582,N_1168);
nor U13612 (N_13612,N_5461,N_1758);
xor U13613 (N_13613,N_643,N_466);
nor U13614 (N_13614,N_6565,N_6967);
nand U13615 (N_13615,N_1188,N_7954);
or U13616 (N_13616,N_7047,N_1981);
xnor U13617 (N_13617,N_2731,N_5615);
nor U13618 (N_13618,N_4911,N_9612);
and U13619 (N_13619,N_834,N_7799);
nor U13620 (N_13620,N_8831,N_8370);
xor U13621 (N_13621,N_8510,N_2610);
nand U13622 (N_13622,N_4187,N_7072);
xnor U13623 (N_13623,N_9514,N_8046);
nand U13624 (N_13624,N_737,N_6267);
and U13625 (N_13625,N_5181,N_5592);
or U13626 (N_13626,N_1788,N_9323);
nand U13627 (N_13627,N_3165,N_3067);
and U13628 (N_13628,N_1448,N_7888);
nand U13629 (N_13629,N_3505,N_6292);
xnor U13630 (N_13630,N_6398,N_9094);
nor U13631 (N_13631,N_5493,N_6361);
and U13632 (N_13632,N_1672,N_2291);
and U13633 (N_13633,N_152,N_3719);
or U13634 (N_13634,N_1175,N_2071);
or U13635 (N_13635,N_5609,N_8738);
xnor U13636 (N_13636,N_9385,N_1821);
nor U13637 (N_13637,N_9600,N_573);
and U13638 (N_13638,N_5002,N_3833);
nand U13639 (N_13639,N_5038,N_8782);
xor U13640 (N_13640,N_6817,N_2701);
and U13641 (N_13641,N_7906,N_8641);
nand U13642 (N_13642,N_5940,N_8145);
or U13643 (N_13643,N_8410,N_2045);
xnor U13644 (N_13644,N_8083,N_1108);
nor U13645 (N_13645,N_7750,N_2590);
xor U13646 (N_13646,N_5042,N_8810);
xor U13647 (N_13647,N_3488,N_5487);
nor U13648 (N_13648,N_4087,N_4253);
and U13649 (N_13649,N_4020,N_8680);
or U13650 (N_13650,N_2833,N_809);
xnor U13651 (N_13651,N_2453,N_8576);
and U13652 (N_13652,N_990,N_9783);
or U13653 (N_13653,N_7837,N_614);
xor U13654 (N_13654,N_8427,N_7809);
nand U13655 (N_13655,N_4405,N_6353);
nand U13656 (N_13656,N_8018,N_3183);
nand U13657 (N_13657,N_8424,N_7036);
nor U13658 (N_13658,N_3687,N_9953);
nand U13659 (N_13659,N_8259,N_2355);
xnor U13660 (N_13660,N_6159,N_1947);
xor U13661 (N_13661,N_431,N_4070);
and U13662 (N_13662,N_4050,N_8549);
or U13663 (N_13663,N_2061,N_6113);
and U13664 (N_13664,N_7611,N_1378);
nor U13665 (N_13665,N_980,N_5251);
xnor U13666 (N_13666,N_9677,N_9142);
or U13667 (N_13667,N_224,N_2688);
and U13668 (N_13668,N_4058,N_9173);
or U13669 (N_13669,N_2847,N_3784);
xor U13670 (N_13670,N_497,N_9879);
nor U13671 (N_13671,N_4130,N_4128);
or U13672 (N_13672,N_800,N_3649);
nand U13673 (N_13673,N_5540,N_6869);
and U13674 (N_13674,N_7999,N_1835);
nor U13675 (N_13675,N_696,N_422);
and U13676 (N_13676,N_1366,N_9782);
or U13677 (N_13677,N_1551,N_878);
nand U13678 (N_13678,N_5557,N_7938);
and U13679 (N_13679,N_1547,N_8591);
nand U13680 (N_13680,N_7500,N_2151);
and U13681 (N_13681,N_7348,N_6774);
xor U13682 (N_13682,N_1397,N_3017);
nand U13683 (N_13683,N_7299,N_8396);
and U13684 (N_13684,N_3276,N_6663);
and U13685 (N_13685,N_4335,N_3628);
or U13686 (N_13686,N_3000,N_8469);
or U13687 (N_13687,N_7086,N_3816);
nand U13688 (N_13688,N_1202,N_1574);
nand U13689 (N_13689,N_6311,N_5357);
nand U13690 (N_13690,N_4802,N_4649);
nand U13691 (N_13691,N_3313,N_5174);
or U13692 (N_13692,N_4023,N_1588);
and U13693 (N_13693,N_9138,N_5646);
and U13694 (N_13694,N_8095,N_7758);
or U13695 (N_13695,N_306,N_9072);
nor U13696 (N_13696,N_8874,N_4310);
nor U13697 (N_13697,N_9126,N_5774);
and U13698 (N_13698,N_6805,N_7893);
xor U13699 (N_13699,N_697,N_4866);
xor U13700 (N_13700,N_1962,N_4346);
and U13701 (N_13701,N_1629,N_4134);
and U13702 (N_13702,N_1591,N_2282);
or U13703 (N_13703,N_9119,N_9712);
nand U13704 (N_13704,N_391,N_4703);
nor U13705 (N_13705,N_9365,N_2735);
nor U13706 (N_13706,N_6475,N_4508);
nor U13707 (N_13707,N_2625,N_3122);
or U13708 (N_13708,N_521,N_7609);
nand U13709 (N_13709,N_1198,N_1286);
nand U13710 (N_13710,N_4531,N_4148);
nand U13711 (N_13711,N_9005,N_6868);
nand U13712 (N_13712,N_1874,N_5286);
nor U13713 (N_13713,N_7586,N_8044);
and U13714 (N_13714,N_1382,N_4613);
nor U13715 (N_13715,N_1597,N_2852);
nand U13716 (N_13716,N_3537,N_624);
nand U13717 (N_13717,N_6651,N_7121);
nand U13718 (N_13718,N_1865,N_8900);
or U13719 (N_13719,N_3690,N_6140);
nand U13720 (N_13720,N_3233,N_7977);
nor U13721 (N_13721,N_3680,N_7369);
or U13722 (N_13722,N_3153,N_5866);
nand U13723 (N_13723,N_8626,N_3129);
and U13724 (N_13724,N_5591,N_6561);
nor U13725 (N_13725,N_1085,N_7032);
nor U13726 (N_13726,N_6086,N_7648);
nand U13727 (N_13727,N_5008,N_8244);
or U13728 (N_13728,N_5350,N_3884);
xor U13729 (N_13729,N_8708,N_4307);
xnor U13730 (N_13730,N_4455,N_8939);
xnor U13731 (N_13731,N_7058,N_8234);
or U13732 (N_13732,N_843,N_8013);
and U13733 (N_13733,N_4108,N_6015);
or U13734 (N_13734,N_4267,N_7212);
or U13735 (N_13735,N_8433,N_961);
or U13736 (N_13736,N_3870,N_8687);
and U13737 (N_13737,N_9015,N_7079);
nand U13738 (N_13738,N_9686,N_1097);
or U13739 (N_13739,N_6082,N_5682);
and U13740 (N_13740,N_1501,N_8768);
xor U13741 (N_13741,N_5355,N_3150);
or U13742 (N_13742,N_4892,N_3050);
xor U13743 (N_13743,N_8318,N_1892);
xor U13744 (N_13744,N_9404,N_5228);
xnor U13745 (N_13745,N_7367,N_7196);
nor U13746 (N_13746,N_1469,N_9275);
and U13747 (N_13747,N_6237,N_3413);
and U13748 (N_13748,N_7202,N_8481);
or U13749 (N_13749,N_9666,N_2512);
nor U13750 (N_13750,N_1716,N_4116);
and U13751 (N_13751,N_7151,N_7602);
and U13752 (N_13752,N_6157,N_5714);
xor U13753 (N_13753,N_9270,N_4046);
nand U13754 (N_13754,N_4614,N_4902);
or U13755 (N_13755,N_6471,N_9538);
nand U13756 (N_13756,N_7259,N_2714);
and U13757 (N_13757,N_3188,N_5832);
or U13758 (N_13758,N_1489,N_3548);
nor U13759 (N_13759,N_6553,N_7787);
or U13760 (N_13760,N_2803,N_8209);
xnor U13761 (N_13761,N_664,N_2725);
nand U13762 (N_13762,N_4301,N_4781);
and U13763 (N_13763,N_2822,N_7381);
or U13764 (N_13764,N_7256,N_4415);
or U13765 (N_13765,N_7373,N_7057);
or U13766 (N_13766,N_6552,N_6517);
nand U13767 (N_13767,N_3976,N_8990);
and U13768 (N_13768,N_7672,N_9735);
and U13769 (N_13769,N_9498,N_3190);
xor U13770 (N_13770,N_8697,N_2079);
or U13771 (N_13771,N_3520,N_9965);
or U13772 (N_13772,N_1722,N_4447);
and U13773 (N_13773,N_6331,N_8627);
and U13774 (N_13774,N_9392,N_8849);
nor U13775 (N_13775,N_5590,N_5401);
nor U13776 (N_13776,N_7410,N_1061);
xor U13777 (N_13777,N_9204,N_2871);
or U13778 (N_13778,N_8301,N_4642);
xnor U13779 (N_13779,N_4857,N_3928);
nand U13780 (N_13780,N_361,N_2793);
and U13781 (N_13781,N_5435,N_2939);
nand U13782 (N_13782,N_6502,N_3662);
xor U13783 (N_13783,N_1318,N_9751);
nor U13784 (N_13784,N_4454,N_5236);
xnor U13785 (N_13785,N_1824,N_9791);
or U13786 (N_13786,N_2055,N_5271);
nand U13787 (N_13787,N_6053,N_7329);
xnor U13788 (N_13788,N_5816,N_698);
nor U13789 (N_13789,N_4066,N_9190);
or U13790 (N_13790,N_3033,N_3696);
and U13791 (N_13791,N_5900,N_1689);
xor U13792 (N_13792,N_6798,N_1323);
and U13793 (N_13793,N_4383,N_5102);
or U13794 (N_13794,N_9828,N_6075);
and U13795 (N_13795,N_4078,N_8997);
nand U13796 (N_13796,N_5934,N_6932);
nor U13797 (N_13797,N_8985,N_1866);
xor U13798 (N_13798,N_6907,N_355);
xnor U13799 (N_13799,N_7252,N_6595);
nor U13800 (N_13800,N_8165,N_3931);
and U13801 (N_13801,N_2100,N_9643);
and U13802 (N_13802,N_9531,N_1799);
and U13803 (N_13803,N_3444,N_7849);
nor U13804 (N_13804,N_377,N_8069);
nand U13805 (N_13805,N_1509,N_3453);
and U13806 (N_13806,N_8924,N_5054);
xnor U13807 (N_13807,N_2998,N_2915);
and U13808 (N_13808,N_6444,N_7897);
nor U13809 (N_13809,N_3750,N_4660);
or U13810 (N_13810,N_3187,N_2223);
or U13811 (N_13811,N_3336,N_76);
nand U13812 (N_13812,N_7484,N_5710);
and U13813 (N_13813,N_3853,N_8260);
nand U13814 (N_13814,N_9068,N_4094);
or U13815 (N_13815,N_9033,N_9760);
nor U13816 (N_13816,N_1052,N_5484);
xnor U13817 (N_13817,N_5790,N_9847);
xor U13818 (N_13818,N_5577,N_9829);
xnor U13819 (N_13819,N_986,N_6162);
or U13820 (N_13820,N_2902,N_7460);
nand U13821 (N_13821,N_5960,N_9035);
xor U13822 (N_13822,N_8432,N_5201);
xnor U13823 (N_13823,N_2245,N_3991);
xor U13824 (N_13824,N_1442,N_9870);
and U13825 (N_13825,N_2257,N_6430);
and U13826 (N_13826,N_1253,N_6451);
or U13827 (N_13827,N_5339,N_6414);
xnor U13828 (N_13828,N_7179,N_2209);
or U13829 (N_13829,N_4591,N_2604);
or U13830 (N_13830,N_5915,N_7613);
nand U13831 (N_13831,N_2857,N_8739);
and U13832 (N_13832,N_260,N_4612);
nor U13833 (N_13833,N_3597,N_5055);
nand U13834 (N_13834,N_7546,N_2723);
nor U13835 (N_13835,N_6638,N_5725);
xor U13836 (N_13836,N_9387,N_6944);
nand U13837 (N_13837,N_6365,N_2429);
nand U13838 (N_13838,N_5930,N_1169);
and U13839 (N_13839,N_5488,N_7307);
xnor U13840 (N_13840,N_2772,N_7385);
xor U13841 (N_13841,N_9017,N_5636);
nand U13842 (N_13842,N_862,N_7238);
nor U13843 (N_13843,N_4025,N_3905);
nand U13844 (N_13844,N_428,N_3443);
and U13845 (N_13845,N_5409,N_9753);
and U13846 (N_13846,N_4037,N_618);
or U13847 (N_13847,N_5463,N_6486);
and U13848 (N_13848,N_2691,N_4117);
xnor U13849 (N_13849,N_3504,N_5962);
nand U13850 (N_13850,N_109,N_185);
xnor U13851 (N_13851,N_9973,N_1196);
or U13852 (N_13852,N_3523,N_6671);
nor U13853 (N_13853,N_5301,N_6018);
or U13854 (N_13854,N_3343,N_2034);
and U13855 (N_13855,N_9558,N_5144);
or U13856 (N_13856,N_3064,N_700);
nor U13857 (N_13857,N_1281,N_9370);
nor U13858 (N_13858,N_385,N_5519);
nand U13859 (N_13859,N_9594,N_6413);
xnor U13860 (N_13860,N_3304,N_4186);
xor U13861 (N_13861,N_6586,N_6679);
and U13862 (N_13862,N_5009,N_1394);
or U13863 (N_13863,N_4929,N_3759);
nand U13864 (N_13864,N_3220,N_400);
nor U13865 (N_13865,N_6694,N_4735);
and U13866 (N_13866,N_8187,N_4835);
and U13867 (N_13867,N_5511,N_4062);
and U13868 (N_13868,N_2356,N_1639);
nand U13869 (N_13869,N_1521,N_3866);
and U13870 (N_13870,N_9774,N_4339);
or U13871 (N_13871,N_1586,N_1871);
xnor U13872 (N_13872,N_4004,N_3764);
and U13873 (N_13873,N_4980,N_5585);
and U13874 (N_13874,N_1136,N_972);
and U13875 (N_13875,N_7901,N_7230);
nand U13876 (N_13876,N_6199,N_5156);
nand U13877 (N_13877,N_134,N_3246);
nand U13878 (N_13878,N_8493,N_5531);
nand U13879 (N_13879,N_3676,N_511);
nand U13880 (N_13880,N_9102,N_5290);
nor U13881 (N_13881,N_8293,N_6065);
or U13882 (N_13882,N_5126,N_9895);
nand U13883 (N_13883,N_9042,N_757);
nor U13884 (N_13884,N_429,N_7206);
xor U13885 (N_13885,N_8324,N_5639);
xor U13886 (N_13886,N_559,N_3725);
and U13887 (N_13887,N_1171,N_1630);
xor U13888 (N_13888,N_3947,N_2510);
nor U13889 (N_13889,N_1080,N_4469);
xor U13890 (N_13890,N_3899,N_8129);
and U13891 (N_13891,N_6843,N_2140);
xor U13892 (N_13892,N_3346,N_577);
xnor U13893 (N_13893,N_8313,N_9038);
or U13894 (N_13894,N_6341,N_4238);
xnor U13895 (N_13895,N_1351,N_1857);
nand U13896 (N_13896,N_754,N_6768);
xor U13897 (N_13897,N_7034,N_9012);
nand U13898 (N_13898,N_1268,N_5137);
or U13899 (N_13899,N_7354,N_3704);
nor U13900 (N_13900,N_9615,N_4360);
nand U13901 (N_13901,N_1079,N_4288);
nor U13902 (N_13902,N_4989,N_674);
nand U13903 (N_13903,N_9504,N_1314);
xor U13904 (N_13904,N_7490,N_9957);
xnor U13905 (N_13905,N_8292,N_4340);
nor U13906 (N_13906,N_7461,N_4748);
nand U13907 (N_13907,N_6312,N_6367);
and U13908 (N_13908,N_5155,N_211);
nand U13909 (N_13909,N_2268,N_9348);
xnor U13910 (N_13910,N_2278,N_1309);
and U13911 (N_13911,N_2446,N_8041);
or U13912 (N_13912,N_9905,N_3186);
nand U13913 (N_13913,N_7964,N_6126);
nor U13914 (N_13914,N_6033,N_4378);
xor U13915 (N_13915,N_8870,N_4767);
nor U13916 (N_13916,N_5224,N_9218);
and U13917 (N_13917,N_1790,N_4089);
nor U13918 (N_13918,N_1334,N_5953);
and U13919 (N_13919,N_5422,N_2361);
or U13920 (N_13920,N_6287,N_2943);
nand U13921 (N_13921,N_6735,N_9346);
nand U13922 (N_13922,N_750,N_3499);
xnor U13923 (N_13923,N_9638,N_6048);
or U13924 (N_13924,N_5064,N_8588);
nand U13925 (N_13925,N_2277,N_5421);
nor U13926 (N_13926,N_4903,N_46);
or U13927 (N_13927,N_9640,N_6356);
nor U13928 (N_13928,N_1385,N_7926);
or U13929 (N_13929,N_7396,N_7113);
nor U13930 (N_13930,N_4446,N_1744);
or U13931 (N_13931,N_3671,N_5800);
xnor U13932 (N_13932,N_2663,N_2366);
nand U13933 (N_13933,N_8008,N_5573);
nor U13934 (N_13934,N_4644,N_9562);
nand U13935 (N_13935,N_7560,N_2672);
xnor U13936 (N_13936,N_4141,N_2671);
and U13937 (N_13937,N_6991,N_3408);
or U13938 (N_13938,N_4290,N_4539);
and U13939 (N_13939,N_3733,N_129);
nand U13940 (N_13940,N_7214,N_312);
or U13941 (N_13941,N_8016,N_7813);
and U13942 (N_13942,N_4086,N_3496);
xor U13943 (N_13943,N_3955,N_7017);
xor U13944 (N_13944,N_7006,N_3236);
nor U13945 (N_13945,N_8961,N_8636);
nand U13946 (N_13946,N_5353,N_9846);
xor U13947 (N_13947,N_1082,N_8199);
nor U13948 (N_13948,N_5803,N_2605);
nand U13949 (N_13949,N_6608,N_4374);
xor U13950 (N_13950,N_3989,N_2897);
nand U13951 (N_13951,N_1237,N_4347);
xor U13952 (N_13952,N_4922,N_9729);
nor U13953 (N_13953,N_6014,N_936);
nand U13954 (N_13954,N_1361,N_2816);
or U13955 (N_13955,N_5465,N_7674);
nand U13956 (N_13956,N_3595,N_1906);
nor U13957 (N_13957,N_8938,N_5300);
nand U13958 (N_13958,N_9454,N_4742);
nand U13959 (N_13959,N_384,N_8638);
nand U13960 (N_13960,N_7973,N_3099);
nand U13961 (N_13961,N_4515,N_1863);
xnor U13962 (N_13962,N_3226,N_4048);
xnor U13963 (N_13963,N_2921,N_8566);
nor U13964 (N_13964,N_9457,N_629);
and U13965 (N_13965,N_2970,N_7181);
and U13966 (N_13966,N_2037,N_8904);
nor U13967 (N_13967,N_764,N_3250);
xor U13968 (N_13968,N_7305,N_2207);
nor U13969 (N_13969,N_8321,N_738);
xor U13970 (N_13970,N_5247,N_652);
xor U13971 (N_13971,N_6731,N_7537);
nand U13972 (N_13972,N_4149,N_5985);
and U13973 (N_13973,N_1648,N_9006);
nor U13974 (N_13974,N_8213,N_6364);
xnor U13975 (N_13975,N_4618,N_5106);
xor U13976 (N_13976,N_4962,N_8540);
xnor U13977 (N_13977,N_7404,N_6952);
xor U13978 (N_13978,N_9693,N_8229);
nor U13979 (N_13979,N_9614,N_7783);
nor U13980 (N_13980,N_9853,N_448);
nor U13981 (N_13981,N_4814,N_3797);
xnor U13982 (N_13982,N_4326,N_2129);
xor U13983 (N_13983,N_8245,N_8771);
and U13984 (N_13984,N_3743,N_4395);
or U13985 (N_13985,N_4874,N_4575);
nand U13986 (N_13986,N_491,N_6603);
nor U13987 (N_13987,N_4357,N_9986);
nand U13988 (N_13988,N_359,N_3757);
nor U13989 (N_13989,N_7495,N_5100);
nand U13990 (N_13990,N_1162,N_930);
xor U13991 (N_13991,N_6987,N_8829);
xnor U13992 (N_13992,N_7757,N_5324);
and U13993 (N_13993,N_6772,N_5306);
and U13994 (N_13994,N_7941,N_5230);
and U13995 (N_13995,N_7959,N_7429);
nand U13996 (N_13996,N_1695,N_519);
and U13997 (N_13997,N_2056,N_9775);
xnor U13998 (N_13998,N_3490,N_6115);
xnor U13999 (N_13999,N_2776,N_7870);
xor U14000 (N_14000,N_5571,N_7649);
and U14001 (N_14001,N_6255,N_8028);
xnor U14002 (N_14002,N_100,N_1214);
nand U14003 (N_14003,N_6598,N_4344);
and U14004 (N_14004,N_7535,N_7608);
nor U14005 (N_14005,N_8668,N_5947);
nor U14006 (N_14006,N_8272,N_8891);
or U14007 (N_14007,N_7481,N_9308);
or U14008 (N_14008,N_6351,N_2265);
and U14009 (N_14009,N_7458,N_2821);
and U14010 (N_14010,N_5217,N_6045);
nor U14011 (N_14011,N_4626,N_6217);
xor U14012 (N_14012,N_7439,N_9637);
nor U14013 (N_14013,N_2114,N_8960);
nor U14014 (N_14014,N_8136,N_8851);
xor U14015 (N_14015,N_9379,N_8278);
xnor U14016 (N_14016,N_3206,N_6922);
nand U14017 (N_14017,N_1715,N_321);
and U14018 (N_14018,N_5607,N_4640);
nand U14019 (N_14019,N_9287,N_7552);
and U14020 (N_14020,N_6614,N_6885);
nand U14021 (N_14021,N_7740,N_6462);
nor U14022 (N_14022,N_4737,N_3069);
and U14023 (N_14023,N_5430,N_4639);
xor U14024 (N_14024,N_5184,N_8249);
nor U14025 (N_14025,N_7049,N_45);
nor U14026 (N_14026,N_6460,N_7028);
or U14027 (N_14027,N_4978,N_3333);
nor U14028 (N_14028,N_6894,N_3808);
and U14029 (N_14029,N_7638,N_8239);
and U14030 (N_14030,N_5892,N_3382);
nor U14031 (N_14031,N_4570,N_669);
and U14032 (N_14032,N_2068,N_2399);
and U14033 (N_14033,N_9801,N_9746);
xnor U14034 (N_14034,N_7050,N_6784);
nand U14035 (N_14035,N_2963,N_1371);
nand U14036 (N_14036,N_9484,N_3357);
and U14037 (N_14037,N_5656,N_2083);
xor U14038 (N_14038,N_6989,N_1601);
nand U14039 (N_14039,N_9697,N_173);
xnor U14040 (N_14040,N_4833,N_7477);
xnor U14041 (N_14041,N_8263,N_9819);
xor U14042 (N_14042,N_9702,N_7194);
xor U14043 (N_14043,N_2526,N_1975);
xor U14044 (N_14044,N_7677,N_8612);
and U14045 (N_14045,N_5747,N_9758);
and U14046 (N_14046,N_5748,N_7018);
xor U14047 (N_14047,N_625,N_6942);
nor U14048 (N_14048,N_1392,N_6544);
and U14049 (N_14049,N_4505,N_1784);
nor U14050 (N_14050,N_4790,N_2357);
or U14051 (N_14051,N_8079,N_2411);
and U14052 (N_14052,N_2631,N_7512);
nand U14053 (N_14053,N_7935,N_8579);
and U14054 (N_14054,N_8434,N_7278);
xnor U14055 (N_14055,N_1937,N_7806);
and U14056 (N_14056,N_258,N_1827);
nand U14057 (N_14057,N_5629,N_6884);
nand U14058 (N_14058,N_8978,N_2928);
nor U14059 (N_14059,N_272,N_9650);
or U14060 (N_14060,N_7098,N_8853);
and U14061 (N_14061,N_7039,N_8719);
and U14062 (N_14062,N_94,N_2216);
or U14063 (N_14063,N_4407,N_7735);
nor U14064 (N_14064,N_6407,N_1570);
or U14065 (N_14065,N_9773,N_8714);
xor U14066 (N_14066,N_1675,N_9318);
nor U14067 (N_14067,N_598,N_8673);
or U14068 (N_14068,N_4262,N_5233);
nor U14069 (N_14069,N_791,N_8120);
or U14070 (N_14070,N_6696,N_2436);
nor U14071 (N_14071,N_3139,N_1958);
or U14072 (N_14072,N_3239,N_9449);
nand U14073 (N_14073,N_7681,N_7453);
nand U14074 (N_14074,N_30,N_4504);
or U14075 (N_14075,N_1759,N_4302);
nor U14076 (N_14076,N_3841,N_2031);
xor U14077 (N_14077,N_9225,N_3563);
and U14078 (N_14078,N_3063,N_3511);
and U14079 (N_14079,N_5801,N_6618);
xnor U14080 (N_14080,N_1042,N_1400);
xor U14081 (N_14081,N_9299,N_6572);
nand U14082 (N_14082,N_7915,N_7182);
nor U14083 (N_14083,N_1265,N_7993);
or U14084 (N_14084,N_2403,N_9353);
nor U14085 (N_14085,N_6491,N_1539);
nor U14086 (N_14086,N_8221,N_9975);
nand U14087 (N_14087,N_1976,N_3131);
or U14088 (N_14088,N_5420,N_7430);
and U14089 (N_14089,N_3442,N_8590);
nand U14090 (N_14090,N_5686,N_4082);
nand U14091 (N_14091,N_4661,N_7334);
and U14092 (N_14092,N_2440,N_4512);
xnor U14093 (N_14093,N_66,N_9996);
xnor U14094 (N_14094,N_1211,N_4961);
xor U14095 (N_14095,N_2914,N_5922);
nor U14096 (N_14096,N_6526,N_4745);
or U14097 (N_14097,N_6171,N_8112);
and U14098 (N_14098,N_3405,N_2820);
nand U14099 (N_14099,N_2878,N_7242);
nand U14100 (N_14100,N_5906,N_9586);
xor U14101 (N_14101,N_1556,N_3415);
nand U14102 (N_14102,N_2508,N_7623);
and U14103 (N_14103,N_9741,N_3491);
or U14104 (N_14104,N_2262,N_3612);
nor U14105 (N_14105,N_9321,N_3199);
xnor U14106 (N_14106,N_77,N_7595);
nor U14107 (N_14107,N_6450,N_2643);
xor U14108 (N_14108,N_5908,N_3340);
or U14109 (N_14109,N_2578,N_9467);
or U14110 (N_14110,N_8033,N_1891);
or U14111 (N_14111,N_6134,N_8451);
nand U14112 (N_14112,N_9480,N_4787);
nor U14113 (N_14113,N_5431,N_5334);
nor U14114 (N_14114,N_5673,N_2315);
nand U14115 (N_14115,N_2706,N_2210);
and U14116 (N_14116,N_4773,N_7981);
or U14117 (N_14117,N_3778,N_9711);
xor U14118 (N_14118,N_1133,N_9245);
nor U14119 (N_14119,N_9855,N_3907);
and U14120 (N_14120,N_7723,N_2880);
or U14121 (N_14121,N_1842,N_4720);
and U14122 (N_14122,N_4373,N_1447);
and U14123 (N_14123,N_5428,N_2444);
nor U14124 (N_14124,N_4323,N_5996);
nor U14125 (N_14125,N_4812,N_3085);
nand U14126 (N_14126,N_969,N_8984);
nand U14127 (N_14127,N_1796,N_7755);
nor U14128 (N_14128,N_8504,N_6545);
nor U14129 (N_14129,N_1808,N_6363);
nor U14130 (N_14130,N_157,N_9170);
or U14131 (N_14131,N_8890,N_9328);
and U14132 (N_14132,N_5974,N_1726);
nor U14133 (N_14133,N_5534,N_1778);
or U14134 (N_14134,N_8102,N_9377);
and U14135 (N_14135,N_2493,N_7693);
and U14136 (N_14136,N_2051,N_8575);
and U14137 (N_14137,N_8294,N_7578);
or U14138 (N_14138,N_7545,N_3558);
or U14139 (N_14139,N_3339,N_1056);
xor U14140 (N_14140,N_6658,N_9950);
nand U14141 (N_14141,N_1275,N_3960);
nand U14142 (N_14142,N_9892,N_2781);
nand U14143 (N_14143,N_6690,N_2101);
xor U14144 (N_14144,N_2764,N_1151);
nand U14145 (N_14145,N_6749,N_9067);
xnor U14146 (N_14146,N_3943,N_9243);
nor U14147 (N_14147,N_6456,N_9901);
xor U14148 (N_14148,N_702,N_5191);
xnor U14149 (N_14149,N_3863,N_5089);
or U14150 (N_14150,N_9494,N_442);
nand U14151 (N_14151,N_2948,N_7075);
nor U14152 (N_14152,N_2917,N_2153);
xnor U14153 (N_14153,N_5661,N_9478);
or U14154 (N_14154,N_8743,N_5738);
nor U14155 (N_14155,N_6002,N_908);
and U14156 (N_14156,N_1118,N_1005);
or U14157 (N_14157,N_4528,N_9960);
nor U14158 (N_14158,N_7670,N_778);
xnor U14159 (N_14159,N_7749,N_1771);
nor U14160 (N_14160,N_8420,N_1650);
and U14161 (N_14161,N_6136,N_998);
nand U14162 (N_14162,N_9663,N_2360);
nand U14163 (N_14163,N_5378,N_1900);
nand U14164 (N_14164,N_5030,N_2785);
nand U14165 (N_14165,N_8466,N_467);
or U14166 (N_14166,N_2812,N_7322);
nor U14167 (N_14167,N_5347,N_1719);
or U14168 (N_14168,N_1413,N_4571);
nor U14169 (N_14169,N_6229,N_7759);
xnor U14170 (N_14170,N_7356,N_5508);
nand U14171 (N_14171,N_2845,N_8040);
nand U14172 (N_14172,N_8220,N_1173);
or U14173 (N_14173,N_369,N_4717);
xor U14174 (N_14174,N_6966,N_4355);
and U14175 (N_14175,N_5660,N_8006);
and U14176 (N_14176,N_493,N_938);
or U14177 (N_14177,N_189,N_8608);
xnor U14178 (N_14178,N_3825,N_7987);
and U14179 (N_14179,N_4016,N_1637);
or U14180 (N_14180,N_7473,N_6275);
xnor U14181 (N_14181,N_6314,N_9424);
nand U14182 (N_14182,N_9845,N_2476);
xnor U14183 (N_14183,N_8682,N_4865);
xor U14184 (N_14184,N_2160,N_4261);
nor U14185 (N_14185,N_3856,N_5553);
or U14186 (N_14186,N_5314,N_7188);
or U14187 (N_14187,N_4379,N_2447);
and U14188 (N_14188,N_9446,N_81);
and U14189 (N_14189,N_9671,N_632);
xnor U14190 (N_14190,N_6996,N_4680);
nand U14191 (N_14191,N_5336,N_6378);
or U14192 (N_14192,N_8595,N_4325);
nor U14193 (N_14193,N_4999,N_128);
and U14194 (N_14194,N_9500,N_9683);
or U14195 (N_14195,N_9143,N_790);
xnor U14196 (N_14196,N_6224,N_1);
nor U14197 (N_14197,N_7853,N_4670);
nor U14198 (N_14198,N_9419,N_4919);
xnor U14199 (N_14199,N_5688,N_661);
nand U14200 (N_14200,N_2200,N_1930);
or U14201 (N_14201,N_1137,N_6370);
and U14202 (N_14202,N_304,N_8953);
and U14203 (N_14203,N_9820,N_2568);
and U14204 (N_14204,N_3983,N_6615);
xor U14205 (N_14205,N_4600,N_3936);
nand U14206 (N_14206,N_971,N_3319);
or U14207 (N_14207,N_8312,N_2759);
xor U14208 (N_14208,N_9968,N_6627);
xnor U14209 (N_14209,N_199,N_3462);
xor U14210 (N_14210,N_3011,N_6632);
nor U14211 (N_14211,N_5496,N_5837);
nand U14212 (N_14212,N_2682,N_8299);
and U14213 (N_14213,N_3894,N_4234);
nor U14214 (N_14214,N_1038,N_6141);
or U14215 (N_14215,N_2783,N_3041);
xor U14216 (N_14216,N_2364,N_2430);
and U14217 (N_14217,N_9014,N_4467);
xnor U14218 (N_14218,N_9178,N_6596);
nor U14219 (N_14219,N_6673,N_4018);
or U14220 (N_14220,N_8905,N_9959);
or U14221 (N_14221,N_6081,N_9064);
nand U14222 (N_14222,N_6016,N_200);
or U14223 (N_14223,N_8109,N_6770);
nand U14224 (N_14224,N_434,N_65);
or U14225 (N_14225,N_8894,N_6274);
xor U14226 (N_14226,N_9623,N_5015);
nor U14227 (N_14227,N_5053,N_9193);
nor U14228 (N_14228,N_7530,N_5059);
nor U14229 (N_14229,N_1984,N_1651);
and U14230 (N_14230,N_5830,N_3823);
nand U14231 (N_14231,N_3263,N_1653);
or U14232 (N_14232,N_4033,N_2457);
nand U14233 (N_14233,N_3677,N_5971);
and U14234 (N_14234,N_353,N_5303);
nor U14235 (N_14235,N_5473,N_9383);
or U14236 (N_14236,N_6009,N_6382);
nand U14237 (N_14237,N_8778,N_5654);
and U14238 (N_14238,N_7020,N_3248);
nor U14239 (N_14239,N_3002,N_1258);
and U14240 (N_14240,N_6736,N_1992);
nand U14241 (N_14241,N_399,N_1032);
or U14242 (N_14242,N_4178,N_9088);
or U14243 (N_14243,N_7626,N_8022);
and U14244 (N_14244,N_2632,N_386);
or U14245 (N_14245,N_5931,N_1468);
and U14246 (N_14246,N_5527,N_6937);
or U14247 (N_14247,N_8364,N_7275);
or U14248 (N_14248,N_9018,N_4457);
nor U14249 (N_14249,N_4747,N_6858);
or U14250 (N_14250,N_772,N_7090);
nand U14251 (N_14251,N_7652,N_7555);
xnor U14252 (N_14252,N_2169,N_7112);
nor U14253 (N_14253,N_2719,N_530);
and U14254 (N_14254,N_2422,N_7734);
nand U14255 (N_14255,N_1248,N_3332);
or U14256 (N_14256,N_2777,N_4371);
xnor U14257 (N_14257,N_6299,N_5775);
and U14258 (N_14258,N_5399,N_1244);
or U14259 (N_14259,N_3144,N_758);
nor U14260 (N_14260,N_4316,N_9409);
and U14261 (N_14261,N_5771,N_1433);
or U14262 (N_14262,N_6087,N_1029);
nor U14263 (N_14263,N_9013,N_2052);
nor U14264 (N_14264,N_7313,N_8350);
nand U14265 (N_14265,N_1149,N_905);
or U14266 (N_14266,N_4723,N_4028);
nor U14267 (N_14267,N_2023,N_237);
or U14268 (N_14268,N_1364,N_5795);
nor U14269 (N_14269,N_9756,N_8649);
nand U14270 (N_14270,N_8237,N_5561);
and U14271 (N_14271,N_9376,N_6318);
and U14272 (N_14272,N_3279,N_7720);
nor U14273 (N_14273,N_4118,N_2416);
nand U14274 (N_14274,N_7792,N_4507);
xnor U14275 (N_14275,N_4501,N_2205);
nand U14276 (N_14276,N_2543,N_7393);
xor U14277 (N_14277,N_760,N_4104);
nand U14278 (N_14278,N_3873,N_5214);
xor U14279 (N_14279,N_3110,N_1235);
nor U14280 (N_14280,N_2563,N_2968);
xor U14281 (N_14281,N_4074,N_4871);
and U14282 (N_14282,N_7644,N_6759);
nand U14283 (N_14283,N_4274,N_9878);
nor U14284 (N_14284,N_622,N_5450);
nor U14285 (N_14285,N_2424,N_6094);
xnor U14286 (N_14286,N_5035,N_5140);
and U14287 (N_14287,N_7661,N_2116);
and U14288 (N_14288,N_4709,N_6241);
and U14289 (N_14289,N_1306,N_9648);
xor U14290 (N_14290,N_7620,N_6350);
and U14291 (N_14291,N_3317,N_5323);
nand U14292 (N_14292,N_3,N_3040);
and U14293 (N_14293,N_9548,N_3727);
nand U14294 (N_14294,N_119,N_1971);
xor U14295 (N_14295,N_8257,N_856);
nand U14296 (N_14296,N_8480,N_4304);
nor U14297 (N_14297,N_6402,N_2115);
and U14298 (N_14298,N_5848,N_110);
and U14299 (N_14299,N_9651,N_6832);
xor U14300 (N_14300,N_9293,N_3576);
xnor U14301 (N_14301,N_1552,N_3030);
and U14302 (N_14302,N_9002,N_720);
nor U14303 (N_14303,N_5510,N_3437);
nand U14304 (N_14304,N_7455,N_2456);
nand U14305 (N_14305,N_1889,N_886);
and U14306 (N_14306,N_8376,N_6465);
nor U14307 (N_14307,N_9222,N_6235);
xnor U14308 (N_14308,N_7074,N_777);
and U14309 (N_14309,N_6532,N_2035);
xor U14310 (N_14310,N_6305,N_5705);
nor U14311 (N_14311,N_8198,N_3141);
and U14312 (N_14312,N_9633,N_2961);
and U14313 (N_14313,N_4609,N_7137);
nand U14314 (N_14314,N_4676,N_6787);
and U14315 (N_14315,N_3815,N_2762);
or U14316 (N_14316,N_7391,N_1957);
and U14317 (N_14317,N_1734,N_7163);
xor U14318 (N_14318,N_9817,N_4268);
nand U14319 (N_14319,N_8323,N_9009);
nor U14320 (N_14320,N_2662,N_515);
or U14321 (N_14321,N_1809,N_5349);
and U14322 (N_14322,N_5547,N_7372);
nand U14323 (N_14323,N_8785,N_3885);
xnor U14324 (N_14324,N_6286,N_8801);
nand U14325 (N_14325,N_8357,N_4526);
nand U14326 (N_14326,N_7636,N_5604);
nand U14327 (N_14327,N_5864,N_8889);
and U14328 (N_14328,N_7472,N_8099);
nor U14329 (N_14329,N_1014,N_2338);
xor U14330 (N_14330,N_5857,N_7269);
xor U14331 (N_14331,N_2462,N_5559);
nand U14332 (N_14332,N_7288,N_2287);
nand U14333 (N_14333,N_7905,N_8750);
xnor U14334 (N_14334,N_9191,N_8368);
and U14335 (N_14335,N_7807,N_1336);
and U14336 (N_14336,N_4690,N_2615);
xnor U14337 (N_14337,N_4367,N_6419);
or U14338 (N_14338,N_5796,N_4831);
and U14339 (N_14339,N_4931,N_6992);
and U14340 (N_14340,N_4611,N_34);
nand U14341 (N_14341,N_9635,N_4184);
nor U14342 (N_14342,N_884,N_4024);
nand U14343 (N_14343,N_2733,N_5752);
nor U14344 (N_14344,N_2879,N_6410);
or U14345 (N_14345,N_1091,N_7068);
and U14346 (N_14346,N_7365,N_3579);
nand U14347 (N_14347,N_9602,N_3532);
nand U14348 (N_14348,N_6842,N_5765);
nand U14349 (N_14349,N_1756,N_4849);
xor U14350 (N_14350,N_658,N_2255);
or U14351 (N_14351,N_51,N_5632);
nand U14352 (N_14352,N_1081,N_9678);
nor U14353 (N_14353,N_8491,N_5394);
or U14354 (N_14354,N_3072,N_7924);
nor U14355 (N_14355,N_522,N_9983);
nor U14356 (N_14356,N_9555,N_5292);
nor U14357 (N_14357,N_8310,N_7975);
xor U14358 (N_14358,N_5956,N_2621);
xnor U14359 (N_14359,N_91,N_2261);
xor U14360 (N_14360,N_4190,N_1698);
or U14361 (N_14361,N_6753,N_9239);
and U14362 (N_14362,N_9603,N_7386);
xnor U14363 (N_14363,N_8094,N_6470);
or U14364 (N_14364,N_3543,N_8651);
and U14365 (N_14365,N_6516,N_1797);
xnor U14366 (N_14366,N_4448,N_4434);
nand U14367 (N_14367,N_7967,N_612);
nand U14368 (N_14368,N_8111,N_2069);
or U14369 (N_14369,N_6559,N_1206);
and U14370 (N_14370,N_8539,N_2609);
and U14371 (N_14371,N_5325,N_3618);
or U14372 (N_14372,N_4163,N_9340);
and U14373 (N_14373,N_6099,N_3383);
or U14374 (N_14374,N_5544,N_8677);
and U14375 (N_14375,N_9145,N_9629);
nand U14376 (N_14376,N_221,N_6576);
and U14377 (N_14377,N_7443,N_8054);
nand U14378 (N_14378,N_9692,N_2983);
nand U14379 (N_14379,N_597,N_7448);
or U14380 (N_14380,N_4293,N_1142);
xor U14381 (N_14381,N_8286,N_1507);
nor U14382 (N_14382,N_6706,N_7432);
nor U14383 (N_14383,N_9564,N_5902);
and U14384 (N_14384,N_7119,N_3059);
nor U14385 (N_14385,N_2906,N_7767);
xnor U14386 (N_14386,N_7001,N_3234);
and U14387 (N_14387,N_928,N_4734);
nor U14388 (N_14388,N_8621,N_9860);
and U14389 (N_14389,N_3811,N_485);
and U14390 (N_14390,N_9869,N_257);
xor U14391 (N_14391,N_9824,N_8164);
and U14392 (N_14392,N_6102,N_9713);
nor U14393 (N_14393,N_8520,N_3076);
or U14394 (N_14394,N_1699,N_7406);
nor U14395 (N_14395,N_6558,N_7441);
nand U14396 (N_14396,N_9395,N_8989);
xor U14397 (N_14397,N_6435,N_5004);
and U14398 (N_14398,N_2142,N_1183);
nand U14399 (N_14399,N_724,N_244);
nor U14400 (N_14400,N_2094,N_7751);
xnor U14401 (N_14401,N_7797,N_8435);
nor U14402 (N_14402,N_1303,N_9515);
and U14403 (N_14403,N_1233,N_2193);
or U14404 (N_14404,N_7606,N_9682);
nor U14405 (N_14405,N_4689,N_1641);
xor U14406 (N_14406,N_3802,N_873);
or U14407 (N_14407,N_3503,N_3119);
nor U14408 (N_14408,N_937,N_3726);
nand U14409 (N_14409,N_4805,N_5262);
nand U14410 (N_14410,N_6662,N_2987);
xnor U14411 (N_14411,N_454,N_4125);
nand U14412 (N_14412,N_528,N_6272);
nand U14413 (N_14413,N_5472,N_8770);
nand U14414 (N_14414,N_7037,N_2066);
and U14415 (N_14415,N_3742,N_7078);
nand U14416 (N_14416,N_8369,N_7777);
nor U14417 (N_14417,N_5740,N_9136);
nand U14418 (N_14418,N_1086,N_5522);
or U14419 (N_14419,N_4054,N_9434);
and U14420 (N_14420,N_84,N_2778);
nand U14421 (N_14421,N_3583,N_4877);
nor U14422 (N_14422,N_5702,N_9601);
or U14423 (N_14423,N_5606,N_7900);
nor U14424 (N_14424,N_1229,N_3482);
nand U14425 (N_14425,N_8987,N_5520);
and U14426 (N_14426,N_4910,N_1463);
nor U14427 (N_14427,N_1197,N_121);
xor U14428 (N_14428,N_5032,N_6054);
and U14429 (N_14429,N_1002,N_450);
or U14430 (N_14430,N_880,N_9280);
nand U14431 (N_14431,N_1322,N_8302);
nor U14432 (N_14432,N_9789,N_6852);
xor U14433 (N_14433,N_2251,N_7320);
nor U14434 (N_14434,N_7907,N_5689);
and U14435 (N_14435,N_9814,N_8447);
nand U14436 (N_14436,N_8530,N_5093);
nand U14437 (N_14437,N_3843,N_7304);
or U14438 (N_14438,N_1836,N_2352);
or U14439 (N_14439,N_6408,N_8393);
nor U14440 (N_14440,N_2040,N_1024);
nor U14441 (N_14441,N_818,N_1907);
xnor U14442 (N_14442,N_3312,N_6202);
and U14443 (N_14443,N_1283,N_4499);
nand U14444 (N_14444,N_213,N_4464);
and U14445 (N_14445,N_1691,N_851);
xnor U14446 (N_14446,N_8789,N_9520);
nor U14447 (N_14447,N_6247,N_506);
or U14448 (N_14448,N_8784,N_8908);
xnor U14449 (N_14449,N_3354,N_516);
and U14450 (N_14450,N_4532,N_5672);
nand U14451 (N_14451,N_5943,N_350);
or U14452 (N_14452,N_1952,N_2120);
nand U14453 (N_14453,N_4704,N_6358);
nor U14454 (N_14454,N_1034,N_7895);
xor U14455 (N_14455,N_770,N_460);
nor U14456 (N_14456,N_6716,N_672);
nor U14457 (N_14457,N_5611,N_3218);
nor U14458 (N_14458,N_2773,N_9361);
or U14459 (N_14459,N_5485,N_5821);
and U14460 (N_14460,N_7243,N_4259);
or U14461 (N_14461,N_765,N_9927);
nand U14462 (N_14462,N_8920,N_2805);
xnor U14463 (N_14463,N_6231,N_7294);
nand U14464 (N_14464,N_140,N_8700);
or U14465 (N_14465,N_8783,N_2455);
xnor U14466 (N_14466,N_501,N_7881);
and U14467 (N_14467,N_8280,N_1850);
or U14468 (N_14468,N_6590,N_1964);
and U14469 (N_14469,N_3573,N_1497);
nand U14470 (N_14470,N_6155,N_2224);
or U14471 (N_14471,N_4075,N_4196);
nand U14472 (N_14472,N_3806,N_2698);
xnor U14473 (N_14473,N_8600,N_5446);
xor U14474 (N_14474,N_9264,N_6979);
or U14475 (N_14475,N_6956,N_1110);
and U14476 (N_14476,N_3180,N_292);
nand U14477 (N_14477,N_819,N_7722);
xor U14478 (N_14478,N_6441,N_242);
and U14479 (N_14479,N_6970,N_9836);
xnor U14480 (N_14480,N_3964,N_3464);
or U14481 (N_14481,N_4441,N_1649);
nand U14482 (N_14482,N_4514,N_3478);
and U14483 (N_14483,N_7600,N_5466);
nor U14484 (N_14484,N_7779,N_4708);
xor U14485 (N_14485,N_7478,N_1729);
nor U14486 (N_14486,N_5703,N_1652);
nand U14487 (N_14487,N_3589,N_1953);
nor U14488 (N_14488,N_2500,N_5016);
xnor U14489 (N_14489,N_4815,N_7544);
nand U14490 (N_14490,N_1909,N_3845);
or U14491 (N_14491,N_3213,N_2594);
and U14492 (N_14492,N_1663,N_4743);
xnor U14493 (N_14493,N_139,N_4706);
or U14494 (N_14494,N_8529,N_2887);
and U14495 (N_14495,N_6717,N_6463);
xor U14496 (N_14496,N_9681,N_1274);
nand U14497 (N_14497,N_118,N_8795);
nor U14498 (N_14498,N_565,N_3788);
nand U14499 (N_14499,N_8378,N_4069);
nand U14500 (N_14500,N_367,N_3533);
and U14501 (N_14501,N_6935,N_8366);
and U14502 (N_14502,N_4488,N_3935);
and U14503 (N_14503,N_1184,N_2941);
xnor U14504 (N_14504,N_2452,N_1536);
nand U14505 (N_14505,N_8289,N_2648);
xor U14506 (N_14506,N_3929,N_979);
xnor U14507 (N_14507,N_5432,N_4009);
and U14508 (N_14508,N_8265,N_67);
xnor U14509 (N_14509,N_6957,N_5679);
nor U14510 (N_14510,N_4653,N_524);
or U14511 (N_14511,N_9157,N_9037);
or U14512 (N_14512,N_7627,N_3772);
or U14513 (N_14513,N_4034,N_2686);
and U14514 (N_14514,N_1877,N_2734);
nand U14515 (N_14515,N_4006,N_3627);
nand U14516 (N_14516,N_8443,N_4438);
nor U14517 (N_14517,N_8916,N_600);
nor U14518 (N_14518,N_9908,N_5080);
nor U14519 (N_14519,N_9583,N_9763);
nor U14520 (N_14520,N_3518,N_9806);
nor U14521 (N_14521,N_1215,N_4506);
and U14522 (N_14522,N_4585,N_8212);
nand U14523 (N_14523,N_6961,N_7566);
or U14524 (N_14524,N_7321,N_9040);
and U14525 (N_14525,N_4602,N_3927);
or U14526 (N_14526,N_3588,N_8314);
nor U14527 (N_14527,N_5021,N_787);
or U14528 (N_14528,N_3909,N_4636);
nand U14529 (N_14529,N_1814,N_5644);
nand U14530 (N_14530,N_4115,N_15);
nor U14531 (N_14531,N_7706,N_6469);
nor U14532 (N_14532,N_9961,N_6779);
and U14533 (N_14533,N_7877,N_2162);
or U14534 (N_14534,N_6027,N_8555);
nor U14535 (N_14535,N_5048,N_2144);
or U14536 (N_14536,N_1020,N_5395);
and U14537 (N_14537,N_5776,N_4938);
xor U14538 (N_14538,N_8174,N_8179);
xor U14539 (N_14539,N_2951,N_83);
nor U14540 (N_14540,N_2524,N_6093);
or U14541 (N_14541,N_4201,N_7717);
nand U14542 (N_14542,N_455,N_1638);
and U14543 (N_14543,N_689,N_5863);
nand U14544 (N_14544,N_3669,N_6124);
xor U14545 (N_14545,N_7175,N_397);
nor U14546 (N_14546,N_6040,N_239);
and U14547 (N_14547,N_36,N_210);
nand U14548 (N_14548,N_2442,N_107);
xor U14549 (N_14549,N_9909,N_1567);
and U14550 (N_14550,N_970,N_9862);
and U14551 (N_14551,N_6755,N_7390);
nand U14552 (N_14552,N_1013,N_7597);
or U14553 (N_14553,N_2170,N_6467);
xnor U14554 (N_14554,N_7925,N_4143);
nand U14555 (N_14555,N_7016,N_9655);
nor U14556 (N_14556,N_8500,N_9725);
xor U14557 (N_14557,N_2840,N_2441);
xnor U14558 (N_14558,N_5145,N_7747);
xor U14559 (N_14559,N_1231,N_5173);
or U14560 (N_14560,N_7204,N_5056);
or U14561 (N_14561,N_1195,N_137);
xor U14562 (N_14562,N_8852,N_5099);
nand U14563 (N_14563,N_1644,N_5206);
or U14564 (N_14564,N_6088,N_9477);
xnor U14565 (N_14565,N_1554,N_5185);
nand U14566 (N_14566,N_9258,N_9990);
xor U14567 (N_14567,N_6634,N_6563);
or U14568 (N_14568,N_250,N_6248);
or U14569 (N_14569,N_5344,N_892);
nor U14570 (N_14570,N_7395,N_111);
or U14571 (N_14571,N_2488,N_7165);
or U14572 (N_14572,N_2384,N_1739);
nand U14573 (N_14573,N_3053,N_1986);
or U14574 (N_14574,N_1172,N_8888);
xor U14575 (N_14575,N_7118,N_8906);
or U14576 (N_14576,N_5135,N_5687);
and U14577 (N_14577,N_5024,N_2468);
or U14578 (N_14578,N_5918,N_1494);
nand U14579 (N_14579,N_9115,N_8544);
nand U14580 (N_14580,N_3896,N_4537);
xnor U14581 (N_14581,N_4673,N_324);
xor U14582 (N_14582,N_6145,N_4837);
nor U14583 (N_14583,N_9019,N_9739);
or U14584 (N_14584,N_5523,N_1411);
nand U14585 (N_14585,N_3670,N_7665);
or U14586 (N_14586,N_8702,N_249);
nand U14587 (N_14587,N_3549,N_2033);
nor U14588 (N_14588,N_2635,N_9505);
nand U14589 (N_14589,N_6950,N_9595);
or U14590 (N_14590,N_9937,N_1010);
xor U14591 (N_14591,N_8585,N_7345);
nor U14592 (N_14592,N_7457,N_1345);
nor U14593 (N_14593,N_8877,N_4123);
or U14594 (N_14594,N_4096,N_4687);
nor U14595 (N_14595,N_8974,N_1918);
xor U14596 (N_14596,N_9177,N_601);
nand U14597 (N_14597,N_4563,N_9852);
or U14598 (N_14598,N_5869,N_3729);
nor U14599 (N_14599,N_7183,N_6537);
xnor U14600 (N_14600,N_3621,N_9167);
and U14601 (N_14601,N_4788,N_2388);
nor U14602 (N_14602,N_3486,N_2438);
and U14603 (N_14603,N_6427,N_4525);
and U14604 (N_14604,N_1036,N_8740);
nand U14605 (N_14605,N_2913,N_1282);
xor U14606 (N_14606,N_4864,N_8183);
or U14607 (N_14607,N_3176,N_841);
and U14608 (N_14608,N_6752,N_2184);
nor U14609 (N_14609,N_5078,N_4652);
and U14610 (N_14610,N_7019,N_755);
nor U14611 (N_14611,N_9134,N_1965);
nor U14612 (N_14612,N_7207,N_8497);
xnor U14613 (N_14613,N_4230,N_6232);
nand U14614 (N_14614,N_660,N_5222);
xnor U14615 (N_14615,N_7729,N_4114);
or U14616 (N_14616,N_2979,N_9792);
or U14617 (N_14617,N_7296,N_8843);
nor U14618 (N_14618,N_2727,N_4521);
or U14619 (N_14619,N_4671,N_3961);
nand U14620 (N_14620,N_9154,N_8813);
xnor U14621 (N_14621,N_4073,N_8110);
or U14622 (N_14622,N_7589,N_4353);
nand U14623 (N_14623,N_2756,N_5195);
xnor U14624 (N_14624,N_6820,N_6786);
xnor U14625 (N_14625,N_6101,N_1812);
or U14626 (N_14626,N_3656,N_6362);
nor U14627 (N_14627,N_2375,N_124);
nand U14628 (N_14628,N_4982,N_5731);
nor U14629 (N_14629,N_7203,N_2027);
nor U14630 (N_14630,N_2576,N_6877);
nor U14631 (N_14631,N_6854,N_9219);
or U14632 (N_14632,N_4110,N_5281);
or U14633 (N_14633,N_5946,N_575);
nand U14634 (N_14634,N_2264,N_5814);
or U14635 (N_14635,N_8936,N_3780);
nand U14636 (N_14636,N_138,N_1212);
or U14637 (N_14637,N_2029,N_2322);
or U14638 (N_14638,N_5150,N_6949);
nor U14639 (N_14639,N_7237,N_2239);
nor U14640 (N_14640,N_60,N_271);
nor U14641 (N_14641,N_7549,N_2238);
nor U14642 (N_14642,N_8819,N_4031);
and U14643 (N_14643,N_7475,N_9624);
and U14644 (N_14644,N_6769,N_4171);
and U14645 (N_14645,N_5458,N_5331);
nand U14646 (N_14646,N_4296,N_7235);
or U14647 (N_14647,N_297,N_5750);
nor U14648 (N_14648,N_264,N_9503);
nand U14649 (N_14649,N_6695,N_8038);
and U14650 (N_14650,N_7178,N_4908);
nor U14651 (N_14651,N_4798,N_5711);
nand U14652 (N_14652,N_3707,N_2054);
nand U14653 (N_14653,N_8227,N_8551);
xnor U14654 (N_14654,N_3694,N_4005);
nand U14655 (N_14655,N_926,N_7276);
and U14656 (N_14656,N_9563,N_117);
or U14657 (N_14657,N_863,N_6103);
or U14658 (N_14658,N_2681,N_3421);
nand U14659 (N_14659,N_1766,N_3200);
and U14660 (N_14660,N_967,N_9970);
nor U14661 (N_14661,N_2689,N_2242);
xor U14662 (N_14662,N_1995,N_3364);
and U14663 (N_14663,N_1553,N_6055);
or U14664 (N_14664,N_8448,N_7336);
and U14665 (N_14665,N_821,N_9298);
nor U14666 (N_14666,N_2246,N_6794);
and U14667 (N_14667,N_6808,N_4740);
nand U14668 (N_14668,N_7814,N_5360);
xor U14669 (N_14669,N_6138,N_323);
nand U14670 (N_14670,N_3817,N_6978);
or U14671 (N_14671,N_7349,N_495);
and U14672 (N_14672,N_5558,N_6551);
or U14673 (N_14673,N_1901,N_4321);
nand U14674 (N_14674,N_4909,N_687);
nor U14675 (N_14675,N_9292,N_9398);
and U14676 (N_14676,N_2358,N_5058);
and U14677 (N_14677,N_9278,N_3906);
and U14678 (N_14678,N_1870,N_3197);
nand U14679 (N_14679,N_8952,N_9566);
nor U14680 (N_14680,N_7470,N_9589);
and U14681 (N_14681,N_9135,N_4014);
nor U14682 (N_14682,N_9848,N_4883);
or U14683 (N_14683,N_2559,N_3977);
or U14684 (N_14684,N_6829,N_4836);
xnor U14685 (N_14685,N_7540,N_2048);
nand U14686 (N_14686,N_4133,N_1985);
or U14687 (N_14687,N_2638,N_5182);
or U14688 (N_14688,N_1899,N_731);
or U14689 (N_14689,N_7618,N_379);
or U14690 (N_14690,N_2145,N_3723);
nor U14691 (N_14691,N_3324,N_6393);
or U14692 (N_14692,N_7682,N_5601);
nand U14693 (N_14693,N_690,N_6383);
xnor U14694 (N_14694,N_4389,N_637);
and U14695 (N_14695,N_3632,N_5398);
xor U14696 (N_14696,N_7997,N_236);
or U14697 (N_14697,N_7394,N_1060);
nand U14698 (N_14698,N_5642,N_4385);
and U14699 (N_14699,N_2179,N_9708);
nand U14700 (N_14700,N_9438,N_1595);
nor U14701 (N_14701,N_8876,N_1853);
and U14702 (N_14702,N_6847,N_6587);
nor U14703 (N_14703,N_6982,N_4944);
nor U14704 (N_14704,N_3948,N_1560);
or U14705 (N_14705,N_5785,N_6539);
and U14706 (N_14706,N_4713,N_1890);
xor U14707 (N_14707,N_4863,N_1284);
nand U14708 (N_14708,N_4167,N_2796);
or U14709 (N_14709,N_1977,N_7534);
or U14710 (N_14710,N_7942,N_178);
nor U14711 (N_14711,N_7859,N_5283);
nand U14712 (N_14712,N_3286,N_7220);
xor U14713 (N_14713,N_8133,N_9569);
xnor U14714 (N_14714,N_8200,N_2829);
or U14715 (N_14715,N_3972,N_1869);
nand U14716 (N_14716,N_9374,N_523);
xnor U14717 (N_14717,N_6958,N_5269);
nor U14718 (N_14718,N_5291,N_6655);
nand U14719 (N_14719,N_5825,N_9727);
nor U14720 (N_14720,N_2289,N_4718);
xor U14721 (N_14721,N_6261,N_1830);
nand U14722 (N_14722,N_6610,N_5512);
nor U14723 (N_14723,N_6525,N_2835);
xnor U14724 (N_14724,N_4311,N_3790);
xnor U14725 (N_14725,N_9389,N_9535);
or U14726 (N_14726,N_2995,N_6567);
or U14727 (N_14727,N_8864,N_2747);
and U14728 (N_14728,N_8098,N_9187);
and U14729 (N_14729,N_4292,N_1124);
and U14730 (N_14730,N_6639,N_7331);
nor U14731 (N_14731,N_1632,N_4634);
nor U14732 (N_14732,N_5226,N_5380);
nor U14733 (N_14733,N_6366,N_808);
nand U14734 (N_14734,N_8409,N_180);
or U14735 (N_14735,N_7684,N_5563);
nor U14736 (N_14736,N_4813,N_9750);
nor U14737 (N_14737,N_3529,N_5811);
or U14738 (N_14738,N_5666,N_1374);
and U14739 (N_14739,N_5082,N_1033);
xor U14740 (N_14740,N_1628,N_5633);
nand U14741 (N_14741,N_4463,N_6116);
and U14742 (N_14742,N_2795,N_3559);
nor U14743 (N_14743,N_4338,N_2705);
or U14744 (N_14744,N_326,N_332);
or U14745 (N_14745,N_4113,N_5655);
xnor U14746 (N_14746,N_7281,N_2496);
xor U14747 (N_14747,N_9573,N_588);
nand U14748 (N_14748,N_196,N_5169);
xor U14749 (N_14749,N_7765,N_5273);
nor U14750 (N_14750,N_7014,N_3792);
nor U14751 (N_14751,N_4635,N_3567);
or U14752 (N_14752,N_1951,N_5073);
xor U14753 (N_14753,N_5261,N_9499);
xnor U14754 (N_14754,N_2674,N_6837);
and U14755 (N_14755,N_6699,N_1914);
nor U14756 (N_14756,N_1495,N_3146);
xnor U14757 (N_14757,N_2514,N_1518);
or U14758 (N_14758,N_6841,N_5742);
xor U14759 (N_14759,N_9251,N_3798);
nand U14760 (N_14760,N_3266,N_1461);
and U14761 (N_14761,N_2502,N_2308);
or U14762 (N_14762,N_1606,N_6579);
nor U14763 (N_14763,N_3800,N_7071);
nor U14764 (N_14764,N_3483,N_1711);
xor U14765 (N_14765,N_3564,N_7871);
nor U14766 (N_14766,N_7056,N_7775);
nand U14767 (N_14767,N_5759,N_5160);
xnor U14768 (N_14768,N_4220,N_9721);
xor U14769 (N_14769,N_3988,N_2642);
nor U14770 (N_14770,N_5375,N_469);
and U14771 (N_14771,N_9277,N_7572);
nor U14772 (N_14772,N_8830,N_3911);
and U14773 (N_14773,N_1955,N_985);
xnor U14774 (N_14774,N_8757,N_3261);
and U14775 (N_14775,N_2232,N_5876);
or U14776 (N_14776,N_3653,N_4265);
nand U14777 (N_14777,N_5209,N_5098);
nor U14778 (N_14778,N_4423,N_3510);
xnor U14779 (N_14779,N_7971,N_3283);
or U14780 (N_14780,N_8605,N_659);
and U14781 (N_14781,N_8594,N_4450);
xor U14782 (N_14782,N_8642,N_7189);
or U14783 (N_14783,N_7647,N_3149);
and U14784 (N_14784,N_858,N_2396);
or U14785 (N_14785,N_5693,N_1346);
nor U14786 (N_14786,N_8029,N_5537);
nor U14787 (N_14787,N_9529,N_5628);
and U14788 (N_14788,N_3301,N_5232);
nand U14789 (N_14789,N_6692,N_4969);
nor U14790 (N_14790,N_8609,N_9041);
or U14791 (N_14791,N_4852,N_896);
or U14792 (N_14792,N_2818,N_8214);
or U14793 (N_14793,N_9055,N_8721);
xor U14794 (N_14794,N_3545,N_8267);
nor U14795 (N_14795,N_3625,N_4666);
and U14796 (N_14796,N_2171,N_512);
nor U14797 (N_14797,N_6192,N_3541);
nand U14798 (N_14798,N_5384,N_294);
or U14799 (N_14799,N_811,N_2443);
xnor U14800 (N_14800,N_461,N_1605);
xnor U14801 (N_14801,N_8701,N_9413);
nand U14802 (N_14802,N_4495,N_6228);
and U14803 (N_14803,N_9875,N_6391);
nand U14804 (N_14804,N_7867,N_6530);
nand U14805 (N_14805,N_864,N_2078);
nor U14806 (N_14806,N_3308,N_6188);
xor U14807 (N_14807,N_4348,N_2434);
and U14808 (N_14808,N_8001,N_4107);
nor U14809 (N_14809,N_7919,N_7197);
or U14810 (N_14810,N_5121,N_9903);
xor U14811 (N_14811,N_8352,N_4714);
nand U14812 (N_14812,N_2343,N_8104);
nor U14813 (N_14813,N_5477,N_5412);
and U14814 (N_14814,N_8944,N_3454);
or U14815 (N_14815,N_4166,N_7297);
or U14816 (N_14816,N_7528,N_9926);
and U14817 (N_14817,N_6549,N_7469);
nor U14818 (N_14818,N_2243,N_6593);
or U14819 (N_14819,N_5977,N_9237);
xnor U14820 (N_14820,N_3640,N_918);
xor U14821 (N_14821,N_3647,N_4257);
nor U14822 (N_14822,N_5670,N_9043);
or U14823 (N_14823,N_9118,N_9400);
or U14824 (N_14824,N_7141,N_8836);
xnor U14825 (N_14825,N_3818,N_8464);
nor U14826 (N_14826,N_3805,N_9330);
nand U14827 (N_14827,N_8142,N_876);
and U14828 (N_14828,N_3973,N_2087);
nor U14829 (N_14829,N_3616,N_5154);
and U14830 (N_14830,N_1816,N_3608);
or U14831 (N_14831,N_3642,N_963);
or U14832 (N_14832,N_8759,N_6165);
nor U14833 (N_14833,N_6848,N_5453);
and U14834 (N_14834,N_8373,N_2633);
nor U14835 (N_14835,N_3968,N_8400);
nor U14836 (N_14836,N_8015,N_6420);
xnor U14837 (N_14837,N_7063,N_9669);
or U14838 (N_14838,N_5377,N_8948);
nand U14839 (N_14839,N_6839,N_7724);
nor U14840 (N_14840,N_8922,N_1817);
and U14841 (N_14841,N_7142,N_7364);
nor U14842 (N_14842,N_9396,N_6195);
nand U14843 (N_14843,N_3148,N_2188);
or U14844 (N_14844,N_3039,N_6976);
nand U14845 (N_14845,N_8980,N_546);
nand U14846 (N_14846,N_7380,N_1921);
nor U14847 (N_14847,N_7833,N_8128);
nor U14848 (N_14848,N_3602,N_8388);
or U14849 (N_14849,N_1009,N_2664);
nand U14850 (N_14850,N_1441,N_8419);
nor U14851 (N_14851,N_458,N_8389);
xor U14852 (N_14852,N_3581,N_2509);
and U14853 (N_14853,N_3026,N_5152);
nand U14854 (N_14854,N_7948,N_2479);
nand U14855 (N_14855,N_1849,N_6037);
xnor U14856 (N_14856,N_7632,N_5694);
xnor U14857 (N_14857,N_9452,N_6347);
nand U14858 (N_14858,N_9604,N_5669);
nand U14859 (N_14859,N_8385,N_3436);
xnor U14860 (N_14860,N_9785,N_4679);
or U14861 (N_14861,N_6654,N_401);
nor U14862 (N_14862,N_5243,N_1506);
and U14863 (N_14863,N_2564,N_4289);
nand U14864 (N_14864,N_4327,N_3513);
nor U14865 (N_14865,N_3639,N_5753);
nand U14866 (N_14866,N_7431,N_2295);
xor U14867 (N_14867,N_7009,N_7440);
nor U14868 (N_14868,N_568,N_1138);
nor U14869 (N_14869,N_6434,N_7215);
xnor U14870 (N_14870,N_1254,N_1330);
xnor U14871 (N_14871,N_2873,N_6853);
and U14872 (N_14872,N_7843,N_2433);
or U14873 (N_14873,N_6677,N_7594);
nand U14874 (N_14874,N_5787,N_7869);
nand U14875 (N_14875,N_8764,N_2965);
or U14876 (N_14876,N_2863,N_3430);
nand U14877 (N_14877,N_2317,N_703);
or U14878 (N_14878,N_734,N_3008);
and U14879 (N_14879,N_3082,N_8644);
or U14880 (N_14880,N_6602,N_6870);
and U14881 (N_14881,N_9849,N_3502);
or U14882 (N_14882,N_2098,N_7766);
or U14883 (N_14883,N_8134,N_3849);
and U14884 (N_14884,N_7082,N_6168);
nand U14885 (N_14885,N_2499,N_6743);
nor U14886 (N_14886,N_1423,N_1679);
nor U14887 (N_14887,N_5535,N_2507);
and U14888 (N_14888,N_4663,N_6813);
nand U14889 (N_14889,N_5723,N_5552);
nand U14890 (N_14890,N_6069,N_8333);
nand U14891 (N_14891,N_2336,N_3684);
and U14892 (N_14892,N_8082,N_8925);
xnor U14893 (N_14893,N_7892,N_1763);
nor U14894 (N_14894,N_5877,N_4099);
and U14895 (N_14895,N_7772,N_7985);
or U14896 (N_14896,N_3807,N_7561);
nand U14897 (N_14897,N_4603,N_1069);
nand U14898 (N_14898,N_3526,N_2665);
nor U14899 (N_14899,N_2167,N_762);
xor U14900 (N_14900,N_6687,N_4440);
nand U14901 (N_14901,N_9076,N_3168);
nand U14902 (N_14902,N_2856,N_1273);
or U14903 (N_14903,N_6073,N_6317);
nand U14904 (N_14904,N_3210,N_1479);
nand U14905 (N_14905,N_3295,N_8275);
or U14906 (N_14906,N_5109,N_1478);
nand U14907 (N_14907,N_2311,N_1388);
xnor U14908 (N_14908,N_7400,N_5899);
xor U14909 (N_14909,N_977,N_162);
nand U14910 (N_14910,N_3607,N_6297);
or U14911 (N_14911,N_916,N_4049);
nor U14912 (N_14912,N_7635,N_2977);
nor U14913 (N_14913,N_5822,N_7810);
or U14914 (N_14914,N_5423,N_8964);
xnor U14915 (N_14915,N_1467,N_1104);
xnor U14916 (N_14916,N_9144,N_641);
nor U14917 (N_14917,N_2808,N_1658);
nand U14918 (N_14918,N_4914,N_251);
nand U14919 (N_14919,N_3284,N_9350);
xor U14920 (N_14920,N_4207,N_9461);
nand U14921 (N_14921,N_4012,N_3035);
xor U14922 (N_14922,N_3887,N_6308);
nor U14923 (N_14923,N_7640,N_9473);
or U14924 (N_14924,N_2739,N_1443);
xor U14925 (N_14925,N_183,N_900);
and U14926 (N_14926,N_17,N_1154);
xnor U14927 (N_14927,N_7522,N_5982);
and U14928 (N_14928,N_1568,N_3682);
or U14929 (N_14929,N_6529,N_426);
nand U14930 (N_14930,N_3419,N_2275);
or U14931 (N_14931,N_1751,N_8928);
nand U14932 (N_14932,N_6071,N_2837);
and U14933 (N_14933,N_3535,N_6862);
or U14934 (N_14934,N_291,N_1470);
and U14935 (N_14935,N_7422,N_2999);
nand U14936 (N_14936,N_826,N_2189);
nor U14937 (N_14937,N_8869,N_4029);
xnor U14938 (N_14938,N_5507,N_5052);
nand U14939 (N_14939,N_1466,N_4215);
or U14940 (N_14940,N_2562,N_7593);
or U14941 (N_14941,N_9951,N_1792);
or U14942 (N_14942,N_9658,N_3876);
xor U14943 (N_14943,N_212,N_8958);
nand U14944 (N_14944,N_4882,N_9942);
xor U14945 (N_14945,N_5393,N_1543);
nor U14946 (N_14946,N_2715,N_850);
xnor U14947 (N_14947,N_2817,N_706);
or U14948 (N_14948,N_161,N_2542);
xnor U14949 (N_14949,N_2538,N_4793);
xnor U14950 (N_14950,N_3762,N_4095);
or U14951 (N_14951,N_1895,N_4543);
nor U14952 (N_14952,N_4368,N_3117);
nor U14953 (N_14953,N_870,N_7986);
nor U14954 (N_14954,N_8507,N_4249);
or U14955 (N_14955,N_931,N_9864);
nand U14956 (N_14956,N_9360,N_7164);
nand U14957 (N_14957,N_5959,N_6096);
and U14958 (N_14958,N_3359,N_3689);
xnor U14959 (N_14959,N_820,N_2414);
and U14960 (N_14960,N_6119,N_7046);
nand U14961 (N_14961,N_2932,N_1811);
or U14962 (N_14962,N_2371,N_4072);
and U14963 (N_14963,N_5067,N_5069);
nand U14964 (N_14964,N_4560,N_5936);
nand U14965 (N_14965,N_3879,N_3980);
and U14966 (N_14966,N_8391,N_4414);
nor U14967 (N_14967,N_9904,N_3517);
or U14968 (N_14968,N_6657,N_9745);
nor U14969 (N_14969,N_5831,N_1708);
xor U14970 (N_14970,N_2811,N_1119);
nand U14971 (N_14971,N_1549,N_1128);
xor U14972 (N_14972,N_3005,N_3015);
and U14973 (N_14973,N_8921,N_5187);
xor U14974 (N_14974,N_7260,N_7104);
xnor U14975 (N_14975,N_6472,N_8556);
nor U14976 (N_14976,N_2593,N_9263);
or U14977 (N_14977,N_1776,N_7476);
nor U14978 (N_14978,N_6500,N_8219);
xnor U14979 (N_14979,N_3098,N_1144);
or U14980 (N_14980,N_3136,N_8252);
nor U14981 (N_14981,N_4727,N_507);
or U14982 (N_14982,N_4819,N_3229);
or U14983 (N_14983,N_6975,N_6453);
nor U14984 (N_14984,N_9738,N_8254);
nand U14985 (N_14985,N_1426,N_3441);
or U14986 (N_14986,N_2004,N_5275);
nand U14987 (N_14987,N_8360,N_3352);
or U14988 (N_14988,N_7150,N_2565);
xnor U14989 (N_14989,N_5894,N_7066);
or U14990 (N_14990,N_4420,N_6034);
nand U14991 (N_14991,N_5220,N_8346);
nand U14992 (N_14992,N_2790,N_5984);
nand U14993 (N_14993,N_3508,N_4179);
or U14994 (N_14994,N_5460,N_9236);
nand U14995 (N_14995,N_57,N_4154);
and U14996 (N_14996,N_5596,N_6010);
xnor U14997 (N_14997,N_7567,N_8586);
nor U14998 (N_14998,N_657,N_8659);
and U14999 (N_14999,N_8264,N_9540);
and U15000 (N_15000,N_5380,N_8105);
or U15001 (N_15001,N_8655,N_8508);
and U15002 (N_15002,N_2875,N_2474);
xor U15003 (N_15003,N_2000,N_9419);
xnor U15004 (N_15004,N_5923,N_6589);
xor U15005 (N_15005,N_1213,N_2054);
xor U15006 (N_15006,N_9629,N_3139);
and U15007 (N_15007,N_7541,N_1714);
or U15008 (N_15008,N_4396,N_3159);
or U15009 (N_15009,N_1822,N_5098);
nand U15010 (N_15010,N_1332,N_9693);
or U15011 (N_15011,N_5230,N_6564);
xor U15012 (N_15012,N_1517,N_5039);
and U15013 (N_15013,N_5913,N_3846);
and U15014 (N_15014,N_2337,N_7217);
nand U15015 (N_15015,N_6826,N_7508);
or U15016 (N_15016,N_7785,N_7852);
or U15017 (N_15017,N_2632,N_3801);
xnor U15018 (N_15018,N_5025,N_7328);
xor U15019 (N_15019,N_8301,N_5969);
xnor U15020 (N_15020,N_3605,N_8283);
and U15021 (N_15021,N_1594,N_7308);
nand U15022 (N_15022,N_2063,N_3092);
and U15023 (N_15023,N_9706,N_8118);
nand U15024 (N_15024,N_309,N_7163);
nand U15025 (N_15025,N_4728,N_1510);
nand U15026 (N_15026,N_3056,N_481);
nor U15027 (N_15027,N_6181,N_4570);
and U15028 (N_15028,N_2396,N_6564);
or U15029 (N_15029,N_4005,N_9607);
nand U15030 (N_15030,N_1964,N_53);
and U15031 (N_15031,N_7299,N_3555);
nand U15032 (N_15032,N_821,N_1492);
or U15033 (N_15033,N_4695,N_2339);
xor U15034 (N_15034,N_8388,N_2590);
nor U15035 (N_15035,N_8864,N_770);
and U15036 (N_15036,N_7254,N_8902);
xor U15037 (N_15037,N_6103,N_6320);
xnor U15038 (N_15038,N_3008,N_2830);
nor U15039 (N_15039,N_8193,N_9333);
and U15040 (N_15040,N_4155,N_2997);
nor U15041 (N_15041,N_6131,N_7644);
xor U15042 (N_15042,N_6077,N_8371);
or U15043 (N_15043,N_539,N_3419);
xnor U15044 (N_15044,N_3049,N_5729);
xor U15045 (N_15045,N_4982,N_9320);
xor U15046 (N_15046,N_8747,N_5765);
nand U15047 (N_15047,N_7584,N_7972);
nand U15048 (N_15048,N_1563,N_4440);
nor U15049 (N_15049,N_7060,N_4163);
or U15050 (N_15050,N_9802,N_8238);
or U15051 (N_15051,N_6985,N_3897);
and U15052 (N_15052,N_1315,N_7731);
or U15053 (N_15053,N_505,N_8872);
xor U15054 (N_15054,N_5364,N_9657);
xnor U15055 (N_15055,N_9414,N_8955);
xor U15056 (N_15056,N_1563,N_3259);
nand U15057 (N_15057,N_1879,N_6847);
or U15058 (N_15058,N_3744,N_2596);
nor U15059 (N_15059,N_8350,N_5717);
nor U15060 (N_15060,N_7080,N_5953);
nor U15061 (N_15061,N_3004,N_5217);
nand U15062 (N_15062,N_1981,N_1098);
nor U15063 (N_15063,N_5877,N_3147);
xnor U15064 (N_15064,N_1638,N_4238);
nand U15065 (N_15065,N_2941,N_2552);
nor U15066 (N_15066,N_8325,N_3404);
and U15067 (N_15067,N_8101,N_2689);
or U15068 (N_15068,N_5514,N_795);
nor U15069 (N_15069,N_1483,N_4844);
nor U15070 (N_15070,N_7287,N_6977);
and U15071 (N_15071,N_5229,N_6376);
nand U15072 (N_15072,N_7766,N_8196);
or U15073 (N_15073,N_4866,N_548);
nor U15074 (N_15074,N_1345,N_94);
xnor U15075 (N_15075,N_9997,N_3466);
and U15076 (N_15076,N_2471,N_5210);
nand U15077 (N_15077,N_4962,N_1698);
nand U15078 (N_15078,N_5682,N_5150);
or U15079 (N_15079,N_4083,N_6101);
nor U15080 (N_15080,N_5175,N_5007);
nor U15081 (N_15081,N_9552,N_2279);
xnor U15082 (N_15082,N_4722,N_6457);
and U15083 (N_15083,N_6132,N_7875);
and U15084 (N_15084,N_9116,N_6435);
xnor U15085 (N_15085,N_3854,N_3293);
xor U15086 (N_15086,N_7102,N_7570);
or U15087 (N_15087,N_9267,N_2317);
and U15088 (N_15088,N_44,N_3480);
xor U15089 (N_15089,N_5502,N_6816);
nand U15090 (N_15090,N_7699,N_4058);
nor U15091 (N_15091,N_8587,N_5440);
nand U15092 (N_15092,N_3327,N_7597);
nor U15093 (N_15093,N_4480,N_9729);
or U15094 (N_15094,N_7738,N_5504);
xor U15095 (N_15095,N_5675,N_2591);
nor U15096 (N_15096,N_4172,N_7094);
nor U15097 (N_15097,N_3820,N_6547);
nor U15098 (N_15098,N_8174,N_2684);
nand U15099 (N_15099,N_2606,N_5536);
nor U15100 (N_15100,N_5914,N_9508);
and U15101 (N_15101,N_9757,N_4002);
and U15102 (N_15102,N_8534,N_4542);
nand U15103 (N_15103,N_9613,N_6345);
xor U15104 (N_15104,N_7787,N_6139);
xnor U15105 (N_15105,N_4037,N_3750);
nand U15106 (N_15106,N_9816,N_9326);
nor U15107 (N_15107,N_3659,N_727);
and U15108 (N_15108,N_960,N_72);
xnor U15109 (N_15109,N_3867,N_7409);
and U15110 (N_15110,N_2851,N_6369);
and U15111 (N_15111,N_694,N_3522);
nand U15112 (N_15112,N_7993,N_5392);
and U15113 (N_15113,N_1960,N_1332);
nor U15114 (N_15114,N_9601,N_7597);
nand U15115 (N_15115,N_234,N_1130);
or U15116 (N_15116,N_1182,N_9706);
xor U15117 (N_15117,N_7772,N_292);
or U15118 (N_15118,N_6959,N_3011);
xnor U15119 (N_15119,N_5121,N_7488);
nand U15120 (N_15120,N_98,N_5617);
and U15121 (N_15121,N_4008,N_1255);
or U15122 (N_15122,N_1470,N_5932);
xnor U15123 (N_15123,N_1634,N_4789);
xor U15124 (N_15124,N_4417,N_5869);
nand U15125 (N_15125,N_9006,N_2598);
nor U15126 (N_15126,N_1430,N_5105);
or U15127 (N_15127,N_558,N_6717);
or U15128 (N_15128,N_8284,N_3531);
nand U15129 (N_15129,N_7171,N_5533);
and U15130 (N_15130,N_1335,N_3567);
nor U15131 (N_15131,N_5767,N_9734);
or U15132 (N_15132,N_237,N_9820);
and U15133 (N_15133,N_4552,N_8008);
and U15134 (N_15134,N_9305,N_6540);
or U15135 (N_15135,N_4491,N_241);
xor U15136 (N_15136,N_9471,N_8743);
xnor U15137 (N_15137,N_1284,N_5381);
or U15138 (N_15138,N_2279,N_1923);
nand U15139 (N_15139,N_7669,N_4018);
nor U15140 (N_15140,N_7827,N_8996);
nand U15141 (N_15141,N_3091,N_6757);
or U15142 (N_15142,N_9033,N_7791);
xor U15143 (N_15143,N_4530,N_5694);
and U15144 (N_15144,N_981,N_557);
and U15145 (N_15145,N_5535,N_5532);
nor U15146 (N_15146,N_1070,N_4786);
xnor U15147 (N_15147,N_2825,N_2547);
nor U15148 (N_15148,N_9399,N_4284);
and U15149 (N_15149,N_9890,N_8366);
and U15150 (N_15150,N_3828,N_5276);
and U15151 (N_15151,N_4182,N_1734);
nor U15152 (N_15152,N_6908,N_6148);
and U15153 (N_15153,N_1071,N_5629);
nor U15154 (N_15154,N_7700,N_6767);
nand U15155 (N_15155,N_598,N_1763);
or U15156 (N_15156,N_8178,N_4346);
and U15157 (N_15157,N_3042,N_340);
xor U15158 (N_15158,N_9709,N_4434);
xnor U15159 (N_15159,N_9479,N_6371);
nand U15160 (N_15160,N_1229,N_8767);
and U15161 (N_15161,N_3016,N_3172);
nand U15162 (N_15162,N_6740,N_2269);
xor U15163 (N_15163,N_6434,N_1004);
xnor U15164 (N_15164,N_175,N_8559);
nand U15165 (N_15165,N_6993,N_7081);
nand U15166 (N_15166,N_2855,N_164);
xor U15167 (N_15167,N_3674,N_8766);
nand U15168 (N_15168,N_7071,N_1266);
nand U15169 (N_15169,N_2838,N_164);
or U15170 (N_15170,N_5068,N_2612);
and U15171 (N_15171,N_3558,N_9382);
nor U15172 (N_15172,N_1080,N_8040);
nor U15173 (N_15173,N_7626,N_2167);
and U15174 (N_15174,N_149,N_7075);
nand U15175 (N_15175,N_6152,N_1774);
nor U15176 (N_15176,N_5762,N_7050);
and U15177 (N_15177,N_8734,N_800);
and U15178 (N_15178,N_7486,N_9396);
or U15179 (N_15179,N_3431,N_8605);
nand U15180 (N_15180,N_7986,N_830);
or U15181 (N_15181,N_7425,N_6814);
xnor U15182 (N_15182,N_1248,N_914);
nand U15183 (N_15183,N_2456,N_1473);
nand U15184 (N_15184,N_7093,N_4584);
and U15185 (N_15185,N_7957,N_1935);
and U15186 (N_15186,N_3319,N_6787);
or U15187 (N_15187,N_5857,N_8237);
xor U15188 (N_15188,N_7252,N_9434);
xor U15189 (N_15189,N_4152,N_7327);
and U15190 (N_15190,N_7502,N_3576);
and U15191 (N_15191,N_9314,N_2195);
nand U15192 (N_15192,N_3480,N_9424);
nand U15193 (N_15193,N_2045,N_1289);
xor U15194 (N_15194,N_6725,N_8948);
and U15195 (N_15195,N_9852,N_2466);
or U15196 (N_15196,N_7343,N_7952);
or U15197 (N_15197,N_1106,N_7980);
nor U15198 (N_15198,N_8637,N_9514);
nor U15199 (N_15199,N_9243,N_5883);
and U15200 (N_15200,N_5750,N_2622);
nand U15201 (N_15201,N_9835,N_16);
or U15202 (N_15202,N_6279,N_8263);
xor U15203 (N_15203,N_1016,N_8337);
and U15204 (N_15204,N_677,N_1229);
xnor U15205 (N_15205,N_6034,N_3095);
xor U15206 (N_15206,N_1379,N_7983);
and U15207 (N_15207,N_9847,N_6032);
and U15208 (N_15208,N_3618,N_8620);
xor U15209 (N_15209,N_4288,N_503);
xor U15210 (N_15210,N_4106,N_9752);
or U15211 (N_15211,N_3908,N_3370);
xnor U15212 (N_15212,N_5976,N_3075);
nor U15213 (N_15213,N_7950,N_2580);
xnor U15214 (N_15214,N_4941,N_3320);
nand U15215 (N_15215,N_3265,N_1434);
nand U15216 (N_15216,N_511,N_6374);
or U15217 (N_15217,N_8625,N_4121);
nand U15218 (N_15218,N_4916,N_7502);
and U15219 (N_15219,N_2164,N_5505);
xnor U15220 (N_15220,N_6081,N_5705);
and U15221 (N_15221,N_5709,N_4725);
or U15222 (N_15222,N_5131,N_7305);
and U15223 (N_15223,N_1287,N_2847);
and U15224 (N_15224,N_9445,N_8871);
and U15225 (N_15225,N_955,N_6141);
xnor U15226 (N_15226,N_8743,N_1299);
nand U15227 (N_15227,N_9721,N_3998);
or U15228 (N_15228,N_2373,N_1245);
or U15229 (N_15229,N_7767,N_7259);
nand U15230 (N_15230,N_8315,N_3843);
nand U15231 (N_15231,N_3507,N_3903);
xnor U15232 (N_15232,N_8031,N_1767);
xor U15233 (N_15233,N_1763,N_2944);
nand U15234 (N_15234,N_6041,N_7823);
or U15235 (N_15235,N_5967,N_3759);
nand U15236 (N_15236,N_9488,N_9769);
nand U15237 (N_15237,N_6375,N_3735);
nor U15238 (N_15238,N_1038,N_8757);
nor U15239 (N_15239,N_9932,N_7954);
and U15240 (N_15240,N_1650,N_8340);
xor U15241 (N_15241,N_7096,N_2071);
nand U15242 (N_15242,N_9140,N_343);
nor U15243 (N_15243,N_1540,N_6113);
and U15244 (N_15244,N_394,N_4641);
nand U15245 (N_15245,N_9181,N_3034);
xor U15246 (N_15246,N_9526,N_8118);
or U15247 (N_15247,N_975,N_7045);
nor U15248 (N_15248,N_7789,N_6921);
xor U15249 (N_15249,N_7177,N_8333);
xor U15250 (N_15250,N_3923,N_9475);
nor U15251 (N_15251,N_4021,N_7779);
nor U15252 (N_15252,N_7962,N_2420);
xnor U15253 (N_15253,N_5508,N_1033);
nor U15254 (N_15254,N_4481,N_255);
nand U15255 (N_15255,N_3959,N_1256);
nor U15256 (N_15256,N_1068,N_1938);
or U15257 (N_15257,N_9589,N_3701);
nand U15258 (N_15258,N_1814,N_710);
nor U15259 (N_15259,N_5687,N_3882);
xor U15260 (N_15260,N_9593,N_6370);
and U15261 (N_15261,N_4473,N_1822);
xor U15262 (N_15262,N_2620,N_5999);
or U15263 (N_15263,N_3433,N_4778);
or U15264 (N_15264,N_4981,N_6864);
nand U15265 (N_15265,N_9055,N_6785);
nand U15266 (N_15266,N_3424,N_4488);
or U15267 (N_15267,N_9418,N_1340);
or U15268 (N_15268,N_3338,N_518);
and U15269 (N_15269,N_3229,N_7634);
nor U15270 (N_15270,N_5299,N_8667);
nor U15271 (N_15271,N_5633,N_131);
or U15272 (N_15272,N_5586,N_8179);
or U15273 (N_15273,N_2457,N_4858);
xnor U15274 (N_15274,N_3135,N_8055);
xnor U15275 (N_15275,N_9901,N_2379);
nand U15276 (N_15276,N_4211,N_9081);
or U15277 (N_15277,N_2411,N_8581);
and U15278 (N_15278,N_4707,N_794);
and U15279 (N_15279,N_121,N_8905);
nor U15280 (N_15280,N_3682,N_3444);
and U15281 (N_15281,N_3148,N_7330);
and U15282 (N_15282,N_6946,N_5472);
or U15283 (N_15283,N_2621,N_912);
nand U15284 (N_15284,N_4232,N_5739);
nor U15285 (N_15285,N_772,N_5107);
xnor U15286 (N_15286,N_7638,N_1907);
nor U15287 (N_15287,N_1105,N_3895);
xor U15288 (N_15288,N_8313,N_8080);
and U15289 (N_15289,N_2865,N_4982);
nand U15290 (N_15290,N_4360,N_4087);
nor U15291 (N_15291,N_7038,N_62);
xnor U15292 (N_15292,N_8130,N_2550);
and U15293 (N_15293,N_9560,N_6191);
nand U15294 (N_15294,N_740,N_6379);
or U15295 (N_15295,N_4320,N_7367);
nor U15296 (N_15296,N_7778,N_7285);
nand U15297 (N_15297,N_3424,N_2730);
nand U15298 (N_15298,N_3533,N_2399);
or U15299 (N_15299,N_2095,N_8081);
xor U15300 (N_15300,N_2186,N_3218);
xor U15301 (N_15301,N_2920,N_5825);
or U15302 (N_15302,N_4792,N_7103);
nor U15303 (N_15303,N_6380,N_6797);
and U15304 (N_15304,N_8612,N_443);
or U15305 (N_15305,N_9742,N_8592);
nand U15306 (N_15306,N_7840,N_6508);
or U15307 (N_15307,N_2650,N_1217);
nor U15308 (N_15308,N_7874,N_2204);
xor U15309 (N_15309,N_1879,N_9262);
nor U15310 (N_15310,N_206,N_4962);
nand U15311 (N_15311,N_3276,N_3496);
xnor U15312 (N_15312,N_8758,N_7053);
or U15313 (N_15313,N_9935,N_4370);
nand U15314 (N_15314,N_8174,N_1633);
xor U15315 (N_15315,N_3773,N_4334);
xnor U15316 (N_15316,N_5770,N_8939);
nand U15317 (N_15317,N_4266,N_7773);
or U15318 (N_15318,N_6635,N_8547);
or U15319 (N_15319,N_1217,N_5335);
nor U15320 (N_15320,N_2271,N_7582);
or U15321 (N_15321,N_4679,N_2044);
nand U15322 (N_15322,N_1434,N_2891);
nand U15323 (N_15323,N_6780,N_8480);
or U15324 (N_15324,N_9195,N_9855);
xor U15325 (N_15325,N_1414,N_6911);
nor U15326 (N_15326,N_854,N_7573);
nand U15327 (N_15327,N_317,N_4539);
nor U15328 (N_15328,N_750,N_2590);
and U15329 (N_15329,N_8025,N_5603);
nor U15330 (N_15330,N_9868,N_6558);
nand U15331 (N_15331,N_7247,N_4788);
nor U15332 (N_15332,N_4363,N_8787);
xnor U15333 (N_15333,N_3677,N_1694);
nor U15334 (N_15334,N_463,N_7659);
or U15335 (N_15335,N_2643,N_9932);
nor U15336 (N_15336,N_6940,N_659);
and U15337 (N_15337,N_4882,N_7465);
or U15338 (N_15338,N_5406,N_2790);
xor U15339 (N_15339,N_5086,N_8386);
or U15340 (N_15340,N_5203,N_9189);
nand U15341 (N_15341,N_4100,N_8336);
or U15342 (N_15342,N_6637,N_3748);
nand U15343 (N_15343,N_2809,N_3685);
nor U15344 (N_15344,N_7441,N_1590);
xor U15345 (N_15345,N_5430,N_8054);
and U15346 (N_15346,N_5329,N_1295);
or U15347 (N_15347,N_22,N_8126);
xor U15348 (N_15348,N_1407,N_3129);
nand U15349 (N_15349,N_7079,N_3125);
and U15350 (N_15350,N_3395,N_1621);
or U15351 (N_15351,N_28,N_5756);
xor U15352 (N_15352,N_1271,N_9470);
nor U15353 (N_15353,N_649,N_3024);
nor U15354 (N_15354,N_7675,N_4453);
nor U15355 (N_15355,N_2114,N_8950);
and U15356 (N_15356,N_7683,N_8350);
and U15357 (N_15357,N_9649,N_9280);
or U15358 (N_15358,N_8323,N_4379);
nor U15359 (N_15359,N_2383,N_6245);
and U15360 (N_15360,N_9235,N_6090);
xor U15361 (N_15361,N_4739,N_2368);
and U15362 (N_15362,N_1906,N_9976);
xnor U15363 (N_15363,N_631,N_1991);
or U15364 (N_15364,N_1359,N_9963);
or U15365 (N_15365,N_8482,N_3771);
nand U15366 (N_15366,N_3560,N_5132);
and U15367 (N_15367,N_5071,N_3220);
nand U15368 (N_15368,N_4396,N_2274);
or U15369 (N_15369,N_5577,N_7773);
and U15370 (N_15370,N_4744,N_2122);
nand U15371 (N_15371,N_1996,N_8139);
or U15372 (N_15372,N_2754,N_2094);
or U15373 (N_15373,N_1170,N_5500);
and U15374 (N_15374,N_8007,N_709);
nand U15375 (N_15375,N_8430,N_703);
nand U15376 (N_15376,N_332,N_7444);
nand U15377 (N_15377,N_7338,N_5993);
xnor U15378 (N_15378,N_8093,N_1935);
and U15379 (N_15379,N_7519,N_4867);
xnor U15380 (N_15380,N_2085,N_950);
and U15381 (N_15381,N_1575,N_2526);
nand U15382 (N_15382,N_9095,N_4049);
or U15383 (N_15383,N_1825,N_4183);
xnor U15384 (N_15384,N_5022,N_2269);
nand U15385 (N_15385,N_7600,N_512);
or U15386 (N_15386,N_5929,N_2333);
xor U15387 (N_15387,N_8050,N_3382);
or U15388 (N_15388,N_3495,N_1192);
nor U15389 (N_15389,N_4980,N_9179);
or U15390 (N_15390,N_2179,N_4491);
xnor U15391 (N_15391,N_5416,N_8436);
xnor U15392 (N_15392,N_1488,N_6964);
nand U15393 (N_15393,N_7385,N_7255);
or U15394 (N_15394,N_8229,N_76);
and U15395 (N_15395,N_2472,N_6494);
nor U15396 (N_15396,N_2758,N_3124);
nand U15397 (N_15397,N_6278,N_9234);
nor U15398 (N_15398,N_9016,N_4909);
or U15399 (N_15399,N_8216,N_4690);
and U15400 (N_15400,N_3161,N_9550);
xor U15401 (N_15401,N_7255,N_4885);
and U15402 (N_15402,N_6533,N_4620);
xor U15403 (N_15403,N_2335,N_8731);
nor U15404 (N_15404,N_6148,N_6833);
or U15405 (N_15405,N_8694,N_3262);
and U15406 (N_15406,N_5678,N_116);
and U15407 (N_15407,N_2891,N_1785);
nand U15408 (N_15408,N_1495,N_2021);
nor U15409 (N_15409,N_4534,N_5777);
and U15410 (N_15410,N_7043,N_7131);
nor U15411 (N_15411,N_9472,N_3906);
nor U15412 (N_15412,N_4478,N_5976);
and U15413 (N_15413,N_4202,N_6757);
xnor U15414 (N_15414,N_6246,N_3661);
or U15415 (N_15415,N_3614,N_598);
and U15416 (N_15416,N_9123,N_3025);
nor U15417 (N_15417,N_9822,N_136);
xnor U15418 (N_15418,N_2580,N_8205);
nor U15419 (N_15419,N_8843,N_5670);
xnor U15420 (N_15420,N_4103,N_8233);
or U15421 (N_15421,N_8098,N_7120);
or U15422 (N_15422,N_4354,N_2987);
or U15423 (N_15423,N_3334,N_8892);
and U15424 (N_15424,N_7028,N_6804);
nand U15425 (N_15425,N_2002,N_4192);
or U15426 (N_15426,N_7462,N_6543);
or U15427 (N_15427,N_3579,N_9208);
nor U15428 (N_15428,N_5465,N_5263);
nor U15429 (N_15429,N_2554,N_4695);
nand U15430 (N_15430,N_667,N_4658);
nand U15431 (N_15431,N_3137,N_874);
nand U15432 (N_15432,N_7677,N_9527);
nor U15433 (N_15433,N_2956,N_4575);
xnor U15434 (N_15434,N_6878,N_9452);
nor U15435 (N_15435,N_6403,N_7205);
nor U15436 (N_15436,N_8091,N_2365);
or U15437 (N_15437,N_6664,N_4198);
nand U15438 (N_15438,N_8295,N_6154);
and U15439 (N_15439,N_2933,N_1551);
nand U15440 (N_15440,N_2294,N_4396);
xor U15441 (N_15441,N_8813,N_556);
nand U15442 (N_15442,N_7207,N_570);
nand U15443 (N_15443,N_6226,N_7003);
and U15444 (N_15444,N_5534,N_119);
nor U15445 (N_15445,N_2618,N_3933);
nand U15446 (N_15446,N_8823,N_2036);
xnor U15447 (N_15447,N_6640,N_5057);
xnor U15448 (N_15448,N_527,N_6560);
nor U15449 (N_15449,N_2931,N_7561);
nand U15450 (N_15450,N_3405,N_5956);
or U15451 (N_15451,N_2568,N_4638);
and U15452 (N_15452,N_4151,N_4068);
nor U15453 (N_15453,N_7971,N_1775);
nor U15454 (N_15454,N_1439,N_145);
nand U15455 (N_15455,N_4059,N_6177);
or U15456 (N_15456,N_7746,N_6028);
xnor U15457 (N_15457,N_1721,N_9191);
and U15458 (N_15458,N_2413,N_7433);
xnor U15459 (N_15459,N_5970,N_865);
xnor U15460 (N_15460,N_1686,N_8237);
and U15461 (N_15461,N_6049,N_1986);
xor U15462 (N_15462,N_4216,N_618);
nand U15463 (N_15463,N_1361,N_2892);
and U15464 (N_15464,N_1852,N_3106);
and U15465 (N_15465,N_7616,N_1858);
or U15466 (N_15466,N_7004,N_3052);
or U15467 (N_15467,N_4079,N_1503);
and U15468 (N_15468,N_3885,N_127);
or U15469 (N_15469,N_8770,N_6271);
nand U15470 (N_15470,N_1725,N_1531);
and U15471 (N_15471,N_3100,N_657);
nand U15472 (N_15472,N_3617,N_1246);
and U15473 (N_15473,N_5307,N_1044);
nand U15474 (N_15474,N_9570,N_4171);
or U15475 (N_15475,N_4083,N_3502);
or U15476 (N_15476,N_4446,N_291);
and U15477 (N_15477,N_35,N_1951);
or U15478 (N_15478,N_5475,N_8177);
or U15479 (N_15479,N_7547,N_7676);
nand U15480 (N_15480,N_3411,N_7117);
or U15481 (N_15481,N_2434,N_7464);
nand U15482 (N_15482,N_5627,N_8431);
nand U15483 (N_15483,N_9021,N_9005);
xor U15484 (N_15484,N_3851,N_7447);
nand U15485 (N_15485,N_1550,N_5515);
nor U15486 (N_15486,N_2575,N_3471);
nand U15487 (N_15487,N_8847,N_9636);
nor U15488 (N_15488,N_6957,N_6237);
and U15489 (N_15489,N_1364,N_2356);
or U15490 (N_15490,N_6035,N_4245);
or U15491 (N_15491,N_7417,N_10);
xor U15492 (N_15492,N_442,N_1203);
and U15493 (N_15493,N_1282,N_6713);
xor U15494 (N_15494,N_9280,N_5852);
or U15495 (N_15495,N_8372,N_8847);
and U15496 (N_15496,N_4432,N_1374);
xnor U15497 (N_15497,N_367,N_4647);
nand U15498 (N_15498,N_4529,N_402);
or U15499 (N_15499,N_3903,N_5110);
nand U15500 (N_15500,N_144,N_7123);
xnor U15501 (N_15501,N_4774,N_3404);
xor U15502 (N_15502,N_7670,N_8860);
and U15503 (N_15503,N_9098,N_8709);
xor U15504 (N_15504,N_3766,N_1447);
and U15505 (N_15505,N_1388,N_5487);
xnor U15506 (N_15506,N_4662,N_188);
nor U15507 (N_15507,N_7954,N_1242);
or U15508 (N_15508,N_376,N_1980);
xnor U15509 (N_15509,N_9494,N_1467);
xor U15510 (N_15510,N_4996,N_1);
nor U15511 (N_15511,N_110,N_9740);
nand U15512 (N_15512,N_1893,N_8075);
nand U15513 (N_15513,N_476,N_2701);
xnor U15514 (N_15514,N_4159,N_4396);
or U15515 (N_15515,N_1577,N_6157);
or U15516 (N_15516,N_8630,N_4722);
and U15517 (N_15517,N_2896,N_3805);
nor U15518 (N_15518,N_2264,N_2940);
nand U15519 (N_15519,N_8755,N_2400);
and U15520 (N_15520,N_7625,N_9705);
and U15521 (N_15521,N_4797,N_7751);
nor U15522 (N_15522,N_7436,N_7739);
or U15523 (N_15523,N_7268,N_1556);
or U15524 (N_15524,N_4252,N_5215);
nor U15525 (N_15525,N_384,N_6879);
or U15526 (N_15526,N_1221,N_3293);
xor U15527 (N_15527,N_1745,N_7431);
nand U15528 (N_15528,N_5958,N_691);
or U15529 (N_15529,N_2475,N_5802);
and U15530 (N_15530,N_226,N_3972);
nand U15531 (N_15531,N_9741,N_1367);
or U15532 (N_15532,N_5833,N_676);
nand U15533 (N_15533,N_3261,N_2818);
and U15534 (N_15534,N_3177,N_8876);
and U15535 (N_15535,N_4808,N_9239);
nor U15536 (N_15536,N_4510,N_3269);
nand U15537 (N_15537,N_1849,N_8816);
xnor U15538 (N_15538,N_9038,N_6311);
nand U15539 (N_15539,N_7181,N_3896);
or U15540 (N_15540,N_4075,N_3584);
xnor U15541 (N_15541,N_621,N_9622);
or U15542 (N_15542,N_7224,N_5925);
xor U15543 (N_15543,N_3884,N_2678);
nand U15544 (N_15544,N_5173,N_1605);
and U15545 (N_15545,N_5123,N_7560);
and U15546 (N_15546,N_9691,N_6970);
or U15547 (N_15547,N_987,N_9014);
xor U15548 (N_15548,N_463,N_5246);
xnor U15549 (N_15549,N_4735,N_7296);
xnor U15550 (N_15550,N_5070,N_2329);
xor U15551 (N_15551,N_1161,N_3568);
and U15552 (N_15552,N_2600,N_2447);
xor U15553 (N_15553,N_6239,N_7180);
xor U15554 (N_15554,N_6901,N_1920);
or U15555 (N_15555,N_6835,N_5732);
or U15556 (N_15556,N_1523,N_7978);
and U15557 (N_15557,N_9552,N_7987);
nor U15558 (N_15558,N_1509,N_6210);
nor U15559 (N_15559,N_9464,N_9665);
xor U15560 (N_15560,N_5776,N_450);
nor U15561 (N_15561,N_5037,N_9639);
or U15562 (N_15562,N_1786,N_5148);
or U15563 (N_15563,N_9465,N_5829);
and U15564 (N_15564,N_7330,N_2778);
and U15565 (N_15565,N_2772,N_6677);
or U15566 (N_15566,N_6316,N_6370);
or U15567 (N_15567,N_6327,N_6491);
and U15568 (N_15568,N_3790,N_396);
or U15569 (N_15569,N_195,N_2518);
xnor U15570 (N_15570,N_6402,N_462);
nor U15571 (N_15571,N_8760,N_5670);
nand U15572 (N_15572,N_9414,N_4991);
nor U15573 (N_15573,N_7979,N_9933);
nor U15574 (N_15574,N_8916,N_3428);
and U15575 (N_15575,N_3586,N_1425);
nor U15576 (N_15576,N_4199,N_1330);
xor U15577 (N_15577,N_1304,N_9855);
and U15578 (N_15578,N_6037,N_4571);
and U15579 (N_15579,N_4422,N_1393);
xor U15580 (N_15580,N_8478,N_1707);
or U15581 (N_15581,N_1979,N_7418);
nor U15582 (N_15582,N_679,N_3135);
and U15583 (N_15583,N_4813,N_8202);
nor U15584 (N_15584,N_7025,N_1461);
and U15585 (N_15585,N_1402,N_5874);
or U15586 (N_15586,N_3609,N_2559);
nand U15587 (N_15587,N_7867,N_6976);
or U15588 (N_15588,N_9965,N_2264);
nand U15589 (N_15589,N_3222,N_6005);
xnor U15590 (N_15590,N_6148,N_688);
xor U15591 (N_15591,N_1615,N_9681);
xor U15592 (N_15592,N_3507,N_1472);
nor U15593 (N_15593,N_6902,N_1540);
nor U15594 (N_15594,N_629,N_5132);
nor U15595 (N_15595,N_8200,N_7472);
or U15596 (N_15596,N_4919,N_8378);
nor U15597 (N_15597,N_410,N_2601);
and U15598 (N_15598,N_6580,N_3296);
or U15599 (N_15599,N_2373,N_6712);
xnor U15600 (N_15600,N_6586,N_7944);
or U15601 (N_15601,N_75,N_1500);
or U15602 (N_15602,N_8321,N_2389);
nor U15603 (N_15603,N_2235,N_9602);
nor U15604 (N_15604,N_280,N_7539);
and U15605 (N_15605,N_4227,N_7489);
xor U15606 (N_15606,N_6554,N_2395);
xor U15607 (N_15607,N_9,N_1928);
nor U15608 (N_15608,N_3293,N_140);
and U15609 (N_15609,N_91,N_7617);
xnor U15610 (N_15610,N_1957,N_1684);
xnor U15611 (N_15611,N_7611,N_9359);
and U15612 (N_15612,N_5961,N_9075);
xnor U15613 (N_15613,N_3701,N_4318);
or U15614 (N_15614,N_5319,N_8225);
nor U15615 (N_15615,N_9515,N_3359);
nand U15616 (N_15616,N_3194,N_521);
and U15617 (N_15617,N_2069,N_840);
and U15618 (N_15618,N_1062,N_6292);
nor U15619 (N_15619,N_4939,N_210);
and U15620 (N_15620,N_5781,N_4482);
xnor U15621 (N_15621,N_7475,N_7850);
xnor U15622 (N_15622,N_4494,N_8350);
and U15623 (N_15623,N_6846,N_4881);
or U15624 (N_15624,N_8717,N_4496);
nor U15625 (N_15625,N_2413,N_1346);
or U15626 (N_15626,N_1197,N_2972);
nor U15627 (N_15627,N_3736,N_9380);
or U15628 (N_15628,N_9592,N_8501);
or U15629 (N_15629,N_2727,N_7354);
xnor U15630 (N_15630,N_5006,N_8009);
nand U15631 (N_15631,N_9936,N_283);
nand U15632 (N_15632,N_8620,N_6716);
or U15633 (N_15633,N_2499,N_8691);
nand U15634 (N_15634,N_3658,N_6966);
xnor U15635 (N_15635,N_794,N_4947);
or U15636 (N_15636,N_3247,N_5802);
nand U15637 (N_15637,N_6712,N_5146);
or U15638 (N_15638,N_3229,N_873);
and U15639 (N_15639,N_8307,N_36);
or U15640 (N_15640,N_524,N_3801);
nand U15641 (N_15641,N_8518,N_4739);
nor U15642 (N_15642,N_4746,N_896);
or U15643 (N_15643,N_4400,N_3624);
nor U15644 (N_15644,N_2702,N_6564);
nor U15645 (N_15645,N_1359,N_9675);
nand U15646 (N_15646,N_3286,N_6633);
and U15647 (N_15647,N_7975,N_3910);
nand U15648 (N_15648,N_5825,N_8788);
or U15649 (N_15649,N_8205,N_2696);
or U15650 (N_15650,N_6561,N_2920);
xor U15651 (N_15651,N_1757,N_1319);
and U15652 (N_15652,N_360,N_6021);
nor U15653 (N_15653,N_2188,N_9587);
and U15654 (N_15654,N_6207,N_3547);
nand U15655 (N_15655,N_6517,N_3300);
and U15656 (N_15656,N_4328,N_4613);
nor U15657 (N_15657,N_1370,N_6281);
nor U15658 (N_15658,N_6300,N_2388);
xor U15659 (N_15659,N_4322,N_4470);
and U15660 (N_15660,N_8273,N_4954);
xnor U15661 (N_15661,N_4048,N_4250);
xor U15662 (N_15662,N_4308,N_505);
xor U15663 (N_15663,N_4373,N_6029);
nand U15664 (N_15664,N_1238,N_1527);
and U15665 (N_15665,N_5412,N_1109);
xor U15666 (N_15666,N_3434,N_9291);
and U15667 (N_15667,N_1112,N_4890);
nor U15668 (N_15668,N_5074,N_6898);
nand U15669 (N_15669,N_9888,N_2232);
nand U15670 (N_15670,N_4458,N_5657);
xor U15671 (N_15671,N_2821,N_1842);
nor U15672 (N_15672,N_9761,N_3404);
and U15673 (N_15673,N_4645,N_5228);
xnor U15674 (N_15674,N_2270,N_4336);
nand U15675 (N_15675,N_8283,N_9708);
and U15676 (N_15676,N_4468,N_9534);
nand U15677 (N_15677,N_3664,N_2089);
nand U15678 (N_15678,N_3524,N_955);
nand U15679 (N_15679,N_1544,N_547);
or U15680 (N_15680,N_7910,N_4487);
xnor U15681 (N_15681,N_8020,N_4625);
and U15682 (N_15682,N_9675,N_531);
nand U15683 (N_15683,N_8741,N_2229);
or U15684 (N_15684,N_4411,N_8026);
nor U15685 (N_15685,N_7684,N_2266);
nor U15686 (N_15686,N_8992,N_8490);
nand U15687 (N_15687,N_7260,N_5337);
nand U15688 (N_15688,N_3567,N_9853);
nor U15689 (N_15689,N_4751,N_1909);
and U15690 (N_15690,N_6815,N_4484);
and U15691 (N_15691,N_5826,N_6945);
xor U15692 (N_15692,N_9053,N_3519);
or U15693 (N_15693,N_8857,N_7048);
or U15694 (N_15694,N_7160,N_5099);
nand U15695 (N_15695,N_7581,N_4731);
or U15696 (N_15696,N_6212,N_2223);
xnor U15697 (N_15697,N_2412,N_5708);
nor U15698 (N_15698,N_1210,N_6943);
xor U15699 (N_15699,N_9335,N_856);
and U15700 (N_15700,N_298,N_1008);
and U15701 (N_15701,N_9327,N_6730);
xnor U15702 (N_15702,N_851,N_2061);
or U15703 (N_15703,N_6832,N_6884);
nor U15704 (N_15704,N_3785,N_4022);
and U15705 (N_15705,N_3323,N_5840);
and U15706 (N_15706,N_2286,N_9341);
or U15707 (N_15707,N_7898,N_5601);
nand U15708 (N_15708,N_9842,N_640);
and U15709 (N_15709,N_7230,N_9198);
or U15710 (N_15710,N_6243,N_462);
nor U15711 (N_15711,N_3831,N_5177);
nor U15712 (N_15712,N_7630,N_6425);
or U15713 (N_15713,N_5747,N_134);
or U15714 (N_15714,N_8098,N_6057);
nand U15715 (N_15715,N_5575,N_9038);
nor U15716 (N_15716,N_7423,N_7194);
nor U15717 (N_15717,N_3671,N_4365);
nand U15718 (N_15718,N_2562,N_9338);
nor U15719 (N_15719,N_2286,N_6152);
and U15720 (N_15720,N_5545,N_6660);
or U15721 (N_15721,N_6023,N_7314);
xnor U15722 (N_15722,N_970,N_806);
and U15723 (N_15723,N_9483,N_6097);
or U15724 (N_15724,N_4568,N_9441);
nand U15725 (N_15725,N_7406,N_81);
nor U15726 (N_15726,N_4284,N_1995);
or U15727 (N_15727,N_6867,N_5329);
or U15728 (N_15728,N_3339,N_4971);
xor U15729 (N_15729,N_3543,N_4633);
xnor U15730 (N_15730,N_4644,N_124);
nand U15731 (N_15731,N_5960,N_231);
nand U15732 (N_15732,N_356,N_2641);
nor U15733 (N_15733,N_8902,N_4470);
and U15734 (N_15734,N_1256,N_1607);
xnor U15735 (N_15735,N_2756,N_6111);
nor U15736 (N_15736,N_2281,N_5669);
and U15737 (N_15737,N_1021,N_8191);
nand U15738 (N_15738,N_2726,N_5638);
xor U15739 (N_15739,N_2005,N_2123);
or U15740 (N_15740,N_8250,N_6764);
xnor U15741 (N_15741,N_800,N_6424);
or U15742 (N_15742,N_8867,N_3547);
or U15743 (N_15743,N_5045,N_7182);
xor U15744 (N_15744,N_4906,N_6601);
nand U15745 (N_15745,N_3930,N_4585);
xnor U15746 (N_15746,N_2863,N_8342);
xor U15747 (N_15747,N_6790,N_6672);
or U15748 (N_15748,N_4673,N_6144);
or U15749 (N_15749,N_4462,N_1566);
nor U15750 (N_15750,N_5973,N_6589);
nand U15751 (N_15751,N_8117,N_3327);
nor U15752 (N_15752,N_9403,N_5939);
nor U15753 (N_15753,N_6746,N_9428);
xor U15754 (N_15754,N_4042,N_2110);
xor U15755 (N_15755,N_3413,N_2827);
nand U15756 (N_15756,N_6999,N_5193);
or U15757 (N_15757,N_3981,N_1001);
xnor U15758 (N_15758,N_9403,N_8544);
and U15759 (N_15759,N_2259,N_4044);
nand U15760 (N_15760,N_3268,N_8920);
or U15761 (N_15761,N_5415,N_698);
xor U15762 (N_15762,N_8267,N_5182);
and U15763 (N_15763,N_329,N_6537);
or U15764 (N_15764,N_1495,N_9800);
nand U15765 (N_15765,N_530,N_2408);
or U15766 (N_15766,N_2193,N_2261);
nand U15767 (N_15767,N_712,N_40);
xnor U15768 (N_15768,N_3307,N_5349);
nor U15769 (N_15769,N_3434,N_1263);
or U15770 (N_15770,N_957,N_4338);
nand U15771 (N_15771,N_2057,N_1495);
nand U15772 (N_15772,N_6018,N_4998);
nor U15773 (N_15773,N_9591,N_7079);
and U15774 (N_15774,N_1353,N_8633);
xor U15775 (N_15775,N_2409,N_5252);
nor U15776 (N_15776,N_7831,N_1277);
xor U15777 (N_15777,N_9355,N_6541);
and U15778 (N_15778,N_9091,N_6269);
and U15779 (N_15779,N_1464,N_8885);
xor U15780 (N_15780,N_6975,N_1026);
and U15781 (N_15781,N_9349,N_9799);
or U15782 (N_15782,N_1064,N_7310);
xnor U15783 (N_15783,N_4230,N_5927);
xnor U15784 (N_15784,N_5130,N_9073);
xor U15785 (N_15785,N_3694,N_7173);
nand U15786 (N_15786,N_6087,N_3111);
xnor U15787 (N_15787,N_2098,N_2636);
and U15788 (N_15788,N_3149,N_1740);
and U15789 (N_15789,N_1433,N_6481);
and U15790 (N_15790,N_6907,N_7691);
nand U15791 (N_15791,N_3466,N_6477);
or U15792 (N_15792,N_2316,N_1461);
nor U15793 (N_15793,N_7253,N_6362);
or U15794 (N_15794,N_9925,N_358);
and U15795 (N_15795,N_8033,N_9629);
or U15796 (N_15796,N_4793,N_911);
and U15797 (N_15797,N_9162,N_2587);
xnor U15798 (N_15798,N_8663,N_6310);
or U15799 (N_15799,N_1777,N_5375);
nand U15800 (N_15800,N_610,N_1670);
nor U15801 (N_15801,N_1983,N_4407);
nor U15802 (N_15802,N_4116,N_6574);
and U15803 (N_15803,N_394,N_6245);
xnor U15804 (N_15804,N_4247,N_6443);
or U15805 (N_15805,N_8637,N_9160);
nand U15806 (N_15806,N_1308,N_1294);
nand U15807 (N_15807,N_2109,N_6829);
xnor U15808 (N_15808,N_5257,N_3370);
or U15809 (N_15809,N_4631,N_7696);
nor U15810 (N_15810,N_4619,N_5343);
xor U15811 (N_15811,N_5420,N_3387);
nand U15812 (N_15812,N_8246,N_7942);
nor U15813 (N_15813,N_4902,N_8664);
and U15814 (N_15814,N_3845,N_6901);
nand U15815 (N_15815,N_4449,N_2370);
and U15816 (N_15816,N_6712,N_3499);
nor U15817 (N_15817,N_6308,N_2429);
or U15818 (N_15818,N_8004,N_2383);
and U15819 (N_15819,N_8497,N_8342);
xnor U15820 (N_15820,N_3080,N_120);
nor U15821 (N_15821,N_6912,N_9028);
nand U15822 (N_15822,N_8077,N_657);
or U15823 (N_15823,N_6909,N_4729);
nand U15824 (N_15824,N_187,N_7923);
xor U15825 (N_15825,N_2714,N_9609);
xnor U15826 (N_15826,N_1608,N_1286);
or U15827 (N_15827,N_2484,N_2017);
nor U15828 (N_15828,N_4481,N_7767);
or U15829 (N_15829,N_5388,N_1609);
nor U15830 (N_15830,N_573,N_4201);
and U15831 (N_15831,N_9938,N_8883);
nand U15832 (N_15832,N_7335,N_4891);
nand U15833 (N_15833,N_9532,N_9844);
and U15834 (N_15834,N_1244,N_4489);
xor U15835 (N_15835,N_6633,N_1475);
xor U15836 (N_15836,N_2128,N_9980);
nand U15837 (N_15837,N_1455,N_1743);
or U15838 (N_15838,N_2027,N_1845);
nor U15839 (N_15839,N_8647,N_592);
xnor U15840 (N_15840,N_8068,N_9777);
nand U15841 (N_15841,N_5783,N_3365);
nor U15842 (N_15842,N_201,N_4706);
or U15843 (N_15843,N_2586,N_7958);
nor U15844 (N_15844,N_8664,N_7337);
nand U15845 (N_15845,N_1822,N_842);
and U15846 (N_15846,N_5933,N_9549);
nor U15847 (N_15847,N_2913,N_8244);
or U15848 (N_15848,N_7681,N_1108);
or U15849 (N_15849,N_9839,N_6658);
nor U15850 (N_15850,N_1143,N_5698);
and U15851 (N_15851,N_1821,N_6189);
nor U15852 (N_15852,N_7076,N_5880);
nor U15853 (N_15853,N_1035,N_289);
and U15854 (N_15854,N_9404,N_9073);
nor U15855 (N_15855,N_3684,N_2839);
or U15856 (N_15856,N_2329,N_4186);
xor U15857 (N_15857,N_9127,N_8852);
nor U15858 (N_15858,N_1831,N_3626);
nor U15859 (N_15859,N_5413,N_8528);
and U15860 (N_15860,N_1374,N_7535);
xor U15861 (N_15861,N_4190,N_4832);
and U15862 (N_15862,N_1827,N_4761);
xnor U15863 (N_15863,N_9327,N_8923);
and U15864 (N_15864,N_5078,N_162);
and U15865 (N_15865,N_9474,N_330);
or U15866 (N_15866,N_8693,N_5041);
xor U15867 (N_15867,N_9333,N_5011);
nand U15868 (N_15868,N_1514,N_6322);
and U15869 (N_15869,N_5237,N_6568);
nand U15870 (N_15870,N_5969,N_8388);
or U15871 (N_15871,N_5647,N_6793);
nand U15872 (N_15872,N_1347,N_2148);
or U15873 (N_15873,N_1140,N_3781);
nor U15874 (N_15874,N_4976,N_1402);
nor U15875 (N_15875,N_6934,N_9135);
nor U15876 (N_15876,N_2861,N_379);
nand U15877 (N_15877,N_3703,N_183);
nor U15878 (N_15878,N_1440,N_6537);
nor U15879 (N_15879,N_4578,N_4967);
xor U15880 (N_15880,N_2304,N_1620);
nor U15881 (N_15881,N_3897,N_8579);
or U15882 (N_15882,N_690,N_7208);
or U15883 (N_15883,N_8730,N_2607);
nor U15884 (N_15884,N_7457,N_9209);
nor U15885 (N_15885,N_7318,N_88);
nand U15886 (N_15886,N_102,N_8948);
nand U15887 (N_15887,N_9526,N_7122);
xor U15888 (N_15888,N_3094,N_1703);
nor U15889 (N_15889,N_6997,N_9824);
nand U15890 (N_15890,N_9552,N_7634);
xor U15891 (N_15891,N_5535,N_5333);
xnor U15892 (N_15892,N_9949,N_7252);
and U15893 (N_15893,N_2015,N_4939);
nand U15894 (N_15894,N_8580,N_717);
xnor U15895 (N_15895,N_7571,N_4999);
nand U15896 (N_15896,N_887,N_3594);
nor U15897 (N_15897,N_8809,N_7354);
nor U15898 (N_15898,N_9043,N_4849);
nor U15899 (N_15899,N_761,N_9188);
nand U15900 (N_15900,N_1404,N_1384);
nor U15901 (N_15901,N_2907,N_1448);
xnor U15902 (N_15902,N_5574,N_7089);
or U15903 (N_15903,N_9133,N_9208);
nor U15904 (N_15904,N_2314,N_8635);
nand U15905 (N_15905,N_6351,N_8368);
and U15906 (N_15906,N_4607,N_3656);
nand U15907 (N_15907,N_2336,N_4104);
nand U15908 (N_15908,N_4805,N_4586);
or U15909 (N_15909,N_8547,N_616);
nand U15910 (N_15910,N_4901,N_1302);
or U15911 (N_15911,N_4697,N_4879);
or U15912 (N_15912,N_6551,N_2615);
or U15913 (N_15913,N_3847,N_3635);
nor U15914 (N_15914,N_4193,N_8002);
xnor U15915 (N_15915,N_4337,N_899);
xnor U15916 (N_15916,N_9465,N_7370);
or U15917 (N_15917,N_3475,N_3714);
or U15918 (N_15918,N_5585,N_131);
and U15919 (N_15919,N_3673,N_9303);
nand U15920 (N_15920,N_3795,N_4649);
and U15921 (N_15921,N_2879,N_6451);
nand U15922 (N_15922,N_7707,N_5782);
nand U15923 (N_15923,N_7771,N_6188);
xnor U15924 (N_15924,N_1077,N_5062);
xnor U15925 (N_15925,N_9221,N_9902);
nand U15926 (N_15926,N_8088,N_1205);
or U15927 (N_15927,N_7369,N_493);
nor U15928 (N_15928,N_9118,N_3152);
or U15929 (N_15929,N_9176,N_9502);
or U15930 (N_15930,N_4957,N_1319);
nand U15931 (N_15931,N_4391,N_194);
nor U15932 (N_15932,N_7366,N_1515);
or U15933 (N_15933,N_8366,N_9176);
nand U15934 (N_15934,N_3285,N_4858);
nand U15935 (N_15935,N_1720,N_5843);
nor U15936 (N_15936,N_9203,N_9190);
or U15937 (N_15937,N_6032,N_5143);
nand U15938 (N_15938,N_4296,N_9002);
or U15939 (N_15939,N_8717,N_3849);
nand U15940 (N_15940,N_171,N_8155);
or U15941 (N_15941,N_2291,N_6399);
nand U15942 (N_15942,N_3968,N_1079);
and U15943 (N_15943,N_1403,N_4728);
nor U15944 (N_15944,N_658,N_8454);
nor U15945 (N_15945,N_6038,N_1601);
and U15946 (N_15946,N_390,N_1313);
nor U15947 (N_15947,N_4729,N_826);
nor U15948 (N_15948,N_208,N_1099);
and U15949 (N_15949,N_3784,N_3447);
or U15950 (N_15950,N_7873,N_7036);
nor U15951 (N_15951,N_1028,N_9901);
xor U15952 (N_15952,N_534,N_2306);
nand U15953 (N_15953,N_9314,N_8090);
or U15954 (N_15954,N_6914,N_5723);
nand U15955 (N_15955,N_5974,N_3109);
nand U15956 (N_15956,N_2748,N_6894);
xor U15957 (N_15957,N_1428,N_9669);
or U15958 (N_15958,N_6273,N_9303);
or U15959 (N_15959,N_2105,N_900);
xnor U15960 (N_15960,N_7041,N_9615);
xnor U15961 (N_15961,N_6143,N_8063);
nand U15962 (N_15962,N_4803,N_3573);
nand U15963 (N_15963,N_5765,N_2384);
and U15964 (N_15964,N_4725,N_7248);
or U15965 (N_15965,N_9298,N_9887);
nor U15966 (N_15966,N_6018,N_3349);
nand U15967 (N_15967,N_3035,N_5010);
nand U15968 (N_15968,N_1660,N_8211);
nor U15969 (N_15969,N_4315,N_4443);
and U15970 (N_15970,N_8296,N_2031);
or U15971 (N_15971,N_5307,N_4402);
and U15972 (N_15972,N_2685,N_5257);
and U15973 (N_15973,N_8013,N_636);
and U15974 (N_15974,N_3297,N_7211);
and U15975 (N_15975,N_1722,N_9641);
and U15976 (N_15976,N_979,N_7074);
xnor U15977 (N_15977,N_6364,N_4581);
xor U15978 (N_15978,N_8711,N_9381);
or U15979 (N_15979,N_9268,N_5986);
and U15980 (N_15980,N_918,N_4115);
and U15981 (N_15981,N_3585,N_6405);
xnor U15982 (N_15982,N_120,N_3439);
nor U15983 (N_15983,N_7544,N_3244);
nor U15984 (N_15984,N_8444,N_1713);
nand U15985 (N_15985,N_2567,N_6103);
or U15986 (N_15986,N_2244,N_9349);
nor U15987 (N_15987,N_6687,N_3881);
xor U15988 (N_15988,N_1651,N_3074);
nand U15989 (N_15989,N_5436,N_6636);
or U15990 (N_15990,N_8360,N_5129);
xnor U15991 (N_15991,N_5692,N_399);
nor U15992 (N_15992,N_6790,N_9022);
xor U15993 (N_15993,N_3694,N_8100);
or U15994 (N_15994,N_3874,N_1266);
or U15995 (N_15995,N_5128,N_9092);
nor U15996 (N_15996,N_2228,N_3690);
or U15997 (N_15997,N_5640,N_1786);
nor U15998 (N_15998,N_6277,N_9427);
nor U15999 (N_15999,N_3100,N_4879);
and U16000 (N_16000,N_2322,N_2034);
and U16001 (N_16001,N_8538,N_7848);
or U16002 (N_16002,N_9967,N_5336);
and U16003 (N_16003,N_6333,N_3120);
and U16004 (N_16004,N_7808,N_8566);
xnor U16005 (N_16005,N_355,N_4064);
or U16006 (N_16006,N_9525,N_9098);
and U16007 (N_16007,N_2,N_8658);
nand U16008 (N_16008,N_7579,N_9376);
nor U16009 (N_16009,N_3510,N_2079);
nand U16010 (N_16010,N_5339,N_4127);
nor U16011 (N_16011,N_7075,N_1294);
or U16012 (N_16012,N_616,N_2317);
nand U16013 (N_16013,N_2452,N_6906);
or U16014 (N_16014,N_1581,N_9546);
nor U16015 (N_16015,N_5260,N_1269);
nand U16016 (N_16016,N_8398,N_9987);
nor U16017 (N_16017,N_836,N_2976);
or U16018 (N_16018,N_9372,N_3017);
xor U16019 (N_16019,N_2237,N_7484);
and U16020 (N_16020,N_7730,N_7364);
and U16021 (N_16021,N_4269,N_173);
nand U16022 (N_16022,N_7981,N_4579);
xnor U16023 (N_16023,N_7065,N_9678);
nand U16024 (N_16024,N_9941,N_400);
nor U16025 (N_16025,N_561,N_7285);
or U16026 (N_16026,N_3667,N_7561);
nor U16027 (N_16027,N_4826,N_5983);
nand U16028 (N_16028,N_1420,N_2522);
xnor U16029 (N_16029,N_9677,N_5956);
xor U16030 (N_16030,N_7066,N_5666);
nor U16031 (N_16031,N_6864,N_6136);
xor U16032 (N_16032,N_3296,N_6666);
nor U16033 (N_16033,N_9959,N_4179);
xnor U16034 (N_16034,N_9635,N_2951);
xor U16035 (N_16035,N_2631,N_9743);
xnor U16036 (N_16036,N_3544,N_8140);
or U16037 (N_16037,N_2597,N_9157);
xnor U16038 (N_16038,N_8389,N_775);
nor U16039 (N_16039,N_977,N_6224);
xor U16040 (N_16040,N_2162,N_3511);
nand U16041 (N_16041,N_5822,N_5395);
nor U16042 (N_16042,N_7291,N_2537);
or U16043 (N_16043,N_9353,N_3496);
nor U16044 (N_16044,N_2200,N_7116);
or U16045 (N_16045,N_6824,N_7558);
nand U16046 (N_16046,N_5499,N_4019);
nor U16047 (N_16047,N_7829,N_2484);
nor U16048 (N_16048,N_9080,N_5882);
or U16049 (N_16049,N_9215,N_1200);
nor U16050 (N_16050,N_1507,N_2105);
and U16051 (N_16051,N_139,N_4580);
nand U16052 (N_16052,N_3189,N_8816);
or U16053 (N_16053,N_7868,N_1321);
and U16054 (N_16054,N_2149,N_9850);
nand U16055 (N_16055,N_812,N_4321);
xnor U16056 (N_16056,N_534,N_9967);
or U16057 (N_16057,N_3941,N_2050);
nor U16058 (N_16058,N_6747,N_3571);
nand U16059 (N_16059,N_7549,N_2808);
or U16060 (N_16060,N_9831,N_8697);
or U16061 (N_16061,N_9996,N_5253);
nor U16062 (N_16062,N_8675,N_5610);
nor U16063 (N_16063,N_523,N_3359);
xnor U16064 (N_16064,N_5448,N_3274);
nand U16065 (N_16065,N_1154,N_283);
or U16066 (N_16066,N_8016,N_5679);
or U16067 (N_16067,N_4624,N_7317);
and U16068 (N_16068,N_1441,N_4294);
nor U16069 (N_16069,N_5782,N_6358);
or U16070 (N_16070,N_5674,N_7947);
nand U16071 (N_16071,N_1671,N_6410);
nor U16072 (N_16072,N_3166,N_8090);
or U16073 (N_16073,N_920,N_2559);
xor U16074 (N_16074,N_4959,N_1888);
and U16075 (N_16075,N_9094,N_906);
or U16076 (N_16076,N_9602,N_9893);
and U16077 (N_16077,N_2758,N_1114);
nand U16078 (N_16078,N_3561,N_8808);
nand U16079 (N_16079,N_9445,N_5860);
nor U16080 (N_16080,N_5109,N_8894);
or U16081 (N_16081,N_3397,N_1343);
and U16082 (N_16082,N_8523,N_4027);
nor U16083 (N_16083,N_6612,N_4049);
nor U16084 (N_16084,N_9272,N_4758);
nor U16085 (N_16085,N_8146,N_7774);
and U16086 (N_16086,N_6753,N_8006);
xor U16087 (N_16087,N_8104,N_5580);
and U16088 (N_16088,N_9844,N_4991);
nor U16089 (N_16089,N_831,N_1312);
or U16090 (N_16090,N_250,N_608);
and U16091 (N_16091,N_3467,N_747);
xor U16092 (N_16092,N_8224,N_1000);
nor U16093 (N_16093,N_5298,N_2179);
or U16094 (N_16094,N_5376,N_1664);
or U16095 (N_16095,N_8486,N_5454);
and U16096 (N_16096,N_9084,N_7983);
or U16097 (N_16097,N_4040,N_9473);
nor U16098 (N_16098,N_4048,N_1928);
nor U16099 (N_16099,N_8045,N_4409);
nor U16100 (N_16100,N_1264,N_6434);
and U16101 (N_16101,N_8501,N_3126);
nand U16102 (N_16102,N_3051,N_7059);
nor U16103 (N_16103,N_5600,N_3337);
nor U16104 (N_16104,N_112,N_7465);
xnor U16105 (N_16105,N_867,N_3205);
nand U16106 (N_16106,N_2857,N_9084);
nand U16107 (N_16107,N_2423,N_1970);
xor U16108 (N_16108,N_4906,N_8807);
xor U16109 (N_16109,N_2680,N_3411);
or U16110 (N_16110,N_4345,N_5263);
nor U16111 (N_16111,N_1505,N_5470);
xnor U16112 (N_16112,N_5095,N_3555);
and U16113 (N_16113,N_4758,N_2582);
xor U16114 (N_16114,N_4164,N_1270);
and U16115 (N_16115,N_6296,N_6994);
nor U16116 (N_16116,N_5621,N_979);
nor U16117 (N_16117,N_2924,N_9613);
xnor U16118 (N_16118,N_7130,N_8289);
nor U16119 (N_16119,N_3757,N_6677);
or U16120 (N_16120,N_8741,N_3630);
xor U16121 (N_16121,N_4810,N_2128);
and U16122 (N_16122,N_2342,N_9400);
nand U16123 (N_16123,N_7621,N_1640);
nor U16124 (N_16124,N_577,N_493);
nor U16125 (N_16125,N_8534,N_5803);
and U16126 (N_16126,N_8112,N_713);
xor U16127 (N_16127,N_8613,N_2054);
or U16128 (N_16128,N_3229,N_5212);
and U16129 (N_16129,N_5196,N_7724);
or U16130 (N_16130,N_2392,N_5579);
nand U16131 (N_16131,N_5408,N_7045);
nand U16132 (N_16132,N_9398,N_5005);
xnor U16133 (N_16133,N_5371,N_4837);
nand U16134 (N_16134,N_4157,N_9227);
or U16135 (N_16135,N_2095,N_8771);
and U16136 (N_16136,N_5746,N_9098);
nand U16137 (N_16137,N_8231,N_9377);
nand U16138 (N_16138,N_9581,N_8676);
nor U16139 (N_16139,N_5767,N_6180);
nor U16140 (N_16140,N_6138,N_5668);
nand U16141 (N_16141,N_3671,N_1579);
and U16142 (N_16142,N_8883,N_8051);
nand U16143 (N_16143,N_727,N_3989);
nor U16144 (N_16144,N_4439,N_2187);
nor U16145 (N_16145,N_922,N_4522);
xnor U16146 (N_16146,N_5831,N_4897);
nor U16147 (N_16147,N_3701,N_5503);
or U16148 (N_16148,N_4300,N_4220);
and U16149 (N_16149,N_5417,N_3843);
or U16150 (N_16150,N_7955,N_6287);
nor U16151 (N_16151,N_8402,N_3617);
nor U16152 (N_16152,N_8155,N_8497);
nand U16153 (N_16153,N_346,N_3589);
and U16154 (N_16154,N_9635,N_4729);
or U16155 (N_16155,N_7397,N_8768);
nor U16156 (N_16156,N_6224,N_6753);
or U16157 (N_16157,N_503,N_9675);
nor U16158 (N_16158,N_5049,N_5163);
nor U16159 (N_16159,N_7217,N_8178);
xnor U16160 (N_16160,N_3864,N_9793);
nand U16161 (N_16161,N_1293,N_9729);
and U16162 (N_16162,N_5184,N_8214);
nor U16163 (N_16163,N_7907,N_4385);
nand U16164 (N_16164,N_7387,N_7757);
xor U16165 (N_16165,N_3418,N_8442);
xnor U16166 (N_16166,N_9396,N_2197);
nor U16167 (N_16167,N_9436,N_732);
nand U16168 (N_16168,N_2008,N_4641);
xnor U16169 (N_16169,N_5077,N_5657);
and U16170 (N_16170,N_5751,N_6112);
and U16171 (N_16171,N_8157,N_9535);
nand U16172 (N_16172,N_5818,N_2402);
or U16173 (N_16173,N_9317,N_4534);
and U16174 (N_16174,N_832,N_5919);
and U16175 (N_16175,N_8380,N_1549);
or U16176 (N_16176,N_6466,N_3055);
or U16177 (N_16177,N_5942,N_5274);
or U16178 (N_16178,N_5681,N_2420);
or U16179 (N_16179,N_4812,N_4446);
or U16180 (N_16180,N_8334,N_6772);
nor U16181 (N_16181,N_5431,N_9587);
nor U16182 (N_16182,N_583,N_9643);
nor U16183 (N_16183,N_9017,N_8802);
nand U16184 (N_16184,N_5189,N_6473);
nor U16185 (N_16185,N_6814,N_2208);
nor U16186 (N_16186,N_5696,N_7610);
or U16187 (N_16187,N_7394,N_5330);
and U16188 (N_16188,N_2354,N_4029);
or U16189 (N_16189,N_1892,N_2575);
nor U16190 (N_16190,N_9010,N_6739);
xor U16191 (N_16191,N_9100,N_9426);
and U16192 (N_16192,N_9809,N_868);
xor U16193 (N_16193,N_3578,N_3756);
nand U16194 (N_16194,N_9628,N_4027);
and U16195 (N_16195,N_9174,N_5451);
or U16196 (N_16196,N_5859,N_5511);
nand U16197 (N_16197,N_7396,N_2480);
or U16198 (N_16198,N_7600,N_9240);
xor U16199 (N_16199,N_5727,N_9307);
xnor U16200 (N_16200,N_6080,N_3847);
nand U16201 (N_16201,N_2079,N_5073);
or U16202 (N_16202,N_214,N_6867);
and U16203 (N_16203,N_2024,N_5425);
xor U16204 (N_16204,N_6493,N_4696);
or U16205 (N_16205,N_667,N_461);
or U16206 (N_16206,N_7170,N_1648);
nor U16207 (N_16207,N_5096,N_4117);
or U16208 (N_16208,N_7057,N_6921);
nor U16209 (N_16209,N_5039,N_4077);
or U16210 (N_16210,N_6597,N_6485);
and U16211 (N_16211,N_7867,N_8167);
and U16212 (N_16212,N_106,N_2617);
or U16213 (N_16213,N_7733,N_8777);
or U16214 (N_16214,N_7841,N_9144);
nand U16215 (N_16215,N_7097,N_1867);
or U16216 (N_16216,N_910,N_2355);
and U16217 (N_16217,N_3210,N_7659);
nand U16218 (N_16218,N_177,N_7313);
and U16219 (N_16219,N_7361,N_5375);
or U16220 (N_16220,N_3517,N_8579);
or U16221 (N_16221,N_1424,N_9689);
nor U16222 (N_16222,N_8180,N_6092);
nor U16223 (N_16223,N_7279,N_3126);
nand U16224 (N_16224,N_1277,N_828);
or U16225 (N_16225,N_5194,N_5643);
nand U16226 (N_16226,N_3225,N_9559);
nand U16227 (N_16227,N_2320,N_4235);
xor U16228 (N_16228,N_663,N_4293);
nor U16229 (N_16229,N_4251,N_7651);
or U16230 (N_16230,N_4787,N_2607);
nand U16231 (N_16231,N_4488,N_8337);
xor U16232 (N_16232,N_1777,N_2125);
nor U16233 (N_16233,N_6973,N_3152);
xor U16234 (N_16234,N_8974,N_2015);
and U16235 (N_16235,N_5056,N_7629);
nor U16236 (N_16236,N_3040,N_5380);
xnor U16237 (N_16237,N_7138,N_1404);
xnor U16238 (N_16238,N_2052,N_962);
xnor U16239 (N_16239,N_54,N_7639);
and U16240 (N_16240,N_9110,N_8507);
and U16241 (N_16241,N_9343,N_4868);
nand U16242 (N_16242,N_7633,N_4941);
nand U16243 (N_16243,N_5758,N_3454);
nor U16244 (N_16244,N_7326,N_6707);
and U16245 (N_16245,N_3119,N_9055);
and U16246 (N_16246,N_9136,N_2860);
nand U16247 (N_16247,N_2124,N_666);
and U16248 (N_16248,N_2343,N_7401);
nor U16249 (N_16249,N_8450,N_9960);
nand U16250 (N_16250,N_7312,N_6705);
and U16251 (N_16251,N_690,N_8966);
and U16252 (N_16252,N_2584,N_1926);
nor U16253 (N_16253,N_8762,N_6726);
nor U16254 (N_16254,N_7792,N_5155);
xnor U16255 (N_16255,N_5590,N_6391);
xnor U16256 (N_16256,N_8045,N_9587);
xor U16257 (N_16257,N_9006,N_3926);
or U16258 (N_16258,N_4541,N_9081);
nor U16259 (N_16259,N_9364,N_7981);
xor U16260 (N_16260,N_7419,N_8625);
and U16261 (N_16261,N_5853,N_1418);
nor U16262 (N_16262,N_5010,N_3464);
nor U16263 (N_16263,N_5643,N_6020);
xnor U16264 (N_16264,N_8184,N_7993);
nand U16265 (N_16265,N_8272,N_6694);
and U16266 (N_16266,N_7606,N_1490);
or U16267 (N_16267,N_7664,N_6683);
and U16268 (N_16268,N_7370,N_5300);
nand U16269 (N_16269,N_6383,N_3452);
nand U16270 (N_16270,N_2505,N_8597);
nand U16271 (N_16271,N_4955,N_4093);
xnor U16272 (N_16272,N_8642,N_7171);
or U16273 (N_16273,N_3008,N_7043);
xor U16274 (N_16274,N_2898,N_1507);
xnor U16275 (N_16275,N_3776,N_7341);
nand U16276 (N_16276,N_7398,N_8663);
nand U16277 (N_16277,N_334,N_1654);
nand U16278 (N_16278,N_4963,N_5928);
or U16279 (N_16279,N_2823,N_5139);
xor U16280 (N_16280,N_8359,N_9435);
nor U16281 (N_16281,N_3794,N_1925);
and U16282 (N_16282,N_8689,N_5639);
nand U16283 (N_16283,N_2352,N_2767);
and U16284 (N_16284,N_5134,N_9441);
or U16285 (N_16285,N_5500,N_2822);
or U16286 (N_16286,N_5665,N_7327);
nand U16287 (N_16287,N_1549,N_4049);
xor U16288 (N_16288,N_5554,N_2461);
or U16289 (N_16289,N_1236,N_6398);
xnor U16290 (N_16290,N_1637,N_1745);
nand U16291 (N_16291,N_9856,N_1957);
nor U16292 (N_16292,N_6273,N_1325);
nor U16293 (N_16293,N_309,N_204);
nor U16294 (N_16294,N_9706,N_4103);
nand U16295 (N_16295,N_8922,N_1291);
xor U16296 (N_16296,N_6056,N_7983);
and U16297 (N_16297,N_4185,N_5512);
and U16298 (N_16298,N_7380,N_859);
and U16299 (N_16299,N_2499,N_2702);
xnor U16300 (N_16300,N_7300,N_2390);
nand U16301 (N_16301,N_7070,N_3266);
nand U16302 (N_16302,N_9994,N_6045);
and U16303 (N_16303,N_7110,N_1536);
and U16304 (N_16304,N_1340,N_3553);
and U16305 (N_16305,N_6181,N_6892);
nand U16306 (N_16306,N_1000,N_1079);
nand U16307 (N_16307,N_2127,N_6464);
nand U16308 (N_16308,N_7365,N_3819);
nor U16309 (N_16309,N_4400,N_1278);
or U16310 (N_16310,N_9937,N_3510);
and U16311 (N_16311,N_4650,N_2195);
nand U16312 (N_16312,N_9296,N_3003);
xor U16313 (N_16313,N_2956,N_1068);
nor U16314 (N_16314,N_7960,N_7526);
nor U16315 (N_16315,N_4401,N_9957);
nand U16316 (N_16316,N_9035,N_1297);
xor U16317 (N_16317,N_2662,N_7298);
nand U16318 (N_16318,N_6947,N_7751);
nor U16319 (N_16319,N_7219,N_1930);
xor U16320 (N_16320,N_5242,N_3017);
or U16321 (N_16321,N_7219,N_9678);
or U16322 (N_16322,N_7787,N_8087);
nand U16323 (N_16323,N_5427,N_6975);
nor U16324 (N_16324,N_9460,N_4920);
xor U16325 (N_16325,N_9381,N_5918);
and U16326 (N_16326,N_1366,N_1031);
xnor U16327 (N_16327,N_3670,N_8646);
nor U16328 (N_16328,N_6763,N_2557);
nand U16329 (N_16329,N_4061,N_9586);
and U16330 (N_16330,N_7118,N_8283);
or U16331 (N_16331,N_8470,N_9518);
and U16332 (N_16332,N_8840,N_799);
and U16333 (N_16333,N_6416,N_1031);
xnor U16334 (N_16334,N_3404,N_5501);
xor U16335 (N_16335,N_5251,N_6894);
nor U16336 (N_16336,N_3346,N_2109);
xnor U16337 (N_16337,N_8687,N_9238);
xor U16338 (N_16338,N_106,N_744);
nand U16339 (N_16339,N_6945,N_4701);
xnor U16340 (N_16340,N_5744,N_4536);
and U16341 (N_16341,N_6202,N_600);
nor U16342 (N_16342,N_657,N_1222);
nor U16343 (N_16343,N_3167,N_1747);
and U16344 (N_16344,N_1883,N_1857);
and U16345 (N_16345,N_8770,N_892);
and U16346 (N_16346,N_7047,N_9096);
xor U16347 (N_16347,N_3393,N_4783);
and U16348 (N_16348,N_790,N_4481);
nor U16349 (N_16349,N_9297,N_4294);
xnor U16350 (N_16350,N_298,N_2532);
or U16351 (N_16351,N_6342,N_9642);
xor U16352 (N_16352,N_7222,N_8469);
nand U16353 (N_16353,N_5497,N_8482);
or U16354 (N_16354,N_9589,N_823);
xor U16355 (N_16355,N_7107,N_9248);
or U16356 (N_16356,N_3446,N_6128);
or U16357 (N_16357,N_9757,N_2329);
and U16358 (N_16358,N_1932,N_3775);
or U16359 (N_16359,N_2573,N_2511);
nand U16360 (N_16360,N_7560,N_218);
and U16361 (N_16361,N_8283,N_7319);
xnor U16362 (N_16362,N_2537,N_88);
or U16363 (N_16363,N_4593,N_413);
nor U16364 (N_16364,N_5006,N_928);
nand U16365 (N_16365,N_9519,N_3934);
and U16366 (N_16366,N_8655,N_9356);
xnor U16367 (N_16367,N_1621,N_3653);
xor U16368 (N_16368,N_688,N_6389);
nor U16369 (N_16369,N_688,N_9597);
or U16370 (N_16370,N_1443,N_4808);
or U16371 (N_16371,N_4965,N_6351);
nand U16372 (N_16372,N_9096,N_7812);
and U16373 (N_16373,N_9373,N_5562);
xor U16374 (N_16374,N_40,N_4589);
or U16375 (N_16375,N_6034,N_4135);
nand U16376 (N_16376,N_6056,N_3964);
nand U16377 (N_16377,N_297,N_918);
nor U16378 (N_16378,N_1260,N_1245);
xor U16379 (N_16379,N_3460,N_675);
and U16380 (N_16380,N_3973,N_8102);
nor U16381 (N_16381,N_9785,N_1311);
xor U16382 (N_16382,N_614,N_8987);
and U16383 (N_16383,N_2967,N_471);
nor U16384 (N_16384,N_326,N_7996);
and U16385 (N_16385,N_5513,N_876);
or U16386 (N_16386,N_1820,N_4522);
or U16387 (N_16387,N_3813,N_2271);
xnor U16388 (N_16388,N_6403,N_7029);
or U16389 (N_16389,N_6625,N_2688);
and U16390 (N_16390,N_9487,N_1906);
nor U16391 (N_16391,N_6591,N_5745);
nor U16392 (N_16392,N_6404,N_7203);
nor U16393 (N_16393,N_3557,N_213);
xor U16394 (N_16394,N_243,N_8279);
xor U16395 (N_16395,N_9961,N_263);
or U16396 (N_16396,N_9169,N_4355);
and U16397 (N_16397,N_6410,N_587);
nand U16398 (N_16398,N_2033,N_4671);
nand U16399 (N_16399,N_387,N_4337);
nand U16400 (N_16400,N_9007,N_2544);
nor U16401 (N_16401,N_6517,N_8481);
xnor U16402 (N_16402,N_9480,N_349);
nor U16403 (N_16403,N_7559,N_2713);
nand U16404 (N_16404,N_3217,N_5227);
xnor U16405 (N_16405,N_739,N_9830);
or U16406 (N_16406,N_9607,N_2153);
nand U16407 (N_16407,N_6626,N_4746);
or U16408 (N_16408,N_5888,N_8270);
or U16409 (N_16409,N_4892,N_9163);
nor U16410 (N_16410,N_4420,N_6662);
and U16411 (N_16411,N_6272,N_3978);
and U16412 (N_16412,N_6721,N_9610);
nand U16413 (N_16413,N_1248,N_3067);
nor U16414 (N_16414,N_380,N_8112);
and U16415 (N_16415,N_6193,N_5670);
xor U16416 (N_16416,N_9741,N_8853);
xor U16417 (N_16417,N_2063,N_694);
nor U16418 (N_16418,N_6497,N_4987);
nor U16419 (N_16419,N_7536,N_2811);
xnor U16420 (N_16420,N_5648,N_3081);
nor U16421 (N_16421,N_3080,N_2608);
nor U16422 (N_16422,N_1515,N_6056);
xor U16423 (N_16423,N_4888,N_7792);
nor U16424 (N_16424,N_7661,N_2713);
and U16425 (N_16425,N_3385,N_7015);
xnor U16426 (N_16426,N_5845,N_1116);
xor U16427 (N_16427,N_209,N_2397);
or U16428 (N_16428,N_5240,N_5831);
or U16429 (N_16429,N_1594,N_4392);
nand U16430 (N_16430,N_381,N_891);
xnor U16431 (N_16431,N_2571,N_9992);
nand U16432 (N_16432,N_8682,N_760);
or U16433 (N_16433,N_2281,N_344);
and U16434 (N_16434,N_4399,N_3897);
or U16435 (N_16435,N_5352,N_3629);
xnor U16436 (N_16436,N_5348,N_2764);
nand U16437 (N_16437,N_3925,N_4190);
and U16438 (N_16438,N_2071,N_5604);
xnor U16439 (N_16439,N_1690,N_6735);
nor U16440 (N_16440,N_9112,N_3804);
xor U16441 (N_16441,N_8350,N_6954);
xor U16442 (N_16442,N_3620,N_551);
nor U16443 (N_16443,N_1536,N_2977);
xnor U16444 (N_16444,N_4822,N_5960);
and U16445 (N_16445,N_9686,N_5177);
or U16446 (N_16446,N_7706,N_3979);
nand U16447 (N_16447,N_2057,N_3156);
and U16448 (N_16448,N_7040,N_9010);
nand U16449 (N_16449,N_1145,N_7723);
xnor U16450 (N_16450,N_389,N_4868);
nor U16451 (N_16451,N_2152,N_3693);
nand U16452 (N_16452,N_6354,N_6415);
nand U16453 (N_16453,N_4219,N_525);
nor U16454 (N_16454,N_7243,N_4283);
nor U16455 (N_16455,N_9031,N_5934);
nor U16456 (N_16456,N_1716,N_9510);
and U16457 (N_16457,N_1560,N_4392);
or U16458 (N_16458,N_3965,N_9609);
nor U16459 (N_16459,N_8668,N_5189);
xor U16460 (N_16460,N_1409,N_1805);
nor U16461 (N_16461,N_911,N_4873);
or U16462 (N_16462,N_1219,N_1041);
and U16463 (N_16463,N_4788,N_2184);
and U16464 (N_16464,N_9233,N_4102);
nor U16465 (N_16465,N_9249,N_5661);
and U16466 (N_16466,N_1216,N_8309);
and U16467 (N_16467,N_3267,N_8014);
and U16468 (N_16468,N_2478,N_3004);
xor U16469 (N_16469,N_3593,N_7506);
xor U16470 (N_16470,N_7838,N_5368);
nor U16471 (N_16471,N_8054,N_4639);
and U16472 (N_16472,N_3929,N_8905);
and U16473 (N_16473,N_5553,N_8321);
nand U16474 (N_16474,N_2893,N_5831);
and U16475 (N_16475,N_287,N_1800);
and U16476 (N_16476,N_5554,N_8683);
or U16477 (N_16477,N_4172,N_8152);
nand U16478 (N_16478,N_8088,N_9684);
nand U16479 (N_16479,N_9083,N_7806);
or U16480 (N_16480,N_6276,N_1986);
and U16481 (N_16481,N_6764,N_898);
or U16482 (N_16482,N_7724,N_5436);
nand U16483 (N_16483,N_31,N_7187);
or U16484 (N_16484,N_9540,N_6169);
nand U16485 (N_16485,N_7037,N_2454);
nor U16486 (N_16486,N_6960,N_8752);
xnor U16487 (N_16487,N_8399,N_2508);
xnor U16488 (N_16488,N_6976,N_9741);
and U16489 (N_16489,N_6450,N_150);
or U16490 (N_16490,N_5608,N_625);
or U16491 (N_16491,N_7829,N_2722);
xnor U16492 (N_16492,N_9487,N_2220);
or U16493 (N_16493,N_9647,N_8658);
xnor U16494 (N_16494,N_6762,N_9414);
xnor U16495 (N_16495,N_4416,N_8719);
or U16496 (N_16496,N_8930,N_4714);
nor U16497 (N_16497,N_3493,N_8592);
and U16498 (N_16498,N_7637,N_168);
xor U16499 (N_16499,N_4324,N_4685);
nand U16500 (N_16500,N_3004,N_2784);
nand U16501 (N_16501,N_4371,N_7219);
xnor U16502 (N_16502,N_4158,N_6307);
and U16503 (N_16503,N_4212,N_3973);
or U16504 (N_16504,N_9330,N_9304);
and U16505 (N_16505,N_4508,N_6058);
and U16506 (N_16506,N_1440,N_8787);
or U16507 (N_16507,N_9336,N_2165);
or U16508 (N_16508,N_1178,N_7524);
nand U16509 (N_16509,N_275,N_1456);
xnor U16510 (N_16510,N_9559,N_5612);
xnor U16511 (N_16511,N_704,N_1242);
nor U16512 (N_16512,N_6412,N_1915);
nand U16513 (N_16513,N_2595,N_6345);
or U16514 (N_16514,N_7029,N_9521);
xor U16515 (N_16515,N_7409,N_1289);
nand U16516 (N_16516,N_5640,N_3503);
nor U16517 (N_16517,N_2709,N_4051);
or U16518 (N_16518,N_5430,N_8854);
nor U16519 (N_16519,N_236,N_8970);
nor U16520 (N_16520,N_5662,N_7714);
nor U16521 (N_16521,N_773,N_8729);
or U16522 (N_16522,N_7540,N_7570);
nor U16523 (N_16523,N_8262,N_3738);
and U16524 (N_16524,N_1627,N_4106);
or U16525 (N_16525,N_374,N_7564);
or U16526 (N_16526,N_6546,N_2433);
or U16527 (N_16527,N_1184,N_6466);
nand U16528 (N_16528,N_1876,N_4486);
or U16529 (N_16529,N_40,N_685);
or U16530 (N_16530,N_2753,N_9604);
xnor U16531 (N_16531,N_1915,N_8959);
xor U16532 (N_16532,N_5774,N_4121);
xnor U16533 (N_16533,N_7584,N_578);
nand U16534 (N_16534,N_2974,N_8894);
or U16535 (N_16535,N_7100,N_2123);
nand U16536 (N_16536,N_2920,N_6990);
nand U16537 (N_16537,N_8510,N_9119);
and U16538 (N_16538,N_6431,N_7348);
and U16539 (N_16539,N_580,N_4305);
nor U16540 (N_16540,N_2373,N_6800);
nand U16541 (N_16541,N_5184,N_5377);
xor U16542 (N_16542,N_3799,N_9728);
xor U16543 (N_16543,N_1526,N_8389);
nand U16544 (N_16544,N_3189,N_8311);
xor U16545 (N_16545,N_6221,N_777);
nor U16546 (N_16546,N_5354,N_6660);
nand U16547 (N_16547,N_4614,N_9048);
nand U16548 (N_16548,N_8277,N_4270);
xnor U16549 (N_16549,N_927,N_2978);
or U16550 (N_16550,N_5613,N_4661);
nand U16551 (N_16551,N_5095,N_6808);
xor U16552 (N_16552,N_8659,N_3780);
and U16553 (N_16553,N_9872,N_9347);
xor U16554 (N_16554,N_8274,N_8581);
or U16555 (N_16555,N_9911,N_9003);
nand U16556 (N_16556,N_1460,N_7625);
and U16557 (N_16557,N_8816,N_7974);
xor U16558 (N_16558,N_2716,N_9934);
and U16559 (N_16559,N_9763,N_7969);
nor U16560 (N_16560,N_6372,N_5221);
and U16561 (N_16561,N_3813,N_5974);
nand U16562 (N_16562,N_6186,N_4164);
nor U16563 (N_16563,N_4390,N_4202);
nand U16564 (N_16564,N_5875,N_2327);
nand U16565 (N_16565,N_1867,N_3931);
or U16566 (N_16566,N_1149,N_9840);
and U16567 (N_16567,N_7232,N_1260);
nor U16568 (N_16568,N_2973,N_2396);
or U16569 (N_16569,N_5633,N_1379);
nor U16570 (N_16570,N_941,N_8485);
xor U16571 (N_16571,N_1513,N_5233);
xor U16572 (N_16572,N_6393,N_514);
xnor U16573 (N_16573,N_1107,N_2407);
xnor U16574 (N_16574,N_6315,N_800);
nand U16575 (N_16575,N_2431,N_9143);
nand U16576 (N_16576,N_7311,N_5316);
xor U16577 (N_16577,N_1607,N_1970);
xnor U16578 (N_16578,N_5458,N_2344);
or U16579 (N_16579,N_2837,N_7414);
or U16580 (N_16580,N_6793,N_9917);
or U16581 (N_16581,N_3958,N_5148);
nand U16582 (N_16582,N_750,N_7098);
nand U16583 (N_16583,N_8329,N_1283);
nand U16584 (N_16584,N_6406,N_8043);
and U16585 (N_16585,N_9548,N_652);
or U16586 (N_16586,N_7279,N_4914);
xor U16587 (N_16587,N_4356,N_331);
xnor U16588 (N_16588,N_4556,N_1803);
nor U16589 (N_16589,N_814,N_9361);
nor U16590 (N_16590,N_7422,N_9987);
xor U16591 (N_16591,N_6526,N_6125);
xor U16592 (N_16592,N_3856,N_5869);
nand U16593 (N_16593,N_3085,N_5240);
or U16594 (N_16594,N_8526,N_8266);
xnor U16595 (N_16595,N_5680,N_9623);
xor U16596 (N_16596,N_1781,N_6659);
xnor U16597 (N_16597,N_3767,N_3207);
nor U16598 (N_16598,N_2396,N_1956);
or U16599 (N_16599,N_6414,N_9646);
nand U16600 (N_16600,N_134,N_9320);
xor U16601 (N_16601,N_6643,N_7160);
and U16602 (N_16602,N_9423,N_8574);
and U16603 (N_16603,N_2507,N_7965);
xor U16604 (N_16604,N_371,N_4839);
nor U16605 (N_16605,N_3809,N_532);
and U16606 (N_16606,N_6227,N_2008);
or U16607 (N_16607,N_4023,N_6073);
xnor U16608 (N_16608,N_4513,N_4433);
or U16609 (N_16609,N_7317,N_1153);
xnor U16610 (N_16610,N_2552,N_7990);
xnor U16611 (N_16611,N_9673,N_8269);
and U16612 (N_16612,N_1374,N_7029);
nor U16613 (N_16613,N_867,N_6442);
or U16614 (N_16614,N_9285,N_6184);
nand U16615 (N_16615,N_5526,N_2581);
nor U16616 (N_16616,N_189,N_1160);
xnor U16617 (N_16617,N_6442,N_5234);
xor U16618 (N_16618,N_7720,N_9072);
and U16619 (N_16619,N_3144,N_8906);
xor U16620 (N_16620,N_5073,N_6224);
nor U16621 (N_16621,N_763,N_4035);
and U16622 (N_16622,N_4591,N_881);
nand U16623 (N_16623,N_3163,N_2236);
and U16624 (N_16624,N_6803,N_7343);
or U16625 (N_16625,N_828,N_8936);
or U16626 (N_16626,N_6500,N_3105);
or U16627 (N_16627,N_4338,N_384);
or U16628 (N_16628,N_7600,N_1512);
and U16629 (N_16629,N_5935,N_4550);
nor U16630 (N_16630,N_305,N_9720);
nor U16631 (N_16631,N_4110,N_6405);
xor U16632 (N_16632,N_8451,N_8210);
and U16633 (N_16633,N_9176,N_6911);
xor U16634 (N_16634,N_5391,N_6796);
nand U16635 (N_16635,N_9637,N_9150);
nor U16636 (N_16636,N_8740,N_518);
or U16637 (N_16637,N_4109,N_3735);
nand U16638 (N_16638,N_4509,N_5976);
nor U16639 (N_16639,N_695,N_2145);
nand U16640 (N_16640,N_755,N_3128);
nor U16641 (N_16641,N_9707,N_9716);
and U16642 (N_16642,N_4912,N_4560);
nand U16643 (N_16643,N_2679,N_4567);
and U16644 (N_16644,N_718,N_1665);
xor U16645 (N_16645,N_131,N_5582);
nand U16646 (N_16646,N_2739,N_8005);
xnor U16647 (N_16647,N_7268,N_8996);
nand U16648 (N_16648,N_7875,N_3030);
and U16649 (N_16649,N_4634,N_1007);
nand U16650 (N_16650,N_7626,N_1615);
nand U16651 (N_16651,N_6153,N_5080);
nor U16652 (N_16652,N_3874,N_575);
nor U16653 (N_16653,N_1953,N_6754);
or U16654 (N_16654,N_2342,N_6657);
or U16655 (N_16655,N_9424,N_4927);
nand U16656 (N_16656,N_1530,N_4348);
or U16657 (N_16657,N_3234,N_4422);
and U16658 (N_16658,N_1587,N_2309);
or U16659 (N_16659,N_7133,N_2032);
and U16660 (N_16660,N_472,N_7959);
xor U16661 (N_16661,N_2147,N_6029);
xor U16662 (N_16662,N_3689,N_8687);
xor U16663 (N_16663,N_2782,N_48);
and U16664 (N_16664,N_4250,N_6764);
xor U16665 (N_16665,N_8778,N_6782);
nor U16666 (N_16666,N_7614,N_9995);
and U16667 (N_16667,N_2114,N_8072);
or U16668 (N_16668,N_9235,N_9097);
nor U16669 (N_16669,N_6172,N_794);
xnor U16670 (N_16670,N_211,N_7433);
nand U16671 (N_16671,N_7467,N_3804);
or U16672 (N_16672,N_8282,N_4915);
nor U16673 (N_16673,N_5279,N_6683);
and U16674 (N_16674,N_6736,N_7730);
xnor U16675 (N_16675,N_3340,N_8353);
and U16676 (N_16676,N_4843,N_6286);
or U16677 (N_16677,N_9859,N_7917);
xor U16678 (N_16678,N_9351,N_9366);
nor U16679 (N_16679,N_989,N_8478);
and U16680 (N_16680,N_4640,N_3005);
xnor U16681 (N_16681,N_1220,N_347);
and U16682 (N_16682,N_76,N_7710);
or U16683 (N_16683,N_9726,N_3397);
and U16684 (N_16684,N_8976,N_940);
and U16685 (N_16685,N_6856,N_6398);
or U16686 (N_16686,N_7082,N_3612);
and U16687 (N_16687,N_8766,N_5599);
nor U16688 (N_16688,N_5006,N_8161);
xnor U16689 (N_16689,N_7646,N_2308);
xor U16690 (N_16690,N_7560,N_2223);
nor U16691 (N_16691,N_9996,N_6021);
and U16692 (N_16692,N_3396,N_6190);
xor U16693 (N_16693,N_5367,N_760);
or U16694 (N_16694,N_593,N_9835);
xnor U16695 (N_16695,N_1682,N_2762);
xnor U16696 (N_16696,N_12,N_3328);
nand U16697 (N_16697,N_8865,N_4989);
nand U16698 (N_16698,N_191,N_676);
xor U16699 (N_16699,N_7860,N_5450);
xnor U16700 (N_16700,N_906,N_540);
nor U16701 (N_16701,N_9232,N_1206);
or U16702 (N_16702,N_3765,N_8790);
nor U16703 (N_16703,N_6011,N_8350);
and U16704 (N_16704,N_8846,N_6897);
nand U16705 (N_16705,N_1597,N_2019);
xor U16706 (N_16706,N_6392,N_4947);
xor U16707 (N_16707,N_4178,N_2499);
or U16708 (N_16708,N_5707,N_6119);
or U16709 (N_16709,N_1547,N_4069);
nand U16710 (N_16710,N_7567,N_3740);
xor U16711 (N_16711,N_7831,N_8778);
xor U16712 (N_16712,N_5558,N_9380);
xor U16713 (N_16713,N_3575,N_5743);
nand U16714 (N_16714,N_5349,N_1999);
xor U16715 (N_16715,N_4988,N_7702);
xnor U16716 (N_16716,N_3013,N_1731);
or U16717 (N_16717,N_2638,N_409);
nand U16718 (N_16718,N_2033,N_5968);
nor U16719 (N_16719,N_4541,N_276);
nor U16720 (N_16720,N_2937,N_8992);
and U16721 (N_16721,N_2752,N_6104);
xor U16722 (N_16722,N_5156,N_8013);
and U16723 (N_16723,N_1072,N_9039);
or U16724 (N_16724,N_653,N_7996);
xnor U16725 (N_16725,N_6002,N_3410);
or U16726 (N_16726,N_7336,N_9272);
xor U16727 (N_16727,N_7470,N_27);
nand U16728 (N_16728,N_5081,N_4855);
nor U16729 (N_16729,N_3532,N_5192);
xor U16730 (N_16730,N_8462,N_8835);
and U16731 (N_16731,N_4571,N_5482);
or U16732 (N_16732,N_247,N_537);
xnor U16733 (N_16733,N_8192,N_312);
xnor U16734 (N_16734,N_235,N_7305);
nor U16735 (N_16735,N_5985,N_3452);
and U16736 (N_16736,N_9248,N_4519);
nor U16737 (N_16737,N_3496,N_183);
nand U16738 (N_16738,N_8095,N_9682);
xor U16739 (N_16739,N_4688,N_7854);
and U16740 (N_16740,N_4482,N_440);
and U16741 (N_16741,N_6856,N_4506);
nand U16742 (N_16742,N_7849,N_3666);
and U16743 (N_16743,N_2899,N_2648);
nor U16744 (N_16744,N_1677,N_8600);
nand U16745 (N_16745,N_9613,N_406);
or U16746 (N_16746,N_7789,N_2906);
xor U16747 (N_16747,N_4995,N_7723);
or U16748 (N_16748,N_768,N_8083);
nand U16749 (N_16749,N_8843,N_900);
or U16750 (N_16750,N_6603,N_7132);
and U16751 (N_16751,N_648,N_4144);
nand U16752 (N_16752,N_3400,N_9556);
or U16753 (N_16753,N_3964,N_4917);
xor U16754 (N_16754,N_5528,N_5210);
nand U16755 (N_16755,N_6055,N_6215);
or U16756 (N_16756,N_6131,N_6132);
nand U16757 (N_16757,N_6874,N_5114);
and U16758 (N_16758,N_6142,N_5801);
and U16759 (N_16759,N_5387,N_8655);
nand U16760 (N_16760,N_6986,N_3863);
and U16761 (N_16761,N_9741,N_8000);
or U16762 (N_16762,N_4603,N_464);
nand U16763 (N_16763,N_4859,N_7119);
xnor U16764 (N_16764,N_2368,N_8374);
xnor U16765 (N_16765,N_1653,N_824);
or U16766 (N_16766,N_8939,N_3643);
xor U16767 (N_16767,N_4997,N_615);
nand U16768 (N_16768,N_820,N_1434);
nor U16769 (N_16769,N_4843,N_1230);
or U16770 (N_16770,N_4209,N_7942);
xnor U16771 (N_16771,N_9132,N_2954);
and U16772 (N_16772,N_3699,N_1617);
xnor U16773 (N_16773,N_9844,N_1630);
or U16774 (N_16774,N_6734,N_2478);
nand U16775 (N_16775,N_2373,N_6994);
and U16776 (N_16776,N_2854,N_2918);
nor U16777 (N_16777,N_27,N_3148);
xnor U16778 (N_16778,N_6740,N_7375);
nor U16779 (N_16779,N_5252,N_3329);
nor U16780 (N_16780,N_867,N_5205);
nand U16781 (N_16781,N_6254,N_5206);
nor U16782 (N_16782,N_5337,N_7385);
xnor U16783 (N_16783,N_7245,N_2019);
or U16784 (N_16784,N_5645,N_4997);
or U16785 (N_16785,N_3670,N_3765);
or U16786 (N_16786,N_9065,N_443);
nor U16787 (N_16787,N_5450,N_5359);
xor U16788 (N_16788,N_129,N_7771);
or U16789 (N_16789,N_5653,N_4872);
nor U16790 (N_16790,N_835,N_3388);
and U16791 (N_16791,N_793,N_9110);
nor U16792 (N_16792,N_3419,N_9519);
nor U16793 (N_16793,N_7582,N_6264);
or U16794 (N_16794,N_278,N_7482);
nand U16795 (N_16795,N_9488,N_5010);
xnor U16796 (N_16796,N_9934,N_2414);
nand U16797 (N_16797,N_8732,N_7123);
or U16798 (N_16798,N_4804,N_2620);
xor U16799 (N_16799,N_9709,N_3299);
nor U16800 (N_16800,N_8157,N_2170);
or U16801 (N_16801,N_4508,N_5024);
and U16802 (N_16802,N_1497,N_9314);
xnor U16803 (N_16803,N_8518,N_2093);
and U16804 (N_16804,N_5471,N_6190);
nor U16805 (N_16805,N_576,N_9625);
nor U16806 (N_16806,N_203,N_3714);
or U16807 (N_16807,N_6921,N_8294);
nor U16808 (N_16808,N_913,N_3190);
nand U16809 (N_16809,N_1085,N_7045);
nand U16810 (N_16810,N_721,N_1930);
xor U16811 (N_16811,N_5383,N_7163);
nor U16812 (N_16812,N_1210,N_1079);
xor U16813 (N_16813,N_1918,N_6024);
nor U16814 (N_16814,N_2822,N_4782);
or U16815 (N_16815,N_6224,N_5352);
and U16816 (N_16816,N_3525,N_9414);
xor U16817 (N_16817,N_8704,N_4759);
and U16818 (N_16818,N_7313,N_6843);
and U16819 (N_16819,N_4464,N_3519);
and U16820 (N_16820,N_3507,N_985);
nor U16821 (N_16821,N_4180,N_7150);
xnor U16822 (N_16822,N_6138,N_2331);
and U16823 (N_16823,N_8411,N_3050);
xnor U16824 (N_16824,N_7804,N_8286);
or U16825 (N_16825,N_6657,N_2845);
or U16826 (N_16826,N_5317,N_1605);
or U16827 (N_16827,N_2030,N_7366);
or U16828 (N_16828,N_2155,N_4768);
and U16829 (N_16829,N_3417,N_8803);
and U16830 (N_16830,N_859,N_3965);
xnor U16831 (N_16831,N_1906,N_7258);
and U16832 (N_16832,N_4780,N_969);
xor U16833 (N_16833,N_314,N_554);
nor U16834 (N_16834,N_8457,N_1391);
or U16835 (N_16835,N_1002,N_9976);
xor U16836 (N_16836,N_4812,N_5254);
xnor U16837 (N_16837,N_3225,N_2016);
or U16838 (N_16838,N_972,N_4402);
nor U16839 (N_16839,N_7671,N_5210);
nor U16840 (N_16840,N_3795,N_6838);
xor U16841 (N_16841,N_8884,N_164);
xor U16842 (N_16842,N_3907,N_2387);
nor U16843 (N_16843,N_1327,N_2980);
xor U16844 (N_16844,N_6879,N_7899);
and U16845 (N_16845,N_5481,N_7630);
and U16846 (N_16846,N_8646,N_4280);
nor U16847 (N_16847,N_3370,N_8140);
or U16848 (N_16848,N_5235,N_3228);
xnor U16849 (N_16849,N_9795,N_6958);
and U16850 (N_16850,N_496,N_7994);
and U16851 (N_16851,N_5904,N_9264);
and U16852 (N_16852,N_530,N_7128);
or U16853 (N_16853,N_1010,N_3067);
xnor U16854 (N_16854,N_8557,N_8635);
or U16855 (N_16855,N_2878,N_8023);
xnor U16856 (N_16856,N_7315,N_4354);
and U16857 (N_16857,N_8916,N_1232);
xor U16858 (N_16858,N_4188,N_3376);
nor U16859 (N_16859,N_3975,N_2783);
nand U16860 (N_16860,N_9290,N_2320);
xor U16861 (N_16861,N_4941,N_4730);
and U16862 (N_16862,N_4627,N_3751);
nor U16863 (N_16863,N_3207,N_8997);
nand U16864 (N_16864,N_623,N_4400);
nor U16865 (N_16865,N_818,N_4617);
and U16866 (N_16866,N_1687,N_1896);
nor U16867 (N_16867,N_9818,N_2022);
nand U16868 (N_16868,N_614,N_555);
and U16869 (N_16869,N_5564,N_9280);
xnor U16870 (N_16870,N_9500,N_8542);
and U16871 (N_16871,N_1166,N_7596);
nor U16872 (N_16872,N_6825,N_9231);
and U16873 (N_16873,N_4311,N_5817);
xor U16874 (N_16874,N_1152,N_1087);
and U16875 (N_16875,N_7350,N_7266);
nand U16876 (N_16876,N_1034,N_4251);
xor U16877 (N_16877,N_5634,N_5998);
nor U16878 (N_16878,N_1472,N_6055);
xnor U16879 (N_16879,N_4764,N_3832);
and U16880 (N_16880,N_8365,N_4007);
or U16881 (N_16881,N_3955,N_3434);
nor U16882 (N_16882,N_7689,N_2504);
xor U16883 (N_16883,N_9850,N_117);
and U16884 (N_16884,N_5020,N_1721);
xor U16885 (N_16885,N_2402,N_2834);
and U16886 (N_16886,N_296,N_7836);
or U16887 (N_16887,N_256,N_8538);
or U16888 (N_16888,N_8913,N_1891);
and U16889 (N_16889,N_8325,N_9252);
nand U16890 (N_16890,N_8822,N_4667);
nor U16891 (N_16891,N_9010,N_6576);
or U16892 (N_16892,N_1074,N_6978);
nand U16893 (N_16893,N_2203,N_8137);
or U16894 (N_16894,N_2147,N_8230);
or U16895 (N_16895,N_7988,N_7623);
or U16896 (N_16896,N_2767,N_110);
nand U16897 (N_16897,N_9666,N_5455);
and U16898 (N_16898,N_5670,N_6413);
or U16899 (N_16899,N_4177,N_8767);
xor U16900 (N_16900,N_9278,N_4958);
or U16901 (N_16901,N_7561,N_5686);
and U16902 (N_16902,N_5423,N_7900);
or U16903 (N_16903,N_1237,N_1715);
or U16904 (N_16904,N_2331,N_5336);
nor U16905 (N_16905,N_7406,N_442);
xor U16906 (N_16906,N_7020,N_6124);
nand U16907 (N_16907,N_8905,N_5225);
and U16908 (N_16908,N_4291,N_4665);
or U16909 (N_16909,N_4730,N_2161);
or U16910 (N_16910,N_1244,N_9007);
nor U16911 (N_16911,N_9532,N_1932);
xnor U16912 (N_16912,N_6548,N_4855);
and U16913 (N_16913,N_454,N_304);
and U16914 (N_16914,N_9234,N_1121);
or U16915 (N_16915,N_9172,N_9157);
nand U16916 (N_16916,N_5907,N_5489);
nand U16917 (N_16917,N_5376,N_1524);
or U16918 (N_16918,N_29,N_8016);
and U16919 (N_16919,N_5358,N_6999);
and U16920 (N_16920,N_1627,N_79);
or U16921 (N_16921,N_6493,N_180);
xnor U16922 (N_16922,N_4711,N_325);
nor U16923 (N_16923,N_7848,N_3714);
and U16924 (N_16924,N_7282,N_5038);
nand U16925 (N_16925,N_8584,N_3919);
and U16926 (N_16926,N_2010,N_3410);
nor U16927 (N_16927,N_6014,N_5173);
nand U16928 (N_16928,N_9933,N_8802);
or U16929 (N_16929,N_7098,N_3939);
nor U16930 (N_16930,N_9083,N_5364);
and U16931 (N_16931,N_7423,N_3376);
or U16932 (N_16932,N_8145,N_1984);
nor U16933 (N_16933,N_9451,N_2864);
and U16934 (N_16934,N_1859,N_7084);
and U16935 (N_16935,N_784,N_9458);
nor U16936 (N_16936,N_3311,N_8167);
and U16937 (N_16937,N_8900,N_9707);
nor U16938 (N_16938,N_5084,N_9230);
nand U16939 (N_16939,N_8786,N_276);
xor U16940 (N_16940,N_8832,N_4632);
and U16941 (N_16941,N_9018,N_2799);
or U16942 (N_16942,N_4263,N_6743);
nand U16943 (N_16943,N_801,N_592);
or U16944 (N_16944,N_3035,N_6353);
and U16945 (N_16945,N_8522,N_7757);
or U16946 (N_16946,N_9967,N_2784);
nor U16947 (N_16947,N_1337,N_8158);
nand U16948 (N_16948,N_2355,N_5728);
nor U16949 (N_16949,N_464,N_4693);
or U16950 (N_16950,N_3026,N_3489);
and U16951 (N_16951,N_6513,N_9421);
xor U16952 (N_16952,N_4952,N_3983);
xor U16953 (N_16953,N_1337,N_7131);
nand U16954 (N_16954,N_7813,N_5726);
or U16955 (N_16955,N_5831,N_112);
or U16956 (N_16956,N_9051,N_9185);
xor U16957 (N_16957,N_6745,N_1424);
nand U16958 (N_16958,N_3549,N_8840);
nand U16959 (N_16959,N_1660,N_4837);
or U16960 (N_16960,N_2385,N_257);
and U16961 (N_16961,N_1004,N_1919);
or U16962 (N_16962,N_5168,N_5300);
xor U16963 (N_16963,N_5693,N_5480);
or U16964 (N_16964,N_271,N_8541);
xor U16965 (N_16965,N_8760,N_5523);
or U16966 (N_16966,N_2220,N_5096);
nand U16967 (N_16967,N_9256,N_6041);
xnor U16968 (N_16968,N_1064,N_178);
nor U16969 (N_16969,N_2294,N_3823);
xor U16970 (N_16970,N_7311,N_4855);
xor U16971 (N_16971,N_2959,N_4822);
nand U16972 (N_16972,N_128,N_9511);
nand U16973 (N_16973,N_6130,N_9396);
nand U16974 (N_16974,N_1277,N_8919);
nor U16975 (N_16975,N_9053,N_2893);
xnor U16976 (N_16976,N_4233,N_9847);
xor U16977 (N_16977,N_8598,N_3848);
nor U16978 (N_16978,N_7068,N_9556);
and U16979 (N_16979,N_4045,N_5627);
nand U16980 (N_16980,N_4638,N_3445);
xnor U16981 (N_16981,N_8107,N_7282);
and U16982 (N_16982,N_2868,N_5449);
xnor U16983 (N_16983,N_9113,N_7921);
nand U16984 (N_16984,N_187,N_8833);
nor U16985 (N_16985,N_6038,N_862);
xor U16986 (N_16986,N_2445,N_8244);
and U16987 (N_16987,N_2055,N_1445);
and U16988 (N_16988,N_9868,N_9085);
xor U16989 (N_16989,N_9170,N_7509);
xor U16990 (N_16990,N_6435,N_2926);
and U16991 (N_16991,N_9452,N_9572);
and U16992 (N_16992,N_2782,N_9518);
and U16993 (N_16993,N_2634,N_8488);
nor U16994 (N_16994,N_3426,N_6159);
xor U16995 (N_16995,N_641,N_195);
nand U16996 (N_16996,N_7580,N_7076);
nor U16997 (N_16997,N_2237,N_3569);
xnor U16998 (N_16998,N_7311,N_2563);
and U16999 (N_16999,N_3758,N_1177);
nand U17000 (N_17000,N_2691,N_6837);
xor U17001 (N_17001,N_5483,N_3345);
and U17002 (N_17002,N_4046,N_9898);
nand U17003 (N_17003,N_8424,N_3323);
xor U17004 (N_17004,N_1841,N_6437);
nand U17005 (N_17005,N_7285,N_9291);
xor U17006 (N_17006,N_7964,N_4980);
nor U17007 (N_17007,N_6163,N_6312);
nand U17008 (N_17008,N_6744,N_1082);
and U17009 (N_17009,N_135,N_8964);
nand U17010 (N_17010,N_3933,N_1904);
or U17011 (N_17011,N_5348,N_3470);
xnor U17012 (N_17012,N_537,N_3053);
or U17013 (N_17013,N_7001,N_4814);
and U17014 (N_17014,N_8911,N_8515);
xor U17015 (N_17015,N_4008,N_261);
nor U17016 (N_17016,N_4072,N_5563);
nand U17017 (N_17017,N_1396,N_490);
nor U17018 (N_17018,N_7413,N_271);
nor U17019 (N_17019,N_9467,N_7802);
and U17020 (N_17020,N_7829,N_743);
nor U17021 (N_17021,N_4397,N_1623);
or U17022 (N_17022,N_292,N_9391);
nor U17023 (N_17023,N_4503,N_6219);
nand U17024 (N_17024,N_7613,N_8078);
nand U17025 (N_17025,N_1302,N_438);
xor U17026 (N_17026,N_6256,N_6794);
xor U17027 (N_17027,N_4374,N_6094);
xnor U17028 (N_17028,N_6754,N_3664);
xor U17029 (N_17029,N_5552,N_1649);
xor U17030 (N_17030,N_8285,N_1505);
or U17031 (N_17031,N_8109,N_2630);
nor U17032 (N_17032,N_1331,N_1251);
nor U17033 (N_17033,N_2966,N_3948);
nor U17034 (N_17034,N_7924,N_101);
xnor U17035 (N_17035,N_5755,N_3032);
and U17036 (N_17036,N_6853,N_6433);
or U17037 (N_17037,N_1208,N_2149);
xor U17038 (N_17038,N_2520,N_7830);
or U17039 (N_17039,N_1385,N_2355);
or U17040 (N_17040,N_1798,N_4890);
xor U17041 (N_17041,N_9520,N_2257);
and U17042 (N_17042,N_6874,N_5393);
nand U17043 (N_17043,N_3605,N_7969);
and U17044 (N_17044,N_8141,N_8964);
xnor U17045 (N_17045,N_565,N_8749);
nand U17046 (N_17046,N_3072,N_794);
or U17047 (N_17047,N_3818,N_4879);
nand U17048 (N_17048,N_7907,N_3895);
and U17049 (N_17049,N_1529,N_9295);
nor U17050 (N_17050,N_694,N_274);
and U17051 (N_17051,N_4884,N_208);
xnor U17052 (N_17052,N_124,N_2763);
nor U17053 (N_17053,N_4570,N_358);
xnor U17054 (N_17054,N_8988,N_4002);
nor U17055 (N_17055,N_4343,N_7022);
and U17056 (N_17056,N_7600,N_5518);
nand U17057 (N_17057,N_6701,N_5659);
nand U17058 (N_17058,N_4556,N_8597);
or U17059 (N_17059,N_5402,N_4137);
and U17060 (N_17060,N_3534,N_6416);
or U17061 (N_17061,N_868,N_5335);
or U17062 (N_17062,N_4476,N_6627);
nor U17063 (N_17063,N_6386,N_9163);
and U17064 (N_17064,N_218,N_3632);
or U17065 (N_17065,N_395,N_2338);
nand U17066 (N_17066,N_7480,N_4946);
nor U17067 (N_17067,N_1080,N_3349);
or U17068 (N_17068,N_1090,N_7348);
xnor U17069 (N_17069,N_2780,N_3652);
xor U17070 (N_17070,N_2122,N_3452);
or U17071 (N_17071,N_5602,N_4598);
nand U17072 (N_17072,N_280,N_633);
or U17073 (N_17073,N_3321,N_420);
or U17074 (N_17074,N_1714,N_4466);
nor U17075 (N_17075,N_6985,N_4778);
xor U17076 (N_17076,N_6763,N_2621);
or U17077 (N_17077,N_9078,N_7381);
xor U17078 (N_17078,N_605,N_3610);
xnor U17079 (N_17079,N_3034,N_1334);
xor U17080 (N_17080,N_7411,N_1626);
nand U17081 (N_17081,N_1263,N_1683);
or U17082 (N_17082,N_2457,N_2127);
and U17083 (N_17083,N_5285,N_4268);
and U17084 (N_17084,N_2240,N_1906);
and U17085 (N_17085,N_6506,N_8875);
and U17086 (N_17086,N_7598,N_8033);
nand U17087 (N_17087,N_9662,N_4603);
or U17088 (N_17088,N_9407,N_2259);
nor U17089 (N_17089,N_2618,N_2165);
nand U17090 (N_17090,N_783,N_3480);
or U17091 (N_17091,N_975,N_1482);
nand U17092 (N_17092,N_3336,N_423);
and U17093 (N_17093,N_673,N_2649);
nor U17094 (N_17094,N_4263,N_7796);
and U17095 (N_17095,N_7197,N_9743);
or U17096 (N_17096,N_6131,N_7418);
nor U17097 (N_17097,N_8748,N_7380);
xnor U17098 (N_17098,N_1543,N_6608);
nand U17099 (N_17099,N_4307,N_2676);
nor U17100 (N_17100,N_183,N_6278);
or U17101 (N_17101,N_1031,N_2621);
nand U17102 (N_17102,N_876,N_2994);
xnor U17103 (N_17103,N_6024,N_417);
and U17104 (N_17104,N_1762,N_5667);
nor U17105 (N_17105,N_4370,N_1502);
xor U17106 (N_17106,N_9577,N_6407);
nand U17107 (N_17107,N_2209,N_4848);
nand U17108 (N_17108,N_6988,N_4503);
nor U17109 (N_17109,N_5939,N_6919);
xnor U17110 (N_17110,N_3513,N_622);
and U17111 (N_17111,N_9907,N_5737);
nor U17112 (N_17112,N_9914,N_6591);
or U17113 (N_17113,N_7029,N_1759);
and U17114 (N_17114,N_4049,N_56);
nand U17115 (N_17115,N_5925,N_91);
and U17116 (N_17116,N_6690,N_4405);
xnor U17117 (N_17117,N_4599,N_5387);
xnor U17118 (N_17118,N_4019,N_8249);
or U17119 (N_17119,N_3844,N_5966);
xor U17120 (N_17120,N_1214,N_2902);
xor U17121 (N_17121,N_4130,N_5208);
nor U17122 (N_17122,N_1231,N_1274);
and U17123 (N_17123,N_6535,N_3662);
and U17124 (N_17124,N_1396,N_8724);
or U17125 (N_17125,N_5329,N_1124);
nor U17126 (N_17126,N_8652,N_1592);
xor U17127 (N_17127,N_1408,N_9876);
nor U17128 (N_17128,N_743,N_8575);
and U17129 (N_17129,N_9396,N_7682);
nand U17130 (N_17130,N_5788,N_290);
xor U17131 (N_17131,N_6522,N_410);
nand U17132 (N_17132,N_6080,N_9784);
nor U17133 (N_17133,N_3597,N_1012);
xnor U17134 (N_17134,N_1134,N_7006);
nand U17135 (N_17135,N_2159,N_8082);
xor U17136 (N_17136,N_7888,N_3594);
nand U17137 (N_17137,N_3350,N_5584);
nand U17138 (N_17138,N_5982,N_7681);
nor U17139 (N_17139,N_1952,N_4097);
xor U17140 (N_17140,N_820,N_9053);
nor U17141 (N_17141,N_1998,N_6197);
nor U17142 (N_17142,N_6764,N_3322);
or U17143 (N_17143,N_1114,N_8379);
and U17144 (N_17144,N_6600,N_3399);
nand U17145 (N_17145,N_1065,N_5301);
xnor U17146 (N_17146,N_2227,N_9679);
xor U17147 (N_17147,N_400,N_1424);
or U17148 (N_17148,N_7907,N_6563);
and U17149 (N_17149,N_9736,N_9059);
or U17150 (N_17150,N_1426,N_6789);
and U17151 (N_17151,N_7652,N_8411);
nor U17152 (N_17152,N_9407,N_3756);
nand U17153 (N_17153,N_6936,N_5404);
nand U17154 (N_17154,N_607,N_3906);
nor U17155 (N_17155,N_4289,N_9248);
nor U17156 (N_17156,N_1215,N_4718);
nor U17157 (N_17157,N_4652,N_3174);
nor U17158 (N_17158,N_3828,N_2996);
or U17159 (N_17159,N_7730,N_5628);
nand U17160 (N_17160,N_3415,N_2806);
nor U17161 (N_17161,N_6289,N_8025);
or U17162 (N_17162,N_3244,N_6357);
or U17163 (N_17163,N_4298,N_7124);
xor U17164 (N_17164,N_882,N_8077);
and U17165 (N_17165,N_8133,N_8900);
nand U17166 (N_17166,N_4499,N_1499);
xor U17167 (N_17167,N_9966,N_1673);
or U17168 (N_17168,N_2331,N_2295);
nand U17169 (N_17169,N_1160,N_9376);
nor U17170 (N_17170,N_5352,N_923);
nand U17171 (N_17171,N_8074,N_3930);
nor U17172 (N_17172,N_2162,N_56);
nand U17173 (N_17173,N_4537,N_1528);
xnor U17174 (N_17174,N_2629,N_5628);
nor U17175 (N_17175,N_1531,N_8813);
or U17176 (N_17176,N_6595,N_448);
xor U17177 (N_17177,N_3943,N_7903);
nor U17178 (N_17178,N_5857,N_1342);
and U17179 (N_17179,N_3209,N_9021);
nand U17180 (N_17180,N_3983,N_6975);
nand U17181 (N_17181,N_6614,N_5861);
nand U17182 (N_17182,N_3052,N_5099);
or U17183 (N_17183,N_5125,N_1097);
xnor U17184 (N_17184,N_3828,N_170);
and U17185 (N_17185,N_9879,N_3190);
or U17186 (N_17186,N_5662,N_4712);
xor U17187 (N_17187,N_2661,N_5313);
and U17188 (N_17188,N_2371,N_922);
nor U17189 (N_17189,N_3150,N_6881);
xor U17190 (N_17190,N_5430,N_3523);
and U17191 (N_17191,N_5194,N_5823);
or U17192 (N_17192,N_1945,N_8276);
nor U17193 (N_17193,N_9586,N_7793);
and U17194 (N_17194,N_5939,N_3724);
and U17195 (N_17195,N_6013,N_1246);
xor U17196 (N_17196,N_7425,N_2690);
or U17197 (N_17197,N_3566,N_1195);
or U17198 (N_17198,N_1963,N_6399);
nor U17199 (N_17199,N_38,N_844);
and U17200 (N_17200,N_7982,N_6850);
nand U17201 (N_17201,N_7440,N_7770);
or U17202 (N_17202,N_4922,N_9908);
nand U17203 (N_17203,N_5696,N_4185);
nor U17204 (N_17204,N_7847,N_9496);
and U17205 (N_17205,N_2104,N_3605);
nand U17206 (N_17206,N_1318,N_9628);
and U17207 (N_17207,N_4298,N_3930);
nor U17208 (N_17208,N_4093,N_1330);
or U17209 (N_17209,N_6661,N_3500);
nor U17210 (N_17210,N_4314,N_5788);
or U17211 (N_17211,N_4804,N_8454);
nor U17212 (N_17212,N_1827,N_7513);
nand U17213 (N_17213,N_859,N_4459);
xnor U17214 (N_17214,N_6292,N_3811);
nand U17215 (N_17215,N_1324,N_5085);
nor U17216 (N_17216,N_8081,N_978);
xnor U17217 (N_17217,N_2131,N_5062);
or U17218 (N_17218,N_2882,N_6305);
and U17219 (N_17219,N_5707,N_7119);
xor U17220 (N_17220,N_2964,N_9476);
nand U17221 (N_17221,N_1582,N_7362);
nor U17222 (N_17222,N_4006,N_7715);
nand U17223 (N_17223,N_1007,N_2644);
or U17224 (N_17224,N_2035,N_5691);
and U17225 (N_17225,N_7891,N_2996);
nand U17226 (N_17226,N_5050,N_4920);
or U17227 (N_17227,N_5679,N_6967);
and U17228 (N_17228,N_4722,N_6508);
and U17229 (N_17229,N_5345,N_7663);
or U17230 (N_17230,N_683,N_6784);
xnor U17231 (N_17231,N_6848,N_27);
nor U17232 (N_17232,N_1434,N_8059);
nand U17233 (N_17233,N_2141,N_387);
nor U17234 (N_17234,N_4219,N_5438);
and U17235 (N_17235,N_9046,N_9765);
nand U17236 (N_17236,N_2137,N_3223);
or U17237 (N_17237,N_9518,N_2593);
nor U17238 (N_17238,N_1098,N_6958);
nor U17239 (N_17239,N_2885,N_2227);
nand U17240 (N_17240,N_4566,N_4716);
and U17241 (N_17241,N_3476,N_1642);
or U17242 (N_17242,N_5263,N_931);
nor U17243 (N_17243,N_8286,N_5006);
xnor U17244 (N_17244,N_9901,N_9929);
or U17245 (N_17245,N_9732,N_7057);
nand U17246 (N_17246,N_2839,N_363);
nand U17247 (N_17247,N_6251,N_4907);
or U17248 (N_17248,N_8019,N_6941);
nand U17249 (N_17249,N_3794,N_1548);
nor U17250 (N_17250,N_5025,N_2082);
or U17251 (N_17251,N_3331,N_7012);
or U17252 (N_17252,N_9786,N_1130);
or U17253 (N_17253,N_9569,N_3865);
nor U17254 (N_17254,N_4952,N_2594);
and U17255 (N_17255,N_8478,N_7103);
nand U17256 (N_17256,N_4738,N_1699);
nand U17257 (N_17257,N_2942,N_9948);
nand U17258 (N_17258,N_1339,N_1550);
or U17259 (N_17259,N_8526,N_94);
xnor U17260 (N_17260,N_5240,N_9808);
or U17261 (N_17261,N_8390,N_2326);
and U17262 (N_17262,N_2950,N_9684);
nand U17263 (N_17263,N_1584,N_8872);
xor U17264 (N_17264,N_5007,N_8638);
nor U17265 (N_17265,N_1354,N_925);
nand U17266 (N_17266,N_9104,N_8376);
xor U17267 (N_17267,N_3258,N_1319);
nand U17268 (N_17268,N_9908,N_182);
nand U17269 (N_17269,N_5334,N_1140);
nor U17270 (N_17270,N_3548,N_8699);
nand U17271 (N_17271,N_2025,N_5071);
xor U17272 (N_17272,N_3784,N_9276);
nand U17273 (N_17273,N_7854,N_2448);
nand U17274 (N_17274,N_8531,N_1722);
or U17275 (N_17275,N_2976,N_1528);
xor U17276 (N_17276,N_4311,N_9782);
or U17277 (N_17277,N_84,N_1954);
and U17278 (N_17278,N_2683,N_6633);
or U17279 (N_17279,N_312,N_2878);
and U17280 (N_17280,N_520,N_2017);
and U17281 (N_17281,N_721,N_4548);
xnor U17282 (N_17282,N_4989,N_249);
and U17283 (N_17283,N_5620,N_3920);
xor U17284 (N_17284,N_6582,N_5876);
nand U17285 (N_17285,N_8771,N_4135);
nor U17286 (N_17286,N_1592,N_1066);
nand U17287 (N_17287,N_3042,N_3596);
nor U17288 (N_17288,N_4005,N_7876);
xnor U17289 (N_17289,N_5104,N_2374);
nand U17290 (N_17290,N_4057,N_4182);
nor U17291 (N_17291,N_4838,N_7808);
or U17292 (N_17292,N_9753,N_6779);
xor U17293 (N_17293,N_3100,N_9042);
nand U17294 (N_17294,N_5804,N_7049);
nor U17295 (N_17295,N_6599,N_3290);
nor U17296 (N_17296,N_6454,N_9723);
nor U17297 (N_17297,N_776,N_3830);
or U17298 (N_17298,N_2506,N_9304);
nand U17299 (N_17299,N_805,N_4065);
or U17300 (N_17300,N_8547,N_2777);
nor U17301 (N_17301,N_2127,N_4676);
nor U17302 (N_17302,N_707,N_6080);
nor U17303 (N_17303,N_2858,N_7926);
nand U17304 (N_17304,N_4594,N_3625);
xnor U17305 (N_17305,N_7533,N_8360);
nand U17306 (N_17306,N_3960,N_6929);
nor U17307 (N_17307,N_9463,N_2563);
nand U17308 (N_17308,N_6857,N_8462);
nor U17309 (N_17309,N_6268,N_228);
and U17310 (N_17310,N_2281,N_6476);
nand U17311 (N_17311,N_625,N_6682);
xor U17312 (N_17312,N_1999,N_7508);
xor U17313 (N_17313,N_3068,N_4);
or U17314 (N_17314,N_5254,N_540);
nor U17315 (N_17315,N_5869,N_1940);
xnor U17316 (N_17316,N_6806,N_3170);
or U17317 (N_17317,N_7483,N_1061);
xor U17318 (N_17318,N_9392,N_8038);
and U17319 (N_17319,N_2406,N_6458);
nor U17320 (N_17320,N_4371,N_9406);
or U17321 (N_17321,N_994,N_1625);
xnor U17322 (N_17322,N_7251,N_7503);
xnor U17323 (N_17323,N_983,N_5635);
or U17324 (N_17324,N_8294,N_6298);
nor U17325 (N_17325,N_7096,N_5103);
and U17326 (N_17326,N_7921,N_1340);
nor U17327 (N_17327,N_969,N_7735);
nor U17328 (N_17328,N_8088,N_6477);
and U17329 (N_17329,N_8722,N_5594);
nand U17330 (N_17330,N_6685,N_2541);
nand U17331 (N_17331,N_6551,N_5892);
xor U17332 (N_17332,N_8064,N_448);
nor U17333 (N_17333,N_1904,N_1647);
nor U17334 (N_17334,N_283,N_4733);
nand U17335 (N_17335,N_4847,N_5208);
and U17336 (N_17336,N_3704,N_8631);
xor U17337 (N_17337,N_6099,N_4911);
or U17338 (N_17338,N_9973,N_1374);
nand U17339 (N_17339,N_951,N_9830);
nor U17340 (N_17340,N_7661,N_8409);
nor U17341 (N_17341,N_4806,N_4844);
and U17342 (N_17342,N_8001,N_8868);
xnor U17343 (N_17343,N_5494,N_4326);
or U17344 (N_17344,N_3727,N_7174);
xnor U17345 (N_17345,N_6873,N_1021);
or U17346 (N_17346,N_1744,N_7781);
xnor U17347 (N_17347,N_4776,N_176);
and U17348 (N_17348,N_7571,N_6095);
nand U17349 (N_17349,N_6744,N_8865);
and U17350 (N_17350,N_4679,N_5611);
nor U17351 (N_17351,N_6686,N_8731);
nor U17352 (N_17352,N_7634,N_3671);
nor U17353 (N_17353,N_9114,N_681);
xor U17354 (N_17354,N_5561,N_5417);
or U17355 (N_17355,N_7350,N_9470);
or U17356 (N_17356,N_5757,N_6491);
nor U17357 (N_17357,N_4380,N_6741);
xor U17358 (N_17358,N_7487,N_2411);
xor U17359 (N_17359,N_3448,N_499);
or U17360 (N_17360,N_538,N_1685);
and U17361 (N_17361,N_3689,N_5405);
or U17362 (N_17362,N_6665,N_5111);
or U17363 (N_17363,N_5830,N_4392);
nor U17364 (N_17364,N_677,N_4796);
or U17365 (N_17365,N_1829,N_4208);
nor U17366 (N_17366,N_2082,N_1713);
and U17367 (N_17367,N_6761,N_4407);
xor U17368 (N_17368,N_1900,N_5669);
xnor U17369 (N_17369,N_9451,N_3126);
nand U17370 (N_17370,N_2285,N_826);
nor U17371 (N_17371,N_3840,N_5059);
and U17372 (N_17372,N_2551,N_3816);
or U17373 (N_17373,N_7356,N_3807);
nand U17374 (N_17374,N_8614,N_1095);
nor U17375 (N_17375,N_5442,N_9868);
nor U17376 (N_17376,N_7077,N_6517);
xor U17377 (N_17377,N_899,N_9808);
nor U17378 (N_17378,N_4659,N_4885);
nand U17379 (N_17379,N_4264,N_8960);
or U17380 (N_17380,N_1452,N_6294);
or U17381 (N_17381,N_4857,N_239);
xnor U17382 (N_17382,N_2129,N_8709);
or U17383 (N_17383,N_925,N_8549);
xor U17384 (N_17384,N_8355,N_1927);
or U17385 (N_17385,N_6337,N_1710);
nor U17386 (N_17386,N_1826,N_2548);
or U17387 (N_17387,N_856,N_9797);
nor U17388 (N_17388,N_4989,N_4060);
and U17389 (N_17389,N_5723,N_6518);
nand U17390 (N_17390,N_3228,N_8469);
and U17391 (N_17391,N_6912,N_9464);
or U17392 (N_17392,N_3226,N_3184);
nand U17393 (N_17393,N_3098,N_7373);
or U17394 (N_17394,N_1443,N_6328);
and U17395 (N_17395,N_6776,N_1045);
nand U17396 (N_17396,N_6806,N_1515);
nor U17397 (N_17397,N_4975,N_1463);
or U17398 (N_17398,N_2095,N_6749);
nor U17399 (N_17399,N_8678,N_5315);
and U17400 (N_17400,N_8414,N_6931);
nor U17401 (N_17401,N_3556,N_5713);
nor U17402 (N_17402,N_1056,N_5109);
and U17403 (N_17403,N_4479,N_4845);
nand U17404 (N_17404,N_4130,N_715);
nor U17405 (N_17405,N_1,N_9658);
nor U17406 (N_17406,N_1899,N_8928);
xor U17407 (N_17407,N_9866,N_6356);
nor U17408 (N_17408,N_8748,N_8459);
and U17409 (N_17409,N_5215,N_8690);
nand U17410 (N_17410,N_3918,N_9791);
or U17411 (N_17411,N_6793,N_6359);
xor U17412 (N_17412,N_3052,N_3763);
nor U17413 (N_17413,N_5941,N_6160);
xnor U17414 (N_17414,N_834,N_8097);
and U17415 (N_17415,N_4475,N_289);
nor U17416 (N_17416,N_949,N_9460);
and U17417 (N_17417,N_4547,N_6310);
nor U17418 (N_17418,N_5811,N_7149);
xor U17419 (N_17419,N_1753,N_5342);
or U17420 (N_17420,N_6546,N_1423);
nand U17421 (N_17421,N_5340,N_7619);
or U17422 (N_17422,N_1550,N_5317);
xor U17423 (N_17423,N_7171,N_3165);
nand U17424 (N_17424,N_2137,N_9554);
and U17425 (N_17425,N_3304,N_7684);
nor U17426 (N_17426,N_2868,N_7665);
nand U17427 (N_17427,N_754,N_3388);
or U17428 (N_17428,N_9875,N_2951);
xnor U17429 (N_17429,N_2860,N_5256);
or U17430 (N_17430,N_1844,N_1448);
nand U17431 (N_17431,N_6866,N_5960);
or U17432 (N_17432,N_7438,N_943);
nor U17433 (N_17433,N_2513,N_3998);
and U17434 (N_17434,N_3685,N_3901);
and U17435 (N_17435,N_118,N_7352);
xor U17436 (N_17436,N_4929,N_8433);
nand U17437 (N_17437,N_2855,N_14);
and U17438 (N_17438,N_6223,N_6442);
and U17439 (N_17439,N_6292,N_4277);
nand U17440 (N_17440,N_8447,N_9732);
nor U17441 (N_17441,N_4571,N_658);
xnor U17442 (N_17442,N_5774,N_7721);
nor U17443 (N_17443,N_7573,N_9293);
and U17444 (N_17444,N_6753,N_1350);
xnor U17445 (N_17445,N_6656,N_6855);
or U17446 (N_17446,N_3968,N_8622);
or U17447 (N_17447,N_2089,N_665);
or U17448 (N_17448,N_6619,N_5433);
xor U17449 (N_17449,N_8352,N_8185);
nand U17450 (N_17450,N_7067,N_4430);
and U17451 (N_17451,N_4958,N_1756);
nor U17452 (N_17452,N_3430,N_7349);
or U17453 (N_17453,N_2724,N_8348);
nand U17454 (N_17454,N_2746,N_5907);
and U17455 (N_17455,N_9186,N_3876);
nor U17456 (N_17456,N_9081,N_2198);
nand U17457 (N_17457,N_9348,N_7434);
and U17458 (N_17458,N_7887,N_3340);
and U17459 (N_17459,N_1945,N_5537);
xor U17460 (N_17460,N_4271,N_393);
and U17461 (N_17461,N_6941,N_6987);
nor U17462 (N_17462,N_5939,N_863);
or U17463 (N_17463,N_6592,N_7123);
xor U17464 (N_17464,N_7184,N_8760);
or U17465 (N_17465,N_9336,N_5790);
and U17466 (N_17466,N_9142,N_9031);
and U17467 (N_17467,N_570,N_2233);
and U17468 (N_17468,N_6169,N_8659);
or U17469 (N_17469,N_6153,N_5066);
nor U17470 (N_17470,N_15,N_383);
or U17471 (N_17471,N_221,N_119);
or U17472 (N_17472,N_6591,N_9683);
nor U17473 (N_17473,N_9963,N_3787);
nand U17474 (N_17474,N_6161,N_5663);
and U17475 (N_17475,N_6630,N_2811);
nor U17476 (N_17476,N_96,N_3858);
and U17477 (N_17477,N_9795,N_9067);
nand U17478 (N_17478,N_4783,N_7079);
nor U17479 (N_17479,N_4028,N_3567);
nor U17480 (N_17480,N_911,N_8581);
nand U17481 (N_17481,N_4645,N_8311);
xor U17482 (N_17482,N_1727,N_3851);
or U17483 (N_17483,N_8167,N_2764);
nor U17484 (N_17484,N_5279,N_932);
nand U17485 (N_17485,N_9564,N_7064);
or U17486 (N_17486,N_6178,N_6962);
and U17487 (N_17487,N_5535,N_603);
xnor U17488 (N_17488,N_9967,N_2436);
nand U17489 (N_17489,N_2336,N_1024);
and U17490 (N_17490,N_1270,N_4590);
xor U17491 (N_17491,N_22,N_5981);
or U17492 (N_17492,N_8648,N_4655);
or U17493 (N_17493,N_4787,N_4891);
nand U17494 (N_17494,N_1136,N_3050);
and U17495 (N_17495,N_7323,N_3152);
nor U17496 (N_17496,N_8603,N_1319);
nand U17497 (N_17497,N_4929,N_3518);
nand U17498 (N_17498,N_4125,N_8183);
xor U17499 (N_17499,N_4980,N_1605);
or U17500 (N_17500,N_5430,N_1524);
and U17501 (N_17501,N_1069,N_3704);
and U17502 (N_17502,N_4555,N_6624);
or U17503 (N_17503,N_3109,N_1152);
or U17504 (N_17504,N_8903,N_9369);
nand U17505 (N_17505,N_2682,N_3172);
nand U17506 (N_17506,N_4684,N_3189);
xnor U17507 (N_17507,N_1036,N_4257);
nand U17508 (N_17508,N_8192,N_5422);
nor U17509 (N_17509,N_5302,N_4299);
or U17510 (N_17510,N_1027,N_675);
xnor U17511 (N_17511,N_3754,N_8535);
and U17512 (N_17512,N_9019,N_5699);
nor U17513 (N_17513,N_2027,N_218);
or U17514 (N_17514,N_2836,N_1537);
xnor U17515 (N_17515,N_4800,N_3619);
nand U17516 (N_17516,N_3,N_5474);
nand U17517 (N_17517,N_8334,N_4433);
nand U17518 (N_17518,N_8314,N_3812);
nor U17519 (N_17519,N_46,N_4351);
xor U17520 (N_17520,N_639,N_1041);
nand U17521 (N_17521,N_6696,N_2722);
and U17522 (N_17522,N_719,N_547);
and U17523 (N_17523,N_3675,N_3934);
nand U17524 (N_17524,N_647,N_5954);
and U17525 (N_17525,N_633,N_8364);
or U17526 (N_17526,N_1328,N_3928);
nor U17527 (N_17527,N_4599,N_5198);
xor U17528 (N_17528,N_9991,N_7815);
xnor U17529 (N_17529,N_733,N_6962);
nor U17530 (N_17530,N_7837,N_6500);
nand U17531 (N_17531,N_7378,N_9654);
nand U17532 (N_17532,N_7238,N_4799);
nand U17533 (N_17533,N_461,N_4993);
and U17534 (N_17534,N_3981,N_9715);
nand U17535 (N_17535,N_2496,N_1801);
xor U17536 (N_17536,N_8616,N_7222);
or U17537 (N_17537,N_6683,N_9717);
or U17538 (N_17538,N_3566,N_8876);
nor U17539 (N_17539,N_8820,N_5734);
xnor U17540 (N_17540,N_2263,N_1186);
nor U17541 (N_17541,N_7247,N_1164);
nand U17542 (N_17542,N_1110,N_6546);
nor U17543 (N_17543,N_4520,N_6203);
nand U17544 (N_17544,N_1660,N_644);
nand U17545 (N_17545,N_9305,N_6712);
and U17546 (N_17546,N_4539,N_2808);
and U17547 (N_17547,N_104,N_7214);
and U17548 (N_17548,N_1493,N_8507);
xnor U17549 (N_17549,N_9960,N_4642);
nor U17550 (N_17550,N_2388,N_3906);
xnor U17551 (N_17551,N_7124,N_5391);
xnor U17552 (N_17552,N_7270,N_5959);
and U17553 (N_17553,N_743,N_4741);
and U17554 (N_17554,N_7035,N_2318);
nand U17555 (N_17555,N_435,N_8055);
and U17556 (N_17556,N_6545,N_3816);
nand U17557 (N_17557,N_5604,N_5313);
nand U17558 (N_17558,N_3436,N_7095);
xnor U17559 (N_17559,N_2073,N_8339);
nor U17560 (N_17560,N_8388,N_9114);
xnor U17561 (N_17561,N_6133,N_8676);
and U17562 (N_17562,N_5991,N_5160);
nand U17563 (N_17563,N_1059,N_5495);
xnor U17564 (N_17564,N_2666,N_1828);
nand U17565 (N_17565,N_4292,N_3714);
nor U17566 (N_17566,N_6109,N_1057);
or U17567 (N_17567,N_4004,N_5499);
xnor U17568 (N_17568,N_6581,N_2645);
and U17569 (N_17569,N_7820,N_9614);
xor U17570 (N_17570,N_5859,N_6923);
or U17571 (N_17571,N_3471,N_6896);
and U17572 (N_17572,N_1556,N_2397);
nor U17573 (N_17573,N_3786,N_2816);
nand U17574 (N_17574,N_6851,N_7412);
nor U17575 (N_17575,N_9248,N_9861);
nor U17576 (N_17576,N_1816,N_8576);
nor U17577 (N_17577,N_6472,N_5916);
nor U17578 (N_17578,N_656,N_1012);
and U17579 (N_17579,N_7163,N_9700);
nand U17580 (N_17580,N_1103,N_9043);
and U17581 (N_17581,N_1268,N_7191);
and U17582 (N_17582,N_8080,N_971);
nand U17583 (N_17583,N_962,N_33);
and U17584 (N_17584,N_352,N_5535);
nand U17585 (N_17585,N_7941,N_3445);
xor U17586 (N_17586,N_464,N_178);
xor U17587 (N_17587,N_4787,N_8388);
nor U17588 (N_17588,N_8659,N_5836);
or U17589 (N_17589,N_3145,N_8741);
nand U17590 (N_17590,N_8595,N_6646);
nand U17591 (N_17591,N_284,N_2358);
and U17592 (N_17592,N_5486,N_7503);
xor U17593 (N_17593,N_9525,N_649);
and U17594 (N_17594,N_2338,N_7197);
and U17595 (N_17595,N_2887,N_5552);
or U17596 (N_17596,N_6445,N_5486);
and U17597 (N_17597,N_9426,N_8383);
or U17598 (N_17598,N_1888,N_4051);
or U17599 (N_17599,N_2916,N_8631);
xnor U17600 (N_17600,N_958,N_5136);
nand U17601 (N_17601,N_8027,N_5109);
and U17602 (N_17602,N_6718,N_8548);
and U17603 (N_17603,N_5084,N_8128);
xnor U17604 (N_17604,N_5302,N_5193);
or U17605 (N_17605,N_909,N_5862);
xnor U17606 (N_17606,N_7412,N_6699);
xor U17607 (N_17607,N_8263,N_2358);
xor U17608 (N_17608,N_9686,N_1799);
nor U17609 (N_17609,N_757,N_3785);
xor U17610 (N_17610,N_896,N_1746);
xor U17611 (N_17611,N_6865,N_1176);
or U17612 (N_17612,N_6912,N_2710);
xor U17613 (N_17613,N_9694,N_1951);
and U17614 (N_17614,N_8898,N_6090);
nand U17615 (N_17615,N_3237,N_2785);
xnor U17616 (N_17616,N_1357,N_7799);
nor U17617 (N_17617,N_3559,N_6777);
nor U17618 (N_17618,N_5814,N_5789);
or U17619 (N_17619,N_7233,N_4688);
nand U17620 (N_17620,N_2460,N_2012);
nor U17621 (N_17621,N_9803,N_5069);
nor U17622 (N_17622,N_9401,N_6551);
xor U17623 (N_17623,N_1317,N_8532);
nand U17624 (N_17624,N_389,N_9902);
xnor U17625 (N_17625,N_5478,N_8244);
xnor U17626 (N_17626,N_8994,N_7211);
nor U17627 (N_17627,N_3931,N_5857);
xnor U17628 (N_17628,N_7723,N_2550);
xnor U17629 (N_17629,N_2743,N_7986);
or U17630 (N_17630,N_8668,N_4415);
or U17631 (N_17631,N_9945,N_9692);
nor U17632 (N_17632,N_890,N_5596);
and U17633 (N_17633,N_3429,N_3782);
nor U17634 (N_17634,N_495,N_6035);
or U17635 (N_17635,N_4278,N_8710);
nand U17636 (N_17636,N_6451,N_8566);
and U17637 (N_17637,N_4205,N_9457);
xnor U17638 (N_17638,N_2164,N_7712);
nand U17639 (N_17639,N_6806,N_30);
or U17640 (N_17640,N_6548,N_8447);
or U17641 (N_17641,N_799,N_9522);
nand U17642 (N_17642,N_4848,N_3531);
and U17643 (N_17643,N_9831,N_4952);
and U17644 (N_17644,N_1751,N_5685);
nand U17645 (N_17645,N_425,N_4021);
and U17646 (N_17646,N_3362,N_9972);
nand U17647 (N_17647,N_7168,N_1528);
xnor U17648 (N_17648,N_1081,N_2365);
xnor U17649 (N_17649,N_396,N_9277);
nand U17650 (N_17650,N_4906,N_4114);
nor U17651 (N_17651,N_605,N_9218);
and U17652 (N_17652,N_8063,N_1797);
nand U17653 (N_17653,N_4519,N_6252);
and U17654 (N_17654,N_8141,N_5611);
xnor U17655 (N_17655,N_1309,N_7778);
xnor U17656 (N_17656,N_7821,N_8597);
or U17657 (N_17657,N_938,N_974);
xor U17658 (N_17658,N_1543,N_3716);
and U17659 (N_17659,N_2785,N_4987);
and U17660 (N_17660,N_4484,N_4069);
and U17661 (N_17661,N_5171,N_5674);
xnor U17662 (N_17662,N_2504,N_5769);
nor U17663 (N_17663,N_6955,N_8481);
and U17664 (N_17664,N_6318,N_3207);
nand U17665 (N_17665,N_2979,N_5127);
xnor U17666 (N_17666,N_242,N_3290);
or U17667 (N_17667,N_7358,N_5248);
or U17668 (N_17668,N_7853,N_1726);
nor U17669 (N_17669,N_4442,N_4587);
or U17670 (N_17670,N_6501,N_7804);
or U17671 (N_17671,N_3062,N_8958);
nand U17672 (N_17672,N_7595,N_2162);
or U17673 (N_17673,N_7277,N_3805);
nor U17674 (N_17674,N_6984,N_2167);
xnor U17675 (N_17675,N_3162,N_2980);
xor U17676 (N_17676,N_8287,N_7121);
or U17677 (N_17677,N_4562,N_9297);
nor U17678 (N_17678,N_5032,N_6804);
and U17679 (N_17679,N_2833,N_7841);
and U17680 (N_17680,N_6413,N_3758);
nor U17681 (N_17681,N_363,N_9780);
nor U17682 (N_17682,N_2161,N_4613);
nor U17683 (N_17683,N_2518,N_9157);
and U17684 (N_17684,N_9959,N_7236);
nor U17685 (N_17685,N_8145,N_7678);
xor U17686 (N_17686,N_8026,N_1664);
xnor U17687 (N_17687,N_2147,N_942);
xnor U17688 (N_17688,N_8241,N_7513);
and U17689 (N_17689,N_2000,N_8902);
or U17690 (N_17690,N_7389,N_8180);
nor U17691 (N_17691,N_3543,N_9392);
and U17692 (N_17692,N_6596,N_5774);
nor U17693 (N_17693,N_7808,N_4828);
nor U17694 (N_17694,N_759,N_976);
xor U17695 (N_17695,N_8976,N_1494);
xor U17696 (N_17696,N_4072,N_2917);
xor U17697 (N_17697,N_786,N_4891);
and U17698 (N_17698,N_364,N_3077);
xnor U17699 (N_17699,N_1066,N_8690);
xor U17700 (N_17700,N_7220,N_9842);
and U17701 (N_17701,N_2816,N_4749);
and U17702 (N_17702,N_4074,N_4992);
xor U17703 (N_17703,N_4935,N_9762);
nand U17704 (N_17704,N_3575,N_8036);
nand U17705 (N_17705,N_6589,N_6542);
xor U17706 (N_17706,N_6426,N_9164);
xor U17707 (N_17707,N_2820,N_6508);
nor U17708 (N_17708,N_208,N_1417);
nand U17709 (N_17709,N_260,N_2051);
xnor U17710 (N_17710,N_412,N_9096);
nand U17711 (N_17711,N_7852,N_3618);
and U17712 (N_17712,N_274,N_8987);
nor U17713 (N_17713,N_7759,N_1943);
and U17714 (N_17714,N_6024,N_7210);
nor U17715 (N_17715,N_1336,N_4141);
nand U17716 (N_17716,N_5516,N_6396);
and U17717 (N_17717,N_9110,N_8184);
or U17718 (N_17718,N_2362,N_6572);
nor U17719 (N_17719,N_4375,N_23);
xor U17720 (N_17720,N_1980,N_6672);
nand U17721 (N_17721,N_8264,N_3302);
nor U17722 (N_17722,N_637,N_6981);
nor U17723 (N_17723,N_5991,N_4191);
xnor U17724 (N_17724,N_8192,N_1976);
or U17725 (N_17725,N_8661,N_3251);
xnor U17726 (N_17726,N_4955,N_7815);
and U17727 (N_17727,N_4102,N_5994);
nand U17728 (N_17728,N_2421,N_3221);
nor U17729 (N_17729,N_8753,N_4266);
nand U17730 (N_17730,N_53,N_3174);
and U17731 (N_17731,N_9461,N_4275);
or U17732 (N_17732,N_1843,N_6061);
nand U17733 (N_17733,N_5387,N_5581);
and U17734 (N_17734,N_9812,N_1503);
xnor U17735 (N_17735,N_7357,N_3282);
nand U17736 (N_17736,N_417,N_6478);
xor U17737 (N_17737,N_5526,N_8385);
and U17738 (N_17738,N_725,N_3369);
nor U17739 (N_17739,N_4394,N_508);
nor U17740 (N_17740,N_5298,N_9173);
nand U17741 (N_17741,N_7399,N_4034);
or U17742 (N_17742,N_5773,N_3041);
or U17743 (N_17743,N_2154,N_3099);
and U17744 (N_17744,N_6945,N_4925);
nor U17745 (N_17745,N_9182,N_3552);
nand U17746 (N_17746,N_6791,N_5665);
or U17747 (N_17747,N_8126,N_6667);
or U17748 (N_17748,N_8896,N_1952);
nand U17749 (N_17749,N_788,N_6008);
nand U17750 (N_17750,N_6067,N_4183);
or U17751 (N_17751,N_9847,N_4604);
xnor U17752 (N_17752,N_9863,N_2329);
nor U17753 (N_17753,N_6664,N_4989);
nor U17754 (N_17754,N_8488,N_9670);
and U17755 (N_17755,N_6803,N_3836);
nand U17756 (N_17756,N_5026,N_9808);
and U17757 (N_17757,N_2652,N_6066);
nor U17758 (N_17758,N_7195,N_1428);
or U17759 (N_17759,N_7185,N_4434);
and U17760 (N_17760,N_7370,N_8572);
nor U17761 (N_17761,N_7997,N_5988);
nor U17762 (N_17762,N_5715,N_6039);
or U17763 (N_17763,N_8203,N_2090);
xnor U17764 (N_17764,N_8154,N_1377);
or U17765 (N_17765,N_9842,N_4466);
or U17766 (N_17766,N_9279,N_4221);
or U17767 (N_17767,N_8591,N_7050);
or U17768 (N_17768,N_2042,N_9520);
nor U17769 (N_17769,N_8167,N_9492);
nand U17770 (N_17770,N_9250,N_2583);
nor U17771 (N_17771,N_1953,N_3018);
nand U17772 (N_17772,N_8702,N_8004);
xnor U17773 (N_17773,N_4370,N_3530);
nand U17774 (N_17774,N_5281,N_8793);
or U17775 (N_17775,N_9804,N_9580);
xor U17776 (N_17776,N_3907,N_3055);
and U17777 (N_17777,N_155,N_5652);
nand U17778 (N_17778,N_7067,N_6376);
nor U17779 (N_17779,N_1768,N_736);
nand U17780 (N_17780,N_9766,N_5661);
or U17781 (N_17781,N_9530,N_1507);
nor U17782 (N_17782,N_8596,N_6253);
and U17783 (N_17783,N_4640,N_8438);
xnor U17784 (N_17784,N_4698,N_3154);
nor U17785 (N_17785,N_2377,N_5749);
nand U17786 (N_17786,N_6167,N_7460);
nor U17787 (N_17787,N_8656,N_6619);
and U17788 (N_17788,N_7380,N_2850);
and U17789 (N_17789,N_330,N_4604);
xor U17790 (N_17790,N_7180,N_5657);
or U17791 (N_17791,N_1002,N_415);
xnor U17792 (N_17792,N_7815,N_527);
and U17793 (N_17793,N_3113,N_6683);
nor U17794 (N_17794,N_2333,N_9790);
or U17795 (N_17795,N_6911,N_1017);
and U17796 (N_17796,N_1951,N_5148);
or U17797 (N_17797,N_5847,N_6228);
nand U17798 (N_17798,N_6005,N_2159);
or U17799 (N_17799,N_8717,N_7580);
nor U17800 (N_17800,N_9092,N_1244);
and U17801 (N_17801,N_7932,N_3543);
nand U17802 (N_17802,N_6239,N_1842);
and U17803 (N_17803,N_7254,N_349);
xor U17804 (N_17804,N_1216,N_9927);
xnor U17805 (N_17805,N_9634,N_2819);
xnor U17806 (N_17806,N_1762,N_8967);
and U17807 (N_17807,N_9483,N_1228);
nand U17808 (N_17808,N_645,N_3381);
and U17809 (N_17809,N_9512,N_4390);
and U17810 (N_17810,N_1698,N_5014);
and U17811 (N_17811,N_6578,N_4959);
and U17812 (N_17812,N_8525,N_7118);
and U17813 (N_17813,N_5603,N_9736);
nor U17814 (N_17814,N_5813,N_4226);
or U17815 (N_17815,N_8238,N_731);
or U17816 (N_17816,N_8862,N_1214);
or U17817 (N_17817,N_1479,N_4978);
or U17818 (N_17818,N_7957,N_3730);
nand U17819 (N_17819,N_7501,N_8361);
nand U17820 (N_17820,N_7179,N_2888);
nand U17821 (N_17821,N_5856,N_8894);
nand U17822 (N_17822,N_8388,N_5673);
xor U17823 (N_17823,N_5428,N_1586);
nor U17824 (N_17824,N_3264,N_1378);
nand U17825 (N_17825,N_1477,N_4824);
or U17826 (N_17826,N_1044,N_1328);
nand U17827 (N_17827,N_256,N_2793);
nand U17828 (N_17828,N_744,N_5972);
xnor U17829 (N_17829,N_1634,N_5006);
xnor U17830 (N_17830,N_6050,N_8700);
and U17831 (N_17831,N_2369,N_122);
or U17832 (N_17832,N_6286,N_9017);
or U17833 (N_17833,N_1246,N_3471);
xnor U17834 (N_17834,N_2840,N_2208);
xor U17835 (N_17835,N_2524,N_6263);
nand U17836 (N_17836,N_2572,N_5696);
or U17837 (N_17837,N_5498,N_9009);
xnor U17838 (N_17838,N_7489,N_8115);
and U17839 (N_17839,N_5352,N_6308);
nor U17840 (N_17840,N_7319,N_5395);
and U17841 (N_17841,N_6071,N_1373);
or U17842 (N_17842,N_9730,N_8306);
and U17843 (N_17843,N_1902,N_8189);
nor U17844 (N_17844,N_9651,N_5977);
xnor U17845 (N_17845,N_4742,N_9008);
xor U17846 (N_17846,N_2121,N_2244);
or U17847 (N_17847,N_1886,N_9382);
and U17848 (N_17848,N_9882,N_8948);
xor U17849 (N_17849,N_7363,N_8155);
and U17850 (N_17850,N_1130,N_7295);
or U17851 (N_17851,N_9391,N_2624);
or U17852 (N_17852,N_5880,N_6457);
xnor U17853 (N_17853,N_3949,N_7101);
nor U17854 (N_17854,N_1317,N_4754);
nand U17855 (N_17855,N_801,N_270);
or U17856 (N_17856,N_1174,N_300);
nor U17857 (N_17857,N_6655,N_3281);
or U17858 (N_17858,N_3704,N_9268);
nor U17859 (N_17859,N_1449,N_2644);
and U17860 (N_17860,N_1210,N_8471);
or U17861 (N_17861,N_1385,N_491);
xnor U17862 (N_17862,N_7036,N_4037);
xor U17863 (N_17863,N_1335,N_8703);
xor U17864 (N_17864,N_7240,N_9705);
and U17865 (N_17865,N_3664,N_6178);
or U17866 (N_17866,N_9999,N_7524);
and U17867 (N_17867,N_8751,N_7699);
nand U17868 (N_17868,N_5069,N_5799);
nand U17869 (N_17869,N_5696,N_3194);
and U17870 (N_17870,N_3382,N_3090);
nor U17871 (N_17871,N_3923,N_933);
nand U17872 (N_17872,N_2495,N_5789);
nor U17873 (N_17873,N_1261,N_2146);
nor U17874 (N_17874,N_1024,N_2807);
and U17875 (N_17875,N_3018,N_2085);
nor U17876 (N_17876,N_871,N_4343);
or U17877 (N_17877,N_3510,N_8585);
xor U17878 (N_17878,N_1025,N_9652);
nand U17879 (N_17879,N_4726,N_9271);
and U17880 (N_17880,N_4429,N_8186);
and U17881 (N_17881,N_3897,N_3488);
nand U17882 (N_17882,N_147,N_4141);
nand U17883 (N_17883,N_151,N_5332);
nor U17884 (N_17884,N_8988,N_1578);
xnor U17885 (N_17885,N_4057,N_4690);
nand U17886 (N_17886,N_1279,N_8220);
xor U17887 (N_17887,N_2167,N_1377);
xnor U17888 (N_17888,N_7446,N_9959);
or U17889 (N_17889,N_1077,N_7085);
nor U17890 (N_17890,N_8756,N_6625);
or U17891 (N_17891,N_5079,N_5694);
or U17892 (N_17892,N_2889,N_3252);
nand U17893 (N_17893,N_5405,N_5392);
or U17894 (N_17894,N_3466,N_6263);
xor U17895 (N_17895,N_644,N_7125);
or U17896 (N_17896,N_1758,N_2590);
xnor U17897 (N_17897,N_9894,N_7266);
or U17898 (N_17898,N_1928,N_4438);
nand U17899 (N_17899,N_3570,N_3376);
and U17900 (N_17900,N_5259,N_845);
and U17901 (N_17901,N_2323,N_4400);
nor U17902 (N_17902,N_853,N_491);
or U17903 (N_17903,N_418,N_9923);
or U17904 (N_17904,N_2058,N_477);
xnor U17905 (N_17905,N_7133,N_8672);
and U17906 (N_17906,N_1273,N_847);
nor U17907 (N_17907,N_6668,N_8551);
nand U17908 (N_17908,N_6286,N_3209);
xnor U17909 (N_17909,N_4811,N_1895);
nor U17910 (N_17910,N_5033,N_6017);
nand U17911 (N_17911,N_4576,N_9744);
and U17912 (N_17912,N_6623,N_262);
nand U17913 (N_17913,N_1989,N_9924);
nand U17914 (N_17914,N_9595,N_5234);
nand U17915 (N_17915,N_8795,N_2239);
nand U17916 (N_17916,N_7556,N_8679);
nand U17917 (N_17917,N_6986,N_1890);
nand U17918 (N_17918,N_7012,N_4380);
xnor U17919 (N_17919,N_2167,N_6319);
nand U17920 (N_17920,N_8180,N_5285);
or U17921 (N_17921,N_5169,N_7768);
and U17922 (N_17922,N_8312,N_7275);
nor U17923 (N_17923,N_4950,N_9767);
or U17924 (N_17924,N_4535,N_4802);
nand U17925 (N_17925,N_4790,N_2306);
and U17926 (N_17926,N_6932,N_2647);
xnor U17927 (N_17927,N_6733,N_3030);
nor U17928 (N_17928,N_4802,N_8587);
xnor U17929 (N_17929,N_1891,N_3398);
nor U17930 (N_17930,N_2299,N_171);
nor U17931 (N_17931,N_2639,N_1960);
or U17932 (N_17932,N_1500,N_9470);
and U17933 (N_17933,N_8549,N_470);
or U17934 (N_17934,N_242,N_6258);
or U17935 (N_17935,N_5441,N_5961);
nand U17936 (N_17936,N_4163,N_9369);
or U17937 (N_17937,N_5240,N_8903);
nor U17938 (N_17938,N_7772,N_2754);
nor U17939 (N_17939,N_6515,N_7707);
and U17940 (N_17940,N_3791,N_4875);
nand U17941 (N_17941,N_9334,N_5512);
nor U17942 (N_17942,N_3660,N_2495);
nand U17943 (N_17943,N_5938,N_1597);
nor U17944 (N_17944,N_4134,N_4317);
nor U17945 (N_17945,N_6793,N_7320);
and U17946 (N_17946,N_3736,N_9178);
nand U17947 (N_17947,N_1502,N_5092);
or U17948 (N_17948,N_891,N_9970);
nand U17949 (N_17949,N_8632,N_2121);
nor U17950 (N_17950,N_3767,N_9673);
nor U17951 (N_17951,N_5856,N_1438);
nor U17952 (N_17952,N_2814,N_411);
or U17953 (N_17953,N_5045,N_9772);
or U17954 (N_17954,N_8095,N_5294);
xnor U17955 (N_17955,N_7466,N_978);
or U17956 (N_17956,N_5206,N_9854);
nand U17957 (N_17957,N_2668,N_6381);
xnor U17958 (N_17958,N_7381,N_2143);
or U17959 (N_17959,N_3809,N_2884);
nor U17960 (N_17960,N_8333,N_5797);
or U17961 (N_17961,N_4933,N_7886);
nor U17962 (N_17962,N_724,N_4622);
and U17963 (N_17963,N_9003,N_8130);
nand U17964 (N_17964,N_9537,N_6080);
xnor U17965 (N_17965,N_7054,N_655);
xor U17966 (N_17966,N_1865,N_7807);
nand U17967 (N_17967,N_2321,N_2039);
nor U17968 (N_17968,N_6605,N_879);
and U17969 (N_17969,N_5625,N_5178);
nor U17970 (N_17970,N_2736,N_7142);
and U17971 (N_17971,N_6461,N_2712);
nand U17972 (N_17972,N_7410,N_3463);
or U17973 (N_17973,N_9604,N_4155);
xnor U17974 (N_17974,N_958,N_6940);
or U17975 (N_17975,N_9571,N_5578);
xor U17976 (N_17976,N_8004,N_2004);
xnor U17977 (N_17977,N_893,N_7190);
and U17978 (N_17978,N_1234,N_9372);
nand U17979 (N_17979,N_2694,N_187);
nor U17980 (N_17980,N_7827,N_9);
and U17981 (N_17981,N_3705,N_6341);
xor U17982 (N_17982,N_5261,N_1744);
nand U17983 (N_17983,N_3173,N_67);
and U17984 (N_17984,N_5641,N_3616);
or U17985 (N_17985,N_2020,N_3557);
nand U17986 (N_17986,N_9777,N_3311);
and U17987 (N_17987,N_1728,N_1082);
nand U17988 (N_17988,N_6016,N_6697);
or U17989 (N_17989,N_8319,N_9811);
xnor U17990 (N_17990,N_6462,N_595);
xnor U17991 (N_17991,N_8073,N_2862);
and U17992 (N_17992,N_8786,N_2537);
xnor U17993 (N_17993,N_7546,N_1724);
nand U17994 (N_17994,N_458,N_1811);
xnor U17995 (N_17995,N_2285,N_8167);
nand U17996 (N_17996,N_8017,N_3512);
xor U17997 (N_17997,N_7698,N_9230);
nor U17998 (N_17998,N_1974,N_8055);
or U17999 (N_17999,N_7411,N_2774);
xor U18000 (N_18000,N_6602,N_2328);
nor U18001 (N_18001,N_600,N_9749);
nand U18002 (N_18002,N_3445,N_4138);
nor U18003 (N_18003,N_287,N_489);
xor U18004 (N_18004,N_5409,N_9571);
or U18005 (N_18005,N_5178,N_4433);
or U18006 (N_18006,N_8906,N_7004);
or U18007 (N_18007,N_856,N_9538);
or U18008 (N_18008,N_4792,N_1006);
xor U18009 (N_18009,N_5396,N_2932);
and U18010 (N_18010,N_2815,N_9868);
xnor U18011 (N_18011,N_587,N_5043);
nand U18012 (N_18012,N_4648,N_1898);
nor U18013 (N_18013,N_5837,N_5236);
nand U18014 (N_18014,N_8329,N_3501);
and U18015 (N_18015,N_3669,N_1036);
or U18016 (N_18016,N_8429,N_2054);
nand U18017 (N_18017,N_2793,N_2416);
nand U18018 (N_18018,N_2150,N_8368);
and U18019 (N_18019,N_8419,N_3178);
nand U18020 (N_18020,N_5396,N_7904);
and U18021 (N_18021,N_9444,N_5485);
xor U18022 (N_18022,N_85,N_1454);
nor U18023 (N_18023,N_9960,N_9142);
nand U18024 (N_18024,N_2530,N_1553);
and U18025 (N_18025,N_3087,N_3115);
nor U18026 (N_18026,N_3408,N_1417);
xor U18027 (N_18027,N_1787,N_5654);
nor U18028 (N_18028,N_5839,N_6744);
and U18029 (N_18029,N_7434,N_3297);
or U18030 (N_18030,N_2905,N_89);
nor U18031 (N_18031,N_1906,N_974);
nor U18032 (N_18032,N_2044,N_824);
nor U18033 (N_18033,N_9709,N_9134);
nand U18034 (N_18034,N_4995,N_6962);
xnor U18035 (N_18035,N_7659,N_7111);
nand U18036 (N_18036,N_850,N_5758);
or U18037 (N_18037,N_5620,N_861);
nand U18038 (N_18038,N_9479,N_3916);
or U18039 (N_18039,N_3778,N_1244);
nor U18040 (N_18040,N_6548,N_7415);
and U18041 (N_18041,N_6424,N_3394);
xnor U18042 (N_18042,N_6745,N_2896);
and U18043 (N_18043,N_2394,N_857);
xor U18044 (N_18044,N_6426,N_6086);
nor U18045 (N_18045,N_2733,N_9388);
nand U18046 (N_18046,N_4502,N_1277);
and U18047 (N_18047,N_3983,N_494);
xor U18048 (N_18048,N_9380,N_8899);
nand U18049 (N_18049,N_9517,N_6669);
nor U18050 (N_18050,N_9247,N_6977);
and U18051 (N_18051,N_9009,N_6162);
xnor U18052 (N_18052,N_4423,N_7300);
or U18053 (N_18053,N_1602,N_3178);
nor U18054 (N_18054,N_286,N_2912);
nor U18055 (N_18055,N_6708,N_7596);
xnor U18056 (N_18056,N_7225,N_9124);
or U18057 (N_18057,N_1342,N_7523);
nand U18058 (N_18058,N_66,N_3325);
and U18059 (N_18059,N_3054,N_7924);
nor U18060 (N_18060,N_8128,N_4062);
nor U18061 (N_18061,N_9511,N_9875);
and U18062 (N_18062,N_5149,N_7743);
and U18063 (N_18063,N_6564,N_4814);
nand U18064 (N_18064,N_1852,N_3923);
and U18065 (N_18065,N_3160,N_3023);
nor U18066 (N_18066,N_2783,N_6182);
and U18067 (N_18067,N_6731,N_262);
or U18068 (N_18068,N_5858,N_583);
nor U18069 (N_18069,N_1856,N_2492);
nand U18070 (N_18070,N_9528,N_5914);
xor U18071 (N_18071,N_4538,N_9480);
and U18072 (N_18072,N_8045,N_7110);
xnor U18073 (N_18073,N_8002,N_3774);
xnor U18074 (N_18074,N_5758,N_9234);
or U18075 (N_18075,N_8931,N_6495);
nand U18076 (N_18076,N_627,N_2981);
xor U18077 (N_18077,N_2650,N_7557);
nand U18078 (N_18078,N_4465,N_8969);
or U18079 (N_18079,N_1555,N_9561);
or U18080 (N_18080,N_7088,N_7705);
nor U18081 (N_18081,N_639,N_386);
nor U18082 (N_18082,N_4255,N_3716);
xor U18083 (N_18083,N_8387,N_8678);
nor U18084 (N_18084,N_9413,N_9412);
nor U18085 (N_18085,N_9662,N_6);
nor U18086 (N_18086,N_2745,N_4203);
nand U18087 (N_18087,N_4383,N_8281);
nor U18088 (N_18088,N_650,N_1530);
and U18089 (N_18089,N_6454,N_7671);
nor U18090 (N_18090,N_317,N_4857);
xnor U18091 (N_18091,N_4498,N_5333);
xnor U18092 (N_18092,N_5511,N_4668);
or U18093 (N_18093,N_1636,N_9022);
nor U18094 (N_18094,N_3049,N_328);
or U18095 (N_18095,N_3841,N_3234);
xor U18096 (N_18096,N_8610,N_2013);
xor U18097 (N_18097,N_8201,N_3059);
or U18098 (N_18098,N_5720,N_7620);
nor U18099 (N_18099,N_1237,N_1206);
nand U18100 (N_18100,N_1029,N_2084);
xnor U18101 (N_18101,N_4539,N_6489);
xnor U18102 (N_18102,N_9783,N_9189);
xnor U18103 (N_18103,N_794,N_3719);
nor U18104 (N_18104,N_856,N_1980);
xor U18105 (N_18105,N_9257,N_622);
nand U18106 (N_18106,N_1407,N_8695);
nor U18107 (N_18107,N_760,N_8251);
and U18108 (N_18108,N_6300,N_3683);
xnor U18109 (N_18109,N_4293,N_4827);
and U18110 (N_18110,N_8621,N_1826);
and U18111 (N_18111,N_8448,N_4282);
nand U18112 (N_18112,N_5265,N_3179);
and U18113 (N_18113,N_8534,N_621);
nor U18114 (N_18114,N_5794,N_7439);
nand U18115 (N_18115,N_3650,N_630);
nor U18116 (N_18116,N_3586,N_6944);
nor U18117 (N_18117,N_648,N_5077);
or U18118 (N_18118,N_4519,N_2150);
and U18119 (N_18119,N_6648,N_412);
xnor U18120 (N_18120,N_9642,N_7703);
nand U18121 (N_18121,N_2362,N_9702);
and U18122 (N_18122,N_114,N_4561);
and U18123 (N_18123,N_6067,N_3883);
nand U18124 (N_18124,N_8109,N_543);
and U18125 (N_18125,N_2744,N_8961);
xor U18126 (N_18126,N_4218,N_3700);
nand U18127 (N_18127,N_4040,N_8602);
xnor U18128 (N_18128,N_5601,N_7435);
xnor U18129 (N_18129,N_7599,N_4404);
nor U18130 (N_18130,N_5637,N_9099);
nand U18131 (N_18131,N_2765,N_7155);
nor U18132 (N_18132,N_7285,N_6915);
and U18133 (N_18133,N_2043,N_7446);
and U18134 (N_18134,N_3689,N_3901);
xnor U18135 (N_18135,N_718,N_4883);
xor U18136 (N_18136,N_3694,N_6551);
or U18137 (N_18137,N_7342,N_8409);
nor U18138 (N_18138,N_3008,N_7853);
nor U18139 (N_18139,N_2178,N_1107);
xor U18140 (N_18140,N_3558,N_1665);
nor U18141 (N_18141,N_1796,N_7355);
or U18142 (N_18142,N_538,N_8058);
and U18143 (N_18143,N_9655,N_941);
xnor U18144 (N_18144,N_9579,N_7839);
or U18145 (N_18145,N_485,N_7272);
and U18146 (N_18146,N_3035,N_8775);
or U18147 (N_18147,N_2649,N_4987);
or U18148 (N_18148,N_4927,N_3934);
nand U18149 (N_18149,N_932,N_1753);
nand U18150 (N_18150,N_5448,N_8281);
or U18151 (N_18151,N_1999,N_7954);
or U18152 (N_18152,N_7221,N_6764);
xnor U18153 (N_18153,N_9383,N_4821);
xnor U18154 (N_18154,N_1804,N_1199);
nand U18155 (N_18155,N_5739,N_3818);
nand U18156 (N_18156,N_5937,N_3484);
and U18157 (N_18157,N_4338,N_1685);
or U18158 (N_18158,N_3224,N_2411);
and U18159 (N_18159,N_2297,N_1337);
nand U18160 (N_18160,N_4580,N_7804);
nor U18161 (N_18161,N_1527,N_9231);
xnor U18162 (N_18162,N_1640,N_5338);
nor U18163 (N_18163,N_7274,N_8291);
xor U18164 (N_18164,N_2377,N_4500);
nand U18165 (N_18165,N_5598,N_3361);
and U18166 (N_18166,N_1834,N_7242);
nand U18167 (N_18167,N_6138,N_9926);
and U18168 (N_18168,N_9721,N_8182);
nor U18169 (N_18169,N_6628,N_2260);
nand U18170 (N_18170,N_9067,N_7967);
and U18171 (N_18171,N_4412,N_3575);
or U18172 (N_18172,N_3835,N_7373);
and U18173 (N_18173,N_7269,N_3577);
and U18174 (N_18174,N_579,N_3696);
nor U18175 (N_18175,N_6065,N_9561);
xor U18176 (N_18176,N_5650,N_6095);
and U18177 (N_18177,N_5309,N_9305);
nand U18178 (N_18178,N_2389,N_4169);
xor U18179 (N_18179,N_8909,N_5748);
nor U18180 (N_18180,N_1972,N_9562);
xnor U18181 (N_18181,N_8522,N_3037);
and U18182 (N_18182,N_9145,N_2914);
nand U18183 (N_18183,N_6651,N_4820);
nor U18184 (N_18184,N_9852,N_5455);
and U18185 (N_18185,N_7963,N_708);
and U18186 (N_18186,N_7163,N_8015);
xnor U18187 (N_18187,N_6895,N_8071);
nor U18188 (N_18188,N_4846,N_4458);
xnor U18189 (N_18189,N_3012,N_8796);
or U18190 (N_18190,N_9717,N_4705);
or U18191 (N_18191,N_4824,N_6268);
or U18192 (N_18192,N_8551,N_6702);
or U18193 (N_18193,N_5443,N_4298);
nor U18194 (N_18194,N_5877,N_6042);
nor U18195 (N_18195,N_313,N_939);
nor U18196 (N_18196,N_7225,N_1470);
nor U18197 (N_18197,N_8969,N_1029);
or U18198 (N_18198,N_190,N_4211);
or U18199 (N_18199,N_3938,N_3425);
xor U18200 (N_18200,N_2088,N_3807);
or U18201 (N_18201,N_5495,N_8481);
nor U18202 (N_18202,N_793,N_8391);
or U18203 (N_18203,N_1586,N_4909);
xnor U18204 (N_18204,N_5555,N_3814);
nand U18205 (N_18205,N_2970,N_4904);
or U18206 (N_18206,N_4868,N_5617);
nor U18207 (N_18207,N_7052,N_3037);
xnor U18208 (N_18208,N_2828,N_3703);
nor U18209 (N_18209,N_1400,N_2144);
and U18210 (N_18210,N_5712,N_1572);
or U18211 (N_18211,N_4616,N_2596);
xnor U18212 (N_18212,N_3303,N_8198);
and U18213 (N_18213,N_1800,N_9726);
nor U18214 (N_18214,N_1169,N_2280);
nor U18215 (N_18215,N_9801,N_8802);
or U18216 (N_18216,N_3801,N_6033);
xnor U18217 (N_18217,N_7419,N_7421);
xor U18218 (N_18218,N_7790,N_6157);
and U18219 (N_18219,N_5475,N_3343);
and U18220 (N_18220,N_625,N_1544);
xnor U18221 (N_18221,N_3748,N_5593);
nor U18222 (N_18222,N_3909,N_5360);
or U18223 (N_18223,N_8998,N_3048);
nand U18224 (N_18224,N_7334,N_6388);
and U18225 (N_18225,N_9619,N_1134);
nor U18226 (N_18226,N_5559,N_3535);
and U18227 (N_18227,N_5791,N_8792);
nand U18228 (N_18228,N_8040,N_947);
and U18229 (N_18229,N_634,N_409);
nand U18230 (N_18230,N_7277,N_7821);
or U18231 (N_18231,N_1509,N_3546);
nand U18232 (N_18232,N_9414,N_649);
or U18233 (N_18233,N_9182,N_6656);
and U18234 (N_18234,N_7967,N_9306);
or U18235 (N_18235,N_9267,N_5849);
nand U18236 (N_18236,N_9721,N_1701);
or U18237 (N_18237,N_5451,N_6399);
and U18238 (N_18238,N_558,N_4712);
xnor U18239 (N_18239,N_1829,N_8769);
nor U18240 (N_18240,N_2864,N_260);
nor U18241 (N_18241,N_2282,N_1223);
xnor U18242 (N_18242,N_8908,N_9846);
nor U18243 (N_18243,N_2562,N_2710);
and U18244 (N_18244,N_1049,N_6009);
xnor U18245 (N_18245,N_5727,N_8522);
nand U18246 (N_18246,N_1866,N_6181);
and U18247 (N_18247,N_5313,N_3693);
nor U18248 (N_18248,N_2078,N_5734);
nor U18249 (N_18249,N_2105,N_2730);
or U18250 (N_18250,N_145,N_5116);
xor U18251 (N_18251,N_1800,N_4399);
and U18252 (N_18252,N_7763,N_2802);
nor U18253 (N_18253,N_6529,N_8399);
xor U18254 (N_18254,N_7233,N_5137);
xor U18255 (N_18255,N_5990,N_6174);
nor U18256 (N_18256,N_369,N_8458);
or U18257 (N_18257,N_576,N_7441);
and U18258 (N_18258,N_6714,N_6691);
xor U18259 (N_18259,N_2412,N_9240);
nand U18260 (N_18260,N_9180,N_3506);
nor U18261 (N_18261,N_6524,N_5462);
nor U18262 (N_18262,N_9423,N_4592);
and U18263 (N_18263,N_1491,N_3887);
or U18264 (N_18264,N_741,N_1321);
nand U18265 (N_18265,N_1934,N_8776);
nor U18266 (N_18266,N_8595,N_9484);
nand U18267 (N_18267,N_931,N_4803);
or U18268 (N_18268,N_2024,N_9401);
or U18269 (N_18269,N_2226,N_4177);
or U18270 (N_18270,N_2227,N_3227);
nand U18271 (N_18271,N_8462,N_9770);
and U18272 (N_18272,N_7101,N_8753);
and U18273 (N_18273,N_1070,N_7071);
xor U18274 (N_18274,N_9093,N_8104);
xnor U18275 (N_18275,N_7060,N_8182);
xor U18276 (N_18276,N_5106,N_7189);
nand U18277 (N_18277,N_3135,N_9141);
and U18278 (N_18278,N_6263,N_9525);
xnor U18279 (N_18279,N_9849,N_1704);
or U18280 (N_18280,N_1434,N_8507);
nand U18281 (N_18281,N_8997,N_4327);
and U18282 (N_18282,N_9414,N_5481);
or U18283 (N_18283,N_5954,N_1904);
nor U18284 (N_18284,N_1348,N_3956);
and U18285 (N_18285,N_1329,N_1222);
nor U18286 (N_18286,N_8635,N_9306);
or U18287 (N_18287,N_627,N_8239);
nand U18288 (N_18288,N_1512,N_1469);
and U18289 (N_18289,N_7472,N_8950);
or U18290 (N_18290,N_5989,N_4734);
xnor U18291 (N_18291,N_1921,N_3876);
nor U18292 (N_18292,N_5300,N_8473);
xor U18293 (N_18293,N_3879,N_7209);
xnor U18294 (N_18294,N_165,N_8177);
or U18295 (N_18295,N_2746,N_2310);
and U18296 (N_18296,N_4897,N_274);
or U18297 (N_18297,N_1012,N_2791);
nand U18298 (N_18298,N_6445,N_634);
xor U18299 (N_18299,N_8094,N_2441);
xor U18300 (N_18300,N_2944,N_6373);
nor U18301 (N_18301,N_4050,N_180);
nand U18302 (N_18302,N_5230,N_8178);
xor U18303 (N_18303,N_167,N_9104);
xor U18304 (N_18304,N_7454,N_3964);
and U18305 (N_18305,N_2206,N_3432);
nand U18306 (N_18306,N_4382,N_2152);
nor U18307 (N_18307,N_6011,N_4990);
xor U18308 (N_18308,N_9930,N_553);
xnor U18309 (N_18309,N_9660,N_3821);
and U18310 (N_18310,N_6229,N_9051);
and U18311 (N_18311,N_9270,N_5951);
nand U18312 (N_18312,N_6788,N_1704);
and U18313 (N_18313,N_758,N_4883);
nor U18314 (N_18314,N_979,N_8984);
or U18315 (N_18315,N_6898,N_9651);
xnor U18316 (N_18316,N_7850,N_5777);
and U18317 (N_18317,N_9916,N_2635);
nand U18318 (N_18318,N_9757,N_9858);
nand U18319 (N_18319,N_3807,N_4964);
and U18320 (N_18320,N_1418,N_685);
and U18321 (N_18321,N_2344,N_2970);
or U18322 (N_18322,N_9452,N_5218);
and U18323 (N_18323,N_3558,N_9019);
nor U18324 (N_18324,N_7879,N_2627);
xor U18325 (N_18325,N_8046,N_4279);
xor U18326 (N_18326,N_2820,N_9159);
nand U18327 (N_18327,N_8602,N_2626);
xor U18328 (N_18328,N_2794,N_8732);
nor U18329 (N_18329,N_4193,N_9039);
or U18330 (N_18330,N_2648,N_6752);
xnor U18331 (N_18331,N_6788,N_4055);
or U18332 (N_18332,N_3133,N_3124);
and U18333 (N_18333,N_5013,N_3061);
xor U18334 (N_18334,N_1847,N_5203);
nand U18335 (N_18335,N_4253,N_465);
nand U18336 (N_18336,N_5400,N_2176);
nor U18337 (N_18337,N_2151,N_495);
xnor U18338 (N_18338,N_5607,N_2247);
nand U18339 (N_18339,N_2452,N_7749);
nor U18340 (N_18340,N_8631,N_4137);
and U18341 (N_18341,N_4742,N_3635);
nor U18342 (N_18342,N_9255,N_7612);
or U18343 (N_18343,N_497,N_5303);
and U18344 (N_18344,N_4339,N_2281);
nor U18345 (N_18345,N_1935,N_568);
or U18346 (N_18346,N_7192,N_7168);
or U18347 (N_18347,N_9449,N_2599);
xnor U18348 (N_18348,N_5357,N_2649);
xor U18349 (N_18349,N_355,N_1528);
and U18350 (N_18350,N_7789,N_6166);
nand U18351 (N_18351,N_1449,N_9734);
xor U18352 (N_18352,N_8751,N_1962);
nor U18353 (N_18353,N_6104,N_100);
or U18354 (N_18354,N_8641,N_2792);
and U18355 (N_18355,N_8945,N_6598);
or U18356 (N_18356,N_432,N_9529);
xor U18357 (N_18357,N_62,N_7938);
xnor U18358 (N_18358,N_6878,N_9031);
nor U18359 (N_18359,N_4167,N_326);
or U18360 (N_18360,N_908,N_5505);
or U18361 (N_18361,N_6426,N_3337);
xor U18362 (N_18362,N_4103,N_9548);
nor U18363 (N_18363,N_7549,N_9320);
and U18364 (N_18364,N_1214,N_1031);
nor U18365 (N_18365,N_3007,N_9567);
nor U18366 (N_18366,N_8747,N_9957);
or U18367 (N_18367,N_9738,N_9541);
xnor U18368 (N_18368,N_5041,N_2378);
nor U18369 (N_18369,N_2416,N_8354);
xnor U18370 (N_18370,N_3711,N_6960);
xnor U18371 (N_18371,N_3536,N_1866);
nor U18372 (N_18372,N_9254,N_8288);
nor U18373 (N_18373,N_7847,N_3221);
nor U18374 (N_18374,N_548,N_6532);
or U18375 (N_18375,N_9037,N_2964);
nand U18376 (N_18376,N_7268,N_2922);
nor U18377 (N_18377,N_8538,N_6521);
and U18378 (N_18378,N_882,N_2471);
nor U18379 (N_18379,N_1919,N_9331);
or U18380 (N_18380,N_4600,N_8833);
nor U18381 (N_18381,N_4845,N_2817);
nand U18382 (N_18382,N_4538,N_3053);
nand U18383 (N_18383,N_610,N_4403);
or U18384 (N_18384,N_1751,N_4234);
and U18385 (N_18385,N_6774,N_7289);
and U18386 (N_18386,N_560,N_8278);
nand U18387 (N_18387,N_9830,N_7290);
nand U18388 (N_18388,N_9552,N_5850);
or U18389 (N_18389,N_8487,N_6979);
nand U18390 (N_18390,N_1106,N_2753);
nor U18391 (N_18391,N_4719,N_4487);
or U18392 (N_18392,N_4723,N_8310);
and U18393 (N_18393,N_6641,N_1098);
xnor U18394 (N_18394,N_7350,N_5897);
and U18395 (N_18395,N_8353,N_6473);
or U18396 (N_18396,N_2683,N_7305);
and U18397 (N_18397,N_5837,N_3602);
nand U18398 (N_18398,N_4273,N_2055);
or U18399 (N_18399,N_6792,N_1223);
xnor U18400 (N_18400,N_7386,N_1850);
xor U18401 (N_18401,N_1249,N_3439);
nand U18402 (N_18402,N_1625,N_6460);
and U18403 (N_18403,N_2131,N_4857);
and U18404 (N_18404,N_4403,N_7866);
nand U18405 (N_18405,N_2967,N_3468);
nand U18406 (N_18406,N_1254,N_64);
nor U18407 (N_18407,N_4792,N_9835);
nand U18408 (N_18408,N_6358,N_7732);
nor U18409 (N_18409,N_483,N_4601);
nand U18410 (N_18410,N_6020,N_8772);
nand U18411 (N_18411,N_964,N_519);
or U18412 (N_18412,N_565,N_6960);
or U18413 (N_18413,N_2104,N_8355);
nor U18414 (N_18414,N_1769,N_7567);
nor U18415 (N_18415,N_6361,N_6809);
nand U18416 (N_18416,N_4316,N_5111);
and U18417 (N_18417,N_2446,N_6271);
nand U18418 (N_18418,N_3756,N_4158);
nand U18419 (N_18419,N_5150,N_6450);
nor U18420 (N_18420,N_5280,N_1688);
xor U18421 (N_18421,N_8321,N_7651);
nand U18422 (N_18422,N_6756,N_5803);
xnor U18423 (N_18423,N_9695,N_3381);
and U18424 (N_18424,N_4987,N_1830);
nand U18425 (N_18425,N_486,N_5605);
nand U18426 (N_18426,N_7221,N_2555);
nand U18427 (N_18427,N_4451,N_4994);
and U18428 (N_18428,N_8868,N_3274);
xnor U18429 (N_18429,N_4550,N_8649);
and U18430 (N_18430,N_8633,N_2287);
nand U18431 (N_18431,N_8628,N_9110);
or U18432 (N_18432,N_8896,N_7018);
or U18433 (N_18433,N_1523,N_7791);
nand U18434 (N_18434,N_2664,N_9814);
xnor U18435 (N_18435,N_6939,N_9268);
or U18436 (N_18436,N_5795,N_8459);
nor U18437 (N_18437,N_7329,N_2847);
and U18438 (N_18438,N_8725,N_5349);
and U18439 (N_18439,N_2621,N_6609);
xor U18440 (N_18440,N_2238,N_4566);
or U18441 (N_18441,N_3761,N_6533);
or U18442 (N_18442,N_4119,N_2549);
or U18443 (N_18443,N_7491,N_4133);
xnor U18444 (N_18444,N_9288,N_7387);
nand U18445 (N_18445,N_1219,N_5522);
or U18446 (N_18446,N_7940,N_3280);
and U18447 (N_18447,N_3778,N_4757);
xnor U18448 (N_18448,N_7017,N_3253);
xor U18449 (N_18449,N_7668,N_194);
or U18450 (N_18450,N_3275,N_1015);
or U18451 (N_18451,N_8851,N_3073);
nand U18452 (N_18452,N_8843,N_5128);
nor U18453 (N_18453,N_3143,N_3151);
xnor U18454 (N_18454,N_247,N_142);
or U18455 (N_18455,N_5290,N_7510);
nor U18456 (N_18456,N_6010,N_2145);
xor U18457 (N_18457,N_1152,N_3334);
nor U18458 (N_18458,N_6712,N_5197);
nand U18459 (N_18459,N_9828,N_3637);
xnor U18460 (N_18460,N_3895,N_1959);
nand U18461 (N_18461,N_2733,N_2266);
nor U18462 (N_18462,N_9442,N_130);
or U18463 (N_18463,N_9048,N_2218);
xnor U18464 (N_18464,N_8753,N_4521);
xnor U18465 (N_18465,N_7906,N_7048);
and U18466 (N_18466,N_4304,N_8832);
or U18467 (N_18467,N_7750,N_418);
nor U18468 (N_18468,N_3540,N_4108);
nor U18469 (N_18469,N_2076,N_8336);
or U18470 (N_18470,N_4694,N_7415);
xnor U18471 (N_18471,N_5032,N_8356);
nand U18472 (N_18472,N_1725,N_3475);
nand U18473 (N_18473,N_7748,N_2381);
xor U18474 (N_18474,N_5875,N_1980);
nand U18475 (N_18475,N_7460,N_4679);
or U18476 (N_18476,N_5083,N_2884);
nand U18477 (N_18477,N_5960,N_3846);
nor U18478 (N_18478,N_9604,N_1112);
nor U18479 (N_18479,N_205,N_768);
or U18480 (N_18480,N_2926,N_5706);
and U18481 (N_18481,N_7503,N_9856);
xnor U18482 (N_18482,N_4206,N_6258);
and U18483 (N_18483,N_2933,N_4566);
xor U18484 (N_18484,N_8060,N_7179);
and U18485 (N_18485,N_1579,N_6298);
or U18486 (N_18486,N_2314,N_908);
or U18487 (N_18487,N_9654,N_4206);
xnor U18488 (N_18488,N_8033,N_9631);
xor U18489 (N_18489,N_2549,N_1467);
and U18490 (N_18490,N_121,N_7576);
nor U18491 (N_18491,N_2177,N_5675);
nor U18492 (N_18492,N_3050,N_1760);
nor U18493 (N_18493,N_5470,N_8357);
xnor U18494 (N_18494,N_3108,N_216);
and U18495 (N_18495,N_9931,N_6347);
xor U18496 (N_18496,N_4623,N_263);
nor U18497 (N_18497,N_7533,N_9577);
nor U18498 (N_18498,N_8919,N_6708);
and U18499 (N_18499,N_6801,N_7703);
xor U18500 (N_18500,N_4899,N_9156);
nand U18501 (N_18501,N_8451,N_2577);
nand U18502 (N_18502,N_8692,N_9831);
or U18503 (N_18503,N_5329,N_8761);
and U18504 (N_18504,N_4173,N_8795);
xor U18505 (N_18505,N_7781,N_8614);
or U18506 (N_18506,N_3914,N_5558);
or U18507 (N_18507,N_5058,N_4299);
nand U18508 (N_18508,N_3564,N_753);
or U18509 (N_18509,N_7837,N_2232);
nand U18510 (N_18510,N_6058,N_2477);
or U18511 (N_18511,N_776,N_2839);
or U18512 (N_18512,N_6963,N_4603);
and U18513 (N_18513,N_7687,N_6369);
or U18514 (N_18514,N_4688,N_7527);
xnor U18515 (N_18515,N_9695,N_8744);
or U18516 (N_18516,N_8895,N_1053);
xnor U18517 (N_18517,N_7851,N_2426);
or U18518 (N_18518,N_61,N_3959);
nor U18519 (N_18519,N_9791,N_3023);
xnor U18520 (N_18520,N_9872,N_463);
nor U18521 (N_18521,N_2829,N_5137);
and U18522 (N_18522,N_8365,N_7075);
nor U18523 (N_18523,N_4635,N_1102);
nor U18524 (N_18524,N_296,N_2140);
nand U18525 (N_18525,N_2343,N_4944);
nand U18526 (N_18526,N_1214,N_3852);
or U18527 (N_18527,N_4089,N_6708);
nand U18528 (N_18528,N_9986,N_8558);
nand U18529 (N_18529,N_1016,N_3143);
and U18530 (N_18530,N_3310,N_2459);
xor U18531 (N_18531,N_7015,N_9813);
nand U18532 (N_18532,N_1831,N_8605);
nor U18533 (N_18533,N_8050,N_7534);
xnor U18534 (N_18534,N_4668,N_3087);
and U18535 (N_18535,N_8795,N_5233);
nand U18536 (N_18536,N_5838,N_5921);
nor U18537 (N_18537,N_4053,N_3027);
nor U18538 (N_18538,N_5817,N_9395);
or U18539 (N_18539,N_1014,N_4611);
nand U18540 (N_18540,N_2497,N_5233);
nor U18541 (N_18541,N_4905,N_7176);
nor U18542 (N_18542,N_9026,N_4133);
or U18543 (N_18543,N_3052,N_9719);
xor U18544 (N_18544,N_9686,N_3035);
xor U18545 (N_18545,N_8763,N_9558);
nand U18546 (N_18546,N_1715,N_4556);
or U18547 (N_18547,N_2838,N_544);
and U18548 (N_18548,N_5994,N_2018);
or U18549 (N_18549,N_4319,N_9234);
nand U18550 (N_18550,N_4477,N_8615);
or U18551 (N_18551,N_8322,N_5210);
or U18552 (N_18552,N_5919,N_9118);
nor U18553 (N_18553,N_3130,N_4700);
or U18554 (N_18554,N_5387,N_3552);
nor U18555 (N_18555,N_8922,N_5851);
and U18556 (N_18556,N_5084,N_7522);
nor U18557 (N_18557,N_4830,N_3671);
xnor U18558 (N_18558,N_2274,N_1875);
nand U18559 (N_18559,N_4909,N_7273);
xor U18560 (N_18560,N_2451,N_9566);
nor U18561 (N_18561,N_2422,N_4799);
or U18562 (N_18562,N_8302,N_3159);
and U18563 (N_18563,N_1890,N_5957);
and U18564 (N_18564,N_2352,N_8440);
and U18565 (N_18565,N_7281,N_6952);
and U18566 (N_18566,N_3623,N_5267);
nor U18567 (N_18567,N_5373,N_3762);
or U18568 (N_18568,N_4304,N_8336);
xnor U18569 (N_18569,N_4627,N_381);
nand U18570 (N_18570,N_362,N_1876);
nor U18571 (N_18571,N_7552,N_2247);
and U18572 (N_18572,N_9354,N_1686);
xnor U18573 (N_18573,N_6993,N_9440);
nor U18574 (N_18574,N_653,N_5636);
or U18575 (N_18575,N_9537,N_4535);
or U18576 (N_18576,N_2913,N_8208);
and U18577 (N_18577,N_3361,N_4878);
or U18578 (N_18578,N_7969,N_1425);
nand U18579 (N_18579,N_990,N_3035);
or U18580 (N_18580,N_6445,N_9471);
and U18581 (N_18581,N_4966,N_2637);
xnor U18582 (N_18582,N_3717,N_5777);
or U18583 (N_18583,N_6381,N_6187);
and U18584 (N_18584,N_1602,N_795);
nand U18585 (N_18585,N_7208,N_4396);
and U18586 (N_18586,N_1471,N_8598);
xor U18587 (N_18587,N_1663,N_1501);
xnor U18588 (N_18588,N_7746,N_1363);
and U18589 (N_18589,N_4002,N_2);
or U18590 (N_18590,N_6802,N_1765);
or U18591 (N_18591,N_4340,N_5732);
xor U18592 (N_18592,N_9944,N_5433);
and U18593 (N_18593,N_9515,N_8470);
or U18594 (N_18594,N_2260,N_1327);
or U18595 (N_18595,N_6762,N_9301);
nand U18596 (N_18596,N_1238,N_1065);
nand U18597 (N_18597,N_9716,N_6702);
nand U18598 (N_18598,N_9171,N_7811);
or U18599 (N_18599,N_1311,N_3787);
xnor U18600 (N_18600,N_4720,N_2719);
nand U18601 (N_18601,N_6276,N_5324);
or U18602 (N_18602,N_5427,N_2635);
and U18603 (N_18603,N_2258,N_12);
and U18604 (N_18604,N_222,N_7545);
and U18605 (N_18605,N_2102,N_1132);
nor U18606 (N_18606,N_8005,N_8987);
or U18607 (N_18607,N_6150,N_5978);
nand U18608 (N_18608,N_4198,N_6682);
nor U18609 (N_18609,N_9185,N_4247);
nand U18610 (N_18610,N_5318,N_8745);
nor U18611 (N_18611,N_8069,N_7891);
or U18612 (N_18612,N_7262,N_8840);
and U18613 (N_18613,N_2639,N_2901);
nor U18614 (N_18614,N_7980,N_9120);
or U18615 (N_18615,N_9110,N_7860);
nor U18616 (N_18616,N_8038,N_3655);
nand U18617 (N_18617,N_1766,N_8182);
or U18618 (N_18618,N_3832,N_8081);
nor U18619 (N_18619,N_6205,N_6343);
xor U18620 (N_18620,N_4283,N_1231);
and U18621 (N_18621,N_3672,N_259);
or U18622 (N_18622,N_9495,N_7553);
nand U18623 (N_18623,N_3536,N_7674);
xnor U18624 (N_18624,N_5214,N_8679);
or U18625 (N_18625,N_4970,N_7539);
xnor U18626 (N_18626,N_2484,N_7504);
nand U18627 (N_18627,N_4790,N_6375);
nand U18628 (N_18628,N_8132,N_8938);
nor U18629 (N_18629,N_6169,N_2701);
and U18630 (N_18630,N_5037,N_5836);
xnor U18631 (N_18631,N_1281,N_4769);
xor U18632 (N_18632,N_3639,N_530);
nor U18633 (N_18633,N_2141,N_8925);
xnor U18634 (N_18634,N_1043,N_1280);
or U18635 (N_18635,N_6467,N_8689);
xor U18636 (N_18636,N_7575,N_2597);
nand U18637 (N_18637,N_2843,N_553);
nor U18638 (N_18638,N_7624,N_8066);
or U18639 (N_18639,N_413,N_4421);
and U18640 (N_18640,N_550,N_8389);
xnor U18641 (N_18641,N_223,N_3320);
nand U18642 (N_18642,N_5710,N_6479);
nand U18643 (N_18643,N_7687,N_5445);
xor U18644 (N_18644,N_8867,N_2321);
nand U18645 (N_18645,N_2144,N_7111);
nand U18646 (N_18646,N_9313,N_7655);
and U18647 (N_18647,N_6574,N_6519);
nor U18648 (N_18648,N_5700,N_3889);
nand U18649 (N_18649,N_4047,N_6982);
nand U18650 (N_18650,N_5605,N_6168);
and U18651 (N_18651,N_6933,N_9527);
xnor U18652 (N_18652,N_3570,N_1178);
nand U18653 (N_18653,N_5138,N_1283);
and U18654 (N_18654,N_5449,N_8272);
nand U18655 (N_18655,N_9287,N_6877);
and U18656 (N_18656,N_3992,N_3475);
nand U18657 (N_18657,N_8786,N_9128);
nand U18658 (N_18658,N_5720,N_762);
and U18659 (N_18659,N_5810,N_9083);
or U18660 (N_18660,N_2239,N_7472);
nand U18661 (N_18661,N_8231,N_7205);
and U18662 (N_18662,N_9813,N_1429);
nor U18663 (N_18663,N_4659,N_8326);
nor U18664 (N_18664,N_926,N_3981);
nor U18665 (N_18665,N_9382,N_7594);
xnor U18666 (N_18666,N_5375,N_7762);
nor U18667 (N_18667,N_2548,N_5227);
and U18668 (N_18668,N_8962,N_1726);
xor U18669 (N_18669,N_831,N_5149);
xor U18670 (N_18670,N_4023,N_1989);
or U18671 (N_18671,N_2061,N_6427);
or U18672 (N_18672,N_481,N_1968);
nand U18673 (N_18673,N_7661,N_8390);
nor U18674 (N_18674,N_9689,N_6803);
nand U18675 (N_18675,N_907,N_259);
and U18676 (N_18676,N_8001,N_4653);
xnor U18677 (N_18677,N_8544,N_7817);
nand U18678 (N_18678,N_3876,N_221);
xnor U18679 (N_18679,N_3834,N_3543);
nand U18680 (N_18680,N_6256,N_475);
and U18681 (N_18681,N_8349,N_1120);
xnor U18682 (N_18682,N_6541,N_3731);
xor U18683 (N_18683,N_1723,N_6003);
xnor U18684 (N_18684,N_9945,N_3900);
nand U18685 (N_18685,N_3778,N_6639);
or U18686 (N_18686,N_5002,N_4170);
xnor U18687 (N_18687,N_5202,N_4439);
xnor U18688 (N_18688,N_5831,N_7362);
or U18689 (N_18689,N_7663,N_8451);
nand U18690 (N_18690,N_4197,N_416);
nand U18691 (N_18691,N_6171,N_5231);
nand U18692 (N_18692,N_1111,N_6419);
xnor U18693 (N_18693,N_1590,N_4771);
and U18694 (N_18694,N_5475,N_2011);
or U18695 (N_18695,N_5233,N_4916);
or U18696 (N_18696,N_794,N_3061);
and U18697 (N_18697,N_2821,N_8595);
and U18698 (N_18698,N_4446,N_4474);
nor U18699 (N_18699,N_329,N_518);
or U18700 (N_18700,N_7053,N_4863);
nand U18701 (N_18701,N_4077,N_7682);
or U18702 (N_18702,N_7788,N_3586);
or U18703 (N_18703,N_6318,N_3680);
and U18704 (N_18704,N_1006,N_8);
xor U18705 (N_18705,N_5760,N_19);
xnor U18706 (N_18706,N_1840,N_1748);
nor U18707 (N_18707,N_9387,N_3191);
nor U18708 (N_18708,N_9968,N_5707);
nor U18709 (N_18709,N_8060,N_1069);
nand U18710 (N_18710,N_8263,N_3339);
xnor U18711 (N_18711,N_6534,N_8229);
and U18712 (N_18712,N_1077,N_9667);
nor U18713 (N_18713,N_4553,N_785);
nand U18714 (N_18714,N_3108,N_2182);
nand U18715 (N_18715,N_3656,N_4981);
xor U18716 (N_18716,N_4132,N_3621);
xnor U18717 (N_18717,N_4697,N_1983);
nand U18718 (N_18718,N_7534,N_1387);
nor U18719 (N_18719,N_2966,N_8634);
and U18720 (N_18720,N_8791,N_7285);
xnor U18721 (N_18721,N_6401,N_7076);
or U18722 (N_18722,N_516,N_2399);
nor U18723 (N_18723,N_2178,N_5347);
xnor U18724 (N_18724,N_1384,N_5911);
or U18725 (N_18725,N_8746,N_3879);
xor U18726 (N_18726,N_4996,N_481);
xnor U18727 (N_18727,N_2114,N_7553);
nor U18728 (N_18728,N_7143,N_2586);
xnor U18729 (N_18729,N_1123,N_8966);
and U18730 (N_18730,N_4836,N_4314);
or U18731 (N_18731,N_6943,N_7983);
and U18732 (N_18732,N_7185,N_772);
nor U18733 (N_18733,N_5093,N_419);
or U18734 (N_18734,N_7674,N_9329);
and U18735 (N_18735,N_6256,N_8345);
xor U18736 (N_18736,N_8826,N_9263);
or U18737 (N_18737,N_2910,N_344);
and U18738 (N_18738,N_2568,N_5680);
nand U18739 (N_18739,N_8066,N_4902);
or U18740 (N_18740,N_6562,N_4659);
xnor U18741 (N_18741,N_6801,N_3457);
xor U18742 (N_18742,N_8405,N_9658);
xor U18743 (N_18743,N_9093,N_9048);
or U18744 (N_18744,N_5993,N_8893);
nand U18745 (N_18745,N_3296,N_2486);
or U18746 (N_18746,N_8177,N_5904);
nand U18747 (N_18747,N_7483,N_7405);
xnor U18748 (N_18748,N_3578,N_9910);
nor U18749 (N_18749,N_3277,N_684);
nand U18750 (N_18750,N_1372,N_5775);
and U18751 (N_18751,N_2342,N_8927);
xnor U18752 (N_18752,N_2771,N_6003);
nor U18753 (N_18753,N_7503,N_8406);
and U18754 (N_18754,N_3198,N_7622);
nand U18755 (N_18755,N_4368,N_9034);
xnor U18756 (N_18756,N_7543,N_6185);
nand U18757 (N_18757,N_6211,N_7493);
or U18758 (N_18758,N_1936,N_2630);
nor U18759 (N_18759,N_5652,N_6349);
and U18760 (N_18760,N_4170,N_516);
or U18761 (N_18761,N_2448,N_5408);
nor U18762 (N_18762,N_957,N_9218);
or U18763 (N_18763,N_6637,N_6982);
and U18764 (N_18764,N_5634,N_5663);
and U18765 (N_18765,N_2450,N_386);
nor U18766 (N_18766,N_2655,N_3952);
nor U18767 (N_18767,N_5464,N_4341);
nand U18768 (N_18768,N_422,N_7616);
and U18769 (N_18769,N_6117,N_1863);
or U18770 (N_18770,N_2623,N_2442);
or U18771 (N_18771,N_5820,N_6161);
nand U18772 (N_18772,N_3707,N_2878);
xor U18773 (N_18773,N_7873,N_3935);
nand U18774 (N_18774,N_7297,N_9655);
xor U18775 (N_18775,N_4455,N_3280);
or U18776 (N_18776,N_8238,N_8857);
nand U18777 (N_18777,N_558,N_5525);
or U18778 (N_18778,N_8969,N_4828);
nand U18779 (N_18779,N_9543,N_9140);
xor U18780 (N_18780,N_9498,N_9250);
nand U18781 (N_18781,N_9496,N_2775);
nand U18782 (N_18782,N_7960,N_7273);
and U18783 (N_18783,N_4341,N_4904);
nand U18784 (N_18784,N_6740,N_6146);
nor U18785 (N_18785,N_8447,N_3040);
nand U18786 (N_18786,N_5337,N_4777);
nor U18787 (N_18787,N_6374,N_2546);
or U18788 (N_18788,N_8589,N_1110);
nand U18789 (N_18789,N_6207,N_2930);
nand U18790 (N_18790,N_9595,N_8752);
and U18791 (N_18791,N_8883,N_296);
and U18792 (N_18792,N_1072,N_8076);
nand U18793 (N_18793,N_4864,N_7177);
nand U18794 (N_18794,N_835,N_7851);
nor U18795 (N_18795,N_4457,N_1044);
nor U18796 (N_18796,N_8312,N_4681);
nand U18797 (N_18797,N_4608,N_3512);
or U18798 (N_18798,N_804,N_5176);
or U18799 (N_18799,N_2876,N_2036);
nand U18800 (N_18800,N_4779,N_8193);
and U18801 (N_18801,N_9273,N_5522);
xor U18802 (N_18802,N_1767,N_6832);
xor U18803 (N_18803,N_7849,N_4714);
xnor U18804 (N_18804,N_4730,N_6111);
or U18805 (N_18805,N_7400,N_999);
or U18806 (N_18806,N_5047,N_8392);
nor U18807 (N_18807,N_8789,N_6840);
nor U18808 (N_18808,N_4584,N_9263);
xor U18809 (N_18809,N_4384,N_6223);
or U18810 (N_18810,N_7532,N_2907);
and U18811 (N_18811,N_9451,N_8098);
or U18812 (N_18812,N_2921,N_5765);
or U18813 (N_18813,N_8575,N_2565);
or U18814 (N_18814,N_495,N_4131);
nand U18815 (N_18815,N_450,N_6469);
xnor U18816 (N_18816,N_6196,N_6716);
nor U18817 (N_18817,N_4719,N_7219);
and U18818 (N_18818,N_5052,N_7216);
xor U18819 (N_18819,N_4610,N_1220);
xnor U18820 (N_18820,N_3182,N_1488);
or U18821 (N_18821,N_5970,N_3149);
nor U18822 (N_18822,N_860,N_2177);
nor U18823 (N_18823,N_642,N_2049);
xor U18824 (N_18824,N_9212,N_3814);
or U18825 (N_18825,N_9403,N_5576);
xnor U18826 (N_18826,N_7064,N_4004);
or U18827 (N_18827,N_8255,N_213);
nor U18828 (N_18828,N_4117,N_5334);
nand U18829 (N_18829,N_4503,N_6725);
nor U18830 (N_18830,N_8407,N_294);
nor U18831 (N_18831,N_933,N_1728);
and U18832 (N_18832,N_2573,N_9987);
or U18833 (N_18833,N_8000,N_8210);
nand U18834 (N_18834,N_6002,N_6246);
or U18835 (N_18835,N_2632,N_284);
xor U18836 (N_18836,N_4492,N_1555);
and U18837 (N_18837,N_5646,N_1180);
and U18838 (N_18838,N_4169,N_7929);
nand U18839 (N_18839,N_6883,N_3022);
xnor U18840 (N_18840,N_9892,N_2764);
or U18841 (N_18841,N_3277,N_8379);
nand U18842 (N_18842,N_9562,N_7352);
nand U18843 (N_18843,N_3105,N_6967);
nand U18844 (N_18844,N_6834,N_2149);
and U18845 (N_18845,N_478,N_697);
nand U18846 (N_18846,N_5206,N_6483);
and U18847 (N_18847,N_1815,N_4146);
nor U18848 (N_18848,N_6164,N_3452);
nand U18849 (N_18849,N_8297,N_1006);
or U18850 (N_18850,N_6408,N_6110);
nand U18851 (N_18851,N_9580,N_819);
and U18852 (N_18852,N_6519,N_9434);
and U18853 (N_18853,N_2275,N_7869);
nand U18854 (N_18854,N_688,N_7678);
or U18855 (N_18855,N_2380,N_2552);
nand U18856 (N_18856,N_5600,N_9600);
xor U18857 (N_18857,N_1928,N_6284);
and U18858 (N_18858,N_4913,N_7754);
nand U18859 (N_18859,N_5164,N_6404);
and U18860 (N_18860,N_6030,N_7733);
or U18861 (N_18861,N_329,N_7827);
or U18862 (N_18862,N_7661,N_93);
xnor U18863 (N_18863,N_7357,N_1020);
nor U18864 (N_18864,N_3104,N_2159);
xor U18865 (N_18865,N_5337,N_3309);
xor U18866 (N_18866,N_1105,N_7163);
or U18867 (N_18867,N_9239,N_1081);
xor U18868 (N_18868,N_4081,N_5935);
or U18869 (N_18869,N_4184,N_15);
and U18870 (N_18870,N_5878,N_3418);
nand U18871 (N_18871,N_7214,N_1112);
xnor U18872 (N_18872,N_5893,N_651);
nand U18873 (N_18873,N_7246,N_5761);
nor U18874 (N_18874,N_8843,N_3806);
xnor U18875 (N_18875,N_4095,N_3361);
or U18876 (N_18876,N_9838,N_6565);
or U18877 (N_18877,N_9536,N_1420);
nor U18878 (N_18878,N_9383,N_7962);
or U18879 (N_18879,N_7346,N_4128);
xor U18880 (N_18880,N_4758,N_433);
nor U18881 (N_18881,N_9003,N_3216);
xnor U18882 (N_18882,N_6746,N_4339);
xnor U18883 (N_18883,N_4224,N_8703);
nor U18884 (N_18884,N_6992,N_307);
nor U18885 (N_18885,N_6976,N_9712);
or U18886 (N_18886,N_4632,N_8206);
or U18887 (N_18887,N_6019,N_9963);
xnor U18888 (N_18888,N_5920,N_5436);
nor U18889 (N_18889,N_9773,N_2829);
xnor U18890 (N_18890,N_8550,N_3648);
xor U18891 (N_18891,N_90,N_7971);
xor U18892 (N_18892,N_5048,N_3847);
or U18893 (N_18893,N_8089,N_3508);
xor U18894 (N_18894,N_9079,N_1057);
and U18895 (N_18895,N_9953,N_2077);
and U18896 (N_18896,N_7056,N_142);
or U18897 (N_18897,N_5161,N_7231);
or U18898 (N_18898,N_3878,N_3190);
nor U18899 (N_18899,N_5212,N_6468);
or U18900 (N_18900,N_4265,N_3781);
xor U18901 (N_18901,N_6263,N_9984);
nor U18902 (N_18902,N_7042,N_8714);
nor U18903 (N_18903,N_9913,N_9249);
nand U18904 (N_18904,N_2735,N_1056);
and U18905 (N_18905,N_4608,N_1526);
xor U18906 (N_18906,N_9097,N_9276);
nand U18907 (N_18907,N_6868,N_2224);
and U18908 (N_18908,N_681,N_1450);
xor U18909 (N_18909,N_6750,N_3516);
nand U18910 (N_18910,N_987,N_309);
nor U18911 (N_18911,N_3786,N_8169);
nand U18912 (N_18912,N_885,N_4843);
or U18913 (N_18913,N_3676,N_9816);
nor U18914 (N_18914,N_5383,N_6281);
or U18915 (N_18915,N_2919,N_8489);
xnor U18916 (N_18916,N_7074,N_8648);
nor U18917 (N_18917,N_8705,N_2987);
xor U18918 (N_18918,N_1021,N_8714);
nor U18919 (N_18919,N_2013,N_797);
and U18920 (N_18920,N_6954,N_73);
and U18921 (N_18921,N_2703,N_6222);
nor U18922 (N_18922,N_9976,N_1288);
nand U18923 (N_18923,N_2196,N_4602);
or U18924 (N_18924,N_1328,N_6293);
or U18925 (N_18925,N_2534,N_6818);
nor U18926 (N_18926,N_9827,N_8310);
nand U18927 (N_18927,N_7470,N_7527);
nand U18928 (N_18928,N_5410,N_6814);
nor U18929 (N_18929,N_819,N_9206);
nor U18930 (N_18930,N_9660,N_1570);
nand U18931 (N_18931,N_8935,N_3480);
xor U18932 (N_18932,N_7973,N_3002);
nand U18933 (N_18933,N_4749,N_8776);
nor U18934 (N_18934,N_7009,N_2460);
or U18935 (N_18935,N_2607,N_4374);
or U18936 (N_18936,N_5532,N_2808);
or U18937 (N_18937,N_5101,N_6502);
nor U18938 (N_18938,N_1496,N_3940);
nor U18939 (N_18939,N_5822,N_2833);
xor U18940 (N_18940,N_135,N_4273);
or U18941 (N_18941,N_8476,N_9824);
nand U18942 (N_18942,N_3699,N_3215);
xnor U18943 (N_18943,N_4011,N_3817);
nand U18944 (N_18944,N_5497,N_7214);
and U18945 (N_18945,N_6000,N_9386);
nand U18946 (N_18946,N_6600,N_1727);
or U18947 (N_18947,N_7271,N_3328);
and U18948 (N_18948,N_3541,N_6649);
nor U18949 (N_18949,N_1648,N_1432);
nor U18950 (N_18950,N_9101,N_5064);
or U18951 (N_18951,N_3309,N_9271);
or U18952 (N_18952,N_5594,N_898);
nand U18953 (N_18953,N_7483,N_2861);
xnor U18954 (N_18954,N_1404,N_8489);
nor U18955 (N_18955,N_4793,N_9636);
nand U18956 (N_18956,N_5962,N_8445);
nand U18957 (N_18957,N_6927,N_489);
nand U18958 (N_18958,N_9813,N_7134);
or U18959 (N_18959,N_7498,N_9048);
or U18960 (N_18960,N_8085,N_1148);
nand U18961 (N_18961,N_3665,N_8808);
nand U18962 (N_18962,N_7901,N_1257);
or U18963 (N_18963,N_1874,N_1752);
and U18964 (N_18964,N_1617,N_9033);
nor U18965 (N_18965,N_6319,N_2425);
or U18966 (N_18966,N_4435,N_6459);
nor U18967 (N_18967,N_4366,N_6555);
or U18968 (N_18968,N_4461,N_4438);
nand U18969 (N_18969,N_8032,N_5560);
xor U18970 (N_18970,N_8703,N_9849);
xnor U18971 (N_18971,N_6269,N_9797);
nand U18972 (N_18972,N_3881,N_6857);
nor U18973 (N_18973,N_4192,N_975);
and U18974 (N_18974,N_5805,N_6416);
nor U18975 (N_18975,N_5621,N_3730);
or U18976 (N_18976,N_2177,N_8984);
xor U18977 (N_18977,N_5608,N_3140);
or U18978 (N_18978,N_3923,N_1235);
or U18979 (N_18979,N_4972,N_221);
nand U18980 (N_18980,N_5534,N_5145);
xor U18981 (N_18981,N_7687,N_6694);
nand U18982 (N_18982,N_859,N_7236);
nor U18983 (N_18983,N_3678,N_8266);
and U18984 (N_18984,N_3958,N_178);
and U18985 (N_18985,N_8169,N_1411);
nor U18986 (N_18986,N_4345,N_4564);
nor U18987 (N_18987,N_8574,N_1969);
nor U18988 (N_18988,N_3258,N_4363);
and U18989 (N_18989,N_2033,N_5952);
nand U18990 (N_18990,N_8247,N_9442);
nor U18991 (N_18991,N_8899,N_2431);
xor U18992 (N_18992,N_9901,N_6190);
nor U18993 (N_18993,N_7264,N_5810);
nor U18994 (N_18994,N_5979,N_4557);
or U18995 (N_18995,N_9661,N_2781);
nand U18996 (N_18996,N_9633,N_865);
or U18997 (N_18997,N_7579,N_8381);
or U18998 (N_18998,N_3606,N_8796);
nor U18999 (N_18999,N_1805,N_7266);
or U19000 (N_19000,N_2003,N_4080);
xnor U19001 (N_19001,N_3427,N_5815);
or U19002 (N_19002,N_6332,N_5283);
nand U19003 (N_19003,N_7086,N_8663);
or U19004 (N_19004,N_46,N_4418);
nor U19005 (N_19005,N_6154,N_8769);
xnor U19006 (N_19006,N_8578,N_5298);
nand U19007 (N_19007,N_7167,N_4172);
or U19008 (N_19008,N_9049,N_379);
xor U19009 (N_19009,N_9906,N_7586);
nand U19010 (N_19010,N_920,N_825);
xnor U19011 (N_19011,N_7571,N_3037);
or U19012 (N_19012,N_8453,N_7588);
nor U19013 (N_19013,N_4775,N_1885);
and U19014 (N_19014,N_1338,N_3351);
nor U19015 (N_19015,N_1033,N_3838);
xnor U19016 (N_19016,N_1116,N_1911);
xnor U19017 (N_19017,N_7606,N_1724);
nand U19018 (N_19018,N_860,N_7617);
nor U19019 (N_19019,N_9073,N_2521);
nand U19020 (N_19020,N_9944,N_1411);
nand U19021 (N_19021,N_7202,N_7644);
nor U19022 (N_19022,N_9233,N_5337);
or U19023 (N_19023,N_207,N_7040);
and U19024 (N_19024,N_5996,N_3314);
and U19025 (N_19025,N_7470,N_7105);
and U19026 (N_19026,N_203,N_7520);
nand U19027 (N_19027,N_4155,N_7461);
nor U19028 (N_19028,N_3666,N_2852);
and U19029 (N_19029,N_1951,N_5876);
nor U19030 (N_19030,N_2008,N_6590);
xor U19031 (N_19031,N_5298,N_6289);
xor U19032 (N_19032,N_3662,N_8397);
xnor U19033 (N_19033,N_3431,N_1189);
nand U19034 (N_19034,N_3515,N_2617);
nor U19035 (N_19035,N_7019,N_8371);
nand U19036 (N_19036,N_8261,N_5427);
xor U19037 (N_19037,N_7108,N_5405);
or U19038 (N_19038,N_5396,N_5730);
xnor U19039 (N_19039,N_7495,N_7852);
xnor U19040 (N_19040,N_187,N_2919);
nand U19041 (N_19041,N_4610,N_1489);
xor U19042 (N_19042,N_5852,N_8078);
nand U19043 (N_19043,N_6979,N_3176);
and U19044 (N_19044,N_2196,N_9436);
xor U19045 (N_19045,N_7053,N_1753);
or U19046 (N_19046,N_8959,N_3028);
and U19047 (N_19047,N_9779,N_3175);
nand U19048 (N_19048,N_5149,N_8093);
or U19049 (N_19049,N_6333,N_152);
and U19050 (N_19050,N_8287,N_7452);
and U19051 (N_19051,N_3233,N_4151);
or U19052 (N_19052,N_9943,N_4338);
nor U19053 (N_19053,N_878,N_8783);
nor U19054 (N_19054,N_388,N_1132);
nand U19055 (N_19055,N_8025,N_6161);
and U19056 (N_19056,N_3774,N_3537);
nor U19057 (N_19057,N_1731,N_137);
nor U19058 (N_19058,N_8817,N_2723);
xnor U19059 (N_19059,N_6390,N_2362);
nor U19060 (N_19060,N_281,N_9146);
and U19061 (N_19061,N_4953,N_9285);
nand U19062 (N_19062,N_7617,N_5837);
nand U19063 (N_19063,N_5857,N_8823);
or U19064 (N_19064,N_334,N_8948);
nor U19065 (N_19065,N_2779,N_5971);
nand U19066 (N_19066,N_2892,N_4864);
xnor U19067 (N_19067,N_3925,N_9451);
nor U19068 (N_19068,N_20,N_5405);
xor U19069 (N_19069,N_3660,N_2195);
xnor U19070 (N_19070,N_4391,N_9264);
xnor U19071 (N_19071,N_6756,N_8791);
nand U19072 (N_19072,N_1142,N_115);
xnor U19073 (N_19073,N_1214,N_6340);
and U19074 (N_19074,N_9232,N_4326);
or U19075 (N_19075,N_2876,N_4545);
and U19076 (N_19076,N_2280,N_5214);
nand U19077 (N_19077,N_4715,N_9357);
nor U19078 (N_19078,N_6047,N_378);
nor U19079 (N_19079,N_8417,N_7077);
nand U19080 (N_19080,N_1798,N_209);
or U19081 (N_19081,N_2321,N_9146);
and U19082 (N_19082,N_4192,N_2169);
and U19083 (N_19083,N_7687,N_2599);
xnor U19084 (N_19084,N_7901,N_8983);
nand U19085 (N_19085,N_3133,N_9140);
xor U19086 (N_19086,N_9944,N_5400);
and U19087 (N_19087,N_6855,N_4271);
or U19088 (N_19088,N_189,N_8353);
nor U19089 (N_19089,N_9373,N_9275);
xnor U19090 (N_19090,N_9750,N_9529);
or U19091 (N_19091,N_7375,N_7796);
xnor U19092 (N_19092,N_7878,N_3815);
and U19093 (N_19093,N_630,N_4137);
or U19094 (N_19094,N_3527,N_4651);
and U19095 (N_19095,N_4553,N_1568);
nor U19096 (N_19096,N_1081,N_683);
nor U19097 (N_19097,N_803,N_4786);
or U19098 (N_19098,N_5934,N_8078);
or U19099 (N_19099,N_2674,N_474);
nor U19100 (N_19100,N_7102,N_1026);
nor U19101 (N_19101,N_4519,N_1075);
or U19102 (N_19102,N_7495,N_6361);
or U19103 (N_19103,N_5301,N_1620);
nand U19104 (N_19104,N_4121,N_5335);
and U19105 (N_19105,N_9093,N_3021);
nor U19106 (N_19106,N_6472,N_1994);
nor U19107 (N_19107,N_5765,N_4576);
and U19108 (N_19108,N_6125,N_5039);
nor U19109 (N_19109,N_3372,N_488);
nor U19110 (N_19110,N_4089,N_1413);
or U19111 (N_19111,N_9689,N_5740);
and U19112 (N_19112,N_3521,N_3382);
and U19113 (N_19113,N_2891,N_6768);
and U19114 (N_19114,N_1094,N_2961);
nor U19115 (N_19115,N_8345,N_10);
nand U19116 (N_19116,N_3413,N_6050);
xnor U19117 (N_19117,N_2350,N_2002);
and U19118 (N_19118,N_8048,N_7090);
xor U19119 (N_19119,N_2086,N_638);
and U19120 (N_19120,N_9980,N_4487);
nand U19121 (N_19121,N_4488,N_2294);
xnor U19122 (N_19122,N_1373,N_648);
xor U19123 (N_19123,N_6986,N_9407);
or U19124 (N_19124,N_2234,N_6444);
and U19125 (N_19125,N_6468,N_1588);
xor U19126 (N_19126,N_1090,N_8133);
nand U19127 (N_19127,N_3605,N_20);
nor U19128 (N_19128,N_6227,N_3382);
nand U19129 (N_19129,N_9214,N_2821);
xnor U19130 (N_19130,N_8864,N_988);
xor U19131 (N_19131,N_7581,N_1195);
xnor U19132 (N_19132,N_6419,N_937);
nor U19133 (N_19133,N_437,N_6891);
or U19134 (N_19134,N_9,N_3759);
nor U19135 (N_19135,N_9159,N_7941);
xor U19136 (N_19136,N_8738,N_7263);
or U19137 (N_19137,N_2482,N_7692);
and U19138 (N_19138,N_9999,N_8785);
or U19139 (N_19139,N_7425,N_8499);
or U19140 (N_19140,N_7249,N_4799);
or U19141 (N_19141,N_8306,N_5453);
nand U19142 (N_19142,N_5257,N_387);
nor U19143 (N_19143,N_8471,N_9989);
nor U19144 (N_19144,N_1080,N_6859);
or U19145 (N_19145,N_1645,N_3323);
or U19146 (N_19146,N_8712,N_3648);
nand U19147 (N_19147,N_369,N_5843);
xnor U19148 (N_19148,N_5499,N_7242);
or U19149 (N_19149,N_7927,N_7544);
nor U19150 (N_19150,N_4139,N_9080);
or U19151 (N_19151,N_8436,N_6858);
xor U19152 (N_19152,N_6739,N_4878);
or U19153 (N_19153,N_2993,N_332);
and U19154 (N_19154,N_1922,N_6577);
or U19155 (N_19155,N_7053,N_2546);
nand U19156 (N_19156,N_6750,N_1543);
xnor U19157 (N_19157,N_7218,N_4213);
nor U19158 (N_19158,N_7178,N_9637);
or U19159 (N_19159,N_7938,N_7718);
xnor U19160 (N_19160,N_1750,N_443);
or U19161 (N_19161,N_6639,N_1538);
nor U19162 (N_19162,N_488,N_6556);
nand U19163 (N_19163,N_1290,N_2218);
xor U19164 (N_19164,N_6785,N_7611);
and U19165 (N_19165,N_4568,N_6546);
nand U19166 (N_19166,N_4443,N_3065);
nand U19167 (N_19167,N_7074,N_3146);
xor U19168 (N_19168,N_5120,N_1789);
nor U19169 (N_19169,N_9753,N_8682);
and U19170 (N_19170,N_1476,N_8671);
xor U19171 (N_19171,N_5987,N_687);
xnor U19172 (N_19172,N_9647,N_6902);
nand U19173 (N_19173,N_1845,N_1618);
or U19174 (N_19174,N_6675,N_8105);
nand U19175 (N_19175,N_1835,N_8989);
or U19176 (N_19176,N_4960,N_6405);
nor U19177 (N_19177,N_9156,N_5505);
nand U19178 (N_19178,N_3564,N_9062);
or U19179 (N_19179,N_1078,N_1604);
and U19180 (N_19180,N_517,N_8598);
nor U19181 (N_19181,N_2472,N_1785);
xnor U19182 (N_19182,N_3151,N_6477);
and U19183 (N_19183,N_7293,N_7135);
or U19184 (N_19184,N_2116,N_1201);
xnor U19185 (N_19185,N_5553,N_7108);
and U19186 (N_19186,N_2022,N_8920);
or U19187 (N_19187,N_6214,N_6201);
nor U19188 (N_19188,N_2435,N_7932);
nand U19189 (N_19189,N_1900,N_5924);
nand U19190 (N_19190,N_3618,N_1216);
nand U19191 (N_19191,N_2775,N_2269);
nor U19192 (N_19192,N_4320,N_1716);
or U19193 (N_19193,N_4261,N_4701);
nand U19194 (N_19194,N_4644,N_7667);
and U19195 (N_19195,N_395,N_7089);
nand U19196 (N_19196,N_8583,N_842);
or U19197 (N_19197,N_1720,N_214);
and U19198 (N_19198,N_5596,N_2552);
xnor U19199 (N_19199,N_9501,N_5341);
nand U19200 (N_19200,N_4795,N_9686);
or U19201 (N_19201,N_9376,N_2136);
and U19202 (N_19202,N_3754,N_7470);
nor U19203 (N_19203,N_4683,N_2145);
and U19204 (N_19204,N_1904,N_9914);
nand U19205 (N_19205,N_7009,N_6846);
and U19206 (N_19206,N_1170,N_8448);
and U19207 (N_19207,N_6093,N_3608);
nor U19208 (N_19208,N_8854,N_5879);
xnor U19209 (N_19209,N_9389,N_7799);
nand U19210 (N_19210,N_9761,N_7959);
and U19211 (N_19211,N_1571,N_2083);
xnor U19212 (N_19212,N_8234,N_1408);
nand U19213 (N_19213,N_7012,N_1323);
nor U19214 (N_19214,N_8278,N_682);
and U19215 (N_19215,N_6775,N_6632);
nand U19216 (N_19216,N_5905,N_4565);
and U19217 (N_19217,N_1225,N_4828);
xor U19218 (N_19218,N_2334,N_9498);
nand U19219 (N_19219,N_8813,N_4130);
xnor U19220 (N_19220,N_6194,N_244);
nand U19221 (N_19221,N_3655,N_519);
xor U19222 (N_19222,N_4968,N_598);
xnor U19223 (N_19223,N_3261,N_1875);
and U19224 (N_19224,N_2615,N_9702);
and U19225 (N_19225,N_3075,N_4637);
xor U19226 (N_19226,N_2765,N_6671);
and U19227 (N_19227,N_4403,N_8399);
nor U19228 (N_19228,N_9278,N_3596);
and U19229 (N_19229,N_5768,N_1427);
nand U19230 (N_19230,N_4534,N_3833);
nor U19231 (N_19231,N_5890,N_5670);
nand U19232 (N_19232,N_2297,N_3218);
nand U19233 (N_19233,N_2049,N_8030);
and U19234 (N_19234,N_7806,N_3215);
and U19235 (N_19235,N_8250,N_8807);
nor U19236 (N_19236,N_9548,N_7334);
nor U19237 (N_19237,N_6436,N_3585);
or U19238 (N_19238,N_8106,N_1270);
nor U19239 (N_19239,N_9626,N_5981);
nand U19240 (N_19240,N_733,N_6183);
or U19241 (N_19241,N_9647,N_1189);
and U19242 (N_19242,N_7061,N_4594);
or U19243 (N_19243,N_7618,N_1751);
nand U19244 (N_19244,N_4207,N_6520);
nor U19245 (N_19245,N_3664,N_3020);
nor U19246 (N_19246,N_5807,N_9353);
xnor U19247 (N_19247,N_2976,N_2862);
xor U19248 (N_19248,N_6406,N_6034);
and U19249 (N_19249,N_1868,N_3431);
or U19250 (N_19250,N_5014,N_6317);
nand U19251 (N_19251,N_2647,N_6855);
or U19252 (N_19252,N_9687,N_728);
and U19253 (N_19253,N_3202,N_7338);
nor U19254 (N_19254,N_2396,N_222);
or U19255 (N_19255,N_3614,N_2737);
nand U19256 (N_19256,N_7454,N_1132);
nand U19257 (N_19257,N_8061,N_1823);
nand U19258 (N_19258,N_1060,N_7650);
and U19259 (N_19259,N_5771,N_7393);
nand U19260 (N_19260,N_1471,N_7742);
xnor U19261 (N_19261,N_6029,N_4837);
xnor U19262 (N_19262,N_3403,N_1736);
xor U19263 (N_19263,N_5658,N_9348);
xnor U19264 (N_19264,N_3166,N_9071);
xnor U19265 (N_19265,N_5432,N_7521);
or U19266 (N_19266,N_8251,N_9458);
nand U19267 (N_19267,N_5025,N_1221);
nand U19268 (N_19268,N_8684,N_4369);
xor U19269 (N_19269,N_1422,N_4994);
nand U19270 (N_19270,N_8082,N_3618);
nor U19271 (N_19271,N_973,N_8272);
nor U19272 (N_19272,N_9417,N_9478);
xor U19273 (N_19273,N_5651,N_6262);
nand U19274 (N_19274,N_3745,N_5736);
nand U19275 (N_19275,N_4717,N_2151);
or U19276 (N_19276,N_3728,N_4283);
nor U19277 (N_19277,N_5990,N_9854);
nor U19278 (N_19278,N_2361,N_9634);
and U19279 (N_19279,N_3602,N_8514);
nor U19280 (N_19280,N_9844,N_1878);
nor U19281 (N_19281,N_8679,N_6196);
and U19282 (N_19282,N_7909,N_6853);
nor U19283 (N_19283,N_6638,N_8914);
xor U19284 (N_19284,N_6923,N_4866);
nor U19285 (N_19285,N_9165,N_2428);
or U19286 (N_19286,N_1166,N_1662);
nor U19287 (N_19287,N_4461,N_7741);
and U19288 (N_19288,N_610,N_8262);
or U19289 (N_19289,N_6030,N_5092);
and U19290 (N_19290,N_5042,N_9211);
nand U19291 (N_19291,N_40,N_2297);
xnor U19292 (N_19292,N_9869,N_8859);
nand U19293 (N_19293,N_3769,N_5223);
nand U19294 (N_19294,N_2509,N_9277);
and U19295 (N_19295,N_3729,N_5027);
xnor U19296 (N_19296,N_7666,N_8528);
xnor U19297 (N_19297,N_1307,N_6722);
xor U19298 (N_19298,N_9128,N_2153);
and U19299 (N_19299,N_7524,N_8755);
nor U19300 (N_19300,N_5666,N_9855);
or U19301 (N_19301,N_8889,N_4217);
or U19302 (N_19302,N_6767,N_3696);
nor U19303 (N_19303,N_3978,N_3877);
nor U19304 (N_19304,N_397,N_1531);
and U19305 (N_19305,N_8878,N_507);
and U19306 (N_19306,N_2285,N_247);
xnor U19307 (N_19307,N_9861,N_2286);
nand U19308 (N_19308,N_8606,N_3501);
xor U19309 (N_19309,N_7160,N_9764);
and U19310 (N_19310,N_1824,N_8399);
nor U19311 (N_19311,N_8430,N_2977);
nor U19312 (N_19312,N_9079,N_6308);
xor U19313 (N_19313,N_4768,N_2027);
nor U19314 (N_19314,N_8469,N_2044);
xor U19315 (N_19315,N_3212,N_1245);
xor U19316 (N_19316,N_9579,N_4251);
nor U19317 (N_19317,N_4040,N_7421);
or U19318 (N_19318,N_818,N_1687);
or U19319 (N_19319,N_3907,N_7877);
nor U19320 (N_19320,N_8416,N_2388);
nor U19321 (N_19321,N_7223,N_27);
and U19322 (N_19322,N_742,N_113);
xor U19323 (N_19323,N_1799,N_2138);
and U19324 (N_19324,N_2000,N_1970);
and U19325 (N_19325,N_1290,N_4514);
or U19326 (N_19326,N_7206,N_7773);
nor U19327 (N_19327,N_7546,N_4844);
nand U19328 (N_19328,N_619,N_2686);
nand U19329 (N_19329,N_3049,N_9107);
or U19330 (N_19330,N_2033,N_9725);
xor U19331 (N_19331,N_3189,N_6616);
or U19332 (N_19332,N_6282,N_6945);
nand U19333 (N_19333,N_8547,N_2433);
nand U19334 (N_19334,N_5414,N_4950);
nor U19335 (N_19335,N_9838,N_142);
nor U19336 (N_19336,N_3715,N_9699);
or U19337 (N_19337,N_1583,N_5504);
and U19338 (N_19338,N_6012,N_3516);
or U19339 (N_19339,N_6364,N_9169);
and U19340 (N_19340,N_2316,N_8640);
nor U19341 (N_19341,N_9538,N_4109);
nand U19342 (N_19342,N_412,N_2226);
or U19343 (N_19343,N_9681,N_5156);
xnor U19344 (N_19344,N_5956,N_3470);
nand U19345 (N_19345,N_7225,N_4396);
xor U19346 (N_19346,N_9798,N_6544);
and U19347 (N_19347,N_890,N_7223);
and U19348 (N_19348,N_7266,N_6127);
and U19349 (N_19349,N_6788,N_3325);
nor U19350 (N_19350,N_5106,N_1536);
nor U19351 (N_19351,N_5705,N_8813);
nor U19352 (N_19352,N_463,N_2411);
or U19353 (N_19353,N_1876,N_1160);
nor U19354 (N_19354,N_2920,N_1702);
xor U19355 (N_19355,N_1825,N_6042);
nor U19356 (N_19356,N_9907,N_5318);
or U19357 (N_19357,N_6957,N_7630);
nand U19358 (N_19358,N_8109,N_4375);
xor U19359 (N_19359,N_4076,N_2657);
xnor U19360 (N_19360,N_1000,N_4144);
nand U19361 (N_19361,N_8168,N_923);
and U19362 (N_19362,N_4816,N_5390);
nand U19363 (N_19363,N_8552,N_7536);
xnor U19364 (N_19364,N_9414,N_1640);
or U19365 (N_19365,N_1340,N_8797);
xor U19366 (N_19366,N_2919,N_3163);
and U19367 (N_19367,N_349,N_19);
or U19368 (N_19368,N_1675,N_2096);
nand U19369 (N_19369,N_4166,N_3940);
xor U19370 (N_19370,N_2092,N_9905);
or U19371 (N_19371,N_2552,N_7910);
nand U19372 (N_19372,N_9465,N_4172);
and U19373 (N_19373,N_2511,N_7721);
xor U19374 (N_19374,N_4539,N_6634);
and U19375 (N_19375,N_6985,N_8294);
nor U19376 (N_19376,N_1898,N_8767);
nand U19377 (N_19377,N_8445,N_4993);
xnor U19378 (N_19378,N_8343,N_8698);
nor U19379 (N_19379,N_5852,N_5248);
or U19380 (N_19380,N_6604,N_1442);
nor U19381 (N_19381,N_3355,N_2152);
nor U19382 (N_19382,N_6438,N_1094);
xor U19383 (N_19383,N_6002,N_6936);
and U19384 (N_19384,N_1431,N_4496);
xnor U19385 (N_19385,N_5028,N_875);
and U19386 (N_19386,N_4121,N_5015);
nand U19387 (N_19387,N_5530,N_5369);
and U19388 (N_19388,N_189,N_9115);
xnor U19389 (N_19389,N_3612,N_8154);
nor U19390 (N_19390,N_68,N_5738);
xor U19391 (N_19391,N_6290,N_1181);
nand U19392 (N_19392,N_7289,N_2843);
nor U19393 (N_19393,N_6502,N_7331);
nand U19394 (N_19394,N_3544,N_3296);
or U19395 (N_19395,N_1016,N_7525);
and U19396 (N_19396,N_9820,N_5254);
xor U19397 (N_19397,N_8093,N_3808);
nor U19398 (N_19398,N_6048,N_9838);
or U19399 (N_19399,N_8524,N_9695);
nor U19400 (N_19400,N_850,N_1891);
and U19401 (N_19401,N_972,N_9599);
nor U19402 (N_19402,N_6099,N_5417);
nand U19403 (N_19403,N_4293,N_5581);
nand U19404 (N_19404,N_4062,N_9324);
nand U19405 (N_19405,N_8525,N_5754);
or U19406 (N_19406,N_4083,N_7160);
or U19407 (N_19407,N_2032,N_4051);
nor U19408 (N_19408,N_9199,N_5102);
nand U19409 (N_19409,N_8695,N_3373);
and U19410 (N_19410,N_6491,N_3096);
nor U19411 (N_19411,N_2914,N_9365);
or U19412 (N_19412,N_9987,N_7296);
nand U19413 (N_19413,N_7259,N_9160);
xnor U19414 (N_19414,N_6140,N_3952);
or U19415 (N_19415,N_6306,N_6264);
nand U19416 (N_19416,N_7660,N_2918);
nor U19417 (N_19417,N_4212,N_511);
or U19418 (N_19418,N_3389,N_6615);
nor U19419 (N_19419,N_9031,N_2188);
nand U19420 (N_19420,N_3732,N_4655);
and U19421 (N_19421,N_5878,N_2945);
and U19422 (N_19422,N_8179,N_5954);
and U19423 (N_19423,N_4296,N_3007);
nor U19424 (N_19424,N_162,N_5202);
nor U19425 (N_19425,N_6079,N_3869);
nand U19426 (N_19426,N_557,N_4832);
nor U19427 (N_19427,N_2730,N_7131);
nand U19428 (N_19428,N_6971,N_7332);
nand U19429 (N_19429,N_9945,N_3391);
or U19430 (N_19430,N_6119,N_424);
and U19431 (N_19431,N_5895,N_6475);
and U19432 (N_19432,N_4367,N_9967);
or U19433 (N_19433,N_9605,N_2623);
xnor U19434 (N_19434,N_5629,N_9038);
or U19435 (N_19435,N_3244,N_8295);
and U19436 (N_19436,N_6965,N_9413);
xor U19437 (N_19437,N_2013,N_953);
nor U19438 (N_19438,N_8998,N_8239);
nand U19439 (N_19439,N_2330,N_6605);
xnor U19440 (N_19440,N_6142,N_695);
xnor U19441 (N_19441,N_7728,N_5146);
and U19442 (N_19442,N_5446,N_6126);
and U19443 (N_19443,N_7670,N_601);
and U19444 (N_19444,N_8675,N_2700);
nand U19445 (N_19445,N_6704,N_2945);
or U19446 (N_19446,N_8023,N_2212);
or U19447 (N_19447,N_4389,N_4949);
xnor U19448 (N_19448,N_5112,N_3930);
nor U19449 (N_19449,N_1713,N_1079);
nor U19450 (N_19450,N_1660,N_4168);
or U19451 (N_19451,N_4356,N_4896);
or U19452 (N_19452,N_5246,N_4334);
and U19453 (N_19453,N_3617,N_3654);
or U19454 (N_19454,N_6585,N_4538);
xnor U19455 (N_19455,N_3328,N_7189);
and U19456 (N_19456,N_2321,N_4354);
nor U19457 (N_19457,N_3682,N_9311);
and U19458 (N_19458,N_3971,N_1014);
nor U19459 (N_19459,N_9704,N_6145);
nand U19460 (N_19460,N_3376,N_4100);
xor U19461 (N_19461,N_7306,N_9974);
or U19462 (N_19462,N_8368,N_6095);
xnor U19463 (N_19463,N_4732,N_6572);
or U19464 (N_19464,N_9395,N_6923);
nand U19465 (N_19465,N_9150,N_1218);
nor U19466 (N_19466,N_4278,N_4898);
or U19467 (N_19467,N_845,N_4300);
nor U19468 (N_19468,N_115,N_4);
xnor U19469 (N_19469,N_5525,N_9842);
nor U19470 (N_19470,N_7121,N_8293);
and U19471 (N_19471,N_6704,N_3438);
nand U19472 (N_19472,N_2816,N_1202);
or U19473 (N_19473,N_4166,N_724);
or U19474 (N_19474,N_4133,N_7046);
xnor U19475 (N_19475,N_5222,N_2972);
xnor U19476 (N_19476,N_3878,N_2813);
nand U19477 (N_19477,N_5938,N_6253);
or U19478 (N_19478,N_2854,N_1930);
and U19479 (N_19479,N_7601,N_1775);
or U19480 (N_19480,N_3149,N_4648);
and U19481 (N_19481,N_1051,N_9030);
xor U19482 (N_19482,N_4344,N_1937);
xnor U19483 (N_19483,N_534,N_6569);
and U19484 (N_19484,N_2936,N_3126);
xor U19485 (N_19485,N_7264,N_4176);
or U19486 (N_19486,N_3607,N_726);
nor U19487 (N_19487,N_4516,N_1688);
xor U19488 (N_19488,N_5856,N_6919);
nor U19489 (N_19489,N_8447,N_6836);
or U19490 (N_19490,N_2672,N_3499);
nand U19491 (N_19491,N_1724,N_7911);
and U19492 (N_19492,N_2427,N_8470);
nor U19493 (N_19493,N_9353,N_404);
and U19494 (N_19494,N_5170,N_888);
nand U19495 (N_19495,N_6924,N_4177);
xor U19496 (N_19496,N_5522,N_1947);
nand U19497 (N_19497,N_1904,N_3198);
or U19498 (N_19498,N_680,N_6408);
nand U19499 (N_19499,N_7734,N_9744);
nand U19500 (N_19500,N_3805,N_1569);
nor U19501 (N_19501,N_7619,N_8881);
nand U19502 (N_19502,N_3784,N_4095);
nor U19503 (N_19503,N_683,N_4586);
or U19504 (N_19504,N_7285,N_9682);
nor U19505 (N_19505,N_8597,N_7167);
and U19506 (N_19506,N_8644,N_7571);
nor U19507 (N_19507,N_823,N_7570);
xor U19508 (N_19508,N_5870,N_2623);
nor U19509 (N_19509,N_9114,N_9249);
xor U19510 (N_19510,N_1785,N_8408);
xnor U19511 (N_19511,N_3054,N_8008);
nor U19512 (N_19512,N_3087,N_1177);
and U19513 (N_19513,N_3796,N_6246);
nand U19514 (N_19514,N_2568,N_5274);
or U19515 (N_19515,N_4604,N_8520);
or U19516 (N_19516,N_2817,N_9793);
and U19517 (N_19517,N_6905,N_3668);
nand U19518 (N_19518,N_9158,N_9166);
or U19519 (N_19519,N_1700,N_9424);
xor U19520 (N_19520,N_8970,N_888);
nor U19521 (N_19521,N_1172,N_4881);
nor U19522 (N_19522,N_6466,N_8472);
nand U19523 (N_19523,N_8828,N_8184);
nor U19524 (N_19524,N_8685,N_1981);
and U19525 (N_19525,N_5309,N_1022);
or U19526 (N_19526,N_3467,N_8082);
or U19527 (N_19527,N_7014,N_3578);
nor U19528 (N_19528,N_9600,N_1081);
nand U19529 (N_19529,N_4011,N_2293);
or U19530 (N_19530,N_3702,N_4406);
and U19531 (N_19531,N_6384,N_9945);
nor U19532 (N_19532,N_644,N_8816);
or U19533 (N_19533,N_6754,N_6742);
or U19534 (N_19534,N_5579,N_3915);
and U19535 (N_19535,N_772,N_9955);
xnor U19536 (N_19536,N_3876,N_2220);
and U19537 (N_19537,N_3477,N_4368);
and U19538 (N_19538,N_7263,N_871);
or U19539 (N_19539,N_6791,N_6988);
xnor U19540 (N_19540,N_1623,N_30);
xnor U19541 (N_19541,N_3946,N_3325);
or U19542 (N_19542,N_9200,N_5903);
and U19543 (N_19543,N_1696,N_6117);
and U19544 (N_19544,N_231,N_6563);
or U19545 (N_19545,N_7226,N_2704);
nand U19546 (N_19546,N_2801,N_8849);
nand U19547 (N_19547,N_4033,N_7163);
xnor U19548 (N_19548,N_6006,N_377);
nand U19549 (N_19549,N_9161,N_3478);
xnor U19550 (N_19550,N_5585,N_2137);
and U19551 (N_19551,N_2993,N_8659);
nand U19552 (N_19552,N_3332,N_6382);
and U19553 (N_19553,N_8234,N_2717);
or U19554 (N_19554,N_1517,N_3220);
xnor U19555 (N_19555,N_4940,N_9980);
and U19556 (N_19556,N_6444,N_1095);
xnor U19557 (N_19557,N_2000,N_1452);
and U19558 (N_19558,N_2373,N_2674);
and U19559 (N_19559,N_4041,N_2489);
xnor U19560 (N_19560,N_3845,N_4792);
and U19561 (N_19561,N_2470,N_7781);
nor U19562 (N_19562,N_6881,N_7573);
and U19563 (N_19563,N_4650,N_6176);
nand U19564 (N_19564,N_889,N_7000);
and U19565 (N_19565,N_4612,N_5800);
or U19566 (N_19566,N_1131,N_7307);
xnor U19567 (N_19567,N_494,N_6908);
and U19568 (N_19568,N_3911,N_3431);
and U19569 (N_19569,N_2628,N_6865);
and U19570 (N_19570,N_5636,N_6153);
nor U19571 (N_19571,N_7838,N_405);
or U19572 (N_19572,N_1068,N_5564);
or U19573 (N_19573,N_1818,N_8989);
nand U19574 (N_19574,N_3018,N_8816);
nor U19575 (N_19575,N_9441,N_1933);
nor U19576 (N_19576,N_2755,N_7973);
or U19577 (N_19577,N_2750,N_9431);
or U19578 (N_19578,N_8108,N_4283);
xor U19579 (N_19579,N_4360,N_5781);
or U19580 (N_19580,N_9372,N_8453);
nor U19581 (N_19581,N_857,N_8187);
or U19582 (N_19582,N_5199,N_5904);
or U19583 (N_19583,N_2749,N_5381);
or U19584 (N_19584,N_1858,N_5573);
and U19585 (N_19585,N_2038,N_6340);
nand U19586 (N_19586,N_3992,N_4420);
and U19587 (N_19587,N_2910,N_9627);
xor U19588 (N_19588,N_6316,N_3133);
and U19589 (N_19589,N_5597,N_425);
or U19590 (N_19590,N_1703,N_9392);
nand U19591 (N_19591,N_4161,N_1434);
xnor U19592 (N_19592,N_8415,N_2103);
nand U19593 (N_19593,N_4296,N_7182);
nor U19594 (N_19594,N_516,N_694);
xnor U19595 (N_19595,N_3469,N_424);
and U19596 (N_19596,N_5369,N_8150);
and U19597 (N_19597,N_3123,N_7207);
or U19598 (N_19598,N_5382,N_7019);
nand U19599 (N_19599,N_8388,N_8409);
xnor U19600 (N_19600,N_1906,N_3989);
nand U19601 (N_19601,N_6392,N_9849);
or U19602 (N_19602,N_9205,N_475);
nand U19603 (N_19603,N_1013,N_4657);
nand U19604 (N_19604,N_6902,N_1196);
nand U19605 (N_19605,N_8168,N_440);
xnor U19606 (N_19606,N_8469,N_569);
xor U19607 (N_19607,N_9426,N_8275);
nor U19608 (N_19608,N_3535,N_3826);
and U19609 (N_19609,N_4751,N_2430);
or U19610 (N_19610,N_1539,N_1078);
nor U19611 (N_19611,N_4980,N_3684);
and U19612 (N_19612,N_3007,N_1133);
or U19613 (N_19613,N_6744,N_8964);
nand U19614 (N_19614,N_5441,N_634);
nand U19615 (N_19615,N_3976,N_2051);
nand U19616 (N_19616,N_7805,N_3917);
xnor U19617 (N_19617,N_7450,N_6525);
nor U19618 (N_19618,N_701,N_6645);
xor U19619 (N_19619,N_1914,N_9008);
and U19620 (N_19620,N_9699,N_768);
nor U19621 (N_19621,N_4041,N_7670);
and U19622 (N_19622,N_456,N_3738);
nor U19623 (N_19623,N_8299,N_6701);
xnor U19624 (N_19624,N_3573,N_2886);
xnor U19625 (N_19625,N_3715,N_8478);
or U19626 (N_19626,N_3898,N_5106);
or U19627 (N_19627,N_8088,N_2455);
nor U19628 (N_19628,N_1481,N_9223);
nor U19629 (N_19629,N_4175,N_7554);
nand U19630 (N_19630,N_572,N_2252);
xor U19631 (N_19631,N_7756,N_7937);
xnor U19632 (N_19632,N_9968,N_8568);
or U19633 (N_19633,N_7745,N_6044);
nor U19634 (N_19634,N_7848,N_9183);
and U19635 (N_19635,N_893,N_1237);
nand U19636 (N_19636,N_7474,N_8415);
xnor U19637 (N_19637,N_2207,N_3746);
xnor U19638 (N_19638,N_4703,N_3622);
or U19639 (N_19639,N_5015,N_7389);
nand U19640 (N_19640,N_6523,N_2022);
nand U19641 (N_19641,N_4728,N_8188);
nand U19642 (N_19642,N_1398,N_7596);
xor U19643 (N_19643,N_173,N_9828);
nor U19644 (N_19644,N_7057,N_7072);
nand U19645 (N_19645,N_3009,N_2545);
nor U19646 (N_19646,N_3288,N_4678);
and U19647 (N_19647,N_9434,N_8559);
xnor U19648 (N_19648,N_6864,N_7203);
nor U19649 (N_19649,N_4949,N_9165);
nand U19650 (N_19650,N_4842,N_7313);
xor U19651 (N_19651,N_488,N_4370);
nor U19652 (N_19652,N_8887,N_776);
nand U19653 (N_19653,N_911,N_1877);
and U19654 (N_19654,N_1183,N_5799);
and U19655 (N_19655,N_9335,N_2477);
and U19656 (N_19656,N_9226,N_1697);
and U19657 (N_19657,N_3402,N_6508);
and U19658 (N_19658,N_79,N_6159);
and U19659 (N_19659,N_4281,N_8361);
xnor U19660 (N_19660,N_3986,N_7749);
nor U19661 (N_19661,N_4895,N_8899);
xor U19662 (N_19662,N_7258,N_2266);
and U19663 (N_19663,N_9856,N_6354);
nand U19664 (N_19664,N_6628,N_8090);
xnor U19665 (N_19665,N_9511,N_3450);
nor U19666 (N_19666,N_8347,N_1134);
or U19667 (N_19667,N_5833,N_5368);
nand U19668 (N_19668,N_7897,N_3584);
xor U19669 (N_19669,N_8515,N_9021);
nor U19670 (N_19670,N_8761,N_3800);
nand U19671 (N_19671,N_5060,N_7762);
nor U19672 (N_19672,N_2129,N_1282);
nor U19673 (N_19673,N_5870,N_2799);
and U19674 (N_19674,N_8523,N_3917);
and U19675 (N_19675,N_668,N_5412);
and U19676 (N_19676,N_5508,N_7699);
and U19677 (N_19677,N_3371,N_1500);
or U19678 (N_19678,N_2756,N_9016);
xnor U19679 (N_19679,N_3924,N_8043);
nor U19680 (N_19680,N_661,N_89);
nor U19681 (N_19681,N_7244,N_2413);
nand U19682 (N_19682,N_7521,N_1974);
nor U19683 (N_19683,N_56,N_2983);
or U19684 (N_19684,N_2830,N_6118);
or U19685 (N_19685,N_352,N_1129);
xnor U19686 (N_19686,N_4060,N_8676);
and U19687 (N_19687,N_2262,N_9696);
or U19688 (N_19688,N_1142,N_4379);
nand U19689 (N_19689,N_6949,N_2489);
xor U19690 (N_19690,N_5327,N_2179);
nand U19691 (N_19691,N_9750,N_6183);
xor U19692 (N_19692,N_2323,N_318);
nand U19693 (N_19693,N_7343,N_134);
nand U19694 (N_19694,N_2363,N_4446);
or U19695 (N_19695,N_408,N_9202);
nand U19696 (N_19696,N_1522,N_8985);
or U19697 (N_19697,N_1646,N_165);
and U19698 (N_19698,N_785,N_924);
and U19699 (N_19699,N_1210,N_6847);
nand U19700 (N_19700,N_4441,N_9151);
and U19701 (N_19701,N_8043,N_4413);
and U19702 (N_19702,N_4387,N_3892);
nor U19703 (N_19703,N_6148,N_3596);
nor U19704 (N_19704,N_693,N_6450);
or U19705 (N_19705,N_9596,N_8047);
or U19706 (N_19706,N_4079,N_4299);
nor U19707 (N_19707,N_451,N_5542);
nor U19708 (N_19708,N_2687,N_9569);
nand U19709 (N_19709,N_1125,N_623);
or U19710 (N_19710,N_5291,N_3543);
nor U19711 (N_19711,N_9333,N_4383);
or U19712 (N_19712,N_3170,N_1066);
nand U19713 (N_19713,N_844,N_1487);
xnor U19714 (N_19714,N_4262,N_2768);
and U19715 (N_19715,N_7010,N_6834);
and U19716 (N_19716,N_9374,N_2274);
nor U19717 (N_19717,N_8347,N_5909);
nand U19718 (N_19718,N_4534,N_3247);
nor U19719 (N_19719,N_845,N_9721);
nand U19720 (N_19720,N_3650,N_3616);
or U19721 (N_19721,N_9055,N_1701);
nand U19722 (N_19722,N_4379,N_1899);
or U19723 (N_19723,N_7384,N_151);
nor U19724 (N_19724,N_8556,N_1355);
or U19725 (N_19725,N_9467,N_3046);
and U19726 (N_19726,N_3269,N_7225);
and U19727 (N_19727,N_2578,N_3867);
xor U19728 (N_19728,N_4845,N_6516);
nand U19729 (N_19729,N_723,N_696);
nand U19730 (N_19730,N_306,N_7621);
nor U19731 (N_19731,N_5515,N_3376);
and U19732 (N_19732,N_875,N_6393);
xor U19733 (N_19733,N_1912,N_6526);
and U19734 (N_19734,N_5782,N_5965);
xor U19735 (N_19735,N_8767,N_7431);
xor U19736 (N_19736,N_5728,N_1511);
nand U19737 (N_19737,N_9590,N_350);
and U19738 (N_19738,N_3139,N_585);
and U19739 (N_19739,N_1874,N_7597);
nand U19740 (N_19740,N_3873,N_1890);
nand U19741 (N_19741,N_4110,N_4523);
xor U19742 (N_19742,N_5874,N_1187);
and U19743 (N_19743,N_1278,N_924);
nand U19744 (N_19744,N_6009,N_4807);
or U19745 (N_19745,N_1800,N_2613);
nor U19746 (N_19746,N_3702,N_9619);
nand U19747 (N_19747,N_6953,N_9242);
and U19748 (N_19748,N_4298,N_3932);
nand U19749 (N_19749,N_2551,N_5799);
and U19750 (N_19750,N_6536,N_8056);
and U19751 (N_19751,N_9836,N_9470);
and U19752 (N_19752,N_1018,N_2436);
nand U19753 (N_19753,N_1399,N_5959);
nand U19754 (N_19754,N_5,N_8522);
nor U19755 (N_19755,N_6991,N_45);
and U19756 (N_19756,N_2954,N_570);
nor U19757 (N_19757,N_5461,N_1895);
xnor U19758 (N_19758,N_6595,N_2914);
or U19759 (N_19759,N_3925,N_2736);
xor U19760 (N_19760,N_7394,N_5588);
and U19761 (N_19761,N_1490,N_8038);
nand U19762 (N_19762,N_6595,N_1502);
xnor U19763 (N_19763,N_9445,N_8098);
and U19764 (N_19764,N_2813,N_9511);
nand U19765 (N_19765,N_184,N_4627);
or U19766 (N_19766,N_7952,N_4098);
or U19767 (N_19767,N_3492,N_4773);
xor U19768 (N_19768,N_8051,N_4639);
xor U19769 (N_19769,N_9701,N_5790);
and U19770 (N_19770,N_2115,N_8469);
nand U19771 (N_19771,N_7132,N_5019);
nand U19772 (N_19772,N_9564,N_271);
nand U19773 (N_19773,N_2761,N_1225);
nor U19774 (N_19774,N_9110,N_6710);
xnor U19775 (N_19775,N_2804,N_1802);
nand U19776 (N_19776,N_1210,N_2747);
nand U19777 (N_19777,N_7037,N_1909);
nand U19778 (N_19778,N_9211,N_382);
or U19779 (N_19779,N_5896,N_1065);
or U19780 (N_19780,N_7374,N_4);
nand U19781 (N_19781,N_3764,N_7987);
and U19782 (N_19782,N_7447,N_3878);
nor U19783 (N_19783,N_5771,N_3257);
nor U19784 (N_19784,N_3971,N_577);
xnor U19785 (N_19785,N_8004,N_8772);
xnor U19786 (N_19786,N_495,N_7740);
xor U19787 (N_19787,N_7774,N_2188);
or U19788 (N_19788,N_1933,N_2212);
or U19789 (N_19789,N_7803,N_2285);
nand U19790 (N_19790,N_5458,N_9733);
xor U19791 (N_19791,N_4171,N_9971);
nand U19792 (N_19792,N_5842,N_4487);
or U19793 (N_19793,N_4196,N_7061);
nand U19794 (N_19794,N_4987,N_2135);
and U19795 (N_19795,N_4059,N_4400);
nand U19796 (N_19796,N_6494,N_8882);
or U19797 (N_19797,N_8171,N_3562);
nand U19798 (N_19798,N_2233,N_4163);
nor U19799 (N_19799,N_1092,N_8531);
xnor U19800 (N_19800,N_9899,N_3707);
nand U19801 (N_19801,N_1212,N_3795);
and U19802 (N_19802,N_6006,N_5756);
xor U19803 (N_19803,N_221,N_1229);
or U19804 (N_19804,N_6141,N_7512);
and U19805 (N_19805,N_5373,N_1140);
and U19806 (N_19806,N_1360,N_809);
nor U19807 (N_19807,N_7205,N_8240);
nor U19808 (N_19808,N_8670,N_9748);
or U19809 (N_19809,N_4754,N_4470);
xnor U19810 (N_19810,N_834,N_7078);
nand U19811 (N_19811,N_1,N_2224);
xnor U19812 (N_19812,N_130,N_6305);
and U19813 (N_19813,N_4426,N_8980);
nand U19814 (N_19814,N_7269,N_485);
xor U19815 (N_19815,N_1304,N_3615);
nor U19816 (N_19816,N_2819,N_3776);
and U19817 (N_19817,N_5835,N_2766);
and U19818 (N_19818,N_6834,N_8085);
or U19819 (N_19819,N_5252,N_5475);
and U19820 (N_19820,N_6175,N_7467);
and U19821 (N_19821,N_7667,N_253);
nand U19822 (N_19822,N_8516,N_7264);
nand U19823 (N_19823,N_9395,N_4443);
or U19824 (N_19824,N_9566,N_4777);
xnor U19825 (N_19825,N_8639,N_2919);
and U19826 (N_19826,N_8831,N_8931);
nand U19827 (N_19827,N_5741,N_2917);
or U19828 (N_19828,N_2120,N_5517);
xor U19829 (N_19829,N_9701,N_1503);
nand U19830 (N_19830,N_8439,N_6271);
and U19831 (N_19831,N_3386,N_6391);
xnor U19832 (N_19832,N_8302,N_3336);
nand U19833 (N_19833,N_2812,N_7650);
and U19834 (N_19834,N_1580,N_969);
nor U19835 (N_19835,N_9975,N_6390);
and U19836 (N_19836,N_5811,N_43);
nor U19837 (N_19837,N_7615,N_735);
and U19838 (N_19838,N_963,N_5428);
nor U19839 (N_19839,N_491,N_1913);
nor U19840 (N_19840,N_3819,N_2053);
and U19841 (N_19841,N_4765,N_7678);
or U19842 (N_19842,N_4910,N_6647);
nand U19843 (N_19843,N_9395,N_1842);
nand U19844 (N_19844,N_6261,N_2672);
nor U19845 (N_19845,N_5778,N_9439);
xnor U19846 (N_19846,N_3009,N_4001);
or U19847 (N_19847,N_9232,N_1080);
xor U19848 (N_19848,N_450,N_3806);
nand U19849 (N_19849,N_9525,N_5992);
or U19850 (N_19850,N_1104,N_9667);
or U19851 (N_19851,N_6513,N_6883);
and U19852 (N_19852,N_1224,N_1187);
or U19853 (N_19853,N_5774,N_9263);
nand U19854 (N_19854,N_2173,N_8448);
nand U19855 (N_19855,N_3988,N_3139);
nor U19856 (N_19856,N_2008,N_9139);
and U19857 (N_19857,N_4444,N_4256);
nor U19858 (N_19858,N_2227,N_6282);
nand U19859 (N_19859,N_9342,N_3367);
or U19860 (N_19860,N_4784,N_5301);
xnor U19861 (N_19861,N_9294,N_4068);
or U19862 (N_19862,N_9961,N_6927);
and U19863 (N_19863,N_4733,N_510);
nand U19864 (N_19864,N_986,N_3204);
nand U19865 (N_19865,N_435,N_5616);
or U19866 (N_19866,N_3248,N_5585);
nor U19867 (N_19867,N_2519,N_7877);
and U19868 (N_19868,N_2983,N_5058);
nand U19869 (N_19869,N_3682,N_532);
or U19870 (N_19870,N_3845,N_6872);
xor U19871 (N_19871,N_2137,N_8231);
nand U19872 (N_19872,N_3236,N_8355);
nor U19873 (N_19873,N_3330,N_9797);
nor U19874 (N_19874,N_2073,N_7797);
xor U19875 (N_19875,N_362,N_7756);
and U19876 (N_19876,N_5690,N_8058);
nand U19877 (N_19877,N_5501,N_3497);
nor U19878 (N_19878,N_9877,N_4365);
and U19879 (N_19879,N_1944,N_5063);
and U19880 (N_19880,N_1721,N_6764);
nor U19881 (N_19881,N_9904,N_9638);
nand U19882 (N_19882,N_1663,N_5807);
nor U19883 (N_19883,N_6168,N_185);
nor U19884 (N_19884,N_9241,N_6733);
or U19885 (N_19885,N_4490,N_4792);
and U19886 (N_19886,N_1479,N_4310);
nor U19887 (N_19887,N_6957,N_7779);
nand U19888 (N_19888,N_5925,N_6372);
nor U19889 (N_19889,N_8620,N_2434);
nand U19890 (N_19890,N_8554,N_9717);
or U19891 (N_19891,N_8295,N_5172);
and U19892 (N_19892,N_5332,N_9306);
and U19893 (N_19893,N_9298,N_4531);
nand U19894 (N_19894,N_236,N_4456);
or U19895 (N_19895,N_4847,N_1983);
xnor U19896 (N_19896,N_5152,N_3075);
nand U19897 (N_19897,N_2813,N_3176);
and U19898 (N_19898,N_5191,N_8745);
nor U19899 (N_19899,N_9183,N_1802);
nand U19900 (N_19900,N_7535,N_8922);
xnor U19901 (N_19901,N_4962,N_4704);
and U19902 (N_19902,N_1412,N_7028);
nor U19903 (N_19903,N_8640,N_4208);
and U19904 (N_19904,N_6120,N_2603);
nor U19905 (N_19905,N_6062,N_8055);
and U19906 (N_19906,N_3909,N_8461);
and U19907 (N_19907,N_4320,N_2587);
nor U19908 (N_19908,N_1679,N_3867);
and U19909 (N_19909,N_8688,N_4443);
nand U19910 (N_19910,N_1444,N_1243);
nand U19911 (N_19911,N_3336,N_7169);
nor U19912 (N_19912,N_9592,N_8862);
and U19913 (N_19913,N_5695,N_2328);
nor U19914 (N_19914,N_4481,N_77);
nand U19915 (N_19915,N_5466,N_1935);
or U19916 (N_19916,N_6176,N_4276);
nor U19917 (N_19917,N_2744,N_8636);
and U19918 (N_19918,N_1527,N_5215);
nor U19919 (N_19919,N_2163,N_1995);
and U19920 (N_19920,N_923,N_8362);
and U19921 (N_19921,N_2829,N_1831);
or U19922 (N_19922,N_7698,N_5450);
and U19923 (N_19923,N_833,N_5514);
xnor U19924 (N_19924,N_1114,N_6704);
or U19925 (N_19925,N_412,N_4559);
xnor U19926 (N_19926,N_4285,N_4446);
xor U19927 (N_19927,N_2748,N_8654);
nor U19928 (N_19928,N_1746,N_8620);
nor U19929 (N_19929,N_5524,N_7805);
and U19930 (N_19930,N_2952,N_5759);
or U19931 (N_19931,N_5107,N_1370);
nand U19932 (N_19932,N_3020,N_8331);
nor U19933 (N_19933,N_5607,N_2170);
or U19934 (N_19934,N_4046,N_9610);
or U19935 (N_19935,N_1318,N_134);
nand U19936 (N_19936,N_7273,N_2082);
nor U19937 (N_19937,N_8157,N_7197);
xnor U19938 (N_19938,N_5896,N_7185);
nor U19939 (N_19939,N_8792,N_4567);
nand U19940 (N_19940,N_7384,N_2244);
and U19941 (N_19941,N_7522,N_1323);
nor U19942 (N_19942,N_4757,N_2841);
and U19943 (N_19943,N_9002,N_2229);
nand U19944 (N_19944,N_2321,N_1947);
nor U19945 (N_19945,N_7298,N_1854);
or U19946 (N_19946,N_1856,N_4637);
and U19947 (N_19947,N_4587,N_1578);
nor U19948 (N_19948,N_7421,N_9742);
xor U19949 (N_19949,N_7266,N_8885);
or U19950 (N_19950,N_9018,N_7547);
xnor U19951 (N_19951,N_4399,N_4483);
nand U19952 (N_19952,N_4752,N_957);
nor U19953 (N_19953,N_3324,N_9554);
xnor U19954 (N_19954,N_8526,N_8451);
and U19955 (N_19955,N_2779,N_3929);
and U19956 (N_19956,N_9968,N_5399);
nor U19957 (N_19957,N_9579,N_6023);
and U19958 (N_19958,N_3900,N_3540);
and U19959 (N_19959,N_5055,N_6349);
nand U19960 (N_19960,N_9420,N_5338);
or U19961 (N_19961,N_4668,N_1929);
and U19962 (N_19962,N_8017,N_3459);
and U19963 (N_19963,N_732,N_8650);
nand U19964 (N_19964,N_5834,N_5034);
or U19965 (N_19965,N_2140,N_6135);
nand U19966 (N_19966,N_9078,N_224);
and U19967 (N_19967,N_8823,N_9594);
and U19968 (N_19968,N_6940,N_3473);
or U19969 (N_19969,N_2427,N_4344);
nor U19970 (N_19970,N_8065,N_5329);
nor U19971 (N_19971,N_284,N_3335);
xnor U19972 (N_19972,N_3555,N_9054);
xnor U19973 (N_19973,N_2986,N_7261);
or U19974 (N_19974,N_6900,N_8071);
or U19975 (N_19975,N_6580,N_516);
and U19976 (N_19976,N_7843,N_3026);
and U19977 (N_19977,N_5912,N_9617);
xor U19978 (N_19978,N_2268,N_5688);
xor U19979 (N_19979,N_7548,N_7312);
or U19980 (N_19980,N_4467,N_6994);
or U19981 (N_19981,N_4719,N_5688);
xor U19982 (N_19982,N_1506,N_6396);
nand U19983 (N_19983,N_747,N_1788);
or U19984 (N_19984,N_2603,N_5587);
nor U19985 (N_19985,N_8935,N_4618);
nor U19986 (N_19986,N_1860,N_5315);
nand U19987 (N_19987,N_1672,N_4957);
and U19988 (N_19988,N_6685,N_6413);
or U19989 (N_19989,N_4283,N_8273);
and U19990 (N_19990,N_7516,N_2156);
xor U19991 (N_19991,N_1631,N_1111);
nor U19992 (N_19992,N_3197,N_9135);
or U19993 (N_19993,N_9526,N_3581);
and U19994 (N_19994,N_3388,N_1884);
nor U19995 (N_19995,N_4881,N_8645);
or U19996 (N_19996,N_9493,N_5798);
nor U19997 (N_19997,N_3965,N_179);
or U19998 (N_19998,N_7201,N_1102);
and U19999 (N_19999,N_8311,N_1452);
and U20000 (N_20000,N_17667,N_15107);
nand U20001 (N_20001,N_13935,N_12310);
xnor U20002 (N_20002,N_10481,N_15148);
nand U20003 (N_20003,N_15787,N_18181);
nand U20004 (N_20004,N_19888,N_13805);
and U20005 (N_20005,N_12529,N_14501);
nand U20006 (N_20006,N_11782,N_18476);
and U20007 (N_20007,N_15513,N_11634);
xnor U20008 (N_20008,N_18091,N_13178);
nand U20009 (N_20009,N_10523,N_14919);
and U20010 (N_20010,N_11661,N_13361);
or U20011 (N_20011,N_19668,N_10841);
or U20012 (N_20012,N_13594,N_16327);
nor U20013 (N_20013,N_10688,N_17446);
and U20014 (N_20014,N_16809,N_11619);
nor U20015 (N_20015,N_17485,N_14455);
or U20016 (N_20016,N_12641,N_13433);
or U20017 (N_20017,N_17101,N_15689);
nor U20018 (N_20018,N_12646,N_18500);
nand U20019 (N_20019,N_17546,N_18225);
nand U20020 (N_20020,N_18932,N_15357);
nor U20021 (N_20021,N_18051,N_10594);
or U20022 (N_20022,N_14130,N_13092);
xnor U20023 (N_20023,N_17879,N_17695);
xor U20024 (N_20024,N_12834,N_18565);
nor U20025 (N_20025,N_15997,N_19617);
nor U20026 (N_20026,N_12260,N_10072);
xor U20027 (N_20027,N_12425,N_17209);
nor U20028 (N_20028,N_15356,N_12986);
xnor U20029 (N_20029,N_11385,N_17480);
xor U20030 (N_20030,N_16708,N_10729);
nor U20031 (N_20031,N_18551,N_10458);
nand U20032 (N_20032,N_15003,N_13014);
nor U20033 (N_20033,N_10805,N_12665);
xnor U20034 (N_20034,N_16016,N_17532);
nor U20035 (N_20035,N_10368,N_17378);
xor U20036 (N_20036,N_10660,N_17720);
nor U20037 (N_20037,N_12824,N_11047);
xor U20038 (N_20038,N_19581,N_12637);
nor U20039 (N_20039,N_16038,N_19071);
xnor U20040 (N_20040,N_18784,N_19164);
xnor U20041 (N_20041,N_13952,N_10727);
and U20042 (N_20042,N_17904,N_14038);
xor U20043 (N_20043,N_10721,N_14494);
xor U20044 (N_20044,N_14562,N_17211);
and U20045 (N_20045,N_18252,N_19009);
nand U20046 (N_20046,N_12912,N_16231);
nor U20047 (N_20047,N_14219,N_17452);
and U20048 (N_20048,N_18077,N_10899);
or U20049 (N_20049,N_16273,N_19502);
and U20050 (N_20050,N_10034,N_13889);
xor U20051 (N_20051,N_11396,N_15273);
nand U20052 (N_20052,N_11110,N_13293);
and U20053 (N_20053,N_13803,N_12569);
nor U20054 (N_20054,N_15136,N_12506);
xor U20055 (N_20055,N_17630,N_18199);
nor U20056 (N_20056,N_10040,N_13714);
or U20057 (N_20057,N_14517,N_14449);
nor U20058 (N_20058,N_17028,N_14350);
and U20059 (N_20059,N_19969,N_15955);
or U20060 (N_20060,N_16101,N_18789);
and U20061 (N_20061,N_17212,N_11698);
or U20062 (N_20062,N_14771,N_19355);
nor U20063 (N_20063,N_10775,N_14278);
nor U20064 (N_20064,N_15945,N_14854);
xnor U20065 (N_20065,N_17748,N_15457);
xnor U20066 (N_20066,N_18674,N_17511);
and U20067 (N_20067,N_16898,N_19674);
and U20068 (N_20068,N_16958,N_11163);
nand U20069 (N_20069,N_14025,N_12890);
nor U20070 (N_20070,N_14031,N_10529);
nand U20071 (N_20071,N_13955,N_15954);
xor U20072 (N_20072,N_13584,N_14266);
xor U20073 (N_20073,N_13601,N_13420);
nor U20074 (N_20074,N_16375,N_13945);
and U20075 (N_20075,N_16578,N_17204);
or U20076 (N_20076,N_12178,N_18765);
and U20077 (N_20077,N_14955,N_11361);
nand U20078 (N_20078,N_17769,N_17268);
or U20079 (N_20079,N_14106,N_12645);
and U20080 (N_20080,N_17289,N_19138);
xor U20081 (N_20081,N_16308,N_19681);
and U20082 (N_20082,N_14186,N_15619);
nand U20083 (N_20083,N_19500,N_13432);
xor U20084 (N_20084,N_14468,N_19191);
or U20085 (N_20085,N_15151,N_17704);
xor U20086 (N_20086,N_18285,N_16936);
nor U20087 (N_20087,N_19454,N_16564);
nand U20088 (N_20088,N_10090,N_10960);
nor U20089 (N_20089,N_16501,N_19889);
xor U20090 (N_20090,N_17399,N_13621);
xor U20091 (N_20091,N_17321,N_14982);
xor U20092 (N_20092,N_11359,N_14704);
or U20093 (N_20093,N_16853,N_15962);
and U20094 (N_20094,N_15564,N_11194);
nand U20095 (N_20095,N_18716,N_19045);
or U20096 (N_20096,N_14333,N_12736);
xnor U20097 (N_20097,N_12317,N_13969);
and U20098 (N_20098,N_15805,N_12988);
xor U20099 (N_20099,N_16609,N_16351);
xnor U20100 (N_20100,N_12672,N_12363);
nor U20101 (N_20101,N_13521,N_18717);
xnor U20102 (N_20102,N_18957,N_12288);
nand U20103 (N_20103,N_17523,N_16746);
and U20104 (N_20104,N_18368,N_12566);
xnor U20105 (N_20105,N_13457,N_13468);
nor U20106 (N_20106,N_17729,N_12617);
nand U20107 (N_20107,N_14353,N_13681);
or U20108 (N_20108,N_12253,N_16493);
nor U20109 (N_20109,N_18188,N_15963);
or U20110 (N_20110,N_11656,N_18652);
nand U20111 (N_20111,N_16703,N_12530);
or U20112 (N_20112,N_16434,N_18012);
or U20113 (N_20113,N_13798,N_11020);
or U20114 (N_20114,N_18136,N_16342);
or U20115 (N_20115,N_19169,N_14240);
and U20116 (N_20116,N_15422,N_14367);
or U20117 (N_20117,N_12698,N_12459);
xor U20118 (N_20118,N_16255,N_14467);
and U20119 (N_20119,N_13400,N_11894);
and U20120 (N_20120,N_16837,N_13698);
nor U20121 (N_20121,N_13831,N_14875);
xnor U20122 (N_20122,N_17730,N_13458);
xor U20123 (N_20123,N_11864,N_10946);
nor U20124 (N_20124,N_13346,N_19086);
nand U20125 (N_20125,N_18171,N_11799);
xnor U20126 (N_20126,N_12446,N_16543);
nor U20127 (N_20127,N_19053,N_12842);
nand U20128 (N_20128,N_19096,N_11990);
and U20129 (N_20129,N_18211,N_17615);
or U20130 (N_20130,N_19363,N_12345);
or U20131 (N_20131,N_12136,N_16668);
nor U20132 (N_20132,N_16435,N_16686);
xor U20133 (N_20133,N_14226,N_10916);
xnor U20134 (N_20134,N_17296,N_10086);
nor U20135 (N_20135,N_14845,N_18631);
xnor U20136 (N_20136,N_17059,N_13058);
nand U20137 (N_20137,N_13970,N_18447);
nor U20138 (N_20138,N_13983,N_11065);
nor U20139 (N_20139,N_10978,N_11810);
nor U20140 (N_20140,N_19115,N_14989);
or U20141 (N_20141,N_11026,N_14580);
nand U20142 (N_20142,N_16863,N_10754);
and U20143 (N_20143,N_18793,N_11477);
or U20144 (N_20144,N_12725,N_16365);
or U20145 (N_20145,N_10622,N_13622);
xnor U20146 (N_20146,N_18248,N_16053);
nand U20147 (N_20147,N_14486,N_14548);
nand U20148 (N_20148,N_11002,N_19923);
xor U20149 (N_20149,N_17120,N_11621);
nor U20150 (N_20150,N_16116,N_16724);
and U20151 (N_20151,N_15669,N_13144);
nor U20152 (N_20152,N_10527,N_18769);
and U20153 (N_20153,N_14934,N_11718);
and U20154 (N_20154,N_11583,N_11560);
nor U20155 (N_20155,N_12657,N_10939);
nor U20156 (N_20156,N_16331,N_18456);
or U20157 (N_20157,N_13909,N_10212);
nor U20158 (N_20158,N_18408,N_11476);
or U20159 (N_20159,N_12972,N_12396);
nand U20160 (N_20160,N_19741,N_18469);
or U20161 (N_20161,N_16326,N_14487);
nand U20162 (N_20162,N_10552,N_13115);
nand U20163 (N_20163,N_13322,N_18223);
nor U20164 (N_20164,N_17562,N_15800);
xor U20165 (N_20165,N_11084,N_18630);
nand U20166 (N_20166,N_19220,N_15578);
nand U20167 (N_20167,N_16887,N_17409);
and U20168 (N_20168,N_10890,N_15705);
or U20169 (N_20169,N_11681,N_17244);
and U20170 (N_20170,N_14034,N_18045);
and U20171 (N_20171,N_15936,N_14198);
xor U20172 (N_20172,N_19544,N_19588);
xor U20173 (N_20173,N_16479,N_11496);
nor U20174 (N_20174,N_10993,N_11165);
and U20175 (N_20175,N_15743,N_11161);
or U20176 (N_20176,N_18217,N_17880);
or U20177 (N_20177,N_17358,N_18909);
nor U20178 (N_20178,N_14066,N_13964);
nand U20179 (N_20179,N_10177,N_11734);
nor U20180 (N_20180,N_13456,N_19409);
or U20181 (N_20181,N_13606,N_17081);
or U20182 (N_20182,N_14737,N_12938);
and U20183 (N_20183,N_12717,N_13228);
or U20184 (N_20184,N_16146,N_12733);
and U20185 (N_20185,N_18926,N_14175);
nand U20186 (N_20186,N_15106,N_18546);
nand U20187 (N_20187,N_14585,N_19628);
nor U20188 (N_20188,N_15629,N_16256);
or U20189 (N_20189,N_18669,N_16183);
nand U20190 (N_20190,N_18907,N_15694);
nand U20191 (N_20191,N_12026,N_10892);
or U20192 (N_20192,N_11828,N_16368);
or U20193 (N_20193,N_14132,N_17586);
and U20194 (N_20194,N_18537,N_10068);
nand U20195 (N_20195,N_17915,N_14702);
and U20196 (N_20196,N_16725,N_17533);
or U20197 (N_20197,N_12847,N_19465);
or U20198 (N_20198,N_17950,N_15056);
xor U20199 (N_20199,N_16426,N_12673);
nand U20200 (N_20200,N_17148,N_12703);
xor U20201 (N_20201,N_10706,N_14250);
nor U20202 (N_20202,N_10346,N_16834);
and U20203 (N_20203,N_12518,N_13286);
and U20204 (N_20204,N_14684,N_16496);
nor U20205 (N_20205,N_15200,N_11048);
or U20206 (N_20206,N_18759,N_15341);
or U20207 (N_20207,N_13929,N_17738);
nor U20208 (N_20208,N_15112,N_12435);
or U20209 (N_20209,N_19898,N_17411);
nand U20210 (N_20210,N_14605,N_11334);
xnor U20211 (N_20211,N_12785,N_13263);
or U20212 (N_20212,N_18421,N_14165);
and U20213 (N_20213,N_12454,N_12831);
or U20214 (N_20214,N_13347,N_10113);
or U20215 (N_20215,N_17080,N_15172);
or U20216 (N_20216,N_17288,N_16645);
nor U20217 (N_20217,N_18756,N_15659);
xor U20218 (N_20218,N_11430,N_16597);
or U20219 (N_20219,N_16133,N_15060);
xor U20220 (N_20220,N_18379,N_10145);
xnor U20221 (N_20221,N_10102,N_16614);
and U20222 (N_20222,N_12587,N_17697);
nor U20223 (N_20223,N_17299,N_16570);
and U20224 (N_20224,N_15114,N_19007);
nand U20225 (N_20225,N_10613,N_14389);
xnor U20226 (N_20226,N_19925,N_14326);
or U20227 (N_20227,N_10653,N_15423);
nor U20228 (N_20228,N_12302,N_19918);
nor U20229 (N_20229,N_12949,N_17518);
xnor U20230 (N_20230,N_19101,N_18676);
xnor U20231 (N_20231,N_16254,N_19715);
or U20232 (N_20232,N_12165,N_11257);
nand U20233 (N_20233,N_19256,N_10907);
and U20234 (N_20234,N_13037,N_13541);
nand U20235 (N_20235,N_17044,N_12947);
nand U20236 (N_20236,N_12577,N_14530);
xnor U20237 (N_20237,N_15517,N_12752);
or U20238 (N_20238,N_14003,N_11957);
and U20239 (N_20239,N_17144,N_11053);
and U20240 (N_20240,N_13990,N_17351);
and U20241 (N_20241,N_15140,N_11001);
xnor U20242 (N_20242,N_19232,N_10099);
or U20243 (N_20243,N_12353,N_18958);
nor U20244 (N_20244,N_10711,N_13630);
nor U20245 (N_20245,N_18415,N_19054);
nor U20246 (N_20246,N_11932,N_18412);
nor U20247 (N_20247,N_13550,N_16923);
nand U20248 (N_20248,N_14414,N_10704);
and U20249 (N_20249,N_14951,N_12203);
nor U20250 (N_20250,N_14541,N_19672);
nand U20251 (N_20251,N_19675,N_11684);
nand U20252 (N_20252,N_16557,N_16820);
nor U20253 (N_20253,N_10741,N_17701);
nand U20254 (N_20254,N_19903,N_12366);
nor U20255 (N_20255,N_12311,N_17319);
or U20256 (N_20256,N_10645,N_19266);
or U20257 (N_20257,N_18267,N_14613);
or U20258 (N_20258,N_10745,N_12862);
and U20259 (N_20259,N_17672,N_18956);
nor U20260 (N_20260,N_15392,N_15053);
nand U20261 (N_20261,N_17669,N_14818);
nor U20262 (N_20262,N_15548,N_10845);
xnor U20263 (N_20263,N_16854,N_16006);
or U20264 (N_20264,N_18228,N_18164);
or U20265 (N_20265,N_14944,N_10384);
nand U20266 (N_20266,N_14298,N_15658);
and U20267 (N_20267,N_17483,N_19388);
xnor U20268 (N_20268,N_18915,N_14911);
nand U20269 (N_20269,N_14412,N_15735);
xor U20270 (N_20270,N_10804,N_13132);
or U20271 (N_20271,N_19439,N_18464);
nand U20272 (N_20272,N_18132,N_15985);
xor U20273 (N_20273,N_12556,N_16465);
xnor U20274 (N_20274,N_12729,N_14608);
nand U20275 (N_20275,N_18617,N_10298);
nand U20276 (N_20276,N_12922,N_16199);
nand U20277 (N_20277,N_13185,N_13069);
xor U20278 (N_20278,N_17257,N_12434);
nor U20279 (N_20279,N_11786,N_13506);
nand U20280 (N_20280,N_19257,N_19076);
or U20281 (N_20281,N_14839,N_11288);
nor U20282 (N_20282,N_10176,N_19719);
nor U20283 (N_20283,N_13476,N_15794);
and U20284 (N_20284,N_10082,N_12299);
nor U20285 (N_20285,N_14206,N_15300);
or U20286 (N_20286,N_14880,N_18999);
nand U20287 (N_20287,N_10553,N_15892);
nor U20288 (N_20288,N_16190,N_13976);
and U20289 (N_20289,N_17414,N_11275);
xor U20290 (N_20290,N_13684,N_14736);
xnor U20291 (N_20291,N_17494,N_16828);
or U20292 (N_20292,N_17371,N_15146);
xor U20293 (N_20293,N_15832,N_10353);
or U20294 (N_20294,N_11501,N_11761);
nor U20295 (N_20295,N_11401,N_12876);
xor U20296 (N_20296,N_10092,N_15228);
and U20297 (N_20297,N_13446,N_11512);
xor U20298 (N_20298,N_16353,N_11032);
or U20299 (N_20299,N_17500,N_16701);
nand U20300 (N_20300,N_14121,N_13159);
xnor U20301 (N_20301,N_19429,N_13104);
xor U20302 (N_20302,N_13135,N_14050);
nand U20303 (N_20303,N_10950,N_13974);
or U20304 (N_20304,N_16730,N_16644);
and U20305 (N_20305,N_13332,N_18362);
nand U20306 (N_20306,N_12830,N_18840);
and U20307 (N_20307,N_18076,N_10784);
or U20308 (N_20308,N_19999,N_10896);
and U20309 (N_20309,N_14103,N_19676);
nor U20310 (N_20310,N_12496,N_13063);
or U20311 (N_20311,N_14232,N_19995);
or U20312 (N_20312,N_18155,N_12067);
nor U20313 (N_20313,N_13150,N_14427);
nand U20314 (N_20314,N_11663,N_19735);
and U20315 (N_20315,N_11788,N_17812);
and U20316 (N_20316,N_11057,N_18080);
and U20317 (N_20317,N_14840,N_10383);
or U20318 (N_20318,N_12009,N_12962);
nand U20319 (N_20319,N_14471,N_17187);
and U20320 (N_20320,N_15309,N_19827);
nand U20321 (N_20321,N_12368,N_12813);
nor U20322 (N_20322,N_19141,N_14531);
xnor U20323 (N_20323,N_18427,N_17974);
nor U20324 (N_20324,N_12534,N_11915);
nor U20325 (N_20325,N_13327,N_12282);
and U20326 (N_20326,N_12559,N_12533);
nor U20327 (N_20327,N_13598,N_19089);
nor U20328 (N_20328,N_13992,N_13140);
or U20329 (N_20329,N_12854,N_10365);
or U20330 (N_20330,N_13398,N_15443);
or U20331 (N_20331,N_18811,N_15968);
xnor U20332 (N_20332,N_18745,N_19954);
and U20333 (N_20333,N_12217,N_14286);
xnor U20334 (N_20334,N_12404,N_17393);
or U20335 (N_20335,N_19847,N_13833);
or U20336 (N_20336,N_12960,N_16604);
or U20337 (N_20337,N_12272,N_16228);
xor U20338 (N_20338,N_12971,N_13816);
and U20339 (N_20339,N_10370,N_11878);
nor U20340 (N_20340,N_16525,N_16343);
nand U20341 (N_20341,N_12380,N_13762);
xnor U20342 (N_20342,N_13891,N_10042);
or U20343 (N_20343,N_15647,N_13657);
nand U20344 (N_20344,N_17646,N_10101);
or U20345 (N_20345,N_19706,N_13100);
or U20346 (N_20346,N_17932,N_11751);
nand U20347 (N_20347,N_19962,N_19655);
or U20348 (N_20348,N_16611,N_14212);
or U20349 (N_20349,N_11499,N_11931);
xor U20350 (N_20350,N_19952,N_10675);
nor U20351 (N_20351,N_19828,N_13326);
and U20352 (N_20352,N_13291,N_15169);
nand U20353 (N_20353,N_13647,N_12924);
xor U20354 (N_20354,N_18397,N_14971);
and U20355 (N_20355,N_17800,N_15662);
or U20356 (N_20356,N_16013,N_11096);
and U20357 (N_20357,N_14921,N_10794);
or U20358 (N_20358,N_16278,N_14281);
nand U20359 (N_20359,N_16558,N_16077);
and U20360 (N_20360,N_14394,N_16941);
and U20361 (N_20361,N_18702,N_17628);
and U20362 (N_20362,N_14368,N_17350);
nand U20363 (N_20363,N_17275,N_18786);
or U20364 (N_20364,N_19566,N_13045);
nor U20365 (N_20365,N_18953,N_18987);
or U20366 (N_20366,N_18879,N_16442);
nor U20367 (N_20367,N_18922,N_18070);
or U20368 (N_20368,N_18954,N_17049);
nor U20369 (N_20369,N_19702,N_13244);
nand U20370 (N_20370,N_15685,N_13838);
nand U20371 (N_20371,N_17717,N_11630);
nand U20372 (N_20372,N_13768,N_15693);
nor U20373 (N_20373,N_15119,N_12359);
nor U20374 (N_20374,N_14214,N_15657);
nand U20375 (N_20375,N_10542,N_19904);
or U20376 (N_20376,N_18140,N_15413);
xnor U20377 (N_20377,N_15759,N_16225);
nand U20378 (N_20378,N_13618,N_16588);
or U20379 (N_20379,N_10551,N_17063);
nor U20380 (N_20380,N_11280,N_18677);
nor U20381 (N_20381,N_11522,N_14963);
nor U20382 (N_20382,N_10392,N_14319);
xnor U20383 (N_20383,N_10686,N_18277);
nor U20384 (N_20384,N_17844,N_15450);
xor U20385 (N_20385,N_19295,N_11193);
nand U20386 (N_20386,N_11654,N_16132);
nor U20387 (N_20387,N_14682,N_14469);
xor U20388 (N_20388,N_14649,N_16106);
and U20389 (N_20389,N_12541,N_19092);
nor U20390 (N_20390,N_12290,N_14127);
xor U20391 (N_20391,N_10669,N_15732);
nand U20392 (N_20392,N_12671,N_18559);
or U20393 (N_20393,N_18835,N_12297);
and U20394 (N_20394,N_12329,N_11825);
and U20395 (N_20395,N_15184,N_17676);
xnor U20396 (N_20396,N_17214,N_10450);
or U20397 (N_20397,N_16583,N_14883);
or U20398 (N_20398,N_19051,N_11484);
and U20399 (N_20399,N_11356,N_13246);
nor U20400 (N_20400,N_16042,N_11870);
and U20401 (N_20401,N_13534,N_17633);
or U20402 (N_20402,N_18417,N_11926);
nand U20403 (N_20403,N_17947,N_11190);
xnor U20404 (N_20404,N_19912,N_15725);
nand U20405 (N_20405,N_13709,N_11982);
nand U20406 (N_20406,N_13189,N_18436);
and U20407 (N_20407,N_13913,N_19484);
or U20408 (N_20408,N_19545,N_11625);
xor U20409 (N_20409,N_10561,N_17708);
nand U20410 (N_20410,N_14488,N_16486);
xor U20411 (N_20411,N_11303,N_19456);
nand U20412 (N_20412,N_18968,N_16034);
nor U20413 (N_20413,N_18874,N_11582);
xnor U20414 (N_20414,N_16388,N_13049);
and U20415 (N_20415,N_11740,N_10828);
or U20416 (N_20416,N_18458,N_11056);
or U20417 (N_20417,N_11814,N_13822);
xnor U20418 (N_20418,N_19350,N_10279);
xnor U20419 (N_20419,N_16807,N_10028);
or U20420 (N_20420,N_14343,N_13072);
nand U20421 (N_20421,N_10199,N_10492);
nor U20422 (N_20422,N_17040,N_14090);
xor U20423 (N_20423,N_14174,N_13911);
and U20424 (N_20424,N_13725,N_17787);
or U20425 (N_20425,N_18242,N_17497);
or U20426 (N_20426,N_11416,N_19507);
or U20427 (N_20427,N_13856,N_12838);
and U20428 (N_20428,N_12444,N_11851);
nor U20429 (N_20429,N_15461,N_16626);
and U20430 (N_20430,N_19337,N_19107);
or U20431 (N_20431,N_10755,N_18731);
and U20432 (N_20432,N_15314,N_12403);
xnor U20433 (N_20433,N_19111,N_14336);
xor U20434 (N_20434,N_11633,N_10426);
xor U20435 (N_20435,N_10697,N_10137);
nor U20436 (N_20436,N_19116,N_11863);
and U20437 (N_20437,N_17791,N_19558);
or U20438 (N_20438,N_18278,N_10484);
or U20439 (N_20439,N_16148,N_12048);
xor U20440 (N_20440,N_16845,N_19633);
or U20441 (N_20441,N_14089,N_13875);
and U20442 (N_20442,N_11922,N_13195);
nor U20443 (N_20443,N_10301,N_18659);
xnor U20444 (N_20444,N_16682,N_19605);
or U20445 (N_20445,N_19953,N_18634);
nand U20446 (N_20446,N_14288,N_10231);
or U20447 (N_20447,N_10373,N_19823);
nand U20448 (N_20448,N_10479,N_15074);
and U20449 (N_20449,N_17184,N_17386);
and U20450 (N_20450,N_19460,N_10297);
nand U20451 (N_20451,N_17711,N_14599);
and U20452 (N_20452,N_12118,N_14681);
nand U20453 (N_20453,N_18385,N_14430);
nor U20454 (N_20454,N_14949,N_16324);
nand U20455 (N_20455,N_17731,N_14860);
nand U20456 (N_20456,N_18026,N_13001);
and U20457 (N_20457,N_15563,N_18883);
and U20458 (N_20458,N_19604,N_12326);
or U20459 (N_20459,N_19155,N_17601);
nand U20460 (N_20460,N_13847,N_14923);
xnor U20461 (N_20461,N_18780,N_15212);
nor U20462 (N_20462,N_17900,N_11132);
nor U20463 (N_20463,N_15400,N_14879);
or U20464 (N_20464,N_16787,N_13297);
nor U20465 (N_20465,N_19578,N_10643);
xor U20466 (N_20466,N_15582,N_13459);
or U20467 (N_20467,N_16386,N_10182);
and U20468 (N_20468,N_12621,N_12227);
nor U20469 (N_20469,N_15522,N_13089);
nand U20470 (N_20470,N_16721,N_10247);
or U20471 (N_20471,N_19529,N_12007);
xnor U20472 (N_20472,N_15957,N_14457);
xnor U20473 (N_20473,N_10194,N_12792);
nand U20474 (N_20474,N_18983,N_12693);
xnor U20475 (N_20475,N_18950,N_16783);
and U20476 (N_20476,N_11309,N_11238);
nand U20477 (N_20477,N_13967,N_14570);
nand U20478 (N_20478,N_12695,N_11896);
and U20479 (N_20479,N_13403,N_18802);
or U20480 (N_20480,N_15057,N_15677);
or U20481 (N_20481,N_14030,N_17116);
nor U20482 (N_20482,N_14596,N_15879);
nand U20483 (N_20483,N_13774,N_14021);
nor U20484 (N_20484,N_12742,N_17180);
nand U20485 (N_20485,N_19657,N_12050);
and U20486 (N_20486,N_13938,N_17690);
or U20487 (N_20487,N_18059,N_14973);
nor U20488 (N_20488,N_16739,N_13500);
nand U20489 (N_20489,N_16226,N_13145);
and U20490 (N_20490,N_11886,N_14434);
and U20491 (N_20491,N_19935,N_12120);
nor U20492 (N_20492,N_13576,N_11085);
nor U20493 (N_20493,N_11234,N_14123);
xnor U20494 (N_20494,N_10480,N_16975);
xor U20495 (N_20495,N_11579,N_14067);
nand U20496 (N_20496,N_16556,N_18259);
nand U20497 (N_20497,N_16980,N_12773);
nand U20498 (N_20498,N_13062,N_15375);
xor U20499 (N_20499,N_18757,N_16723);
and U20500 (N_20500,N_16024,N_13066);
or U20501 (N_20501,N_14375,N_11242);
nor U20502 (N_20502,N_14566,N_14903);
and U20503 (N_20503,N_14622,N_11314);
nor U20504 (N_20504,N_17119,N_17907);
xor U20505 (N_20505,N_11246,N_13133);
nor U20506 (N_20506,N_12800,N_19293);
and U20507 (N_20507,N_12371,N_10872);
nor U20508 (N_20508,N_11599,N_16498);
nor U20509 (N_20509,N_17761,N_15626);
nand U20510 (N_20510,N_16976,N_19165);
or U20511 (N_20511,N_10121,N_19095);
nand U20512 (N_20512,N_10602,N_19127);
xor U20513 (N_20513,N_19983,N_17894);
nor U20514 (N_20514,N_16418,N_17034);
or U20515 (N_20515,N_13465,N_12235);
xnor U20516 (N_20516,N_18826,N_10041);
and U20517 (N_20517,N_16429,N_11366);
and U20518 (N_20518,N_17805,N_13790);
and U20519 (N_20519,N_17343,N_18925);
xnor U20520 (N_20520,N_11622,N_13442);
nand U20521 (N_20521,N_14112,N_12114);
nand U20522 (N_20522,N_13312,N_13424);
nand U20523 (N_20523,N_13003,N_18625);
xnor U20524 (N_20524,N_14043,N_19928);
and U20525 (N_20525,N_15084,N_10577);
nor U20526 (N_20526,N_10283,N_15766);
or U20527 (N_20527,N_17970,N_13695);
and U20528 (N_20528,N_16584,N_12386);
nand U20529 (N_20529,N_11629,N_14421);
xor U20530 (N_20530,N_11175,N_12954);
nand U20531 (N_20531,N_15546,N_11265);
or U20532 (N_20532,N_19589,N_12886);
or U20533 (N_20533,N_13158,N_13096);
nor U20534 (N_20534,N_11382,N_14521);
and U20535 (N_20535,N_16953,N_13397);
and U20536 (N_20536,N_14954,N_16371);
xor U20537 (N_20537,N_19226,N_14722);
xnor U20538 (N_20538,N_17236,N_15460);
nor U20539 (N_20539,N_17890,N_11299);
xor U20540 (N_20540,N_10761,N_12941);
or U20541 (N_20541,N_12826,N_11724);
or U20542 (N_20542,N_17867,N_18577);
nand U20543 (N_20543,N_12746,N_10749);
and U20544 (N_20544,N_13812,N_15904);
xor U20545 (N_20545,N_18605,N_10820);
nor U20546 (N_20546,N_19058,N_10519);
nor U20547 (N_20547,N_10214,N_13120);
or U20548 (N_20548,N_13041,N_16428);
nand U20549 (N_20549,N_10238,N_17394);
nand U20550 (N_20550,N_14223,N_12083);
and U20551 (N_20551,N_17495,N_11789);
nor U20552 (N_20552,N_15394,N_15286);
nand U20553 (N_20553,N_17931,N_18291);
or U20554 (N_20554,N_19725,N_15977);
xor U20555 (N_20555,N_15008,N_15308);
or U20556 (N_20556,N_18633,N_12228);
nor U20557 (N_20557,N_19538,N_10106);
nand U20558 (N_20558,N_15750,N_12953);
xor U20559 (N_20559,N_11022,N_14947);
xnor U20560 (N_20560,N_19273,N_11727);
xnor U20561 (N_20561,N_16048,N_10225);
nor U20562 (N_20562,N_19185,N_18976);
and U20563 (N_20563,N_13167,N_16135);
nand U20564 (N_20564,N_11224,N_17839);
xnor U20565 (N_20565,N_15967,N_15839);
xor U20566 (N_20566,N_16112,N_19731);
or U20567 (N_20567,N_19428,N_12806);
nor U20568 (N_20568,N_11997,N_12883);
or U20569 (N_20569,N_14134,N_16781);
xor U20570 (N_20570,N_14314,N_13203);
and U20571 (N_20571,N_15950,N_19550);
or U20572 (N_20572,N_14002,N_12913);
nor U20573 (N_20573,N_15698,N_17131);
or U20574 (N_20574,N_19880,N_10436);
nand U20575 (N_20575,N_14027,N_14504);
xnor U20576 (N_20576,N_12040,N_10171);
xor U20577 (N_20577,N_14378,N_17143);
or U20578 (N_20578,N_19343,N_13575);
and U20579 (N_20579,N_13979,N_12833);
and U20580 (N_20580,N_16194,N_15757);
xor U20581 (N_20581,N_19422,N_15621);
nor U20582 (N_20582,N_10652,N_17764);
nand U20583 (N_20583,N_15686,N_16534);
xnor U20584 (N_20584,N_19313,N_16063);
and U20585 (N_20585,N_14833,N_12472);
nand U20586 (N_20586,N_12304,N_12821);
xor U20587 (N_20587,N_15246,N_14609);
or U20588 (N_20588,N_15820,N_14731);
or U20589 (N_20589,N_11790,N_11942);
or U20590 (N_20590,N_10539,N_17280);
nand U20591 (N_20591,N_14586,N_14346);
nand U20592 (N_20592,N_12015,N_16599);
and U20593 (N_20593,N_15791,N_14646);
nor U20594 (N_20594,N_18416,N_13881);
nand U20595 (N_20595,N_19892,N_16483);
and U20596 (N_20596,N_11052,N_12680);
nand U20597 (N_20597,N_18850,N_18018);
or U20598 (N_20598,N_15948,N_14689);
nand U20599 (N_20599,N_19136,N_14320);
or U20600 (N_20600,N_10886,N_15242);
or U20601 (N_20601,N_18039,N_15016);
and U20602 (N_20602,N_17152,N_19793);
or U20603 (N_20603,N_13517,N_17538);
xnor U20604 (N_20604,N_17614,N_11146);
nand U20605 (N_20605,N_16959,N_16873);
and U20606 (N_20606,N_19213,N_19598);
nor U20607 (N_20607,N_10289,N_11548);
nor U20608 (N_20608,N_10531,N_14076);
nand U20609 (N_20609,N_19993,N_16270);
and U20610 (N_20610,N_18475,N_19901);
xor U20611 (N_20611,N_15381,N_14166);
nand U20612 (N_20612,N_17906,N_14992);
nand U20613 (N_20613,N_10513,N_19252);
xnor U20614 (N_20614,N_13520,N_17387);
nor U20615 (N_20615,N_11542,N_10617);
nand U20616 (N_20616,N_16852,N_17759);
and U20617 (N_20617,N_15093,N_16185);
and U20618 (N_20618,N_13491,N_17025);
xor U20619 (N_20619,N_15448,N_18779);
or U20620 (N_20620,N_11614,N_12889);
nand U20621 (N_20621,N_18548,N_14766);
nor U20622 (N_20622,N_19697,N_14745);
nand U20623 (N_20623,N_10646,N_14936);
and U20624 (N_20624,N_15361,N_19099);
and U20625 (N_20625,N_10300,N_15480);
or U20626 (N_20626,N_10466,N_16196);
nor U20627 (N_20627,N_13091,N_16698);
nand U20628 (N_20628,N_15736,N_10511);
nor U20629 (N_20629,N_14489,N_17468);
and U20630 (N_20630,N_11586,N_13352);
or U20631 (N_20631,N_19365,N_13843);
or U20632 (N_20632,N_11192,N_15537);
nor U20633 (N_20633,N_13863,N_19461);
nor U20634 (N_20634,N_10567,N_12241);
xor U20635 (N_20635,N_11254,N_16844);
nand U20636 (N_20636,N_17579,N_18109);
and U20637 (N_20637,N_10839,N_15065);
and U20638 (N_20638,N_10022,N_13226);
and U20639 (N_20639,N_11766,N_17898);
nor U20640 (N_20640,N_12959,N_14685);
xor U20641 (N_20641,N_19025,N_18216);
or U20642 (N_20642,N_16999,N_17607);
or U20643 (N_20643,N_16860,N_16843);
xor U20644 (N_20644,N_16111,N_12745);
xor U20645 (N_20645,N_13260,N_18860);
or U20646 (N_20646,N_19268,N_18079);
or U20647 (N_20647,N_10391,N_15555);
nand U20648 (N_20648,N_15344,N_13006);
or U20649 (N_20649,N_12866,N_10662);
or U20650 (N_20650,N_16870,N_11691);
xnor U20651 (N_20651,N_18226,N_11114);
or U20652 (N_20652,N_18167,N_11543);
nor U20653 (N_20653,N_15185,N_10433);
and U20654 (N_20654,N_18839,N_11726);
nor U20655 (N_20655,N_18927,N_11744);
nand U20656 (N_20656,N_15739,N_10204);
or U20657 (N_20657,N_17589,N_19018);
nand U20658 (N_20658,N_16469,N_12069);
nor U20659 (N_20659,N_18345,N_17810);
xnor U20660 (N_20660,N_17254,N_11803);
nand U20661 (N_20661,N_12981,N_11332);
or U20662 (N_20662,N_19354,N_14492);
xnor U20663 (N_20663,N_11717,N_17905);
nand U20664 (N_20664,N_11898,N_10259);
and U20665 (N_20665,N_15605,N_10550);
nor U20666 (N_20666,N_18297,N_17273);
xnor U20667 (N_20667,N_17985,N_12471);
nand U20668 (N_20668,N_14210,N_18229);
or U20669 (N_20669,N_14914,N_10060);
or U20670 (N_20670,N_13275,N_12181);
nor U20671 (N_20671,N_16076,N_18536);
xor U20672 (N_20672,N_17576,N_14891);
and U20673 (N_20673,N_12521,N_16875);
xor U20674 (N_20674,N_19767,N_14590);
nand U20675 (N_20675,N_19539,N_16772);
and U20676 (N_20676,N_17834,N_13222);
or U20677 (N_20677,N_10439,N_18616);
and U20678 (N_20678,N_13645,N_13883);
and U20679 (N_20679,N_11911,N_17946);
nand U20680 (N_20680,N_10654,N_16744);
nor U20681 (N_20681,N_15597,N_12375);
and U20682 (N_20682,N_15403,N_16167);
nand U20683 (N_20683,N_12442,N_11594);
nand U20684 (N_20684,N_18053,N_17431);
xor U20685 (N_20685,N_14876,N_12497);
or U20686 (N_20686,N_10340,N_16956);
nor U20687 (N_20687,N_17685,N_14287);
or U20688 (N_20688,N_17692,N_10104);
xnor U20689 (N_20689,N_18897,N_10879);
nor U20690 (N_20690,N_11709,N_10299);
or U20691 (N_20691,N_15944,N_10585);
or U20692 (N_20692,N_14484,N_18234);
and U20693 (N_20693,N_13761,N_12432);
or U20694 (N_20694,N_13836,N_14755);
and U20695 (N_20695,N_19929,N_14717);
nor U20696 (N_20696,N_10263,N_11443);
nor U20697 (N_20697,N_14322,N_10483);
nor U20698 (N_20698,N_10722,N_10810);
xnor U20699 (N_20699,N_18206,N_12426);
and U20700 (N_20700,N_13131,N_17189);
and U20701 (N_20701,N_14713,N_10943);
and U20702 (N_20702,N_16335,N_11236);
and U20703 (N_20703,N_10374,N_17582);
or U20704 (N_20704,N_19229,N_14694);
nand U20705 (N_20705,N_15201,N_14432);
nand U20706 (N_20706,N_11688,N_18202);
nor U20707 (N_20707,N_16674,N_15644);
or U20708 (N_20708,N_12236,N_11974);
nand U20709 (N_20709,N_17113,N_17927);
nand U20710 (N_20710,N_11747,N_10728);
or U20711 (N_20711,N_11506,N_17136);
nor U20712 (N_20712,N_16021,N_12553);
nand U20713 (N_20713,N_13837,N_12421);
and U20714 (N_20714,N_12567,N_17266);
nand U20715 (N_20715,N_17334,N_18710);
nand U20716 (N_20716,N_11472,N_17829);
or U20717 (N_20717,N_14498,N_15063);
xor U20718 (N_20718,N_17491,N_19831);
xor U20719 (N_20719,N_13245,N_15158);
nand U20720 (N_20720,N_12601,N_19885);
and U20721 (N_20721,N_19299,N_12480);
xnor U20722 (N_20722,N_11039,N_14479);
and U20723 (N_20723,N_11587,N_12798);
nor U20724 (N_20724,N_16089,N_12920);
nor U20725 (N_20725,N_13088,N_18177);
nor U20726 (N_20726,N_19342,N_15260);
and U20727 (N_20727,N_16913,N_16729);
or U20728 (N_20728,N_13284,N_16302);
or U20729 (N_20729,N_12003,N_12025);
nor U20730 (N_20730,N_12406,N_14996);
or U20731 (N_20731,N_14377,N_19120);
xnor U20732 (N_20732,N_16768,N_12429);
and U20733 (N_20733,N_15130,N_15029);
nor U20734 (N_20734,N_16045,N_16079);
nor U20735 (N_20735,N_16118,N_11978);
nand U20736 (N_20736,N_17219,N_13385);
nand U20737 (N_20737,N_18318,N_19951);
xor U20738 (N_20738,N_11824,N_11769);
and U20739 (N_20739,N_16177,N_12845);
xor U20740 (N_20740,N_12882,N_18808);
and U20741 (N_20741,N_16306,N_12708);
and U20742 (N_20742,N_12334,N_11079);
xnor U20743 (N_20743,N_19711,N_13679);
and U20744 (N_20744,N_11200,N_18124);
and U20745 (N_20745,N_10187,N_17134);
nand U20746 (N_20746,N_13887,N_18134);
and U20747 (N_20747,N_13113,N_18365);
nor U20748 (N_20748,N_14045,N_14643);
xor U20749 (N_20749,N_18560,N_18878);
nor U20750 (N_20750,N_18063,N_17372);
xnor U20751 (N_20751,N_17929,N_10673);
nand U20752 (N_20752,N_13729,N_19455);
xor U20753 (N_20753,N_17109,N_10951);
xor U20754 (N_20754,N_12644,N_17373);
nand U20755 (N_20755,N_12606,N_14159);
nor U20756 (N_20756,N_13194,N_19085);
or U20757 (N_20757,N_19480,N_17952);
nor U20758 (N_20758,N_19934,N_18042);
xor U20759 (N_20759,N_16246,N_10827);
and U20760 (N_20760,N_11440,N_15406);
xnor U20761 (N_20761,N_18485,N_14553);
and U20762 (N_20762,N_13231,N_14556);
nor U20763 (N_20763,N_18393,N_17313);
xor U20764 (N_20764,N_16792,N_15465);
or U20765 (N_20765,N_11804,N_18270);
xor U20766 (N_20766,N_15680,N_19317);
nand U20767 (N_20767,N_16964,N_11464);
nand U20768 (N_20768,N_18303,N_16039);
and U20769 (N_20769,N_10149,N_10915);
xnor U20770 (N_20770,N_14096,N_14933);
or U20771 (N_20771,N_13213,N_11491);
and U20772 (N_20772,N_17087,N_14765);
nor U20773 (N_20773,N_10339,N_18127);
nand U20774 (N_20774,N_15263,N_10142);
and U20775 (N_20775,N_16221,N_17145);
xor U20776 (N_20776,N_16876,N_17996);
nor U20777 (N_20777,N_13543,N_15227);
nor U20778 (N_20778,N_19867,N_18971);
or U20779 (N_20779,N_17969,N_11983);
nand U20780 (N_20780,N_16453,N_11258);
nand U20781 (N_20781,N_11276,N_12214);
and U20782 (N_20782,N_16950,N_10456);
nor U20783 (N_20783,N_11796,N_15482);
nor U20784 (N_20784,N_12184,N_19069);
nand U20785 (N_20785,N_13035,N_12554);
nand U20786 (N_20786,N_13560,N_18642);
xor U20787 (N_20787,N_16510,N_12542);
and U20788 (N_20788,N_10753,N_17757);
xnor U20789 (N_20789,N_12723,N_18174);
nand U20790 (N_20790,N_11167,N_12877);
and U20791 (N_20791,N_13080,N_14991);
nand U20792 (N_20792,N_14307,N_19703);
or U20793 (N_20793,N_16840,N_18187);
nand U20794 (N_20794,N_16675,N_15366);
nor U20795 (N_20795,N_10193,N_19569);
nand U20796 (N_20796,N_17465,N_17315);
or U20797 (N_20797,N_16696,N_14900);
or U20798 (N_20798,N_17926,N_18873);
xnor U20799 (N_20799,N_16097,N_17634);
and U20800 (N_20800,N_15025,N_13590);
or U20801 (N_20801,N_10170,N_17205);
nor U20802 (N_20802,N_11271,N_10495);
nand U20803 (N_20803,N_13274,N_19491);
xor U20804 (N_20804,N_14211,N_10179);
and U20805 (N_20805,N_15002,N_15625);
nor U20806 (N_20806,N_19642,N_19521);
nor U20807 (N_20807,N_11713,N_15472);
nor U20808 (N_20808,N_14932,N_15981);
nor U20809 (N_20809,N_19301,N_17865);
nand U20810 (N_20810,N_11142,N_19636);
nand U20811 (N_20811,N_13048,N_10073);
nand U20812 (N_20812,N_18369,N_13261);
nor U20813 (N_20813,N_12580,N_14750);
nand U20814 (N_20814,N_14190,N_13249);
nor U20815 (N_20815,N_17295,N_12775);
and U20816 (N_20816,N_15171,N_12138);
or U20817 (N_20817,N_19159,N_16234);
and U20818 (N_20818,N_13706,N_13777);
or U20819 (N_20819,N_14273,N_10064);
or U20820 (N_20820,N_14928,N_17308);
nor U20821 (N_20821,N_17489,N_14109);
nor U20822 (N_20822,N_19052,N_15027);
xor U20823 (N_20823,N_14835,N_13097);
xnor U20824 (N_20824,N_16692,N_13116);
and U20825 (N_20825,N_11301,N_18495);
or U20826 (N_20826,N_18590,N_12173);
nor U20827 (N_20827,N_12230,N_16312);
xor U20828 (N_20828,N_17556,N_15864);
nand U20829 (N_20829,N_13202,N_13666);
nor U20830 (N_20830,N_12549,N_14440);
xor U20831 (N_20831,N_17285,N_17941);
nor U20832 (N_20832,N_19608,N_16047);
and U20833 (N_20833,N_10437,N_17366);
nand U20834 (N_20834,N_13928,N_15607);
xor U20835 (N_20835,N_17569,N_10707);
xor U20836 (N_20836,N_18220,N_17377);
and U20837 (N_20837,N_13399,N_12597);
and U20838 (N_20838,N_17797,N_12844);
and U20839 (N_20839,N_10284,N_14386);
nand U20840 (N_20840,N_19297,N_18939);
nand U20841 (N_20841,N_18477,N_14321);
nand U20842 (N_20842,N_18723,N_14253);
xnor U20843 (N_20843,N_18744,N_12797);
or U20844 (N_20844,N_18982,N_12231);
or U20845 (N_20845,N_13616,N_10449);
nor U20846 (N_20846,N_14160,N_14419);
nor U20847 (N_20847,N_10010,N_16181);
or U20848 (N_20848,N_14505,N_12027);
nand U20849 (N_20849,N_17311,N_13658);
and U20850 (N_20850,N_18276,N_15653);
or U20851 (N_20851,N_16374,N_10593);
xor U20852 (N_20852,N_17725,N_19695);
xnor U20853 (N_20853,N_13034,N_19199);
nand U20854 (N_20854,N_18882,N_16836);
or U20855 (N_20855,N_12056,N_17978);
xor U20856 (N_20856,N_14804,N_16172);
and U20857 (N_20857,N_13778,N_10795);
nand U20858 (N_20858,N_12818,N_19875);
xor U20859 (N_20859,N_12001,N_15208);
and U20860 (N_20860,N_19351,N_13247);
xnor U20861 (N_20861,N_16188,N_19145);
and U20862 (N_20862,N_19870,N_15066);
xnor U20863 (N_20863,N_17547,N_11598);
nor U20864 (N_20864,N_17045,N_16023);
or U20865 (N_20865,N_17564,N_15305);
and U20866 (N_20866,N_12724,N_15747);
or U20867 (N_20867,N_15360,N_18479);
nor U20868 (N_20868,N_16735,N_16345);
or U20869 (N_20869,N_17151,N_14708);
nand U20870 (N_20870,N_16279,N_18010);
and U20871 (N_20871,N_10877,N_10315);
nor U20872 (N_20872,N_17075,N_16314);
xnor U20873 (N_20873,N_10160,N_19181);
nand U20874 (N_20874,N_18531,N_13467);
nor U20875 (N_20875,N_19385,N_11973);
xor U20876 (N_20876,N_16075,N_12408);
and U20877 (N_20877,N_11918,N_13455);
nand U20878 (N_20878,N_17526,N_10568);
nor U20879 (N_20879,N_15996,N_10847);
nor U20880 (N_20880,N_17210,N_15306);
xnor U20881 (N_20881,N_12832,N_15101);
nand U20882 (N_20882,N_13441,N_13830);
or U20883 (N_20883,N_10823,N_14459);
xor U20884 (N_20884,N_18911,N_13958);
xnor U20885 (N_20885,N_17332,N_13216);
nand U20886 (N_20886,N_18656,N_18526);
xor U20887 (N_20887,N_18146,N_18773);
nor U20888 (N_20888,N_15570,N_16987);
or U20889 (N_20889,N_12452,N_15319);
nor U20890 (N_20890,N_16651,N_14380);
nand U20891 (N_20891,N_15298,N_19856);
nand U20892 (N_20892,N_10131,N_10504);
xnor U20893 (N_20893,N_17629,N_16869);
nand U20894 (N_20894,N_14341,N_17792);
or U20895 (N_20895,N_11036,N_14759);
nand U20896 (N_20896,N_19390,N_16137);
and U20897 (N_20897,N_15568,N_17462);
or U20898 (N_20898,N_15953,N_19651);
nor U20899 (N_20899,N_11893,N_17486);
or U20900 (N_20900,N_17403,N_14442);
or U20901 (N_20901,N_17675,N_15155);
and U20902 (N_20902,N_11674,N_14237);
nand U20903 (N_20903,N_18827,N_12762);
or U20904 (N_20904,N_13209,N_10731);
nand U20905 (N_20905,N_15692,N_18342);
nor U20906 (N_20906,N_18843,N_18348);
nor U20907 (N_20907,N_14503,N_13693);
and U20908 (N_20908,N_13596,N_14817);
or U20909 (N_20909,N_16711,N_14470);
nor U20910 (N_20910,N_11887,N_14957);
nand U20911 (N_20911,N_12820,N_11351);
xnor U20912 (N_20912,N_19773,N_14931);
xor U20913 (N_20913,N_18024,N_19258);
nor U20914 (N_20914,N_15588,N_18742);
xor U20915 (N_20915,N_10607,N_17762);
nor U20916 (N_20916,N_17191,N_14594);
and U20917 (N_20917,N_15267,N_19883);
nor U20918 (N_20918,N_10831,N_11149);
xor U20919 (N_20919,N_18314,N_14615);
xor U20920 (N_20920,N_12090,N_15921);
and U20921 (N_20921,N_19124,N_16549);
xnor U20922 (N_20922,N_11304,N_13718);
and U20923 (N_20923,N_17930,N_10764);
and U20924 (N_20924,N_14551,N_10575);
or U20925 (N_20925,N_13129,N_19812);
nor U20926 (N_20926,N_14020,N_17750);
and U20927 (N_20927,N_12242,N_19004);
and U20928 (N_20928,N_10515,N_17790);
xnor U20929 (N_20929,N_15205,N_12764);
xnor U20930 (N_20930,N_11610,N_19048);
or U20931 (N_20931,N_17159,N_19790);
nand U20932 (N_20932,N_11235,N_16414);
or U20933 (N_20933,N_16805,N_18316);
or U20934 (N_20934,N_16091,N_13174);
nor U20935 (N_20935,N_12410,N_16275);
nor U20936 (N_20936,N_17741,N_18478);
and U20937 (N_20937,N_10955,N_18162);
or U20938 (N_20938,N_19858,N_19783);
or U20939 (N_20939,N_18011,N_17683);
xnor U20940 (N_20940,N_15176,N_11287);
xor U20941 (N_20941,N_14848,N_14740);
and U20942 (N_20942,N_17565,N_15869);
xnor U20943 (N_20943,N_12560,N_19068);
or U20944 (N_20944,N_14347,N_10412);
nand U20945 (N_20945,N_17115,N_13325);
nor U20946 (N_20946,N_11527,N_10703);
or U20947 (N_20947,N_11651,N_16733);
and U20948 (N_20948,N_16949,N_11780);
or U20949 (N_20949,N_11071,N_11116);
or U20950 (N_20950,N_16685,N_15830);
nand U20951 (N_20951,N_16271,N_14888);
nand U20952 (N_20952,N_19862,N_12650);
nand U20953 (N_20953,N_18857,N_15111);
xor U20954 (N_20954,N_18349,N_10465);
nor U20955 (N_20955,N_12370,N_10661);
or U20956 (N_20956,N_15021,N_15980);
and U20957 (N_20957,N_14005,N_12466);
and U20958 (N_20958,N_16839,N_16424);
nand U20959 (N_20959,N_15156,N_15415);
nor U20960 (N_20960,N_19401,N_18803);
xor U20961 (N_20961,N_10959,N_13671);
nand U20962 (N_20962,N_13732,N_16041);
or U20963 (N_20963,N_17092,N_15104);
or U20964 (N_20964,N_16057,N_10404);
nor U20965 (N_20965,N_17560,N_19863);
nand U20966 (N_20966,N_13558,N_19525);
or U20967 (N_20967,N_18561,N_18628);
or U20968 (N_20968,N_15956,N_11871);
nand U20969 (N_20969,N_17391,N_10861);
xor U20970 (N_20970,N_16657,N_14499);
and U20971 (N_20971,N_17613,N_15919);
xor U20972 (N_20972,N_12583,N_18597);
nor U20973 (N_20973,N_10705,N_10573);
nand U20974 (N_20974,N_11044,N_10798);
nand U20975 (N_20975,N_19118,N_17847);
and U20976 (N_20976,N_17866,N_16594);
nor U20977 (N_20977,N_12322,N_17779);
xnor U20978 (N_20978,N_11697,N_12291);
nand U20979 (N_20979,N_14664,N_11445);
nand U20980 (N_20980,N_12266,N_12836);
nand U20981 (N_20981,N_13612,N_10777);
nand U20982 (N_20982,N_13406,N_14009);
nand U20983 (N_20983,N_10027,N_17073);
nand U20984 (N_20984,N_15230,N_16816);
and U20985 (N_20985,N_19501,N_15684);
nor U20986 (N_20986,N_10571,N_10304);
nor U20987 (N_20987,N_11554,N_11868);
or U20988 (N_20988,N_11693,N_18761);
or U20989 (N_20989,N_12205,N_16937);
or U20990 (N_20990,N_11355,N_11538);
nand U20991 (N_20991,N_12760,N_18335);
nor U20992 (N_20992,N_11524,N_14256);
and U20993 (N_20993,N_17971,N_19505);
nor U20994 (N_20994,N_12757,N_16003);
xnor U20995 (N_20995,N_17514,N_14535);
nand U20996 (N_20996,N_19614,N_12358);
xor U20997 (N_20997,N_19606,N_12632);
and U20998 (N_20998,N_10272,N_10969);
nor U20999 (N_20999,N_19376,N_18302);
or U21000 (N_21000,N_15240,N_14899);
nor U21001 (N_21001,N_18425,N_12917);
or U21002 (N_21002,N_15675,N_15473);
xnor U21003 (N_21003,N_15601,N_19522);
or U21004 (N_21004,N_19367,N_19173);
nand U21005 (N_21005,N_12540,N_18734);
and U21006 (N_21006,N_15531,N_15131);
or U21007 (N_21007,N_16452,N_13722);
nor U21008 (N_21008,N_14150,N_17706);
nor U21009 (N_21009,N_19849,N_10663);
nand U21010 (N_21010,N_12880,N_15872);
or U21011 (N_21011,N_18977,N_12692);
or U21012 (N_21012,N_15197,N_10569);
and U21013 (N_21013,N_15730,N_18336);
xnor U21014 (N_21014,N_17142,N_16596);
or U21015 (N_21015,N_18106,N_11247);
nor U21016 (N_21016,N_13372,N_12571);
xnor U21017 (N_21017,N_17818,N_15850);
and U21018 (N_21018,N_11914,N_13437);
nor U21019 (N_21019,N_17840,N_12937);
nand U21020 (N_21020,N_16008,N_12850);
or U21021 (N_21021,N_10889,N_12612);
nor U21022 (N_21022,N_17022,N_13619);
nand U21023 (N_21023,N_12407,N_11339);
nor U21024 (N_21024,N_19132,N_18131);
nor U21025 (N_21025,N_19580,N_12629);
and U21026 (N_21026,N_18884,N_17798);
or U21027 (N_21027,N_14558,N_15525);
nand U21028 (N_21028,N_16404,N_19634);
xnor U21029 (N_21029,N_13054,N_19265);
xnor U21030 (N_21030,N_19217,N_13524);
and U21031 (N_21031,N_15648,N_12870);
and U21032 (N_21032,N_18194,N_14626);
and U21033 (N_21033,N_11830,N_17442);
and U21034 (N_21034,N_14168,N_18876);
nand U21035 (N_21035,N_10408,N_13980);
xnor U21036 (N_21036,N_15115,N_14075);
or U21037 (N_21037,N_16009,N_18846);
nand U21038 (N_21038,N_19768,N_14733);
or U21039 (N_21039,N_10748,N_16533);
xor U21040 (N_21040,N_10267,N_11298);
nand U21041 (N_21041,N_14534,N_10885);
or U21042 (N_21042,N_16459,N_17069);
xor U21043 (N_21043,N_18836,N_12598);
and U21044 (N_21044,N_13719,N_16589);
nand U21045 (N_21045,N_12361,N_15590);
nand U21046 (N_21046,N_13737,N_17988);
and U21047 (N_21047,N_13353,N_10888);
or U21048 (N_21048,N_18418,N_15302);
nand U21049 (N_21049,N_14428,N_14406);
nor U21050 (N_21050,N_19602,N_16896);
and U21051 (N_21051,N_15720,N_12839);
nand U21052 (N_21052,N_13850,N_12400);
nand U21053 (N_21053,N_18823,N_19871);
and U21054 (N_21054,N_14793,N_14588);
or U21055 (N_21055,N_13343,N_11683);
nand U21056 (N_21056,N_18308,N_18441);
or U21057 (N_21057,N_18973,N_11029);
nor U21058 (N_21058,N_18908,N_16109);
and U21059 (N_21059,N_14508,N_13886);
xor U21060 (N_21060,N_16206,N_17747);
nor U21061 (N_21061,N_16187,N_15405);
xor U21062 (N_21062,N_15338,N_18864);
xnor U21063 (N_21063,N_10580,N_16202);
nand U21064 (N_21064,N_11214,N_15277);
or U21065 (N_21065,N_10059,N_18711);
xor U21066 (N_21066,N_11779,N_14436);
xnor U21067 (N_21067,N_14351,N_16258);
nand U21068 (N_21068,N_14033,N_10342);
xor U21069 (N_21069,N_18816,N_12987);
nand U21070 (N_21070,N_15528,N_15177);
nand U21071 (N_21071,N_11067,N_11007);
nand U21072 (N_21072,N_13333,N_10687);
xnor U21073 (N_21073,N_14830,N_19809);
nand U21074 (N_21074,N_10808,N_11009);
and U21075 (N_21075,N_17235,N_14511);
nor U21076 (N_21076,N_18090,N_10031);
or U21077 (N_21077,N_12055,N_19964);
nor U21078 (N_21078,N_14283,N_12823);
and U21079 (N_21079,N_17234,N_16245);
and U21080 (N_21080,N_18459,N_12483);
and U21081 (N_21081,N_14811,N_16236);
nand U21082 (N_21082,N_12771,N_16149);
xnor U21083 (N_21083,N_19405,N_11350);
and U21084 (N_21084,N_11479,N_10174);
nand U21085 (N_21085,N_16992,N_16186);
or U21086 (N_21086,N_13933,N_19816);
nor U21087 (N_21087,N_19349,N_14064);
and U21088 (N_21088,N_15802,N_16994);
or U21089 (N_21089,N_13462,N_16338);
nand U21090 (N_21090,N_11173,N_14142);
and U21091 (N_21091,N_16738,N_14035);
nand U21092 (N_21092,N_16249,N_10909);
nand U21093 (N_21093,N_11676,N_11748);
or U21094 (N_21094,N_14819,N_19209);
xor U21095 (N_21095,N_10345,N_13298);
and U21096 (N_21096,N_12995,N_17043);
nor U21097 (N_21097,N_11721,N_17433);
nor U21098 (N_21098,N_14629,N_16262);
or U21099 (N_21099,N_18192,N_11647);
or U21100 (N_21100,N_10599,N_18161);
and U21101 (N_21101,N_11107,N_12591);
nor U21102 (N_21102,N_16794,N_13469);
nor U21103 (N_21103,N_11652,N_12903);
nand U21104 (N_21104,N_15876,N_11584);
xor U21105 (N_21105,N_10363,N_17535);
nor U21106 (N_21106,N_13180,N_14433);
and U21107 (N_21107,N_17398,N_17604);
nor U21108 (N_21108,N_16568,N_13278);
xor U21109 (N_21109,N_12215,N_12613);
nand U21110 (N_21110,N_18179,N_12656);
or U21111 (N_21111,N_11735,N_14644);
nand U21112 (N_21112,N_11869,N_14113);
nand U21113 (N_21113,N_13486,N_16051);
or U21114 (N_21114,N_14392,N_13545);
or U21115 (N_21115,N_13920,N_11597);
nand U21116 (N_21116,N_15603,N_12799);
nand U21117 (N_21117,N_12037,N_14178);
nor U21118 (N_21118,N_10424,N_17110);
nand U21119 (N_21119,N_13791,N_15299);
and U21120 (N_21120,N_11088,N_17023);
xnor U21121 (N_21121,N_18650,N_13081);
nor U21122 (N_21122,N_18073,N_16029);
nand U21123 (N_21123,N_16067,N_15054);
or U21124 (N_21124,N_11480,N_18098);
xor U21125 (N_21125,N_11189,N_12902);
or U21126 (N_21126,N_19483,N_13533);
nand U21127 (N_21127,N_10032,N_12450);
nor U21128 (N_21128,N_13417,N_10572);
xnor U21129 (N_21129,N_19551,N_12573);
and U21130 (N_21130,N_11123,N_15594);
nor U21131 (N_21131,N_11203,N_18554);
nor U21132 (N_21132,N_18358,N_10257);
or U21133 (N_21133,N_17083,N_11818);
nor U21134 (N_21134,N_14801,N_16033);
nor U21135 (N_21135,N_14205,N_19078);
or U21136 (N_21136,N_17689,N_19677);
and U21137 (N_21137,N_17309,N_19666);
nor U21138 (N_21138,N_16832,N_12223);
or U21139 (N_21139,N_12513,N_17540);
xnor U21140 (N_21140,N_19341,N_16173);
nand U21141 (N_21141,N_12763,N_18699);
nor U21142 (N_21142,N_15471,N_10931);
nor U21143 (N_21143,N_19347,N_17674);
nand U21144 (N_21144,N_15910,N_12318);
and U21145 (N_21145,N_18896,N_14369);
or U21146 (N_21146,N_14095,N_12722);
xor U21147 (N_21147,N_17482,N_18409);
xnor U21148 (N_21148,N_18566,N_13893);
nand U21149 (N_21149,N_18311,N_12191);
or U21150 (N_21150,N_13702,N_10510);
nand U21151 (N_21151,N_14062,N_11960);
nand U21152 (N_21152,N_11023,N_18929);
and U21153 (N_21153,N_19727,N_15828);
and U21154 (N_21154,N_18612,N_18776);
nor U21155 (N_21155,N_12051,N_17061);
and U21156 (N_21156,N_18568,N_14686);
nand U21157 (N_21157,N_13817,N_19227);
nor U21158 (N_21158,N_11854,N_11278);
or U21159 (N_21159,N_19091,N_10597);
xor U21160 (N_21160,N_16758,N_19648);
xnor U21161 (N_21161,N_15627,N_18214);
xnor U21162 (N_21162,N_16136,N_14604);
xnor U21163 (N_21163,N_19097,N_18795);
nor U21164 (N_21164,N_18841,N_10937);
nor U21165 (N_21165,N_18320,N_17195);
nand U21166 (N_21166,N_15812,N_15922);
xnor U21167 (N_21167,N_15081,N_14986);
and U21168 (N_21168,N_16910,N_10485);
nand U21169 (N_21169,N_15377,N_10934);
and U21170 (N_21170,N_19014,N_11537);
nor U21171 (N_21171,N_18889,N_11437);
or U21172 (N_21172,N_10053,N_17178);
nor U21173 (N_21173,N_19001,N_10029);
xor U21174 (N_21174,N_19195,N_13797);
and U21175 (N_21175,N_14907,N_10229);
nor U21176 (N_21176,N_17338,N_19176);
and U21177 (N_21177,N_16694,N_16184);
and U21178 (N_21178,N_17330,N_13978);
nor U21179 (N_21179,N_18439,N_12616);
and U21180 (N_21180,N_19251,N_16743);
xnor U21181 (N_21181,N_18542,N_13306);
nand U21182 (N_21182,N_16357,N_17478);
or U21183 (N_21183,N_12381,N_17416);
nand U21184 (N_21184,N_15970,N_11600);
or U21185 (N_21185,N_17426,N_13864);
and U21186 (N_21186,N_14557,N_17005);
or U21187 (N_21187,N_17661,N_11802);
and U21188 (N_21188,N_17650,N_10725);
nand U21189 (N_21189,N_15793,N_12028);
or U21190 (N_21190,N_19908,N_12338);
xor U21191 (N_21191,N_17071,N_11925);
and U21192 (N_21192,N_10358,N_19006);
xor U21193 (N_21193,N_11346,N_11220);
and U21194 (N_21194,N_15661,N_10952);
nand U21195 (N_21195,N_11935,N_17997);
or U21196 (N_21196,N_10197,N_17327);
nand U21197 (N_21197,N_17522,N_19326);
nor U21198 (N_21198,N_19729,N_18741);
and U21199 (N_21199,N_17220,N_14905);
nor U21200 (N_21200,N_19035,N_10649);
xor U21201 (N_21201,N_10015,N_12325);
xor U21202 (N_21202,N_13804,N_16947);
or U21203 (N_21203,N_16751,N_13808);
nand U21204 (N_21204,N_15436,N_12627);
xnor U21205 (N_21205,N_18553,N_17967);
nand U21206 (N_21206,N_15501,N_15801);
xnor U21207 (N_21207,N_15269,N_13782);
and U21208 (N_21208,N_12720,N_18774);
or U21209 (N_21209,N_17552,N_19822);
and U21210 (N_21210,N_19061,N_15700);
xnor U21211 (N_21211,N_14312,N_17111);
and U21212 (N_21212,N_16529,N_12579);
xnor U21213 (N_21213,N_17949,N_11517);
nor U21214 (N_21214,N_18254,N_10209);
nand U21215 (N_21215,N_17167,N_18156);
nand U21216 (N_21216,N_13449,N_18544);
xor U21217 (N_21217,N_12098,N_18377);
and U21218 (N_21218,N_11295,N_11943);
nand U21219 (N_21219,N_14703,N_14831);
and U21220 (N_21220,N_13530,N_17513);
nand U21221 (N_21221,N_17238,N_18321);
and U21222 (N_21222,N_19452,N_19868);
and U21223 (N_21223,N_11903,N_10008);
or U21224 (N_21224,N_14995,N_14565);
or U21225 (N_21225,N_15129,N_12032);
and U21226 (N_21226,N_19631,N_12374);
or U21227 (N_21227,N_13175,N_16530);
and U21228 (N_21228,N_19160,N_15434);
nand U21229 (N_21229,N_19296,N_12638);
xnor U21230 (N_21230,N_17945,N_11505);
nor U21231 (N_21231,N_13894,N_11669);
and U21232 (N_21232,N_17539,N_14082);
and U21233 (N_21233,N_10685,N_10608);
nor U21234 (N_21234,N_12207,N_12980);
nand U21235 (N_21235,N_16970,N_18430);
and U21236 (N_21236,N_19153,N_13942);
xor U21237 (N_21237,N_16082,N_18596);
xor U21238 (N_21238,N_16998,N_18328);
and U21239 (N_21239,N_18948,N_14241);
nor U21240 (N_21240,N_18118,N_14855);
xnor U21241 (N_21241,N_13901,N_10739);
nand U21242 (N_21242,N_14204,N_15988);
or U21243 (N_21243,N_16760,N_18578);
and U21244 (N_21244,N_18651,N_18869);
nand U21245 (N_21245,N_10198,N_16575);
nand U21246 (N_21246,N_18715,N_14014);
and U21247 (N_21247,N_10565,N_15295);
nand U21248 (N_21248,N_18359,N_19891);
nand U21249 (N_21249,N_13494,N_13656);
or U21250 (N_21250,N_16040,N_16954);
xor U21251 (N_21251,N_18533,N_12576);
nand U21252 (N_21252,N_13099,N_10007);
nand U21253 (N_21253,N_18906,N_19547);
nand U21254 (N_21254,N_18919,N_17128);
xor U21255 (N_21255,N_12409,N_11529);
nor U21256 (N_21256,N_12753,N_13391);
nor U21257 (N_21257,N_14805,N_12284);
nor U21258 (N_21258,N_16400,N_14543);
xor U21259 (N_21259,N_19887,N_19906);
xnor U21260 (N_21260,N_12082,N_19167);
nor U21261 (N_21261,N_17434,N_19511);
nor U21262 (N_21262,N_10819,N_18833);
nor U21263 (N_21263,N_12170,N_10881);
and U21264 (N_21264,N_15646,N_19670);
nor U21265 (N_21265,N_10533,N_16362);
and U21266 (N_21266,N_13789,N_19457);
xnor U21267 (N_21267,N_11286,N_17458);
nor U21268 (N_21268,N_10148,N_16318);
and U21269 (N_21269,N_16849,N_15035);
xor U21270 (N_21270,N_19212,N_17541);
nand U21271 (N_21271,N_14225,N_18209);
nand U21272 (N_21272,N_10791,N_10967);
and U21273 (N_21273,N_10744,N_18732);
and U21274 (N_21274,N_18463,N_16266);
xor U21275 (N_21275,N_12901,N_17631);
and U21276 (N_21276,N_16304,N_12875);
xor U21277 (N_21277,N_16102,N_14292);
nand U21278 (N_21278,N_16741,N_12305);
or U21279 (N_21279,N_15071,N_19040);
and U21280 (N_21280,N_15280,N_15817);
xor U21281 (N_21281,N_14920,N_18768);
nor U21282 (N_21282,N_18392,N_13288);
or U21283 (N_21283,N_16142,N_17502);
and U21284 (N_21284,N_13265,N_15386);
nand U21285 (N_21285,N_15432,N_13264);
nand U21286 (N_21286,N_10014,N_11125);
nand U21287 (N_21287,N_12900,N_10026);
nor U21288 (N_21288,N_11251,N_10111);
and U21289 (N_21289,N_10835,N_19180);
or U21290 (N_21290,N_19845,N_15311);
and U21291 (N_21291,N_13826,N_16750);
and U21292 (N_21292,N_18310,N_10140);
and U21293 (N_21293,N_12129,N_16403);
nor U21294 (N_21294,N_13636,N_11153);
nand U21295 (N_21295,N_17550,N_11849);
or U21296 (N_21296,N_16383,N_17297);
nor U21297 (N_21297,N_17104,N_17893);
xor U21298 (N_21298,N_17006,N_17598);
nor U21299 (N_21299,N_12183,N_19276);
xnor U21300 (N_21300,N_16191,N_10175);
xnor U21301 (N_21301,N_11335,N_17388);
nor U21302 (N_21302,N_13171,N_12653);
or U21303 (N_21303,N_19627,N_19665);
nor U21304 (N_21304,N_13471,N_12805);
and U21305 (N_21305,N_12333,N_10435);
or U21306 (N_21306,N_12263,N_18771);
xnor U21307 (N_21307,N_12943,N_12104);
nand U21308 (N_21308,N_13674,N_13839);
and U21309 (N_21309,N_13483,N_15760);
nand U21310 (N_21310,N_18052,N_19747);
nand U21311 (N_21311,N_12896,N_10524);
xor U21312 (N_21312,N_14083,N_12761);
nand U21313 (N_21313,N_11148,N_15575);
and U21314 (N_21314,N_16165,N_16916);
xnor U21315 (N_21315,N_11119,N_10329);
and U21316 (N_21316,N_13892,N_12113);
nand U21317 (N_21317,N_13678,N_14153);
nand U21318 (N_21318,N_13240,N_10942);
and U21319 (N_21319,N_14004,N_11518);
and U21320 (N_21320,N_12137,N_17258);
nand U21321 (N_21321,N_17333,N_16879);
nor U21322 (N_21322,N_14772,N_19207);
and U21323 (N_21323,N_11530,N_15167);
or U21324 (N_21324,N_15553,N_14705);
or U21325 (N_21325,N_19618,N_11969);
nand U21326 (N_21326,N_11101,N_19664);
xnor U21327 (N_21327,N_18969,N_17037);
and U21328 (N_21328,N_10570,N_15303);
and U21329 (N_21329,N_13061,N_16643);
nor U21330 (N_21330,N_13179,N_12373);
nand U21331 (N_21331,N_10874,N_15734);
nand U21332 (N_21332,N_11736,N_18271);
xor U21333 (N_21333,N_15499,N_11532);
nor U21334 (N_21334,N_12099,N_14984);
xor U21335 (N_21335,N_13537,N_16545);
and U21336 (N_21336,N_15399,N_13661);
nand U21337 (N_21337,N_14814,N_19330);
nand U21338 (N_21338,N_17157,N_10001);
nor U21339 (N_21339,N_13236,N_13697);
nor U21340 (N_21340,N_17207,N_11317);
or U21341 (N_21341,N_19391,N_16573);
nor U21342 (N_21342,N_17637,N_11777);
xnor U21343 (N_21343,N_13926,N_15486);
or U21344 (N_21344,N_13921,N_12501);
xor U21345 (N_21345,N_19114,N_12734);
xnor U21346 (N_21346,N_14600,N_16782);
nor U21347 (N_21347,N_13813,N_10812);
nand U21348 (N_21348,N_10098,N_17780);
and U21349 (N_21349,N_16164,N_12611);
nand U21350 (N_21350,N_16988,N_15173);
nand U21351 (N_21351,N_10641,N_18492);
and U21352 (N_21352,N_16592,N_19613);
and U21353 (N_21353,N_10440,N_19102);
xor U21354 (N_21354,N_19468,N_18727);
or U21355 (N_21355,N_13153,N_15214);
or U21356 (N_21356,N_16989,N_12109);
xor U21357 (N_21357,N_15778,N_17477);
or U21358 (N_21358,N_19027,N_11805);
or U21359 (N_21359,N_14918,N_17470);
nor U21360 (N_21360,N_11449,N_14332);
nor U21361 (N_21361,N_14295,N_13141);
xnor U21362 (N_21362,N_14220,N_13095);
or U21363 (N_21363,N_19037,N_14218);
xnor U21364 (N_21364,N_10786,N_16776);
nor U21365 (N_21365,N_15408,N_19561);
xor U21366 (N_21366,N_17781,N_15362);
xnor U21367 (N_21367,N_19030,N_17265);
xor U21368 (N_21368,N_10679,N_18097);
nand U21369 (N_21369,N_18527,N_16381);
nand U21370 (N_21370,N_18125,N_15335);
or U21371 (N_21371,N_15633,N_14555);
nand U21372 (N_21372,N_11511,N_16847);
nand U21373 (N_21373,N_11495,N_14983);
and U21374 (N_21374,N_18437,N_12936);
and U21375 (N_21375,N_11390,N_14061);
nor U21376 (N_21376,N_14723,N_15010);
and U21377 (N_21377,N_14764,N_17239);
nor U21378 (N_21378,N_14006,N_17174);
xor U21379 (N_21379,N_10096,N_16147);
and U21380 (N_21380,N_18363,N_18593);
and U21381 (N_21381,N_12463,N_11929);
nor U21382 (N_21382,N_12490,N_18587);
or U21383 (N_21383,N_19811,N_10117);
nor U21384 (N_21384,N_14315,N_15583);
nand U21385 (N_21385,N_14672,N_11345);
and U21386 (N_21386,N_14362,N_19059);
nand U21387 (N_21387,N_17801,N_11040);
nor U21388 (N_21388,N_19481,N_18613);
and U21389 (N_21389,N_16608,N_10469);
nor U21390 (N_21390,N_10587,N_14423);
and U21391 (N_21391,N_19635,N_16918);
and U21392 (N_21392,N_19344,N_11533);
or U21393 (N_21393,N_12243,N_15446);
xnor U21394 (N_21394,N_11702,N_13071);
or U21395 (N_21395,N_19944,N_11992);
nand U21396 (N_21396,N_15440,N_15373);
xnor U21397 (N_21397,N_15026,N_10076);
or U21398 (N_21398,N_17754,N_18972);
nand U21399 (N_21399,N_14847,N_16296);
nor U21400 (N_21400,N_17621,N_17440);
and U21401 (N_21401,N_16340,N_18030);
nand U21402 (N_21402,N_13304,N_13715);
nor U21403 (N_21403,N_13154,N_15807);
nor U21404 (N_21404,N_15144,N_16595);
xnor U21405 (N_21405,N_11671,N_11602);
nor U21406 (N_21406,N_16248,N_15756);
xnor U21407 (N_21407,N_19399,N_11571);
and U21408 (N_21408,N_16930,N_14564);
nand U21409 (N_21409,N_15454,N_10817);
or U21410 (N_21410,N_17292,N_16361);
xor U21411 (N_21411,N_19687,N_11859);
nand U21412 (N_21412,N_11482,N_10234);
and U21413 (N_21413,N_17281,N_10477);
and U21414 (N_21414,N_11791,N_18505);
and U21415 (N_21415,N_10012,N_13234);
nor U21416 (N_21416,N_13818,N_14262);
xor U21417 (N_21417,N_17843,N_17817);
xnor U21418 (N_21418,N_11950,N_19329);
and U21419 (N_21419,N_19308,N_12819);
and U21420 (N_21420,N_15105,N_12259);
or U21421 (N_21421,N_12062,N_12285);
or U21422 (N_21422,N_10803,N_13597);
nor U21423 (N_21423,N_17177,N_11775);
nand U21424 (N_21424,N_16687,N_10146);
xor U21425 (N_21425,N_11763,N_10095);
and U21426 (N_21426,N_18736,N_17444);
xor U21427 (N_21427,N_15050,N_19063);
and U21428 (N_21428,N_18074,N_12551);
nand U21429 (N_21429,N_14474,N_16295);
and U21430 (N_21430,N_12778,N_18516);
or U21431 (N_21431,N_19306,N_13557);
nand U21432 (N_21432,N_12365,N_17318);
or U21433 (N_21433,N_19742,N_14790);
nor U21434 (N_21434,N_19981,N_16157);
xnor U21435 (N_21435,N_18096,N_10164);
nand U21436 (N_21436,N_15363,N_12254);
nor U21437 (N_21437,N_19791,N_19794);
or U21438 (N_21438,N_13861,N_15946);
xor U21439 (N_21439,N_13017,N_11219);
xnor U21440 (N_21440,N_13409,N_14977);
nor U21441 (N_21441,N_19495,N_18455);
nand U21442 (N_21442,N_16624,N_17147);
or U21443 (N_21443,N_19335,N_12011);
nor U21444 (N_21444,N_17877,N_17196);
nand U21445 (N_21445,N_14852,N_10288);
xnor U21446 (N_21446,N_19267,N_17578);
and U21447 (N_21447,N_14768,N_14099);
and U21448 (N_21448,N_18033,N_19806);
nor U21449 (N_21449,N_17112,N_10328);
or U21450 (N_21450,N_12308,N_18200);
and U21451 (N_21451,N_13386,N_10600);
or U21452 (N_21452,N_18585,N_17051);
and U21453 (N_21453,N_17549,N_14641);
nand U21454 (N_21454,N_14909,N_19305);
and U21455 (N_21455,N_12985,N_14746);
xor U21456 (N_21456,N_18871,N_10020);
nor U21457 (N_21457,N_19074,N_15958);
xnor U21458 (N_21458,N_14037,N_11589);
or U21459 (N_21459,N_10019,N_13599);
and U21460 (N_21460,N_15764,N_13005);
nand U21461 (N_21461,N_10964,N_13895);
nand U21462 (N_21462,N_17074,N_15718);
or U21463 (N_21463,N_11708,N_17626);
and U21464 (N_21464,N_12087,N_15877);
xor U21465 (N_21465,N_18454,N_18000);
nand U21466 (N_21466,N_13461,N_16382);
and U21467 (N_21467,N_14670,N_15243);
or U21468 (N_21468,N_17871,N_14271);
xor U21469 (N_21469,N_18657,N_13255);
and U21470 (N_21470,N_11100,N_15875);
nor U21471 (N_21471,N_10156,N_10489);
xnor U21472 (N_21472,N_12440,N_12931);
xor U21473 (N_21473,N_11041,N_11410);
xor U21474 (N_21474,N_13013,N_11872);
xor U21475 (N_21475,N_12219,N_18974);
xnor U21476 (N_21476,N_15901,N_12789);
xnor U21477 (N_21477,N_13801,N_12388);
xor U21478 (N_21478,N_18712,N_10487);
xor U21479 (N_21479,N_17326,N_11014);
xor U21480 (N_21480,N_18204,N_17135);
xor U21481 (N_21481,N_15383,N_18325);
xor U21482 (N_21482,N_14391,N_17182);
xnor U21483 (N_21483,N_13604,N_19098);
nand U21484 (N_21484,N_10509,N_10938);
and U21485 (N_21485,N_11471,N_12159);
nand U21486 (N_21486,N_17778,N_16179);
nand U21487 (N_21487,N_14465,N_13200);
xor U21488 (N_21488,N_19470,N_12898);
nor U21489 (N_21489,N_13305,N_10349);
nor U21490 (N_21490,N_17245,N_19154);
xor U21491 (N_21491,N_10854,N_18360);
or U21492 (N_21492,N_19818,N_12929);
nor U21493 (N_21493,N_14668,N_15430);
and U21494 (N_21494,N_16265,N_12852);
and U21495 (N_21495,N_18113,N_16037);
nor U21496 (N_21496,N_12071,N_16704);
or U21497 (N_21497,N_19304,N_15708);
or U21498 (N_21498,N_11231,N_17307);
or U21499 (N_21499,N_18946,N_11378);
and U21500 (N_21500,N_17663,N_15435);
and U21501 (N_21501,N_16263,N_16859);
xnor U21502 (N_21502,N_19042,N_10977);
xnor U21503 (N_21503,N_18641,N_17305);
or U21504 (N_21504,N_15011,N_13595);
and U21505 (N_21505,N_18834,N_13254);
xor U21506 (N_21506,N_18274,N_12992);
and U21507 (N_21507,N_12066,N_10191);
xor U21508 (N_21508,N_19973,N_16623);
and U21509 (N_21509,N_15420,N_12044);
nand U21510 (N_21510,N_19134,N_11438);
nand U21511 (N_21511,N_19397,N_11981);
nand U21512 (N_21512,N_14080,N_16114);
xor U21513 (N_21513,N_14577,N_19269);
xor U21514 (N_21514,N_10589,N_14478);
nor U21515 (N_21515,N_16346,N_15458);
nor U21516 (N_21516,N_13766,N_17250);
xor U21517 (N_21517,N_14125,N_12786);
nor U21518 (N_21518,N_12122,N_10320);
or U21519 (N_21519,N_14773,N_12527);
nand U21520 (N_21520,N_16369,N_11357);
xor U21521 (N_21521,N_14425,N_10858);
xnor U21522 (N_21522,N_10759,N_17686);
nand U21523 (N_21523,N_16093,N_11420);
xnor U21524 (N_21524,N_14904,N_13452);
and U21525 (N_21525,N_12324,N_16445);
xnor U21526 (N_21526,N_19988,N_13857);
nand U21527 (N_21527,N_17654,N_14892);
and U21528 (N_21528,N_11781,N_18965);
nor U21529 (N_21529,N_17602,N_13359);
nor U21530 (N_21530,N_12251,N_16973);
or U21531 (N_21531,N_14573,N_11150);
nor U21532 (N_21532,N_16138,N_13512);
nand U21533 (N_21533,N_17760,N_16899);
and U21534 (N_21534,N_15530,N_12697);
xnor U21535 (N_21535,N_14472,N_18532);
nor U21536 (N_21536,N_13068,N_16150);
or U21537 (N_21537,N_11711,N_14837);
and U21538 (N_21538,N_11182,N_12744);
nand U21539 (N_21539,N_19298,N_13954);
or U21540 (N_21540,N_16376,N_13948);
nand U21541 (N_21541,N_17990,N_19902);
or U21542 (N_21542,N_11027,N_15380);
xnor U21543 (N_21543,N_13351,N_12133);
and U21544 (N_21544,N_11076,N_11169);
xor U21545 (N_21545,N_18550,N_11503);
or U21546 (N_21546,N_18215,N_14917);
and U21547 (N_21547,N_18880,N_19654);
nand U21548 (N_21548,N_12320,N_13299);
or U21549 (N_21549,N_17487,N_10984);
xor U21550 (N_21550,N_15174,N_18729);
nor U21551 (N_21551,N_12619,N_16672);
nand U21552 (N_21552,N_11109,N_15890);
xor U21553 (N_21553,N_17527,N_18916);
xnor U21554 (N_21554,N_12702,N_13806);
and U21555 (N_21555,N_17067,N_17165);
or U21556 (N_21556,N_15976,N_16514);
or U21557 (N_21557,N_14047,N_10855);
or U21558 (N_21558,N_14719,N_16716);
nand U21559 (N_21559,N_11285,N_13739);
nand U21560 (N_21560,N_15152,N_10584);
nor U21561 (N_21561,N_19438,N_18269);
and U21562 (N_21562,N_13272,N_18404);
xor U21563 (N_21563,N_14257,N_14128);
nor U21564 (N_21564,N_12351,N_16699);
nand U21565 (N_21565,N_11639,N_17114);
nor U21566 (N_21566,N_12966,N_18402);
or U21567 (N_21567,N_11592,N_15070);
and U21568 (N_21568,N_13906,N_15088);
nor U21569 (N_21569,N_15437,N_19060);
nand U21570 (N_21570,N_19909,N_17055);
or U21571 (N_21571,N_10413,N_12216);
nor U21572 (N_21572,N_17545,N_13019);
and U21573 (N_21573,N_12925,N_16454);
xor U21574 (N_21574,N_10677,N_19436);
xnor U21575 (N_21575,N_11964,N_12687);
xnor U21576 (N_21576,N_15033,N_13764);
or U21577 (N_21577,N_19292,N_16621);
or U21578 (N_21578,N_18448,N_18720);
and U21579 (N_21579,N_12274,N_12602);
and U21580 (N_21580,N_17645,N_16833);
and U21581 (N_21581,N_11140,N_15580);
nand U21582 (N_21582,N_15325,N_14081);
nand U21583 (N_21583,N_11611,N_16022);
or U21584 (N_21584,N_11374,N_12669);
nand U21585 (N_21585,N_16961,N_17558);
and U21586 (N_21586,N_14017,N_10940);
or U21587 (N_21587,N_15039,N_14661);
and U21588 (N_21588,N_18380,N_17751);
xor U21589 (N_21589,N_11564,N_16712);
xnor U21590 (N_21590,N_18726,N_13328);
and U21591 (N_21591,N_12398,N_10743);
or U21592 (N_21592,N_13329,N_13490);
or U21593 (N_21593,N_19270,N_15052);
or U21594 (N_21594,N_15843,N_11470);
xnor U21595 (N_21595,N_11187,N_14008);
nor U21596 (N_21596,N_15971,N_17146);
and U21597 (N_21597,N_15345,N_10935);
xor U21598 (N_21598,N_14255,N_18868);
or U21599 (N_21599,N_15815,N_13064);
or U21600 (N_21600,N_10537,N_11344);
or U21601 (N_21601,N_17271,N_18406);
nand U21602 (N_21602,N_19792,N_11856);
nor U21603 (N_21603,N_17976,N_19382);
or U21604 (N_21604,N_11967,N_19359);
and U21605 (N_21605,N_12655,N_12293);
nor U21606 (N_21606,N_11848,N_15896);
nor U21607 (N_21607,N_10525,N_12143);
or U21608 (N_21608,N_11016,N_11852);
and U21609 (N_21609,N_18798,N_16650);
and U21610 (N_21610,N_18089,N_18583);
nand U21611 (N_21611,N_11865,N_18592);
nor U21612 (N_21612,N_16272,N_18696);
and U21613 (N_21613,N_14754,N_15650);
nand U21614 (N_21614,N_17936,N_10462);
nor U21615 (N_21615,N_16842,N_13571);
xor U21616 (N_21616,N_14715,N_10266);
or U21617 (N_21617,N_14561,N_19360);
nor U21618 (N_21618,N_11196,N_16804);
or U21619 (N_21619,N_19803,N_12738);
nor U21620 (N_21620,N_14086,N_17928);
xnor U21621 (N_21621,N_14710,N_19288);
nor U21622 (N_21622,N_12856,N_16874);
and U21623 (N_21623,N_14583,N_12298);
nor U21624 (N_21624,N_12963,N_16830);
or U21625 (N_21625,N_19780,N_19997);
nor U21626 (N_21626,N_13393,N_10948);
or U21627 (N_21627,N_18027,N_14863);
and U21628 (N_21628,N_16218,N_13078);
nor U21629 (N_21629,N_16352,N_19065);
and U21630 (N_21630,N_11012,N_10302);
and U21631 (N_21631,N_18523,N_16763);
nand U21632 (N_21632,N_14001,N_10591);
nand U21633 (N_21633,N_15777,N_19469);
and U21634 (N_21634,N_13743,N_16139);
nor U21635 (N_21635,N_16439,N_12161);
nor U21636 (N_21636,N_11080,N_12840);
xnor U21637 (N_21637,N_18608,N_13477);
or U21638 (N_21638,N_11397,N_11297);
and U21639 (N_21639,N_14177,N_14669);
or U21640 (N_21640,N_15318,N_19824);
xor U21641 (N_21641,N_14263,N_17756);
xnor U21642 (N_21642,N_13112,N_13800);
or U21643 (N_21643,N_16785,N_10866);
xnor U21644 (N_21644,N_14642,N_19442);
xnor U21645 (N_21645,N_14396,N_17183);
xor U21646 (N_21646,N_19543,N_15742);
xor U21647 (N_21647,N_11979,N_16579);
or U21648 (N_21648,N_11507,N_14587);
xor U21649 (N_21649,N_18307,N_11038);
nand U21650 (N_21650,N_15951,N_18121);
or U21651 (N_21651,N_13503,N_14725);
nand U21652 (N_21652,N_16201,N_16499);
and U21653 (N_21653,N_12713,N_19963);
and U21654 (N_21654,N_14728,N_15737);
or U21655 (N_21655,N_11906,N_17476);
nor U21656 (N_21656,N_18655,N_16620);
nor U21657 (N_21657,N_18646,N_17162);
nand U21658 (N_21658,N_10612,N_17855);
or U21659 (N_21659,N_13262,N_16684);
nor U21660 (N_21660,N_15949,N_15194);
nor U21661 (N_21661,N_17397,N_11073);
xor U21662 (N_21662,N_10260,N_11987);
xor U21663 (N_21663,N_13237,N_15037);
or U21664 (N_21664,N_19108,N_19509);
nand U21665 (N_21665,N_16864,N_19418);
or U21666 (N_21666,N_10488,N_11609);
and U21667 (N_21667,N_15765,N_19459);
and U21668 (N_21668,N_17863,N_17557);
nand U21669 (N_21669,N_16755,N_19926);
or U21670 (N_21670,N_12385,N_18366);
nor U21671 (N_21671,N_18116,N_13905);
nor U21672 (N_21672,N_13623,N_11994);
and U21673 (N_21673,N_16775,N_15206);
or U21674 (N_21674,N_12776,N_16463);
nand U21675 (N_21675,N_15125,N_11130);
nand U21676 (N_21676,N_14595,N_15903);
nand U21677 (N_21677,N_16280,N_17031);
and U21678 (N_21678,N_17799,N_17348);
or U21679 (N_21679,N_15547,N_12714);
and U21680 (N_21680,N_19744,N_14403);
and U21681 (N_21681,N_14084,N_11070);
nand U21682 (N_21682,N_17655,N_13919);
xnor U21683 (N_21683,N_16563,N_16151);
and U21684 (N_21684,N_17380,N_12200);
or U21685 (N_21685,N_14305,N_10455);
and U21686 (N_21686,N_13196,N_11569);
or U21687 (N_21687,N_13507,N_12156);
or U21688 (N_21688,N_10085,N_19328);
or U21689 (N_21689,N_15496,N_16577);
or U21690 (N_21690,N_17301,N_14395);
nand U21691 (N_21691,N_13538,N_13835);
and U21692 (N_21692,N_17284,N_12172);
nor U21693 (N_21693,N_17856,N_13946);
nand U21694 (N_21694,N_15451,N_15878);
xnor U21695 (N_21695,N_10045,N_15419);
xnor U21696 (N_21696,N_19913,N_14980);
nand U21697 (N_21697,N_18571,N_13139);
xor U21698 (N_21698,N_18460,N_13415);
and U21699 (N_21699,N_16747,N_16517);
nand U21700 (N_21700,N_14946,N_11270);
nand U21701 (N_21701,N_11426,N_18996);
nor U21702 (N_21702,N_18807,N_18435);
nand U21703 (N_21703,N_17484,N_18353);
nor U21704 (N_21704,N_12328,N_12245);
xor U21705 (N_21705,N_18017,N_13910);
or U21706 (N_21706,N_19896,N_18955);
xnor U21707 (N_21707,N_11729,N_14318);
xor U21708 (N_21708,N_10359,N_16546);
nor U21709 (N_21709,N_17121,N_13559);
and U21710 (N_21710,N_16078,N_12507);
nand U21711 (N_21711,N_11675,N_17294);
nand U21712 (N_21712,N_15558,N_17253);
nand U21713 (N_21713,N_17251,N_19149);
and U21714 (N_21714,N_16653,N_12154);
or U21715 (N_21715,N_15250,N_16247);
xor U21716 (N_21716,N_18885,N_12244);
xor U21717 (N_21717,N_11696,N_17891);
xnor U21718 (N_21718,N_15385,N_11516);
or U21719 (N_21719,N_15225,N_15337);
xnor U21720 (N_21720,N_13730,N_17681);
or U21721 (N_21721,N_13827,N_14525);
nand U21722 (N_21722,N_14567,N_15738);
nor U21723 (N_21723,N_15516,N_17009);
nor U21724 (N_21724,N_12088,N_11835);
nand U21725 (N_21725,N_13565,N_16299);
nor U21726 (N_21726,N_19336,N_15199);
and U21727 (N_21727,N_11033,N_12663);
xnor U21728 (N_21728,N_17881,N_17772);
nand U21729 (N_21729,N_18581,N_10281);
xnor U21730 (N_21730,N_10405,N_15086);
nand U21731 (N_21731,N_17528,N_14865);
nor U21732 (N_21732,N_10789,N_15098);
nor U21733 (N_21733,N_11144,N_11776);
and U21734 (N_21734,N_16793,N_19738);
or U21735 (N_21735,N_16656,N_12468);
and U21736 (N_21736,N_12589,N_18195);
or U21737 (N_21737,N_19375,N_16395);
xor U21738 (N_21738,N_16154,N_16786);
nor U21739 (N_21739,N_10999,N_12837);
nor U21740 (N_21740,N_14878,N_11113);
xnor U21741 (N_21741,N_10230,N_13197);
or U21742 (N_21742,N_13580,N_10025);
nand U21743 (N_21743,N_16363,N_14151);
nand U21744 (N_21744,N_14245,N_10213);
xor U21745 (N_21745,N_19764,N_15475);
nand U21746 (N_21746,N_14834,N_15543);
xor U21747 (N_21747,N_14795,N_13810);
and U21748 (N_21748,N_11544,N_14462);
xnor U21749 (N_21749,N_13869,N_12220);
and U21750 (N_21750,N_19607,N_14411);
xnor U21751 (N_21751,N_16796,N_16425);
or U21752 (N_21752,N_15089,N_13727);
nand U21753 (N_21753,N_14975,N_10419);
nor U21754 (N_21754,N_12072,N_10737);
nor U21755 (N_21755,N_16430,N_14602);
xnor U21756 (N_21756,N_18461,N_16325);
and U21757 (N_21757,N_19041,N_10464);
nand U21758 (N_21758,N_14279,N_18294);
nor U21759 (N_21759,N_12075,N_13230);
or U21760 (N_21760,N_19230,N_16025);
or U21761 (N_21761,N_17573,N_17218);
or U21762 (N_21762,N_12588,N_14267);
nand U21763 (N_21763,N_16903,N_17875);
xnor U21764 (N_21764,N_10205,N_14815);
nand U21765 (N_21765,N_10996,N_13292);
or U21766 (N_21766,N_15153,N_18111);
nor U21767 (N_21767,N_10502,N_16448);
nand U21768 (N_21768,N_12473,N_18264);
nand U21769 (N_21769,N_13635,N_16503);
and U21770 (N_21770,N_15204,N_17804);
xnor U21771 (N_21771,N_17349,N_10618);
and U21772 (N_21772,N_14209,N_13779);
or U21773 (N_21773,N_11386,N_19516);
nand U21774 (N_21774,N_12618,N_18707);
or U21775 (N_21775,N_15894,N_13998);
nor U21776 (N_21776,N_11439,N_17264);
xor U21777 (N_21777,N_19206,N_17561);
and U21778 (N_21778,N_18557,N_12595);
nand U21779 (N_21779,N_14806,N_10255);
and U21780 (N_21780,N_13514,N_16759);
or U21781 (N_21781,N_11880,N_15560);
nand U21782 (N_21782,N_16193,N_10884);
nor U21783 (N_21783,N_14700,N_16691);
nand U21784 (N_21784,N_13548,N_16232);
nand U21785 (N_21785,N_19800,N_18015);
or U21786 (N_21786,N_17198,N_13205);
and U21787 (N_21787,N_15928,N_18367);
and U21788 (N_21788,N_12347,N_16055);
and U21789 (N_21789,N_13107,N_14507);
xnor U21790 (N_21790,N_10797,N_16742);
or U21791 (N_21791,N_11343,N_13294);
nor U21792 (N_21792,N_12265,N_15897);
nor U21793 (N_21793,N_11277,N_16087);
xor U21794 (N_21794,N_19563,N_10381);
xor U21795 (N_21795,N_12416,N_10355);
and U21796 (N_21796,N_19848,N_15608);
or U21797 (N_21797,N_17381,N_17329);
or U21798 (N_21798,N_18108,N_12754);
nand U21799 (N_21799,N_10958,N_13434);
nor U21800 (N_21800,N_18700,N_14942);
xor U21801 (N_21801,N_17665,N_11122);
and U21802 (N_21802,N_17344,N_15304);
and U21803 (N_21803,N_16094,N_15425);
nand U21804 (N_21804,N_18582,N_16064);
or U21805 (N_21805,N_15382,N_16707);
xor U21806 (N_21806,N_17953,N_15975);
nand U21807 (N_21807,N_10046,N_19629);
nand U21808 (N_21808,N_15371,N_13547);
nand U21809 (N_21809,N_19782,N_16767);
nand U21810 (N_21810,N_13338,N_19259);
xnor U21811 (N_21811,N_11924,N_19784);
and U21812 (N_21812,N_19535,N_11492);
or U21813 (N_21813,N_12018,N_10070);
xor U21814 (N_21814,N_15087,N_10720);
nor U21815 (N_21815,N_14866,N_18329);
and U21816 (N_21816,N_18290,N_13160);
nand U21817 (N_21817,N_15519,N_11486);
or U21818 (N_21818,N_11658,N_14724);
or U21819 (N_21819,N_17129,N_18040);
or U21820 (N_21820,N_17588,N_11588);
nand U21821 (N_21821,N_15541,N_17955);
or U21822 (N_21822,N_13758,N_13676);
nor U21823 (N_21823,N_19532,N_14721);
nand U21824 (N_21824,N_11272,N_18739);
nand U21825 (N_21825,N_18815,N_12448);
nand U21826 (N_21826,N_10128,N_17794);
or U21827 (N_21827,N_18250,N_16827);
nand U21828 (N_21828,N_15891,N_15581);
nor U21829 (N_21829,N_19467,N_19593);
or U21830 (N_21830,N_14536,N_16103);
or U21831 (N_21831,N_15470,N_13736);
and U21832 (N_21832,N_13528,N_18300);
and U21833 (N_21833,N_17141,N_13870);
or U21834 (N_21834,N_16240,N_12766);
or U21835 (N_21835,N_18104,N_13844);
nand U21836 (N_21836,N_13638,N_16402);
or U21837 (N_21837,N_15550,N_10366);
nor U21838 (N_21838,N_11831,N_17825);
nor U21839 (N_21839,N_16855,N_11131);
nand U21840 (N_21840,N_10021,N_17933);
and U21841 (N_21841,N_19284,N_19785);
nor U21842 (N_21842,N_13281,N_12509);
xor U21843 (N_21843,N_16977,N_15703);
or U21844 (N_21844,N_10451,N_15888);
xor U21845 (N_21845,N_19294,N_10724);
nand U21846 (N_21846,N_17543,N_19044);
nor U21847 (N_21847,N_18914,N_11704);
and U21848 (N_21848,N_15678,N_13056);
nand U21849 (N_21849,N_13470,N_14850);
xnor U21850 (N_21850,N_10508,N_12063);
and U21851 (N_21851,N_11934,N_19024);
nor U21852 (N_21852,N_18375,N_16019);
nor U21853 (N_21853,N_18142,N_14791);
xor U21854 (N_21854,N_12747,N_12519);
and U21855 (N_21855,N_18144,N_13103);
nor U21856 (N_21856,N_19246,N_19332);
nor U21857 (N_21857,N_17088,N_18019);
nor U21858 (N_21858,N_17846,N_19771);
nand U21859 (N_21859,N_13561,N_13221);
or U21860 (N_21860,N_19113,N_15353);
nor U21861 (N_21861,N_18449,N_19632);
nand U21862 (N_21862,N_16012,N_11966);
nor U21863 (N_21863,N_12008,N_13256);
xor U21864 (N_21864,N_14523,N_15252);
nor U21865 (N_21865,N_17965,N_11502);
nand U21866 (N_21866,N_19175,N_13377);
nand U21867 (N_21867,N_14152,N_13169);
and U21868 (N_21868,N_18951,N_11487);
and U21869 (N_21869,N_16241,N_16566);
xor U21870 (N_21870,N_10218,N_13532);
and U21871 (N_21871,N_12748,N_13008);
xnor U21872 (N_21872,N_16261,N_18247);
xnor U21873 (N_21873,N_17571,N_13917);
nand U21874 (N_21874,N_12978,N_10087);
nor U21875 (N_21875,N_18679,N_13253);
nand U21876 (N_21876,N_13463,N_16580);
nand U21877 (N_21877,N_15889,N_12735);
or U21878 (N_21878,N_14693,N_13845);
xnor U21879 (N_21879,N_18825,N_18904);
xnor U21880 (N_21880,N_12043,N_19279);
nand U21881 (N_21881,N_17716,N_18851);
xnor U21882 (N_21882,N_15825,N_14450);
and U21883 (N_21883,N_19842,N_16881);
nor U21884 (N_21884,N_11555,N_18201);
nand U21885 (N_21885,N_12331,N_19646);
nor U21886 (N_21886,N_11063,N_14019);
or U21887 (N_21887,N_10322,N_16678);
xor U21888 (N_21888,N_17580,N_19763);
nor U21889 (N_21889,N_19955,N_18503);
nand U21890 (N_21890,N_15047,N_12859);
and U21891 (N_21891,N_14796,N_10684);
nand U21892 (N_21892,N_10714,N_19591);
nand U21893 (N_21893,N_15163,N_10134);
xor U21894 (N_21894,N_15769,N_11510);
or U21895 (N_21895,N_15873,N_10501);
or U21896 (N_21896,N_11322,N_12511);
and U21897 (N_21897,N_18007,N_16778);
nor U21898 (N_21898,N_19017,N_17407);
nand U21899 (N_21899,N_17512,N_14870);
xnor U21900 (N_21900,N_10242,N_11128);
nor U21901 (N_21901,N_13663,N_16083);
nor U21902 (N_21902,N_17610,N_14143);
and U21903 (N_21903,N_17243,N_19253);
and U21904 (N_21904,N_10422,N_16419);
nand U21905 (N_21905,N_12914,N_15731);
nor U21906 (N_21906,N_17784,N_13440);
or U21907 (N_21907,N_13031,N_15166);
nor U21908 (N_21908,N_18970,N_13950);
xnor U21909 (N_21909,N_17740,N_11399);
and U21910 (N_21910,N_19989,N_12013);
and U21911 (N_21911,N_17739,N_12134);
or U21912 (N_21912,N_14431,N_16061);
xnor U21913 (N_21913,N_19814,N_14500);
xnor U21914 (N_21914,N_14617,N_15282);
and U21915 (N_21915,N_15851,N_15523);
or U21916 (N_21916,N_19487,N_13086);
nand U21917 (N_21917,N_11595,N_19215);
and U21918 (N_21918,N_14345,N_10135);
nand U21919 (N_21919,N_15835,N_16161);
or U21920 (N_21920,N_16700,N_11060);
or U21921 (N_21921,N_11218,N_18755);
nor U21922 (N_21922,N_14370,N_17194);
nand U21923 (N_21923,N_11677,N_12111);
nor U21924 (N_21924,N_17226,N_15238);
xnor U21925 (N_21925,N_14485,N_11444);
nor U21926 (N_21926,N_16276,N_18534);
or U21927 (N_21927,N_18467,N_10278);
nand U21928 (N_21928,N_17197,N_11797);
and U21929 (N_21929,N_10486,N_18094);
or U21930 (N_21930,N_10418,N_18275);
nor U21931 (N_21931,N_14544,N_11333);
nor U21932 (N_21932,N_12780,N_17448);
xnor U21933 (N_21933,N_14011,N_11626);
nor U21934 (N_21934,N_17035,N_18280);
nor U21935 (N_21935,N_10292,N_13673);
and U21936 (N_21936,N_19319,N_10185);
nand U21937 (N_21937,N_13077,N_19728);
nor U21938 (N_21938,N_16007,N_15265);
or U21939 (N_21939,N_13637,N_15674);
and U21940 (N_21940,N_13829,N_14619);
nor U21941 (N_21941,N_19026,N_11798);
or U21942 (N_21942,N_17687,N_13223);
and U21943 (N_21943,N_12495,N_19056);
nor U21944 (N_21944,N_13018,N_12271);
nor U21945 (N_21945,N_15180,N_11290);
xor U21946 (N_21946,N_11936,N_15804);
or U21947 (N_21947,N_19701,N_13639);
xnor U21948 (N_21948,N_17404,N_14792);
nand U21949 (N_21949,N_13607,N_16655);
nand U21950 (N_21950,N_14418,N_18638);
nor U21951 (N_21951,N_10905,N_17026);
nor U21952 (N_21952,N_16330,N_10926);
or U21953 (N_21953,N_10742,N_12144);
or U21954 (N_21954,N_16384,N_19714);
or U21955 (N_21955,N_14189,N_13991);
xnor U21956 (N_21956,N_16519,N_12545);
nor U21957 (N_21957,N_15989,N_15666);
nand U21958 (N_21958,N_13716,N_19974);
and U21959 (N_21959,N_14800,N_16972);
xor U21960 (N_21960,N_17376,N_15076);
and U21961 (N_21961,N_14650,N_17827);
and U21962 (N_21962,N_11352,N_12169);
xnor U21963 (N_21963,N_10838,N_15061);
nand U21964 (N_21964,N_18251,N_15867);
and U21965 (N_21965,N_18598,N_17982);
xor U21966 (N_21966,N_10406,N_13161);
or U21967 (N_21967,N_19877,N_11659);
nor U21968 (N_21968,N_11557,N_19372);
nand U21969 (N_21969,N_13191,N_17175);
nand U21970 (N_21970,N_18831,N_11876);
or U21971 (N_21971,N_19622,N_10071);
nand U21972 (N_21972,N_15556,N_12103);
or U21973 (N_21973,N_10048,N_16616);
xor U21974 (N_21974,N_10332,N_11829);
and U21975 (N_21975,N_16518,N_12102);
and U21976 (N_21976,N_10664,N_10766);
or U21977 (N_21977,N_18445,N_16722);
xor U21978 (N_21978,N_15929,N_15154);
xor U21979 (N_21979,N_16443,N_10385);
nand U21980 (N_21980,N_14058,N_19795);
or U21981 (N_21981,N_19023,N_12369);
or U21982 (N_21982,N_14738,N_12683);
and U21983 (N_21983,N_18635,N_12630);
and U21984 (N_21984,N_19726,N_18236);
nand U21985 (N_21985,N_14147,N_17231);
and U21986 (N_21986,N_12921,N_13430);
nor U21987 (N_21987,N_16398,N_17382);
and U21988 (N_21988,N_14887,N_15251);
and U21989 (N_21989,N_18182,N_15814);
and U21990 (N_21990,N_15938,N_14299);
nand U21991 (N_21991,N_12675,N_19003);
xnor U21992 (N_21992,N_17766,N_18411);
nor U21993 (N_21993,N_14188,N_15456);
nor U21994 (N_21994,N_11572,N_14172);
nand U21995 (N_21995,N_11778,N_19402);
xor U21996 (N_21996,N_11962,N_19260);
nor U21997 (N_21997,N_11646,N_17423);
nor U21998 (N_21998,N_13307,N_16355);
xnor U21999 (N_21999,N_19612,N_13055);
and U22000 (N_22000,N_14252,N_18150);
nand U22001 (N_22001,N_15974,N_14102);
and U22002 (N_22002,N_17176,N_11792);
nor U22003 (N_22003,N_12415,N_17320);
or U22004 (N_22004,N_19733,N_13668);
xor U22005 (N_22005,N_17062,N_13648);
nand U22006 (N_22006,N_11837,N_17241);
and U22007 (N_22007,N_13241,N_12148);
xnor U22008 (N_22008,N_18330,N_13036);
xnor U22009 (N_22009,N_14039,N_19374);
or U22010 (N_22010,N_19474,N_15842);
xor U22011 (N_22011,N_14614,N_10514);
nand U22012 (N_22012,N_17341,N_16867);
or U22013 (N_22013,N_14520,N_10147);
or U22014 (N_22014,N_14164,N_12872);
nand U22015 (N_22015,N_10650,N_18978);
and U22016 (N_22016,N_11211,N_15536);
nand U22017 (N_22017,N_17744,N_18703);
xnor U22018 (N_22018,N_15681,N_10976);
nor U22019 (N_22019,N_19348,N_15495);
and U22020 (N_22020,N_11662,N_17252);
nor U22021 (N_22021,N_14779,N_12301);
or U22022 (N_22022,N_17357,N_13485);
nand U22023 (N_22023,N_18627,N_15288);
and U22024 (N_22024,N_13940,N_15202);
nor U22025 (N_22025,N_13219,N_14607);
xnor U22026 (N_22026,N_18405,N_14654);
nor U22027 (N_22027,N_14229,N_13276);
or U22028 (N_22028,N_12999,N_14712);
nor U22029 (N_22029,N_14634,N_10824);
and U22030 (N_22030,N_15639,N_12221);
and U22031 (N_22031,N_17019,N_18143);
and U22032 (N_22032,N_16906,N_12287);
and U22033 (N_22033,N_10473,N_16938);
xor U22034 (N_22034,N_10180,N_19774);
and U22035 (N_22035,N_17944,N_18266);
nor U22036 (N_22036,N_17237,N_18661);
or U22037 (N_22037,N_10982,N_18513);
or U22038 (N_22038,N_19072,N_12871);
xnor U22039 (N_22039,N_15283,N_17255);
or U22040 (N_22040,N_15697,N_11015);
and U22041 (N_22041,N_19837,N_19394);
nand U22042 (N_22042,N_11223,N_10244);
nor U22043 (N_22043,N_10500,N_12965);
or U22044 (N_22044,N_13860,N_14405);
or U22045 (N_22045,N_18624,N_14268);
and U22046 (N_22046,N_10018,N_15058);
and U22047 (N_22047,N_18506,N_17758);
and U22048 (N_22048,N_17247,N_19876);
nor U22049 (N_22049,N_17753,N_14572);
xnor U22050 (N_22050,N_10296,N_10864);
nor U22051 (N_22051,N_10084,N_11456);
and U22052 (N_22052,N_10208,N_19956);
nand U22053 (N_22053,N_11166,N_10139);
nor U22054 (N_22054,N_12557,N_17137);
or U22055 (N_22055,N_12874,N_14823);
nor U22056 (N_22056,N_15679,N_17912);
and U22057 (N_22057,N_19032,N_18295);
nor U22058 (N_22058,N_15987,N_19526);
nor U22059 (N_22059,N_18967,N_14782);
xor U22060 (N_22060,N_17599,N_12915);
xor U22061 (N_22061,N_14475,N_15959);
nand U22062 (N_22062,N_10360,N_10166);
nor U22063 (N_22063,N_12390,N_15905);
nand U22064 (N_22064,N_16203,N_15854);
xor U22065 (N_22065,N_17261,N_15907);
and U22066 (N_22066,N_17574,N_12447);
nand U22067 (N_22067,N_11379,N_19957);
nor U22068 (N_22068,N_14677,N_15256);
nand U22069 (N_22069,N_12068,N_18664);
nor U22070 (N_22070,N_16933,N_18750);
xor U22071 (N_22071,N_10604,N_16628);
nor U22072 (N_22072,N_10269,N_15143);
nand U22073 (N_22073,N_18491,N_16618);
and U22074 (N_22074,N_14426,N_11451);
or U22075 (N_22075,N_16665,N_16555);
xor U22076 (N_22076,N_19189,N_15939);
nand U22077 (N_22077,N_16380,N_15224);
and U22078 (N_22078,N_10323,N_14606);
or U22079 (N_22079,N_10206,N_15979);
nand U22080 (N_22080,N_17460,N_19541);
nor U22081 (N_22081,N_11927,N_14401);
xnor U22082 (N_22082,N_16561,N_10361);
and U22083 (N_22083,N_15947,N_19496);
nand U22084 (N_22084,N_13395,N_13900);
nand U22085 (N_22085,N_14673,N_12198);
or U22086 (N_22086,N_19625,N_17896);
and U22087 (N_22087,N_18709,N_14578);
and U22088 (N_22088,N_10626,N_11907);
nand U22089 (N_22089,N_11099,N_10162);
and U22090 (N_22090,N_18766,N_16689);
or U22091 (N_22091,N_13497,N_14306);
xnor U22092 (N_22092,N_11815,N_11547);
nor U22093 (N_22093,N_16174,N_11031);
or U22094 (N_22094,N_11895,N_11255);
nand U22095 (N_22095,N_16485,N_10733);
nor U22096 (N_22096,N_13445,N_19777);
and U22097 (N_22097,N_12659,N_15236);
nand U22098 (N_22098,N_14884,N_15696);
or U22099 (N_22099,N_10226,N_12417);
and U22100 (N_22100,N_15813,N_13357);
nor U22101 (N_22101,N_15317,N_12718);
xor U22102 (N_22102,N_18496,N_15218);
xor U22103 (N_22103,N_19083,N_15616);
and U22104 (N_22104,N_11811,N_13444);
nand U22105 (N_22105,N_18166,N_13915);
or U22106 (N_22106,N_16761,N_16627);
nand U22107 (N_22107,N_12383,N_14616);
and U22108 (N_22108,N_15034,N_15390);
nor U22109 (N_22109,N_12163,N_17096);
or U22110 (N_22110,N_16567,N_14196);
and U22111 (N_22111,N_14456,N_12343);
and U22112 (N_22112,N_17461,N_16389);
or U22113 (N_22113,N_15467,N_12647);
nor U22114 (N_22114,N_13319,N_17957);
nand U22115 (N_22115,N_15776,N_19907);
nand U22116 (N_22116,N_13376,N_16890);
or U22117 (N_22117,N_12240,N_11340);
or U22118 (N_22118,N_10319,N_19919);
xnor U22119 (N_22119,N_16405,N_12942);
xnor U22120 (N_22120,N_17596,N_19821);
nand U22121 (N_22121,N_15749,N_17789);
and U22122 (N_22122,N_13024,N_13973);
xnor U22123 (N_22123,N_19838,N_16512);
nand U22124 (N_22124,N_13680,N_15902);
nand U22125 (N_22125,N_11003,N_13504);
nand U22126 (N_22126,N_14628,N_15223);
or U22127 (N_22127,N_18579,N_19339);
or U22128 (N_22128,N_13614,N_16951);
nand U22129 (N_22129,N_13122,N_16283);
and U22130 (N_22130,N_18072,N_18515);
or U22131 (N_22131,N_16646,N_15264);
nor U22132 (N_22132,N_15441,N_11112);
and U22133 (N_22133,N_14966,N_19853);
or U22134 (N_22134,N_11841,N_14309);
xor U22135 (N_22135,N_18570,N_13079);
or U22136 (N_22136,N_19718,N_13510);
and U22137 (N_22137,N_18898,N_17998);
or U22138 (N_22138,N_14329,N_15893);
xnor U22139 (N_22139,N_15262,N_10403);
xnor U22140 (N_22140,N_10088,N_10994);
and U22141 (N_22141,N_11731,N_16944);
or U22142 (N_22142,N_14184,N_19586);
and U22143 (N_22143,N_12926,N_18754);
or U22144 (N_22144,N_19057,N_14827);
xnor U22145 (N_22145,N_16586,N_13187);
and U22146 (N_22146,N_17279,N_12514);
xnor U22147 (N_22147,N_11473,N_12993);
or U22148 (N_22148,N_18539,N_10773);
xor U22149 (N_22149,N_15645,N_17076);
xnor U22150 (N_22150,N_10172,N_19990);
or U22151 (N_22151,N_19789,N_16819);
nor U22152 (N_22152,N_17509,N_16366);
xor U22153 (N_22153,N_11108,N_10044);
xnor U22154 (N_22154,N_19202,N_15445);
and U22155 (N_22155,N_13057,N_17702);
nand U22156 (N_22156,N_12696,N_11306);
xor U22157 (N_22157,N_11770,N_13519);
and U22158 (N_22158,N_13369,N_11904);
or U22159 (N_22159,N_14429,N_10344);
xor U22160 (N_22160,N_19850,N_18981);
xnor U22161 (N_22161,N_13815,N_12815);
and U22162 (N_22162,N_17948,N_14228);
and U22163 (N_22163,N_13982,N_19224);
xor U22164 (N_22164,N_14036,N_16922);
nor U22165 (N_22165,N_15409,N_13364);
xnor U22166 (N_22166,N_14131,N_10388);
xnor U22167 (N_22167,N_16633,N_14799);
or U22168 (N_22168,N_19587,N_13118);
and U22169 (N_22169,N_13414,N_12550);
xor U22170 (N_22170,N_12107,N_10734);
and U22171 (N_22171,N_10830,N_19287);
and U22172 (N_22172,N_10752,N_11325);
or U22173 (N_22173,N_14714,N_10639);
or U22174 (N_22174,N_11844,N_12767);
and U22175 (N_22175,N_16521,N_16311);
or U22176 (N_22176,N_12662,N_18262);
nand U22177 (N_22177,N_12089,N_18451);
and U22178 (N_22178,N_18748,N_16749);
or U22179 (N_22179,N_11089,N_19201);
xor U22180 (N_22180,N_18381,N_13025);
nor U22181 (N_22181,N_13712,N_16462);
and U22182 (N_22182,N_13874,N_13853);
xnor U22183 (N_22183,N_15579,N_19582);
and U22184 (N_22184,N_13515,N_14743);
or U22185 (N_22185,N_19694,N_12313);
and U22186 (N_22186,N_12042,N_19652);
or U22187 (N_22187,N_18249,N_19620);
xor U22188 (N_22188,N_15535,N_10988);
xor U22189 (N_22189,N_17763,N_19302);
and U22190 (N_22190,N_14945,N_15498);
or U22191 (N_22191,N_15097,N_18931);
nand U22192 (N_22192,N_18256,N_12257);
or U22193 (N_22193,N_19645,N_14571);
nor U22194 (N_22194,N_14816,N_18801);
nand U22195 (N_22195,N_18357,N_12829);
nand U22196 (N_22196,N_12141,N_11424);
xnor U22197 (N_22197,N_16532,N_19590);
or U22198 (N_22198,N_18959,N_13339);
xor U22199 (N_22199,N_16542,N_13082);
or U22200 (N_22200,N_16550,N_17774);
and U22201 (N_22201,N_16471,N_16504);
xor U22202 (N_22202,N_18694,N_16818);
and U22203 (N_22203,N_16637,N_17078);
nand U22204 (N_22204,N_15376,N_15203);
or U22205 (N_22205,N_13577,N_14539);
nand U22206 (N_22206,N_17897,N_10769);
and U22207 (N_22207,N_12002,N_12268);
nand U22208 (N_22208,N_17475,N_19519);
or U22209 (N_22209,N_13662,N_17820);
or U22210 (N_22210,N_16491,N_17038);
xnor U22211 (N_22211,N_17317,N_10023);
or U22212 (N_22212,N_10401,N_11750);
xor U22213 (N_22213,N_15797,N_16264);
or U22214 (N_22214,N_14639,N_13210);
nor U22215 (N_22215,N_14409,N_19497);
and U22216 (N_22216,N_14680,N_19900);
or U22217 (N_22217,N_13786,N_11912);
nor U22218 (N_22218,N_19161,N_11843);
or U22219 (N_22219,N_11450,N_15369);
and U22220 (N_22220,N_17085,N_16658);
and U22221 (N_22221,N_15514,N_14647);
and U22222 (N_22222,N_19396,N_11030);
and U22223 (N_22223,N_13613,N_17942);
and U22224 (N_22224,N_18758,N_11360);
nor U22225 (N_22225,N_12809,N_17392);
and U22226 (N_22226,N_11905,N_12642);
and U22227 (N_22227,N_10498,N_19802);
nand U22228 (N_22228,N_19758,N_18601);
and U22229 (N_22229,N_15031,N_10394);
xnor U22230 (N_22230,N_17300,N_15490);
nor U22231 (N_22231,N_19135,N_15998);
and U22232 (N_22232,N_10592,N_16457);
and U22233 (N_22233,N_17525,N_19239);
nor U22234 (N_22234,N_13773,N_13108);
nand U22235 (N_22235,N_12402,N_11570);
and U22236 (N_22236,N_13615,N_14756);
xnor U22237 (N_22237,N_15378,N_16670);
xor U22238 (N_22238,N_19750,N_18844);
nand U22239 (N_22239,N_19960,N_15881);
nand U22240 (N_22240,N_18685,N_11273);
or U22241 (N_22241,N_14611,N_17192);
xor U22242 (N_22242,N_19638,N_19234);
nor U22243 (N_22243,N_16598,N_12946);
nor U22244 (N_22244,N_19571,N_10058);
and U22245 (N_22245,N_11092,N_14180);
and U22246 (N_22246,N_15164,N_16745);
xor U22247 (N_22247,N_10066,N_15157);
xnor U22248 (N_22248,N_16281,N_15774);
nand U22249 (N_22249,N_15290,N_15506);
xor U22250 (N_22250,N_13501,N_10224);
xnor U22251 (N_22251,N_10560,N_14926);
nand U22252 (N_22252,N_10579,N_15798);
xnor U22253 (N_22253,N_14788,N_14453);
or U22254 (N_22254,N_12354,N_15110);
nor U22255 (N_22255,N_18273,N_13495);
xnor U22256 (N_22256,N_14631,N_11890);
nand U22257 (N_22257,N_13972,N_13067);
and U22258 (N_22258,N_18413,N_10656);
and U22259 (N_22259,N_18227,N_18604);
nand U22260 (N_22260,N_19917,N_13784);
xnor U22261 (N_22261,N_11615,N_18805);
nand U22262 (N_22262,N_11300,N_16495);
nand U22263 (N_22263,N_13044,N_12537);
nor U22264 (N_22264,N_10293,N_10695);
or U22265 (N_22265,N_17733,N_14592);
and U22266 (N_22266,N_10069,N_15709);
nand U22267 (N_22267,N_17454,N_14882);
and U22268 (N_22268,N_10979,N_11066);
nand U22269 (N_22269,N_10089,N_19021);
xnor U22270 (N_22270,N_19829,N_17335);
nand U22271 (N_22271,N_13966,N_15209);
nor U22272 (N_22272,N_15012,N_12211);
nor U22273 (N_22273,N_12229,N_15297);
nor U22274 (N_22274,N_16017,N_15602);
xnor U22275 (N_22275,N_11526,N_11184);
and U22276 (N_22276,N_18103,N_12049);
nor U22277 (N_22277,N_13300,N_18887);
or U22278 (N_22278,N_10610,N_10846);
and U22279 (N_22279,N_11862,N_14052);
or U22280 (N_22280,N_12609,N_15339);
nand U22281 (N_22281,N_12439,N_18714);
and U22282 (N_22282,N_19392,N_13152);
or U22283 (N_22283,N_11168,N_15134);
or U22284 (N_22284,N_12336,N_10124);
and U22285 (N_22285,N_17920,N_14051);
or U22286 (N_22286,N_13711,N_16260);
or U22287 (N_22287,N_16993,N_15132);
nand U22288 (N_22288,N_10420,N_16316);
nor U22289 (N_22289,N_14524,N_18205);
xor U22290 (N_22290,N_18724,N_19046);
xor U22291 (N_22291,N_15673,N_19404);
and U22292 (N_22292,N_14269,N_10730);
xnor U22293 (N_22293,N_11435,N_12105);
or U22294 (N_22294,N_15069,N_10918);
or U22295 (N_22295,N_11217,N_14822);
or U22296 (N_22296,N_15226,N_13653);
xnor U22297 (N_22297,N_13944,N_12863);
and U22298 (N_22298,N_14399,N_11086);
or U22299 (N_22299,N_15367,N_16934);
nor U22300 (N_22300,N_12499,N_18618);
and U22301 (N_22301,N_13114,N_19766);
xor U22302 (N_22302,N_12793,N_17983);
nor U22303 (N_22303,N_10699,N_16925);
nor U22304 (N_22304,N_17479,N_12649);
nor U22305 (N_22305,N_19749,N_11467);
and U22306 (N_22306,N_12073,N_15272);
xnor U22307 (N_22307,N_12193,N_13059);
nor U22308 (N_22308,N_11279,N_13076);
nand U22309 (N_22309,N_14527,N_15866);
or U22310 (N_22310,N_17671,N_12004);
nor U22311 (N_22311,N_10700,N_16649);
nor U22312 (N_22312,N_18332,N_12225);
xnor U22313 (N_22313,N_10240,N_19575);
and U22314 (N_22314,N_16005,N_18333);
and U22315 (N_22315,N_13323,N_14864);
or U22316 (N_22316,N_12035,N_10878);
or U22317 (N_22317,N_14970,N_10423);
nor U22318 (N_22318,N_10397,N_11817);
or U22319 (N_22319,N_13756,N_12475);
and U22320 (N_22320,N_15418,N_10428);
nand U22321 (N_22321,N_19395,N_14506);
xnor U22322 (N_22322,N_14012,N_12676);
nand U22323 (N_22323,N_14120,N_14094);
xor U22324 (N_22324,N_13654,N_16349);
or U22325 (N_22325,N_18025,N_17595);
or U22326 (N_22326,N_12093,N_19518);
nand U22327 (N_22327,N_15717,N_15239);
nand U22328 (N_22328,N_18020,N_19458);
nor U22329 (N_22329,N_18087,N_18567);
or U22330 (N_22330,N_19778,N_18688);
nor U22331 (N_22331,N_15085,N_13128);
or U22332 (N_22332,N_13552,N_11977);
xor U22333 (N_22333,N_19307,N_12116);
and U22334 (N_22334,N_12905,N_12190);
xnor U22335 (N_22335,N_11694,N_19150);
nor U22336 (N_22336,N_11372,N_10126);
nor U22337 (N_22337,N_14114,N_17125);
and U22338 (N_22338,N_11673,N_19623);
or U22339 (N_22339,N_19751,N_18804);
or U22340 (N_22340,N_13481,N_11075);
nand U22341 (N_22341,N_19559,N_13279);
nor U22342 (N_22342,N_10716,N_13650);
or U22343 (N_22343,N_16476,N_12168);
nor U22344 (N_22344,N_15438,N_15379);
nand U22345 (N_22345,N_17278,N_15013);
or U22346 (N_22346,N_14158,N_13771);
or U22347 (N_22347,N_12772,N_11391);
or U22348 (N_22348,N_15727,N_11928);
nor U22349 (N_22349,N_11657,N_19745);
nand U22350 (N_22350,N_17435,N_17989);
nor U22351 (N_22351,N_16387,N_13605);
nor U22352 (N_22352,N_18034,N_11749);
nand U22353 (N_22353,N_11715,N_13375);
xnor U22354 (N_22354,N_18552,N_13600);
xnor U22355 (N_22355,N_19691,N_15231);
nor U22356 (N_22356,N_16884,N_15489);
nor U22357 (N_22357,N_16332,N_10006);
xnor U22358 (N_22358,N_19508,N_12631);
nand U22359 (N_22359,N_15055,N_17934);
or U22360 (N_22360,N_14390,N_18468);
nor U22361 (N_22361,N_18767,N_19427);
nand U22362 (N_22362,N_10287,N_19499);
and U22363 (N_22363,N_15469,N_15313);
or U22364 (N_22364,N_12935,N_19693);
nand U22365 (N_22365,N_10986,N_13536);
and U22366 (N_22366,N_11292,N_11263);
xnor U22367 (N_22367,N_16056,N_15188);
or U22368 (N_22368,N_10962,N_15916);
nand U22369 (N_22369,N_19417,N_10767);
and U22370 (N_22370,N_18746,N_14939);
xnor U22371 (N_22371,N_15792,N_12600);
and U22372 (N_22372,N_19851,N_15296);
and U22373 (N_22373,N_11620,N_12199);
and U22374 (N_22374,N_10980,N_17272);
nor U22375 (N_22375,N_11042,N_11855);
xor U22376 (N_22376,N_10183,N_17924);
and U22377 (N_22377,N_17015,N_16617);
and U22378 (N_22378,N_12572,N_17445);
nand U22379 (N_22379,N_14355,N_19240);
nor U22380 (N_22380,N_18054,N_12547);
nor U22381 (N_22381,N_15834,N_13585);
nand U22382 (N_22382,N_14784,N_11226);
and U22383 (N_22383,N_10249,N_19463);
nor U22384 (N_22384,N_17773,N_19062);
and U22385 (N_22385,N_18810,N_11466);
and U22386 (N_22386,N_13214,N_15258);
nor U22387 (N_22387,N_15370,N_18573);
nand U22388 (N_22388,N_11836,N_16971);
nand U22389 (N_22389,N_13643,N_19724);
or U22390 (N_22390,N_13717,N_18510);
nor U22391 (N_22391,N_16754,N_18993);
or U22392 (N_22392,N_13204,N_11458);
nand U22393 (N_22393,N_15906,N_17737);
nor U22394 (N_22394,N_18178,N_18782);
nor U22395 (N_22395,N_18115,N_16986);
and U22396 (N_22396,N_10616,N_10815);
and U22397 (N_22397,N_17822,N_18673);
nor U22398 (N_22398,N_15494,N_15117);
nand U22399 (N_22399,N_19028,N_19377);
nand U22400 (N_22400,N_11010,N_14098);
and U22401 (N_22401,N_19512,N_17216);
and U22402 (N_22402,N_19996,N_17056);
xor U22403 (N_22403,N_10017,N_13124);
or U22404 (N_22404,N_16908,N_12791);
xor U22405 (N_22405,N_17100,N_14129);
nand U22406 (N_22406,N_10696,N_11946);
and U22407 (N_22407,N_16290,N_14568);
or U22408 (N_22408,N_18854,N_18847);
nor U22409 (N_22409,N_17336,N_19013);
or U22410 (N_22410,N_14748,N_16158);
nand U22411 (N_22411,N_14761,N_14697);
nand U22412 (N_22412,N_16505,N_16939);
nand U22413 (N_22413,N_17094,N_12086);
nand U22414 (N_22414,N_14549,N_10251);
and U22415 (N_22415,N_17625,N_14115);
and U22416 (N_22416,N_14545,N_12908);
xor U22417 (N_22417,N_12933,N_16734);
and U22418 (N_22418,N_15271,N_10264);
nor U22419 (N_22419,N_19133,N_18740);
nor U22420 (N_22420,N_16515,N_19819);
and U22421 (N_22421,N_16800,N_13227);
or U22422 (N_22422,N_12740,N_17024);
and U22423 (N_22423,N_19514,N_19504);
nor U22424 (N_22424,N_13439,N_12590);
xnor U22425 (N_22425,N_14496,N_10351);
or U22426 (N_22426,N_18168,N_18105);
or U22427 (N_22427,N_18068,N_11268);
xor U22428 (N_22428,N_14627,N_17432);
and U22429 (N_22429,N_11500,N_14461);
or U22430 (N_22430,N_13155,N_18530);
nand U22431 (N_22431,N_12774,N_17516);
or U22432 (N_22432,N_10410,N_10644);
and U22433 (N_22433,N_19277,N_19932);
nand U22434 (N_22434,N_16632,N_18309);
or U22435 (N_22435,N_11422,N_17474);
xor U22436 (N_22436,N_16748,N_17726);
xnor U22437 (N_22437,N_19093,N_11425);
or U22438 (N_22438,N_11037,N_15799);
and U22439 (N_22439,N_13050,N_15840);
and U22440 (N_22440,N_17360,N_12081);
xnor U22441 (N_22441,N_17668,N_11901);
or U22442 (N_22442,N_14789,N_11585);
nor U22443 (N_22443,N_14678,N_17836);
nand U22444 (N_22444,N_18708,N_19361);
or U22445 (N_22445,N_18752,N_16912);
nand U22446 (N_22446,N_15030,N_15931);
nor U22447 (N_22447,N_10123,N_15726);
or U22448 (N_22448,N_11062,N_11746);
nand U22449 (N_22449,N_10220,N_14747);
and U22450 (N_22450,N_15447,N_18240);
xor U22451 (N_22451,N_19689,N_11857);
and U22452 (N_22452,N_11885,N_14618);
nor U22453 (N_22453,N_19852,N_13511);
nand U22454 (N_22454,N_12391,N_13335);
nor U22455 (N_22455,N_14063,N_19414);
nand U22456 (N_22456,N_10202,N_15077);
xor U22457 (N_22457,N_15048,N_11819);
nor U22458 (N_22458,N_17242,N_13042);
nor U22459 (N_22459,N_17481,N_17385);
nor U22460 (N_22460,N_18376,N_12096);
and U22461 (N_22461,N_18787,N_17260);
xor U22462 (N_22462,N_13030,N_13138);
and U22463 (N_22463,N_17833,N_18680);
nor U22464 (N_22464,N_14965,N_16450);
nand U22465 (N_22465,N_12453,N_17036);
or U22466 (N_22466,N_10030,N_13419);
or U22467 (N_22467,N_18175,N_10595);
and U22468 (N_22468,N_14137,N_13988);
and U22469 (N_22469,N_19534,N_16891);
xnor U22470 (N_22470,N_11021,N_18778);
and U22471 (N_22471,N_16423,N_13796);
nand U22472 (N_22472,N_10811,N_13010);
or U22473 (N_22473,N_16420,N_19583);
and U22474 (N_22474,N_17027,N_13755);
nand U22475 (N_22475,N_13733,N_14929);
and U22476 (N_22476,N_18061,N_15491);
nor U22477 (N_22477,N_16878,N_19371);
nor U22478 (N_22478,N_18472,N_10372);
and U22479 (N_22479,N_16105,N_18830);
nand U22480 (N_22480,N_19430,N_12209);
and U22481 (N_22481,N_12652,N_10290);
nand U22482 (N_22482,N_14666,N_11758);
xnor U22483 (N_22483,N_12857,N_15634);
nand U22484 (N_22484,N_13311,N_12195);
nand U22485 (N_22485,N_18818,N_13134);
nand U22486 (N_22486,N_15711,N_15874);
or U22487 (N_22487,N_16152,N_10157);
nor U22488 (N_22488,N_13436,N_15836);
nor U22489 (N_22489,N_15870,N_17064);
xor U22490 (N_22490,N_11605,N_14912);
nand U22491 (N_22491,N_17885,N_13188);
and U22492 (N_22492,N_14366,N_12843);
xnor U22493 (N_22493,N_16705,N_17316);
nor U22494 (N_22494,N_10115,N_18706);
and U22495 (N_22495,N_12256,N_10963);
nand U22496 (N_22496,N_15109,N_19471);
nor U22497 (N_22497,N_19411,N_16693);
nand U22498 (N_22498,N_12167,N_12378);
xnor U22499 (N_22499,N_16808,N_18260);
and U22500 (N_22500,N_18535,N_14183);
xor U22501 (N_22501,N_14344,N_18041);
or U22502 (N_22502,N_19931,N_16905);
or U22503 (N_22503,N_18842,N_13412);
xor U22504 (N_22504,N_10778,N_19255);
xor U22505 (N_22505,N_15285,N_17229);
or U22506 (N_22506,N_16128,N_12208);
and U22507 (N_22507,N_16433,N_16108);
and U22508 (N_22508,N_16851,N_19055);
or U22509 (N_22509,N_11049,N_16506);
or U22510 (N_22510,N_10634,N_11540);
nand U22511 (N_22511,N_18862,N_18160);
nor U22512 (N_22512,N_14890,N_12811);
or U22513 (N_22513,N_15346,N_13151);
nor U22514 (N_22514,N_13285,N_14233);
nand U22515 (N_22515,N_12492,N_12721);
or U22516 (N_22516,N_14908,N_10611);
nor U22517 (N_22517,N_17084,N_18903);
or U22518 (N_22518,N_13690,N_13508);
nand U22519 (N_22519,N_12517,N_15404);
nor U22520 (N_22520,N_17017,N_15853);
nor U22521 (N_22521,N_11565,N_14994);
and U22522 (N_22522,N_10549,N_13513);
xor U22523 (N_22523,N_11353,N_15160);
xor U22524 (N_22524,N_15257,N_16732);
xnor U22525 (N_22525,N_13665,N_14739);
or U22526 (N_22526,N_14397,N_19431);
nand U22527 (N_22527,N_17705,N_19490);
nor U22528 (N_22528,N_11222,N_13388);
and U22529 (N_22529,N_14138,N_14985);
nor U22530 (N_22530,N_13873,N_15593);
or U22531 (N_22531,N_18944,N_17591);
xnor U22532 (N_22532,N_18629,N_19967);
nor U22533 (N_22533,N_17520,N_15395);
nand U22534 (N_22534,N_11264,N_13367);
or U22535 (N_22535,N_12750,N_18525);
nand U22536 (N_22536,N_15559,N_17420);
nor U22537 (N_22537,N_16155,N_16244);
nor U22538 (N_22538,N_10779,N_10409);
nand U22539 (N_22539,N_17921,N_18721);
xnor U22540 (N_22540,N_11985,N_10851);
xor U22541 (N_22541,N_17649,N_10676);
and U22542 (N_22542,N_12867,N_12975);
nand U22543 (N_22543,N_14007,N_12927);
nand U22544 (N_22544,N_19242,N_19696);
nand U22545 (N_22545,N_18173,N_12974);
nor U22546 (N_22546,N_13321,N_14111);
xnor U22547 (N_22547,N_11820,N_18370);
nor U22548 (N_22548,N_15216,N_16554);
and U22549 (N_22549,N_14978,N_18036);
nor U22550 (N_22550,N_11916,N_17029);
nand U22551 (N_22551,N_11581,N_16823);
xor U22552 (N_22552,N_16455,N_10740);
or U22553 (N_22553,N_19237,N_14701);
and U22554 (N_22554,N_10248,N_16237);
nor U22555 (N_22555,N_17021,N_13957);
and U22556 (N_22556,N_13724,N_19233);
nand U22557 (N_22557,N_11018,N_11327);
or U22558 (N_22558,N_11494,N_10776);
nand U22559 (N_22559,N_19922,N_11434);
and U22560 (N_22560,N_10232,N_15270);
nand U22561 (N_22561,N_17814,N_14234);
nand U22562 (N_22562,N_11892,N_14974);
nand U22563 (N_22563,N_16210,N_13689);
nor U22564 (N_22564,N_18346,N_12667);
and U22565 (N_22565,N_15761,N_12948);
xor U22566 (N_22566,N_12726,N_18352);
and U22567 (N_22567,N_15331,N_15641);
nand U22568 (N_22568,N_19473,N_16965);
nand U22569 (N_22569,N_15991,N_12021);
and U22570 (N_22570,N_11631,N_18222);
or U22571 (N_22571,N_10271,N_18279);
nor U22572 (N_22572,N_19669,N_14447);
or U22573 (N_22573,N_11772,N_13750);
and U22574 (N_22574,N_10806,N_10586);
nor U22575 (N_22575,N_10601,N_13396);
nor U22576 (N_22576,N_17383,N_19353);
nand U22577 (N_22577,N_15744,N_12769);
nor U22578 (N_22578,N_10680,N_13721);
nor U22579 (N_22579,N_12224,N_18665);
or U22580 (N_22580,N_15278,N_18465);
and U22581 (N_22581,N_11561,N_13229);
and U22582 (N_22582,N_10788,N_16829);
nor U22583 (N_22583,N_15783,N_18002);
and U22584 (N_22584,N_14149,N_12341);
nand U22585 (N_22585,N_18003,N_18689);
xnor U22586 (N_22586,N_10252,N_17181);
xor U22587 (N_22587,N_16695,N_18684);
nand U22588 (N_22588,N_19756,N_12149);
nand U22589 (N_22589,N_10438,N_18378);
or U22590 (N_22590,N_14280,N_12957);
and U22591 (N_22591,N_14526,N_17624);
xor U22592 (N_22592,N_11685,N_10445);
or U22593 (N_22593,N_15245,N_19437);
xor U22594 (N_22594,N_15808,N_17657);
nor U22595 (N_22595,N_13407,N_16235);
and U22596 (N_22596,N_11883,N_12969);
or U22597 (N_22597,N_12520,N_12934);
nor U22598 (N_22598,N_15617,N_12950);
nor U22599 (N_22599,N_10122,N_11995);
or U22600 (N_22600,N_11902,N_13405);
xnor U22601 (N_22601,N_18935,N_16539);
or U22602 (N_22602,N_17095,N_19985);
nand U22603 (N_22603,N_11320,N_10563);
or U22604 (N_22604,N_19151,N_19379);
nand U22605 (N_22605,N_16215,N_13632);
or U22606 (N_22606,N_15324,N_18083);
xnor U22607 (N_22607,N_16123,N_13872);
or U22608 (N_22608,N_14901,N_14124);
and U22609 (N_22609,N_17868,N_19700);
or U22610 (N_22610,N_10452,N_11478);
and U22611 (N_22611,N_11838,N_16289);
nor U22612 (N_22612,N_15411,N_11509);
xnor U22613 (N_22613,N_16777,N_17201);
and U22614 (N_22614,N_19346,N_11371);
xor U22615 (N_22615,N_17277,N_18558);
xnor U22616 (N_22616,N_13101,N_15001);
xnor U22617 (N_22617,N_15009,N_17884);
or U22618 (N_22618,N_10689,N_13696);
nand U22619 (N_22619,N_11201,N_13119);
and U22620 (N_22620,N_15789,N_12979);
xor U22621 (N_22621,N_15587,N_10079);
xor U22622 (N_22622,N_18319,N_14532);
and U22623 (N_22623,N_10624,N_10133);
nor U22624 (N_22624,N_14495,N_10543);
nand U22625 (N_22625,N_19311,N_16162);
and U22626 (N_22626,N_19911,N_10713);
nor U22627 (N_22627,N_17108,N_11937);
and U22628 (N_22628,N_19182,N_14593);
or U22629 (N_22629,N_16407,N_12292);
xor U22630 (N_22630,N_10520,N_13429);
or U22631 (N_22631,N_10556,N_12020);
nor U22632 (N_22632,N_19156,N_10143);
and U22633 (N_22633,N_10065,N_19920);
nand U22634 (N_22634,N_13381,N_19597);
nand U22635 (N_22635,N_18952,N_14832);
xor U22636 (N_22636,N_14916,N_15780);
or U22637 (N_22637,N_13971,N_12575);
or U22638 (N_22638,N_13660,N_17170);
xor U22639 (N_22639,N_14662,N_17874);
nand U22640 (N_22640,N_15431,N_11369);
or U22641 (N_22641,N_13923,N_19893);
xor U22642 (N_22642,N_15145,N_18942);
nor U22643 (N_22643,N_12428,N_17984);
nor U22644 (N_22644,N_16441,N_10640);
nand U22645 (N_22645,N_15387,N_10475);
nor U22646 (N_22646,N_15294,N_18753);
and U22647 (N_22647,N_18517,N_12804);
or U22648 (N_22648,N_17600,N_17419);
or U22649 (N_22649,N_13999,N_11574);
xnor U22650 (N_22650,N_12512,N_10217);
xor U22651 (N_22651,N_16336,N_14637);
and U22652 (N_22652,N_10375,N_12608);
or U22653 (N_22653,N_11137,N_12101);
xor U22654 (N_22654,N_12132,N_17734);
and U22655 (N_22655,N_16619,N_14041);
nor U22656 (N_22656,N_14480,N_15755);
or U22657 (N_22657,N_13795,N_16321);
or U22658 (N_22658,N_17091,N_18663);
xnor U22659 (N_22659,N_13527,N_16850);
and U22660 (N_22660,N_10154,N_16081);
nand U22661 (N_22661,N_16520,N_15609);
xnor U22662 (N_22662,N_12451,N_15064);
xor U22663 (N_22663,N_13242,N_19214);
xnor U22664 (N_22664,N_11908,N_18913);
nor U22665 (N_22665,N_19565,N_10468);
nand U22666 (N_22666,N_19564,N_17072);
xor U22667 (N_22667,N_15222,N_16285);
xor U22668 (N_22668,N_13570,N_19855);
and U22669 (N_22669,N_14464,N_13235);
nand U22670 (N_22670,N_16378,N_13345);
nand U22671 (N_22671,N_13233,N_14439);
or U22672 (N_22672,N_11415,N_15186);
nor U22673 (N_22673,N_16004,N_19080);
nor U22674 (N_22674,N_19599,N_14612);
or U22675 (N_22675,N_11627,N_15289);
xor U22676 (N_22676,N_18001,N_18545);
or U22677 (N_22677,N_14696,N_19805);
nand U22678 (N_22678,N_11293,N_13371);
nand U22679 (N_22679,N_11139,N_10526);
or U22680 (N_22680,N_16212,N_12568);
and U22681 (N_22681,N_18158,N_11794);
or U22682 (N_22682,N_11305,N_18263);
xor U22683 (N_22683,N_19131,N_14621);
nor U22684 (N_22684,N_19520,N_16432);
or U22685 (N_22685,N_10581,N_15672);
xor U22686 (N_22686,N_18994,N_14699);
and U22687 (N_22687,N_10605,N_10906);
and U22688 (N_22688,N_12247,N_12849);
nand U22689 (N_22689,N_17887,N_16406);
nor U22690 (N_22690,N_18832,N_17172);
and U22691 (N_22691,N_18433,N_14871);
nor U22692 (N_22692,N_11972,N_18607);
nand U22693 (N_22693,N_19660,N_15667);
and U22694 (N_22694,N_13867,N_17902);
and U22695 (N_22695,N_11134,N_11074);
nor U22696 (N_22696,N_16018,N_16054);
nand U22697 (N_22697,N_12670,N_15995);
or U22698 (N_22698,N_12261,N_17688);
or U22699 (N_22699,N_12707,N_12342);
or U22700 (N_22700,N_19011,N_18028);
or U22701 (N_22701,N_10129,N_19624);
or U22702 (N_22702,N_18219,N_10651);
nand U22703 (N_22703,N_15343,N_11559);
nor U22704 (N_22704,N_18008,N_17597);
nor U22705 (N_22705,N_14192,N_16673);
nor U22706 (N_22706,N_15505,N_11207);
xor U22707 (N_22707,N_11156,N_14331);
nand U22708 (N_22708,N_12794,N_16474);
or U22709 (N_22709,N_17508,N_12958);
xor U22710 (N_22710,N_16799,N_13177);
nor U22711 (N_22711,N_19709,N_19314);
xnor U22712 (N_22712,N_16569,N_15195);
nand U22713 (N_22713,N_16866,N_12445);
nand U22714 (N_22714,N_14145,N_17869);
xor U22715 (N_22715,N_13093,N_10949);
nor U22716 (N_22716,N_17666,N_10868);
nand U22717 (N_22717,N_19410,N_16991);
xnor U22718 (N_22718,N_13825,N_18261);
nand U22719 (N_22719,N_18985,N_17457);
nor U22720 (N_22720,N_15038,N_16294);
nor U22721 (N_22721,N_18388,N_16892);
xor U22722 (N_22722,N_18686,N_15266);
or U22723 (N_22723,N_17673,N_18520);
or U22724 (N_22724,N_19776,N_14653);
nor U22725 (N_22725,N_13516,N_11241);
nand U22726 (N_22726,N_13184,N_12801);
nand U22727 (N_22727,N_19010,N_10116);
and U22728 (N_22728,N_11111,N_10682);
and U22729 (N_22729,N_13085,N_18374);
or U22730 (N_22730,N_19704,N_15914);
nand U22731 (N_22731,N_12807,N_17506);
nand U22732 (N_22732,N_10973,N_18086);
nor U22733 (N_22733,N_13413,N_19686);
nor U22734 (N_22734,N_17097,N_14896);
or U22735 (N_22735,N_11783,N_10668);
nor U22736 (N_22736,N_17488,N_11984);
nand U22737 (N_22737,N_11179,N_13239);
xnor U22738 (N_22738,N_11947,N_14437);
nand U22739 (N_22739,N_18733,N_17007);
or U22740 (N_22740,N_13649,N_19760);
nor U22741 (N_22741,N_10690,N_16422);
xnor U22742 (N_22742,N_13793,N_15175);
nand U22743 (N_22743,N_16676,N_19574);
nor U22744 (N_22744,N_19073,N_13832);
or U22745 (N_22745,N_18938,N_16347);
or U22746 (N_22746,N_18170,N_15630);
or U22747 (N_22747,N_15596,N_17994);
or U22748 (N_22748,N_16315,N_14207);
nand U22749 (N_22749,N_16250,N_15821);
nand U22750 (N_22750,N_13888,N_10666);
and U22751 (N_22751,N_16593,N_16544);
nand U22752 (N_22752,N_10223,N_13301);
nor U22753 (N_22753,N_10583,N_14179);
or U22754 (N_22754,N_16629,N_16894);
or U22755 (N_22755,N_12994,N_19611);
nor U22756 (N_22756,N_15137,N_13211);
and U22757 (N_22757,N_15758,N_13794);
nand U22758 (N_22758,N_10822,N_16182);
and U22759 (N_22759,N_17728,N_17721);
or U22760 (N_22760,N_13930,N_10000);
or U22761 (N_22761,N_18489,N_16709);
nor U22762 (N_22762,N_13780,N_18139);
or U22763 (N_22763,N_13840,N_19140);
nor U22764 (N_22764,N_11433,N_10870);
xnor U22765 (N_22765,N_13127,N_16813);
nor U22766 (N_22766,N_12327,N_10389);
or U22767 (N_22767,N_13033,N_13916);
xor U22768 (N_22768,N_16488,N_13854);
and U22769 (N_22769,N_14842,N_16582);
nor U22770 (N_22770,N_16551,N_14139);
and U22771 (N_22771,N_11059,N_12340);
nand U22772 (N_22772,N_17293,N_14844);
nand U22773 (N_22773,N_13581,N_17079);
xnor U22774 (N_22774,N_17012,N_10303);
or U22775 (N_22775,N_15682,N_13337);
or U22776 (N_22776,N_17910,N_13267);
nor U22777 (N_22777,N_18894,N_12841);
xor U22778 (N_22778,N_19943,N_17291);
or U22779 (N_22779,N_13149,N_12449);
or U22780 (N_22780,N_16963,N_12029);
or U22781 (N_22781,N_19894,N_13106);
or U22782 (N_22782,N_10518,N_14323);
xnor U22783 (N_22783,N_18331,N_16010);
or U22784 (N_22784,N_17913,N_11556);
xor U22785 (N_22785,N_14540,N_13738);
xor U22786 (N_22786,N_16014,N_13148);
nor U22787 (N_22787,N_15433,N_16068);
nor U22788 (N_22788,N_12166,N_18305);
xnor U22789 (N_22789,N_19720,N_17161);
and U22790 (N_22790,N_14176,N_18050);
and U22791 (N_22791,N_12273,N_12210);
nand U22792 (N_22792,N_12295,N_16990);
and U22793 (N_22793,N_10169,N_18322);
and U22794 (N_22794,N_10305,N_19475);
nand U22795 (N_22795,N_19291,N_16654);
or U22796 (N_22796,N_16303,N_12715);
nand U22797 (N_22797,N_16727,N_15961);
nor U22798 (N_22798,N_16791,N_15926);
nor U22799 (N_22799,N_17259,N_11566);
or U22800 (N_22800,N_11475,N_10336);
and U22801 (N_22801,N_15398,N_10491);
and U22802 (N_22802,N_10920,N_14502);
nand U22803 (N_22803,N_12012,N_16522);
and U22804 (N_22804,N_12123,N_11945);
xor U22805 (N_22805,N_12119,N_15592);
xnor U22806 (N_22806,N_16697,N_14065);
and U22807 (N_22807,N_16436,N_17232);
or U22808 (N_22808,N_15908,N_12816);
or U22809 (N_22809,N_18979,N_19423);
nand U22810 (N_22810,N_15927,N_11988);
and U22811 (N_22811,N_15771,N_14476);
and U22812 (N_22812,N_12278,N_15841);
and U22813 (N_22813,N_14156,N_13173);
nor U22814 (N_22814,N_18653,N_16615);
xor U22815 (N_22815,N_15247,N_18498);
nand U22816 (N_22816,N_10446,N_11624);
or U22817 (N_22817,N_10127,N_11395);
xnor U22818 (N_22818,N_18232,N_17240);
nand U22819 (N_22819,N_15886,N_12523);
nor U22820 (N_22820,N_13225,N_17919);
and U22821 (N_22821,N_12712,N_17510);
or U22822 (N_22822,N_12596,N_17459);
nand U22823 (N_22823,N_13102,N_12853);
and U22824 (N_22824,N_14316,N_18775);
or U22825 (N_22825,N_10107,N_19203);
nand U22826 (N_22826,N_14874,N_16197);
xnor U22827 (N_22827,N_13626,N_12039);
and U22828 (N_22828,N_18777,N_17126);
nand U22829 (N_22829,N_11274,N_10411);
nor U22830 (N_22830,N_18945,N_13021);
or U22831 (N_22831,N_18212,N_19616);
nor U22832 (N_22832,N_19249,N_19801);
nor U22833 (N_22833,N_17374,N_17490);
and U22834 (N_22834,N_11180,N_16121);
nand U22835 (N_22835,N_15182,N_17171);
nand U22836 (N_22836,N_19966,N_18391);
xnor U22837 (N_22837,N_13350,N_15293);
and U22838 (N_22838,N_15096,N_16050);
xnor U22839 (N_22839,N_15397,N_18603);
nand U22840 (N_22840,N_13342,N_10215);
nand U22841 (N_22841,N_12036,N_13199);
or U22842 (N_22842,N_12057,N_19610);
or U22843 (N_22843,N_11228,N_14010);
nor U22844 (N_22844,N_12469,N_18912);
nor U22845 (N_22845,N_13587,N_12582);
xnor U22846 (N_22846,N_18988,N_16460);
or U22847 (N_22847,N_11640,N_17709);
nor U22848 (N_22848,N_17256,N_12817);
and U22849 (N_22849,N_15019,N_15942);
or U22850 (N_22850,N_19874,N_14781);
or U22851 (N_22851,N_12689,N_15847);
xor U22852 (N_22852,N_15729,N_12005);
nor U22853 (N_22853,N_16356,N_11384);
or U22854 (N_22854,N_14625,N_12465);
and U22855 (N_22855,N_12164,N_18838);
nor U22856 (N_22856,N_19524,N_14950);
or U22857 (N_22857,N_14763,N_12570);
nor U22858 (N_22858,N_15652,N_12787);
nand U22859 (N_22859,N_11414,N_13896);
nor U22860 (N_22860,N_17795,N_17168);
xor U22861 (N_22861,N_14940,N_15542);
or U22862 (N_22862,N_11284,N_10221);
nand U22863 (N_22863,N_16909,N_13740);
nor U22864 (N_22864,N_18799,N_12858);
and U22865 (N_22865,N_13672,N_15871);
nand U22866 (N_22866,N_14683,N_18662);
or U22867 (N_22867,N_13243,N_16788);
nand U22868 (N_22868,N_16494,N_18286);
nor U22869 (N_22869,N_10774,N_17568);
nor U22870 (N_22870,N_12552,N_16413);
nand U22871 (N_22871,N_16124,N_10506);
or U22872 (N_22872,N_17542,N_19398);
and U22873 (N_22873,N_13474,N_14858);
or U22874 (N_22874,N_14441,N_10932);
xor U22875 (N_22875,N_11454,N_16065);
xor U22876 (N_22876,N_18918,N_13747);
and U22877 (N_22877,N_14424,N_16168);
nand U22878 (N_22878,N_10083,N_13248);
nor U22879 (N_22879,N_15863,N_15332);
or U22880 (N_22880,N_15391,N_15775);
xor U22881 (N_22881,N_17693,N_12531);
and U22882 (N_22882,N_17923,N_16287);
nor U22883 (N_22883,N_14640,N_14786);
and U22884 (N_22884,N_10159,N_10246);
nor U22885 (N_22885,N_13627,N_11753);
nand U22886 (N_22886,N_16127,N_12462);
xnor U22887 (N_22887,N_18056,N_12674);
nor U22888 (N_22888,N_11833,N_14690);
and U22889 (N_22889,N_14776,N_19366);
or U22890 (N_22890,N_19100,N_12892);
nand U22891 (N_22891,N_12795,N_11389);
or U22892 (N_22892,N_11822,N_11553);
or U22893 (N_22893,N_15511,N_17303);
or U22894 (N_22894,N_15123,N_13208);
and U22895 (N_22895,N_17339,N_13282);
nor U22896 (N_22896,N_14167,N_18268);
or U22897 (N_22897,N_16044,N_13309);
nor U22898 (N_22898,N_15827,N_16508);
or U22899 (N_22899,N_11368,N_16288);
nor U22900 (N_22900,N_15952,N_10233);
or U22901 (N_22901,N_10965,N_10497);
nand U22902 (N_22902,N_14825,N_12124);
nor U22903 (N_22903,N_18235,N_16141);
and U22904 (N_22904,N_10103,N_19368);
nor U22905 (N_22905,N_18004,N_11212);
xnor U22906 (N_22906,N_14651,N_19820);
or U22907 (N_22907,N_16841,N_10981);
nand U22908 (N_22908,N_14194,N_18895);
xnor U22909 (N_22909,N_11045,N_19857);
and U22910 (N_22910,N_13772,N_10395);
and U22911 (N_22911,N_17467,N_11121);
xor U22912 (N_22912,N_10163,N_19786);
and U22913 (N_22913,N_13956,N_18660);
and U22914 (N_22914,N_17962,N_19139);
xor U22915 (N_22915,N_19699,N_10620);
nand U22916 (N_22916,N_11157,N_13686);
xnor U22917 (N_22917,N_11853,N_10228);
nand U22918 (N_22918,N_18117,N_10623);
and U22919 (N_22919,N_17537,N_18176);
and U22920 (N_22920,N_10036,N_11719);
nand U22921 (N_22921,N_11965,N_18133);
nor U22922 (N_22922,N_16243,N_10168);
or U22923 (N_22923,N_10052,N_12828);
nand U22924 (N_22924,N_19022,N_16502);
nor U22925 (N_22925,N_19673,N_19464);
xnor U22926 (N_22926,N_13047,N_15220);
nand U22927 (N_22927,N_15416,N_13043);
nand U22928 (N_22928,N_12636,N_18586);
nand U22929 (N_22929,N_10911,N_17939);
or U22930 (N_22930,N_17830,N_16229);
and U22931 (N_22931,N_12339,N_11861);
nor U22932 (N_22932,N_10941,N_16664);
and U22933 (N_22933,N_14935,N_18783);
xor U22934 (N_22934,N_12522,N_19413);
and U22935 (N_22935,N_11213,N_15179);
and U22936 (N_22936,N_12456,N_10262);
xnor U22937 (N_22937,N_18055,N_10256);
nor U22938 (N_22938,N_11970,N_16341);
or U22939 (N_22939,N_10535,N_18386);
xnor U22940 (N_22940,N_14620,N_17742);
or U22941 (N_22941,N_11170,N_13610);
and U22942 (N_22942,N_11590,N_12182);
nor U22943 (N_22943,N_15920,N_13378);
nor U22944 (N_22944,N_10867,N_16180);
xnor U22945 (N_22945,N_19419,N_12951);
nor U22946 (N_22946,N_18165,N_13783);
nand U22947 (N_22947,N_15540,N_15818);
nand U22948 (N_22948,N_14692,N_19890);
nand U22949 (N_22949,N_19476,N_16771);
nor U22950 (N_22950,N_16239,N_10517);
nor U22951 (N_22951,N_11221,N_19109);
and U22952 (N_22952,N_16932,N_17437);
or U22953 (N_22953,N_12851,N_13707);
nor U22954 (N_22954,N_19218,N_12461);
or U22955 (N_22955,N_19649,N_15388);
xor U22956 (N_22956,N_13878,N_19370);
nand U22957 (N_22957,N_17389,N_16548);
and U22958 (N_22958,N_14787,N_13912);
nor U22959 (N_22959,N_16901,N_13628);
or U22960 (N_22960,N_19002,N_12213);
xnor U22961 (N_22961,N_17521,N_16189);
xor U22962 (N_22962,N_16000,N_12175);
nand U22963 (N_22963,N_15426,N_17499);
nand U22964 (N_22964,N_18678,N_18917);
xor U22965 (N_22965,N_11077,N_13075);
and U22966 (N_22966,N_19692,N_18190);
or U22967 (N_22967,N_10161,N_14023);
or U22968 (N_22968,N_15183,N_15020);
and U22969 (N_22969,N_15623,N_16297);
or U22970 (N_22970,N_18474,N_15589);
and U22971 (N_22971,N_13742,N_11245);
or U22972 (N_22972,N_19075,N_18095);
or U22973 (N_22973,N_19088,N_15452);
or U22974 (N_22974,N_15930,N_17831);
or U22975 (N_22975,N_14726,N_19859);
nor U22976 (N_22976,N_11465,N_15102);
and U22977 (N_22977,N_12034,N_17054);
nor U22978 (N_22978,N_10326,N_16659);
nand U22979 (N_22979,N_18395,N_18501);
or U22980 (N_22980,N_16996,N_10528);
or U22981 (N_22981,N_19685,N_11124);
xnor U22982 (N_22982,N_10243,N_15417);
or U22983 (N_22983,N_12964,N_15150);
and U22984 (N_22984,N_17886,N_17283);
or U22985 (N_22985,N_16373,N_15713);
or U22986 (N_22986,N_11723,N_19865);
or U22987 (N_22987,N_10369,N_17057);
nor U22988 (N_22988,N_18785,N_10927);
and U22989 (N_22989,N_12586,N_18934);
nor U22990 (N_22990,N_11742,N_17290);
xor U22991 (N_22991,N_16920,N_14317);
or U22992 (N_22992,N_10840,N_15483);
nand U22993 (N_22993,N_11174,N_17302);
nor U22994 (N_22994,N_12592,N_19797);
or U22995 (N_22995,N_16952,N_19241);
xor U22996 (N_22996,N_11216,N_16967);
and U22997 (N_22997,N_16984,N_12998);
xor U22998 (N_22998,N_10390,N_12603);
or U22999 (N_22999,N_18419,N_15810);
nand U23000 (N_23000,N_15746,N_16416);
nand U23001 (N_23001,N_17584,N_14136);
nor U23002 (N_23002,N_16779,N_16143);
nand U23003 (N_23003,N_18044,N_10512);
xor U23004 (N_23004,N_12157,N_13943);
xnor U23005 (N_23005,N_14400,N_13157);
nand U23006 (N_23006,N_16824,N_18738);
nor U23007 (N_23007,N_19179,N_15529);
nor U23008 (N_23008,N_13760,N_13692);
and U23009 (N_23009,N_17375,N_17643);
and U23010 (N_23010,N_15414,N_19079);
nand U23011 (N_23011,N_18691,N_17352);
or U23012 (N_23012,N_10957,N_15407);
nand U23013 (N_23013,N_18821,N_18574);
and U23014 (N_23014,N_12204,N_16411);
xor U23015 (N_23015,N_17852,N_14711);
xnor U23016 (N_23016,N_19421,N_14729);
nor U23017 (N_23017,N_13012,N_13130);
or U23018 (N_23018,N_14028,N_10499);
and U23019 (N_23019,N_19325,N_13198);
xnor U23020 (N_23020,N_17223,N_13315);
nor U23021 (N_23021,N_16209,N_17413);
or U23022 (N_23022,N_13416,N_13775);
nand U23023 (N_23023,N_15075,N_13664);
xor U23024 (N_23024,N_17179,N_10619);
nand U23025 (N_23025,N_13238,N_13583);
nand U23026 (N_23026,N_19183,N_11785);
xnor U23027 (N_23027,N_13431,N_15984);
xor U23028 (N_23028,N_15210,N_15557);
nor U23029 (N_23029,N_19594,N_16291);
or U23030 (N_23030,N_10970,N_14108);
and U23031 (N_23031,N_15671,N_12092);
or U23032 (N_23032,N_15323,N_12825);
nor U23033 (N_23033,N_11313,N_17980);
or U23034 (N_23034,N_18667,N_17501);
and U23035 (N_23035,N_10844,N_11545);
and U23036 (N_23036,N_13602,N_14821);
and U23037 (N_23037,N_15754,N_16032);
xor U23038 (N_23038,N_18507,N_11406);
xor U23039 (N_23039,N_16385,N_14348);
nand U23040 (N_23040,N_19864,N_19503);
xor U23041 (N_23041,N_14671,N_17956);
nand U23042 (N_23042,N_19736,N_17065);
and U23043 (N_23043,N_10751,N_10574);
and U23044 (N_23044,N_12158,N_16680);
and U23045 (N_23045,N_17848,N_13453);
and U23046 (N_23046,N_17362,N_19188);
and U23047 (N_23047,N_19000,N_14938);
xnor U23048 (N_23048,N_18038,N_14849);
and U23049 (N_23049,N_19315,N_10621);
or U23050 (N_23050,N_15782,N_13165);
nand U23051 (N_23051,N_14941,N_15372);
nand U23052 (N_23052,N_13480,N_11281);
nand U23053 (N_23053,N_13876,N_15654);
nor U23054 (N_23054,N_17806,N_19162);
or U23055 (N_23055,N_10521,N_16070);
nor U23056 (N_23056,N_16393,N_10860);
xor U23057 (N_23057,N_13579,N_12564);
or U23058 (N_23058,N_11800,N_14327);
nor U23059 (N_23059,N_19424,N_11485);
xor U23060 (N_23060,N_14144,N_14119);
nor U23061 (N_23061,N_16242,N_14820);
or U23062 (N_23062,N_17815,N_16635);
and U23063 (N_23063,N_18893,N_17749);
nand U23064 (N_23064,N_12162,N_19844);
xnor U23065 (N_23065,N_12515,N_15040);
nand U23066 (N_23066,N_12491,N_14349);
and U23067 (N_23067,N_19976,N_11795);
xor U23068 (N_23068,N_14513,N_10454);
xnor U23069 (N_23069,N_18339,N_19050);
nand U23070 (N_23070,N_17359,N_10630);
and U23071 (N_23071,N_14092,N_13809);
and U23072 (N_23072,N_13941,N_18855);
or U23073 (N_23073,N_10295,N_10614);
nor U23074 (N_23074,N_19662,N_10913);
nor U23075 (N_23075,N_17047,N_18649);
or U23076 (N_23076,N_18891,N_10254);
or U23077 (N_23077,N_12192,N_14187);
or U23078 (N_23078,N_15141,N_18930);
nor U23079 (N_23079,N_15192,N_15858);
nand U23080 (N_23080,N_19144,N_13868);
xnor U23081 (N_23081,N_16216,N_14812);
xor U23082 (N_23082,N_15943,N_13039);
xor U23083 (N_23083,N_10534,N_16713);
or U23084 (N_23084,N_14861,N_10338);
nor U23085 (N_23085,N_12685,N_10291);
and U23086 (N_23086,N_10929,N_16924);
xnor U23087 (N_23087,N_11706,N_14393);
nand U23088 (N_23088,N_14828,N_14867);
or U23089 (N_23089,N_12010,N_13478);
nand U23090 (N_23090,N_14972,N_19942);
xor U23091 (N_23091,N_16888,N_14185);
or U23092 (N_23092,N_10362,N_17263);
nor U23093 (N_23093,N_19882,N_15993);
nand U23094 (N_23094,N_15213,N_19222);
nor U23095 (N_23095,N_11103,N_13751);
xor U23096 (N_23096,N_15584,N_13016);
nand U23097 (N_23097,N_14537,N_15503);
xnor U23098 (N_23098,N_18237,N_13734);
or U23099 (N_23099,N_12019,N_16131);
nand U23100 (N_23100,N_12078,N_12664);
xnor U23101 (N_23101,N_18845,N_19472);
nor U23102 (N_23102,N_12289,N_11809);
and U23103 (N_23103,N_13683,N_12376);
nand U23104 (N_23104,N_14410,N_19386);
xor U23105 (N_23105,N_11690,N_15000);
nand U23106 (N_23106,N_17870,N_13296);
xnor U23107 (N_23107,N_17365,N_17872);
xnor U23108 (N_23108,N_12270,N_11210);
or U23109 (N_23109,N_11381,N_18682);
nand U23110 (N_23110,N_18186,N_15788);
or U23111 (N_23111,N_12952,N_13000);
or U23112 (N_23112,N_18504,N_16011);
or U23113 (N_23113,N_14242,N_10991);
xnor U23114 (N_23114,N_17594,N_14533);
nand U23115 (N_23115,N_19187,N_12730);
nand U23116 (N_23116,N_19231,N_10947);
xor U23117 (N_23117,N_18563,N_17003);
xnor U23118 (N_23118,N_11447,N_10002);
nand U23119 (N_23119,N_12622,N_13767);
or U23120 (N_23120,N_17287,N_11227);
xor U23121 (N_23121,N_10629,N_12516);
nor U23122 (N_23122,N_11923,N_17188);
and U23123 (N_23123,N_15165,N_15322);
and U23124 (N_23124,N_17364,N_16528);
nor U23125 (N_23125,N_11787,N_19403);
or U23126 (N_23126,N_10434,N_12377);
nor U23127 (N_23127,N_13334,N_10109);
nor U23128 (N_23128,N_19275,N_16978);
or U23129 (N_23129,N_11370,N_10325);
nand U23130 (N_23130,N_16983,N_17882);
xor U23131 (N_23131,N_12411,N_12779);
and U23132 (N_23132,N_14154,N_12894);
and U23133 (N_23133,N_13360,N_11948);
or U23134 (N_23134,N_14077,N_11953);
xor U23135 (N_23135,N_16877,N_17082);
xor U23136 (N_23136,N_18058,N_13792);
nand U23137 (N_23137,N_11250,N_14364);
and U23138 (N_23138,N_12405,N_11801);
xnor U23139 (N_23139,N_17802,N_17014);
and U23140 (N_23140,N_10314,N_12944);
nand U23141 (N_23141,N_12930,N_16313);
xor U23142 (N_23142,N_19106,N_12932);
and U23143 (N_23143,N_19174,N_14652);
and U23144 (N_23144,N_16507,N_13168);
xor U23145 (N_23145,N_11118,N_18632);
and U23146 (N_23146,N_16612,N_11008);
or U23147 (N_23147,N_16467,N_14046);
or U23148 (N_23148,N_10080,N_17200);
xnor U23149 (N_23149,N_17020,N_18645);
and U23150 (N_23150,N_12923,N_12705);
nand U23151 (N_23151,N_13569,N_19970);
nor U23152 (N_23152,N_11432,N_13392);
nor U23153 (N_23153,N_18648,N_16846);
and U23154 (N_23154,N_15091,N_10548);
nor U23155 (N_23155,N_16797,N_13963);
and U23156 (N_23156,N_18082,N_10011);
nand U23157 (N_23157,N_19449,N_12682);
and U23158 (N_23158,N_12835,N_14182);
and U23159 (N_23159,N_14140,N_18183);
nand U23160 (N_23160,N_16509,N_16960);
nand U23161 (N_23161,N_11405,N_18355);
or U23162 (N_23162,N_11011,N_11441);
or U23163 (N_23163,N_13344,N_12419);
or U23164 (N_23164,N_11576,N_19748);
nand U23165 (N_23165,N_19835,N_16417);
nor U23166 (N_23166,N_17262,N_15576);
and U23167 (N_23167,N_14999,N_10636);
or U23168 (N_23168,N_16669,N_11643);
nor U23169 (N_23169,N_16409,N_12610);
and U23170 (N_23170,N_15911,N_18185);
or U23171 (N_23171,N_18407,N_14720);
nand U23172 (N_23172,N_14072,N_15615);
nor U23173 (N_23173,N_12189,N_11813);
and U23174 (N_23174,N_16773,N_16397);
nand U23175 (N_23175,N_14251,N_13701);
nor U23176 (N_23176,N_17328,N_18394);
and U23177 (N_23177,N_14512,N_19510);
xor U23178 (N_23178,N_10414,N_19453);
xor U23179 (N_23179,N_19384,N_10894);
nand U23180 (N_23180,N_13460,N_16871);
xnor U23181 (N_23181,N_10923,N_15533);
nand U23182 (N_23182,N_17340,N_13146);
and U23183 (N_23183,N_10632,N_15215);
and U23184 (N_23184,N_17000,N_15051);
nor U23185 (N_23185,N_15565,N_14181);
or U23186 (N_23186,N_13083,N_14246);
nor U23187 (N_23187,N_14325,N_10848);
xnor U23188 (N_23188,N_10173,N_18135);
and U23189 (N_23189,N_10936,N_11429);
or U23190 (N_23190,N_19992,N_10598);
nand U23191 (N_23191,N_16145,N_11606);
or U23192 (N_23192,N_12280,N_11329);
or U23193 (N_23193,N_16641,N_11956);
nor U23194 (N_23194,N_15196,N_13324);
xnor U23195 (N_23195,N_19536,N_11628);
and U23196 (N_23196,N_16421,N_19950);
and U23197 (N_23197,N_11733,N_17841);
nand U23198 (N_23198,N_11866,N_19289);
or U23199 (N_23199,N_15007,N_12194);
nor U23200 (N_23200,N_11204,N_15606);
xor U23201 (N_23201,N_12085,N_14422);
nand U23202 (N_23202,N_11240,N_12584);
and U23203 (N_23203,N_19303,N_15526);
nor U23204 (N_23204,N_18265,N_13387);
and U23205 (N_23205,N_18029,N_10258);
or U23206 (N_23206,N_17132,N_12232);
and U23207 (N_23207,N_19171,N_18992);
or U23208 (N_23208,N_11705,N_11954);
nor U23209 (N_23209,N_18924,N_15585);
nor U23210 (N_23210,N_10207,N_19444);
and U23211 (N_23211,N_14635,N_10367);
nor U23212 (N_23212,N_18065,N_17346);
nand U23213 (N_23213,N_11913,N_15365);
and U23214 (N_23214,N_15396,N_15898);
nor U23215 (N_23215,N_13473,N_11308);
or U23216 (N_23216,N_12218,N_19373);
or U23217 (N_23217,N_14055,N_14987);
nand U23218 (N_23218,N_17623,N_12860);
xnor U23219 (N_23219,N_11568,N_14829);
xor U23220 (N_23220,N_19129,N_15253);
nand U23221 (N_23221,N_12759,N_18426);
and U23222 (N_23222,N_19192,N_11686);
xor U23223 (N_23223,N_19210,N_13425);
nand U23224 (N_23224,N_14079,N_14193);
xnor U23225 (N_23225,N_14824,N_12482);
and U23226 (N_23226,N_12781,N_15181);
and U23227 (N_23227,N_16683,N_10286);
or U23228 (N_23228,N_10648,N_10416);
nand U23229 (N_23229,N_16942,N_15507);
xor U23230 (N_23230,N_10313,N_16477);
or U23231 (N_23231,N_11760,N_16170);
nor U23232 (N_23232,N_14272,N_11563);
nor U23233 (N_23233,N_16642,N_18193);
and U23234 (N_23234,N_17940,N_18481);
nor U23235 (N_23235,N_15883,N_15023);
xor U23236 (N_23236,N_15015,N_19595);
or U23237 (N_23237,N_19579,N_17353);
and U23238 (N_23238,N_13564,N_10966);
or U23239 (N_23239,N_14582,N_14853);
nand U23240 (N_23240,N_10037,N_13374);
nor U23241 (N_23241,N_10829,N_12286);
or U23242 (N_23242,N_12188,N_10837);
and U23243 (N_23243,N_18440,N_15187);
xnor U23244 (N_23244,N_17632,N_19619);
nor U23245 (N_23245,N_18198,N_15745);
xnor U23246 (N_23246,N_13217,N_11483);
nor U23247 (N_23247,N_16688,N_19263);
nand U23248 (N_23248,N_16238,N_10559);
xor U23249 (N_23249,N_18432,N_10200);
nor U23250 (N_23250,N_11302,N_19722);
and U23251 (N_23251,N_13053,N_17832);
xnor U23252 (N_23252,N_18046,N_19972);
xor U23253 (N_23253,N_15221,N_10024);
nand U23254 (N_23254,N_13368,N_12393);
xnor U23255 (N_23255,N_18293,N_10038);
and U23256 (N_23256,N_17854,N_14633);
or U23257 (N_23257,N_12581,N_13156);
and U23258 (N_23258,N_14105,N_15449);
nor U23259 (N_23259,N_10118,N_17715);
and U23260 (N_23260,N_13421,N_10708);
nand U23261 (N_23261,N_10578,N_13502);
or U23262 (N_23262,N_19184,N_15349);
nor U23263 (N_23263,N_11741,N_17587);
xnor U23264 (N_23264,N_12620,N_18610);
or U23265 (N_23265,N_13182,N_15723);
nor U23266 (N_23266,N_12812,N_16559);
and U23267 (N_23267,N_19861,N_12307);
and U23268 (N_23268,N_16030,N_14104);
nor U23269 (N_23269,N_15358,N_14162);
nor U23270 (N_23270,N_19740,N_12503);
nor U23271 (N_23271,N_13568,N_19264);
or U23272 (N_23272,N_15829,N_15856);
nand U23273 (N_23273,N_15292,N_13687);
or U23274 (N_23274,N_14998,N_14203);
xnor U23275 (N_23275,N_19039,N_10781);
nor U23276 (N_23276,N_13410,N_13603);
xor U23277 (N_23277,N_10698,N_19166);
and U23278 (N_23278,N_13578,N_15162);
or U23279 (N_23279,N_16613,N_18636);
or U23280 (N_23280,N_10253,N_13710);
or U23281 (N_23281,N_18154,N_18519);
xor U23282 (N_23282,N_17453,N_15733);
and U23283 (N_23283,N_18283,N_18128);
nand U23284 (N_23284,N_11952,N_10637);
nand U23285 (N_23285,N_11393,N_15848);
or U23286 (N_23286,N_19389,N_15532);
xnor U23287 (N_23287,N_14749,N_16536);
xnor U23288 (N_23288,N_14402,N_14013);
nor U23289 (N_23289,N_15073,N_14230);
xor U23290 (N_23290,N_14215,N_15249);
or U23291 (N_23291,N_13341,N_11519);
xnor U23292 (N_23292,N_10658,N_19186);
and U23293 (N_23293,N_16848,N_18292);
and U23294 (N_23294,N_11678,N_14070);
and U23295 (N_23295,N_19684,N_19680);
or U23296 (N_23296,N_19327,N_10516);
and U23297 (N_23297,N_14603,N_17158);
nand U23298 (N_23298,N_13535,N_12330);
and U23299 (N_23299,N_10463,N_10633);
or U23300 (N_23300,N_19515,N_19717);
and U23301 (N_23301,N_14997,N_12441);
and U23302 (N_23302,N_10398,N_15687);
xnor U23303 (N_23303,N_15752,N_18933);
or U23304 (N_23304,N_19448,N_16780);
nand U23305 (N_23305,N_13212,N_13384);
xor U23306 (N_23306,N_17117,N_18246);
or U23307 (N_23307,N_17544,N_11017);
nor U23308 (N_23308,N_14981,N_11515);
nor U23309 (N_23309,N_18037,N_19770);
or U23310 (N_23310,N_16602,N_13181);
xnor U23311 (N_23311,N_19796,N_18683);
or U23312 (N_23312,N_19772,N_16886);
and U23313 (N_23313,N_11127,N_13475);
nand U23314 (N_23314,N_10718,N_12574);
nand U23315 (N_23315,N_19860,N_10050);
nand U23316 (N_23316,N_15334,N_16935);
nand U23317 (N_23317,N_15707,N_15442);
xnor U23318 (N_23318,N_11650,N_11337);
xnor U23319 (N_23319,N_14438,N_17504);
nand U23320 (N_23320,N_16639,N_18169);
nor U23321 (N_23321,N_11081,N_17077);
or U23322 (N_23322,N_13646,N_16858);
and U23323 (N_23323,N_18522,N_11054);
and U23324 (N_23324,N_16224,N_18852);
nor U23325 (N_23325,N_10505,N_12688);
and U23326 (N_23326,N_10642,N_17248);
nand U23327 (N_23327,N_18210,N_12006);
and U23328 (N_23328,N_15368,N_12940);
nand U23329 (N_23329,N_19178,N_17770);
or U23330 (N_23330,N_14930,N_19916);
nand U23331 (N_23331,N_13995,N_19656);
xnor U23332 (N_23332,N_19924,N_12485);
nand U23333 (N_23333,N_13232,N_10201);
nor U23334 (N_23334,N_10311,N_19949);
nor U23335 (N_23335,N_14359,N_18147);
and U23336 (N_23336,N_11930,N_15598);
and U23337 (N_23337,N_11050,N_16415);
nand U23338 (N_23338,N_15670,N_14300);
nand U23339 (N_23339,N_10151,N_13143);
or U23340 (N_23340,N_17937,N_10625);
xor U23341 (N_23341,N_16765,N_14780);
nand U23342 (N_23342,N_16667,N_19352);
and U23343 (N_23343,N_10371,N_15638);
nor U23344 (N_23344,N_18299,N_17139);
nor U23345 (N_23345,N_18751,N_19754);
nand U23346 (N_23346,N_17228,N_19250);
or U23347 (N_23347,N_12392,N_15934);
xor U23348 (N_23348,N_13566,N_13968);
nor U23349 (N_23349,N_16456,N_11732);
nand U23350 (N_23350,N_15612,N_10992);
xor U23351 (N_23351,N_13699,N_19271);
and U23352 (N_23352,N_18867,N_11151);
xnor U23353 (N_23353,N_18814,N_16175);
or U23354 (N_23354,N_10235,N_13277);
nand U23355 (N_23355,N_12041,N_11239);
and U23356 (N_23356,N_10407,N_14741);
nor U23357 (N_23357,N_18208,N_13259);
xnor U23358 (N_23358,N_15768,N_19112);
nand U23359 (N_23359,N_15655,N_19945);
and U23360 (N_23360,N_16835,N_11858);
nor U23361 (N_23361,N_14988,N_14851);
xnor U23362 (N_23362,N_18428,N_10832);
xor U23363 (N_23363,N_14116,N_11452);
nand U23364 (N_23364,N_15857,N_12802);
or U23365 (N_23365,N_19426,N_16320);
and U23366 (N_23366,N_14575,N_15604);
nand U23367 (N_23367,N_15479,N_15342);
or U23368 (N_23368,N_11436,N_17746);
nand U23369 (N_23369,N_16472,N_15855);
xor U23370 (N_23370,N_14054,N_16821);
xor U23371 (N_23371,N_12145,N_14169);
nor U23372 (N_23372,N_19034,N_19286);
nor U23373 (N_23373,N_13218,N_17553);
nor U23374 (N_23374,N_16214,N_14563);
nand U23375 (N_23375,N_15241,N_19238);
and U23376 (N_23376,N_17609,N_11699);
nand U23377 (N_23377,N_19356,N_11493);
nor U23378 (N_23378,N_16060,N_17106);
nor U23379 (N_23379,N_15992,N_12046);
or U23380 (N_23380,N_13859,N_15554);
xnor U23381 (N_23381,N_17123,N_18284);
or U23382 (N_23382,N_13961,N_18401);
and U23383 (N_23383,N_17788,N_11198);
nor U23384 (N_23384,N_14636,N_14383);
and U23385 (N_23385,N_14141,N_16344);
nand U23386 (N_23386,N_14510,N_19678);
or U23387 (N_23387,N_19193,N_18364);
nand U23388 (N_23388,N_15964,N_11534);
and U23389 (N_23389,N_17684,N_13147);
or U23390 (N_23390,N_17551,N_12196);
nor U23391 (N_23391,N_14758,N_17786);
and U23392 (N_23392,N_12281,N_16831);
and U23393 (N_23393,N_10631,N_12238);
xnor U23394 (N_23394,N_15347,N_11126);
nand U23395 (N_23395,N_11975,N_11604);
nor U23396 (N_23396,N_13544,N_14074);
and U23397 (N_23397,N_10316,N_12294);
and U23398 (N_23398,N_11580,N_12625);
xnor U23399 (N_23399,N_15424,N_11497);
xnor U23400 (N_23400,N_11846,N_10715);
xor U23401 (N_23401,N_14857,N_12684);
nand U23402 (N_23402,N_16492,N_10472);
xor U23403 (N_23403,N_11774,N_19064);
xnor U23404 (N_23404,N_17620,N_16119);
or U23405 (N_23405,N_19836,N_19148);
nand U23406 (N_23406,N_15453,N_16305);
xnor U23407 (N_23407,N_12970,N_19991);
and U23408 (N_23408,N_17707,N_19556);
nor U23409 (N_23409,N_13899,N_18114);
and U23410 (N_23410,N_17463,N_12768);
or U23411 (N_23411,N_13925,N_18622);
or U23412 (N_23412,N_19119,N_14559);
nor U23413 (N_23413,N_16140,N_17370);
and U23414 (N_23414,N_12758,N_17572);
xnor U23415 (N_23415,N_10119,N_16893);
and U23416 (N_23416,N_18819,N_16926);
and U23417 (N_23417,N_15276,N_14407);
xnor U23418 (N_23418,N_11448,N_15067);
xnor U23419 (N_23419,N_17438,N_13363);
nor U23420 (N_23420,N_15439,N_12316);
xor U23421 (N_23421,N_15999,N_14665);
xor U23422 (N_23422,N_19168,N_16438);
xnor U23423 (N_23423,N_10379,N_14335);
nor U23424 (N_23424,N_11888,N_11827);
nand U23425 (N_23425,N_14674,N_14757);
and U23426 (N_23426,N_15268,N_16104);
or U23427 (N_23427,N_16122,N_18621);
nand U23428 (N_23428,N_17345,N_13273);
nor U23429 (N_23429,N_17938,N_19445);
nor U23430 (N_23430,N_17401,N_10141);
and U23431 (N_23431,N_14088,N_11459);
xor U23432 (N_23432,N_15790,N_16473);
and U23433 (N_23433,N_13849,N_18991);
xnor U23434 (N_23434,N_19235,N_18403);
xor U23435 (N_23435,N_19152,N_18420);
or U23436 (N_23436,N_10665,N_16458);
or U23437 (N_23437,N_10609,N_18693);
nor U23438 (N_23438,N_15549,N_18681);
and U23439 (N_23439,N_13625,N_13090);
xor U23440 (N_23440,N_17782,N_11603);
xor U23441 (N_23441,N_19621,N_11767);
or U23442 (N_23442,N_15229,N_18312);
or U23443 (N_23443,N_14087,N_18960);
nand U23444 (N_23444,N_15307,N_17436);
and U23445 (N_23445,N_15722,N_11738);
or U23446 (N_23446,N_19753,N_17156);
nor U23447 (N_23447,N_19190,N_11136);
nor U23448 (N_23448,N_13027,N_13051);
or U23449 (N_23449,N_16134,N_18910);
nand U23450 (N_23450,N_11664,N_10853);
or U23451 (N_23451,N_12248,N_19600);
or U23452 (N_23452,N_16464,N_11757);
and U23453 (N_23453,N_17622,N_10833);
xnor U23454 (N_23454,N_16298,N_16661);
nand U23455 (N_23455,N_11330,N_10880);
or U23456 (N_23456,N_19552,N_16516);
xor U23457 (N_23457,N_18499,N_11577);
or U23458 (N_23458,N_15811,N_19553);
and U23459 (N_23459,N_13932,N_14943);
and U23460 (N_23460,N_11206,N_13757);
nor U23461 (N_23461,N_11874,N_11737);
xnor U23462 (N_23462,N_15990,N_15784);
nor U23463 (N_23463,N_13251,N_12607);
and U23464 (N_23464,N_14838,N_15127);
or U23465 (N_23465,N_13960,N_18410);
or U23466 (N_23466,N_19081,N_14352);
nand U23467 (N_23467,N_18856,N_16857);
or U23468 (N_23468,N_10033,N_18371);
or U23469 (N_23469,N_12967,N_12431);
and U23470 (N_23470,N_15427,N_12487);
nand U23471 (N_23471,N_11093,N_19732);
and U23472 (N_23472,N_19494,N_17154);
and U23473 (N_23473,N_12185,N_16394);
nand U23474 (N_23474,N_18698,N_14624);
nand U23475 (N_23475,N_14413,N_16144);
nor U23476 (N_23476,N_15699,N_13002);
nand U23477 (N_23477,N_13435,N_11541);
xnor U23478 (N_23478,N_10897,N_11680);
or U23479 (N_23479,N_16328,N_12526);
and U23480 (N_23480,N_17430,N_15972);
nand U23481 (N_23481,N_15082,N_17732);
or U23482 (N_23482,N_12437,N_14990);
nand U23483 (N_23483,N_19788,N_19961);
xnor U23484 (N_23484,N_13370,N_18141);
nand U23485 (N_23485,N_12593,N_19833);
xor U23486 (N_23486,N_11531,N_14126);
and U23487 (N_23487,N_12084,N_14163);
nand U23488 (N_23488,N_18304,N_12648);
nand U23489 (N_23489,N_15147,N_16475);
nor U23490 (N_23490,N_12047,N_15401);
and U23491 (N_23491,N_18351,N_11752);
nand U23492 (N_23492,N_17208,N_10335);
xnor U23493 (N_23493,N_18961,N_12276);
and U23494 (N_23494,N_10261,N_17450);
or U23495 (N_23495,N_18639,N_15062);
xor U23496 (N_23496,N_13624,N_16904);
or U23497 (N_23497,N_18203,N_17325);
nand U23498 (N_23498,N_12239,N_13314);
and U23499 (N_23499,N_13937,N_12956);
nand U23500 (N_23500,N_15348,N_18594);
and U23501 (N_23501,N_16461,N_11046);
or U23502 (N_23502,N_11535,N_12983);
and U23503 (N_23503,N_11324,N_10799);
xor U23504 (N_23504,N_19601,N_13220);
xnor U23505 (N_23505,N_16484,N_11933);
nand U23506 (N_23506,N_10674,N_11195);
and U23507 (N_23507,N_14775,N_14968);
or U23508 (N_23508,N_11117,N_13807);
or U23509 (N_23509,N_12418,N_18343);
xnor U23510 (N_23510,N_11513,N_13908);
xnor U23511 (N_23511,N_10343,N_15287);
or U23512 (N_23512,N_13004,N_13675);
or U23513 (N_23513,N_14361,N_15714);
nor U23514 (N_23514,N_14340,N_14284);
xor U23515 (N_23515,N_13884,N_15328);
nor U23516 (N_23516,N_19698,N_19387);
nor U23517 (N_23517,N_13380,N_11225);
nor U23518 (N_23518,N_11944,N_17903);
xnor U23519 (N_23519,N_17429,N_13907);
and U23520 (N_23520,N_12479,N_17048);
nor U23521 (N_23521,N_10756,N_13539);
nor U23522 (N_23522,N_17973,N_16208);
nand U23523 (N_23523,N_19443,N_16348);
nor U23524 (N_23524,N_11311,N_11980);
xnor U23525 (N_23525,N_19947,N_12976);
or U23526 (N_23526,N_12357,N_19225);
and U23527 (N_23527,N_15628,N_10039);
xor U23528 (N_23528,N_15823,N_18760);
or U23529 (N_23529,N_10816,N_17640);
nor U23530 (N_23530,N_16801,N_15691);
or U23531 (N_23531,N_17227,N_16764);
xor U23532 (N_23532,N_15632,N_11407);
or U23533 (N_23533,N_19219,N_15539);
nor U23534 (N_23534,N_15773,N_15664);
xnor U23535 (N_23535,N_14338,N_16606);
and U23536 (N_23536,N_15770,N_15852);
nand U23537 (N_23537,N_11695,N_10441);
and U23538 (N_23538,N_17217,N_18006);
nand U23539 (N_23539,N_18749,N_13356);
nor U23540 (N_23540,N_13531,N_12727);
and U23541 (N_23541,N_18589,N_10701);
xnor U23542 (N_23542,N_11289,N_14663);
nand U23543 (N_23543,N_10902,N_10158);
and U23544 (N_23544,N_17899,N_10236);
nand U23545 (N_23545,N_13745,N_15510);
nor U23546 (N_23546,N_13032,N_18940);
nand U23547 (N_23547,N_13065,N_16603);
and U23548 (N_23548,N_10350,N_17424);
nor U23549 (N_23549,N_16027,N_18863);
or U23550 (N_23550,N_13070,N_13588);
xor U23551 (N_23551,N_13820,N_11682);
xor U23552 (N_23552,N_13529,N_10444);
and U23553 (N_23553,N_11710,N_10442);
and U23554 (N_23554,N_18241,N_19630);
nand U23555 (N_23555,N_10671,N_13879);
or U23556 (N_23556,N_10532,N_15072);
nor U23557 (N_23557,N_14224,N_17888);
and U23558 (N_23558,N_10308,N_17922);
or U23559 (N_23559,N_11955,N_19425);
nand U23560 (N_23560,N_18110,N_16625);
xnor U23561 (N_23561,N_16217,N_13038);
nor U23562 (N_23562,N_17164,N_16036);
nand U23563 (N_23563,N_19626,N_10842);
nand U23564 (N_23564,N_15508,N_17206);
nor U23565 (N_23565,N_10005,N_12464);
and U23566 (N_23566,N_10110,N_16364);
xnor U23567 (N_23567,N_18905,N_15978);
nand U23568 (N_23568,N_11338,N_13349);
nor U23569 (N_23569,N_19878,N_10834);
or U23570 (N_23570,N_15359,N_19682);
or U23571 (N_23571,N_13852,N_17286);
xnor U23572 (N_23572,N_11094,N_19688);
and U23573 (N_23573,N_18859,N_17451);
or U23574 (N_23574,N_15715,N_16211);
nand U23575 (N_23575,N_16066,N_13074);
or U23576 (N_23576,N_17068,N_12279);
and U23577 (N_23577,N_17472,N_14841);
nand U23578 (N_23578,N_12679,N_16086);
xor U23579 (N_23579,N_12427,N_10130);
and U23580 (N_23580,N_17783,N_19679);
nor U23581 (N_23581,N_10241,N_11900);
nor U23582 (N_23582,N_11408,N_19533);
xor U23583 (N_23583,N_10801,N_13303);
and U23584 (N_23584,N_19357,N_19948);
or U23585 (N_23585,N_14915,N_18032);
nand U23586 (N_23586,N_15045,N_16679);
nor U23587 (N_23587,N_11668,N_16334);
nand U23588 (N_23588,N_11660,N_18672);
and U23589 (N_23589,N_12565,N_19369);
and U23590 (N_23590,N_19528,N_13418);
and U23591 (N_23591,N_17548,N_17222);
and U23592 (N_23592,N_13642,N_13977);
nor U23593 (N_23593,N_17041,N_10196);
or U23594 (N_23594,N_14762,N_12918);
or U23595 (N_23595,N_15688,N_12349);
xor U23596 (N_23596,N_17449,N_12770);
and U23597 (N_23597,N_16883,N_13121);
nor U23598 (N_23598,N_19640,N_14610);
xnor U23599 (N_23599,N_13428,N_16293);
nand U23600 (N_23600,N_13362,N_13379);
xor U23601 (N_23601,N_17086,N_16784);
and U23602 (N_23602,N_17803,N_11632);
or U23603 (N_23603,N_15083,N_10930);
and U23604 (N_23604,N_19223,N_11342);
nand U23605 (N_23605,N_15384,N_19609);
xnor U23606 (N_23606,N_17771,N_11612);
xor U23607 (N_23607,N_11608,N_15816);
xor U23608 (N_23608,N_14601,N_14042);
nor U23609 (N_23609,N_11635,N_16153);
or U23610 (N_23610,N_13268,N_15364);
xor U23611 (N_23611,N_15668,N_16440);
and U23612 (N_23612,N_18640,N_16862);
xnor U23613 (N_23613,N_13555,N_17138);
and U23614 (N_23614,N_13799,N_13670);
nand U23615 (N_23615,N_18704,N_15090);
nor U23616 (N_23616,N_10628,N_11312);
nand U23617 (N_23617,N_12315,N_11412);
xor U23618 (N_23618,N_17743,N_12202);
nand U23619 (N_23619,N_13123,N_19975);
xnor U23620 (N_23620,N_13280,N_12395);
or U23621 (N_23621,N_11319,N_12079);
or U23622 (N_23622,N_14843,N_18890);
nor U23623 (N_23623,N_14598,N_17718);
nor U23624 (N_23624,N_17592,N_10013);
nor U23625 (N_23625,N_16717,N_19274);
or U23626 (N_23626,N_19658,N_19084);
xor U23627 (N_23627,N_12335,N_18875);
nor U23628 (N_23628,N_14477,N_18287);
or U23629 (N_23629,N_17824,N_19450);
nor U23630 (N_23630,N_14239,N_19393);
nand U23631 (N_23631,N_15484,N_12796);
and U23632 (N_23632,N_10219,N_18373);
nor U23633 (N_23633,N_19036,N_13073);
xnor U23634 (N_23634,N_11689,N_11266);
nor U23635 (N_23635,N_15103,N_13862);
nor U23636 (N_23636,N_10364,N_15340);
nand U23637 (N_23637,N_18695,N_13186);
nor U23638 (N_23638,N_15336,N_18334);
nand U23639 (N_23639,N_13882,N_19807);
or U23640 (N_23640,N_15573,N_12115);
or U23641 (N_23641,N_13553,N_15844);
nor U23642 (N_23642,N_14249,N_14925);
nand U23643 (N_23643,N_14473,N_15515);
or U23644 (N_23644,N_18151,N_11259);
nand U23645 (N_23645,N_18078,N_12869);
nand U23646 (N_23646,N_19312,N_10091);
nor U23647 (N_23647,N_12544,N_13193);
and U23648 (N_23648,N_11377,N_17892);
nand U23649 (N_23649,N_12961,N_14446);
and U23650 (N_23650,N_18126,N_17153);
or U23651 (N_23651,N_16600,N_19708);
xnor U23652 (N_23652,N_15572,N_14294);
nand U23653 (N_23653,N_12599,N_19787);
nand U23654 (N_23654,N_17249,N_13404);
and U23655 (N_23655,N_17828,N_12884);
and U23656 (N_23656,N_19841,N_14730);
and U23657 (N_23657,N_11520,N_10919);
or U23658 (N_23658,N_10882,N_18569);
xor U23659 (N_23659,N_19489,N_17916);
nor U23660 (N_23660,N_12187,N_12489);
nor U23661 (N_23661,N_18486,N_13451);
xor U23662 (N_23662,N_10108,N_10474);
or U23663 (N_23663,N_17911,N_12314);
and U23664 (N_23664,N_17858,N_17838);
nand U23665 (N_23665,N_11261,N_18423);
nor U23666 (N_23666,N_18902,N_13087);
xnor U23667 (N_23667,N_19170,N_13994);
nand U23668 (N_23668,N_11178,N_11186);
nor U23669 (N_23669,N_15193,N_10239);
and U23670 (N_23670,N_12467,N_12061);
xnor U23671 (N_23671,N_17583,N_11158);
xor U23672 (N_23672,N_11388,N_15466);
or U23673 (N_23673,N_18326,N_10971);
and U23674 (N_23674,N_16757,N_14769);
nand U23675 (N_23675,N_10387,N_14910);
xor U23676 (N_23676,N_14952,N_11536);
and U23677 (N_23677,N_18014,N_16391);
xor U23678 (N_23678,N_15459,N_10055);
nor U23679 (N_23679,N_17853,N_19994);
and U23680 (N_23680,N_12412,N_15487);
nor U23681 (N_23681,N_16572,N_13593);
nand U23682 (N_23682,N_12312,N_12128);
or U23683 (N_23683,N_19493,N_12790);
or U23684 (N_23684,N_12264,N_17563);
nand U23685 (N_23685,N_19309,N_13028);
xor U23686 (N_23686,N_16535,N_14270);
nor U23687 (N_23687,N_11402,N_15217);
nor U23688 (N_23688,N_17355,N_15254);
nand U23689 (N_23689,N_13720,N_16622);
nand U23690 (N_23690,N_13382,N_13266);
and U23691 (N_23691,N_17842,N_18289);
or U23692 (N_23692,N_11897,N_10546);
and U23693 (N_23693,N_11468,N_14623);
or U23694 (N_23694,N_11971,N_13317);
nand U23695 (N_23695,N_16538,N_10285);
nor U23696 (N_23696,N_19334,N_13634);
nor U23697 (N_23697,N_19211,N_13316);
and U23698 (N_23698,N_17369,N_18354);
or U23699 (N_23699,N_19584,N_16166);
nand U23700 (N_23700,N_16178,N_12749);
nand U23701 (N_23701,N_16360,N_16092);
and U23702 (N_23702,N_14516,N_14073);
or U23703 (N_23703,N_17954,N_13563);
xnor U23704 (N_23704,N_13383,N_14859);
nor U23705 (N_23705,N_15122,N_11446);
nand U23706 (N_23706,N_14481,N_14889);
and U23707 (N_23707,N_12614,N_11755);
and U23708 (N_23708,N_11821,N_18947);
and U23709 (N_23709,N_12474,N_18936);
and U23710 (N_23710,N_17736,N_11418);
or U23711 (N_23711,N_17724,N_19128);
xor U23712 (N_23712,N_11164,N_15232);
or U23713 (N_23713,N_10457,N_13688);
and U23714 (N_23714,N_18901,N_13819);
xnor U23715 (N_23715,N_18865,N_11645);
nand U23716 (N_23716,N_18488,N_14275);
and U23717 (N_23717,N_16946,N_11419);
or U23718 (N_23718,N_10709,N_17536);
or U23719 (N_23719,N_10178,N_14258);
and U23720 (N_23720,N_12640,N_15481);
and U23721 (N_23721,N_15014,N_13046);
nand U23722 (N_23722,N_14458,N_14554);
xnor U23723 (N_23723,N_16981,N_19946);
and U23724 (N_23724,N_11208,N_14200);
and U23725 (N_23725,N_13489,N_12578);
and U23726 (N_23726,N_15004,N_17883);
nor U23727 (N_23727,N_12234,N_14872);
and U23728 (N_23728,N_19280,N_11596);
xor U23729 (N_23729,N_14836,N_17813);
xnor U23730 (N_23730,N_19530,N_19548);
and U23731 (N_23731,N_19486,N_15940);
and U23732 (N_23732,N_14161,N_18022);
or U23733 (N_23733,N_12074,N_19433);
or U23734 (N_23734,N_11546,N_16408);
nand U23735 (N_23735,N_11881,N_14660);
and U23736 (N_23736,N_16449,N_16125);
nor U23737 (N_23737,N_19333,N_11637);
xnor U23738 (N_23738,N_16541,N_18218);
nor U23739 (N_23739,N_18043,N_13987);
xnor U23740 (N_23740,N_13022,N_19815);
or U23741 (N_23741,N_14339,N_13726);
or U23742 (N_23742,N_18788,N_14213);
nor U23743 (N_23743,N_12142,N_14282);
nor U23744 (N_23744,N_14869,N_18737);
nand U23745 (N_23745,N_12719,N_17616);
xor U23746 (N_23746,N_12525,N_16766);
or U23747 (N_23747,N_14924,N_12861);
or U23748 (N_23748,N_15233,N_17647);
xnor U23749 (N_23749,N_10912,N_15900);
nand U23750 (N_23750,N_11573,N_10693);
xnor U23751 (N_23751,N_12654,N_13705);
or U23752 (N_23752,N_13546,N_13904);
and U23753 (N_23753,N_16035,N_14444);
nor U23754 (N_23754,N_13354,N_12535);
nor U23755 (N_23755,N_13824,N_10331);
nor U23756 (N_23756,N_13313,N_18858);
or U23757 (N_23757,N_16020,N_13207);
xnor U23758 (N_23758,N_16806,N_17861);
and U23759 (N_23759,N_11523,N_17368);
and U23760 (N_23760,N_16752,N_17680);
xnor U23761 (N_23761,N_17066,N_12140);
xor U23762 (N_23762,N_12017,N_12865);
and U23763 (N_23763,N_15941,N_15969);
xnor U23764 (N_23764,N_14363,N_10763);
and U23765 (N_23765,N_11383,N_10891);
and U23766 (N_23766,N_19103,N_16129);
xor U23767 (N_23767,N_18062,N_18384);
nand U23768 (N_23768,N_17682,N_16095);
xnor U23769 (N_23769,N_11716,N_12543);
nor U23770 (N_23770,N_14798,N_18482);
and U23771 (N_23771,N_13111,N_11058);
xor U23772 (N_23772,N_16269,N_11035);
nand U23773 (N_23773,N_19082,N_18238);
or U23774 (N_23774,N_17456,N_17765);
nor U23775 (N_23775,N_17755,N_12355);
xor U23776 (N_23776,N_15509,N_11722);
nand U23777 (N_23777,N_12130,N_15402);
xnor U23778 (N_23778,N_12563,N_11958);
or U23779 (N_23779,N_18480,N_19012);
nor U23780 (N_23780,N_13903,N_10895);
and U23781 (N_23781,N_19094,N_18647);
or U23782 (N_23782,N_14416,N_10557);
nor U23783 (N_23783,N_13408,N_10150);
nor U23784 (N_23784,N_18541,N_13040);
nand U23785 (N_23785,N_18872,N_17107);
nand U23786 (N_23786,N_10900,N_16120);
and U23787 (N_23787,N_19927,N_13841);
xnor U23788 (N_23788,N_19143,N_15462);
or U23789 (N_23789,N_16107,N_16929);
nand U23790 (N_23790,N_14785,N_10352);
nand U23791 (N_23791,N_18728,N_10144);
nand U23792 (N_23792,N_14110,N_10125);
or U23793 (N_23793,N_18921,N_17356);
nor U23794 (N_23794,N_17519,N_13975);
nor U23795 (N_23795,N_16826,N_13523);
nand U23796 (N_23796,N_11269,N_18892);
nor U23797 (N_23797,N_11188,N_11394);
nor U23798 (N_23798,N_13201,N_13959);
nor U23799 (N_23799,N_16540,N_12982);
nand U23800 (N_23800,N_19531,N_17322);
nand U23801 (N_23801,N_15552,N_17710);
nand U23802 (N_23802,N_17466,N_14463);
and U23803 (N_23803,N_18514,N_14342);
nand U23804 (N_23804,N_18016,N_17395);
and U23805 (N_23805,N_14451,N_16085);
nand U23806 (N_23806,N_14519,N_19813);
nor U23807 (N_23807,N_10825,N_11823);
and U23808 (N_23808,N_17441,N_18414);
or U23809 (N_23809,N_16803,N_16169);
nand U23810 (N_23810,N_17796,N_15862);
or U23811 (N_23811,N_16446,N_15591);
nor U23812 (N_23812,N_18575,N_18555);
xnor U23813 (N_23813,N_19743,N_18658);
xor U23814 (N_23814,N_12873,N_17876);
nor U23815 (N_23815,N_15120,N_12848);
and U23816 (N_23816,N_14581,N_19905);
or U23817 (N_23817,N_18763,N_18438);
and U23818 (N_23818,N_11771,N_16812);
and U23819 (N_23819,N_14358,N_14415);
and U23820 (N_23820,N_18701,N_16666);
xor U23821 (N_23821,N_17058,N_18671);
nor U23822 (N_23822,N_18064,N_10544);
nor U23823 (N_23823,N_16585,N_10997);
and U23824 (N_23824,N_14687,N_13823);
xor U23825 (N_23825,N_10726,N_14056);
nand U23826 (N_23826,N_11160,N_14445);
xor U23827 (N_23827,N_19245,N_13871);
and U23828 (N_23828,N_19557,N_11882);
or U23829 (N_23829,N_17276,N_12433);
or U23830 (N_23830,N_11521,N_15121);
nand U23831 (N_23831,N_14744,N_15611);
nor U23832 (N_23832,N_11155,N_10386);
nand U23833 (N_23833,N_11806,N_17864);
xor U23834 (N_23834,N_16333,N_18623);
nand U23835 (N_23835,N_14387,N_19659);
nor U23836 (N_23836,N_11469,N_19762);
or U23837 (N_23837,N_10093,N_10453);
or U23838 (N_23838,N_18719,N_18543);
xor U23839 (N_23839,N_11773,N_14311);
nand U23840 (N_23840,N_12810,N_19879);
or U23841 (N_23841,N_12060,N_13617);
nor U23842 (N_23842,N_17618,N_17439);
xnor U23843 (N_23843,N_18713,N_17331);
or U23844 (N_23844,N_14443,N_19432);
nor U23845 (N_23845,N_17053,N_15142);
nor U23846 (N_23846,N_18344,N_18615);
nand U23847 (N_23847,N_16547,N_17306);
xnor U23848 (N_23848,N_12053,N_18021);
or U23849 (N_23849,N_13700,N_18796);
or U23850 (N_23850,N_10203,N_14365);
or U23851 (N_23851,N_11403,N_13472);
nor U23852 (N_23852,N_14964,N_13192);
xor U23853 (N_23853,N_17961,N_15837);
xnor U23854 (N_23854,N_17662,N_15374);
or U23855 (N_23855,N_11976,N_13295);
nor U23856 (N_23856,N_10494,N_12539);
xor U23857 (N_23857,N_15080,N_11098);
nand U23858 (N_23858,N_11679,N_13989);
xor U23859 (N_23859,N_10447,N_13986);
xor U23860 (N_23860,N_17400,N_19939);
or U23861 (N_23861,N_18112,N_18069);
nor U23862 (N_23862,N_19936,N_15068);
or U23863 (N_23863,N_15108,N_11055);
or U23864 (N_23864,N_15913,N_18817);
xnor U23865 (N_23865,N_14091,N_19713);
xor U23866 (N_23866,N_12233,N_10917);
and U23867 (N_23867,N_18943,N_14155);
nor U23868 (N_23868,N_18009,N_19290);
xor U23869 (N_23869,N_14735,N_14707);
nor U23870 (N_23870,N_16489,N_16795);
nand U23871 (N_23871,N_19197,N_15923);
and U23872 (N_23872,N_11551,N_10871);
nor U23873 (N_23873,N_12585,N_11409);
or U23874 (N_23874,N_10035,N_10983);
nand U23875 (N_23875,N_18966,N_14727);
and U23876 (N_23876,N_18606,N_13962);
nand U23877 (N_23877,N_12367,N_19941);
or U23878 (N_23878,N_10376,N_10294);
nor U23879 (N_23879,N_14960,N_10710);
and U23880 (N_23880,N_13126,N_12635);
or U23881 (N_23881,N_11364,N_11427);
or U23882 (N_23882,N_15310,N_19466);
nand U23883 (N_23883,N_18600,N_11481);
xor U23884 (N_23884,N_16565,N_16802);
nand U23885 (N_23885,N_11623,N_14497);
or U23886 (N_23886,N_16610,N_19873);
and U23887 (N_23887,N_10190,N_12822);
and U23888 (N_23888,N_13885,N_15899);
and U23889 (N_23889,N_15478,N_14264);
nor U23890 (N_23890,N_10074,N_14546);
and U23891 (N_23891,N_16468,N_17566);
nand U23892 (N_23892,N_11348,N_13752);
xor U23893 (N_23893,N_13290,N_12686);
nand U23894 (N_23894,N_15493,N_15965);
xor U23895 (N_23895,N_13318,N_14679);
xor U23896 (N_23896,N_15544,N_12151);
nor U23897 (N_23897,N_19663,N_17696);
and U23898 (N_23898,N_11461,N_11951);
or U23899 (N_23899,N_11462,N_11613);
or U23900 (N_23900,N_11185,N_14937);
or U23901 (N_23901,N_15845,N_15463);
xnor U23902 (N_23902,N_19016,N_13682);
and U23903 (N_23903,N_15512,N_12996);
and U23904 (N_23904,N_13394,N_12222);
and U23905 (N_23905,N_17908,N_15211);
nor U23906 (N_23906,N_12356,N_12246);
nand U23907 (N_23907,N_10540,N_15960);
or U23908 (N_23908,N_10538,N_13252);
xnor U23909 (N_23909,N_15772,N_19408);
or U23910 (N_23910,N_17999,N_11392);
or U23911 (N_23911,N_16257,N_19310);
nand U23912 (N_23912,N_10277,N_17821);
nand U23913 (N_23913,N_17282,N_12484);
nand U23914 (N_23914,N_10922,N_15665);
nor U23915 (N_23915,N_13308,N_17727);
nor U23916 (N_23916,N_14290,N_13984);
or U23917 (N_23917,N_12808,N_18191);
and U23918 (N_23918,N_18997,N_12457);
nand U23919 (N_23919,N_17699,N_16377);
xnor U23920 (N_23920,N_17033,N_11728);
xor U23921 (N_23921,N_18429,N_19705);
and U23922 (N_23922,N_19779,N_18372);
nand U23923 (N_23923,N_10836,N_15099);
xor U23924 (N_23924,N_17140,N_10975);
xnor U23925 (N_23925,N_14953,N_19158);
xnor U23926 (N_23926,N_17670,N_10282);
or U23927 (N_23927,N_10152,N_12095);
or U23928 (N_23928,N_12094,N_16562);
xor U23929 (N_23929,N_18637,N_16447);
nand U23930 (N_23930,N_10849,N_17700);
xor U23931 (N_23931,N_14752,N_13936);
nor U23932 (N_23932,N_16880,N_13572);
and U23933 (N_23933,N_15281,N_13608);
and U23934 (N_23934,N_13611,N_14330);
or U23935 (N_23935,N_15354,N_10672);
or U23936 (N_23936,N_10768,N_12997);
nor U23937 (N_23937,N_11842,N_18718);
nand U23938 (N_23938,N_10347,N_11826);
nor U23939 (N_23939,N_11986,N_11616);
or U23940 (N_23940,N_15521,N_19142);
and U23941 (N_23941,N_11138,N_18980);
and U23942 (N_23942,N_12127,N_18399);
and U23943 (N_23943,N_14742,N_14491);
nor U23944 (N_23944,N_15248,N_11764);
and U23945 (N_23945,N_16268,N_13166);
or U23946 (N_23946,N_14959,N_12080);
nand U23947 (N_23947,N_16252,N_19492);
or U23948 (N_23948,N_11875,N_19321);
nor U23949 (N_23949,N_14069,N_15683);
and U23950 (N_23950,N_18473,N_16810);
nor U23951 (N_23951,N_17105,N_13631);
and U23952 (N_23952,N_17664,N_19585);
or U23953 (N_23953,N_17679,N_17641);
and U23954 (N_23954,N_19015,N_15170);
nand U23955 (N_23955,N_17627,N_15428);
or U23956 (N_23956,N_13855,N_17570);
nand U23957 (N_23957,N_14117,N_13677);
nand U23958 (N_23958,N_17656,N_17099);
and U23959 (N_23959,N_11375,N_17859);
or U23960 (N_23960,N_11367,N_10954);
and U23961 (N_23961,N_15393,N_13443);
or U23962 (N_23962,N_12160,N_18085);
xnor U23963 (N_23963,N_18149,N_14877);
and U23964 (N_23964,N_18184,N_11358);
nor U23965 (N_23965,N_11884,N_16897);
nand U23966 (N_23966,N_10670,N_10307);
nor U23967 (N_23967,N_10762,N_14248);
or U23968 (N_23968,N_17895,N_16015);
xor U23969 (N_23969,N_18067,N_10723);
nor U23970 (N_23970,N_17270,N_16814);
xor U23971 (N_23971,N_11949,N_19488);
or U23972 (N_23972,N_15741,N_13250);
xor U23973 (N_23973,N_11550,N_12476);
nand U23974 (N_23974,N_12633,N_13842);
or U23975 (N_23975,N_18888,N_16367);
nor U23976 (N_23976,N_11700,N_18483);
or U23977 (N_23977,N_19644,N_16638);
nand U23978 (N_23978,N_12269,N_14894);
xor U23979 (N_23979,N_14420,N_17559);
or U23980 (N_23980,N_18298,N_17752);
xor U23981 (N_23981,N_12743,N_13423);
and U23982 (N_23982,N_19765,N_11638);
xnor U23983 (N_23983,N_13518,N_16274);
xor U23984 (N_23984,N_15918,N_13898);
or U23985 (N_23985,N_16957,N_16080);
nor U23986 (N_23986,N_15476,N_19248);
nand U23987 (N_23987,N_15779,N_18989);
or U23988 (N_23988,N_11202,N_15046);
and U23989 (N_23989,N_10995,N_19683);
and U23990 (N_23990,N_17651,N_10627);
and U23991 (N_23991,N_10165,N_13851);
nor U23992 (N_23992,N_16220,N_18327);
or U23993 (N_23993,N_12350,N_10925);
xor U23994 (N_23994,N_17851,N_19872);
xor U23995 (N_23995,N_19216,N_15139);
nand U23996 (N_23996,N_17991,N_10582);
and U23997 (N_23997,N_16204,N_17312);
nor U23998 (N_23998,N_13723,N_18611);
or U23999 (N_23999,N_16490,N_18431);
nand U24000 (N_24000,N_14774,N_11006);
xor U24001 (N_24001,N_14675,N_14235);
or U24002 (N_24002,N_16323,N_11765);
nor U24003 (N_24003,N_13641,N_16571);
nor U24004 (N_24004,N_12765,N_10771);
or U24005 (N_24005,N_13746,N_11097);
or U24006 (N_24006,N_15569,N_12916);
or U24007 (N_24007,N_10310,N_15329);
or U24008 (N_24008,N_18047,N_12422);
nor U24009 (N_24009,N_10461,N_10826);
or U24010 (N_24010,N_18071,N_16789);
nand U24011 (N_24011,N_10493,N_14902);
nor U24012 (N_24012,N_14337,N_12275);
xor U24013 (N_24013,N_18487,N_12562);
nor U24014 (N_24014,N_19915,N_12694);
or U24015 (N_24015,N_14221,N_15350);
and U24016 (N_24016,N_19262,N_18743);
or U24017 (N_24017,N_14927,N_13589);
nand U24018 (N_24018,N_17703,N_11141);
xor U24019 (N_24019,N_11759,N_19899);
nand U24020 (N_24020,N_19560,N_12594);
or U24021 (N_24021,N_12643,N_15191);
nand U24022 (N_24022,N_17224,N_16198);
or U24023 (N_24023,N_16753,N_10883);
xor U24024 (N_24024,N_14078,N_11999);
or U24025 (N_24025,N_15327,N_18521);
or U24026 (N_24026,N_13918,N_12504);
nand U24027 (N_24027,N_18317,N_10155);
and U24028 (N_24028,N_18564,N_13190);
nand U24029 (N_24029,N_17190,N_11380);
xnor U24030 (N_24030,N_15562,N_13496);
or U24031 (N_24031,N_18005,N_17473);
nand U24032 (N_24032,N_12555,N_12546);
and U24033 (N_24033,N_14691,N_15566);
nand U24034 (N_24034,N_16329,N_17819);
nor U24035 (N_24035,N_17722,N_13540);
nand U24036 (N_24036,N_10638,N_13981);
or U24037 (N_24037,N_15937,N_18099);
nor U24038 (N_24038,N_17202,N_11090);
nor U24039 (N_24039,N_17793,N_11102);
nand U24040 (N_24040,N_16046,N_18812);
nor U24041 (N_24041,N_19506,N_11363);
nand U24042 (N_24042,N_10887,N_18221);
xor U24043 (N_24043,N_12968,N_13136);
nor U24044 (N_24044,N_12126,N_12139);
nor U24045 (N_24045,N_12458,N_10989);
or U24046 (N_24046,N_18792,N_15865);
xnor U24047 (N_24047,N_15613,N_18457);
xnor U24048 (N_24048,N_10341,N_18584);
nor U24049 (N_24049,N_17492,N_15168);
nor U24050 (N_24050,N_10421,N_14197);
and U24051 (N_24051,N_10097,N_13549);
xor U24052 (N_24052,N_19730,N_17694);
nor U24053 (N_24053,N_16979,N_10490);
or U24054 (N_24054,N_18306,N_11323);
nor U24055 (N_24055,N_19958,N_13934);
or U24056 (N_24056,N_16605,N_11069);
nand U24057 (N_24057,N_17691,N_11607);
nand U24058 (N_24058,N_16401,N_19661);
xor U24059 (N_24059,N_11354,N_17619);
nor U24060 (N_24060,N_11807,N_10470);
or U24061 (N_24061,N_15728,N_19930);
and U24062 (N_24062,N_12893,N_10985);
xnor U24063 (N_24063,N_16372,N_19572);
and U24064 (N_24064,N_12150,N_11455);
and U24065 (N_24065,N_16817,N_19406);
or U24066 (N_24066,N_14238,N_10746);
xnor U24067 (N_24067,N_11839,N_17186);
and U24068 (N_24068,N_15695,N_10914);
xor U24069 (N_24069,N_12615,N_12372);
xnor U24070 (N_24070,N_13479,N_10606);
xnor U24071 (N_24071,N_10112,N_14100);
nor U24072 (N_24072,N_10933,N_12135);
and U24073 (N_24073,N_11504,N_12097);
nor U24074 (N_24074,N_13172,N_14216);
or U24075 (N_24075,N_16636,N_15915);
nand U24076 (N_24076,N_17039,N_18347);
or U24077 (N_24077,N_16798,N_15631);
nor U24078 (N_24078,N_11115,N_15485);
nor U24079 (N_24079,N_13289,N_16822);
nor U24080 (N_24080,N_16940,N_11205);
xor U24081 (N_24081,N_15455,N_11816);
or U24082 (N_24082,N_12296,N_17816);
and U24083 (N_24083,N_16919,N_12389);
nand U24084 (N_24084,N_16310,N_12397);
nor U24085 (N_24085,N_10333,N_13586);
or U24086 (N_24086,N_11336,N_18450);
nor U24087 (N_24087,N_15049,N_18145);
nor U24088 (N_24088,N_10327,N_13713);
or U24089 (N_24089,N_15861,N_15622);
nor U24090 (N_24090,N_12014,N_12212);
nand U24091 (N_24091,N_16731,N_17274);
or U24092 (N_24092,N_11867,N_14454);
xnor U24093 (N_24093,N_13939,N_19826);
nand U24094 (N_24094,N_11171,N_16300);
and U24095 (N_24095,N_11248,N_11365);
nand U24096 (N_24096,N_18101,N_13749);
nor U24097 (N_24097,N_14529,N_14381);
xor U24098 (N_24098,N_13464,N_10576);
xor U24099 (N_24099,N_10945,N_16560);
nor U24100 (N_24100,N_10378,N_14659);
nand U24101 (N_24101,N_14303,N_12186);
nor U24102 (N_24102,N_11034,N_17118);
or U24103 (N_24103,N_14310,N_11463);
and U24104 (N_24104,N_18066,N_18900);
xor U24105 (N_24105,N_10961,N_19567);
and U24106 (N_24106,N_18654,N_10275);
xor U24107 (N_24107,N_17443,N_14490);
and U24108 (N_24108,N_19407,N_13993);
nand U24109 (N_24109,N_15803,N_16968);
nor U24110 (N_24110,N_16156,N_10910);
nor U24111 (N_24111,N_17230,N_14259);
nand U24112 (N_24112,N_17155,N_11768);
xor U24113 (N_24113,N_13996,N_10181);
and U24114 (N_24114,N_10478,N_13770);
and U24115 (N_24115,N_14579,N_12739);
nor U24116 (N_24116,N_11552,N_10430);
nand U24117 (N_24117,N_15785,N_18494);
nand U24118 (N_24118,N_13592,N_18790);
and U24119 (N_24119,N_11457,N_18493);
nand U24120 (N_24120,N_19769,N_10541);
nand U24121 (N_24121,N_15237,N_10274);
and U24122 (N_24122,N_17050,N_17347);
xnor U24123 (N_24123,N_14732,N_17046);
or U24124 (N_24124,N_11687,N_17093);
xor U24125 (N_24125,N_12846,N_17354);
nand U24126 (N_24126,N_11730,N_17149);
nor U24127 (N_24127,N_19447,N_15244);
or U24128 (N_24128,N_19261,N_14569);
and U24129 (N_24129,N_15982,N_13331);
or U24130 (N_24130,N_11296,N_15520);
xor U24131 (N_24131,N_19498,N_14550);
xor U24132 (N_24132,N_17464,N_10924);
nor U24133 (N_24133,N_19441,N_19358);
nor U24134 (N_24134,N_14435,N_15128);
nand U24135 (N_24135,N_14276,N_16470);
or U24136 (N_24136,N_16072,N_17010);
nor U24137 (N_24137,N_15983,N_14808);
or U24138 (N_24138,N_13215,N_15500);
or U24139 (N_24139,N_10814,N_11043);
nor U24140 (N_24140,N_17993,N_17030);
nor U24141 (N_24141,N_11244,N_16790);
xor U24142 (N_24142,N_14993,N_13787);
or U24143 (N_24143,N_15330,N_12346);
or U24144 (N_24144,N_14382,N_19381);
nor U24145 (N_24145,N_14291,N_16997);
and U24146 (N_24146,N_18434,N_10077);
xor U24147 (N_24147,N_16309,N_17402);
nand U24148 (N_24148,N_18964,N_19125);
nor U24149 (N_24149,N_19710,N_13556);
or U24150 (N_24150,N_10270,N_15966);
nor U24151 (N_24151,N_17013,N_19775);
nand U24152 (N_24152,N_10536,N_12510);
and U24153 (N_24153,N_16895,N_13401);
or U24154 (N_24154,N_16286,N_15488);
xnor U24155 (N_24155,N_16001,N_18313);
or U24156 (N_24156,N_19759,N_12038);
and U24157 (N_24157,N_13858,N_19840);
or U24158 (N_24158,N_19228,N_14048);
nor U24159 (N_24159,N_12436,N_19647);
or U24160 (N_24160,N_16885,N_17396);
xnor U24161 (N_24161,N_17714,N_10547);
or U24162 (N_24162,N_16392,N_13390);
nand U24163 (N_24163,N_17032,N_12626);
and U24164 (N_24164,N_18341,N_15895);
xor U24165 (N_24165,N_11941,N_17004);
or U24166 (N_24166,N_17992,N_17845);
xnor U24167 (N_24167,N_14122,N_12277);
nor U24168 (N_24168,N_17314,N_15859);
xnor U24169 (N_24169,N_19984,N_16917);
or U24170 (N_24170,N_11834,N_16715);
and U24171 (N_24171,N_15614,N_18152);
nand U24172 (N_24172,N_10009,N_18747);
nor U24173 (N_24173,N_15092,N_16444);
or U24174 (N_24174,N_17390,N_13865);
or U24175 (N_24175,N_10324,N_10476);
or U24176 (N_24176,N_15567,N_19047);
and U24177 (N_24177,N_13902,N_17987);
or U24178 (N_24178,N_18060,N_13644);
xnor U24179 (N_24179,N_13609,N_19451);
nor U24180 (N_24180,N_18837,N_11159);
or U24181 (N_24181,N_19650,N_16207);
and U24182 (N_24182,N_17493,N_17835);
nor U24183 (N_24183,N_19123,N_15651);
and U24184 (N_24184,N_18813,N_18157);
and U24185 (N_24185,N_18963,N_19937);
nor U24186 (N_24186,N_15909,N_14133);
nand U24187 (N_24187,N_15036,N_19979);
and U24188 (N_24188,N_14302,N_13652);
and U24189 (N_24189,N_11525,N_10312);
nand U24190 (N_24190,N_17122,N_10770);
or U24191 (N_24191,N_12661,N_12070);
nor U24192 (N_24192,N_12024,N_12323);
or U24193 (N_24193,N_17878,N_11064);
or U24194 (N_24194,N_17575,N_13949);
or U24195 (N_24195,N_13505,N_16902);
xor U24196 (N_24196,N_16223,N_16702);
and U24197 (N_24197,N_12891,N_17966);
or U24198 (N_24198,N_19959,N_16028);
or U24199 (N_24199,N_18692,N_12704);
and U24200 (N_24200,N_10530,N_16379);
nor U24201 (N_24201,N_11328,N_18137);
nor U24202 (N_24202,N_18035,N_16526);
nor U24203 (N_24203,N_11105,N_13728);
nor U24204 (N_24204,N_10357,N_10309);
and U24205 (N_24205,N_19643,N_18387);
nand U24206 (N_24206,N_13651,N_15781);
nor U24207 (N_24207,N_12561,N_16663);
nor U24208 (N_24208,N_11567,N_17421);
nand U24209 (N_24209,N_10843,N_12179);
nor U24210 (N_24210,N_10921,N_10448);
nand U24211 (N_24211,N_15018,N_10545);
nor U24212 (N_24212,N_11558,N_15599);
or U24213 (N_24213,N_12147,N_16130);
nand U24214 (N_24214,N_16431,N_11593);
xnor U24215 (N_24215,N_12878,N_11961);
xnor U24216 (N_24216,N_18396,N_17124);
or U24217 (N_24217,N_12176,N_17018);
and U24218 (N_24218,N_13765,N_17660);
nand U24219 (N_24219,N_15924,N_16253);
and U24220 (N_24220,N_14868,N_15932);
nand U24221 (N_24221,N_12045,N_19804);
nor U24222 (N_24222,N_16482,N_11910);
xnor U24223 (N_24223,N_16531,N_15429);
nor U24224 (N_24224,N_10227,N_12605);
or U24225 (N_24225,N_18899,N_11004);
nand U24226 (N_24226,N_15649,N_12309);
and U24227 (N_24227,N_10467,N_10647);
or U24228 (N_24228,N_17524,N_12262);
or U24229 (N_24229,N_18528,N_14274);
nand U24230 (N_24230,N_11191,N_12508);
xnor U24231 (N_24231,N_15636,N_18995);
xor U24232 (N_24232,N_18258,N_17678);
or U24233 (N_24233,N_19987,N_15538);
or U24234 (N_24234,N_13788,N_19808);
nand U24235 (N_24235,N_15316,N_10330);
xnor U24236 (N_24236,N_12907,N_19653);
nor U24237 (N_24237,N_17185,N_11720);
xor U24238 (N_24238,N_17977,N_12623);
nor U24239 (N_24239,N_17427,N_17361);
nor U24240 (N_24240,N_11106,N_11183);
nor U24241 (N_24241,N_18230,N_18614);
and U24242 (N_24242,N_15024,N_10603);
nor U24243 (N_24243,N_18148,N_17808);
and U24244 (N_24244,N_18130,N_19243);
and U24245 (N_24245,N_19322,N_11919);
nand U24246 (N_24246,N_10691,N_17785);
nor U24247 (N_24247,N_16126,N_10782);
xnor U24248 (N_24248,N_13105,N_19562);
and U24249 (N_24249,N_13880,N_19485);
xnor U24250 (N_24250,N_12782,N_16662);
xnor U24251 (N_24251,N_18159,N_10813);
nor U24252 (N_24252,N_16513,N_14060);
xnor U24253 (N_24253,N_19895,N_10138);
nor U24254 (N_24254,N_12110,N_10787);
or U24255 (N_24255,N_14718,N_14862);
or U24256 (N_24256,N_16889,N_18870);
xor U24257 (N_24257,N_19090,N_14107);
nand U24258 (N_24258,N_15660,N_18626);
or U24259 (N_24259,N_11618,N_17712);
and U24260 (N_24260,N_11879,N_18975);
or U24261 (N_24261,N_16176,N_14886);
nand U24262 (N_24262,N_17807,N_16159);
nor U24263 (N_24263,N_17918,N_14285);
nor U24264 (N_24264,N_10901,N_13640);
xor U24265 (N_24265,N_16412,N_13176);
and U24266 (N_24266,N_13269,N_14658);
xor U24267 (N_24267,N_15819,N_13731);
or U24268 (N_24268,N_12984,N_14906);
and U24269 (N_24269,N_17901,N_16096);
or U24270 (N_24270,N_12382,N_11909);
nor U24271 (N_24271,N_17130,N_18088);
xor U24272 (N_24272,N_17221,N_12494);
and U24273 (N_24273,N_16284,N_17160);
xor U24274 (N_24274,N_10471,N_10056);
and U24275 (N_24275,N_15444,N_12237);
nor U24276 (N_24276,N_19121,N_11147);
nand U24277 (N_24277,N_16059,N_12728);
or U24278 (N_24278,N_17943,N_18984);
nor U24279 (N_24279,N_15042,N_12666);
nor U24280 (N_24280,N_13011,N_19781);
and U24281 (N_24281,N_11283,N_18466);
xnor U24282 (N_24282,N_10807,N_18735);
xnor U24283 (N_24283,N_15321,N_10276);
xnor U24284 (N_24284,N_12394,N_11417);
nor U24285 (N_24285,N_18998,N_17612);
nor U24286 (N_24286,N_12477,N_18282);
or U24287 (N_24287,N_13029,N_12864);
xor U24288 (N_24288,N_11899,N_19029);
nor U24289 (N_24289,N_15721,N_10863);
nand U24290 (N_24290,N_17567,N_15255);
nand U24291 (N_24291,N_11347,N_10712);
and U24292 (N_24292,N_12155,N_19537);
or U24293 (N_24293,N_10415,N_14148);
or U24294 (N_24294,N_19477,N_10998);
nand U24295 (N_24295,N_16171,N_14813);
nor U24296 (N_24296,N_15421,N_15352);
xnor U24297 (N_24297,N_14452,N_18580);
nor U24298 (N_24298,N_14509,N_14057);
nor U24299 (N_24299,N_18092,N_18422);
xor U24300 (N_24300,N_16911,N_17412);
and U24301 (N_24301,N_19320,N_13125);
or U24302 (N_24302,N_11349,N_10953);
nor U24303 (N_24303,N_12928,N_17379);
nand U24304 (N_24304,N_12344,N_10427);
xnor U24305 (N_24305,N_11739,N_15884);
and U24306 (N_24306,N_11215,N_16098);
nor U24307 (N_24307,N_16945,N_15235);
or U24308 (N_24308,N_11176,N_10195);
nor U24309 (N_24309,N_18828,N_12108);
nand U24310 (N_24310,N_16915,N_10054);
or U24311 (N_24311,N_11578,N_19380);
and U24312 (N_24312,N_19884,N_12076);
or U24313 (N_24313,N_16466,N_17269);
or U24314 (N_24314,N_16282,N_14217);
xnor U24315 (N_24315,N_14807,N_14032);
nor U24316 (N_24316,N_14171,N_15006);
or U24317 (N_24317,N_14667,N_18849);
nor U24318 (N_24318,N_17408,N_14374);
and U24319 (N_24319,N_12868,N_12379);
and U24320 (N_24320,N_19200,N_18794);
or U24321 (N_24321,N_11784,N_14049);
or U24322 (N_24322,N_17635,N_12054);
or U24323 (N_24323,N_15135,N_12031);
nor U24324 (N_24324,N_13487,N_11847);
or U24325 (N_24325,N_11104,N_10876);
xnor U24326 (N_24326,N_11665,N_16590);
nand U24327 (N_24327,N_19435,N_13052);
xor U24328 (N_24328,N_11145,N_13525);
and U24329 (N_24329,N_18224,N_15786);
xnor U24330 (N_24330,N_18820,N_11413);
nand U24331 (N_24331,N_14751,N_13781);
and U24332 (N_24332,N_12364,N_19446);
or U24333 (N_24333,N_17554,N_19157);
or U24334 (N_24334,N_17193,N_14885);
nand U24335 (N_24335,N_16213,N_17698);
and U24336 (N_24336,N_16576,N_13448);
or U24337 (N_24337,N_18213,N_10908);
nor U24338 (N_24338,N_12904,N_11172);
or U24339 (N_24339,N_16090,N_15118);
nor U24340 (N_24340,N_17455,N_16487);
nand U24341 (N_24341,N_19977,N_15620);
or U24342 (N_24342,N_10719,N_15041);
or U24343 (N_24343,N_13785,N_16928);
xor U24344 (N_24344,N_12639,N_12197);
nor U24345 (N_24345,N_13498,N_10566);
or U24346 (N_24346,N_12899,N_16640);
nor U24347 (N_24347,N_10348,N_16115);
nor U24348 (N_24348,N_12691,N_17267);
nand U24349 (N_24349,N_18509,N_16339);
nand U24350 (N_24350,N_14695,N_11282);
or U24351 (N_24351,N_18123,N_13142);
xnor U24352 (N_24352,N_10306,N_13271);
nor U24353 (N_24353,N_18102,N_14547);
xor U24354 (N_24354,N_14093,N_18272);
xor U24355 (N_24355,N_12973,N_16233);
or U24356 (N_24356,N_18881,N_12887);
nor U24357 (N_24357,N_19603,N_12741);
or U24358 (N_24358,N_12536,N_10153);
nand U24359 (N_24359,N_14398,N_12206);
or U24360 (N_24360,N_19570,N_13877);
xnor U24361 (N_24361,N_12624,N_14261);
and U24362 (N_24362,N_13567,N_19712);
xor U24363 (N_24363,N_11133,N_13814);
nand U24364 (N_24364,N_19810,N_10736);
or U24365 (N_24365,N_14716,N_11940);
and U24366 (N_24366,N_18049,N_10425);
xor U24367 (N_24367,N_13629,N_14514);
or U24368 (N_24368,N_12486,N_13655);
nor U24369 (N_24369,N_11701,N_19221);
xnor U24370 (N_24370,N_12737,N_18540);
nand U24371 (N_24371,N_19324,N_16117);
nand U24372 (N_24372,N_14576,N_18323);
xor U24373 (N_24373,N_12909,N_13834);
nor U24374 (N_24374,N_10459,N_14260);
and U24375 (N_24375,N_16359,N_12332);
or U24376 (N_24376,N_19345,N_11508);
nor U24377 (N_24377,N_15100,N_11642);
xnor U24378 (N_24378,N_10780,N_16948);
xnor U24379 (N_24379,N_14515,N_14777);
and U24380 (N_24380,N_16026,N_19549);
and U24381 (N_24381,N_11575,N_10132);
and U24382 (N_24382,N_12283,N_17410);
nand U24383 (N_24383,N_19832,N_13759);
nor U24384 (N_24384,N_11636,N_14247);
nand U24385 (N_24385,N_16062,N_16222);
nand U24386 (N_24386,N_10987,N_13447);
or U24387 (N_24387,N_11850,N_19077);
xnor U24388 (N_24388,N_13522,N_10245);
or U24389 (N_24389,N_14810,N_16553);
and U24390 (N_24390,N_19971,N_10120);
xor U24391 (N_24391,N_17052,N_14000);
xor U24392 (N_24392,N_18697,N_19020);
xnor U24393 (N_24393,N_10635,N_16710);
or U24394 (N_24394,N_11845,N_12751);
nor U24395 (N_24395,N_19440,N_17169);
nand U24396 (N_24396,N_10694,N_13573);
nor U24397 (N_24397,N_11840,N_16728);
or U24398 (N_24398,N_10809,N_12911);
xnor U24399 (N_24399,N_12628,N_16921);
xor U24400 (N_24400,N_18424,N_12064);
nand U24401 (N_24401,N_17418,N_18644);
nand U24402 (N_24402,N_17581,N_14026);
and U24403 (N_24403,N_19163,N_19721);
nor U24404 (N_24404,N_13811,N_15551);
xor U24405 (N_24405,N_12180,N_14417);
xor U24406 (N_24406,N_15831,N_18453);
or U24407 (N_24407,N_12177,N_14201);
nand U24408 (N_24408,N_18572,N_15600);
or U24409 (N_24409,N_12125,N_12814);
nand U24410 (N_24410,N_16943,N_14482);
nor U24411 (N_24411,N_19122,N_17652);
nor U24412 (N_24412,N_12401,N_11087);
and U24413 (N_24413,N_14448,N_15701);
or U24414 (N_24414,N_13026,N_19331);
xnor U24415 (N_24415,N_18231,N_10250);
or U24416 (N_24416,N_13922,N_14922);
and U24417 (N_24417,N_11991,N_14466);
xor U24418 (N_24418,N_15716,N_15161);
or U24419 (N_24419,N_11917,N_14522);
nand U24420 (N_24420,N_12668,N_12678);
or U24421 (N_24421,N_15846,N_14357);
xor U24422 (N_24422,N_15712,N_17653);
nor U24423 (N_24423,N_19592,N_15275);
or U24424 (N_24424,N_17367,N_13454);
nand U24425 (N_24425,N_15574,N_19126);
nand U24426 (N_24426,N_18547,N_15912);
xor U24427 (N_24427,N_14170,N_19196);
or U24428 (N_24428,N_18470,N_15207);
xor U24429 (N_24429,N_17981,N_15860);
xnor U24430 (N_24430,N_14770,N_16049);
xnor U24431 (N_24431,N_14334,N_14528);
nand U24432 (N_24432,N_16354,N_17719);
and U24433 (N_24433,N_11197,N_11082);
nor U24434 (N_24434,N_11326,N_16982);
and U24435 (N_24435,N_12319,N_17060);
xor U24436 (N_24436,N_17585,N_12201);
and U24437 (N_24437,N_12478,N_14202);
nand U24438 (N_24438,N_19825,N_10655);
xor U24439 (N_24439,N_13866,N_19087);
nand U24440 (N_24440,N_17642,N_15635);
xor U24441 (N_24441,N_13846,N_18928);
xor U24442 (N_24442,N_12677,N_19690);
nand U24443 (N_24443,N_14552,N_12023);
or U24444 (N_24444,N_17809,N_16774);
nand U24445 (N_24445,N_12112,N_11648);
xor U24446 (N_24446,N_15748,N_12362);
nand U24447 (N_24447,N_17964,N_19839);
or U24448 (N_24448,N_14881,N_17496);
nor U24449 (N_24449,N_19420,N_12538);
or U24450 (N_24450,N_12106,N_18861);
and U24451 (N_24451,N_19272,N_13744);
or U24452 (N_24452,N_14760,N_10765);
or U24453 (N_24453,N_13735,N_12065);
and U24454 (N_24454,N_15410,N_17011);
and U24455 (N_24455,N_13953,N_17042);
or U24456 (N_24456,N_15351,N_14157);
and U24457 (N_24457,N_17298,N_18549);
nand U24458 (N_24458,N_11921,N_15094);
and U24459 (N_24459,N_14656,N_16497);
xor U24460 (N_24460,N_19412,N_12991);
and U24461 (N_24461,N_12414,N_18853);
xor U24462 (N_24462,N_16690,N_15159);
and U24463 (N_24463,N_19596,N_16607);
or U24464 (N_24464,N_17098,N_19568);
nor U24465 (N_24465,N_13402,N_12413);
nand U24466 (N_24466,N_15032,N_19716);
nor U24467 (N_24467,N_15504,N_16740);
or U24468 (N_24468,N_13110,N_10875);
or U24469 (N_24469,N_14236,N_19204);
nor U24470 (N_24470,N_10956,N_14015);
nand U24471 (N_24471,N_19980,N_12171);
nor U24472 (N_24472,N_19205,N_12803);
or U24473 (N_24473,N_10004,N_16319);
nand U24474 (N_24474,N_16969,N_17133);
nor U24475 (N_24475,N_15849,N_13526);
xnor U24476 (N_24476,N_16737,N_12897);
nor U24477 (N_24477,N_12100,N_16706);
nor U24478 (N_24478,N_11756,N_19479);
and U24479 (N_24479,N_13694,N_15261);
xor U24480 (N_24480,N_12303,N_19998);
xnor U24481 (N_24481,N_10417,N_16882);
nor U24482 (N_24482,N_10615,N_15751);
xnor U24483 (N_24483,N_13438,N_13482);
nand U24484 (N_24484,N_11083,N_18129);
or U24485 (N_24485,N_12755,N_13007);
xnor U24486 (N_24486,N_10944,N_13060);
nand U24487 (N_24487,N_18153,N_16074);
nand U24488 (N_24488,N_11307,N_13554);
xnor U24489 (N_24489,N_12784,N_16872);
xor U24490 (N_24490,N_17001,N_18107);
and U24491 (N_24491,N_17203,N_18806);
xor U24492 (N_24492,N_15610,N_17735);
or U24493 (N_24493,N_12424,N_16451);
or U24494 (N_24494,N_10443,N_14802);
and U24495 (N_24495,N_18705,N_12481);
or U24496 (N_24496,N_11237,N_18781);
nor U24497 (N_24497,N_12700,N_18990);
xor U24498 (N_24498,N_15642,N_19400);
nor U24499 (N_24499,N_16770,N_10210);
xnor U24500 (N_24500,N_17975,N_12399);
and U24501 (N_24501,N_14371,N_17860);
nand U24502 (N_24502,N_13183,N_13094);
or U24503 (N_24503,N_16099,N_15044);
xnor U24504 (N_24504,N_17498,N_15124);
nor U24505 (N_24505,N_15198,N_15724);
nor U24506 (N_24506,N_18462,N_14753);
xor U24507 (N_24507,N_18770,N_12250);
nor U24508 (N_24508,N_14191,N_11199);
nor U24509 (N_24509,N_18389,N_14244);
and U24510 (N_24510,N_15333,N_12879);
or U24511 (N_24511,N_15043,N_14895);
or U24512 (N_24512,N_14372,N_10016);
or U24513 (N_24513,N_12352,N_19986);
nand U24514 (N_24514,N_18255,N_16811);
nor U24515 (N_24515,N_11143,N_19177);
nor U24516 (N_24516,N_14893,N_11025);
xor U24517 (N_24517,N_14783,N_10757);
xor U24518 (N_24518,N_14676,N_14044);
nand U24519 (N_24519,N_13985,N_19364);
xnor U24520 (N_24520,N_12321,N_17951);
and U24521 (N_24521,N_12777,N_15753);
nor U24522 (N_24522,N_10496,N_19318);
or U24523 (N_24523,N_18764,N_11996);
xnor U24524 (N_24524,N_16480,N_17960);
or U24525 (N_24525,N_15502,N_10859);
nand U24526 (N_24526,N_18382,N_19737);
and U24527 (N_24527,N_11601,N_14289);
xor U24528 (N_24528,N_12488,N_19323);
or U24529 (N_24529,N_13997,N_17310);
and U24530 (N_24530,N_17593,N_16856);
xnor U24531 (N_24531,N_12059,N_16437);
or U24532 (N_24532,N_10237,N_16205);
xnor U24533 (N_24533,N_15767,N_14632);
or U24534 (N_24534,N_14254,N_14379);
xnor U24535 (N_24535,N_16230,N_10334);
or U24536 (N_24536,N_14313,N_14979);
nand U24537 (N_24537,N_12121,N_16069);
xnor U24538 (N_24538,N_16719,N_11423);
nor U24539 (N_24539,N_14195,N_10460);
and U24540 (N_24540,N_15887,N_18518);
nor U24541 (N_24541,N_15326,N_15719);
nand U24542 (N_24542,N_15079,N_10063);
and U24543 (N_24543,N_18511,N_13551);
xor U24544 (N_24544,N_19067,N_12788);
xor U24545 (N_24545,N_19285,N_16396);
nand U24546 (N_24546,N_10396,N_11498);
nor U24547 (N_24547,N_17577,N_14301);
xor U24548 (N_24548,N_19283,N_11670);
nor U24549 (N_24549,N_11315,N_14222);
xor U24550 (N_24550,N_12634,N_18609);
xnor U24551 (N_24551,N_18057,N_11072);
or U24552 (N_24552,N_14384,N_10800);
and U24553 (N_24553,N_11000,N_13389);
nand U24554 (N_24554,N_19340,N_16113);
xnor U24555 (N_24555,N_19798,N_19799);
nor U24556 (N_24556,N_12052,N_15291);
and U24557 (N_24557,N_15312,N_13620);
and U24558 (N_24558,N_16500,N_13509);
nor U24559 (N_24559,N_16601,N_11291);
xor U24560 (N_24560,N_14018,N_16358);
nor U24561 (N_24561,N_11421,N_17363);
nor U24562 (N_24562,N_13748,N_13164);
nand U24563 (N_24563,N_16718,N_18668);
nor U24564 (N_24564,N_10596,N_14296);
xnor U24565 (N_24565,N_19254,N_10057);
nor U24566 (N_24566,N_17233,N_10903);
or U24567 (N_24567,N_15126,N_18576);
xor U24568 (N_24568,N_15935,N_11267);
xnor U24569 (N_24569,N_16581,N_18120);
or U24570 (N_24570,N_11490,N_12022);
and U24571 (N_24571,N_15524,N_18244);
nand U24572 (N_24572,N_11963,N_19517);
nor U24573 (N_24573,N_15740,N_19117);
nand U24574 (N_24574,N_17531,N_17590);
nor U24575 (N_24575,N_10503,N_15492);
or U24576 (N_24576,N_11745,N_19244);
nand U24577 (N_24577,N_16071,N_18324);
nor U24578 (N_24578,N_11209,N_19146);
nand U24579 (N_24579,N_19723,N_11442);
nor U24580 (N_24580,N_12493,N_10667);
nor U24581 (N_24581,N_17323,N_18023);
and U24582 (N_24582,N_15477,N_10659);
nor U24583 (N_24583,N_12360,N_15274);
and U24584 (N_24584,N_10717,N_19739);
nand U24585 (N_24585,N_19236,N_17163);
or U24586 (N_24586,N_12016,N_14897);
xnor U24587 (N_24587,N_18239,N_18643);
xor U24588 (N_24588,N_11655,N_19137);
nand U24589 (N_24589,N_14199,N_19755);
nor U24590 (N_24590,N_14059,N_19540);
nand U24591 (N_24591,N_12502,N_10273);
and U24592 (N_24592,N_18081,N_16587);
nor U24593 (N_24593,N_16966,N_16762);
and U24594 (N_24594,N_16267,N_17070);
nand U24595 (N_24595,N_11428,N_14709);
xnor U24596 (N_24596,N_16350,N_15190);
nor U24597 (N_24597,N_11318,N_17405);
nor U24598 (N_24598,N_18886,N_12731);
nand U24599 (N_24599,N_11762,N_11398);
nor U24600 (N_24600,N_12058,N_16647);
nor U24601 (N_24601,N_12690,N_17775);
xnor U24602 (N_24602,N_16648,N_13669);
and U24603 (N_24603,N_15880,N_13206);
xor U24604 (N_24604,N_17016,N_10760);
and U24605 (N_24605,N_18243,N_14969);
or U24606 (N_24606,N_11488,N_16292);
or U24607 (N_24607,N_15643,N_17837);
nor U24608 (N_24608,N_17342,N_16652);
nand U24609 (N_24609,N_13426,N_17849);
and U24610 (N_24610,N_16756,N_12706);
xor U24611 (N_24611,N_14376,N_13704);
and U24612 (N_24612,N_15259,N_15809);
and U24613 (N_24613,N_14657,N_10280);
nand U24614 (N_24614,N_16671,N_18138);
and U24615 (N_24615,N_16160,N_18602);
and U24616 (N_24616,N_16100,N_10893);
or U24617 (N_24617,N_15933,N_18620);
and U24618 (N_24618,N_14913,N_12077);
nand U24619 (N_24619,N_19208,N_14146);
or U24620 (N_24620,N_17909,N_12660);
nor U24621 (N_24621,N_15833,N_11968);
and U24622 (N_24622,N_18562,N_15994);
nor U24623 (N_24623,N_18502,N_12337);
nand U24624 (N_24624,N_18877,N_12249);
and U24625 (N_24625,N_11373,N_11431);
nor U24626 (N_24626,N_17658,N_14101);
and U24627 (N_24627,N_16219,N_19338);
nand U24628 (N_24628,N_17644,N_15796);
or U24629 (N_24629,N_11993,N_15022);
xnor U24630 (N_24630,N_14591,N_10852);
nand U24631 (N_24631,N_13951,N_14797);
and U24632 (N_24632,N_19415,N_17767);
nor U24633 (N_24633,N_18824,N_10222);
xnor U24634 (N_24634,N_13287,N_12430);
nor U24635 (N_24635,N_18937,N_16427);
nand U24636 (N_24636,N_12701,N_12827);
nor U24637 (N_24637,N_13336,N_16631);
nand U24638 (N_24638,N_18690,N_19527);
nand U24639 (N_24639,N_17745,N_10657);
and U24640 (N_24640,N_15468,N_11249);
nand U24641 (N_24641,N_19378,N_16900);
nor U24642 (N_24642,N_12505,N_14118);
or U24643 (N_24643,N_13769,N_10683);
or U24644 (N_24644,N_15885,N_14574);
or U24645 (N_24645,N_12919,N_18122);
xnor U24646 (N_24646,N_13302,N_12716);
nand U24647 (N_24647,N_17972,N_13492);
or U24648 (N_24648,N_17917,N_10904);
xnor U24649 (N_24649,N_12255,N_11891);
nand U24650 (N_24650,N_17246,N_18180);
or U24651 (N_24651,N_10865,N_19482);
or U24652 (N_24652,N_11078,N_18866);
nand U24653 (N_24653,N_15095,N_15806);
nor U24654 (N_24654,N_15762,N_17605);
nand U24655 (N_24655,N_11013,N_17958);
nand U24656 (N_24656,N_16720,N_14173);
nand U24657 (N_24657,N_16481,N_19866);
nand U24658 (N_24658,N_18398,N_14356);
and U24659 (N_24659,N_12881,N_13776);
nor U24660 (N_24660,N_11162,N_15474);
and U24661 (N_24661,N_18301,N_15690);
nor U24662 (N_24662,N_11453,N_17422);
nor U24663 (N_24663,N_16907,N_10758);
and U24664 (N_24664,N_14265,N_17823);
or U24665 (N_24665,N_12528,N_14630);
or U24666 (N_24666,N_11714,N_16163);
or U24667 (N_24667,N_14029,N_13257);
xnor U24668 (N_24668,N_17102,N_17776);
and U24669 (N_24669,N_18725,N_16192);
xnor U24670 (N_24670,N_11489,N_18350);
or U24671 (N_24671,N_12267,N_15676);
nand U24672 (N_24672,N_14698,N_12306);
nor U24673 (N_24673,N_18591,N_12910);
or U24674 (N_24674,N_12091,N_16927);
nor U24675 (N_24675,N_15315,N_10393);
nor U24676 (N_24676,N_18245,N_17515);
nor U24677 (N_24677,N_19513,N_16825);
nor U24678 (N_24678,N_15219,N_11591);
or U24679 (N_24679,N_12906,N_13366);
and U24680 (N_24680,N_13310,N_12033);
nand U24681 (N_24681,N_15320,N_12443);
xnor U24682 (N_24682,N_19300,N_13320);
xor U24683 (N_24683,N_11754,N_18920);
or U24684 (N_24684,N_11667,N_16370);
xnor U24685 (N_24685,N_17768,N_17826);
or U24686 (N_24686,N_17862,N_13582);
nand U24687 (N_24687,N_18497,N_19757);
nor U24688 (N_24688,N_10790,N_15637);
nor U24689 (N_24689,N_19910,N_16052);
xor U24690 (N_24690,N_19316,N_13330);
nand U24691 (N_24691,N_16277,N_19038);
nor U24692 (N_24692,N_14898,N_10192);
nor U24693 (N_24693,N_10081,N_14846);
xnor U24694 (N_24694,N_14385,N_19542);
and U24695 (N_24695,N_18196,N_10564);
nand U24696 (N_24696,N_12710,N_18197);
nand U24697 (N_24697,N_16399,N_16537);
and U24698 (N_24698,N_13741,N_19282);
nor U24699 (N_24699,N_19639,N_10382);
nand U24700 (N_24700,N_10802,N_14948);
and U24701 (N_24701,N_11376,N_17428);
or U24702 (N_24702,N_16058,N_13484);
xor U24703 (N_24703,N_11889,N_15822);
nand U24704 (N_24704,N_18452,N_14208);
xnor U24705 (N_24705,N_19641,N_14097);
nand U24706 (N_24706,N_10482,N_10265);
or U24707 (N_24707,N_11666,N_19198);
nand U24708 (N_24708,N_12498,N_12783);
nor U24709 (N_24709,N_11528,N_18848);
and U24710 (N_24710,N_14324,N_11005);
nand U24711 (N_24711,N_18257,N_19615);
xnor U24712 (N_24712,N_19066,N_13422);
nand U24713 (N_24713,N_12348,N_15706);
nor U24714 (N_24714,N_14293,N_11707);
nand U24715 (N_24715,N_15595,N_17935);
nor U24716 (N_24716,N_18941,N_13365);
or U24717 (N_24717,N_13754,N_10402);
and U24718 (N_24718,N_19746,N_15133);
or U24719 (N_24719,N_19105,N_18048);
or U24720 (N_24720,N_16410,N_19834);
and U24721 (N_24721,N_18986,N_18538);
nand U24722 (N_24722,N_11703,N_14826);
xor U24723 (N_24723,N_16002,N_13685);
or U24724 (N_24724,N_10873,N_17979);
nor U24725 (N_24725,N_19846,N_14277);
and U24726 (N_24726,N_18809,N_11812);
nand U24727 (N_24727,N_16200,N_12558);
xnor U24728 (N_24728,N_13411,N_15518);
or U24729 (N_24729,N_13015,N_15138);
nand U24730 (N_24730,N_16714,N_13427);
or U24731 (N_24731,N_10862,N_14767);
and U24732 (N_24732,N_14483,N_14778);
xnor U24733 (N_24733,N_14408,N_16591);
and U24734 (N_24734,N_14227,N_17507);
or U24735 (N_24735,N_10354,N_14024);
nor U24736 (N_24736,N_16511,N_12000);
xor U24737 (N_24737,N_18512,N_14645);
xnor U24738 (N_24738,N_14809,N_18529);
nand U24739 (N_24739,N_10928,N_15389);
and U24740 (N_24740,N_12681,N_10507);
and U24741 (N_24741,N_15545,N_16337);
xor U24742 (N_24742,N_12977,N_10268);
xor U24743 (N_24743,N_10075,N_19830);
xnor U24744 (N_24744,N_17611,N_13109);
nor U24745 (N_24745,N_13340,N_10399);
nand U24746 (N_24746,N_13763,N_12548);
nand U24747 (N_24747,N_19281,N_10184);
and U24748 (N_24748,N_11230,N_10432);
nor U24749 (N_24749,N_18670,N_13947);
nor U24750 (N_24750,N_12438,N_17530);
or U24751 (N_24751,N_10968,N_17517);
xnor U24752 (N_24752,N_14022,N_12699);
and U24753 (N_24753,N_19478,N_19554);
or U24754 (N_24754,N_15234,N_13258);
nor U24755 (N_24755,N_15795,N_10796);
nand U24756 (N_24756,N_16322,N_12152);
xnor U24757 (N_24757,N_14794,N_14589);
nand U24758 (N_24758,N_10047,N_18730);
xnor U24759 (N_24759,N_17959,N_10793);
nand U24760 (N_24760,N_10590,N_11873);
nor U24761 (N_24761,N_11644,N_16195);
nor U24762 (N_24762,N_13162,N_16227);
and U24763 (N_24763,N_11793,N_10318);
xnor U24764 (N_24764,N_10990,N_10100);
and U24765 (N_24765,N_16317,N_10105);
and U24766 (N_24766,N_11252,N_13137);
xor U24767 (N_24767,N_17324,N_19869);
nand U24768 (N_24768,N_18797,N_13020);
nor U24769 (N_24769,N_19462,N_19881);
nor U24770 (N_24770,N_15571,N_19110);
nor U24771 (N_24771,N_18772,N_18722);
or U24772 (N_24772,N_10062,N_18233);
xor U24773 (N_24773,N_15059,N_13170);
xor U24774 (N_24774,N_19921,N_19978);
xor U24775 (N_24775,N_14958,N_16523);
nor U24776 (N_24776,N_13931,N_18163);
xnor U24777 (N_24777,N_13283,N_17215);
xnor U24778 (N_24778,N_17713,N_16736);
xor U24779 (N_24779,N_10747,N_16974);
nand U24780 (N_24780,N_17002,N_18443);
nand U24781 (N_24781,N_15624,N_16955);
xnor U24782 (N_24782,N_14231,N_10216);
xor U24783 (N_24783,N_15618,N_10702);
xor U24784 (N_24784,N_12252,N_13358);
xnor U24785 (N_24785,N_10772,N_15078);
and U24786 (N_24786,N_19523,N_11832);
nand U24787 (N_24787,N_12500,N_14803);
xor U24788 (N_24788,N_16660,N_11387);
and U24789 (N_24789,N_16681,N_18315);
nand U24790 (N_24790,N_13373,N_12532);
and U24791 (N_24791,N_14068,N_18829);
or U24792 (N_24792,N_17986,N_15824);
nand U24793 (N_24793,N_14560,N_12300);
and U24794 (N_24794,N_19843,N_17090);
xnor U24795 (N_24795,N_19049,N_12030);
nor U24796 (N_24796,N_11743,N_16307);
xnor U24797 (N_24797,N_19172,N_13708);
or U24798 (N_24798,N_18762,N_19416);
nand U24799 (N_24799,N_10735,N_17873);
nand U24800 (N_24800,N_14542,N_19886);
nand U24801 (N_24801,N_18666,N_19031);
or U24802 (N_24802,N_17213,N_16769);
nand U24803 (N_24803,N_11362,N_11998);
xor U24804 (N_24804,N_12732,N_14961);
or U24805 (N_24805,N_18524,N_16043);
or U24806 (N_24806,N_18675,N_10186);
or U24807 (N_24807,N_14328,N_17103);
xnor U24808 (N_24808,N_16677,N_11712);
nand U24809 (N_24809,N_12387,N_12888);
or U24810 (N_24810,N_11243,N_10067);
and U24811 (N_24811,N_15412,N_11672);
nor U24812 (N_24812,N_13897,N_18013);
or U24813 (N_24813,N_18442,N_17889);
nand U24814 (N_24814,N_17425,N_14135);
or U24815 (N_24815,N_18093,N_16914);
and U24816 (N_24816,N_10043,N_11938);
nor U24817 (N_24817,N_19104,N_14460);
nor U24818 (N_24818,N_14962,N_15763);
or U24819 (N_24819,N_12855,N_11019);
xnor U24820 (N_24820,N_16861,N_13499);
nor U24821 (N_24821,N_14071,N_14976);
nor U24822 (N_24822,N_17636,N_12885);
or U24823 (N_24823,N_15710,N_13450);
xor U24824 (N_24824,N_12258,N_12455);
and U24825 (N_24825,N_15640,N_17963);
xor U24826 (N_24826,N_15355,N_15973);
nor U24827 (N_24827,N_16931,N_17447);
nor U24828 (N_24828,N_17304,N_12384);
and U24829 (N_24829,N_11653,N_11028);
or U24830 (N_24830,N_14040,N_18296);
nand U24831 (N_24831,N_16031,N_15704);
nand U24832 (N_24832,N_10049,N_18923);
and U24833 (N_24833,N_17638,N_14655);
nand U24834 (N_24834,N_17008,N_10136);
and U24835 (N_24835,N_18556,N_16301);
and U24836 (N_24836,N_14304,N_11256);
nor U24837 (N_24837,N_19194,N_13802);
xor U24838 (N_24838,N_15917,N_14354);
xnor U24839 (N_24839,N_13691,N_13965);
or U24840 (N_24840,N_16838,N_10869);
xnor U24841 (N_24841,N_10522,N_15017);
xor U24842 (N_24842,N_16995,N_18822);
xnor U24843 (N_24843,N_19043,N_13117);
and U24844 (N_24844,N_19752,N_12153);
and U24845 (N_24845,N_19555,N_19576);
or U24846 (N_24846,N_17089,N_11262);
or U24847 (N_24847,N_11959,N_18340);
nor U24848 (N_24848,N_17471,N_17173);
or U24849 (N_24849,N_16073,N_17639);
or U24850 (N_24850,N_12651,N_11400);
nor U24851 (N_24851,N_10051,N_12939);
nor U24852 (N_24852,N_13914,N_15577);
or U24853 (N_24853,N_12131,N_12945);
nand U24854 (N_24854,N_15656,N_15149);
xnor U24855 (N_24855,N_10857,N_19982);
nor U24856 (N_24856,N_10783,N_16865);
nand U24857 (N_24857,N_13493,N_15301);
or U24858 (N_24858,N_10555,N_19546);
nand U24859 (N_24859,N_17603,N_18338);
nor U24860 (N_24860,N_13927,N_18390);
nand U24861 (N_24861,N_19278,N_10377);
and U24862 (N_24862,N_19940,N_18207);
xor U24863 (N_24863,N_18490,N_14053);
nor U24864 (N_24864,N_17166,N_18687);
and U24865 (N_24865,N_13753,N_19671);
nand U24866 (N_24866,N_15986,N_14873);
and U24867 (N_24867,N_16630,N_14243);
nand U24868 (N_24868,N_18595,N_11808);
or U24869 (N_24869,N_13355,N_18588);
nand U24870 (N_24870,N_18253,N_13542);
or U24871 (N_24871,N_19914,N_12226);
nor U24872 (N_24872,N_17995,N_15279);
nor U24873 (N_24873,N_17150,N_16985);
or U24874 (N_24874,N_18119,N_10974);
nor U24875 (N_24875,N_12460,N_19434);
nand U24876 (N_24876,N_13488,N_10692);
xnor U24877 (N_24877,N_10678,N_11649);
xor U24878 (N_24878,N_18281,N_17617);
or U24879 (N_24879,N_15925,N_15868);
or U24880 (N_24880,N_19854,N_14648);
and U24881 (N_24881,N_12604,N_10431);
nor U24882 (N_24882,N_11152,N_14956);
nand U24883 (N_24883,N_14706,N_14493);
or U24884 (N_24884,N_11939,N_11232);
xnor U24885 (N_24885,N_18084,N_13633);
nor U24886 (N_24886,N_18075,N_10898);
xor U24887 (N_24887,N_17606,N_15663);
nor U24888 (N_24888,N_19362,N_17469);
or U24889 (N_24889,N_19577,N_11989);
or U24890 (N_24890,N_18471,N_16815);
xor U24891 (N_24891,N_17415,N_19933);
nor U24892 (N_24892,N_12709,N_13890);
nand U24893 (N_24893,N_17384,N_14016);
or U24894 (N_24894,N_10321,N_10094);
or U24895 (N_24895,N_13574,N_11331);
and U24896 (N_24896,N_17406,N_12990);
nand U24897 (N_24897,N_11310,N_13703);
nand U24898 (N_24898,N_15826,N_17850);
nor U24899 (N_24899,N_14388,N_11260);
or U24900 (N_24900,N_17914,N_16084);
and U24901 (N_24901,N_15189,N_13023);
xnor U24902 (N_24902,N_14584,N_19008);
nand U24903 (N_24903,N_17608,N_18400);
nand U24904 (N_24904,N_13828,N_17723);
xnor U24905 (N_24905,N_11474,N_14856);
nor U24906 (N_24906,N_15561,N_17199);
nand U24907 (N_24907,N_10337,N_18949);
and U24908 (N_24908,N_10792,N_19965);
and U24909 (N_24909,N_10850,N_19383);
nand U24910 (N_24910,N_16259,N_19033);
xor U24911 (N_24911,N_12524,N_18288);
nor U24912 (N_24912,N_14638,N_12955);
nor U24913 (N_24913,N_13224,N_11135);
nand U24914 (N_24914,N_17857,N_18962);
or U24915 (N_24915,N_11316,N_16088);
and U24916 (N_24916,N_17659,N_10972);
xnor U24917 (N_24917,N_10188,N_11181);
or U24918 (N_24918,N_11725,N_10356);
xor U24919 (N_24919,N_18031,N_18800);
nand U24920 (N_24920,N_10821,N_10738);
nor U24921 (N_24921,N_11233,N_11514);
and U24922 (N_24922,N_11229,N_17337);
nand U24923 (N_24923,N_13667,N_13659);
nand U24924 (N_24924,N_18172,N_11253);
xor U24925 (N_24925,N_16726,N_13163);
xor U24926 (N_24926,N_11177,N_17534);
nand U24927 (N_24927,N_18337,N_12711);
and U24928 (N_24928,N_11617,N_13348);
xnor U24929 (N_24929,N_10562,N_10380);
nor U24930 (N_24930,N_14597,N_11051);
and U24931 (N_24931,N_18508,N_19247);
or U24932 (N_24932,N_18444,N_19019);
nor U24933 (N_24933,N_14360,N_18484);
nand U24934 (N_24934,N_18446,N_14373);
nand U24935 (N_24935,N_11692,N_12989);
or U24936 (N_24936,N_10588,N_10078);
and U24937 (N_24937,N_19817,N_19637);
and U24938 (N_24938,N_14308,N_19761);
nand U24939 (N_24939,N_17677,N_10732);
xor U24940 (N_24940,N_11641,N_11061);
or U24941 (N_24941,N_16634,N_12895);
xnor U24942 (N_24942,N_15882,N_16574);
nor U24943 (N_24943,N_18383,N_11404);
and U24944 (N_24944,N_10750,N_11549);
xnor U24945 (N_24945,N_16524,N_15113);
and U24946 (N_24946,N_10554,N_19573);
xor U24947 (N_24947,N_18189,N_11091);
nor U24948 (N_24948,N_11539,N_14688);
xor U24949 (N_24949,N_17555,N_15116);
nor U24950 (N_24950,N_10429,N_18619);
xor U24951 (N_24951,N_19005,N_12423);
nand U24952 (N_24952,N_11321,N_17503);
xnor U24953 (N_24953,N_11024,N_15028);
and U24954 (N_24954,N_13821,N_18100);
or U24955 (N_24955,N_12117,N_17505);
or U24956 (N_24956,N_15534,N_11154);
or U24957 (N_24957,N_16527,N_14085);
nand U24958 (N_24958,N_15497,N_11411);
nor U24959 (N_24959,N_10785,N_19734);
nor U24960 (N_24960,N_16478,N_12658);
xor U24961 (N_24961,N_13270,N_10167);
or U24962 (N_24962,N_11294,N_15178);
xnor U24963 (N_24963,N_15702,N_10681);
nor U24964 (N_24964,N_14297,N_16251);
and U24965 (N_24965,N_11860,N_11068);
nand U24966 (N_24966,N_19707,N_11129);
xor U24967 (N_24967,N_14734,N_16110);
and U24968 (N_24968,N_19897,N_11341);
or U24969 (N_24969,N_13098,N_12174);
nand U24970 (N_24970,N_10856,N_14404);
and U24971 (N_24971,N_13084,N_11562);
xnor U24972 (N_24972,N_10211,N_17925);
nor U24973 (N_24973,N_13562,N_14518);
nor U24974 (N_24974,N_17811,N_10114);
nor U24975 (N_24975,N_19667,N_13924);
or U24976 (N_24976,N_15284,N_10558);
xnor U24977 (N_24977,N_16390,N_15005);
or U24978 (N_24978,N_10061,N_19938);
xor U24979 (N_24979,N_11120,N_19070);
nand U24980 (N_24980,N_14967,N_17648);
nand U24981 (N_24981,N_16868,N_15464);
xnor U24982 (N_24982,N_11877,N_18791);
xor U24983 (N_24983,N_12756,N_10317);
xor U24984 (N_24984,N_18599,N_17968);
and U24985 (N_24985,N_10818,N_16962);
and U24986 (N_24986,N_15527,N_19968);
or U24987 (N_24987,N_17529,N_14538);
and U24988 (N_24988,N_12420,N_18361);
or U24989 (N_24989,N_17777,N_12146);
nor U24990 (N_24990,N_17225,N_15586);
nor U24991 (N_24991,N_12470,N_11095);
and U24992 (N_24992,N_17127,N_13009);
nor U24993 (N_24993,N_13466,N_10003);
nor U24994 (N_24994,N_17417,N_16552);
nor U24995 (N_24995,N_13848,N_11920);
or U24996 (N_24996,N_18356,N_19130);
nand U24997 (N_24997,N_13591,N_19147);
or U24998 (N_24998,N_15838,N_10400);
or U24999 (N_24999,N_11460,N_10189);
xor U25000 (N_25000,N_11772,N_12904);
nand U25001 (N_25001,N_19786,N_17892);
or U25002 (N_25002,N_13617,N_12862);
nand U25003 (N_25003,N_11502,N_17332);
and U25004 (N_25004,N_18744,N_12770);
and U25005 (N_25005,N_19508,N_16804);
nand U25006 (N_25006,N_17037,N_10911);
or U25007 (N_25007,N_12756,N_17826);
and U25008 (N_25008,N_15035,N_16329);
nor U25009 (N_25009,N_13844,N_13690);
or U25010 (N_25010,N_12802,N_17704);
and U25011 (N_25011,N_13767,N_16190);
xor U25012 (N_25012,N_15364,N_16363);
xnor U25013 (N_25013,N_16820,N_15805);
and U25014 (N_25014,N_10582,N_13764);
xor U25015 (N_25015,N_19600,N_12814);
and U25016 (N_25016,N_10999,N_12755);
or U25017 (N_25017,N_18700,N_13280);
and U25018 (N_25018,N_18069,N_19321);
nand U25019 (N_25019,N_10740,N_13588);
nor U25020 (N_25020,N_14539,N_13167);
or U25021 (N_25021,N_16171,N_16241);
xnor U25022 (N_25022,N_13315,N_13498);
or U25023 (N_25023,N_13573,N_13804);
nor U25024 (N_25024,N_12550,N_14157);
nor U25025 (N_25025,N_15928,N_11227);
and U25026 (N_25026,N_12957,N_14405);
nor U25027 (N_25027,N_10232,N_19666);
nand U25028 (N_25028,N_15151,N_12790);
nor U25029 (N_25029,N_12008,N_11985);
nor U25030 (N_25030,N_10241,N_15844);
xnor U25031 (N_25031,N_18736,N_11612);
or U25032 (N_25032,N_10493,N_18817);
nor U25033 (N_25033,N_19735,N_10780);
nor U25034 (N_25034,N_16275,N_14514);
nor U25035 (N_25035,N_17034,N_13096);
xor U25036 (N_25036,N_10060,N_12408);
or U25037 (N_25037,N_19479,N_14795);
xor U25038 (N_25038,N_16318,N_14870);
nor U25039 (N_25039,N_19893,N_14496);
xor U25040 (N_25040,N_19368,N_11866);
nand U25041 (N_25041,N_17788,N_11284);
nand U25042 (N_25042,N_16116,N_18690);
or U25043 (N_25043,N_12233,N_16069);
xnor U25044 (N_25044,N_10972,N_17820);
or U25045 (N_25045,N_17756,N_15884);
nor U25046 (N_25046,N_17329,N_15680);
or U25047 (N_25047,N_11144,N_18270);
and U25048 (N_25048,N_13082,N_10892);
xnor U25049 (N_25049,N_13167,N_18578);
or U25050 (N_25050,N_10511,N_12090);
and U25051 (N_25051,N_19849,N_11403);
or U25052 (N_25052,N_15279,N_15881);
nor U25053 (N_25053,N_10084,N_10492);
and U25054 (N_25054,N_14429,N_16425);
xnor U25055 (N_25055,N_13117,N_13439);
xnor U25056 (N_25056,N_15965,N_13669);
xor U25057 (N_25057,N_18185,N_13500);
or U25058 (N_25058,N_12065,N_12307);
nand U25059 (N_25059,N_11793,N_16792);
nor U25060 (N_25060,N_15605,N_15768);
or U25061 (N_25061,N_12382,N_19698);
or U25062 (N_25062,N_10457,N_19291);
and U25063 (N_25063,N_19136,N_17433);
xnor U25064 (N_25064,N_12789,N_15557);
and U25065 (N_25065,N_18325,N_14734);
and U25066 (N_25066,N_15885,N_18670);
nand U25067 (N_25067,N_14085,N_18857);
or U25068 (N_25068,N_18937,N_14598);
xnor U25069 (N_25069,N_19553,N_13558);
or U25070 (N_25070,N_11697,N_12410);
or U25071 (N_25071,N_12302,N_19688);
nor U25072 (N_25072,N_15074,N_18645);
or U25073 (N_25073,N_16163,N_16950);
and U25074 (N_25074,N_10152,N_14608);
or U25075 (N_25075,N_19024,N_10866);
nor U25076 (N_25076,N_17263,N_14614);
nor U25077 (N_25077,N_15320,N_16736);
nor U25078 (N_25078,N_18647,N_15219);
nor U25079 (N_25079,N_17347,N_13330);
nor U25080 (N_25080,N_14433,N_10931);
xnor U25081 (N_25081,N_16501,N_17759);
xnor U25082 (N_25082,N_19754,N_11815);
and U25083 (N_25083,N_17932,N_10475);
or U25084 (N_25084,N_10135,N_11900);
or U25085 (N_25085,N_12180,N_11487);
nor U25086 (N_25086,N_15230,N_18227);
or U25087 (N_25087,N_13729,N_12010);
and U25088 (N_25088,N_10030,N_11283);
xnor U25089 (N_25089,N_10828,N_13021);
or U25090 (N_25090,N_16119,N_15406);
or U25091 (N_25091,N_11728,N_19550);
nand U25092 (N_25092,N_10819,N_16039);
nand U25093 (N_25093,N_17531,N_17878);
nand U25094 (N_25094,N_12765,N_12070);
nor U25095 (N_25095,N_18508,N_18784);
xor U25096 (N_25096,N_13309,N_19461);
nor U25097 (N_25097,N_15972,N_11454);
nand U25098 (N_25098,N_13404,N_19256);
xor U25099 (N_25099,N_12028,N_16835);
or U25100 (N_25100,N_13795,N_11514);
or U25101 (N_25101,N_14169,N_19492);
and U25102 (N_25102,N_17201,N_16131);
xnor U25103 (N_25103,N_17758,N_17250);
xnor U25104 (N_25104,N_15206,N_10103);
nand U25105 (N_25105,N_12303,N_11839);
or U25106 (N_25106,N_10596,N_10095);
nor U25107 (N_25107,N_14845,N_16568);
and U25108 (N_25108,N_16078,N_10472);
nor U25109 (N_25109,N_12758,N_11999);
nand U25110 (N_25110,N_11650,N_11030);
and U25111 (N_25111,N_10940,N_15263);
or U25112 (N_25112,N_18077,N_12724);
nor U25113 (N_25113,N_19882,N_13644);
nand U25114 (N_25114,N_15882,N_12246);
xnor U25115 (N_25115,N_18482,N_12587);
or U25116 (N_25116,N_18848,N_12723);
xor U25117 (N_25117,N_17398,N_18019);
and U25118 (N_25118,N_18933,N_15241);
nor U25119 (N_25119,N_13156,N_11184);
nor U25120 (N_25120,N_14398,N_18561);
and U25121 (N_25121,N_15191,N_17657);
nor U25122 (N_25122,N_13317,N_10657);
or U25123 (N_25123,N_13916,N_18913);
and U25124 (N_25124,N_19140,N_10110);
or U25125 (N_25125,N_17891,N_15368);
nand U25126 (N_25126,N_10701,N_14533);
and U25127 (N_25127,N_16089,N_15532);
nand U25128 (N_25128,N_17828,N_15961);
or U25129 (N_25129,N_18619,N_13597);
nand U25130 (N_25130,N_11640,N_18711);
or U25131 (N_25131,N_15953,N_13637);
nand U25132 (N_25132,N_17121,N_15128);
xor U25133 (N_25133,N_14719,N_17950);
or U25134 (N_25134,N_10997,N_17474);
xnor U25135 (N_25135,N_11563,N_13985);
or U25136 (N_25136,N_12839,N_10861);
and U25137 (N_25137,N_15029,N_10542);
nor U25138 (N_25138,N_14595,N_13055);
and U25139 (N_25139,N_10980,N_14538);
nor U25140 (N_25140,N_14589,N_17021);
xor U25141 (N_25141,N_18390,N_16534);
and U25142 (N_25142,N_11846,N_18041);
and U25143 (N_25143,N_17273,N_11724);
nand U25144 (N_25144,N_10824,N_11188);
or U25145 (N_25145,N_10763,N_10581);
or U25146 (N_25146,N_18043,N_19061);
or U25147 (N_25147,N_11212,N_11935);
nand U25148 (N_25148,N_14553,N_12843);
or U25149 (N_25149,N_13932,N_13398);
xnor U25150 (N_25150,N_11999,N_19880);
and U25151 (N_25151,N_14571,N_12463);
nor U25152 (N_25152,N_19344,N_12443);
or U25153 (N_25153,N_12605,N_13165);
and U25154 (N_25154,N_12421,N_14292);
nor U25155 (N_25155,N_11902,N_16991);
nor U25156 (N_25156,N_19359,N_12656);
or U25157 (N_25157,N_11268,N_17662);
nand U25158 (N_25158,N_16426,N_13374);
or U25159 (N_25159,N_12606,N_14925);
and U25160 (N_25160,N_18619,N_18405);
nand U25161 (N_25161,N_19402,N_17253);
or U25162 (N_25162,N_17127,N_18478);
and U25163 (N_25163,N_15157,N_15958);
or U25164 (N_25164,N_13758,N_14454);
nor U25165 (N_25165,N_19010,N_11438);
nand U25166 (N_25166,N_16429,N_15239);
nand U25167 (N_25167,N_18949,N_11273);
xor U25168 (N_25168,N_12701,N_18078);
xor U25169 (N_25169,N_15237,N_12085);
nand U25170 (N_25170,N_12275,N_17013);
or U25171 (N_25171,N_11079,N_10190);
or U25172 (N_25172,N_15556,N_14577);
xor U25173 (N_25173,N_14838,N_15996);
or U25174 (N_25174,N_19554,N_17373);
xor U25175 (N_25175,N_17321,N_16068);
nor U25176 (N_25176,N_19223,N_14898);
and U25177 (N_25177,N_12542,N_13927);
nand U25178 (N_25178,N_12321,N_10187);
and U25179 (N_25179,N_19522,N_15469);
and U25180 (N_25180,N_12227,N_10058);
xnor U25181 (N_25181,N_16558,N_16486);
or U25182 (N_25182,N_14085,N_15800);
and U25183 (N_25183,N_19591,N_10498);
nor U25184 (N_25184,N_12550,N_17618);
nor U25185 (N_25185,N_18652,N_19861);
nor U25186 (N_25186,N_11821,N_15294);
or U25187 (N_25187,N_14117,N_18892);
or U25188 (N_25188,N_18249,N_17027);
or U25189 (N_25189,N_16870,N_12264);
nor U25190 (N_25190,N_11957,N_14581);
xnor U25191 (N_25191,N_15623,N_19558);
or U25192 (N_25192,N_10690,N_15938);
nand U25193 (N_25193,N_14161,N_12121);
nor U25194 (N_25194,N_17006,N_16643);
nor U25195 (N_25195,N_14454,N_17217);
or U25196 (N_25196,N_18856,N_16016);
xnor U25197 (N_25197,N_17922,N_13438);
or U25198 (N_25198,N_12174,N_18042);
and U25199 (N_25199,N_17738,N_10170);
xor U25200 (N_25200,N_12248,N_12146);
nand U25201 (N_25201,N_15629,N_19415);
or U25202 (N_25202,N_18189,N_13983);
nand U25203 (N_25203,N_17571,N_15644);
or U25204 (N_25204,N_10111,N_18510);
xor U25205 (N_25205,N_11785,N_13812);
nor U25206 (N_25206,N_12948,N_18842);
nand U25207 (N_25207,N_14469,N_16466);
nand U25208 (N_25208,N_11173,N_16614);
and U25209 (N_25209,N_12459,N_12736);
or U25210 (N_25210,N_13900,N_11497);
nor U25211 (N_25211,N_12239,N_12304);
or U25212 (N_25212,N_13119,N_15776);
nor U25213 (N_25213,N_12019,N_17781);
xnor U25214 (N_25214,N_16750,N_19456);
xnor U25215 (N_25215,N_14532,N_10776);
and U25216 (N_25216,N_19088,N_15554);
nand U25217 (N_25217,N_12987,N_14107);
nor U25218 (N_25218,N_16307,N_11066);
or U25219 (N_25219,N_12301,N_11364);
nor U25220 (N_25220,N_13030,N_10122);
nor U25221 (N_25221,N_19544,N_17586);
and U25222 (N_25222,N_19720,N_17987);
and U25223 (N_25223,N_12241,N_12481);
or U25224 (N_25224,N_19744,N_15643);
nor U25225 (N_25225,N_16833,N_14735);
and U25226 (N_25226,N_17030,N_11426);
and U25227 (N_25227,N_15472,N_18535);
and U25228 (N_25228,N_14008,N_19082);
nand U25229 (N_25229,N_15869,N_17622);
and U25230 (N_25230,N_10800,N_10177);
or U25231 (N_25231,N_13040,N_11125);
and U25232 (N_25232,N_13140,N_16695);
or U25233 (N_25233,N_18840,N_18313);
nand U25234 (N_25234,N_13084,N_14881);
nand U25235 (N_25235,N_13759,N_19868);
nand U25236 (N_25236,N_14560,N_18803);
nand U25237 (N_25237,N_16373,N_17876);
nand U25238 (N_25238,N_19088,N_12760);
nor U25239 (N_25239,N_14406,N_17759);
nand U25240 (N_25240,N_10452,N_15786);
xnor U25241 (N_25241,N_10496,N_14101);
or U25242 (N_25242,N_10069,N_12008);
xnor U25243 (N_25243,N_13409,N_13770);
or U25244 (N_25244,N_16755,N_18679);
xnor U25245 (N_25245,N_19198,N_17454);
nand U25246 (N_25246,N_19419,N_15206);
and U25247 (N_25247,N_18551,N_19570);
and U25248 (N_25248,N_17870,N_16596);
and U25249 (N_25249,N_14670,N_16449);
and U25250 (N_25250,N_18411,N_12821);
or U25251 (N_25251,N_12688,N_10594);
nor U25252 (N_25252,N_18829,N_18763);
xor U25253 (N_25253,N_11404,N_14972);
nor U25254 (N_25254,N_13462,N_15707);
xor U25255 (N_25255,N_12859,N_14595);
xnor U25256 (N_25256,N_18085,N_14637);
or U25257 (N_25257,N_12060,N_19084);
and U25258 (N_25258,N_12058,N_14189);
and U25259 (N_25259,N_12584,N_14667);
or U25260 (N_25260,N_18496,N_10689);
nor U25261 (N_25261,N_11019,N_15242);
xor U25262 (N_25262,N_15839,N_17184);
xor U25263 (N_25263,N_19298,N_18975);
nor U25264 (N_25264,N_16278,N_15786);
xor U25265 (N_25265,N_15477,N_12468);
xor U25266 (N_25266,N_15296,N_15665);
xor U25267 (N_25267,N_11592,N_18488);
or U25268 (N_25268,N_11211,N_15539);
nand U25269 (N_25269,N_14789,N_10214);
and U25270 (N_25270,N_11599,N_18402);
or U25271 (N_25271,N_13802,N_14039);
xnor U25272 (N_25272,N_12859,N_17214);
xor U25273 (N_25273,N_17573,N_18549);
or U25274 (N_25274,N_10025,N_19515);
nand U25275 (N_25275,N_19741,N_19760);
and U25276 (N_25276,N_19591,N_14543);
nand U25277 (N_25277,N_19072,N_18230);
xnor U25278 (N_25278,N_10210,N_13345);
xor U25279 (N_25279,N_16702,N_18408);
nand U25280 (N_25280,N_19311,N_10345);
xor U25281 (N_25281,N_19083,N_16741);
and U25282 (N_25282,N_12381,N_16448);
xnor U25283 (N_25283,N_14295,N_10190);
xor U25284 (N_25284,N_16505,N_11336);
nor U25285 (N_25285,N_18219,N_19326);
and U25286 (N_25286,N_12896,N_13341);
or U25287 (N_25287,N_17596,N_10270);
nand U25288 (N_25288,N_13654,N_15322);
or U25289 (N_25289,N_17096,N_19402);
xnor U25290 (N_25290,N_16180,N_13882);
nor U25291 (N_25291,N_15708,N_13146);
nand U25292 (N_25292,N_16676,N_16758);
xnor U25293 (N_25293,N_16004,N_18468);
or U25294 (N_25294,N_19457,N_17856);
and U25295 (N_25295,N_12712,N_19087);
nand U25296 (N_25296,N_16435,N_18127);
and U25297 (N_25297,N_13791,N_13795);
and U25298 (N_25298,N_19293,N_10026);
xor U25299 (N_25299,N_19523,N_17056);
and U25300 (N_25300,N_13394,N_15858);
nor U25301 (N_25301,N_18210,N_18338);
nand U25302 (N_25302,N_13135,N_16352);
or U25303 (N_25303,N_19521,N_10663);
or U25304 (N_25304,N_17383,N_10802);
xor U25305 (N_25305,N_15424,N_13931);
nand U25306 (N_25306,N_16475,N_18322);
nand U25307 (N_25307,N_10733,N_12293);
and U25308 (N_25308,N_11115,N_17065);
or U25309 (N_25309,N_12873,N_15947);
or U25310 (N_25310,N_13772,N_19551);
and U25311 (N_25311,N_11571,N_18580);
nand U25312 (N_25312,N_19587,N_10668);
and U25313 (N_25313,N_16801,N_15091);
nor U25314 (N_25314,N_16633,N_18999);
and U25315 (N_25315,N_14477,N_16049);
xnor U25316 (N_25316,N_13207,N_15845);
or U25317 (N_25317,N_15853,N_13132);
xor U25318 (N_25318,N_14829,N_13503);
nor U25319 (N_25319,N_18861,N_15298);
nand U25320 (N_25320,N_15756,N_18653);
and U25321 (N_25321,N_13694,N_10509);
xor U25322 (N_25322,N_13607,N_14677);
nand U25323 (N_25323,N_11442,N_14257);
or U25324 (N_25324,N_15463,N_12698);
nand U25325 (N_25325,N_18384,N_18450);
xnor U25326 (N_25326,N_14573,N_14980);
or U25327 (N_25327,N_15577,N_15718);
nand U25328 (N_25328,N_18178,N_16809);
nor U25329 (N_25329,N_15496,N_11253);
or U25330 (N_25330,N_13411,N_17284);
nand U25331 (N_25331,N_16651,N_11820);
or U25332 (N_25332,N_15430,N_10052);
xnor U25333 (N_25333,N_11021,N_12565);
nor U25334 (N_25334,N_12253,N_17509);
or U25335 (N_25335,N_14319,N_11029);
nor U25336 (N_25336,N_18846,N_12325);
nand U25337 (N_25337,N_10966,N_18199);
or U25338 (N_25338,N_14159,N_16948);
nor U25339 (N_25339,N_12024,N_15105);
xor U25340 (N_25340,N_17927,N_17679);
xor U25341 (N_25341,N_12931,N_14149);
xor U25342 (N_25342,N_11884,N_15715);
nand U25343 (N_25343,N_11739,N_19722);
xnor U25344 (N_25344,N_15096,N_12223);
or U25345 (N_25345,N_13536,N_13609);
or U25346 (N_25346,N_19439,N_18625);
and U25347 (N_25347,N_14451,N_11401);
nor U25348 (N_25348,N_13948,N_15749);
xor U25349 (N_25349,N_13328,N_18558);
nor U25350 (N_25350,N_13966,N_14922);
xnor U25351 (N_25351,N_10162,N_19916);
nand U25352 (N_25352,N_11051,N_13250);
nor U25353 (N_25353,N_13526,N_11034);
nand U25354 (N_25354,N_10999,N_13939);
xnor U25355 (N_25355,N_17024,N_12293);
nor U25356 (N_25356,N_17784,N_11663);
and U25357 (N_25357,N_16450,N_12505);
xor U25358 (N_25358,N_17615,N_15874);
or U25359 (N_25359,N_17894,N_19406);
xnor U25360 (N_25360,N_10914,N_18134);
nor U25361 (N_25361,N_12965,N_17765);
nand U25362 (N_25362,N_10628,N_13330);
xnor U25363 (N_25363,N_13906,N_11211);
xor U25364 (N_25364,N_14670,N_11139);
nor U25365 (N_25365,N_18022,N_18347);
or U25366 (N_25366,N_16118,N_10503);
xnor U25367 (N_25367,N_16263,N_16065);
or U25368 (N_25368,N_17177,N_18665);
or U25369 (N_25369,N_10768,N_13526);
xor U25370 (N_25370,N_13971,N_17119);
xor U25371 (N_25371,N_19456,N_14474);
and U25372 (N_25372,N_11403,N_15935);
nor U25373 (N_25373,N_11500,N_10745);
nand U25374 (N_25374,N_13437,N_13043);
nor U25375 (N_25375,N_18361,N_15526);
or U25376 (N_25376,N_16931,N_11542);
or U25377 (N_25377,N_17998,N_16794);
nand U25378 (N_25378,N_12720,N_11279);
or U25379 (N_25379,N_12418,N_11299);
nand U25380 (N_25380,N_12015,N_17996);
xnor U25381 (N_25381,N_13911,N_18820);
xnor U25382 (N_25382,N_11498,N_19042);
and U25383 (N_25383,N_19537,N_17268);
or U25384 (N_25384,N_11424,N_10488);
or U25385 (N_25385,N_17165,N_18094);
or U25386 (N_25386,N_14503,N_19149);
or U25387 (N_25387,N_11091,N_18022);
nor U25388 (N_25388,N_10908,N_19290);
xor U25389 (N_25389,N_11707,N_11276);
or U25390 (N_25390,N_11304,N_16514);
nor U25391 (N_25391,N_14357,N_14411);
or U25392 (N_25392,N_16819,N_15363);
and U25393 (N_25393,N_11096,N_18761);
or U25394 (N_25394,N_16852,N_14064);
or U25395 (N_25395,N_18012,N_16364);
and U25396 (N_25396,N_13999,N_18629);
and U25397 (N_25397,N_19783,N_12696);
xor U25398 (N_25398,N_12103,N_12008);
nor U25399 (N_25399,N_17874,N_14544);
and U25400 (N_25400,N_19918,N_13536);
or U25401 (N_25401,N_17978,N_12287);
nand U25402 (N_25402,N_18673,N_18406);
nor U25403 (N_25403,N_19052,N_18577);
or U25404 (N_25404,N_16082,N_17057);
or U25405 (N_25405,N_15344,N_11287);
nor U25406 (N_25406,N_16077,N_10419);
or U25407 (N_25407,N_17362,N_13890);
nand U25408 (N_25408,N_17312,N_13579);
and U25409 (N_25409,N_11446,N_13314);
nand U25410 (N_25410,N_18736,N_15810);
nor U25411 (N_25411,N_15037,N_12998);
or U25412 (N_25412,N_19318,N_12082);
and U25413 (N_25413,N_12862,N_16774);
and U25414 (N_25414,N_19098,N_16380);
nor U25415 (N_25415,N_12839,N_11054);
or U25416 (N_25416,N_15503,N_12724);
nand U25417 (N_25417,N_16766,N_16488);
nor U25418 (N_25418,N_10429,N_10271);
xor U25419 (N_25419,N_17035,N_16175);
nand U25420 (N_25420,N_18878,N_12864);
nor U25421 (N_25421,N_12452,N_11411);
nand U25422 (N_25422,N_12706,N_13022);
nor U25423 (N_25423,N_19427,N_13758);
or U25424 (N_25424,N_16604,N_19233);
or U25425 (N_25425,N_11879,N_18295);
nor U25426 (N_25426,N_11793,N_15210);
nor U25427 (N_25427,N_16134,N_14925);
xor U25428 (N_25428,N_15757,N_10990);
and U25429 (N_25429,N_11693,N_16229);
or U25430 (N_25430,N_15045,N_11047);
and U25431 (N_25431,N_13529,N_18058);
nor U25432 (N_25432,N_11635,N_17035);
or U25433 (N_25433,N_16014,N_16226);
or U25434 (N_25434,N_11686,N_16947);
xor U25435 (N_25435,N_13296,N_19627);
and U25436 (N_25436,N_10774,N_16238);
or U25437 (N_25437,N_17818,N_17855);
nand U25438 (N_25438,N_18136,N_12903);
nand U25439 (N_25439,N_15594,N_10567);
xnor U25440 (N_25440,N_11875,N_15479);
or U25441 (N_25441,N_14793,N_18164);
nand U25442 (N_25442,N_19130,N_18109);
nor U25443 (N_25443,N_18783,N_13420);
or U25444 (N_25444,N_17450,N_18010);
xnor U25445 (N_25445,N_11132,N_15380);
and U25446 (N_25446,N_10778,N_10743);
or U25447 (N_25447,N_14210,N_11554);
xnor U25448 (N_25448,N_15828,N_18913);
or U25449 (N_25449,N_17746,N_18233);
and U25450 (N_25450,N_13517,N_12596);
and U25451 (N_25451,N_16981,N_11847);
nand U25452 (N_25452,N_14403,N_12188);
nor U25453 (N_25453,N_11894,N_10449);
nor U25454 (N_25454,N_13333,N_19699);
xor U25455 (N_25455,N_12290,N_17785);
and U25456 (N_25456,N_10404,N_17649);
and U25457 (N_25457,N_19927,N_18919);
or U25458 (N_25458,N_11379,N_11109);
and U25459 (N_25459,N_18456,N_11535);
or U25460 (N_25460,N_18963,N_15097);
nand U25461 (N_25461,N_19362,N_16255);
nor U25462 (N_25462,N_17308,N_14679);
nor U25463 (N_25463,N_14282,N_10062);
and U25464 (N_25464,N_10520,N_15879);
nor U25465 (N_25465,N_14621,N_18238);
or U25466 (N_25466,N_17536,N_12889);
nand U25467 (N_25467,N_11488,N_10062);
or U25468 (N_25468,N_14505,N_11505);
nor U25469 (N_25469,N_18549,N_12251);
nand U25470 (N_25470,N_14592,N_19493);
and U25471 (N_25471,N_13988,N_15204);
or U25472 (N_25472,N_12641,N_17897);
nand U25473 (N_25473,N_18462,N_16517);
nor U25474 (N_25474,N_11730,N_18110);
nor U25475 (N_25475,N_12440,N_12028);
nor U25476 (N_25476,N_10977,N_14602);
nor U25477 (N_25477,N_13952,N_12176);
nand U25478 (N_25478,N_14676,N_13871);
nor U25479 (N_25479,N_19852,N_19438);
nor U25480 (N_25480,N_13825,N_16464);
and U25481 (N_25481,N_15422,N_18223);
nand U25482 (N_25482,N_15688,N_12236);
nand U25483 (N_25483,N_14681,N_17250);
xnor U25484 (N_25484,N_13101,N_13689);
or U25485 (N_25485,N_10613,N_16689);
or U25486 (N_25486,N_18896,N_16188);
or U25487 (N_25487,N_19810,N_17919);
nand U25488 (N_25488,N_14369,N_18389);
nor U25489 (N_25489,N_12994,N_15931);
or U25490 (N_25490,N_13797,N_18287);
and U25491 (N_25491,N_17762,N_12872);
xor U25492 (N_25492,N_16157,N_12085);
xor U25493 (N_25493,N_12142,N_19700);
xnor U25494 (N_25494,N_19381,N_11509);
nand U25495 (N_25495,N_13622,N_19637);
or U25496 (N_25496,N_11430,N_18567);
or U25497 (N_25497,N_17016,N_19295);
nor U25498 (N_25498,N_15361,N_11795);
nand U25499 (N_25499,N_19370,N_10335);
nor U25500 (N_25500,N_10765,N_11926);
nand U25501 (N_25501,N_11159,N_12832);
nor U25502 (N_25502,N_14584,N_18084);
and U25503 (N_25503,N_17241,N_13557);
nor U25504 (N_25504,N_15574,N_18135);
nor U25505 (N_25505,N_16538,N_15936);
nor U25506 (N_25506,N_13161,N_19849);
xor U25507 (N_25507,N_18029,N_18094);
nand U25508 (N_25508,N_10849,N_17766);
nand U25509 (N_25509,N_14310,N_14559);
xnor U25510 (N_25510,N_18372,N_14696);
or U25511 (N_25511,N_11243,N_15660);
and U25512 (N_25512,N_10154,N_15624);
or U25513 (N_25513,N_10603,N_14235);
nand U25514 (N_25514,N_15851,N_18749);
xor U25515 (N_25515,N_15053,N_10504);
and U25516 (N_25516,N_10381,N_16926);
nand U25517 (N_25517,N_15766,N_16495);
or U25518 (N_25518,N_10164,N_14636);
nor U25519 (N_25519,N_11406,N_16313);
nand U25520 (N_25520,N_17167,N_19538);
nor U25521 (N_25521,N_12087,N_19007);
or U25522 (N_25522,N_12808,N_15489);
nand U25523 (N_25523,N_16514,N_13078);
xor U25524 (N_25524,N_17040,N_17031);
nand U25525 (N_25525,N_16141,N_18365);
nor U25526 (N_25526,N_13259,N_12769);
xor U25527 (N_25527,N_13915,N_14375);
and U25528 (N_25528,N_10859,N_15576);
nor U25529 (N_25529,N_13580,N_18474);
nand U25530 (N_25530,N_18781,N_16546);
xor U25531 (N_25531,N_15070,N_17110);
xor U25532 (N_25532,N_15329,N_13254);
nor U25533 (N_25533,N_19699,N_16232);
and U25534 (N_25534,N_19542,N_16835);
and U25535 (N_25535,N_14898,N_11847);
xnor U25536 (N_25536,N_17866,N_19384);
or U25537 (N_25537,N_18543,N_10385);
xnor U25538 (N_25538,N_16014,N_17818);
nor U25539 (N_25539,N_12097,N_17318);
nand U25540 (N_25540,N_16642,N_10450);
or U25541 (N_25541,N_16166,N_18364);
and U25542 (N_25542,N_12328,N_12351);
nor U25543 (N_25543,N_12470,N_11171);
nor U25544 (N_25544,N_18645,N_17547);
or U25545 (N_25545,N_19166,N_10273);
and U25546 (N_25546,N_12082,N_10498);
nor U25547 (N_25547,N_18150,N_10172);
or U25548 (N_25548,N_17594,N_16921);
xor U25549 (N_25549,N_11003,N_16255);
xor U25550 (N_25550,N_12724,N_12710);
xor U25551 (N_25551,N_18849,N_10812);
nor U25552 (N_25552,N_10055,N_15334);
or U25553 (N_25553,N_17041,N_14816);
or U25554 (N_25554,N_11471,N_13748);
nor U25555 (N_25555,N_12837,N_14486);
nand U25556 (N_25556,N_14089,N_15229);
or U25557 (N_25557,N_10824,N_12141);
xnor U25558 (N_25558,N_10100,N_15521);
nand U25559 (N_25559,N_11605,N_11053);
or U25560 (N_25560,N_19919,N_16239);
xnor U25561 (N_25561,N_14056,N_11666);
nand U25562 (N_25562,N_16023,N_18882);
nor U25563 (N_25563,N_15500,N_19978);
and U25564 (N_25564,N_14695,N_13380);
and U25565 (N_25565,N_10240,N_10154);
nand U25566 (N_25566,N_15048,N_14149);
or U25567 (N_25567,N_10481,N_16676);
nand U25568 (N_25568,N_11870,N_10418);
or U25569 (N_25569,N_10360,N_15146);
and U25570 (N_25570,N_10665,N_11095);
or U25571 (N_25571,N_11491,N_10166);
nand U25572 (N_25572,N_10673,N_11973);
and U25573 (N_25573,N_17548,N_11772);
or U25574 (N_25574,N_14758,N_14175);
xnor U25575 (N_25575,N_15071,N_10439);
or U25576 (N_25576,N_13543,N_14651);
and U25577 (N_25577,N_14363,N_12312);
xor U25578 (N_25578,N_14503,N_10705);
or U25579 (N_25579,N_12903,N_11210);
nor U25580 (N_25580,N_13757,N_19208);
or U25581 (N_25581,N_15578,N_11255);
and U25582 (N_25582,N_11462,N_16730);
nand U25583 (N_25583,N_17351,N_18557);
and U25584 (N_25584,N_12166,N_14073);
nand U25585 (N_25585,N_13687,N_14857);
nand U25586 (N_25586,N_15815,N_12759);
or U25587 (N_25587,N_11243,N_17845);
nand U25588 (N_25588,N_11441,N_15209);
nor U25589 (N_25589,N_19521,N_19689);
and U25590 (N_25590,N_18677,N_14903);
xnor U25591 (N_25591,N_14815,N_11596);
or U25592 (N_25592,N_10427,N_12610);
nand U25593 (N_25593,N_14337,N_10733);
or U25594 (N_25594,N_13694,N_18535);
nor U25595 (N_25595,N_17573,N_17307);
xnor U25596 (N_25596,N_18315,N_12043);
nor U25597 (N_25597,N_14273,N_13240);
nand U25598 (N_25598,N_13398,N_12652);
or U25599 (N_25599,N_17194,N_13986);
nor U25600 (N_25600,N_19367,N_10893);
xnor U25601 (N_25601,N_10633,N_19325);
nor U25602 (N_25602,N_17940,N_12503);
or U25603 (N_25603,N_15523,N_17154);
nand U25604 (N_25604,N_17358,N_17513);
nor U25605 (N_25605,N_18967,N_12903);
nor U25606 (N_25606,N_13450,N_10209);
xor U25607 (N_25607,N_14525,N_14594);
or U25608 (N_25608,N_18137,N_11884);
or U25609 (N_25609,N_11423,N_11619);
nor U25610 (N_25610,N_19124,N_11194);
nor U25611 (N_25611,N_15261,N_15868);
nor U25612 (N_25612,N_10609,N_12393);
and U25613 (N_25613,N_18117,N_15937);
nand U25614 (N_25614,N_18524,N_19932);
or U25615 (N_25615,N_17973,N_19066);
and U25616 (N_25616,N_10585,N_14584);
or U25617 (N_25617,N_12176,N_15387);
nand U25618 (N_25618,N_11648,N_18302);
or U25619 (N_25619,N_16234,N_12240);
xor U25620 (N_25620,N_19076,N_15512);
nand U25621 (N_25621,N_19034,N_15334);
nand U25622 (N_25622,N_12688,N_19848);
nand U25623 (N_25623,N_11632,N_13564);
or U25624 (N_25624,N_16358,N_16061);
nand U25625 (N_25625,N_11403,N_19213);
xor U25626 (N_25626,N_18245,N_13197);
xnor U25627 (N_25627,N_10504,N_11515);
xnor U25628 (N_25628,N_15980,N_10962);
nor U25629 (N_25629,N_12863,N_18879);
and U25630 (N_25630,N_13851,N_12815);
xnor U25631 (N_25631,N_13123,N_10352);
and U25632 (N_25632,N_14519,N_14363);
xor U25633 (N_25633,N_12037,N_15390);
nor U25634 (N_25634,N_12365,N_18803);
or U25635 (N_25635,N_16682,N_14552);
and U25636 (N_25636,N_16907,N_18059);
nand U25637 (N_25637,N_11371,N_19788);
or U25638 (N_25638,N_12257,N_16914);
or U25639 (N_25639,N_11805,N_17081);
nor U25640 (N_25640,N_10337,N_17128);
and U25641 (N_25641,N_18885,N_19702);
xor U25642 (N_25642,N_10878,N_11191);
or U25643 (N_25643,N_13463,N_18727);
or U25644 (N_25644,N_13477,N_17289);
or U25645 (N_25645,N_19787,N_11727);
and U25646 (N_25646,N_10636,N_17551);
nand U25647 (N_25647,N_19835,N_16015);
or U25648 (N_25648,N_13939,N_19707);
nand U25649 (N_25649,N_12925,N_17555);
and U25650 (N_25650,N_10426,N_16700);
nand U25651 (N_25651,N_19249,N_17200);
xor U25652 (N_25652,N_19727,N_10727);
nand U25653 (N_25653,N_16157,N_13461);
xor U25654 (N_25654,N_18522,N_17433);
and U25655 (N_25655,N_12172,N_11160);
xnor U25656 (N_25656,N_10581,N_12831);
nor U25657 (N_25657,N_18259,N_17585);
nor U25658 (N_25658,N_15341,N_14724);
and U25659 (N_25659,N_16772,N_11656);
xor U25660 (N_25660,N_16804,N_19197);
and U25661 (N_25661,N_12769,N_18837);
nor U25662 (N_25662,N_12429,N_12476);
nor U25663 (N_25663,N_12481,N_14528);
or U25664 (N_25664,N_12564,N_17648);
and U25665 (N_25665,N_12859,N_12168);
and U25666 (N_25666,N_10514,N_14412);
or U25667 (N_25667,N_16316,N_16014);
nand U25668 (N_25668,N_18876,N_18830);
xor U25669 (N_25669,N_16487,N_18704);
nor U25670 (N_25670,N_12578,N_17837);
and U25671 (N_25671,N_17628,N_16999);
xor U25672 (N_25672,N_10749,N_15776);
nor U25673 (N_25673,N_13268,N_16253);
or U25674 (N_25674,N_11145,N_19551);
or U25675 (N_25675,N_18531,N_11434);
xor U25676 (N_25676,N_17869,N_16533);
xor U25677 (N_25677,N_12773,N_14587);
nand U25678 (N_25678,N_10626,N_10178);
and U25679 (N_25679,N_16744,N_19100);
or U25680 (N_25680,N_10934,N_17643);
and U25681 (N_25681,N_12424,N_16091);
nand U25682 (N_25682,N_11159,N_16774);
or U25683 (N_25683,N_12944,N_13093);
nand U25684 (N_25684,N_17034,N_16227);
and U25685 (N_25685,N_12259,N_19252);
or U25686 (N_25686,N_17370,N_18309);
nor U25687 (N_25687,N_15475,N_18849);
or U25688 (N_25688,N_14914,N_19961);
or U25689 (N_25689,N_14710,N_16682);
nand U25690 (N_25690,N_10865,N_10717);
and U25691 (N_25691,N_15262,N_15962);
or U25692 (N_25692,N_15198,N_13260);
and U25693 (N_25693,N_10520,N_13391);
or U25694 (N_25694,N_15795,N_15768);
nor U25695 (N_25695,N_11322,N_17186);
xnor U25696 (N_25696,N_11572,N_15597);
xnor U25697 (N_25697,N_14042,N_11874);
xnor U25698 (N_25698,N_11319,N_12187);
or U25699 (N_25699,N_11393,N_11417);
and U25700 (N_25700,N_13457,N_15126);
nand U25701 (N_25701,N_11357,N_16045);
and U25702 (N_25702,N_13174,N_18235);
or U25703 (N_25703,N_14812,N_16669);
nand U25704 (N_25704,N_16627,N_11418);
xor U25705 (N_25705,N_19623,N_11711);
or U25706 (N_25706,N_14256,N_12407);
or U25707 (N_25707,N_14249,N_15905);
or U25708 (N_25708,N_14486,N_11450);
and U25709 (N_25709,N_16737,N_14266);
xor U25710 (N_25710,N_12780,N_19303);
xnor U25711 (N_25711,N_12981,N_15696);
and U25712 (N_25712,N_13203,N_17902);
nand U25713 (N_25713,N_19854,N_14553);
nand U25714 (N_25714,N_19828,N_15656);
and U25715 (N_25715,N_11525,N_17167);
and U25716 (N_25716,N_10928,N_16167);
xnor U25717 (N_25717,N_17519,N_12688);
nand U25718 (N_25718,N_18692,N_14344);
xor U25719 (N_25719,N_18053,N_18914);
or U25720 (N_25720,N_15357,N_16421);
and U25721 (N_25721,N_13462,N_13714);
nor U25722 (N_25722,N_19229,N_18686);
nor U25723 (N_25723,N_10796,N_15657);
or U25724 (N_25724,N_18158,N_10100);
nand U25725 (N_25725,N_19261,N_12814);
xor U25726 (N_25726,N_14277,N_16382);
and U25727 (N_25727,N_15358,N_16987);
nor U25728 (N_25728,N_16540,N_14260);
xnor U25729 (N_25729,N_12753,N_14316);
nand U25730 (N_25730,N_16307,N_15738);
nor U25731 (N_25731,N_14064,N_17374);
nor U25732 (N_25732,N_15437,N_16569);
nor U25733 (N_25733,N_13944,N_14730);
or U25734 (N_25734,N_13232,N_17138);
nand U25735 (N_25735,N_18566,N_16849);
nand U25736 (N_25736,N_17505,N_14678);
and U25737 (N_25737,N_19645,N_15427);
nor U25738 (N_25738,N_16182,N_10655);
and U25739 (N_25739,N_17625,N_11689);
xnor U25740 (N_25740,N_13969,N_12342);
and U25741 (N_25741,N_19280,N_15768);
xor U25742 (N_25742,N_12098,N_16389);
or U25743 (N_25743,N_19153,N_19819);
or U25744 (N_25744,N_10938,N_13981);
and U25745 (N_25745,N_12253,N_13306);
nand U25746 (N_25746,N_15317,N_10015);
or U25747 (N_25747,N_13375,N_14964);
or U25748 (N_25748,N_10119,N_15380);
nand U25749 (N_25749,N_17731,N_14943);
xnor U25750 (N_25750,N_18986,N_10766);
nand U25751 (N_25751,N_14323,N_19198);
xor U25752 (N_25752,N_16731,N_17228);
xor U25753 (N_25753,N_12372,N_18597);
xnor U25754 (N_25754,N_12394,N_17406);
xnor U25755 (N_25755,N_17122,N_17629);
nand U25756 (N_25756,N_15358,N_15552);
and U25757 (N_25757,N_17419,N_15446);
xnor U25758 (N_25758,N_13321,N_11578);
and U25759 (N_25759,N_13783,N_13475);
or U25760 (N_25760,N_14285,N_19594);
and U25761 (N_25761,N_11695,N_10620);
nor U25762 (N_25762,N_12345,N_13539);
nand U25763 (N_25763,N_10449,N_19911);
xnor U25764 (N_25764,N_19547,N_10898);
and U25765 (N_25765,N_15235,N_11632);
nor U25766 (N_25766,N_19887,N_14596);
nor U25767 (N_25767,N_19159,N_15430);
nor U25768 (N_25768,N_18788,N_16934);
nand U25769 (N_25769,N_18487,N_14237);
or U25770 (N_25770,N_14663,N_19729);
nand U25771 (N_25771,N_18055,N_19000);
and U25772 (N_25772,N_12013,N_17406);
xnor U25773 (N_25773,N_14197,N_17789);
nand U25774 (N_25774,N_12965,N_15938);
xnor U25775 (N_25775,N_16562,N_19489);
or U25776 (N_25776,N_19904,N_19030);
nand U25777 (N_25777,N_10890,N_11451);
xor U25778 (N_25778,N_12070,N_16512);
or U25779 (N_25779,N_14670,N_18755);
nor U25780 (N_25780,N_11732,N_18735);
nand U25781 (N_25781,N_11346,N_19980);
nand U25782 (N_25782,N_11743,N_14509);
xor U25783 (N_25783,N_16949,N_13166);
and U25784 (N_25784,N_10017,N_17944);
nor U25785 (N_25785,N_18319,N_13678);
nand U25786 (N_25786,N_14459,N_19412);
and U25787 (N_25787,N_13884,N_11386);
nand U25788 (N_25788,N_17602,N_19009);
xor U25789 (N_25789,N_12878,N_17868);
xnor U25790 (N_25790,N_19321,N_12791);
or U25791 (N_25791,N_16710,N_13142);
xor U25792 (N_25792,N_19454,N_18963);
nand U25793 (N_25793,N_11784,N_15185);
nand U25794 (N_25794,N_12940,N_15181);
and U25795 (N_25795,N_14027,N_19953);
nor U25796 (N_25796,N_17256,N_18126);
or U25797 (N_25797,N_14345,N_13238);
and U25798 (N_25798,N_10634,N_16365);
nand U25799 (N_25799,N_18745,N_10711);
or U25800 (N_25800,N_13117,N_15287);
xor U25801 (N_25801,N_12556,N_18132);
nand U25802 (N_25802,N_15287,N_15270);
nand U25803 (N_25803,N_13252,N_19211);
and U25804 (N_25804,N_19129,N_14837);
nand U25805 (N_25805,N_14804,N_14271);
or U25806 (N_25806,N_10486,N_10813);
nand U25807 (N_25807,N_17870,N_10177);
or U25808 (N_25808,N_18189,N_17346);
nand U25809 (N_25809,N_12170,N_19990);
or U25810 (N_25810,N_18056,N_11114);
nand U25811 (N_25811,N_15492,N_14439);
nand U25812 (N_25812,N_11218,N_10880);
and U25813 (N_25813,N_11543,N_17923);
or U25814 (N_25814,N_17936,N_11869);
xor U25815 (N_25815,N_18972,N_16452);
nand U25816 (N_25816,N_12055,N_16311);
nor U25817 (N_25817,N_19802,N_12152);
xnor U25818 (N_25818,N_19734,N_16832);
and U25819 (N_25819,N_16430,N_10734);
nand U25820 (N_25820,N_14766,N_11377);
nor U25821 (N_25821,N_16654,N_13178);
or U25822 (N_25822,N_19872,N_10448);
or U25823 (N_25823,N_15220,N_12178);
nor U25824 (N_25824,N_17247,N_13016);
nor U25825 (N_25825,N_11924,N_16688);
nand U25826 (N_25826,N_18285,N_16552);
or U25827 (N_25827,N_19592,N_18906);
nor U25828 (N_25828,N_18366,N_13267);
or U25829 (N_25829,N_13620,N_14907);
or U25830 (N_25830,N_10424,N_16770);
nor U25831 (N_25831,N_11609,N_18627);
nor U25832 (N_25832,N_10444,N_13429);
xor U25833 (N_25833,N_12726,N_16545);
nor U25834 (N_25834,N_14591,N_12499);
nand U25835 (N_25835,N_17239,N_12794);
and U25836 (N_25836,N_15557,N_17953);
and U25837 (N_25837,N_19210,N_15824);
xor U25838 (N_25838,N_10362,N_18449);
xnor U25839 (N_25839,N_13960,N_16809);
or U25840 (N_25840,N_11106,N_11012);
nand U25841 (N_25841,N_15950,N_13814);
nand U25842 (N_25842,N_10882,N_18477);
and U25843 (N_25843,N_15145,N_17752);
or U25844 (N_25844,N_18237,N_10085);
nand U25845 (N_25845,N_16706,N_11040);
xnor U25846 (N_25846,N_19936,N_10956);
nand U25847 (N_25847,N_14244,N_17616);
nor U25848 (N_25848,N_17124,N_13860);
nand U25849 (N_25849,N_12067,N_11940);
or U25850 (N_25850,N_11344,N_11071);
and U25851 (N_25851,N_11791,N_14841);
nand U25852 (N_25852,N_11909,N_10346);
and U25853 (N_25853,N_18407,N_12200);
or U25854 (N_25854,N_16652,N_13453);
nor U25855 (N_25855,N_14955,N_11395);
nand U25856 (N_25856,N_10179,N_18717);
and U25857 (N_25857,N_16315,N_10235);
nor U25858 (N_25858,N_12554,N_11749);
xor U25859 (N_25859,N_19059,N_14976);
or U25860 (N_25860,N_10003,N_11934);
and U25861 (N_25861,N_14186,N_11855);
or U25862 (N_25862,N_19798,N_17197);
xnor U25863 (N_25863,N_17645,N_19033);
xor U25864 (N_25864,N_18782,N_16970);
or U25865 (N_25865,N_11335,N_19098);
nor U25866 (N_25866,N_18934,N_16824);
or U25867 (N_25867,N_13857,N_12726);
nor U25868 (N_25868,N_13775,N_13043);
or U25869 (N_25869,N_12887,N_10752);
nor U25870 (N_25870,N_17004,N_18141);
and U25871 (N_25871,N_11253,N_11502);
and U25872 (N_25872,N_12311,N_14192);
or U25873 (N_25873,N_16787,N_18335);
nand U25874 (N_25874,N_12716,N_14437);
nand U25875 (N_25875,N_17545,N_12473);
xor U25876 (N_25876,N_17459,N_10146);
or U25877 (N_25877,N_19005,N_14198);
xor U25878 (N_25878,N_10357,N_13567);
and U25879 (N_25879,N_16906,N_14397);
or U25880 (N_25880,N_14877,N_16072);
xnor U25881 (N_25881,N_17238,N_15238);
or U25882 (N_25882,N_19049,N_13179);
nor U25883 (N_25883,N_19197,N_16382);
nor U25884 (N_25884,N_17994,N_14939);
nand U25885 (N_25885,N_14718,N_15344);
nand U25886 (N_25886,N_15764,N_19494);
xnor U25887 (N_25887,N_14759,N_17232);
nand U25888 (N_25888,N_17721,N_19251);
nor U25889 (N_25889,N_14083,N_16655);
or U25890 (N_25890,N_19091,N_16881);
nand U25891 (N_25891,N_19678,N_10037);
and U25892 (N_25892,N_17535,N_11052);
xnor U25893 (N_25893,N_12901,N_14888);
nand U25894 (N_25894,N_11830,N_14763);
and U25895 (N_25895,N_16575,N_15384);
xnor U25896 (N_25896,N_16167,N_13916);
nand U25897 (N_25897,N_15587,N_18974);
and U25898 (N_25898,N_12938,N_15652);
nor U25899 (N_25899,N_16236,N_19185);
xor U25900 (N_25900,N_16743,N_16546);
xor U25901 (N_25901,N_16395,N_10939);
and U25902 (N_25902,N_11613,N_11623);
and U25903 (N_25903,N_15197,N_18467);
and U25904 (N_25904,N_11922,N_11548);
or U25905 (N_25905,N_13958,N_18393);
xor U25906 (N_25906,N_10390,N_11640);
or U25907 (N_25907,N_12475,N_13276);
xor U25908 (N_25908,N_16684,N_18592);
nand U25909 (N_25909,N_17644,N_15493);
and U25910 (N_25910,N_18131,N_10892);
xor U25911 (N_25911,N_12447,N_15418);
nor U25912 (N_25912,N_14899,N_17496);
and U25913 (N_25913,N_16979,N_15808);
or U25914 (N_25914,N_14233,N_16445);
or U25915 (N_25915,N_11126,N_11781);
nor U25916 (N_25916,N_15970,N_17496);
nor U25917 (N_25917,N_18408,N_18519);
or U25918 (N_25918,N_17115,N_14845);
xnor U25919 (N_25919,N_19894,N_19183);
nand U25920 (N_25920,N_10520,N_12204);
nor U25921 (N_25921,N_12654,N_10110);
and U25922 (N_25922,N_19497,N_14118);
nand U25923 (N_25923,N_12117,N_16004);
nand U25924 (N_25924,N_15163,N_19072);
or U25925 (N_25925,N_12343,N_16914);
or U25926 (N_25926,N_12911,N_13199);
and U25927 (N_25927,N_19101,N_16081);
and U25928 (N_25928,N_15566,N_13390);
xor U25929 (N_25929,N_15560,N_13140);
nor U25930 (N_25930,N_18187,N_13031);
or U25931 (N_25931,N_17197,N_16071);
xor U25932 (N_25932,N_18589,N_18212);
nor U25933 (N_25933,N_19252,N_16216);
and U25934 (N_25934,N_18014,N_10717);
xor U25935 (N_25935,N_17102,N_17374);
and U25936 (N_25936,N_10675,N_14308);
or U25937 (N_25937,N_14194,N_10785);
xor U25938 (N_25938,N_19489,N_13316);
nand U25939 (N_25939,N_15311,N_14962);
nand U25940 (N_25940,N_12114,N_19746);
xnor U25941 (N_25941,N_18782,N_15904);
and U25942 (N_25942,N_14075,N_14705);
nand U25943 (N_25943,N_19250,N_11237);
nor U25944 (N_25944,N_13706,N_19126);
nor U25945 (N_25945,N_17861,N_19876);
xnor U25946 (N_25946,N_15842,N_19204);
nand U25947 (N_25947,N_19306,N_11415);
or U25948 (N_25948,N_18237,N_12233);
xnor U25949 (N_25949,N_14137,N_15180);
xnor U25950 (N_25950,N_13968,N_18843);
xor U25951 (N_25951,N_14159,N_18298);
nand U25952 (N_25952,N_12525,N_12438);
and U25953 (N_25953,N_15436,N_14434);
nor U25954 (N_25954,N_15944,N_15517);
xor U25955 (N_25955,N_15812,N_14883);
or U25956 (N_25956,N_18519,N_18534);
nor U25957 (N_25957,N_11305,N_19212);
xor U25958 (N_25958,N_18504,N_19106);
and U25959 (N_25959,N_16606,N_14322);
or U25960 (N_25960,N_14538,N_11547);
or U25961 (N_25961,N_18579,N_15534);
xor U25962 (N_25962,N_18189,N_19971);
and U25963 (N_25963,N_12777,N_15829);
xnor U25964 (N_25964,N_14892,N_14439);
and U25965 (N_25965,N_17125,N_14029);
and U25966 (N_25966,N_10782,N_13103);
nor U25967 (N_25967,N_15069,N_19214);
nor U25968 (N_25968,N_14908,N_14982);
and U25969 (N_25969,N_11865,N_10232);
or U25970 (N_25970,N_13330,N_16851);
or U25971 (N_25971,N_12102,N_16768);
and U25972 (N_25972,N_12682,N_18301);
nand U25973 (N_25973,N_10122,N_13195);
nand U25974 (N_25974,N_17533,N_13344);
nor U25975 (N_25975,N_14545,N_10246);
or U25976 (N_25976,N_12314,N_10092);
nor U25977 (N_25977,N_10819,N_17345);
and U25978 (N_25978,N_17022,N_12163);
or U25979 (N_25979,N_16258,N_15180);
or U25980 (N_25980,N_10597,N_17154);
nor U25981 (N_25981,N_15608,N_17961);
xor U25982 (N_25982,N_12758,N_11812);
and U25983 (N_25983,N_15392,N_12251);
xnor U25984 (N_25984,N_11210,N_13217);
nor U25985 (N_25985,N_14989,N_13403);
or U25986 (N_25986,N_19047,N_18712);
or U25987 (N_25987,N_17320,N_19319);
xnor U25988 (N_25988,N_18160,N_17017);
or U25989 (N_25989,N_14904,N_13026);
nand U25990 (N_25990,N_18005,N_16564);
xnor U25991 (N_25991,N_11325,N_18727);
or U25992 (N_25992,N_18739,N_14588);
nor U25993 (N_25993,N_19967,N_15255);
and U25994 (N_25994,N_17006,N_12777);
xor U25995 (N_25995,N_16135,N_13866);
nor U25996 (N_25996,N_11977,N_14850);
nor U25997 (N_25997,N_13659,N_14435);
xor U25998 (N_25998,N_13098,N_14786);
or U25999 (N_25999,N_14106,N_10507);
nand U26000 (N_26000,N_12075,N_11143);
or U26001 (N_26001,N_15623,N_19513);
xnor U26002 (N_26002,N_13005,N_10243);
and U26003 (N_26003,N_11555,N_12439);
xnor U26004 (N_26004,N_11911,N_11103);
and U26005 (N_26005,N_14760,N_19615);
nand U26006 (N_26006,N_18853,N_14969);
nand U26007 (N_26007,N_17898,N_19981);
nor U26008 (N_26008,N_16223,N_12827);
and U26009 (N_26009,N_12208,N_15461);
nand U26010 (N_26010,N_18624,N_10595);
or U26011 (N_26011,N_18113,N_15609);
nor U26012 (N_26012,N_10358,N_15278);
xnor U26013 (N_26013,N_14727,N_12634);
and U26014 (N_26014,N_15788,N_14566);
nor U26015 (N_26015,N_10792,N_10694);
nor U26016 (N_26016,N_15226,N_15576);
nand U26017 (N_26017,N_18130,N_17865);
xor U26018 (N_26018,N_10938,N_16659);
xnor U26019 (N_26019,N_17825,N_18089);
nand U26020 (N_26020,N_10518,N_18381);
or U26021 (N_26021,N_18680,N_18289);
nor U26022 (N_26022,N_15238,N_19966);
and U26023 (N_26023,N_16744,N_12135);
xnor U26024 (N_26024,N_18634,N_13418);
and U26025 (N_26025,N_10968,N_13642);
or U26026 (N_26026,N_16176,N_17166);
xor U26027 (N_26027,N_15815,N_16385);
nor U26028 (N_26028,N_11264,N_14406);
nor U26029 (N_26029,N_19649,N_18145);
and U26030 (N_26030,N_13800,N_10197);
xor U26031 (N_26031,N_14855,N_15806);
or U26032 (N_26032,N_14581,N_15461);
or U26033 (N_26033,N_19023,N_13779);
and U26034 (N_26034,N_18168,N_13672);
or U26035 (N_26035,N_16589,N_12134);
nor U26036 (N_26036,N_14701,N_12101);
or U26037 (N_26037,N_16786,N_16167);
nand U26038 (N_26038,N_15163,N_17086);
nand U26039 (N_26039,N_10086,N_12445);
xor U26040 (N_26040,N_14820,N_16778);
and U26041 (N_26041,N_19946,N_19231);
or U26042 (N_26042,N_14139,N_19510);
and U26043 (N_26043,N_18625,N_13762);
nor U26044 (N_26044,N_18687,N_16414);
and U26045 (N_26045,N_16204,N_13613);
nand U26046 (N_26046,N_12908,N_11881);
xor U26047 (N_26047,N_13243,N_12321);
and U26048 (N_26048,N_12937,N_10753);
nand U26049 (N_26049,N_13173,N_11035);
and U26050 (N_26050,N_19520,N_10228);
nor U26051 (N_26051,N_10054,N_17838);
nand U26052 (N_26052,N_11972,N_13636);
and U26053 (N_26053,N_11162,N_18583);
xor U26054 (N_26054,N_13238,N_18112);
or U26055 (N_26055,N_13560,N_13854);
and U26056 (N_26056,N_15342,N_14726);
xnor U26057 (N_26057,N_19618,N_17508);
xor U26058 (N_26058,N_12451,N_12343);
and U26059 (N_26059,N_18166,N_14132);
nor U26060 (N_26060,N_16647,N_14978);
xor U26061 (N_26061,N_19143,N_18143);
and U26062 (N_26062,N_14618,N_18308);
xor U26063 (N_26063,N_11957,N_14659);
or U26064 (N_26064,N_17805,N_18274);
and U26065 (N_26065,N_14582,N_16887);
and U26066 (N_26066,N_15249,N_13917);
or U26067 (N_26067,N_15694,N_16729);
or U26068 (N_26068,N_19025,N_18096);
or U26069 (N_26069,N_19398,N_13355);
nor U26070 (N_26070,N_15814,N_18875);
nand U26071 (N_26071,N_13883,N_11231);
nand U26072 (N_26072,N_15868,N_17500);
and U26073 (N_26073,N_16686,N_19807);
or U26074 (N_26074,N_17692,N_11322);
xnor U26075 (N_26075,N_15135,N_19514);
xnor U26076 (N_26076,N_19697,N_15672);
nor U26077 (N_26077,N_10246,N_11528);
xnor U26078 (N_26078,N_18609,N_13861);
xnor U26079 (N_26079,N_18873,N_15170);
nand U26080 (N_26080,N_14135,N_12764);
or U26081 (N_26081,N_11649,N_17716);
xnor U26082 (N_26082,N_15450,N_12940);
nor U26083 (N_26083,N_17546,N_18120);
and U26084 (N_26084,N_12224,N_13896);
nand U26085 (N_26085,N_14821,N_10182);
or U26086 (N_26086,N_16342,N_19603);
or U26087 (N_26087,N_17388,N_15148);
xor U26088 (N_26088,N_13967,N_11278);
or U26089 (N_26089,N_15621,N_12894);
or U26090 (N_26090,N_11378,N_16122);
nor U26091 (N_26091,N_15172,N_14519);
xnor U26092 (N_26092,N_12938,N_18059);
and U26093 (N_26093,N_18880,N_12375);
or U26094 (N_26094,N_19889,N_14767);
xor U26095 (N_26095,N_17506,N_15958);
nand U26096 (N_26096,N_18143,N_10222);
or U26097 (N_26097,N_14766,N_15716);
nor U26098 (N_26098,N_15768,N_13652);
or U26099 (N_26099,N_17686,N_11681);
and U26100 (N_26100,N_17554,N_16862);
and U26101 (N_26101,N_17672,N_14802);
and U26102 (N_26102,N_12071,N_15945);
or U26103 (N_26103,N_15492,N_13169);
xnor U26104 (N_26104,N_14401,N_12991);
or U26105 (N_26105,N_12532,N_19513);
or U26106 (N_26106,N_14568,N_13117);
and U26107 (N_26107,N_10276,N_16782);
xor U26108 (N_26108,N_10661,N_15651);
and U26109 (N_26109,N_13725,N_14721);
nand U26110 (N_26110,N_13198,N_17522);
xnor U26111 (N_26111,N_17860,N_10536);
or U26112 (N_26112,N_11507,N_16185);
nand U26113 (N_26113,N_13859,N_14800);
or U26114 (N_26114,N_12792,N_18433);
or U26115 (N_26115,N_16568,N_14495);
or U26116 (N_26116,N_13684,N_10505);
and U26117 (N_26117,N_16720,N_13433);
and U26118 (N_26118,N_14768,N_12177);
and U26119 (N_26119,N_13130,N_14478);
nand U26120 (N_26120,N_13991,N_16342);
and U26121 (N_26121,N_15374,N_14129);
nand U26122 (N_26122,N_12321,N_18457);
xnor U26123 (N_26123,N_17292,N_18522);
nor U26124 (N_26124,N_17347,N_18073);
or U26125 (N_26125,N_11325,N_11686);
and U26126 (N_26126,N_16952,N_14872);
and U26127 (N_26127,N_15994,N_19450);
nand U26128 (N_26128,N_19136,N_19962);
nand U26129 (N_26129,N_13816,N_12930);
nand U26130 (N_26130,N_15350,N_12915);
or U26131 (N_26131,N_19749,N_15966);
nor U26132 (N_26132,N_12562,N_15310);
and U26133 (N_26133,N_18395,N_17263);
or U26134 (N_26134,N_10678,N_16437);
xor U26135 (N_26135,N_16135,N_19370);
xnor U26136 (N_26136,N_15357,N_16554);
and U26137 (N_26137,N_19602,N_16733);
nand U26138 (N_26138,N_16041,N_13704);
nand U26139 (N_26139,N_18491,N_13783);
and U26140 (N_26140,N_10125,N_19704);
xnor U26141 (N_26141,N_16107,N_12052);
and U26142 (N_26142,N_17995,N_12349);
nand U26143 (N_26143,N_12873,N_16431);
nand U26144 (N_26144,N_16334,N_11050);
nor U26145 (N_26145,N_18825,N_13217);
or U26146 (N_26146,N_15246,N_19738);
and U26147 (N_26147,N_10390,N_10701);
nor U26148 (N_26148,N_19646,N_11257);
or U26149 (N_26149,N_19411,N_14149);
and U26150 (N_26150,N_19463,N_18706);
and U26151 (N_26151,N_16008,N_19846);
and U26152 (N_26152,N_19798,N_18338);
or U26153 (N_26153,N_12902,N_15852);
nand U26154 (N_26154,N_18133,N_17396);
nand U26155 (N_26155,N_19872,N_17405);
nand U26156 (N_26156,N_16049,N_14911);
or U26157 (N_26157,N_13628,N_15231);
nor U26158 (N_26158,N_15557,N_16424);
or U26159 (N_26159,N_10649,N_17394);
nand U26160 (N_26160,N_19903,N_17813);
or U26161 (N_26161,N_14499,N_15668);
nand U26162 (N_26162,N_11515,N_10694);
xnor U26163 (N_26163,N_13259,N_12420);
or U26164 (N_26164,N_19317,N_13588);
and U26165 (N_26165,N_12883,N_13967);
and U26166 (N_26166,N_16581,N_17719);
nand U26167 (N_26167,N_19632,N_10374);
or U26168 (N_26168,N_17599,N_16746);
nor U26169 (N_26169,N_18007,N_15701);
xnor U26170 (N_26170,N_14730,N_11106);
nand U26171 (N_26171,N_19572,N_15314);
or U26172 (N_26172,N_19108,N_17018);
nor U26173 (N_26173,N_18587,N_14443);
and U26174 (N_26174,N_10164,N_15955);
nor U26175 (N_26175,N_19597,N_16926);
xnor U26176 (N_26176,N_15876,N_18494);
and U26177 (N_26177,N_11922,N_14104);
nor U26178 (N_26178,N_15427,N_11184);
nor U26179 (N_26179,N_18348,N_17771);
or U26180 (N_26180,N_10269,N_11270);
xnor U26181 (N_26181,N_13426,N_15931);
and U26182 (N_26182,N_13682,N_19368);
xor U26183 (N_26183,N_13511,N_18675);
xnor U26184 (N_26184,N_17716,N_14642);
nand U26185 (N_26185,N_14451,N_15582);
nor U26186 (N_26186,N_12590,N_18153);
or U26187 (N_26187,N_18158,N_14237);
nand U26188 (N_26188,N_19854,N_10786);
nor U26189 (N_26189,N_12790,N_10253);
nand U26190 (N_26190,N_16587,N_16748);
nand U26191 (N_26191,N_16888,N_16191);
nor U26192 (N_26192,N_11345,N_11867);
and U26193 (N_26193,N_14209,N_18519);
or U26194 (N_26194,N_10009,N_18077);
or U26195 (N_26195,N_17930,N_10901);
nor U26196 (N_26196,N_12589,N_18885);
xnor U26197 (N_26197,N_17823,N_18238);
nor U26198 (N_26198,N_16894,N_15727);
xnor U26199 (N_26199,N_10548,N_10143);
xnor U26200 (N_26200,N_19705,N_10045);
xor U26201 (N_26201,N_12422,N_11097);
nor U26202 (N_26202,N_13277,N_11243);
or U26203 (N_26203,N_14765,N_12101);
xnor U26204 (N_26204,N_16825,N_16958);
xnor U26205 (N_26205,N_18089,N_12132);
nand U26206 (N_26206,N_17472,N_13858);
nand U26207 (N_26207,N_18641,N_11960);
nor U26208 (N_26208,N_11042,N_18796);
nand U26209 (N_26209,N_15618,N_12969);
xor U26210 (N_26210,N_11822,N_10695);
or U26211 (N_26211,N_13567,N_14985);
xnor U26212 (N_26212,N_11706,N_13226);
and U26213 (N_26213,N_12950,N_16326);
and U26214 (N_26214,N_17633,N_11078);
or U26215 (N_26215,N_18914,N_11961);
nand U26216 (N_26216,N_11587,N_12117);
xor U26217 (N_26217,N_18085,N_14749);
nand U26218 (N_26218,N_10901,N_10708);
xnor U26219 (N_26219,N_11004,N_15065);
nor U26220 (N_26220,N_11125,N_16965);
xnor U26221 (N_26221,N_18110,N_16206);
nand U26222 (N_26222,N_12697,N_17741);
xnor U26223 (N_26223,N_14999,N_11884);
nand U26224 (N_26224,N_15303,N_10385);
or U26225 (N_26225,N_16755,N_13946);
and U26226 (N_26226,N_16828,N_18480);
xor U26227 (N_26227,N_14266,N_10126);
and U26228 (N_26228,N_14003,N_10829);
nor U26229 (N_26229,N_18230,N_18250);
nor U26230 (N_26230,N_13564,N_10482);
and U26231 (N_26231,N_19494,N_13136);
xnor U26232 (N_26232,N_11239,N_13155);
xnor U26233 (N_26233,N_17343,N_13737);
nand U26234 (N_26234,N_16344,N_12482);
nand U26235 (N_26235,N_15225,N_18122);
xor U26236 (N_26236,N_11506,N_11261);
nor U26237 (N_26237,N_19892,N_19587);
and U26238 (N_26238,N_14826,N_18901);
nor U26239 (N_26239,N_15947,N_19831);
nor U26240 (N_26240,N_18989,N_13770);
and U26241 (N_26241,N_19382,N_12528);
nand U26242 (N_26242,N_18142,N_11570);
xnor U26243 (N_26243,N_17438,N_11858);
nand U26244 (N_26244,N_10621,N_13658);
nand U26245 (N_26245,N_16354,N_14558);
and U26246 (N_26246,N_10135,N_12319);
nor U26247 (N_26247,N_16803,N_16609);
nor U26248 (N_26248,N_11739,N_13226);
nand U26249 (N_26249,N_14654,N_19076);
and U26250 (N_26250,N_11047,N_11578);
xnor U26251 (N_26251,N_13874,N_14158);
nand U26252 (N_26252,N_11738,N_18578);
or U26253 (N_26253,N_19726,N_10955);
and U26254 (N_26254,N_15446,N_19722);
nand U26255 (N_26255,N_13867,N_16701);
and U26256 (N_26256,N_13975,N_19300);
xor U26257 (N_26257,N_11193,N_17498);
or U26258 (N_26258,N_17355,N_19173);
nand U26259 (N_26259,N_10546,N_15339);
and U26260 (N_26260,N_17048,N_14316);
nor U26261 (N_26261,N_17781,N_16251);
and U26262 (N_26262,N_10799,N_13988);
xnor U26263 (N_26263,N_15855,N_15851);
nor U26264 (N_26264,N_14197,N_16733);
or U26265 (N_26265,N_13592,N_19372);
nand U26266 (N_26266,N_13526,N_18688);
nand U26267 (N_26267,N_10722,N_11631);
or U26268 (N_26268,N_12159,N_11420);
and U26269 (N_26269,N_11351,N_19287);
nor U26270 (N_26270,N_11879,N_18834);
nor U26271 (N_26271,N_10451,N_18513);
nand U26272 (N_26272,N_19807,N_16738);
and U26273 (N_26273,N_18443,N_15868);
xor U26274 (N_26274,N_16654,N_16218);
xnor U26275 (N_26275,N_18193,N_14402);
and U26276 (N_26276,N_16003,N_18946);
nand U26277 (N_26277,N_10616,N_10911);
xnor U26278 (N_26278,N_18974,N_13122);
nand U26279 (N_26279,N_15853,N_16473);
xnor U26280 (N_26280,N_11976,N_14532);
nand U26281 (N_26281,N_19581,N_11220);
and U26282 (N_26282,N_17315,N_13732);
nand U26283 (N_26283,N_12460,N_12500);
xor U26284 (N_26284,N_18937,N_14793);
or U26285 (N_26285,N_14913,N_19298);
or U26286 (N_26286,N_11624,N_18265);
xnor U26287 (N_26287,N_14275,N_19415);
xor U26288 (N_26288,N_19692,N_10374);
or U26289 (N_26289,N_16631,N_18233);
nand U26290 (N_26290,N_16535,N_19330);
nor U26291 (N_26291,N_17450,N_11010);
and U26292 (N_26292,N_16602,N_15048);
and U26293 (N_26293,N_12576,N_15946);
and U26294 (N_26294,N_10701,N_13033);
and U26295 (N_26295,N_12924,N_18940);
xnor U26296 (N_26296,N_11451,N_14075);
or U26297 (N_26297,N_11034,N_15784);
nor U26298 (N_26298,N_17620,N_11034);
and U26299 (N_26299,N_10719,N_18083);
nand U26300 (N_26300,N_19561,N_13922);
xnor U26301 (N_26301,N_12205,N_14027);
xor U26302 (N_26302,N_18152,N_18284);
or U26303 (N_26303,N_14313,N_18643);
and U26304 (N_26304,N_17972,N_15727);
xnor U26305 (N_26305,N_17263,N_13645);
nor U26306 (N_26306,N_10634,N_18541);
xnor U26307 (N_26307,N_15376,N_12896);
or U26308 (N_26308,N_12663,N_12316);
nor U26309 (N_26309,N_18598,N_11403);
nand U26310 (N_26310,N_17825,N_19246);
xnor U26311 (N_26311,N_12678,N_10030);
or U26312 (N_26312,N_18150,N_15159);
or U26313 (N_26313,N_10829,N_10674);
xor U26314 (N_26314,N_11383,N_18292);
nand U26315 (N_26315,N_17683,N_10287);
and U26316 (N_26316,N_14669,N_17038);
nor U26317 (N_26317,N_10361,N_12316);
nand U26318 (N_26318,N_10353,N_18602);
and U26319 (N_26319,N_16929,N_10808);
or U26320 (N_26320,N_13699,N_16317);
or U26321 (N_26321,N_17960,N_14988);
or U26322 (N_26322,N_15956,N_11275);
nand U26323 (N_26323,N_11332,N_19408);
nand U26324 (N_26324,N_10817,N_19538);
and U26325 (N_26325,N_17969,N_10457);
and U26326 (N_26326,N_14784,N_12452);
or U26327 (N_26327,N_14767,N_11989);
nand U26328 (N_26328,N_11180,N_12949);
and U26329 (N_26329,N_14543,N_17147);
nand U26330 (N_26330,N_18061,N_11570);
nand U26331 (N_26331,N_17904,N_10347);
or U26332 (N_26332,N_17096,N_11609);
nand U26333 (N_26333,N_13719,N_16261);
xnor U26334 (N_26334,N_14425,N_11772);
or U26335 (N_26335,N_10899,N_11772);
nand U26336 (N_26336,N_16716,N_19822);
or U26337 (N_26337,N_18576,N_18898);
nand U26338 (N_26338,N_18170,N_10403);
xnor U26339 (N_26339,N_14240,N_17653);
and U26340 (N_26340,N_11682,N_11172);
or U26341 (N_26341,N_16773,N_16997);
xnor U26342 (N_26342,N_10702,N_13769);
nand U26343 (N_26343,N_19481,N_19534);
nor U26344 (N_26344,N_11186,N_14246);
xnor U26345 (N_26345,N_19990,N_14206);
xnor U26346 (N_26346,N_14720,N_19416);
nor U26347 (N_26347,N_15212,N_13259);
nor U26348 (N_26348,N_10380,N_16188);
nor U26349 (N_26349,N_16287,N_12844);
and U26350 (N_26350,N_17723,N_17248);
and U26351 (N_26351,N_19608,N_16196);
nor U26352 (N_26352,N_11132,N_11304);
nor U26353 (N_26353,N_13293,N_14122);
and U26354 (N_26354,N_19336,N_14586);
or U26355 (N_26355,N_18064,N_19171);
or U26356 (N_26356,N_17108,N_18933);
xnor U26357 (N_26357,N_16979,N_18334);
nand U26358 (N_26358,N_11894,N_16175);
or U26359 (N_26359,N_11423,N_13220);
or U26360 (N_26360,N_19757,N_19936);
nor U26361 (N_26361,N_12204,N_19294);
and U26362 (N_26362,N_19175,N_17263);
nor U26363 (N_26363,N_18459,N_13129);
xor U26364 (N_26364,N_17639,N_16291);
nand U26365 (N_26365,N_19533,N_10898);
or U26366 (N_26366,N_16013,N_18270);
nor U26367 (N_26367,N_17990,N_19361);
nor U26368 (N_26368,N_14415,N_13397);
xor U26369 (N_26369,N_14239,N_17407);
nor U26370 (N_26370,N_17079,N_12419);
nand U26371 (N_26371,N_16308,N_19107);
or U26372 (N_26372,N_11104,N_17004);
xor U26373 (N_26373,N_19605,N_10524);
or U26374 (N_26374,N_10864,N_17331);
nand U26375 (N_26375,N_18716,N_10164);
nor U26376 (N_26376,N_13574,N_13811);
xor U26377 (N_26377,N_11938,N_18108);
xor U26378 (N_26378,N_18294,N_13193);
xnor U26379 (N_26379,N_17471,N_10598);
nor U26380 (N_26380,N_19587,N_10868);
xor U26381 (N_26381,N_19181,N_12534);
nand U26382 (N_26382,N_16939,N_13026);
and U26383 (N_26383,N_18298,N_19101);
nand U26384 (N_26384,N_19115,N_14958);
and U26385 (N_26385,N_11784,N_15326);
xnor U26386 (N_26386,N_11388,N_10287);
nor U26387 (N_26387,N_12754,N_10808);
nor U26388 (N_26388,N_15389,N_10282);
xor U26389 (N_26389,N_15985,N_17984);
and U26390 (N_26390,N_12621,N_19954);
or U26391 (N_26391,N_13893,N_11491);
nor U26392 (N_26392,N_10310,N_16870);
or U26393 (N_26393,N_19684,N_15841);
and U26394 (N_26394,N_11199,N_13228);
and U26395 (N_26395,N_13576,N_10091);
or U26396 (N_26396,N_13858,N_12267);
and U26397 (N_26397,N_17343,N_13808);
xor U26398 (N_26398,N_13437,N_11030);
and U26399 (N_26399,N_18016,N_17953);
and U26400 (N_26400,N_17913,N_12810);
or U26401 (N_26401,N_15166,N_10189);
and U26402 (N_26402,N_11404,N_19885);
and U26403 (N_26403,N_13606,N_13821);
xor U26404 (N_26404,N_11551,N_16910);
nand U26405 (N_26405,N_18159,N_19731);
nor U26406 (N_26406,N_15299,N_13319);
xnor U26407 (N_26407,N_12971,N_14074);
and U26408 (N_26408,N_19472,N_10240);
or U26409 (N_26409,N_15320,N_10879);
nand U26410 (N_26410,N_17484,N_14431);
xor U26411 (N_26411,N_15420,N_11240);
nor U26412 (N_26412,N_15502,N_19928);
nor U26413 (N_26413,N_14294,N_16284);
or U26414 (N_26414,N_17988,N_10326);
or U26415 (N_26415,N_16254,N_11631);
nor U26416 (N_26416,N_15898,N_10178);
nor U26417 (N_26417,N_16751,N_18256);
nand U26418 (N_26418,N_14126,N_11841);
or U26419 (N_26419,N_11464,N_16631);
nand U26420 (N_26420,N_16906,N_11821);
and U26421 (N_26421,N_13452,N_12190);
nor U26422 (N_26422,N_14494,N_18945);
nand U26423 (N_26423,N_17755,N_17994);
nor U26424 (N_26424,N_15431,N_15427);
xnor U26425 (N_26425,N_10557,N_15360);
and U26426 (N_26426,N_12117,N_17619);
or U26427 (N_26427,N_13725,N_13819);
or U26428 (N_26428,N_19820,N_10224);
or U26429 (N_26429,N_12184,N_14348);
nand U26430 (N_26430,N_10260,N_10254);
or U26431 (N_26431,N_12751,N_11550);
and U26432 (N_26432,N_18005,N_12236);
nor U26433 (N_26433,N_17126,N_12081);
nand U26434 (N_26434,N_18834,N_16246);
nand U26435 (N_26435,N_12289,N_15502);
xor U26436 (N_26436,N_16565,N_14773);
nor U26437 (N_26437,N_11938,N_19976);
nor U26438 (N_26438,N_11096,N_13449);
nor U26439 (N_26439,N_10196,N_10132);
nor U26440 (N_26440,N_18527,N_15132);
xnor U26441 (N_26441,N_12039,N_14232);
and U26442 (N_26442,N_11384,N_16978);
nor U26443 (N_26443,N_15265,N_18428);
nand U26444 (N_26444,N_10234,N_10428);
nand U26445 (N_26445,N_18437,N_15675);
nor U26446 (N_26446,N_12695,N_14324);
nor U26447 (N_26447,N_11305,N_16903);
and U26448 (N_26448,N_16922,N_15173);
or U26449 (N_26449,N_12205,N_18934);
or U26450 (N_26450,N_16211,N_18829);
or U26451 (N_26451,N_11104,N_15348);
or U26452 (N_26452,N_10751,N_13949);
nand U26453 (N_26453,N_16280,N_19068);
or U26454 (N_26454,N_10170,N_16298);
or U26455 (N_26455,N_11279,N_11115);
nand U26456 (N_26456,N_10785,N_19789);
xnor U26457 (N_26457,N_11645,N_16536);
nor U26458 (N_26458,N_18877,N_12722);
and U26459 (N_26459,N_11604,N_16092);
and U26460 (N_26460,N_19276,N_18501);
and U26461 (N_26461,N_11927,N_10022);
and U26462 (N_26462,N_17232,N_10280);
and U26463 (N_26463,N_19945,N_15615);
or U26464 (N_26464,N_12321,N_16275);
xor U26465 (N_26465,N_15238,N_19388);
or U26466 (N_26466,N_10569,N_11957);
nor U26467 (N_26467,N_14860,N_11379);
nand U26468 (N_26468,N_10628,N_15119);
or U26469 (N_26469,N_10015,N_13930);
nor U26470 (N_26470,N_19081,N_14229);
and U26471 (N_26471,N_17515,N_15198);
or U26472 (N_26472,N_19976,N_12720);
nor U26473 (N_26473,N_13052,N_18441);
and U26474 (N_26474,N_16916,N_11334);
or U26475 (N_26475,N_15959,N_18085);
xor U26476 (N_26476,N_11111,N_15266);
or U26477 (N_26477,N_14241,N_10306);
nand U26478 (N_26478,N_12800,N_17216);
and U26479 (N_26479,N_16909,N_10037);
nor U26480 (N_26480,N_13476,N_15415);
or U26481 (N_26481,N_15686,N_14882);
nand U26482 (N_26482,N_12461,N_18450);
nor U26483 (N_26483,N_15299,N_11140);
and U26484 (N_26484,N_18622,N_18422);
and U26485 (N_26485,N_16884,N_18200);
or U26486 (N_26486,N_13034,N_11053);
or U26487 (N_26487,N_19070,N_12879);
or U26488 (N_26488,N_13123,N_14549);
nor U26489 (N_26489,N_10312,N_14942);
nor U26490 (N_26490,N_19599,N_14553);
or U26491 (N_26491,N_17901,N_14718);
and U26492 (N_26492,N_15704,N_15509);
nand U26493 (N_26493,N_13548,N_11681);
nor U26494 (N_26494,N_12746,N_17131);
or U26495 (N_26495,N_15401,N_13344);
or U26496 (N_26496,N_17791,N_15161);
and U26497 (N_26497,N_19857,N_14766);
nor U26498 (N_26498,N_17969,N_15944);
nand U26499 (N_26499,N_18142,N_19270);
or U26500 (N_26500,N_12084,N_17428);
xnor U26501 (N_26501,N_10974,N_10247);
and U26502 (N_26502,N_15312,N_17077);
nand U26503 (N_26503,N_15637,N_12646);
xnor U26504 (N_26504,N_15139,N_11029);
nand U26505 (N_26505,N_11712,N_10425);
or U26506 (N_26506,N_12718,N_14163);
nand U26507 (N_26507,N_19918,N_12337);
xnor U26508 (N_26508,N_17169,N_12975);
nand U26509 (N_26509,N_15179,N_16873);
and U26510 (N_26510,N_16488,N_16997);
or U26511 (N_26511,N_17236,N_17474);
or U26512 (N_26512,N_10800,N_16604);
and U26513 (N_26513,N_15058,N_16940);
nor U26514 (N_26514,N_15084,N_12137);
or U26515 (N_26515,N_11125,N_10937);
or U26516 (N_26516,N_16284,N_14858);
xor U26517 (N_26517,N_12549,N_17605);
xor U26518 (N_26518,N_16128,N_16614);
nor U26519 (N_26519,N_14272,N_18961);
and U26520 (N_26520,N_14713,N_13306);
and U26521 (N_26521,N_13952,N_16611);
nor U26522 (N_26522,N_18334,N_15643);
and U26523 (N_26523,N_12254,N_15085);
or U26524 (N_26524,N_13369,N_13372);
nand U26525 (N_26525,N_16983,N_12857);
xnor U26526 (N_26526,N_18232,N_12978);
nor U26527 (N_26527,N_12786,N_10581);
nand U26528 (N_26528,N_19433,N_18488);
or U26529 (N_26529,N_12978,N_12687);
nand U26530 (N_26530,N_18349,N_16859);
and U26531 (N_26531,N_15305,N_12103);
or U26532 (N_26532,N_10228,N_10009);
xnor U26533 (N_26533,N_12620,N_14268);
and U26534 (N_26534,N_18727,N_17472);
and U26535 (N_26535,N_18970,N_18870);
xor U26536 (N_26536,N_13749,N_19703);
or U26537 (N_26537,N_15893,N_14029);
nor U26538 (N_26538,N_19658,N_11306);
xnor U26539 (N_26539,N_10781,N_19618);
or U26540 (N_26540,N_12541,N_15965);
or U26541 (N_26541,N_10631,N_19921);
and U26542 (N_26542,N_12477,N_14237);
nand U26543 (N_26543,N_19647,N_12611);
or U26544 (N_26544,N_12657,N_14629);
and U26545 (N_26545,N_18478,N_10423);
or U26546 (N_26546,N_10272,N_10618);
xor U26547 (N_26547,N_13600,N_10683);
nor U26548 (N_26548,N_18074,N_17192);
or U26549 (N_26549,N_13110,N_14128);
or U26550 (N_26550,N_16463,N_13363);
or U26551 (N_26551,N_15246,N_18088);
nor U26552 (N_26552,N_16729,N_13813);
nand U26553 (N_26553,N_19461,N_19147);
nor U26554 (N_26554,N_17587,N_13279);
and U26555 (N_26555,N_10584,N_14828);
and U26556 (N_26556,N_18105,N_15998);
xor U26557 (N_26557,N_12471,N_11027);
nand U26558 (N_26558,N_19589,N_19479);
nor U26559 (N_26559,N_11291,N_12105);
nand U26560 (N_26560,N_10033,N_18995);
nor U26561 (N_26561,N_12667,N_13119);
and U26562 (N_26562,N_10352,N_13211);
nand U26563 (N_26563,N_18797,N_13559);
nand U26564 (N_26564,N_11308,N_18129);
nand U26565 (N_26565,N_12401,N_13034);
or U26566 (N_26566,N_17861,N_16593);
and U26567 (N_26567,N_13655,N_15144);
and U26568 (N_26568,N_16656,N_11767);
or U26569 (N_26569,N_14845,N_19780);
nor U26570 (N_26570,N_14553,N_10379);
nand U26571 (N_26571,N_18083,N_16305);
nor U26572 (N_26572,N_14348,N_17026);
nor U26573 (N_26573,N_16695,N_10889);
and U26574 (N_26574,N_10833,N_13597);
nor U26575 (N_26575,N_10020,N_10722);
and U26576 (N_26576,N_10732,N_12298);
xor U26577 (N_26577,N_17910,N_12390);
nand U26578 (N_26578,N_14519,N_15879);
and U26579 (N_26579,N_11965,N_13702);
xnor U26580 (N_26580,N_13080,N_14133);
nand U26581 (N_26581,N_16031,N_13910);
and U26582 (N_26582,N_11443,N_11463);
and U26583 (N_26583,N_10061,N_11433);
nand U26584 (N_26584,N_10697,N_10508);
or U26585 (N_26585,N_13401,N_11632);
xnor U26586 (N_26586,N_14638,N_18870);
nand U26587 (N_26587,N_18284,N_17286);
xnor U26588 (N_26588,N_15729,N_17920);
xor U26589 (N_26589,N_19577,N_18141);
and U26590 (N_26590,N_18492,N_19797);
xor U26591 (N_26591,N_17745,N_17375);
xor U26592 (N_26592,N_18336,N_17566);
xnor U26593 (N_26593,N_17276,N_15664);
nand U26594 (N_26594,N_17751,N_10131);
xnor U26595 (N_26595,N_12109,N_14663);
or U26596 (N_26596,N_10997,N_15144);
nor U26597 (N_26597,N_16301,N_16133);
or U26598 (N_26598,N_13799,N_14325);
or U26599 (N_26599,N_19879,N_16779);
nor U26600 (N_26600,N_11915,N_18453);
or U26601 (N_26601,N_19397,N_12867);
and U26602 (N_26602,N_19084,N_10511);
or U26603 (N_26603,N_18309,N_10748);
or U26604 (N_26604,N_13889,N_12944);
and U26605 (N_26605,N_17536,N_10488);
nor U26606 (N_26606,N_13346,N_15711);
and U26607 (N_26607,N_14118,N_12475);
nand U26608 (N_26608,N_16038,N_10611);
nand U26609 (N_26609,N_16712,N_16681);
xor U26610 (N_26610,N_15269,N_14337);
or U26611 (N_26611,N_18704,N_16107);
nor U26612 (N_26612,N_10540,N_10808);
or U26613 (N_26613,N_13739,N_13798);
and U26614 (N_26614,N_19442,N_19797);
xor U26615 (N_26615,N_12876,N_17439);
nand U26616 (N_26616,N_12943,N_16216);
nand U26617 (N_26617,N_18868,N_19980);
and U26618 (N_26618,N_12835,N_16510);
nand U26619 (N_26619,N_12248,N_12413);
or U26620 (N_26620,N_14515,N_17077);
xnor U26621 (N_26621,N_17079,N_12914);
xnor U26622 (N_26622,N_10198,N_15644);
xor U26623 (N_26623,N_11973,N_17117);
xor U26624 (N_26624,N_19290,N_13561);
nand U26625 (N_26625,N_18946,N_11221);
or U26626 (N_26626,N_11180,N_19626);
and U26627 (N_26627,N_14843,N_14808);
nand U26628 (N_26628,N_11644,N_16863);
nor U26629 (N_26629,N_13575,N_10745);
nand U26630 (N_26630,N_12644,N_11314);
nor U26631 (N_26631,N_11863,N_10798);
xnor U26632 (N_26632,N_13158,N_19213);
nand U26633 (N_26633,N_11144,N_12219);
and U26634 (N_26634,N_11980,N_19952);
or U26635 (N_26635,N_15545,N_10397);
nor U26636 (N_26636,N_14284,N_14008);
nor U26637 (N_26637,N_15300,N_11225);
and U26638 (N_26638,N_10802,N_16154);
and U26639 (N_26639,N_19072,N_19549);
xnor U26640 (N_26640,N_19668,N_14899);
nor U26641 (N_26641,N_12667,N_14485);
and U26642 (N_26642,N_18308,N_18927);
xor U26643 (N_26643,N_11060,N_19392);
nor U26644 (N_26644,N_16555,N_11701);
and U26645 (N_26645,N_11295,N_19037);
and U26646 (N_26646,N_17415,N_10837);
xnor U26647 (N_26647,N_15462,N_12000);
xor U26648 (N_26648,N_17765,N_15787);
nor U26649 (N_26649,N_14666,N_10563);
xor U26650 (N_26650,N_18153,N_11794);
xor U26651 (N_26651,N_17840,N_15735);
nor U26652 (N_26652,N_19216,N_17520);
xor U26653 (N_26653,N_12505,N_14574);
nor U26654 (N_26654,N_11188,N_17051);
xnor U26655 (N_26655,N_15002,N_16663);
nand U26656 (N_26656,N_15817,N_19428);
nor U26657 (N_26657,N_14118,N_15295);
nand U26658 (N_26658,N_13635,N_13987);
nor U26659 (N_26659,N_12575,N_17169);
and U26660 (N_26660,N_19848,N_10547);
and U26661 (N_26661,N_10540,N_18808);
or U26662 (N_26662,N_15095,N_10465);
and U26663 (N_26663,N_18430,N_14224);
or U26664 (N_26664,N_13728,N_12645);
or U26665 (N_26665,N_14506,N_10421);
nand U26666 (N_26666,N_10053,N_13625);
xnor U26667 (N_26667,N_19280,N_13810);
xor U26668 (N_26668,N_19762,N_11502);
or U26669 (N_26669,N_14276,N_17061);
or U26670 (N_26670,N_17554,N_11891);
nand U26671 (N_26671,N_18405,N_16003);
xnor U26672 (N_26672,N_13067,N_17128);
or U26673 (N_26673,N_12969,N_13918);
or U26674 (N_26674,N_14797,N_19406);
nand U26675 (N_26675,N_18265,N_15594);
nand U26676 (N_26676,N_16626,N_15563);
nor U26677 (N_26677,N_17169,N_18825);
and U26678 (N_26678,N_13646,N_17340);
nand U26679 (N_26679,N_17192,N_13638);
nor U26680 (N_26680,N_16037,N_10834);
or U26681 (N_26681,N_17849,N_13785);
and U26682 (N_26682,N_19125,N_13633);
nand U26683 (N_26683,N_14802,N_13767);
nand U26684 (N_26684,N_17460,N_11165);
xnor U26685 (N_26685,N_17476,N_14964);
nor U26686 (N_26686,N_16275,N_18152);
or U26687 (N_26687,N_11459,N_12410);
nand U26688 (N_26688,N_12905,N_13228);
and U26689 (N_26689,N_14467,N_17013);
and U26690 (N_26690,N_19226,N_11618);
and U26691 (N_26691,N_11875,N_12013);
xnor U26692 (N_26692,N_18080,N_12049);
nand U26693 (N_26693,N_13051,N_14086);
nand U26694 (N_26694,N_18196,N_19038);
xor U26695 (N_26695,N_10103,N_19915);
nand U26696 (N_26696,N_10922,N_17627);
or U26697 (N_26697,N_12288,N_17895);
or U26698 (N_26698,N_19418,N_14548);
and U26699 (N_26699,N_16511,N_12422);
xnor U26700 (N_26700,N_11541,N_15367);
nor U26701 (N_26701,N_18989,N_19687);
nor U26702 (N_26702,N_17740,N_13168);
or U26703 (N_26703,N_11675,N_17461);
or U26704 (N_26704,N_18666,N_14538);
nor U26705 (N_26705,N_16938,N_18243);
xor U26706 (N_26706,N_13201,N_13847);
xnor U26707 (N_26707,N_16466,N_11997);
or U26708 (N_26708,N_17202,N_10748);
xnor U26709 (N_26709,N_19378,N_17033);
xor U26710 (N_26710,N_13212,N_11887);
xor U26711 (N_26711,N_15498,N_14119);
or U26712 (N_26712,N_13603,N_14844);
nor U26713 (N_26713,N_16332,N_12891);
and U26714 (N_26714,N_11896,N_12994);
nand U26715 (N_26715,N_16595,N_15289);
and U26716 (N_26716,N_18866,N_15707);
or U26717 (N_26717,N_15746,N_15968);
and U26718 (N_26718,N_18741,N_12398);
xor U26719 (N_26719,N_10213,N_17660);
nand U26720 (N_26720,N_11681,N_11524);
xnor U26721 (N_26721,N_14531,N_19917);
and U26722 (N_26722,N_13276,N_19706);
and U26723 (N_26723,N_11522,N_15951);
nor U26724 (N_26724,N_17488,N_19055);
nand U26725 (N_26725,N_14995,N_12774);
nand U26726 (N_26726,N_17064,N_16583);
nand U26727 (N_26727,N_18889,N_13353);
or U26728 (N_26728,N_14410,N_19400);
and U26729 (N_26729,N_16741,N_11086);
nand U26730 (N_26730,N_10861,N_12029);
nand U26731 (N_26731,N_15442,N_10322);
or U26732 (N_26732,N_16218,N_10491);
nor U26733 (N_26733,N_13179,N_10758);
nand U26734 (N_26734,N_16112,N_18382);
nand U26735 (N_26735,N_18843,N_17990);
nand U26736 (N_26736,N_15776,N_12386);
or U26737 (N_26737,N_12944,N_11399);
nand U26738 (N_26738,N_17822,N_12784);
nor U26739 (N_26739,N_11770,N_18697);
or U26740 (N_26740,N_12467,N_11647);
and U26741 (N_26741,N_18028,N_13175);
nor U26742 (N_26742,N_13509,N_16695);
and U26743 (N_26743,N_13532,N_10475);
nand U26744 (N_26744,N_13972,N_11899);
nand U26745 (N_26745,N_11494,N_19920);
and U26746 (N_26746,N_11515,N_11135);
nand U26747 (N_26747,N_14959,N_19730);
and U26748 (N_26748,N_19129,N_18212);
and U26749 (N_26749,N_10432,N_10722);
and U26750 (N_26750,N_14384,N_11182);
nor U26751 (N_26751,N_17070,N_14173);
nor U26752 (N_26752,N_10763,N_16431);
nand U26753 (N_26753,N_15220,N_19943);
and U26754 (N_26754,N_14484,N_16038);
nor U26755 (N_26755,N_13222,N_13053);
and U26756 (N_26756,N_14010,N_15789);
nand U26757 (N_26757,N_15204,N_13133);
and U26758 (N_26758,N_13978,N_18347);
and U26759 (N_26759,N_16820,N_11415);
and U26760 (N_26760,N_15185,N_13133);
nor U26761 (N_26761,N_11393,N_18066);
nand U26762 (N_26762,N_15558,N_13107);
and U26763 (N_26763,N_19181,N_15794);
nand U26764 (N_26764,N_11720,N_18914);
nand U26765 (N_26765,N_17648,N_19613);
nand U26766 (N_26766,N_18411,N_17813);
or U26767 (N_26767,N_17537,N_15732);
or U26768 (N_26768,N_13830,N_13342);
nor U26769 (N_26769,N_12035,N_14944);
and U26770 (N_26770,N_16935,N_12457);
or U26771 (N_26771,N_14744,N_12324);
nor U26772 (N_26772,N_16833,N_12591);
nor U26773 (N_26773,N_11929,N_19394);
nand U26774 (N_26774,N_19937,N_19274);
nor U26775 (N_26775,N_14067,N_16945);
and U26776 (N_26776,N_13423,N_11857);
nor U26777 (N_26777,N_16044,N_10418);
nand U26778 (N_26778,N_13790,N_11166);
xor U26779 (N_26779,N_13544,N_11183);
xnor U26780 (N_26780,N_11974,N_17062);
nor U26781 (N_26781,N_15295,N_14731);
xor U26782 (N_26782,N_11314,N_19390);
nand U26783 (N_26783,N_13237,N_16183);
nor U26784 (N_26784,N_16195,N_17720);
or U26785 (N_26785,N_19512,N_16353);
nand U26786 (N_26786,N_10035,N_13610);
or U26787 (N_26787,N_14811,N_15777);
and U26788 (N_26788,N_18332,N_18380);
nand U26789 (N_26789,N_16333,N_10105);
and U26790 (N_26790,N_16477,N_14008);
or U26791 (N_26791,N_11707,N_17254);
xnor U26792 (N_26792,N_12610,N_12695);
nor U26793 (N_26793,N_14975,N_11827);
and U26794 (N_26794,N_10508,N_17175);
xor U26795 (N_26795,N_10412,N_12865);
and U26796 (N_26796,N_12048,N_14956);
nor U26797 (N_26797,N_12281,N_17284);
nand U26798 (N_26798,N_15278,N_10955);
and U26799 (N_26799,N_12090,N_19532);
and U26800 (N_26800,N_19344,N_11847);
nor U26801 (N_26801,N_17734,N_16015);
nor U26802 (N_26802,N_19141,N_15307);
nor U26803 (N_26803,N_10024,N_17923);
nand U26804 (N_26804,N_13156,N_17502);
nor U26805 (N_26805,N_10996,N_11305);
and U26806 (N_26806,N_11776,N_14672);
or U26807 (N_26807,N_17459,N_19687);
nor U26808 (N_26808,N_12032,N_11561);
and U26809 (N_26809,N_16286,N_10517);
xor U26810 (N_26810,N_17820,N_13980);
or U26811 (N_26811,N_19567,N_18267);
nor U26812 (N_26812,N_14818,N_17528);
nor U26813 (N_26813,N_15130,N_15101);
nand U26814 (N_26814,N_15727,N_17954);
xnor U26815 (N_26815,N_13928,N_19959);
nor U26816 (N_26816,N_18846,N_11520);
or U26817 (N_26817,N_10410,N_15762);
nor U26818 (N_26818,N_17903,N_15165);
and U26819 (N_26819,N_18968,N_18809);
nor U26820 (N_26820,N_10214,N_18006);
nand U26821 (N_26821,N_13871,N_19744);
or U26822 (N_26822,N_13807,N_19262);
nor U26823 (N_26823,N_17865,N_18468);
and U26824 (N_26824,N_16684,N_19835);
xor U26825 (N_26825,N_13832,N_12331);
nand U26826 (N_26826,N_10966,N_18969);
xor U26827 (N_26827,N_15276,N_18531);
nand U26828 (N_26828,N_14802,N_10452);
nor U26829 (N_26829,N_16540,N_11163);
nor U26830 (N_26830,N_19890,N_17023);
or U26831 (N_26831,N_16388,N_19010);
and U26832 (N_26832,N_15455,N_16780);
and U26833 (N_26833,N_17929,N_16076);
and U26834 (N_26834,N_15802,N_19357);
xnor U26835 (N_26835,N_17974,N_11881);
nor U26836 (N_26836,N_16250,N_18553);
nand U26837 (N_26837,N_17395,N_14643);
or U26838 (N_26838,N_19131,N_11867);
xor U26839 (N_26839,N_18744,N_14753);
or U26840 (N_26840,N_18304,N_12751);
or U26841 (N_26841,N_13784,N_18616);
or U26842 (N_26842,N_16807,N_17565);
or U26843 (N_26843,N_16441,N_11495);
or U26844 (N_26844,N_17146,N_15806);
xnor U26845 (N_26845,N_11117,N_12068);
xnor U26846 (N_26846,N_15539,N_16547);
nor U26847 (N_26847,N_14680,N_17067);
nand U26848 (N_26848,N_11229,N_15215);
and U26849 (N_26849,N_17385,N_12026);
nor U26850 (N_26850,N_14299,N_14452);
nand U26851 (N_26851,N_18461,N_11035);
nor U26852 (N_26852,N_19265,N_13341);
and U26853 (N_26853,N_10137,N_19203);
nand U26854 (N_26854,N_11854,N_14024);
nor U26855 (N_26855,N_14415,N_11117);
nor U26856 (N_26856,N_13686,N_13484);
and U26857 (N_26857,N_13570,N_19293);
and U26858 (N_26858,N_19938,N_15738);
nor U26859 (N_26859,N_19551,N_16461);
xnor U26860 (N_26860,N_18181,N_10294);
nand U26861 (N_26861,N_18481,N_10967);
and U26862 (N_26862,N_10587,N_16249);
xnor U26863 (N_26863,N_10509,N_18794);
or U26864 (N_26864,N_12439,N_18481);
and U26865 (N_26865,N_17373,N_12855);
or U26866 (N_26866,N_12299,N_12003);
nand U26867 (N_26867,N_16826,N_14381);
nand U26868 (N_26868,N_12420,N_14363);
nand U26869 (N_26869,N_11730,N_15847);
xor U26870 (N_26870,N_13719,N_10575);
or U26871 (N_26871,N_16608,N_11937);
nand U26872 (N_26872,N_18026,N_10541);
and U26873 (N_26873,N_12708,N_15846);
nand U26874 (N_26874,N_13808,N_19787);
xnor U26875 (N_26875,N_17859,N_12702);
nand U26876 (N_26876,N_19210,N_18781);
nor U26877 (N_26877,N_16317,N_14016);
xor U26878 (N_26878,N_13887,N_12987);
xor U26879 (N_26879,N_18703,N_11954);
or U26880 (N_26880,N_11702,N_16916);
or U26881 (N_26881,N_18951,N_18985);
nand U26882 (N_26882,N_17269,N_15338);
nand U26883 (N_26883,N_16714,N_16986);
nand U26884 (N_26884,N_15694,N_15361);
nand U26885 (N_26885,N_17186,N_11197);
nand U26886 (N_26886,N_17654,N_11751);
xor U26887 (N_26887,N_17393,N_13560);
or U26888 (N_26888,N_14920,N_18648);
and U26889 (N_26889,N_16894,N_16235);
and U26890 (N_26890,N_10800,N_17532);
xnor U26891 (N_26891,N_15389,N_10294);
or U26892 (N_26892,N_10692,N_14857);
or U26893 (N_26893,N_17303,N_16607);
nand U26894 (N_26894,N_10140,N_12098);
xnor U26895 (N_26895,N_19107,N_14373);
xnor U26896 (N_26896,N_14818,N_19320);
nand U26897 (N_26897,N_10265,N_11952);
nand U26898 (N_26898,N_15606,N_16106);
xnor U26899 (N_26899,N_17727,N_10884);
nor U26900 (N_26900,N_12707,N_14521);
nor U26901 (N_26901,N_16194,N_10373);
and U26902 (N_26902,N_16164,N_15010);
nand U26903 (N_26903,N_18901,N_11170);
or U26904 (N_26904,N_13498,N_12383);
nand U26905 (N_26905,N_11757,N_16801);
nor U26906 (N_26906,N_16230,N_11942);
xnor U26907 (N_26907,N_13769,N_13574);
nor U26908 (N_26908,N_18805,N_19402);
or U26909 (N_26909,N_15186,N_11609);
xor U26910 (N_26910,N_16067,N_17835);
xor U26911 (N_26911,N_11787,N_12847);
nor U26912 (N_26912,N_17338,N_15818);
and U26913 (N_26913,N_16117,N_13416);
and U26914 (N_26914,N_16709,N_16055);
nand U26915 (N_26915,N_12345,N_19256);
xnor U26916 (N_26916,N_19554,N_14452);
nand U26917 (N_26917,N_14198,N_15202);
and U26918 (N_26918,N_15732,N_14469);
nand U26919 (N_26919,N_17438,N_13325);
xnor U26920 (N_26920,N_14046,N_16592);
nor U26921 (N_26921,N_11319,N_17927);
nor U26922 (N_26922,N_18509,N_16060);
or U26923 (N_26923,N_17365,N_12421);
xor U26924 (N_26924,N_15759,N_16885);
xnor U26925 (N_26925,N_13438,N_12959);
xnor U26926 (N_26926,N_17702,N_16196);
or U26927 (N_26927,N_13743,N_10354);
xnor U26928 (N_26928,N_17376,N_15945);
or U26929 (N_26929,N_10558,N_10519);
nand U26930 (N_26930,N_17861,N_15900);
nand U26931 (N_26931,N_11274,N_16879);
and U26932 (N_26932,N_17770,N_15737);
or U26933 (N_26933,N_18098,N_15691);
nand U26934 (N_26934,N_18108,N_13728);
nand U26935 (N_26935,N_14240,N_10767);
xor U26936 (N_26936,N_15284,N_14997);
nor U26937 (N_26937,N_18048,N_10229);
nand U26938 (N_26938,N_10249,N_12255);
nor U26939 (N_26939,N_14141,N_13178);
and U26940 (N_26940,N_17274,N_15745);
nand U26941 (N_26941,N_13491,N_12415);
xnor U26942 (N_26942,N_15347,N_12944);
nor U26943 (N_26943,N_12819,N_16176);
nand U26944 (N_26944,N_11878,N_19704);
nor U26945 (N_26945,N_17385,N_17260);
nand U26946 (N_26946,N_14786,N_19523);
xor U26947 (N_26947,N_10217,N_14961);
or U26948 (N_26948,N_15579,N_16798);
xnor U26949 (N_26949,N_10836,N_11820);
nor U26950 (N_26950,N_12448,N_11607);
nor U26951 (N_26951,N_12728,N_12715);
or U26952 (N_26952,N_12948,N_14827);
and U26953 (N_26953,N_11734,N_11114);
xor U26954 (N_26954,N_13720,N_16662);
nor U26955 (N_26955,N_15967,N_18383);
or U26956 (N_26956,N_11227,N_11564);
nor U26957 (N_26957,N_15444,N_15001);
nor U26958 (N_26958,N_19396,N_16461);
xor U26959 (N_26959,N_18219,N_10954);
nand U26960 (N_26960,N_12702,N_14700);
nor U26961 (N_26961,N_14755,N_10452);
and U26962 (N_26962,N_16202,N_17169);
xnor U26963 (N_26963,N_19821,N_15303);
nand U26964 (N_26964,N_14529,N_18912);
and U26965 (N_26965,N_16170,N_10289);
and U26966 (N_26966,N_12335,N_15900);
xnor U26967 (N_26967,N_12610,N_14916);
nor U26968 (N_26968,N_11932,N_17910);
nor U26969 (N_26969,N_13770,N_17224);
or U26970 (N_26970,N_13861,N_11710);
xor U26971 (N_26971,N_13238,N_13045);
nor U26972 (N_26972,N_11948,N_10462);
nand U26973 (N_26973,N_17281,N_19244);
nor U26974 (N_26974,N_16890,N_11768);
nor U26975 (N_26975,N_19192,N_16241);
xnor U26976 (N_26976,N_14907,N_18625);
nand U26977 (N_26977,N_15186,N_16711);
xnor U26978 (N_26978,N_10806,N_13262);
and U26979 (N_26979,N_16652,N_13615);
nand U26980 (N_26980,N_15986,N_18216);
xnor U26981 (N_26981,N_17383,N_19955);
and U26982 (N_26982,N_14913,N_11861);
nor U26983 (N_26983,N_13954,N_17997);
and U26984 (N_26984,N_18711,N_18305);
nand U26985 (N_26985,N_17283,N_18328);
nor U26986 (N_26986,N_17523,N_13603);
or U26987 (N_26987,N_16412,N_12628);
or U26988 (N_26988,N_11787,N_13072);
or U26989 (N_26989,N_11113,N_16733);
and U26990 (N_26990,N_11001,N_11916);
or U26991 (N_26991,N_14480,N_12027);
or U26992 (N_26992,N_16935,N_14436);
or U26993 (N_26993,N_13545,N_19713);
nor U26994 (N_26994,N_14624,N_14273);
nand U26995 (N_26995,N_19273,N_12863);
and U26996 (N_26996,N_19732,N_10554);
or U26997 (N_26997,N_13016,N_17152);
nand U26998 (N_26998,N_14476,N_14334);
or U26999 (N_26999,N_16693,N_17446);
nor U27000 (N_27000,N_17598,N_13376);
nand U27001 (N_27001,N_19691,N_12536);
xor U27002 (N_27002,N_12789,N_12875);
xor U27003 (N_27003,N_10299,N_12847);
and U27004 (N_27004,N_16741,N_14415);
xor U27005 (N_27005,N_15543,N_19214);
nor U27006 (N_27006,N_18057,N_14965);
and U27007 (N_27007,N_11146,N_12345);
nand U27008 (N_27008,N_13117,N_13849);
and U27009 (N_27009,N_15536,N_13950);
xnor U27010 (N_27010,N_13827,N_19273);
or U27011 (N_27011,N_17536,N_17648);
or U27012 (N_27012,N_10476,N_13838);
nand U27013 (N_27013,N_18310,N_16512);
or U27014 (N_27014,N_19709,N_17785);
nand U27015 (N_27015,N_11582,N_18678);
or U27016 (N_27016,N_17513,N_13315);
nand U27017 (N_27017,N_10073,N_19447);
nor U27018 (N_27018,N_11708,N_14452);
nor U27019 (N_27019,N_10619,N_12281);
xnor U27020 (N_27020,N_16676,N_15387);
xor U27021 (N_27021,N_11244,N_13849);
xnor U27022 (N_27022,N_18913,N_14503);
or U27023 (N_27023,N_11996,N_16156);
nor U27024 (N_27024,N_14530,N_10944);
or U27025 (N_27025,N_17247,N_13363);
xor U27026 (N_27026,N_18876,N_13283);
xor U27027 (N_27027,N_13900,N_12879);
and U27028 (N_27028,N_12272,N_19868);
nand U27029 (N_27029,N_10009,N_13313);
and U27030 (N_27030,N_13208,N_14571);
or U27031 (N_27031,N_15427,N_17907);
and U27032 (N_27032,N_15327,N_14196);
nand U27033 (N_27033,N_11883,N_17423);
or U27034 (N_27034,N_13119,N_17718);
nor U27035 (N_27035,N_15409,N_11331);
nand U27036 (N_27036,N_19030,N_10710);
nor U27037 (N_27037,N_13869,N_12792);
or U27038 (N_27038,N_18551,N_11789);
nand U27039 (N_27039,N_19437,N_19914);
nand U27040 (N_27040,N_18119,N_12374);
nand U27041 (N_27041,N_12031,N_13577);
or U27042 (N_27042,N_17378,N_16921);
xnor U27043 (N_27043,N_11223,N_14342);
xnor U27044 (N_27044,N_14483,N_10012);
and U27045 (N_27045,N_14032,N_12632);
nor U27046 (N_27046,N_12016,N_15456);
nand U27047 (N_27047,N_15300,N_16107);
and U27048 (N_27048,N_19302,N_12170);
and U27049 (N_27049,N_15072,N_11664);
or U27050 (N_27050,N_13186,N_18833);
xor U27051 (N_27051,N_19531,N_11768);
and U27052 (N_27052,N_19268,N_11782);
nor U27053 (N_27053,N_13991,N_18922);
or U27054 (N_27054,N_10831,N_13473);
or U27055 (N_27055,N_10641,N_12968);
and U27056 (N_27056,N_13199,N_12648);
nand U27057 (N_27057,N_12388,N_16135);
nand U27058 (N_27058,N_13200,N_13261);
and U27059 (N_27059,N_19913,N_19576);
or U27060 (N_27060,N_14443,N_18410);
and U27061 (N_27061,N_16483,N_13157);
xor U27062 (N_27062,N_12607,N_10754);
and U27063 (N_27063,N_11420,N_16121);
nor U27064 (N_27064,N_19551,N_13308);
nand U27065 (N_27065,N_18216,N_12556);
or U27066 (N_27066,N_17952,N_10577);
and U27067 (N_27067,N_11976,N_17257);
nand U27068 (N_27068,N_19006,N_18333);
or U27069 (N_27069,N_11127,N_13720);
xor U27070 (N_27070,N_10911,N_18093);
nand U27071 (N_27071,N_19249,N_10308);
and U27072 (N_27072,N_16550,N_16782);
nand U27073 (N_27073,N_15582,N_19180);
and U27074 (N_27074,N_12705,N_13358);
nand U27075 (N_27075,N_14792,N_16479);
nor U27076 (N_27076,N_19987,N_12691);
xnor U27077 (N_27077,N_11597,N_18443);
nor U27078 (N_27078,N_13335,N_17908);
xor U27079 (N_27079,N_18825,N_18312);
and U27080 (N_27080,N_17927,N_11933);
or U27081 (N_27081,N_16326,N_14817);
and U27082 (N_27082,N_19434,N_17668);
xnor U27083 (N_27083,N_11488,N_14512);
nand U27084 (N_27084,N_14594,N_19418);
nor U27085 (N_27085,N_15021,N_11405);
or U27086 (N_27086,N_12359,N_12859);
or U27087 (N_27087,N_18961,N_12080);
or U27088 (N_27088,N_18583,N_11604);
nor U27089 (N_27089,N_18745,N_19323);
and U27090 (N_27090,N_13064,N_14910);
xor U27091 (N_27091,N_15481,N_16508);
nand U27092 (N_27092,N_16981,N_17812);
and U27093 (N_27093,N_16534,N_16843);
nor U27094 (N_27094,N_18002,N_14413);
or U27095 (N_27095,N_16436,N_19767);
or U27096 (N_27096,N_18378,N_11648);
or U27097 (N_27097,N_13880,N_15534);
and U27098 (N_27098,N_15505,N_12316);
nor U27099 (N_27099,N_19603,N_10328);
nor U27100 (N_27100,N_11226,N_16246);
or U27101 (N_27101,N_16565,N_14907);
xnor U27102 (N_27102,N_17799,N_15359);
nand U27103 (N_27103,N_14635,N_18152);
nand U27104 (N_27104,N_13989,N_16000);
or U27105 (N_27105,N_19982,N_10369);
and U27106 (N_27106,N_19025,N_16032);
xnor U27107 (N_27107,N_17561,N_11568);
or U27108 (N_27108,N_10659,N_13852);
or U27109 (N_27109,N_15729,N_11215);
nor U27110 (N_27110,N_13380,N_13851);
xnor U27111 (N_27111,N_12018,N_14595);
or U27112 (N_27112,N_19855,N_13093);
xor U27113 (N_27113,N_14278,N_15179);
and U27114 (N_27114,N_18134,N_17603);
nor U27115 (N_27115,N_16865,N_18303);
and U27116 (N_27116,N_10904,N_17163);
nand U27117 (N_27117,N_17568,N_11637);
nand U27118 (N_27118,N_16473,N_17356);
nor U27119 (N_27119,N_16396,N_16618);
xnor U27120 (N_27120,N_12287,N_18732);
nor U27121 (N_27121,N_14539,N_19743);
xnor U27122 (N_27122,N_19083,N_16439);
and U27123 (N_27123,N_15759,N_18001);
nand U27124 (N_27124,N_14811,N_17788);
or U27125 (N_27125,N_13243,N_15486);
xor U27126 (N_27126,N_10650,N_14463);
or U27127 (N_27127,N_17967,N_19378);
and U27128 (N_27128,N_11570,N_10972);
nor U27129 (N_27129,N_16818,N_19195);
nand U27130 (N_27130,N_12733,N_12329);
nor U27131 (N_27131,N_10861,N_17411);
or U27132 (N_27132,N_17990,N_14919);
nor U27133 (N_27133,N_18312,N_18278);
xnor U27134 (N_27134,N_19364,N_10173);
or U27135 (N_27135,N_10956,N_14948);
nand U27136 (N_27136,N_15935,N_19277);
xor U27137 (N_27137,N_17502,N_14263);
and U27138 (N_27138,N_16709,N_14936);
or U27139 (N_27139,N_18589,N_17658);
or U27140 (N_27140,N_17275,N_11181);
or U27141 (N_27141,N_17883,N_18288);
nand U27142 (N_27142,N_15093,N_12941);
nor U27143 (N_27143,N_10166,N_10640);
and U27144 (N_27144,N_14505,N_15796);
nand U27145 (N_27145,N_19628,N_16159);
xnor U27146 (N_27146,N_12123,N_16714);
nor U27147 (N_27147,N_19010,N_11110);
and U27148 (N_27148,N_19296,N_13349);
nor U27149 (N_27149,N_11368,N_16645);
or U27150 (N_27150,N_10343,N_14454);
or U27151 (N_27151,N_11577,N_13840);
xnor U27152 (N_27152,N_11034,N_19852);
or U27153 (N_27153,N_17202,N_15268);
or U27154 (N_27154,N_10311,N_12763);
and U27155 (N_27155,N_11598,N_12017);
xnor U27156 (N_27156,N_19079,N_17743);
and U27157 (N_27157,N_15128,N_12844);
or U27158 (N_27158,N_15875,N_19782);
nand U27159 (N_27159,N_18082,N_18300);
and U27160 (N_27160,N_14632,N_16091);
nand U27161 (N_27161,N_17990,N_11364);
nand U27162 (N_27162,N_17144,N_16258);
xnor U27163 (N_27163,N_16707,N_14547);
nor U27164 (N_27164,N_17375,N_10403);
or U27165 (N_27165,N_14339,N_14896);
or U27166 (N_27166,N_10109,N_15398);
nand U27167 (N_27167,N_16839,N_16048);
or U27168 (N_27168,N_16507,N_10457);
or U27169 (N_27169,N_16331,N_19922);
xnor U27170 (N_27170,N_13136,N_10127);
and U27171 (N_27171,N_18381,N_17893);
nand U27172 (N_27172,N_16251,N_19985);
nor U27173 (N_27173,N_15622,N_19382);
or U27174 (N_27174,N_15833,N_16396);
nand U27175 (N_27175,N_14911,N_13044);
xor U27176 (N_27176,N_17572,N_17618);
xor U27177 (N_27177,N_19069,N_15361);
or U27178 (N_27178,N_10487,N_17004);
and U27179 (N_27179,N_11795,N_19064);
or U27180 (N_27180,N_19162,N_13232);
nand U27181 (N_27181,N_13048,N_15121);
and U27182 (N_27182,N_14806,N_12934);
nand U27183 (N_27183,N_11768,N_19583);
or U27184 (N_27184,N_14372,N_18270);
or U27185 (N_27185,N_19580,N_12340);
nor U27186 (N_27186,N_10090,N_10253);
nand U27187 (N_27187,N_13603,N_12512);
and U27188 (N_27188,N_18744,N_15076);
nand U27189 (N_27189,N_10081,N_15457);
or U27190 (N_27190,N_13122,N_17355);
and U27191 (N_27191,N_18824,N_19569);
and U27192 (N_27192,N_12394,N_17025);
nor U27193 (N_27193,N_15311,N_16287);
xnor U27194 (N_27194,N_13690,N_16072);
and U27195 (N_27195,N_11936,N_19548);
or U27196 (N_27196,N_18585,N_12937);
and U27197 (N_27197,N_19683,N_18436);
nand U27198 (N_27198,N_11649,N_14866);
and U27199 (N_27199,N_14176,N_11328);
xor U27200 (N_27200,N_19329,N_10478);
nand U27201 (N_27201,N_19178,N_17231);
or U27202 (N_27202,N_17129,N_11656);
and U27203 (N_27203,N_14996,N_16255);
or U27204 (N_27204,N_13589,N_16573);
nor U27205 (N_27205,N_13700,N_11870);
xnor U27206 (N_27206,N_17089,N_15451);
or U27207 (N_27207,N_10741,N_16667);
or U27208 (N_27208,N_17023,N_10258);
nand U27209 (N_27209,N_19355,N_14514);
nand U27210 (N_27210,N_18046,N_12233);
nand U27211 (N_27211,N_10814,N_17794);
xor U27212 (N_27212,N_17932,N_16867);
nand U27213 (N_27213,N_15489,N_11065);
and U27214 (N_27214,N_14548,N_19972);
xor U27215 (N_27215,N_16525,N_14595);
or U27216 (N_27216,N_10968,N_13585);
and U27217 (N_27217,N_15585,N_10885);
or U27218 (N_27218,N_17655,N_13931);
or U27219 (N_27219,N_19930,N_10833);
nand U27220 (N_27220,N_18607,N_13593);
nor U27221 (N_27221,N_18007,N_17105);
and U27222 (N_27222,N_15800,N_15267);
and U27223 (N_27223,N_19863,N_10386);
or U27224 (N_27224,N_16551,N_19241);
nand U27225 (N_27225,N_13100,N_13321);
and U27226 (N_27226,N_12003,N_14173);
or U27227 (N_27227,N_16513,N_14441);
and U27228 (N_27228,N_16283,N_12662);
xnor U27229 (N_27229,N_15695,N_11905);
or U27230 (N_27230,N_14772,N_15662);
nand U27231 (N_27231,N_17161,N_14600);
and U27232 (N_27232,N_15533,N_19894);
or U27233 (N_27233,N_11426,N_17508);
and U27234 (N_27234,N_18869,N_10181);
nand U27235 (N_27235,N_17755,N_11995);
xnor U27236 (N_27236,N_15889,N_16449);
and U27237 (N_27237,N_12144,N_18068);
nand U27238 (N_27238,N_15360,N_10545);
and U27239 (N_27239,N_15999,N_11198);
or U27240 (N_27240,N_14213,N_17254);
xor U27241 (N_27241,N_12228,N_10526);
and U27242 (N_27242,N_19292,N_15929);
or U27243 (N_27243,N_10045,N_10921);
xor U27244 (N_27244,N_15338,N_12914);
xor U27245 (N_27245,N_16224,N_14515);
and U27246 (N_27246,N_14534,N_12707);
or U27247 (N_27247,N_11003,N_16185);
and U27248 (N_27248,N_16871,N_19789);
or U27249 (N_27249,N_19943,N_19646);
or U27250 (N_27250,N_15262,N_13799);
nor U27251 (N_27251,N_16562,N_16387);
xnor U27252 (N_27252,N_12698,N_16198);
nor U27253 (N_27253,N_14943,N_18352);
nor U27254 (N_27254,N_17647,N_10264);
xor U27255 (N_27255,N_15365,N_14676);
nor U27256 (N_27256,N_15539,N_13226);
and U27257 (N_27257,N_17207,N_13170);
nor U27258 (N_27258,N_13835,N_10474);
nor U27259 (N_27259,N_10010,N_12019);
xor U27260 (N_27260,N_19531,N_19501);
nand U27261 (N_27261,N_18776,N_10250);
or U27262 (N_27262,N_17494,N_18810);
nand U27263 (N_27263,N_19686,N_19157);
nand U27264 (N_27264,N_15577,N_14825);
xor U27265 (N_27265,N_18275,N_19729);
and U27266 (N_27266,N_13273,N_14007);
or U27267 (N_27267,N_13521,N_19022);
and U27268 (N_27268,N_13779,N_12867);
and U27269 (N_27269,N_10666,N_15758);
and U27270 (N_27270,N_13499,N_19439);
or U27271 (N_27271,N_18630,N_11672);
xnor U27272 (N_27272,N_11878,N_11004);
nand U27273 (N_27273,N_18630,N_14790);
xnor U27274 (N_27274,N_10194,N_13307);
and U27275 (N_27275,N_11486,N_10813);
xnor U27276 (N_27276,N_14695,N_10388);
nand U27277 (N_27277,N_11386,N_11331);
nand U27278 (N_27278,N_14729,N_11179);
or U27279 (N_27279,N_15149,N_17299);
and U27280 (N_27280,N_13375,N_13706);
xnor U27281 (N_27281,N_15193,N_19988);
nor U27282 (N_27282,N_16055,N_16862);
and U27283 (N_27283,N_17575,N_13202);
nand U27284 (N_27284,N_15772,N_13239);
xnor U27285 (N_27285,N_19938,N_11617);
and U27286 (N_27286,N_15705,N_17939);
and U27287 (N_27287,N_11859,N_13273);
or U27288 (N_27288,N_10581,N_12929);
nor U27289 (N_27289,N_19751,N_16552);
or U27290 (N_27290,N_14988,N_12310);
nor U27291 (N_27291,N_15110,N_10099);
nor U27292 (N_27292,N_13775,N_10276);
or U27293 (N_27293,N_19420,N_13608);
nand U27294 (N_27294,N_13906,N_11362);
nor U27295 (N_27295,N_16753,N_12427);
nor U27296 (N_27296,N_15722,N_18011);
nand U27297 (N_27297,N_13421,N_11955);
and U27298 (N_27298,N_14442,N_15657);
xnor U27299 (N_27299,N_17306,N_12503);
or U27300 (N_27300,N_12708,N_15780);
nand U27301 (N_27301,N_15132,N_14701);
or U27302 (N_27302,N_15269,N_18239);
nor U27303 (N_27303,N_18245,N_10620);
or U27304 (N_27304,N_12595,N_14498);
nor U27305 (N_27305,N_11314,N_12741);
or U27306 (N_27306,N_17346,N_12565);
xor U27307 (N_27307,N_19913,N_11231);
or U27308 (N_27308,N_13714,N_12408);
xnor U27309 (N_27309,N_14970,N_17463);
xnor U27310 (N_27310,N_17496,N_16564);
nand U27311 (N_27311,N_11873,N_17220);
or U27312 (N_27312,N_19284,N_16388);
or U27313 (N_27313,N_18612,N_15630);
nand U27314 (N_27314,N_10548,N_17377);
nand U27315 (N_27315,N_19256,N_16792);
xnor U27316 (N_27316,N_16228,N_12591);
nor U27317 (N_27317,N_12257,N_13047);
nor U27318 (N_27318,N_13842,N_12260);
or U27319 (N_27319,N_10698,N_14160);
nor U27320 (N_27320,N_18771,N_14584);
or U27321 (N_27321,N_17721,N_17935);
nand U27322 (N_27322,N_15667,N_17711);
and U27323 (N_27323,N_13856,N_14615);
or U27324 (N_27324,N_16367,N_17532);
and U27325 (N_27325,N_12709,N_16114);
nor U27326 (N_27326,N_16071,N_11713);
or U27327 (N_27327,N_10217,N_17892);
nand U27328 (N_27328,N_17324,N_16580);
nor U27329 (N_27329,N_12485,N_15219);
and U27330 (N_27330,N_14959,N_18852);
and U27331 (N_27331,N_18628,N_19217);
or U27332 (N_27332,N_12174,N_19385);
xor U27333 (N_27333,N_17720,N_10954);
nand U27334 (N_27334,N_16382,N_18024);
and U27335 (N_27335,N_19817,N_10135);
or U27336 (N_27336,N_16960,N_13602);
nor U27337 (N_27337,N_15420,N_14367);
nor U27338 (N_27338,N_12934,N_18711);
and U27339 (N_27339,N_11347,N_18628);
and U27340 (N_27340,N_13430,N_15919);
xnor U27341 (N_27341,N_19160,N_19167);
or U27342 (N_27342,N_14811,N_13800);
and U27343 (N_27343,N_16780,N_18288);
and U27344 (N_27344,N_11820,N_15196);
or U27345 (N_27345,N_10341,N_19107);
nand U27346 (N_27346,N_19052,N_18755);
nand U27347 (N_27347,N_13190,N_19275);
or U27348 (N_27348,N_13608,N_10278);
xnor U27349 (N_27349,N_18977,N_18500);
or U27350 (N_27350,N_17526,N_14519);
or U27351 (N_27351,N_17288,N_14955);
nor U27352 (N_27352,N_12301,N_19996);
nor U27353 (N_27353,N_13473,N_14451);
and U27354 (N_27354,N_14563,N_10470);
nand U27355 (N_27355,N_10085,N_17798);
nand U27356 (N_27356,N_10806,N_14036);
or U27357 (N_27357,N_12326,N_14773);
nor U27358 (N_27358,N_10744,N_16447);
or U27359 (N_27359,N_11210,N_12826);
nor U27360 (N_27360,N_14994,N_11620);
nor U27361 (N_27361,N_11064,N_14742);
or U27362 (N_27362,N_18762,N_10270);
or U27363 (N_27363,N_10404,N_12444);
nor U27364 (N_27364,N_17290,N_17918);
nand U27365 (N_27365,N_12866,N_14889);
xnor U27366 (N_27366,N_16070,N_16057);
or U27367 (N_27367,N_10170,N_19765);
or U27368 (N_27368,N_12928,N_13339);
and U27369 (N_27369,N_13643,N_12239);
xor U27370 (N_27370,N_16473,N_13012);
xor U27371 (N_27371,N_11202,N_19368);
nand U27372 (N_27372,N_17227,N_18013);
and U27373 (N_27373,N_12927,N_13079);
or U27374 (N_27374,N_13175,N_12213);
or U27375 (N_27375,N_12478,N_11482);
or U27376 (N_27376,N_10211,N_18251);
xnor U27377 (N_27377,N_13342,N_16157);
xor U27378 (N_27378,N_15454,N_10177);
or U27379 (N_27379,N_11454,N_16538);
xor U27380 (N_27380,N_17092,N_10896);
and U27381 (N_27381,N_13195,N_11959);
nand U27382 (N_27382,N_14772,N_14555);
xnor U27383 (N_27383,N_13369,N_14087);
or U27384 (N_27384,N_11090,N_15231);
xnor U27385 (N_27385,N_10306,N_18117);
or U27386 (N_27386,N_14745,N_15150);
nand U27387 (N_27387,N_15684,N_14286);
nand U27388 (N_27388,N_19433,N_17795);
or U27389 (N_27389,N_10642,N_14974);
and U27390 (N_27390,N_12001,N_10668);
and U27391 (N_27391,N_11892,N_19044);
nor U27392 (N_27392,N_18438,N_11707);
nor U27393 (N_27393,N_16137,N_16784);
nand U27394 (N_27394,N_13193,N_10980);
nor U27395 (N_27395,N_13328,N_16535);
nand U27396 (N_27396,N_19236,N_13453);
nor U27397 (N_27397,N_14154,N_17216);
nand U27398 (N_27398,N_15098,N_12131);
and U27399 (N_27399,N_15791,N_18461);
nand U27400 (N_27400,N_13108,N_19426);
nand U27401 (N_27401,N_18684,N_14249);
nor U27402 (N_27402,N_11803,N_16588);
or U27403 (N_27403,N_14172,N_10007);
nor U27404 (N_27404,N_12883,N_15030);
or U27405 (N_27405,N_14011,N_15315);
nor U27406 (N_27406,N_10398,N_17306);
or U27407 (N_27407,N_19237,N_14083);
nand U27408 (N_27408,N_19918,N_14329);
and U27409 (N_27409,N_12620,N_19278);
xnor U27410 (N_27410,N_10859,N_14217);
and U27411 (N_27411,N_11204,N_15120);
xnor U27412 (N_27412,N_17737,N_18548);
and U27413 (N_27413,N_19473,N_17340);
nor U27414 (N_27414,N_18449,N_10591);
xor U27415 (N_27415,N_11707,N_13187);
or U27416 (N_27416,N_14508,N_11544);
xor U27417 (N_27417,N_10290,N_19195);
and U27418 (N_27418,N_18364,N_18830);
xnor U27419 (N_27419,N_11415,N_14774);
and U27420 (N_27420,N_17936,N_16714);
or U27421 (N_27421,N_17512,N_19601);
nand U27422 (N_27422,N_18701,N_19556);
and U27423 (N_27423,N_12837,N_14503);
nor U27424 (N_27424,N_19194,N_18061);
or U27425 (N_27425,N_16049,N_14101);
and U27426 (N_27426,N_14993,N_13235);
xor U27427 (N_27427,N_15806,N_12669);
nor U27428 (N_27428,N_19647,N_19374);
nor U27429 (N_27429,N_12702,N_19142);
nand U27430 (N_27430,N_14965,N_16456);
xnor U27431 (N_27431,N_11083,N_14835);
and U27432 (N_27432,N_14266,N_12577);
nor U27433 (N_27433,N_16596,N_10862);
or U27434 (N_27434,N_13955,N_10284);
nor U27435 (N_27435,N_15412,N_16190);
nor U27436 (N_27436,N_15393,N_13472);
and U27437 (N_27437,N_17464,N_14936);
nor U27438 (N_27438,N_16518,N_11852);
and U27439 (N_27439,N_19325,N_10964);
xnor U27440 (N_27440,N_19463,N_18136);
nand U27441 (N_27441,N_13504,N_15238);
nor U27442 (N_27442,N_12373,N_12614);
and U27443 (N_27443,N_18386,N_11176);
or U27444 (N_27444,N_18500,N_12064);
or U27445 (N_27445,N_19310,N_18498);
nand U27446 (N_27446,N_18888,N_19236);
nand U27447 (N_27447,N_12382,N_17332);
xnor U27448 (N_27448,N_10665,N_15064);
xnor U27449 (N_27449,N_17642,N_12114);
xor U27450 (N_27450,N_15833,N_13012);
and U27451 (N_27451,N_19644,N_16440);
xor U27452 (N_27452,N_18682,N_11357);
nor U27453 (N_27453,N_12054,N_10596);
nor U27454 (N_27454,N_14823,N_15343);
nor U27455 (N_27455,N_14741,N_17200);
nor U27456 (N_27456,N_13686,N_18269);
and U27457 (N_27457,N_16376,N_15725);
or U27458 (N_27458,N_10833,N_12648);
xor U27459 (N_27459,N_17810,N_17980);
nand U27460 (N_27460,N_18557,N_10813);
or U27461 (N_27461,N_14112,N_10200);
or U27462 (N_27462,N_17178,N_15515);
nor U27463 (N_27463,N_14776,N_18149);
nand U27464 (N_27464,N_16648,N_10726);
xor U27465 (N_27465,N_19226,N_13855);
xor U27466 (N_27466,N_12979,N_13607);
and U27467 (N_27467,N_13069,N_17322);
or U27468 (N_27468,N_13068,N_17704);
nor U27469 (N_27469,N_16600,N_12587);
nand U27470 (N_27470,N_19974,N_16970);
nand U27471 (N_27471,N_13414,N_15489);
or U27472 (N_27472,N_10053,N_12571);
and U27473 (N_27473,N_16675,N_14807);
xnor U27474 (N_27474,N_14196,N_15138);
nand U27475 (N_27475,N_18705,N_10664);
or U27476 (N_27476,N_15186,N_16365);
or U27477 (N_27477,N_11831,N_14002);
and U27478 (N_27478,N_10476,N_14745);
or U27479 (N_27479,N_15937,N_16790);
nand U27480 (N_27480,N_19997,N_15102);
nor U27481 (N_27481,N_13915,N_11755);
or U27482 (N_27482,N_10178,N_14087);
nand U27483 (N_27483,N_13030,N_12730);
or U27484 (N_27484,N_14452,N_17577);
or U27485 (N_27485,N_10667,N_15596);
and U27486 (N_27486,N_12441,N_11864);
nand U27487 (N_27487,N_14866,N_17938);
nor U27488 (N_27488,N_10712,N_14250);
nor U27489 (N_27489,N_12703,N_17794);
nor U27490 (N_27490,N_12333,N_12032);
nand U27491 (N_27491,N_16786,N_16174);
or U27492 (N_27492,N_10060,N_16686);
nor U27493 (N_27493,N_15940,N_17240);
nor U27494 (N_27494,N_10617,N_14630);
and U27495 (N_27495,N_18483,N_14410);
nand U27496 (N_27496,N_15213,N_15066);
nor U27497 (N_27497,N_15152,N_10912);
and U27498 (N_27498,N_19162,N_17801);
nand U27499 (N_27499,N_17697,N_16790);
nor U27500 (N_27500,N_13386,N_19237);
or U27501 (N_27501,N_14242,N_15747);
or U27502 (N_27502,N_10492,N_15600);
or U27503 (N_27503,N_12658,N_13304);
and U27504 (N_27504,N_18715,N_15820);
nand U27505 (N_27505,N_11017,N_12851);
nor U27506 (N_27506,N_12236,N_11298);
or U27507 (N_27507,N_12351,N_14328);
nor U27508 (N_27508,N_14079,N_13695);
nand U27509 (N_27509,N_19769,N_12202);
or U27510 (N_27510,N_14954,N_12495);
xor U27511 (N_27511,N_19226,N_14253);
xnor U27512 (N_27512,N_12613,N_17927);
xnor U27513 (N_27513,N_12518,N_19450);
nand U27514 (N_27514,N_17625,N_13381);
xnor U27515 (N_27515,N_14852,N_15912);
nand U27516 (N_27516,N_18928,N_13222);
or U27517 (N_27517,N_12885,N_12048);
nand U27518 (N_27518,N_12003,N_11547);
nor U27519 (N_27519,N_17926,N_11163);
xor U27520 (N_27520,N_19166,N_14931);
or U27521 (N_27521,N_13248,N_12132);
xnor U27522 (N_27522,N_15208,N_12649);
and U27523 (N_27523,N_19608,N_18143);
nor U27524 (N_27524,N_12857,N_10284);
and U27525 (N_27525,N_15287,N_12578);
and U27526 (N_27526,N_16467,N_14869);
nand U27527 (N_27527,N_11524,N_14467);
nand U27528 (N_27528,N_11054,N_11765);
and U27529 (N_27529,N_10937,N_11959);
or U27530 (N_27530,N_19937,N_13351);
xnor U27531 (N_27531,N_15653,N_18898);
nor U27532 (N_27532,N_18971,N_10814);
xor U27533 (N_27533,N_15268,N_19583);
or U27534 (N_27534,N_15219,N_11625);
nor U27535 (N_27535,N_11721,N_14103);
and U27536 (N_27536,N_19214,N_16962);
nor U27537 (N_27537,N_17632,N_17706);
nor U27538 (N_27538,N_10477,N_18584);
nor U27539 (N_27539,N_17428,N_19336);
nor U27540 (N_27540,N_19917,N_19368);
nand U27541 (N_27541,N_18370,N_14363);
nor U27542 (N_27542,N_15442,N_18290);
nor U27543 (N_27543,N_11171,N_15732);
xnor U27544 (N_27544,N_10527,N_15726);
nor U27545 (N_27545,N_17536,N_14259);
nor U27546 (N_27546,N_10774,N_18095);
xor U27547 (N_27547,N_10870,N_14028);
nand U27548 (N_27548,N_10063,N_17455);
and U27549 (N_27549,N_13859,N_11790);
xor U27550 (N_27550,N_17262,N_13398);
nor U27551 (N_27551,N_13824,N_17547);
and U27552 (N_27552,N_12618,N_13158);
nor U27553 (N_27553,N_10483,N_11253);
xnor U27554 (N_27554,N_15080,N_12478);
nor U27555 (N_27555,N_19022,N_19751);
nand U27556 (N_27556,N_14250,N_18067);
or U27557 (N_27557,N_11307,N_17898);
nand U27558 (N_27558,N_19598,N_14779);
nand U27559 (N_27559,N_16806,N_12631);
xor U27560 (N_27560,N_19407,N_15071);
xor U27561 (N_27561,N_19021,N_17250);
nand U27562 (N_27562,N_11222,N_10844);
and U27563 (N_27563,N_10406,N_10637);
or U27564 (N_27564,N_14971,N_16567);
xor U27565 (N_27565,N_13397,N_16193);
or U27566 (N_27566,N_19075,N_19770);
nand U27567 (N_27567,N_12638,N_11367);
or U27568 (N_27568,N_10687,N_14769);
and U27569 (N_27569,N_14615,N_12118);
nor U27570 (N_27570,N_19366,N_19535);
and U27571 (N_27571,N_13119,N_16111);
xnor U27572 (N_27572,N_15193,N_12259);
and U27573 (N_27573,N_11638,N_19002);
xor U27574 (N_27574,N_15156,N_13484);
or U27575 (N_27575,N_17512,N_18150);
and U27576 (N_27576,N_15149,N_14482);
xnor U27577 (N_27577,N_16893,N_16929);
nor U27578 (N_27578,N_10212,N_18950);
and U27579 (N_27579,N_12042,N_11844);
nand U27580 (N_27580,N_14315,N_12947);
nand U27581 (N_27581,N_16510,N_12791);
xnor U27582 (N_27582,N_14532,N_10433);
nand U27583 (N_27583,N_10358,N_10407);
nand U27584 (N_27584,N_14495,N_18519);
nand U27585 (N_27585,N_18748,N_19049);
xnor U27586 (N_27586,N_17035,N_12515);
or U27587 (N_27587,N_12818,N_15345);
nand U27588 (N_27588,N_16039,N_13115);
nor U27589 (N_27589,N_13294,N_11164);
and U27590 (N_27590,N_16975,N_13676);
xor U27591 (N_27591,N_13404,N_13893);
nor U27592 (N_27592,N_17274,N_13344);
xor U27593 (N_27593,N_12107,N_12930);
xor U27594 (N_27594,N_17708,N_19539);
xor U27595 (N_27595,N_18887,N_13216);
nor U27596 (N_27596,N_10858,N_10799);
and U27597 (N_27597,N_11833,N_14209);
xor U27598 (N_27598,N_16241,N_15259);
xnor U27599 (N_27599,N_12217,N_17559);
nand U27600 (N_27600,N_17041,N_10387);
nand U27601 (N_27601,N_12990,N_17421);
nand U27602 (N_27602,N_10656,N_12818);
or U27603 (N_27603,N_17756,N_13725);
and U27604 (N_27604,N_13205,N_19603);
and U27605 (N_27605,N_13460,N_19840);
xnor U27606 (N_27606,N_11858,N_16022);
xor U27607 (N_27607,N_14797,N_18143);
and U27608 (N_27608,N_17544,N_13304);
nor U27609 (N_27609,N_10764,N_18423);
xor U27610 (N_27610,N_16085,N_17348);
nor U27611 (N_27611,N_15022,N_18524);
nor U27612 (N_27612,N_17482,N_16907);
xor U27613 (N_27613,N_15336,N_13435);
nand U27614 (N_27614,N_13208,N_14492);
nor U27615 (N_27615,N_10408,N_18470);
and U27616 (N_27616,N_11026,N_15221);
or U27617 (N_27617,N_15543,N_16551);
xor U27618 (N_27618,N_16371,N_19750);
nor U27619 (N_27619,N_10029,N_12240);
nor U27620 (N_27620,N_11511,N_10716);
xor U27621 (N_27621,N_15481,N_11423);
nor U27622 (N_27622,N_17103,N_10759);
nor U27623 (N_27623,N_17923,N_12973);
nor U27624 (N_27624,N_18695,N_14552);
nand U27625 (N_27625,N_17345,N_19173);
nand U27626 (N_27626,N_12405,N_18576);
xor U27627 (N_27627,N_12126,N_17702);
or U27628 (N_27628,N_16101,N_16113);
xnor U27629 (N_27629,N_13482,N_18468);
xor U27630 (N_27630,N_10124,N_18095);
or U27631 (N_27631,N_17818,N_19545);
and U27632 (N_27632,N_18242,N_10838);
or U27633 (N_27633,N_10939,N_12329);
nand U27634 (N_27634,N_17920,N_11730);
nor U27635 (N_27635,N_14401,N_18761);
nand U27636 (N_27636,N_14301,N_15780);
and U27637 (N_27637,N_14689,N_13647);
nor U27638 (N_27638,N_14934,N_15057);
nor U27639 (N_27639,N_10129,N_12130);
or U27640 (N_27640,N_14959,N_11927);
and U27641 (N_27641,N_13023,N_17880);
or U27642 (N_27642,N_10391,N_17467);
and U27643 (N_27643,N_17699,N_19129);
or U27644 (N_27644,N_10967,N_10495);
or U27645 (N_27645,N_17844,N_19088);
nor U27646 (N_27646,N_14883,N_17431);
or U27647 (N_27647,N_17481,N_11655);
or U27648 (N_27648,N_13234,N_14177);
nand U27649 (N_27649,N_18051,N_18142);
xor U27650 (N_27650,N_12728,N_14815);
xor U27651 (N_27651,N_15984,N_10330);
and U27652 (N_27652,N_17644,N_13613);
nor U27653 (N_27653,N_10462,N_13184);
and U27654 (N_27654,N_13463,N_17615);
xor U27655 (N_27655,N_14872,N_10647);
nor U27656 (N_27656,N_10334,N_16523);
nor U27657 (N_27657,N_19658,N_16251);
or U27658 (N_27658,N_19296,N_18672);
or U27659 (N_27659,N_14503,N_11710);
nand U27660 (N_27660,N_16278,N_15937);
and U27661 (N_27661,N_11111,N_14371);
xnor U27662 (N_27662,N_16133,N_13987);
and U27663 (N_27663,N_12147,N_13306);
and U27664 (N_27664,N_14040,N_18956);
nor U27665 (N_27665,N_15733,N_19233);
nand U27666 (N_27666,N_15484,N_16930);
and U27667 (N_27667,N_17354,N_12885);
or U27668 (N_27668,N_14555,N_16576);
and U27669 (N_27669,N_17875,N_14030);
xor U27670 (N_27670,N_17652,N_16133);
and U27671 (N_27671,N_11102,N_13627);
nor U27672 (N_27672,N_10524,N_16532);
or U27673 (N_27673,N_13720,N_19814);
and U27674 (N_27674,N_15296,N_19894);
xnor U27675 (N_27675,N_12030,N_10360);
nor U27676 (N_27676,N_12442,N_10533);
nor U27677 (N_27677,N_11702,N_12325);
or U27678 (N_27678,N_17403,N_17128);
and U27679 (N_27679,N_13538,N_12269);
nor U27680 (N_27680,N_14263,N_13365);
nor U27681 (N_27681,N_12132,N_10207);
nand U27682 (N_27682,N_12899,N_15408);
nor U27683 (N_27683,N_10619,N_10757);
and U27684 (N_27684,N_19638,N_12405);
nor U27685 (N_27685,N_14543,N_10077);
nor U27686 (N_27686,N_14752,N_13092);
xor U27687 (N_27687,N_12569,N_17825);
xor U27688 (N_27688,N_11801,N_14292);
and U27689 (N_27689,N_11219,N_19942);
or U27690 (N_27690,N_18550,N_15549);
nand U27691 (N_27691,N_12621,N_12857);
nor U27692 (N_27692,N_10364,N_11349);
xor U27693 (N_27693,N_17353,N_19530);
nand U27694 (N_27694,N_10474,N_16974);
and U27695 (N_27695,N_12365,N_11554);
xor U27696 (N_27696,N_13123,N_13082);
xor U27697 (N_27697,N_19975,N_13203);
nor U27698 (N_27698,N_12292,N_11925);
nand U27699 (N_27699,N_14303,N_19304);
nor U27700 (N_27700,N_11519,N_19953);
nor U27701 (N_27701,N_18486,N_10213);
and U27702 (N_27702,N_11967,N_14349);
xor U27703 (N_27703,N_10478,N_15568);
nand U27704 (N_27704,N_17996,N_12032);
nand U27705 (N_27705,N_13066,N_19376);
nor U27706 (N_27706,N_19622,N_19953);
nand U27707 (N_27707,N_18465,N_17459);
xnor U27708 (N_27708,N_13618,N_16560);
nand U27709 (N_27709,N_15351,N_13571);
or U27710 (N_27710,N_17307,N_18139);
nand U27711 (N_27711,N_11287,N_18280);
nor U27712 (N_27712,N_13793,N_14850);
nor U27713 (N_27713,N_14965,N_15373);
xor U27714 (N_27714,N_10655,N_13208);
or U27715 (N_27715,N_14900,N_11235);
nor U27716 (N_27716,N_13338,N_19584);
or U27717 (N_27717,N_19751,N_17829);
nor U27718 (N_27718,N_15448,N_12532);
nor U27719 (N_27719,N_12041,N_19190);
nor U27720 (N_27720,N_16672,N_13711);
xor U27721 (N_27721,N_10356,N_15928);
and U27722 (N_27722,N_18602,N_12079);
xnor U27723 (N_27723,N_16848,N_10519);
nor U27724 (N_27724,N_17949,N_16019);
or U27725 (N_27725,N_11415,N_17063);
nand U27726 (N_27726,N_12251,N_12086);
nor U27727 (N_27727,N_10237,N_11567);
or U27728 (N_27728,N_10761,N_19328);
or U27729 (N_27729,N_16511,N_12360);
nor U27730 (N_27730,N_11202,N_17574);
nand U27731 (N_27731,N_14545,N_11522);
xnor U27732 (N_27732,N_17920,N_18855);
nand U27733 (N_27733,N_13358,N_15715);
or U27734 (N_27734,N_10994,N_14866);
and U27735 (N_27735,N_14838,N_14842);
xnor U27736 (N_27736,N_15561,N_17244);
nand U27737 (N_27737,N_14730,N_10976);
or U27738 (N_27738,N_10325,N_19893);
xor U27739 (N_27739,N_11082,N_14476);
xor U27740 (N_27740,N_14540,N_12011);
or U27741 (N_27741,N_14605,N_10085);
or U27742 (N_27742,N_15651,N_17281);
or U27743 (N_27743,N_11057,N_11130);
nand U27744 (N_27744,N_14847,N_19483);
nand U27745 (N_27745,N_14160,N_14035);
xnor U27746 (N_27746,N_16627,N_15494);
and U27747 (N_27747,N_14017,N_17213);
and U27748 (N_27748,N_14689,N_11506);
nor U27749 (N_27749,N_14457,N_18440);
nand U27750 (N_27750,N_12804,N_19749);
nand U27751 (N_27751,N_10024,N_16585);
xnor U27752 (N_27752,N_15012,N_11790);
nor U27753 (N_27753,N_16408,N_15893);
nor U27754 (N_27754,N_14781,N_12193);
and U27755 (N_27755,N_15999,N_11425);
and U27756 (N_27756,N_14279,N_18810);
and U27757 (N_27757,N_16387,N_11993);
and U27758 (N_27758,N_13985,N_12147);
nand U27759 (N_27759,N_11545,N_18452);
xor U27760 (N_27760,N_10434,N_15903);
nand U27761 (N_27761,N_12069,N_18105);
nand U27762 (N_27762,N_11998,N_13571);
nor U27763 (N_27763,N_10841,N_11542);
or U27764 (N_27764,N_17096,N_11075);
nor U27765 (N_27765,N_15148,N_19094);
or U27766 (N_27766,N_16294,N_11463);
xor U27767 (N_27767,N_17615,N_15658);
or U27768 (N_27768,N_15134,N_19052);
nor U27769 (N_27769,N_15086,N_16506);
or U27770 (N_27770,N_16678,N_16774);
nor U27771 (N_27771,N_16870,N_17884);
and U27772 (N_27772,N_14062,N_19050);
or U27773 (N_27773,N_18187,N_15661);
and U27774 (N_27774,N_18240,N_13467);
xnor U27775 (N_27775,N_19859,N_18942);
or U27776 (N_27776,N_17055,N_13864);
nor U27777 (N_27777,N_11845,N_14063);
and U27778 (N_27778,N_15206,N_10502);
and U27779 (N_27779,N_11160,N_11449);
and U27780 (N_27780,N_11412,N_16209);
or U27781 (N_27781,N_10384,N_17874);
xnor U27782 (N_27782,N_19264,N_13883);
or U27783 (N_27783,N_11142,N_10236);
or U27784 (N_27784,N_16976,N_16444);
and U27785 (N_27785,N_18358,N_13331);
xor U27786 (N_27786,N_19255,N_11904);
xnor U27787 (N_27787,N_10749,N_11701);
nor U27788 (N_27788,N_18640,N_16900);
or U27789 (N_27789,N_11872,N_14181);
and U27790 (N_27790,N_16455,N_10137);
nor U27791 (N_27791,N_18739,N_16614);
and U27792 (N_27792,N_18014,N_13850);
nand U27793 (N_27793,N_10854,N_19714);
nor U27794 (N_27794,N_19370,N_14371);
nand U27795 (N_27795,N_17686,N_17010);
or U27796 (N_27796,N_12592,N_10216);
nor U27797 (N_27797,N_16994,N_14807);
nand U27798 (N_27798,N_19825,N_10952);
nand U27799 (N_27799,N_11182,N_10533);
nor U27800 (N_27800,N_18395,N_16004);
and U27801 (N_27801,N_15860,N_14777);
nand U27802 (N_27802,N_18685,N_18083);
xor U27803 (N_27803,N_17832,N_15332);
and U27804 (N_27804,N_14092,N_15048);
or U27805 (N_27805,N_15010,N_16881);
xor U27806 (N_27806,N_17232,N_15372);
and U27807 (N_27807,N_14654,N_15616);
and U27808 (N_27808,N_15884,N_10725);
and U27809 (N_27809,N_12727,N_12182);
nor U27810 (N_27810,N_13889,N_17409);
xnor U27811 (N_27811,N_18984,N_14885);
xor U27812 (N_27812,N_19731,N_11605);
nand U27813 (N_27813,N_19124,N_13089);
and U27814 (N_27814,N_13368,N_11065);
nand U27815 (N_27815,N_10500,N_19322);
nand U27816 (N_27816,N_17100,N_18631);
and U27817 (N_27817,N_18831,N_19525);
or U27818 (N_27818,N_16405,N_14177);
and U27819 (N_27819,N_15676,N_16160);
nor U27820 (N_27820,N_12044,N_18880);
or U27821 (N_27821,N_18348,N_18490);
nor U27822 (N_27822,N_18519,N_19416);
nand U27823 (N_27823,N_10268,N_10940);
nor U27824 (N_27824,N_16836,N_11395);
nand U27825 (N_27825,N_11804,N_14378);
or U27826 (N_27826,N_13157,N_10045);
xor U27827 (N_27827,N_19436,N_15800);
or U27828 (N_27828,N_16329,N_11858);
and U27829 (N_27829,N_15998,N_18183);
or U27830 (N_27830,N_16314,N_12626);
and U27831 (N_27831,N_14138,N_17541);
xor U27832 (N_27832,N_17619,N_13533);
xor U27833 (N_27833,N_17865,N_15399);
nand U27834 (N_27834,N_19560,N_12467);
or U27835 (N_27835,N_14512,N_15569);
xor U27836 (N_27836,N_14023,N_14566);
and U27837 (N_27837,N_19728,N_13370);
xor U27838 (N_27838,N_14018,N_13049);
nor U27839 (N_27839,N_13480,N_19805);
or U27840 (N_27840,N_12891,N_11701);
nor U27841 (N_27841,N_16755,N_13495);
nand U27842 (N_27842,N_10840,N_17678);
nor U27843 (N_27843,N_17700,N_10015);
nand U27844 (N_27844,N_18645,N_11586);
nor U27845 (N_27845,N_11475,N_18496);
nand U27846 (N_27846,N_18742,N_18292);
and U27847 (N_27847,N_15233,N_13604);
or U27848 (N_27848,N_12743,N_19784);
xnor U27849 (N_27849,N_15394,N_19869);
nor U27850 (N_27850,N_10826,N_19050);
nand U27851 (N_27851,N_18069,N_19859);
xor U27852 (N_27852,N_18098,N_17022);
nand U27853 (N_27853,N_12090,N_17302);
nor U27854 (N_27854,N_14045,N_17957);
and U27855 (N_27855,N_10633,N_13360);
nand U27856 (N_27856,N_17653,N_19816);
and U27857 (N_27857,N_10307,N_12584);
nand U27858 (N_27858,N_19814,N_17907);
and U27859 (N_27859,N_12604,N_15185);
and U27860 (N_27860,N_17904,N_16600);
xor U27861 (N_27861,N_10709,N_15536);
or U27862 (N_27862,N_12742,N_15946);
xor U27863 (N_27863,N_14193,N_12455);
xor U27864 (N_27864,N_19242,N_19205);
xnor U27865 (N_27865,N_17011,N_18541);
nor U27866 (N_27866,N_15160,N_15032);
nand U27867 (N_27867,N_10206,N_14639);
and U27868 (N_27868,N_15314,N_12255);
or U27869 (N_27869,N_12695,N_14892);
nand U27870 (N_27870,N_13551,N_11356);
or U27871 (N_27871,N_17116,N_11812);
nand U27872 (N_27872,N_19273,N_12262);
and U27873 (N_27873,N_16480,N_16761);
and U27874 (N_27874,N_16701,N_19451);
nor U27875 (N_27875,N_15693,N_12127);
and U27876 (N_27876,N_14319,N_15753);
nand U27877 (N_27877,N_15091,N_12950);
nor U27878 (N_27878,N_18734,N_16518);
nor U27879 (N_27879,N_16287,N_19668);
nand U27880 (N_27880,N_17274,N_17663);
or U27881 (N_27881,N_16979,N_18113);
or U27882 (N_27882,N_17317,N_17852);
nand U27883 (N_27883,N_19721,N_15414);
and U27884 (N_27884,N_13854,N_15959);
or U27885 (N_27885,N_15715,N_16584);
and U27886 (N_27886,N_18134,N_14362);
nor U27887 (N_27887,N_18596,N_15276);
nor U27888 (N_27888,N_16707,N_19674);
or U27889 (N_27889,N_17099,N_19263);
or U27890 (N_27890,N_12895,N_18892);
and U27891 (N_27891,N_12357,N_14170);
nand U27892 (N_27892,N_18718,N_19293);
xor U27893 (N_27893,N_14836,N_19201);
and U27894 (N_27894,N_12507,N_15885);
xor U27895 (N_27895,N_10103,N_10350);
xor U27896 (N_27896,N_12910,N_18259);
or U27897 (N_27897,N_15715,N_12381);
xor U27898 (N_27898,N_16129,N_14772);
or U27899 (N_27899,N_17197,N_13402);
nand U27900 (N_27900,N_14678,N_10304);
nor U27901 (N_27901,N_14623,N_14432);
and U27902 (N_27902,N_12707,N_11192);
and U27903 (N_27903,N_13361,N_15868);
nand U27904 (N_27904,N_10723,N_16769);
xnor U27905 (N_27905,N_18229,N_10416);
nand U27906 (N_27906,N_15074,N_17516);
and U27907 (N_27907,N_11879,N_17780);
and U27908 (N_27908,N_19726,N_15809);
xnor U27909 (N_27909,N_17028,N_10787);
nand U27910 (N_27910,N_13859,N_10165);
nor U27911 (N_27911,N_11310,N_11077);
nand U27912 (N_27912,N_14854,N_19350);
xnor U27913 (N_27913,N_19645,N_19440);
nor U27914 (N_27914,N_13906,N_12505);
or U27915 (N_27915,N_13226,N_16176);
and U27916 (N_27916,N_19106,N_17358);
nor U27917 (N_27917,N_10588,N_19863);
nor U27918 (N_27918,N_10004,N_14786);
nor U27919 (N_27919,N_19931,N_14946);
and U27920 (N_27920,N_14692,N_19406);
nand U27921 (N_27921,N_15450,N_19105);
and U27922 (N_27922,N_19002,N_16072);
nor U27923 (N_27923,N_14042,N_13724);
or U27924 (N_27924,N_16305,N_16463);
and U27925 (N_27925,N_14577,N_10021);
and U27926 (N_27926,N_12881,N_15923);
and U27927 (N_27927,N_19251,N_18895);
or U27928 (N_27928,N_17813,N_17625);
xnor U27929 (N_27929,N_11340,N_13427);
or U27930 (N_27930,N_11744,N_11851);
nor U27931 (N_27931,N_16687,N_16396);
nand U27932 (N_27932,N_19134,N_14432);
nor U27933 (N_27933,N_17053,N_19969);
and U27934 (N_27934,N_16110,N_12481);
nor U27935 (N_27935,N_18981,N_12254);
xor U27936 (N_27936,N_19399,N_12678);
nand U27937 (N_27937,N_19097,N_15482);
nor U27938 (N_27938,N_19451,N_11307);
nand U27939 (N_27939,N_19023,N_13115);
nor U27940 (N_27940,N_19861,N_13225);
xor U27941 (N_27941,N_13315,N_18525);
xor U27942 (N_27942,N_15517,N_18996);
nor U27943 (N_27943,N_10868,N_10821);
or U27944 (N_27944,N_12287,N_14794);
xor U27945 (N_27945,N_11224,N_11028);
xnor U27946 (N_27946,N_15644,N_12432);
nor U27947 (N_27947,N_10313,N_18112);
nor U27948 (N_27948,N_13959,N_17920);
nand U27949 (N_27949,N_18587,N_12749);
xnor U27950 (N_27950,N_13237,N_14278);
nand U27951 (N_27951,N_18792,N_18659);
and U27952 (N_27952,N_18648,N_14846);
xor U27953 (N_27953,N_16483,N_13913);
xor U27954 (N_27954,N_11489,N_16304);
nor U27955 (N_27955,N_14830,N_14306);
xor U27956 (N_27956,N_18116,N_12255);
nand U27957 (N_27957,N_15013,N_14991);
or U27958 (N_27958,N_18052,N_12621);
nand U27959 (N_27959,N_11421,N_12558);
xor U27960 (N_27960,N_11990,N_11608);
nand U27961 (N_27961,N_15109,N_18468);
or U27962 (N_27962,N_12456,N_18485);
and U27963 (N_27963,N_12576,N_18995);
nor U27964 (N_27964,N_15358,N_13130);
or U27965 (N_27965,N_11492,N_11088);
or U27966 (N_27966,N_17835,N_18624);
or U27967 (N_27967,N_13225,N_10603);
or U27968 (N_27968,N_10932,N_16900);
nor U27969 (N_27969,N_16059,N_19349);
and U27970 (N_27970,N_11570,N_18489);
or U27971 (N_27971,N_19966,N_13115);
xor U27972 (N_27972,N_13687,N_16436);
nand U27973 (N_27973,N_18108,N_19763);
nand U27974 (N_27974,N_19036,N_16169);
or U27975 (N_27975,N_17978,N_14690);
xor U27976 (N_27976,N_19580,N_13985);
xor U27977 (N_27977,N_19282,N_16519);
nor U27978 (N_27978,N_18428,N_19838);
and U27979 (N_27979,N_15041,N_10161);
or U27980 (N_27980,N_11165,N_14518);
or U27981 (N_27981,N_17448,N_13191);
nand U27982 (N_27982,N_17301,N_18866);
nor U27983 (N_27983,N_10863,N_17345);
xnor U27984 (N_27984,N_12250,N_19247);
nor U27985 (N_27985,N_15640,N_15629);
and U27986 (N_27986,N_11261,N_15500);
or U27987 (N_27987,N_14004,N_12273);
xnor U27988 (N_27988,N_12911,N_10397);
xnor U27989 (N_27989,N_11219,N_13774);
or U27990 (N_27990,N_13327,N_18406);
and U27991 (N_27991,N_15600,N_14317);
nor U27992 (N_27992,N_19373,N_10394);
or U27993 (N_27993,N_17326,N_11412);
or U27994 (N_27994,N_11466,N_18306);
xnor U27995 (N_27995,N_11505,N_19801);
xor U27996 (N_27996,N_18076,N_12366);
xnor U27997 (N_27997,N_19314,N_12792);
xor U27998 (N_27998,N_12891,N_19510);
or U27999 (N_27999,N_13406,N_11737);
nand U28000 (N_28000,N_18273,N_17080);
nor U28001 (N_28001,N_12864,N_17932);
or U28002 (N_28002,N_15389,N_18521);
nor U28003 (N_28003,N_14776,N_12485);
nand U28004 (N_28004,N_13604,N_14476);
or U28005 (N_28005,N_16426,N_13657);
nand U28006 (N_28006,N_15773,N_19711);
and U28007 (N_28007,N_14754,N_19857);
nor U28008 (N_28008,N_14724,N_17456);
and U28009 (N_28009,N_12545,N_11492);
or U28010 (N_28010,N_11564,N_13573);
or U28011 (N_28011,N_17650,N_12229);
and U28012 (N_28012,N_16760,N_15719);
nand U28013 (N_28013,N_16307,N_15392);
and U28014 (N_28014,N_13716,N_17621);
or U28015 (N_28015,N_17261,N_18686);
or U28016 (N_28016,N_15234,N_18376);
or U28017 (N_28017,N_11349,N_12161);
nand U28018 (N_28018,N_13964,N_13410);
or U28019 (N_28019,N_14774,N_11653);
or U28020 (N_28020,N_19336,N_15968);
or U28021 (N_28021,N_11545,N_17013);
xor U28022 (N_28022,N_10406,N_14627);
and U28023 (N_28023,N_10036,N_11517);
nor U28024 (N_28024,N_14348,N_11177);
xnor U28025 (N_28025,N_18074,N_16428);
nor U28026 (N_28026,N_14850,N_17452);
or U28027 (N_28027,N_11619,N_14354);
nor U28028 (N_28028,N_18201,N_18278);
and U28029 (N_28029,N_16214,N_14988);
or U28030 (N_28030,N_19379,N_17994);
or U28031 (N_28031,N_12694,N_12425);
and U28032 (N_28032,N_19688,N_17051);
nand U28033 (N_28033,N_13220,N_13520);
xor U28034 (N_28034,N_10464,N_17864);
nand U28035 (N_28035,N_15190,N_18623);
nor U28036 (N_28036,N_14125,N_15768);
nand U28037 (N_28037,N_15926,N_15886);
xor U28038 (N_28038,N_15097,N_13937);
nor U28039 (N_28039,N_10718,N_14408);
and U28040 (N_28040,N_10342,N_10556);
or U28041 (N_28041,N_13690,N_12700);
nor U28042 (N_28042,N_17441,N_15175);
xnor U28043 (N_28043,N_16943,N_11403);
or U28044 (N_28044,N_18504,N_12119);
nand U28045 (N_28045,N_19710,N_15020);
or U28046 (N_28046,N_12483,N_15910);
or U28047 (N_28047,N_14185,N_17192);
and U28048 (N_28048,N_12662,N_12334);
or U28049 (N_28049,N_12740,N_15380);
nand U28050 (N_28050,N_19803,N_16031);
nand U28051 (N_28051,N_10983,N_17849);
and U28052 (N_28052,N_18937,N_10215);
and U28053 (N_28053,N_13812,N_19777);
nand U28054 (N_28054,N_13863,N_16743);
nor U28055 (N_28055,N_12090,N_19849);
nor U28056 (N_28056,N_17023,N_19434);
nand U28057 (N_28057,N_12915,N_19566);
nand U28058 (N_28058,N_14562,N_14008);
nor U28059 (N_28059,N_15988,N_19581);
and U28060 (N_28060,N_10463,N_12794);
xnor U28061 (N_28061,N_17278,N_10425);
xnor U28062 (N_28062,N_17401,N_16392);
xnor U28063 (N_28063,N_16676,N_11108);
and U28064 (N_28064,N_17898,N_17420);
and U28065 (N_28065,N_18460,N_11765);
or U28066 (N_28066,N_16631,N_12621);
or U28067 (N_28067,N_11786,N_19980);
nor U28068 (N_28068,N_14152,N_12144);
nand U28069 (N_28069,N_18866,N_12991);
xor U28070 (N_28070,N_11506,N_17450);
and U28071 (N_28071,N_12065,N_17466);
nor U28072 (N_28072,N_15726,N_18576);
nor U28073 (N_28073,N_17706,N_18833);
and U28074 (N_28074,N_12271,N_18266);
xnor U28075 (N_28075,N_14401,N_18061);
or U28076 (N_28076,N_18243,N_16739);
nor U28077 (N_28077,N_12456,N_16265);
nor U28078 (N_28078,N_12567,N_13772);
xnor U28079 (N_28079,N_14699,N_13554);
xor U28080 (N_28080,N_10856,N_12881);
nand U28081 (N_28081,N_11995,N_12672);
xnor U28082 (N_28082,N_10920,N_17642);
and U28083 (N_28083,N_18664,N_13197);
nand U28084 (N_28084,N_12675,N_18516);
nand U28085 (N_28085,N_17504,N_15323);
xnor U28086 (N_28086,N_13498,N_18478);
nor U28087 (N_28087,N_19963,N_16746);
xnor U28088 (N_28088,N_15670,N_11642);
nor U28089 (N_28089,N_17049,N_15769);
and U28090 (N_28090,N_13523,N_15208);
xnor U28091 (N_28091,N_18134,N_16807);
nand U28092 (N_28092,N_14930,N_18629);
or U28093 (N_28093,N_18298,N_16012);
and U28094 (N_28094,N_12626,N_11246);
nor U28095 (N_28095,N_17955,N_17986);
nor U28096 (N_28096,N_15797,N_10862);
and U28097 (N_28097,N_14938,N_15273);
xor U28098 (N_28098,N_12232,N_11579);
nand U28099 (N_28099,N_18011,N_11954);
xor U28100 (N_28100,N_17803,N_11177);
xnor U28101 (N_28101,N_10224,N_12346);
or U28102 (N_28102,N_17473,N_17622);
or U28103 (N_28103,N_19616,N_13206);
or U28104 (N_28104,N_14725,N_18651);
xor U28105 (N_28105,N_17289,N_17146);
or U28106 (N_28106,N_18027,N_16471);
xnor U28107 (N_28107,N_14956,N_13972);
or U28108 (N_28108,N_18686,N_11545);
nor U28109 (N_28109,N_14359,N_13323);
or U28110 (N_28110,N_10636,N_12860);
nor U28111 (N_28111,N_14397,N_17849);
or U28112 (N_28112,N_10268,N_12233);
xnor U28113 (N_28113,N_12408,N_12637);
and U28114 (N_28114,N_10802,N_15335);
xor U28115 (N_28115,N_16567,N_18482);
nand U28116 (N_28116,N_17192,N_17468);
nand U28117 (N_28117,N_19409,N_19439);
nor U28118 (N_28118,N_13870,N_14011);
nand U28119 (N_28119,N_12298,N_17265);
and U28120 (N_28120,N_13493,N_18264);
or U28121 (N_28121,N_15943,N_15601);
and U28122 (N_28122,N_15006,N_13827);
and U28123 (N_28123,N_16261,N_13240);
and U28124 (N_28124,N_15347,N_11790);
nand U28125 (N_28125,N_12808,N_17159);
nand U28126 (N_28126,N_10109,N_19440);
nor U28127 (N_28127,N_18513,N_12372);
nand U28128 (N_28128,N_18677,N_15964);
and U28129 (N_28129,N_17523,N_16842);
xor U28130 (N_28130,N_12670,N_15724);
and U28131 (N_28131,N_15877,N_10760);
or U28132 (N_28132,N_17795,N_10487);
and U28133 (N_28133,N_10148,N_11952);
or U28134 (N_28134,N_17498,N_13275);
or U28135 (N_28135,N_16112,N_19754);
xor U28136 (N_28136,N_12671,N_11767);
and U28137 (N_28137,N_19399,N_16397);
and U28138 (N_28138,N_19460,N_10774);
or U28139 (N_28139,N_16181,N_13403);
nand U28140 (N_28140,N_17361,N_17337);
xnor U28141 (N_28141,N_13366,N_16939);
and U28142 (N_28142,N_19372,N_12208);
nor U28143 (N_28143,N_15971,N_14839);
xor U28144 (N_28144,N_15512,N_15588);
and U28145 (N_28145,N_13724,N_16692);
nor U28146 (N_28146,N_11142,N_15913);
nand U28147 (N_28147,N_14854,N_11248);
and U28148 (N_28148,N_15939,N_14326);
and U28149 (N_28149,N_11240,N_11887);
nor U28150 (N_28150,N_19024,N_16723);
xor U28151 (N_28151,N_14135,N_10000);
nand U28152 (N_28152,N_15837,N_18407);
nor U28153 (N_28153,N_16386,N_13366);
xnor U28154 (N_28154,N_10931,N_15385);
or U28155 (N_28155,N_13669,N_18425);
xor U28156 (N_28156,N_14572,N_18225);
or U28157 (N_28157,N_16567,N_12613);
or U28158 (N_28158,N_13824,N_18868);
or U28159 (N_28159,N_11372,N_16372);
nand U28160 (N_28160,N_10839,N_18128);
nand U28161 (N_28161,N_15403,N_15950);
or U28162 (N_28162,N_16467,N_11275);
or U28163 (N_28163,N_16400,N_11693);
nor U28164 (N_28164,N_10909,N_18104);
nor U28165 (N_28165,N_17742,N_13265);
or U28166 (N_28166,N_15913,N_14627);
nor U28167 (N_28167,N_18194,N_18369);
nand U28168 (N_28168,N_16818,N_12358);
nand U28169 (N_28169,N_11425,N_10756);
or U28170 (N_28170,N_19189,N_14318);
nor U28171 (N_28171,N_14426,N_17908);
xnor U28172 (N_28172,N_14944,N_11657);
and U28173 (N_28173,N_11702,N_10679);
nand U28174 (N_28174,N_14110,N_15829);
or U28175 (N_28175,N_19764,N_13034);
xor U28176 (N_28176,N_18447,N_11058);
and U28177 (N_28177,N_18398,N_14241);
and U28178 (N_28178,N_10605,N_12569);
or U28179 (N_28179,N_15871,N_17247);
nor U28180 (N_28180,N_10969,N_19655);
nor U28181 (N_28181,N_13089,N_10026);
or U28182 (N_28182,N_12451,N_17191);
or U28183 (N_28183,N_12074,N_14255);
nand U28184 (N_28184,N_16236,N_10603);
xnor U28185 (N_28185,N_16242,N_11742);
xor U28186 (N_28186,N_19823,N_13174);
xor U28187 (N_28187,N_14608,N_19311);
and U28188 (N_28188,N_17010,N_11756);
or U28189 (N_28189,N_17115,N_15321);
xor U28190 (N_28190,N_10230,N_10801);
or U28191 (N_28191,N_14302,N_15950);
and U28192 (N_28192,N_19909,N_11350);
and U28193 (N_28193,N_12245,N_10125);
or U28194 (N_28194,N_10573,N_10259);
nand U28195 (N_28195,N_19355,N_14043);
xor U28196 (N_28196,N_18029,N_12947);
and U28197 (N_28197,N_15990,N_19831);
and U28198 (N_28198,N_18786,N_14519);
xor U28199 (N_28199,N_12335,N_19772);
nand U28200 (N_28200,N_18749,N_19743);
or U28201 (N_28201,N_16414,N_10336);
xnor U28202 (N_28202,N_14886,N_19684);
and U28203 (N_28203,N_16533,N_12929);
and U28204 (N_28204,N_19644,N_19716);
nand U28205 (N_28205,N_16553,N_11494);
nor U28206 (N_28206,N_14736,N_14066);
xor U28207 (N_28207,N_14073,N_13768);
nor U28208 (N_28208,N_10189,N_15154);
or U28209 (N_28209,N_13856,N_10583);
and U28210 (N_28210,N_10197,N_19014);
or U28211 (N_28211,N_15648,N_14836);
nand U28212 (N_28212,N_13853,N_17436);
nor U28213 (N_28213,N_19549,N_13124);
nor U28214 (N_28214,N_19030,N_16733);
or U28215 (N_28215,N_11087,N_12882);
xor U28216 (N_28216,N_19486,N_18626);
and U28217 (N_28217,N_17078,N_13632);
nor U28218 (N_28218,N_12404,N_16672);
nand U28219 (N_28219,N_17393,N_10065);
or U28220 (N_28220,N_19045,N_11279);
xnor U28221 (N_28221,N_16054,N_14259);
nor U28222 (N_28222,N_10931,N_15008);
and U28223 (N_28223,N_13412,N_10032);
or U28224 (N_28224,N_10346,N_19276);
nor U28225 (N_28225,N_12125,N_10349);
and U28226 (N_28226,N_11277,N_19007);
and U28227 (N_28227,N_12416,N_11331);
or U28228 (N_28228,N_17752,N_10327);
and U28229 (N_28229,N_19237,N_11429);
nand U28230 (N_28230,N_14276,N_13763);
and U28231 (N_28231,N_10212,N_16736);
and U28232 (N_28232,N_14043,N_11437);
and U28233 (N_28233,N_10936,N_11568);
nand U28234 (N_28234,N_17343,N_18095);
or U28235 (N_28235,N_17872,N_15136);
xor U28236 (N_28236,N_19231,N_16846);
xor U28237 (N_28237,N_18905,N_14155);
and U28238 (N_28238,N_18084,N_19510);
or U28239 (N_28239,N_12055,N_13330);
nand U28240 (N_28240,N_11533,N_19171);
xor U28241 (N_28241,N_18833,N_13921);
xor U28242 (N_28242,N_10542,N_10851);
nand U28243 (N_28243,N_11315,N_12981);
and U28244 (N_28244,N_18493,N_12846);
or U28245 (N_28245,N_13296,N_17331);
and U28246 (N_28246,N_16268,N_10730);
nor U28247 (N_28247,N_13759,N_19799);
nor U28248 (N_28248,N_15042,N_12847);
and U28249 (N_28249,N_15186,N_16596);
nor U28250 (N_28250,N_15812,N_12393);
and U28251 (N_28251,N_17431,N_12072);
xnor U28252 (N_28252,N_19743,N_14289);
nand U28253 (N_28253,N_10020,N_11504);
nor U28254 (N_28254,N_14341,N_12052);
nor U28255 (N_28255,N_11096,N_11823);
nor U28256 (N_28256,N_14449,N_17023);
xnor U28257 (N_28257,N_17370,N_15573);
xor U28258 (N_28258,N_17511,N_19915);
nor U28259 (N_28259,N_18493,N_17292);
nor U28260 (N_28260,N_11643,N_19441);
xor U28261 (N_28261,N_18532,N_11507);
or U28262 (N_28262,N_15684,N_10181);
nor U28263 (N_28263,N_11079,N_10918);
or U28264 (N_28264,N_12470,N_16827);
or U28265 (N_28265,N_13812,N_18390);
nand U28266 (N_28266,N_18567,N_14838);
xnor U28267 (N_28267,N_13419,N_13537);
or U28268 (N_28268,N_12044,N_15065);
nor U28269 (N_28269,N_16353,N_11644);
or U28270 (N_28270,N_15464,N_13789);
nor U28271 (N_28271,N_15419,N_12165);
or U28272 (N_28272,N_18890,N_12677);
xor U28273 (N_28273,N_17751,N_19484);
and U28274 (N_28274,N_19908,N_14394);
or U28275 (N_28275,N_13283,N_16101);
nor U28276 (N_28276,N_16342,N_15536);
and U28277 (N_28277,N_10604,N_18906);
nand U28278 (N_28278,N_15128,N_10653);
nand U28279 (N_28279,N_10178,N_14599);
or U28280 (N_28280,N_12110,N_11499);
or U28281 (N_28281,N_13105,N_13066);
and U28282 (N_28282,N_16554,N_12795);
or U28283 (N_28283,N_15037,N_10723);
or U28284 (N_28284,N_15915,N_17690);
xor U28285 (N_28285,N_17189,N_17121);
xor U28286 (N_28286,N_10474,N_12489);
nand U28287 (N_28287,N_15873,N_11651);
nor U28288 (N_28288,N_15679,N_19288);
xor U28289 (N_28289,N_17749,N_19680);
nand U28290 (N_28290,N_14098,N_15956);
or U28291 (N_28291,N_16223,N_14842);
and U28292 (N_28292,N_13673,N_17809);
and U28293 (N_28293,N_17553,N_19209);
xor U28294 (N_28294,N_11793,N_19400);
nor U28295 (N_28295,N_14542,N_12691);
xnor U28296 (N_28296,N_16617,N_18802);
nor U28297 (N_28297,N_17215,N_11318);
nand U28298 (N_28298,N_13801,N_10968);
nand U28299 (N_28299,N_15251,N_17831);
nand U28300 (N_28300,N_13650,N_19356);
and U28301 (N_28301,N_12734,N_18422);
or U28302 (N_28302,N_13669,N_14624);
nor U28303 (N_28303,N_16513,N_16094);
or U28304 (N_28304,N_16652,N_10279);
xnor U28305 (N_28305,N_11952,N_17938);
and U28306 (N_28306,N_12038,N_18173);
and U28307 (N_28307,N_12800,N_17641);
and U28308 (N_28308,N_10292,N_17837);
and U28309 (N_28309,N_11118,N_14541);
nor U28310 (N_28310,N_18821,N_17352);
nand U28311 (N_28311,N_19963,N_12540);
xnor U28312 (N_28312,N_13750,N_16626);
or U28313 (N_28313,N_14810,N_10836);
nand U28314 (N_28314,N_15965,N_10684);
nand U28315 (N_28315,N_15981,N_16310);
and U28316 (N_28316,N_11468,N_13467);
nand U28317 (N_28317,N_10355,N_12726);
nor U28318 (N_28318,N_14063,N_19268);
xor U28319 (N_28319,N_11686,N_12028);
and U28320 (N_28320,N_17218,N_12142);
and U28321 (N_28321,N_18247,N_11008);
and U28322 (N_28322,N_12146,N_17811);
and U28323 (N_28323,N_10567,N_10735);
xnor U28324 (N_28324,N_11469,N_10964);
xor U28325 (N_28325,N_10403,N_12638);
or U28326 (N_28326,N_18801,N_10495);
nor U28327 (N_28327,N_16624,N_14540);
nand U28328 (N_28328,N_16287,N_10057);
nand U28329 (N_28329,N_17016,N_13897);
nor U28330 (N_28330,N_12788,N_19624);
nor U28331 (N_28331,N_18633,N_10022);
xor U28332 (N_28332,N_11031,N_15561);
xnor U28333 (N_28333,N_13938,N_18361);
and U28334 (N_28334,N_19894,N_14478);
nand U28335 (N_28335,N_16251,N_10442);
xor U28336 (N_28336,N_13193,N_12222);
or U28337 (N_28337,N_11072,N_11663);
nor U28338 (N_28338,N_11808,N_18396);
or U28339 (N_28339,N_19830,N_16665);
or U28340 (N_28340,N_10524,N_13305);
xor U28341 (N_28341,N_11558,N_14861);
and U28342 (N_28342,N_18418,N_18050);
nor U28343 (N_28343,N_19978,N_15854);
or U28344 (N_28344,N_18804,N_17566);
or U28345 (N_28345,N_19901,N_10492);
or U28346 (N_28346,N_16630,N_19123);
and U28347 (N_28347,N_19007,N_18881);
nand U28348 (N_28348,N_19925,N_12428);
or U28349 (N_28349,N_14712,N_10866);
or U28350 (N_28350,N_10781,N_15861);
and U28351 (N_28351,N_19755,N_16553);
or U28352 (N_28352,N_18471,N_13831);
and U28353 (N_28353,N_16513,N_17411);
or U28354 (N_28354,N_13453,N_10695);
nand U28355 (N_28355,N_16588,N_18963);
and U28356 (N_28356,N_19341,N_16011);
and U28357 (N_28357,N_12290,N_17553);
or U28358 (N_28358,N_18404,N_12345);
or U28359 (N_28359,N_16868,N_17261);
xor U28360 (N_28360,N_16475,N_15380);
xnor U28361 (N_28361,N_11227,N_15035);
and U28362 (N_28362,N_18492,N_17729);
xnor U28363 (N_28363,N_17207,N_17896);
nand U28364 (N_28364,N_18555,N_17462);
xor U28365 (N_28365,N_18846,N_11688);
or U28366 (N_28366,N_11378,N_19686);
xnor U28367 (N_28367,N_17290,N_18813);
xnor U28368 (N_28368,N_18889,N_10748);
or U28369 (N_28369,N_17126,N_16332);
xor U28370 (N_28370,N_15726,N_19121);
and U28371 (N_28371,N_11965,N_11223);
or U28372 (N_28372,N_19780,N_19805);
nand U28373 (N_28373,N_17445,N_16055);
and U28374 (N_28374,N_19257,N_14564);
nand U28375 (N_28375,N_13722,N_16677);
and U28376 (N_28376,N_15382,N_11788);
nor U28377 (N_28377,N_14657,N_19554);
xor U28378 (N_28378,N_13181,N_19654);
or U28379 (N_28379,N_12733,N_14732);
nand U28380 (N_28380,N_19936,N_15435);
nand U28381 (N_28381,N_15503,N_18785);
nand U28382 (N_28382,N_11682,N_18884);
nor U28383 (N_28383,N_17640,N_16922);
or U28384 (N_28384,N_18849,N_12908);
nor U28385 (N_28385,N_12676,N_16791);
nand U28386 (N_28386,N_12265,N_16676);
nand U28387 (N_28387,N_17880,N_15378);
or U28388 (N_28388,N_17881,N_15827);
and U28389 (N_28389,N_16246,N_11432);
or U28390 (N_28390,N_14068,N_19553);
or U28391 (N_28391,N_14118,N_13164);
and U28392 (N_28392,N_13764,N_19054);
xnor U28393 (N_28393,N_13188,N_19784);
nand U28394 (N_28394,N_13907,N_15051);
nor U28395 (N_28395,N_19240,N_11279);
xor U28396 (N_28396,N_10414,N_10420);
nor U28397 (N_28397,N_14941,N_14443);
and U28398 (N_28398,N_11135,N_15929);
nand U28399 (N_28399,N_19135,N_19336);
nand U28400 (N_28400,N_15373,N_13655);
and U28401 (N_28401,N_16264,N_11833);
xor U28402 (N_28402,N_19451,N_19246);
nor U28403 (N_28403,N_10924,N_18960);
nand U28404 (N_28404,N_14512,N_18122);
xnor U28405 (N_28405,N_11920,N_12655);
xor U28406 (N_28406,N_11352,N_14631);
xnor U28407 (N_28407,N_10348,N_17776);
nor U28408 (N_28408,N_16004,N_11632);
and U28409 (N_28409,N_13195,N_13931);
xnor U28410 (N_28410,N_14044,N_18454);
or U28411 (N_28411,N_16518,N_16926);
or U28412 (N_28412,N_12320,N_17766);
nand U28413 (N_28413,N_12848,N_19253);
and U28414 (N_28414,N_18077,N_15399);
and U28415 (N_28415,N_19145,N_18054);
or U28416 (N_28416,N_12192,N_14029);
xor U28417 (N_28417,N_11033,N_11402);
or U28418 (N_28418,N_10173,N_17195);
nor U28419 (N_28419,N_12713,N_10469);
xor U28420 (N_28420,N_18776,N_15420);
and U28421 (N_28421,N_13132,N_14068);
and U28422 (N_28422,N_10410,N_14531);
xor U28423 (N_28423,N_11028,N_11429);
and U28424 (N_28424,N_18167,N_11135);
nor U28425 (N_28425,N_13794,N_14309);
or U28426 (N_28426,N_14446,N_16530);
or U28427 (N_28427,N_17419,N_12736);
nand U28428 (N_28428,N_14646,N_15624);
nor U28429 (N_28429,N_13934,N_14257);
nand U28430 (N_28430,N_13709,N_18304);
nor U28431 (N_28431,N_15920,N_16089);
nand U28432 (N_28432,N_10440,N_19422);
and U28433 (N_28433,N_19434,N_10421);
xor U28434 (N_28434,N_18543,N_12742);
or U28435 (N_28435,N_10090,N_17491);
nor U28436 (N_28436,N_15555,N_16733);
nor U28437 (N_28437,N_15250,N_11644);
nand U28438 (N_28438,N_11966,N_13391);
and U28439 (N_28439,N_13982,N_12556);
and U28440 (N_28440,N_16614,N_17436);
nor U28441 (N_28441,N_10202,N_14073);
nand U28442 (N_28442,N_18397,N_15309);
nor U28443 (N_28443,N_10805,N_15078);
nand U28444 (N_28444,N_17779,N_19555);
and U28445 (N_28445,N_16694,N_12825);
xnor U28446 (N_28446,N_17420,N_19894);
and U28447 (N_28447,N_15256,N_15417);
xnor U28448 (N_28448,N_11532,N_15726);
or U28449 (N_28449,N_11293,N_16629);
or U28450 (N_28450,N_12678,N_11929);
or U28451 (N_28451,N_16804,N_19585);
xnor U28452 (N_28452,N_15020,N_12315);
xnor U28453 (N_28453,N_16944,N_16286);
xor U28454 (N_28454,N_11031,N_14653);
or U28455 (N_28455,N_16938,N_15147);
or U28456 (N_28456,N_16042,N_14435);
xor U28457 (N_28457,N_16863,N_10980);
nor U28458 (N_28458,N_18057,N_10282);
or U28459 (N_28459,N_18684,N_14983);
or U28460 (N_28460,N_15895,N_16967);
xor U28461 (N_28461,N_18432,N_11541);
and U28462 (N_28462,N_18239,N_10241);
xor U28463 (N_28463,N_14533,N_19168);
nand U28464 (N_28464,N_11883,N_13183);
or U28465 (N_28465,N_13955,N_15868);
nor U28466 (N_28466,N_18619,N_13897);
nor U28467 (N_28467,N_19376,N_11416);
xor U28468 (N_28468,N_10883,N_19144);
nand U28469 (N_28469,N_17471,N_19162);
or U28470 (N_28470,N_13705,N_14491);
and U28471 (N_28471,N_12199,N_19760);
nor U28472 (N_28472,N_12841,N_12770);
xor U28473 (N_28473,N_13712,N_11025);
and U28474 (N_28474,N_15935,N_15520);
or U28475 (N_28475,N_18618,N_10159);
nor U28476 (N_28476,N_18126,N_13977);
or U28477 (N_28477,N_13623,N_18759);
xnor U28478 (N_28478,N_15618,N_11017);
nor U28479 (N_28479,N_16189,N_16951);
xnor U28480 (N_28480,N_18214,N_18627);
and U28481 (N_28481,N_12988,N_10255);
and U28482 (N_28482,N_11267,N_18148);
xnor U28483 (N_28483,N_17040,N_13818);
nor U28484 (N_28484,N_18854,N_18642);
nor U28485 (N_28485,N_13465,N_11552);
and U28486 (N_28486,N_19970,N_17714);
and U28487 (N_28487,N_17761,N_11096);
nand U28488 (N_28488,N_18491,N_12728);
nand U28489 (N_28489,N_19384,N_15686);
nor U28490 (N_28490,N_15329,N_16467);
and U28491 (N_28491,N_11609,N_10148);
xor U28492 (N_28492,N_19854,N_15291);
nand U28493 (N_28493,N_17232,N_19320);
or U28494 (N_28494,N_15904,N_15321);
or U28495 (N_28495,N_15397,N_12996);
xnor U28496 (N_28496,N_12433,N_12181);
nor U28497 (N_28497,N_11324,N_19462);
and U28498 (N_28498,N_17154,N_10450);
nor U28499 (N_28499,N_19417,N_18388);
xor U28500 (N_28500,N_18454,N_13638);
nor U28501 (N_28501,N_15121,N_17568);
or U28502 (N_28502,N_12651,N_17531);
xnor U28503 (N_28503,N_17047,N_18873);
xnor U28504 (N_28504,N_13554,N_12930);
nand U28505 (N_28505,N_13795,N_19692);
nor U28506 (N_28506,N_16687,N_19786);
nand U28507 (N_28507,N_15426,N_17715);
and U28508 (N_28508,N_17433,N_10972);
xnor U28509 (N_28509,N_15277,N_18402);
nor U28510 (N_28510,N_16964,N_19777);
and U28511 (N_28511,N_11916,N_13714);
nor U28512 (N_28512,N_19214,N_13845);
or U28513 (N_28513,N_18590,N_14803);
nand U28514 (N_28514,N_10119,N_11712);
or U28515 (N_28515,N_11674,N_14628);
xnor U28516 (N_28516,N_15834,N_12653);
xnor U28517 (N_28517,N_16621,N_12172);
nand U28518 (N_28518,N_12349,N_19748);
nand U28519 (N_28519,N_15965,N_14133);
nor U28520 (N_28520,N_15677,N_18656);
nor U28521 (N_28521,N_12290,N_18272);
or U28522 (N_28522,N_19280,N_12682);
and U28523 (N_28523,N_10087,N_15357);
or U28524 (N_28524,N_11957,N_19419);
nor U28525 (N_28525,N_11834,N_11659);
and U28526 (N_28526,N_16534,N_14525);
nand U28527 (N_28527,N_13154,N_15463);
nand U28528 (N_28528,N_17090,N_11484);
nand U28529 (N_28529,N_15949,N_19909);
nor U28530 (N_28530,N_13235,N_12926);
or U28531 (N_28531,N_10346,N_13455);
and U28532 (N_28532,N_12630,N_10479);
and U28533 (N_28533,N_17864,N_19086);
xor U28534 (N_28534,N_14676,N_17713);
or U28535 (N_28535,N_17133,N_11986);
nand U28536 (N_28536,N_11044,N_19564);
xor U28537 (N_28537,N_11296,N_10000);
nor U28538 (N_28538,N_11746,N_19958);
and U28539 (N_28539,N_19854,N_18535);
nor U28540 (N_28540,N_17426,N_18077);
nand U28541 (N_28541,N_11973,N_18849);
and U28542 (N_28542,N_13217,N_17021);
and U28543 (N_28543,N_16675,N_12067);
or U28544 (N_28544,N_17755,N_14885);
nand U28545 (N_28545,N_11353,N_13587);
or U28546 (N_28546,N_12078,N_10088);
or U28547 (N_28547,N_16359,N_13555);
nor U28548 (N_28548,N_11170,N_15052);
and U28549 (N_28549,N_12874,N_13684);
nor U28550 (N_28550,N_10695,N_11065);
and U28551 (N_28551,N_19720,N_13006);
xnor U28552 (N_28552,N_13076,N_19710);
and U28553 (N_28553,N_15904,N_12416);
and U28554 (N_28554,N_13598,N_16813);
nand U28555 (N_28555,N_17703,N_10925);
or U28556 (N_28556,N_19291,N_17692);
nand U28557 (N_28557,N_14878,N_16240);
nand U28558 (N_28558,N_12509,N_15081);
and U28559 (N_28559,N_19980,N_13544);
and U28560 (N_28560,N_18522,N_12437);
nor U28561 (N_28561,N_15059,N_11607);
nand U28562 (N_28562,N_11248,N_17396);
or U28563 (N_28563,N_17969,N_15976);
xnor U28564 (N_28564,N_14990,N_13229);
and U28565 (N_28565,N_19829,N_15048);
nand U28566 (N_28566,N_16140,N_19368);
or U28567 (N_28567,N_11428,N_16250);
and U28568 (N_28568,N_12572,N_18985);
or U28569 (N_28569,N_14024,N_12164);
and U28570 (N_28570,N_12296,N_10258);
or U28571 (N_28571,N_17616,N_11194);
or U28572 (N_28572,N_17380,N_11910);
nand U28573 (N_28573,N_17214,N_11248);
nor U28574 (N_28574,N_15121,N_12875);
and U28575 (N_28575,N_13163,N_15962);
or U28576 (N_28576,N_11362,N_17644);
and U28577 (N_28577,N_11034,N_14194);
xnor U28578 (N_28578,N_15331,N_11624);
xor U28579 (N_28579,N_19230,N_16919);
nand U28580 (N_28580,N_12234,N_13757);
xnor U28581 (N_28581,N_14127,N_17925);
nor U28582 (N_28582,N_14587,N_12606);
and U28583 (N_28583,N_11415,N_13392);
nor U28584 (N_28584,N_18398,N_11526);
and U28585 (N_28585,N_18443,N_14940);
nor U28586 (N_28586,N_12680,N_13773);
xor U28587 (N_28587,N_12645,N_17164);
and U28588 (N_28588,N_11214,N_16312);
nand U28589 (N_28589,N_17239,N_12065);
xor U28590 (N_28590,N_17935,N_16375);
nor U28591 (N_28591,N_19775,N_11296);
or U28592 (N_28592,N_13680,N_16533);
xnor U28593 (N_28593,N_16686,N_10081);
nand U28594 (N_28594,N_17972,N_19196);
nand U28595 (N_28595,N_13470,N_17412);
and U28596 (N_28596,N_14672,N_19597);
and U28597 (N_28597,N_16788,N_17100);
and U28598 (N_28598,N_11544,N_19706);
nand U28599 (N_28599,N_12632,N_14962);
or U28600 (N_28600,N_16249,N_16526);
and U28601 (N_28601,N_12881,N_19610);
and U28602 (N_28602,N_13298,N_13625);
nand U28603 (N_28603,N_12159,N_13220);
or U28604 (N_28604,N_15053,N_19079);
xnor U28605 (N_28605,N_15965,N_16786);
nor U28606 (N_28606,N_14355,N_16589);
and U28607 (N_28607,N_17686,N_19816);
or U28608 (N_28608,N_19388,N_11170);
xnor U28609 (N_28609,N_10798,N_10875);
and U28610 (N_28610,N_14485,N_12976);
nor U28611 (N_28611,N_19662,N_16820);
nand U28612 (N_28612,N_17889,N_18338);
xnor U28613 (N_28613,N_13899,N_12358);
nand U28614 (N_28614,N_19187,N_17697);
nand U28615 (N_28615,N_18266,N_10781);
and U28616 (N_28616,N_13083,N_17650);
nand U28617 (N_28617,N_11204,N_12227);
nand U28618 (N_28618,N_11912,N_13446);
nor U28619 (N_28619,N_15906,N_10453);
xor U28620 (N_28620,N_10232,N_12213);
nand U28621 (N_28621,N_11972,N_10383);
nor U28622 (N_28622,N_10471,N_13189);
nand U28623 (N_28623,N_10387,N_15509);
xnor U28624 (N_28624,N_10778,N_10549);
nand U28625 (N_28625,N_12139,N_13506);
xor U28626 (N_28626,N_14077,N_11168);
xor U28627 (N_28627,N_12629,N_11580);
xor U28628 (N_28628,N_16868,N_19949);
and U28629 (N_28629,N_13199,N_18306);
nor U28630 (N_28630,N_19065,N_10554);
nor U28631 (N_28631,N_13669,N_17341);
and U28632 (N_28632,N_13479,N_12478);
or U28633 (N_28633,N_13970,N_11475);
nand U28634 (N_28634,N_16049,N_19741);
xor U28635 (N_28635,N_13261,N_13323);
nand U28636 (N_28636,N_16736,N_18154);
and U28637 (N_28637,N_16263,N_13296);
and U28638 (N_28638,N_18780,N_14815);
and U28639 (N_28639,N_11507,N_18840);
nand U28640 (N_28640,N_10449,N_19640);
xor U28641 (N_28641,N_19865,N_14054);
xor U28642 (N_28642,N_15765,N_13097);
xor U28643 (N_28643,N_12747,N_19195);
and U28644 (N_28644,N_16527,N_13068);
xor U28645 (N_28645,N_15335,N_15036);
nand U28646 (N_28646,N_15069,N_11113);
nor U28647 (N_28647,N_10021,N_13629);
nor U28648 (N_28648,N_18897,N_17292);
or U28649 (N_28649,N_15448,N_11527);
xor U28650 (N_28650,N_16753,N_10258);
or U28651 (N_28651,N_13604,N_14305);
nor U28652 (N_28652,N_14167,N_18080);
nor U28653 (N_28653,N_13965,N_16972);
nor U28654 (N_28654,N_11049,N_15358);
nor U28655 (N_28655,N_12505,N_11442);
xor U28656 (N_28656,N_15677,N_14395);
or U28657 (N_28657,N_13718,N_11531);
or U28658 (N_28658,N_11848,N_15509);
xor U28659 (N_28659,N_12409,N_17178);
or U28660 (N_28660,N_16743,N_18845);
nand U28661 (N_28661,N_16592,N_19223);
xnor U28662 (N_28662,N_19244,N_17199);
nand U28663 (N_28663,N_15198,N_19043);
nor U28664 (N_28664,N_15006,N_11922);
nor U28665 (N_28665,N_12529,N_18004);
and U28666 (N_28666,N_19399,N_17812);
nand U28667 (N_28667,N_11301,N_13717);
or U28668 (N_28668,N_14986,N_11815);
nor U28669 (N_28669,N_11991,N_17411);
nand U28670 (N_28670,N_15770,N_12656);
and U28671 (N_28671,N_14814,N_17859);
or U28672 (N_28672,N_16991,N_17626);
nor U28673 (N_28673,N_13104,N_13448);
nand U28674 (N_28674,N_13402,N_10829);
nor U28675 (N_28675,N_18615,N_14262);
or U28676 (N_28676,N_16468,N_16198);
nand U28677 (N_28677,N_10683,N_16576);
or U28678 (N_28678,N_10987,N_16979);
nand U28679 (N_28679,N_12017,N_15573);
xor U28680 (N_28680,N_12003,N_13675);
nor U28681 (N_28681,N_18250,N_12989);
xor U28682 (N_28682,N_16866,N_14652);
or U28683 (N_28683,N_14198,N_10934);
and U28684 (N_28684,N_17577,N_10570);
and U28685 (N_28685,N_13750,N_17950);
and U28686 (N_28686,N_12148,N_18796);
xnor U28687 (N_28687,N_13442,N_10343);
nor U28688 (N_28688,N_19709,N_18025);
and U28689 (N_28689,N_17779,N_17157);
or U28690 (N_28690,N_11987,N_15776);
and U28691 (N_28691,N_18208,N_17287);
and U28692 (N_28692,N_11181,N_11768);
or U28693 (N_28693,N_12393,N_14465);
or U28694 (N_28694,N_19218,N_13852);
or U28695 (N_28695,N_11910,N_14832);
xor U28696 (N_28696,N_12827,N_16342);
xor U28697 (N_28697,N_11062,N_19557);
xnor U28698 (N_28698,N_15685,N_14416);
and U28699 (N_28699,N_18500,N_13285);
and U28700 (N_28700,N_16197,N_12833);
or U28701 (N_28701,N_10041,N_18569);
nand U28702 (N_28702,N_13562,N_19002);
nand U28703 (N_28703,N_14401,N_14663);
and U28704 (N_28704,N_15989,N_11392);
nor U28705 (N_28705,N_16591,N_13396);
or U28706 (N_28706,N_10192,N_13452);
and U28707 (N_28707,N_13567,N_13518);
xnor U28708 (N_28708,N_14848,N_15673);
and U28709 (N_28709,N_14105,N_17172);
or U28710 (N_28710,N_10221,N_18690);
or U28711 (N_28711,N_19150,N_14629);
and U28712 (N_28712,N_11891,N_17432);
and U28713 (N_28713,N_17158,N_16788);
nor U28714 (N_28714,N_13494,N_14199);
nor U28715 (N_28715,N_15072,N_18484);
nand U28716 (N_28716,N_12888,N_10877);
and U28717 (N_28717,N_12287,N_15895);
xor U28718 (N_28718,N_17723,N_16373);
xor U28719 (N_28719,N_16122,N_16697);
nand U28720 (N_28720,N_18225,N_11229);
nor U28721 (N_28721,N_18424,N_14930);
xor U28722 (N_28722,N_10614,N_10351);
xnor U28723 (N_28723,N_15673,N_13795);
or U28724 (N_28724,N_19983,N_11133);
nand U28725 (N_28725,N_11202,N_11363);
nand U28726 (N_28726,N_17374,N_19101);
or U28727 (N_28727,N_13864,N_19423);
nand U28728 (N_28728,N_14539,N_19336);
nand U28729 (N_28729,N_16548,N_15599);
nand U28730 (N_28730,N_15216,N_19512);
xor U28731 (N_28731,N_17566,N_13291);
and U28732 (N_28732,N_10624,N_15212);
or U28733 (N_28733,N_19728,N_17990);
or U28734 (N_28734,N_19262,N_13120);
nor U28735 (N_28735,N_17451,N_12918);
and U28736 (N_28736,N_19710,N_12027);
and U28737 (N_28737,N_10089,N_14452);
nor U28738 (N_28738,N_14830,N_18817);
or U28739 (N_28739,N_16991,N_18322);
xor U28740 (N_28740,N_10756,N_16928);
nor U28741 (N_28741,N_13097,N_11997);
nand U28742 (N_28742,N_12991,N_11972);
nand U28743 (N_28743,N_16663,N_18510);
xnor U28744 (N_28744,N_11025,N_15937);
xnor U28745 (N_28745,N_19237,N_19668);
or U28746 (N_28746,N_18025,N_13420);
nand U28747 (N_28747,N_10668,N_17474);
or U28748 (N_28748,N_11581,N_17319);
nor U28749 (N_28749,N_16613,N_19341);
nor U28750 (N_28750,N_10612,N_11369);
xor U28751 (N_28751,N_19813,N_12010);
nor U28752 (N_28752,N_15613,N_13682);
nor U28753 (N_28753,N_14118,N_18702);
and U28754 (N_28754,N_17376,N_16159);
nand U28755 (N_28755,N_13254,N_12176);
xor U28756 (N_28756,N_18631,N_18621);
nand U28757 (N_28757,N_11415,N_15752);
nand U28758 (N_28758,N_10448,N_15128);
xor U28759 (N_28759,N_19508,N_17084);
xnor U28760 (N_28760,N_18152,N_17194);
nand U28761 (N_28761,N_19045,N_10220);
nor U28762 (N_28762,N_16281,N_17158);
or U28763 (N_28763,N_12942,N_12653);
xnor U28764 (N_28764,N_14505,N_11372);
or U28765 (N_28765,N_14816,N_19554);
nand U28766 (N_28766,N_19403,N_18803);
nor U28767 (N_28767,N_12410,N_11517);
nand U28768 (N_28768,N_14626,N_11424);
nand U28769 (N_28769,N_17149,N_17039);
nand U28770 (N_28770,N_17041,N_15454);
or U28771 (N_28771,N_15748,N_19518);
nand U28772 (N_28772,N_12722,N_17778);
or U28773 (N_28773,N_11313,N_17581);
and U28774 (N_28774,N_10221,N_18075);
or U28775 (N_28775,N_11070,N_16713);
nor U28776 (N_28776,N_10873,N_18084);
xnor U28777 (N_28777,N_14187,N_14664);
nand U28778 (N_28778,N_19119,N_17678);
nand U28779 (N_28779,N_15876,N_10609);
or U28780 (N_28780,N_14320,N_18820);
and U28781 (N_28781,N_14109,N_18343);
and U28782 (N_28782,N_15017,N_11581);
and U28783 (N_28783,N_14292,N_17654);
nor U28784 (N_28784,N_10419,N_14833);
or U28785 (N_28785,N_12510,N_12639);
nor U28786 (N_28786,N_14220,N_12790);
or U28787 (N_28787,N_19441,N_12626);
and U28788 (N_28788,N_16924,N_14800);
xor U28789 (N_28789,N_11777,N_12718);
nor U28790 (N_28790,N_11028,N_10567);
xor U28791 (N_28791,N_17373,N_10135);
xnor U28792 (N_28792,N_16584,N_16683);
nor U28793 (N_28793,N_14171,N_10583);
xor U28794 (N_28794,N_16127,N_13824);
or U28795 (N_28795,N_13002,N_18598);
or U28796 (N_28796,N_11183,N_17938);
or U28797 (N_28797,N_12665,N_11723);
xor U28798 (N_28798,N_14344,N_12535);
nand U28799 (N_28799,N_12463,N_19466);
or U28800 (N_28800,N_16672,N_19321);
and U28801 (N_28801,N_13196,N_17039);
xor U28802 (N_28802,N_11621,N_12466);
nand U28803 (N_28803,N_12457,N_11646);
xor U28804 (N_28804,N_16008,N_10944);
and U28805 (N_28805,N_11476,N_17086);
or U28806 (N_28806,N_17532,N_17296);
xor U28807 (N_28807,N_10993,N_16487);
or U28808 (N_28808,N_17588,N_11618);
nor U28809 (N_28809,N_15455,N_17362);
and U28810 (N_28810,N_18561,N_15248);
or U28811 (N_28811,N_10303,N_16096);
or U28812 (N_28812,N_16187,N_19416);
and U28813 (N_28813,N_12965,N_18747);
nand U28814 (N_28814,N_17949,N_13471);
nand U28815 (N_28815,N_16698,N_16408);
xnor U28816 (N_28816,N_11588,N_14384);
or U28817 (N_28817,N_11657,N_13595);
nand U28818 (N_28818,N_14717,N_18169);
xnor U28819 (N_28819,N_19215,N_15833);
and U28820 (N_28820,N_10588,N_12638);
nand U28821 (N_28821,N_16620,N_15868);
nand U28822 (N_28822,N_19759,N_13029);
xor U28823 (N_28823,N_17350,N_13421);
nor U28824 (N_28824,N_10711,N_13566);
nor U28825 (N_28825,N_11406,N_16092);
or U28826 (N_28826,N_12273,N_12276);
nand U28827 (N_28827,N_16776,N_13500);
xor U28828 (N_28828,N_11797,N_19020);
and U28829 (N_28829,N_10857,N_14595);
or U28830 (N_28830,N_17754,N_11836);
xnor U28831 (N_28831,N_14229,N_10901);
nand U28832 (N_28832,N_18109,N_15256);
nand U28833 (N_28833,N_15773,N_15826);
xnor U28834 (N_28834,N_10274,N_17958);
or U28835 (N_28835,N_18830,N_17989);
nand U28836 (N_28836,N_17456,N_19424);
nor U28837 (N_28837,N_10986,N_19875);
nor U28838 (N_28838,N_12883,N_13586);
or U28839 (N_28839,N_13359,N_15593);
nor U28840 (N_28840,N_12143,N_10585);
nand U28841 (N_28841,N_15041,N_15642);
and U28842 (N_28842,N_14796,N_18034);
nor U28843 (N_28843,N_11181,N_12780);
xnor U28844 (N_28844,N_14256,N_13187);
xnor U28845 (N_28845,N_18608,N_10639);
xnor U28846 (N_28846,N_15968,N_13720);
nor U28847 (N_28847,N_14644,N_12331);
xor U28848 (N_28848,N_19673,N_19926);
nand U28849 (N_28849,N_18277,N_16837);
xnor U28850 (N_28850,N_17756,N_19467);
and U28851 (N_28851,N_17471,N_15674);
nand U28852 (N_28852,N_11884,N_12380);
and U28853 (N_28853,N_17707,N_18349);
and U28854 (N_28854,N_19355,N_13509);
or U28855 (N_28855,N_15180,N_11009);
nor U28856 (N_28856,N_13792,N_14815);
nor U28857 (N_28857,N_12249,N_11291);
xor U28858 (N_28858,N_17857,N_11153);
nand U28859 (N_28859,N_14773,N_18577);
and U28860 (N_28860,N_11186,N_12512);
xor U28861 (N_28861,N_10924,N_15345);
nor U28862 (N_28862,N_14683,N_13377);
and U28863 (N_28863,N_12252,N_19068);
nor U28864 (N_28864,N_18531,N_12100);
nor U28865 (N_28865,N_11426,N_11943);
nand U28866 (N_28866,N_12415,N_16441);
nor U28867 (N_28867,N_17704,N_15642);
nor U28868 (N_28868,N_16384,N_18299);
xnor U28869 (N_28869,N_14938,N_12914);
nand U28870 (N_28870,N_12192,N_19049);
xor U28871 (N_28871,N_13252,N_10270);
nor U28872 (N_28872,N_15498,N_12531);
xor U28873 (N_28873,N_13040,N_13284);
or U28874 (N_28874,N_18190,N_16039);
xnor U28875 (N_28875,N_11667,N_13842);
xnor U28876 (N_28876,N_19002,N_13929);
or U28877 (N_28877,N_14603,N_18096);
xor U28878 (N_28878,N_11472,N_18419);
or U28879 (N_28879,N_11775,N_15134);
xor U28880 (N_28880,N_19177,N_12131);
or U28881 (N_28881,N_11489,N_14118);
xor U28882 (N_28882,N_11541,N_18681);
nand U28883 (N_28883,N_11168,N_11990);
nor U28884 (N_28884,N_10866,N_16221);
nand U28885 (N_28885,N_16131,N_17739);
xnor U28886 (N_28886,N_11187,N_13741);
or U28887 (N_28887,N_15917,N_14322);
and U28888 (N_28888,N_16135,N_11022);
nor U28889 (N_28889,N_19225,N_14797);
nand U28890 (N_28890,N_14830,N_14781);
nand U28891 (N_28891,N_10586,N_11317);
nor U28892 (N_28892,N_10601,N_11827);
nor U28893 (N_28893,N_11873,N_15596);
xor U28894 (N_28894,N_10895,N_13348);
or U28895 (N_28895,N_14501,N_16856);
nand U28896 (N_28896,N_15367,N_13486);
or U28897 (N_28897,N_18622,N_16082);
and U28898 (N_28898,N_11213,N_14846);
nor U28899 (N_28899,N_19915,N_16253);
xor U28900 (N_28900,N_10611,N_17798);
and U28901 (N_28901,N_14469,N_19700);
nor U28902 (N_28902,N_12366,N_17406);
xor U28903 (N_28903,N_18542,N_11018);
or U28904 (N_28904,N_15490,N_19218);
nand U28905 (N_28905,N_16759,N_17696);
nor U28906 (N_28906,N_17315,N_11283);
xor U28907 (N_28907,N_11073,N_16593);
and U28908 (N_28908,N_12925,N_17829);
and U28909 (N_28909,N_19708,N_15059);
xnor U28910 (N_28910,N_15179,N_18412);
xor U28911 (N_28911,N_10886,N_14325);
xor U28912 (N_28912,N_17645,N_10643);
xor U28913 (N_28913,N_13031,N_19712);
nand U28914 (N_28914,N_10211,N_17200);
and U28915 (N_28915,N_13196,N_16113);
and U28916 (N_28916,N_10772,N_14206);
nor U28917 (N_28917,N_16816,N_19687);
xnor U28918 (N_28918,N_11028,N_10521);
and U28919 (N_28919,N_16837,N_17687);
xnor U28920 (N_28920,N_15547,N_17811);
nand U28921 (N_28921,N_13991,N_19003);
and U28922 (N_28922,N_15043,N_19633);
and U28923 (N_28923,N_15417,N_15160);
nor U28924 (N_28924,N_12108,N_11453);
nor U28925 (N_28925,N_15038,N_14242);
nand U28926 (N_28926,N_10594,N_18496);
xnor U28927 (N_28927,N_13944,N_15898);
xnor U28928 (N_28928,N_17894,N_11924);
and U28929 (N_28929,N_18158,N_18268);
xor U28930 (N_28930,N_12265,N_17113);
or U28931 (N_28931,N_11562,N_16898);
nor U28932 (N_28932,N_13827,N_13342);
nor U28933 (N_28933,N_16724,N_10870);
or U28934 (N_28934,N_13484,N_18524);
and U28935 (N_28935,N_17103,N_17793);
nand U28936 (N_28936,N_15632,N_10364);
xor U28937 (N_28937,N_16341,N_18631);
nor U28938 (N_28938,N_10219,N_18295);
nor U28939 (N_28939,N_14501,N_13590);
nand U28940 (N_28940,N_13834,N_18036);
xor U28941 (N_28941,N_13150,N_12440);
and U28942 (N_28942,N_14837,N_15161);
or U28943 (N_28943,N_12472,N_17871);
xor U28944 (N_28944,N_15594,N_11640);
and U28945 (N_28945,N_10172,N_14487);
xor U28946 (N_28946,N_18903,N_16248);
nand U28947 (N_28947,N_14813,N_12757);
xor U28948 (N_28948,N_14606,N_13847);
xor U28949 (N_28949,N_14555,N_17774);
or U28950 (N_28950,N_16332,N_17370);
xor U28951 (N_28951,N_13669,N_11223);
nor U28952 (N_28952,N_15831,N_11486);
and U28953 (N_28953,N_11385,N_15227);
and U28954 (N_28954,N_14226,N_17050);
or U28955 (N_28955,N_15630,N_16791);
nand U28956 (N_28956,N_15241,N_18461);
nor U28957 (N_28957,N_16601,N_11746);
or U28958 (N_28958,N_10898,N_16917);
nor U28959 (N_28959,N_17306,N_12788);
xnor U28960 (N_28960,N_19815,N_15898);
nor U28961 (N_28961,N_14746,N_17267);
xor U28962 (N_28962,N_15869,N_18946);
nand U28963 (N_28963,N_19178,N_14162);
xor U28964 (N_28964,N_11588,N_14778);
xnor U28965 (N_28965,N_18545,N_19970);
xor U28966 (N_28966,N_14343,N_13077);
nand U28967 (N_28967,N_18660,N_11675);
nand U28968 (N_28968,N_10082,N_19667);
xor U28969 (N_28969,N_11232,N_14528);
nor U28970 (N_28970,N_17261,N_18997);
and U28971 (N_28971,N_19543,N_18889);
nand U28972 (N_28972,N_19024,N_11032);
nand U28973 (N_28973,N_14636,N_10037);
nand U28974 (N_28974,N_10521,N_19094);
and U28975 (N_28975,N_11093,N_17774);
nor U28976 (N_28976,N_16033,N_14913);
nand U28977 (N_28977,N_11055,N_19507);
or U28978 (N_28978,N_10506,N_11990);
or U28979 (N_28979,N_12602,N_19211);
xnor U28980 (N_28980,N_12103,N_19100);
nor U28981 (N_28981,N_13820,N_11074);
and U28982 (N_28982,N_11812,N_16091);
nor U28983 (N_28983,N_18499,N_18107);
nor U28984 (N_28984,N_13025,N_16811);
xnor U28985 (N_28985,N_13248,N_17837);
or U28986 (N_28986,N_10395,N_14223);
or U28987 (N_28987,N_11505,N_14548);
xor U28988 (N_28988,N_19695,N_16963);
nor U28989 (N_28989,N_12351,N_11394);
or U28990 (N_28990,N_14085,N_13395);
or U28991 (N_28991,N_12900,N_15137);
or U28992 (N_28992,N_12681,N_16127);
nand U28993 (N_28993,N_11798,N_12956);
nor U28994 (N_28994,N_17071,N_17162);
nor U28995 (N_28995,N_17422,N_17546);
and U28996 (N_28996,N_18075,N_10280);
xor U28997 (N_28997,N_19598,N_14403);
or U28998 (N_28998,N_10074,N_10640);
xor U28999 (N_28999,N_13780,N_18471);
nor U29000 (N_29000,N_15936,N_16096);
nand U29001 (N_29001,N_15685,N_19138);
xnor U29002 (N_29002,N_16582,N_17722);
nand U29003 (N_29003,N_16023,N_12142);
nand U29004 (N_29004,N_10569,N_13761);
and U29005 (N_29005,N_10197,N_18921);
and U29006 (N_29006,N_16943,N_18211);
xnor U29007 (N_29007,N_13074,N_16965);
xnor U29008 (N_29008,N_12670,N_19521);
nand U29009 (N_29009,N_10196,N_13673);
nand U29010 (N_29010,N_14527,N_18563);
nand U29011 (N_29011,N_18710,N_15593);
nor U29012 (N_29012,N_11417,N_11895);
and U29013 (N_29013,N_15887,N_19530);
xnor U29014 (N_29014,N_17591,N_15338);
and U29015 (N_29015,N_16253,N_13281);
and U29016 (N_29016,N_16254,N_18763);
nor U29017 (N_29017,N_11718,N_10492);
and U29018 (N_29018,N_11886,N_11794);
or U29019 (N_29019,N_11396,N_17963);
nand U29020 (N_29020,N_17167,N_11308);
and U29021 (N_29021,N_12244,N_10567);
xnor U29022 (N_29022,N_18286,N_12370);
and U29023 (N_29023,N_15922,N_10158);
or U29024 (N_29024,N_18035,N_16635);
nand U29025 (N_29025,N_19589,N_19162);
nand U29026 (N_29026,N_19999,N_16092);
nand U29027 (N_29027,N_15096,N_11194);
or U29028 (N_29028,N_19439,N_14285);
and U29029 (N_29029,N_17985,N_12780);
and U29030 (N_29030,N_16299,N_12317);
nand U29031 (N_29031,N_14740,N_12381);
nand U29032 (N_29032,N_18936,N_19992);
xor U29033 (N_29033,N_14536,N_13191);
or U29034 (N_29034,N_16086,N_10785);
nor U29035 (N_29035,N_18410,N_12641);
and U29036 (N_29036,N_12535,N_17675);
nand U29037 (N_29037,N_13804,N_18078);
or U29038 (N_29038,N_12987,N_12763);
nor U29039 (N_29039,N_14051,N_15514);
and U29040 (N_29040,N_12927,N_14065);
nand U29041 (N_29041,N_18048,N_18261);
and U29042 (N_29042,N_19539,N_16144);
or U29043 (N_29043,N_10651,N_13948);
and U29044 (N_29044,N_17572,N_16372);
or U29045 (N_29045,N_10469,N_14919);
xor U29046 (N_29046,N_12859,N_14935);
and U29047 (N_29047,N_18738,N_10224);
and U29048 (N_29048,N_17572,N_12827);
nand U29049 (N_29049,N_16221,N_11989);
xnor U29050 (N_29050,N_14616,N_16204);
nor U29051 (N_29051,N_17436,N_12040);
and U29052 (N_29052,N_15600,N_11608);
and U29053 (N_29053,N_12484,N_11997);
xor U29054 (N_29054,N_10324,N_17389);
nor U29055 (N_29055,N_10146,N_14023);
or U29056 (N_29056,N_10577,N_18174);
nand U29057 (N_29057,N_10033,N_13719);
nor U29058 (N_29058,N_17483,N_17082);
and U29059 (N_29059,N_19721,N_12148);
nor U29060 (N_29060,N_14831,N_11277);
and U29061 (N_29061,N_12608,N_14892);
nand U29062 (N_29062,N_13350,N_13227);
and U29063 (N_29063,N_11879,N_11642);
nor U29064 (N_29064,N_17179,N_17132);
nand U29065 (N_29065,N_12224,N_12251);
nand U29066 (N_29066,N_16893,N_17427);
xnor U29067 (N_29067,N_16925,N_10535);
xor U29068 (N_29068,N_11359,N_19612);
or U29069 (N_29069,N_18685,N_16096);
and U29070 (N_29070,N_11136,N_11842);
nor U29071 (N_29071,N_10440,N_14332);
or U29072 (N_29072,N_10118,N_18632);
nor U29073 (N_29073,N_11299,N_13451);
nand U29074 (N_29074,N_10750,N_14302);
or U29075 (N_29075,N_19868,N_15313);
nand U29076 (N_29076,N_12582,N_18964);
nand U29077 (N_29077,N_15281,N_15664);
and U29078 (N_29078,N_11611,N_16348);
or U29079 (N_29079,N_19323,N_13788);
xor U29080 (N_29080,N_11092,N_16933);
or U29081 (N_29081,N_16113,N_17860);
and U29082 (N_29082,N_18811,N_19816);
xor U29083 (N_29083,N_15310,N_11287);
and U29084 (N_29084,N_19041,N_14420);
and U29085 (N_29085,N_15143,N_15660);
nor U29086 (N_29086,N_18741,N_19312);
nand U29087 (N_29087,N_10458,N_16176);
nor U29088 (N_29088,N_17922,N_10168);
nand U29089 (N_29089,N_12776,N_17708);
and U29090 (N_29090,N_18019,N_16560);
nand U29091 (N_29091,N_18630,N_11989);
xnor U29092 (N_29092,N_14858,N_17970);
nor U29093 (N_29093,N_15808,N_10512);
or U29094 (N_29094,N_13073,N_15362);
and U29095 (N_29095,N_18078,N_15725);
or U29096 (N_29096,N_19805,N_19189);
and U29097 (N_29097,N_15490,N_19880);
and U29098 (N_29098,N_12076,N_15051);
nand U29099 (N_29099,N_15041,N_15696);
nor U29100 (N_29100,N_11409,N_16197);
or U29101 (N_29101,N_15847,N_14705);
xnor U29102 (N_29102,N_18320,N_18343);
nand U29103 (N_29103,N_18452,N_17577);
xnor U29104 (N_29104,N_13556,N_10941);
or U29105 (N_29105,N_16403,N_17923);
xnor U29106 (N_29106,N_17532,N_18364);
nor U29107 (N_29107,N_18028,N_16358);
nand U29108 (N_29108,N_10948,N_16211);
xor U29109 (N_29109,N_18734,N_18062);
nand U29110 (N_29110,N_18007,N_11494);
or U29111 (N_29111,N_19789,N_13716);
xnor U29112 (N_29112,N_11498,N_18209);
xnor U29113 (N_29113,N_18477,N_14479);
xnor U29114 (N_29114,N_15575,N_16386);
nor U29115 (N_29115,N_14034,N_18909);
nor U29116 (N_29116,N_17883,N_18211);
nand U29117 (N_29117,N_18118,N_15845);
nand U29118 (N_29118,N_19248,N_18878);
or U29119 (N_29119,N_11704,N_11732);
nand U29120 (N_29120,N_10315,N_15835);
xnor U29121 (N_29121,N_17842,N_12072);
nand U29122 (N_29122,N_18973,N_10674);
nand U29123 (N_29123,N_17466,N_14289);
or U29124 (N_29124,N_17344,N_12440);
xnor U29125 (N_29125,N_10407,N_10664);
or U29126 (N_29126,N_15020,N_12135);
or U29127 (N_29127,N_13713,N_12048);
nor U29128 (N_29128,N_10094,N_15618);
and U29129 (N_29129,N_16250,N_18017);
xor U29130 (N_29130,N_15150,N_12562);
and U29131 (N_29131,N_18931,N_18350);
and U29132 (N_29132,N_13371,N_11352);
and U29133 (N_29133,N_18123,N_13573);
nor U29134 (N_29134,N_17954,N_18192);
xnor U29135 (N_29135,N_16375,N_19233);
or U29136 (N_29136,N_11120,N_17831);
nand U29137 (N_29137,N_14885,N_14568);
nor U29138 (N_29138,N_10617,N_12236);
nand U29139 (N_29139,N_18614,N_15668);
and U29140 (N_29140,N_16325,N_13284);
nand U29141 (N_29141,N_18048,N_19375);
nor U29142 (N_29142,N_18158,N_12609);
nor U29143 (N_29143,N_15098,N_19653);
nor U29144 (N_29144,N_14675,N_15249);
xnor U29145 (N_29145,N_14532,N_10666);
or U29146 (N_29146,N_17625,N_13330);
or U29147 (N_29147,N_11996,N_12046);
nor U29148 (N_29148,N_14067,N_12745);
or U29149 (N_29149,N_11163,N_11073);
nand U29150 (N_29150,N_11904,N_11175);
nor U29151 (N_29151,N_11048,N_13600);
nor U29152 (N_29152,N_18288,N_14088);
or U29153 (N_29153,N_16473,N_10371);
nand U29154 (N_29154,N_18075,N_12217);
and U29155 (N_29155,N_15811,N_19973);
or U29156 (N_29156,N_19244,N_14663);
xnor U29157 (N_29157,N_12935,N_13634);
or U29158 (N_29158,N_18524,N_12463);
xor U29159 (N_29159,N_15158,N_11381);
xor U29160 (N_29160,N_12965,N_17119);
xor U29161 (N_29161,N_13808,N_11463);
or U29162 (N_29162,N_19954,N_19169);
nor U29163 (N_29163,N_11505,N_17002);
and U29164 (N_29164,N_18772,N_14890);
or U29165 (N_29165,N_14332,N_15866);
nor U29166 (N_29166,N_15549,N_11436);
nand U29167 (N_29167,N_19803,N_16785);
xnor U29168 (N_29168,N_11896,N_13521);
or U29169 (N_29169,N_14461,N_16537);
and U29170 (N_29170,N_19079,N_18636);
or U29171 (N_29171,N_17515,N_18681);
or U29172 (N_29172,N_14479,N_17756);
and U29173 (N_29173,N_15037,N_17008);
or U29174 (N_29174,N_13821,N_11144);
and U29175 (N_29175,N_10996,N_15743);
nor U29176 (N_29176,N_11482,N_13366);
nor U29177 (N_29177,N_10613,N_17137);
nor U29178 (N_29178,N_15728,N_19173);
nor U29179 (N_29179,N_16823,N_19882);
and U29180 (N_29180,N_14859,N_14467);
nand U29181 (N_29181,N_18446,N_16627);
or U29182 (N_29182,N_14213,N_17013);
xnor U29183 (N_29183,N_18917,N_15039);
nand U29184 (N_29184,N_13014,N_11104);
xor U29185 (N_29185,N_18962,N_12590);
and U29186 (N_29186,N_16068,N_10803);
xnor U29187 (N_29187,N_19802,N_12201);
nand U29188 (N_29188,N_10767,N_13277);
nand U29189 (N_29189,N_13609,N_15124);
nor U29190 (N_29190,N_15544,N_19444);
or U29191 (N_29191,N_15855,N_17288);
and U29192 (N_29192,N_11264,N_12621);
or U29193 (N_29193,N_18330,N_18793);
and U29194 (N_29194,N_18768,N_13456);
nand U29195 (N_29195,N_18628,N_13122);
and U29196 (N_29196,N_15697,N_19534);
or U29197 (N_29197,N_13697,N_19874);
xnor U29198 (N_29198,N_17868,N_16741);
nand U29199 (N_29199,N_10892,N_13322);
nand U29200 (N_29200,N_16622,N_15233);
xnor U29201 (N_29201,N_17147,N_17921);
xnor U29202 (N_29202,N_18078,N_10809);
or U29203 (N_29203,N_16185,N_18231);
or U29204 (N_29204,N_14527,N_10581);
nand U29205 (N_29205,N_16385,N_17609);
nor U29206 (N_29206,N_18871,N_12525);
or U29207 (N_29207,N_15244,N_10431);
or U29208 (N_29208,N_14418,N_13904);
and U29209 (N_29209,N_17980,N_10400);
nor U29210 (N_29210,N_11956,N_19944);
xnor U29211 (N_29211,N_18603,N_10064);
or U29212 (N_29212,N_11545,N_13094);
xor U29213 (N_29213,N_15298,N_19295);
nor U29214 (N_29214,N_15443,N_13226);
and U29215 (N_29215,N_11447,N_11034);
nor U29216 (N_29216,N_11323,N_18455);
xnor U29217 (N_29217,N_18836,N_12899);
or U29218 (N_29218,N_15097,N_19368);
and U29219 (N_29219,N_12881,N_11690);
nor U29220 (N_29220,N_10276,N_13903);
xnor U29221 (N_29221,N_11319,N_16472);
nor U29222 (N_29222,N_14098,N_14882);
nand U29223 (N_29223,N_10541,N_17259);
xor U29224 (N_29224,N_19023,N_11499);
xnor U29225 (N_29225,N_15825,N_19021);
and U29226 (N_29226,N_10281,N_16370);
and U29227 (N_29227,N_14444,N_15117);
xnor U29228 (N_29228,N_18219,N_11516);
xnor U29229 (N_29229,N_18247,N_13899);
and U29230 (N_29230,N_19692,N_11927);
and U29231 (N_29231,N_15172,N_18822);
nand U29232 (N_29232,N_14709,N_16398);
and U29233 (N_29233,N_17653,N_18744);
or U29234 (N_29234,N_19392,N_16811);
nand U29235 (N_29235,N_15395,N_17174);
nor U29236 (N_29236,N_12326,N_13964);
nand U29237 (N_29237,N_13401,N_11217);
xnor U29238 (N_29238,N_18218,N_10117);
xor U29239 (N_29239,N_14940,N_14492);
or U29240 (N_29240,N_18368,N_17764);
and U29241 (N_29241,N_12473,N_17360);
and U29242 (N_29242,N_12738,N_17271);
nor U29243 (N_29243,N_19299,N_14251);
and U29244 (N_29244,N_11066,N_14436);
xor U29245 (N_29245,N_19921,N_11389);
or U29246 (N_29246,N_19593,N_15702);
and U29247 (N_29247,N_17922,N_16582);
nor U29248 (N_29248,N_16183,N_18730);
nor U29249 (N_29249,N_14186,N_13166);
and U29250 (N_29250,N_11024,N_14747);
or U29251 (N_29251,N_17828,N_15832);
or U29252 (N_29252,N_17923,N_15776);
and U29253 (N_29253,N_12633,N_19114);
and U29254 (N_29254,N_18536,N_17033);
xnor U29255 (N_29255,N_16973,N_11578);
nand U29256 (N_29256,N_17556,N_12316);
or U29257 (N_29257,N_16259,N_13067);
or U29258 (N_29258,N_19906,N_15676);
and U29259 (N_29259,N_10603,N_14028);
and U29260 (N_29260,N_15988,N_19930);
and U29261 (N_29261,N_16064,N_18120);
or U29262 (N_29262,N_17222,N_14318);
nand U29263 (N_29263,N_19577,N_13249);
nor U29264 (N_29264,N_13430,N_11970);
nand U29265 (N_29265,N_13579,N_12256);
nor U29266 (N_29266,N_13311,N_11206);
or U29267 (N_29267,N_16896,N_15894);
or U29268 (N_29268,N_18899,N_12743);
nand U29269 (N_29269,N_13570,N_18688);
nor U29270 (N_29270,N_14047,N_18844);
nor U29271 (N_29271,N_16138,N_17762);
and U29272 (N_29272,N_18474,N_17119);
nand U29273 (N_29273,N_11678,N_10656);
or U29274 (N_29274,N_16066,N_12768);
xnor U29275 (N_29275,N_13384,N_11630);
and U29276 (N_29276,N_11931,N_16868);
xor U29277 (N_29277,N_11025,N_10727);
or U29278 (N_29278,N_11223,N_17158);
nand U29279 (N_29279,N_15001,N_14078);
and U29280 (N_29280,N_10401,N_15487);
and U29281 (N_29281,N_10202,N_14721);
and U29282 (N_29282,N_16732,N_16905);
nor U29283 (N_29283,N_10466,N_19224);
and U29284 (N_29284,N_15210,N_11459);
xor U29285 (N_29285,N_11540,N_15798);
xor U29286 (N_29286,N_10490,N_10532);
nand U29287 (N_29287,N_10502,N_15939);
nor U29288 (N_29288,N_11342,N_19073);
and U29289 (N_29289,N_12128,N_16283);
nor U29290 (N_29290,N_10470,N_11657);
nand U29291 (N_29291,N_17409,N_18832);
nand U29292 (N_29292,N_15706,N_11819);
nand U29293 (N_29293,N_13176,N_17115);
nor U29294 (N_29294,N_13260,N_16150);
nand U29295 (N_29295,N_17577,N_17283);
and U29296 (N_29296,N_13487,N_16997);
nand U29297 (N_29297,N_11765,N_10057);
nand U29298 (N_29298,N_11678,N_11028);
xnor U29299 (N_29299,N_15715,N_12591);
and U29300 (N_29300,N_10288,N_11594);
xor U29301 (N_29301,N_18186,N_18442);
xnor U29302 (N_29302,N_13780,N_11331);
nor U29303 (N_29303,N_14450,N_19433);
or U29304 (N_29304,N_17046,N_11670);
xor U29305 (N_29305,N_13515,N_18646);
nor U29306 (N_29306,N_14109,N_17237);
or U29307 (N_29307,N_13512,N_18915);
nor U29308 (N_29308,N_11004,N_13209);
xnor U29309 (N_29309,N_13563,N_18574);
xnor U29310 (N_29310,N_18759,N_12729);
nand U29311 (N_29311,N_13212,N_17764);
nor U29312 (N_29312,N_12957,N_16302);
nand U29313 (N_29313,N_13749,N_11600);
xor U29314 (N_29314,N_11878,N_15819);
nand U29315 (N_29315,N_19965,N_11076);
nor U29316 (N_29316,N_16553,N_17725);
nor U29317 (N_29317,N_13103,N_13142);
or U29318 (N_29318,N_18176,N_19738);
or U29319 (N_29319,N_10397,N_15735);
or U29320 (N_29320,N_15209,N_14809);
and U29321 (N_29321,N_14067,N_18341);
xor U29322 (N_29322,N_11733,N_13086);
and U29323 (N_29323,N_19839,N_19038);
and U29324 (N_29324,N_19662,N_11741);
xnor U29325 (N_29325,N_10252,N_16173);
xnor U29326 (N_29326,N_13601,N_12437);
and U29327 (N_29327,N_14639,N_11574);
nand U29328 (N_29328,N_16112,N_10920);
xor U29329 (N_29329,N_13298,N_15886);
and U29330 (N_29330,N_16120,N_10743);
nor U29331 (N_29331,N_16704,N_17701);
nor U29332 (N_29332,N_19519,N_11476);
nor U29333 (N_29333,N_10901,N_12058);
and U29334 (N_29334,N_12044,N_16005);
and U29335 (N_29335,N_10652,N_19504);
and U29336 (N_29336,N_11997,N_13895);
and U29337 (N_29337,N_11927,N_16007);
or U29338 (N_29338,N_18971,N_10284);
xor U29339 (N_29339,N_13348,N_16490);
or U29340 (N_29340,N_16230,N_11911);
or U29341 (N_29341,N_19542,N_17931);
and U29342 (N_29342,N_10492,N_15029);
and U29343 (N_29343,N_11510,N_15678);
xor U29344 (N_29344,N_19395,N_14219);
nand U29345 (N_29345,N_10896,N_12424);
and U29346 (N_29346,N_10064,N_13982);
nor U29347 (N_29347,N_10394,N_10319);
or U29348 (N_29348,N_12380,N_10238);
and U29349 (N_29349,N_16106,N_14254);
and U29350 (N_29350,N_13772,N_14740);
nand U29351 (N_29351,N_16740,N_14155);
or U29352 (N_29352,N_19170,N_19513);
nand U29353 (N_29353,N_19325,N_14920);
nor U29354 (N_29354,N_19029,N_19979);
nor U29355 (N_29355,N_11979,N_16728);
or U29356 (N_29356,N_10767,N_14790);
and U29357 (N_29357,N_10648,N_19351);
nor U29358 (N_29358,N_19897,N_13144);
xnor U29359 (N_29359,N_19248,N_17806);
nor U29360 (N_29360,N_17773,N_19084);
nor U29361 (N_29361,N_12148,N_16964);
or U29362 (N_29362,N_12578,N_11977);
nor U29363 (N_29363,N_17665,N_13612);
or U29364 (N_29364,N_13877,N_12405);
xor U29365 (N_29365,N_15652,N_17909);
nor U29366 (N_29366,N_13852,N_18130);
nor U29367 (N_29367,N_12393,N_10213);
or U29368 (N_29368,N_14099,N_16692);
and U29369 (N_29369,N_19657,N_16997);
nand U29370 (N_29370,N_12290,N_17264);
xnor U29371 (N_29371,N_19373,N_10441);
nand U29372 (N_29372,N_17700,N_18710);
and U29373 (N_29373,N_14909,N_13768);
and U29374 (N_29374,N_11083,N_13334);
nor U29375 (N_29375,N_16645,N_10070);
nand U29376 (N_29376,N_18979,N_18925);
and U29377 (N_29377,N_19777,N_11387);
nand U29378 (N_29378,N_17560,N_19594);
nor U29379 (N_29379,N_11986,N_15562);
and U29380 (N_29380,N_10418,N_18739);
nor U29381 (N_29381,N_19409,N_17639);
nand U29382 (N_29382,N_13848,N_11479);
xor U29383 (N_29383,N_18074,N_13097);
nand U29384 (N_29384,N_11993,N_18700);
nand U29385 (N_29385,N_11410,N_16519);
xor U29386 (N_29386,N_14007,N_17811);
or U29387 (N_29387,N_11996,N_19387);
nand U29388 (N_29388,N_19969,N_15822);
nand U29389 (N_29389,N_16941,N_11018);
and U29390 (N_29390,N_17270,N_18750);
and U29391 (N_29391,N_11366,N_19516);
nor U29392 (N_29392,N_11624,N_15274);
and U29393 (N_29393,N_18983,N_12130);
and U29394 (N_29394,N_14088,N_10832);
or U29395 (N_29395,N_14282,N_12621);
nor U29396 (N_29396,N_11675,N_11442);
or U29397 (N_29397,N_14455,N_18843);
nor U29398 (N_29398,N_10999,N_14010);
nand U29399 (N_29399,N_15384,N_12869);
nand U29400 (N_29400,N_17624,N_15559);
nand U29401 (N_29401,N_12572,N_11166);
or U29402 (N_29402,N_14488,N_11197);
and U29403 (N_29403,N_10599,N_10380);
xnor U29404 (N_29404,N_11618,N_14198);
and U29405 (N_29405,N_13153,N_17271);
or U29406 (N_29406,N_13471,N_12898);
nand U29407 (N_29407,N_13903,N_11938);
nor U29408 (N_29408,N_17999,N_18187);
nand U29409 (N_29409,N_14548,N_17497);
nand U29410 (N_29410,N_13728,N_16983);
or U29411 (N_29411,N_15323,N_11877);
or U29412 (N_29412,N_16589,N_15338);
and U29413 (N_29413,N_19615,N_14521);
or U29414 (N_29414,N_16379,N_12867);
xnor U29415 (N_29415,N_10949,N_16083);
nor U29416 (N_29416,N_18994,N_13507);
nor U29417 (N_29417,N_16917,N_16412);
nand U29418 (N_29418,N_10790,N_16736);
or U29419 (N_29419,N_15731,N_14634);
nand U29420 (N_29420,N_10509,N_19471);
xnor U29421 (N_29421,N_19815,N_13823);
nor U29422 (N_29422,N_14282,N_11952);
nor U29423 (N_29423,N_11942,N_15380);
and U29424 (N_29424,N_14978,N_10804);
and U29425 (N_29425,N_18861,N_11471);
and U29426 (N_29426,N_18681,N_18482);
nor U29427 (N_29427,N_13884,N_15319);
xnor U29428 (N_29428,N_14687,N_14428);
xor U29429 (N_29429,N_13969,N_19471);
and U29430 (N_29430,N_18082,N_10302);
and U29431 (N_29431,N_16658,N_12339);
and U29432 (N_29432,N_17087,N_15112);
xnor U29433 (N_29433,N_12058,N_12230);
nand U29434 (N_29434,N_12124,N_17377);
and U29435 (N_29435,N_12507,N_17031);
nor U29436 (N_29436,N_12230,N_16438);
xor U29437 (N_29437,N_12163,N_18560);
and U29438 (N_29438,N_10518,N_19313);
or U29439 (N_29439,N_14315,N_15669);
nor U29440 (N_29440,N_15849,N_10877);
and U29441 (N_29441,N_15363,N_16135);
nand U29442 (N_29442,N_10862,N_15847);
nor U29443 (N_29443,N_16169,N_12232);
or U29444 (N_29444,N_17375,N_13908);
or U29445 (N_29445,N_11845,N_13593);
xor U29446 (N_29446,N_11081,N_18952);
nand U29447 (N_29447,N_16058,N_16897);
and U29448 (N_29448,N_15320,N_19353);
or U29449 (N_29449,N_15505,N_12388);
and U29450 (N_29450,N_19450,N_15814);
nor U29451 (N_29451,N_11332,N_13633);
nor U29452 (N_29452,N_14595,N_12452);
and U29453 (N_29453,N_18216,N_16557);
nand U29454 (N_29454,N_15461,N_16009);
nand U29455 (N_29455,N_16648,N_14534);
nand U29456 (N_29456,N_15508,N_17463);
and U29457 (N_29457,N_19659,N_12362);
nor U29458 (N_29458,N_13397,N_14735);
or U29459 (N_29459,N_11686,N_15233);
nand U29460 (N_29460,N_19215,N_17071);
nor U29461 (N_29461,N_17663,N_14906);
and U29462 (N_29462,N_13850,N_11403);
xnor U29463 (N_29463,N_19147,N_18759);
and U29464 (N_29464,N_16526,N_17322);
nand U29465 (N_29465,N_10093,N_18047);
xor U29466 (N_29466,N_16670,N_11412);
nor U29467 (N_29467,N_15469,N_13415);
or U29468 (N_29468,N_18497,N_19675);
or U29469 (N_29469,N_19021,N_17493);
nor U29470 (N_29470,N_16088,N_18879);
nand U29471 (N_29471,N_17125,N_12573);
xnor U29472 (N_29472,N_18259,N_14482);
xor U29473 (N_29473,N_17135,N_10011);
or U29474 (N_29474,N_13973,N_17261);
nand U29475 (N_29475,N_17065,N_11287);
or U29476 (N_29476,N_13769,N_16915);
nand U29477 (N_29477,N_19587,N_17075);
nor U29478 (N_29478,N_10538,N_16534);
xnor U29479 (N_29479,N_12344,N_16990);
or U29480 (N_29480,N_11122,N_17799);
or U29481 (N_29481,N_14823,N_14766);
xor U29482 (N_29482,N_12430,N_13003);
xor U29483 (N_29483,N_13119,N_13011);
and U29484 (N_29484,N_17225,N_13263);
or U29485 (N_29485,N_11747,N_10717);
or U29486 (N_29486,N_13049,N_15683);
xor U29487 (N_29487,N_15740,N_11651);
and U29488 (N_29488,N_16667,N_15011);
xor U29489 (N_29489,N_17732,N_14531);
nor U29490 (N_29490,N_19096,N_17496);
or U29491 (N_29491,N_18168,N_17563);
nand U29492 (N_29492,N_14947,N_17946);
nor U29493 (N_29493,N_17584,N_10581);
xnor U29494 (N_29494,N_11758,N_17949);
and U29495 (N_29495,N_19524,N_16648);
xnor U29496 (N_29496,N_10873,N_12888);
nand U29497 (N_29497,N_16153,N_19217);
xnor U29498 (N_29498,N_14405,N_13801);
nor U29499 (N_29499,N_16861,N_13667);
nor U29500 (N_29500,N_14205,N_17757);
xor U29501 (N_29501,N_19643,N_16722);
xnor U29502 (N_29502,N_14870,N_11376);
nand U29503 (N_29503,N_12010,N_11456);
nor U29504 (N_29504,N_16920,N_13193);
nor U29505 (N_29505,N_12853,N_19641);
or U29506 (N_29506,N_18906,N_19883);
xnor U29507 (N_29507,N_18685,N_14180);
and U29508 (N_29508,N_19629,N_12529);
xnor U29509 (N_29509,N_18044,N_19210);
or U29510 (N_29510,N_14927,N_17695);
or U29511 (N_29511,N_11881,N_11365);
or U29512 (N_29512,N_19711,N_19947);
xnor U29513 (N_29513,N_10554,N_12968);
and U29514 (N_29514,N_16155,N_13473);
xnor U29515 (N_29515,N_12932,N_15008);
and U29516 (N_29516,N_17383,N_19688);
and U29517 (N_29517,N_16209,N_10805);
xnor U29518 (N_29518,N_18312,N_16193);
nor U29519 (N_29519,N_14205,N_10373);
and U29520 (N_29520,N_10790,N_12425);
or U29521 (N_29521,N_15158,N_15908);
nand U29522 (N_29522,N_10000,N_15972);
and U29523 (N_29523,N_10669,N_12936);
or U29524 (N_29524,N_18738,N_15474);
xnor U29525 (N_29525,N_11353,N_18578);
nand U29526 (N_29526,N_13047,N_10246);
nand U29527 (N_29527,N_13505,N_12117);
nor U29528 (N_29528,N_19107,N_15058);
nand U29529 (N_29529,N_15147,N_13448);
and U29530 (N_29530,N_15039,N_17297);
xnor U29531 (N_29531,N_11064,N_11134);
xor U29532 (N_29532,N_17689,N_18049);
xnor U29533 (N_29533,N_19743,N_15573);
xnor U29534 (N_29534,N_14280,N_18368);
and U29535 (N_29535,N_11597,N_12410);
or U29536 (N_29536,N_17460,N_13507);
xnor U29537 (N_29537,N_18251,N_12144);
xnor U29538 (N_29538,N_13293,N_14454);
nand U29539 (N_29539,N_18494,N_14440);
xor U29540 (N_29540,N_13061,N_12985);
or U29541 (N_29541,N_19817,N_13370);
or U29542 (N_29542,N_13688,N_12993);
nor U29543 (N_29543,N_15604,N_14221);
nand U29544 (N_29544,N_13572,N_18835);
xnor U29545 (N_29545,N_17669,N_12419);
nor U29546 (N_29546,N_12976,N_17449);
nand U29547 (N_29547,N_17477,N_13787);
and U29548 (N_29548,N_11646,N_19063);
nand U29549 (N_29549,N_16199,N_19188);
or U29550 (N_29550,N_19196,N_11134);
nor U29551 (N_29551,N_14958,N_19538);
and U29552 (N_29552,N_10800,N_13129);
and U29553 (N_29553,N_17513,N_12644);
xnor U29554 (N_29554,N_18645,N_12736);
or U29555 (N_29555,N_10601,N_15018);
xnor U29556 (N_29556,N_15886,N_10933);
nand U29557 (N_29557,N_18790,N_19892);
nand U29558 (N_29558,N_13030,N_18810);
and U29559 (N_29559,N_17597,N_11914);
nor U29560 (N_29560,N_13185,N_13396);
nor U29561 (N_29561,N_19121,N_12584);
and U29562 (N_29562,N_18517,N_13814);
nor U29563 (N_29563,N_15725,N_11762);
or U29564 (N_29564,N_12020,N_10387);
nand U29565 (N_29565,N_17856,N_13234);
or U29566 (N_29566,N_11684,N_14260);
nor U29567 (N_29567,N_12866,N_13901);
xor U29568 (N_29568,N_16962,N_18100);
xor U29569 (N_29569,N_18142,N_17788);
nor U29570 (N_29570,N_16332,N_11752);
xnor U29571 (N_29571,N_19908,N_10066);
nor U29572 (N_29572,N_13073,N_12468);
and U29573 (N_29573,N_15805,N_17190);
and U29574 (N_29574,N_15498,N_13130);
xor U29575 (N_29575,N_12638,N_11206);
and U29576 (N_29576,N_16887,N_18688);
xnor U29577 (N_29577,N_18486,N_14868);
or U29578 (N_29578,N_14818,N_16345);
xnor U29579 (N_29579,N_18925,N_14236);
xor U29580 (N_29580,N_18785,N_19402);
or U29581 (N_29581,N_19719,N_12544);
and U29582 (N_29582,N_10543,N_11206);
and U29583 (N_29583,N_14168,N_17637);
nor U29584 (N_29584,N_14310,N_13402);
or U29585 (N_29585,N_12913,N_10987);
nand U29586 (N_29586,N_11721,N_19678);
xnor U29587 (N_29587,N_12761,N_16959);
xnor U29588 (N_29588,N_11785,N_12433);
xnor U29589 (N_29589,N_19583,N_19475);
or U29590 (N_29590,N_12049,N_15501);
nor U29591 (N_29591,N_15716,N_19068);
xnor U29592 (N_29592,N_14944,N_19201);
xor U29593 (N_29593,N_10255,N_13740);
and U29594 (N_29594,N_16523,N_14906);
and U29595 (N_29595,N_18750,N_13769);
and U29596 (N_29596,N_17861,N_14942);
and U29597 (N_29597,N_19252,N_11470);
nand U29598 (N_29598,N_17609,N_11398);
or U29599 (N_29599,N_13779,N_19976);
and U29600 (N_29600,N_15274,N_13292);
or U29601 (N_29601,N_18099,N_19490);
and U29602 (N_29602,N_11568,N_11063);
xnor U29603 (N_29603,N_18486,N_11490);
nand U29604 (N_29604,N_12160,N_19863);
nand U29605 (N_29605,N_18616,N_12782);
xnor U29606 (N_29606,N_19648,N_11220);
xor U29607 (N_29607,N_17536,N_18357);
or U29608 (N_29608,N_11920,N_19586);
or U29609 (N_29609,N_14478,N_15695);
nand U29610 (N_29610,N_11350,N_10509);
nor U29611 (N_29611,N_14025,N_15709);
nor U29612 (N_29612,N_16847,N_11645);
nor U29613 (N_29613,N_19702,N_10749);
nand U29614 (N_29614,N_10317,N_14043);
xnor U29615 (N_29615,N_11773,N_19314);
nand U29616 (N_29616,N_15298,N_15415);
nor U29617 (N_29617,N_10181,N_13752);
or U29618 (N_29618,N_19979,N_12900);
nor U29619 (N_29619,N_18567,N_10117);
xnor U29620 (N_29620,N_14442,N_11315);
or U29621 (N_29621,N_16379,N_16217);
xor U29622 (N_29622,N_17529,N_12716);
xnor U29623 (N_29623,N_12078,N_11076);
nor U29624 (N_29624,N_14663,N_15787);
and U29625 (N_29625,N_15216,N_11967);
nor U29626 (N_29626,N_12895,N_10324);
nand U29627 (N_29627,N_18462,N_17936);
and U29628 (N_29628,N_19229,N_18154);
nor U29629 (N_29629,N_16502,N_19889);
or U29630 (N_29630,N_11009,N_15468);
nand U29631 (N_29631,N_11563,N_11909);
xnor U29632 (N_29632,N_10010,N_11876);
nand U29633 (N_29633,N_13097,N_18277);
nor U29634 (N_29634,N_16186,N_13162);
nor U29635 (N_29635,N_12442,N_13362);
nand U29636 (N_29636,N_14419,N_13713);
nor U29637 (N_29637,N_11647,N_19635);
xor U29638 (N_29638,N_13593,N_14366);
xor U29639 (N_29639,N_18586,N_15964);
nand U29640 (N_29640,N_12548,N_16367);
nor U29641 (N_29641,N_19201,N_18806);
nand U29642 (N_29642,N_16614,N_10313);
and U29643 (N_29643,N_12384,N_11696);
nor U29644 (N_29644,N_11224,N_10795);
nor U29645 (N_29645,N_14669,N_19629);
nor U29646 (N_29646,N_12474,N_10848);
and U29647 (N_29647,N_10174,N_12221);
nor U29648 (N_29648,N_18537,N_15525);
and U29649 (N_29649,N_18625,N_15583);
or U29650 (N_29650,N_19002,N_15647);
or U29651 (N_29651,N_15780,N_12726);
xor U29652 (N_29652,N_17792,N_15317);
and U29653 (N_29653,N_19182,N_12159);
xnor U29654 (N_29654,N_13802,N_10223);
and U29655 (N_29655,N_17314,N_15036);
nand U29656 (N_29656,N_10351,N_14691);
or U29657 (N_29657,N_10252,N_19934);
and U29658 (N_29658,N_18767,N_18158);
nor U29659 (N_29659,N_18070,N_19894);
nand U29660 (N_29660,N_11024,N_19322);
nor U29661 (N_29661,N_11289,N_16209);
xnor U29662 (N_29662,N_14648,N_17078);
xnor U29663 (N_29663,N_18421,N_13475);
or U29664 (N_29664,N_12869,N_15876);
xnor U29665 (N_29665,N_19005,N_19024);
nor U29666 (N_29666,N_10675,N_19882);
or U29667 (N_29667,N_14433,N_13389);
or U29668 (N_29668,N_18251,N_14903);
xor U29669 (N_29669,N_15075,N_14868);
nand U29670 (N_29670,N_19600,N_11119);
or U29671 (N_29671,N_19100,N_12894);
nand U29672 (N_29672,N_17257,N_11951);
xnor U29673 (N_29673,N_13018,N_11461);
xor U29674 (N_29674,N_16510,N_16627);
nor U29675 (N_29675,N_19004,N_12992);
or U29676 (N_29676,N_11221,N_16153);
nand U29677 (N_29677,N_13710,N_13404);
and U29678 (N_29678,N_10353,N_10214);
nand U29679 (N_29679,N_16973,N_11991);
xnor U29680 (N_29680,N_16750,N_13533);
or U29681 (N_29681,N_17404,N_15550);
or U29682 (N_29682,N_15065,N_18898);
nand U29683 (N_29683,N_17279,N_17995);
nand U29684 (N_29684,N_10437,N_14380);
xor U29685 (N_29685,N_10384,N_10529);
and U29686 (N_29686,N_18325,N_16795);
or U29687 (N_29687,N_15424,N_13026);
and U29688 (N_29688,N_14787,N_11517);
nand U29689 (N_29689,N_14450,N_16312);
nand U29690 (N_29690,N_13474,N_19436);
and U29691 (N_29691,N_12345,N_16137);
and U29692 (N_29692,N_13741,N_18661);
nand U29693 (N_29693,N_16707,N_10886);
nor U29694 (N_29694,N_18926,N_12142);
or U29695 (N_29695,N_11392,N_14121);
nand U29696 (N_29696,N_12862,N_19370);
and U29697 (N_29697,N_12508,N_13958);
nor U29698 (N_29698,N_15411,N_17074);
nor U29699 (N_29699,N_13573,N_16187);
and U29700 (N_29700,N_19645,N_18281);
nand U29701 (N_29701,N_15802,N_18290);
or U29702 (N_29702,N_12134,N_12507);
and U29703 (N_29703,N_14139,N_14374);
nor U29704 (N_29704,N_11476,N_10580);
and U29705 (N_29705,N_11097,N_14790);
and U29706 (N_29706,N_19471,N_12658);
and U29707 (N_29707,N_12202,N_12865);
nand U29708 (N_29708,N_19737,N_11563);
xnor U29709 (N_29709,N_11414,N_11378);
and U29710 (N_29710,N_18563,N_17453);
nor U29711 (N_29711,N_12470,N_15178);
and U29712 (N_29712,N_12498,N_16272);
nor U29713 (N_29713,N_14941,N_18716);
and U29714 (N_29714,N_10594,N_19089);
nor U29715 (N_29715,N_15116,N_11965);
and U29716 (N_29716,N_10455,N_14204);
or U29717 (N_29717,N_14753,N_18046);
xnor U29718 (N_29718,N_16414,N_16010);
nand U29719 (N_29719,N_12323,N_18054);
xnor U29720 (N_29720,N_11649,N_16410);
nor U29721 (N_29721,N_16285,N_16215);
nor U29722 (N_29722,N_11104,N_19482);
xnor U29723 (N_29723,N_19928,N_11325);
nand U29724 (N_29724,N_15454,N_14472);
or U29725 (N_29725,N_10873,N_11999);
xor U29726 (N_29726,N_12508,N_13740);
nor U29727 (N_29727,N_19609,N_12969);
nand U29728 (N_29728,N_16043,N_18825);
and U29729 (N_29729,N_19728,N_16630);
or U29730 (N_29730,N_10462,N_16890);
nor U29731 (N_29731,N_16757,N_14255);
nor U29732 (N_29732,N_11595,N_11967);
nand U29733 (N_29733,N_12805,N_15520);
and U29734 (N_29734,N_13759,N_18509);
or U29735 (N_29735,N_10190,N_16552);
xnor U29736 (N_29736,N_11230,N_14406);
or U29737 (N_29737,N_19470,N_16998);
or U29738 (N_29738,N_18171,N_10178);
xor U29739 (N_29739,N_14083,N_13075);
and U29740 (N_29740,N_13330,N_13922);
or U29741 (N_29741,N_12424,N_12776);
or U29742 (N_29742,N_13951,N_18159);
nand U29743 (N_29743,N_14394,N_11453);
nand U29744 (N_29744,N_12164,N_10904);
nand U29745 (N_29745,N_19176,N_12737);
xnor U29746 (N_29746,N_18979,N_15400);
xor U29747 (N_29747,N_10673,N_11574);
or U29748 (N_29748,N_10142,N_11044);
or U29749 (N_29749,N_18387,N_17046);
or U29750 (N_29750,N_17122,N_10738);
and U29751 (N_29751,N_15549,N_12976);
xnor U29752 (N_29752,N_14632,N_13200);
or U29753 (N_29753,N_11089,N_15552);
xor U29754 (N_29754,N_15483,N_12005);
and U29755 (N_29755,N_19837,N_10019);
xor U29756 (N_29756,N_11247,N_14582);
nor U29757 (N_29757,N_14953,N_19668);
or U29758 (N_29758,N_14223,N_18828);
nand U29759 (N_29759,N_19457,N_12469);
and U29760 (N_29760,N_18056,N_15489);
xor U29761 (N_29761,N_10000,N_16788);
nor U29762 (N_29762,N_12253,N_14529);
xnor U29763 (N_29763,N_17758,N_11087);
nor U29764 (N_29764,N_18937,N_10770);
xnor U29765 (N_29765,N_11734,N_14661);
xor U29766 (N_29766,N_15193,N_16503);
xor U29767 (N_29767,N_11991,N_19738);
xor U29768 (N_29768,N_18554,N_17466);
or U29769 (N_29769,N_19141,N_16692);
or U29770 (N_29770,N_18678,N_10920);
xnor U29771 (N_29771,N_10127,N_13404);
nand U29772 (N_29772,N_18316,N_19252);
xor U29773 (N_29773,N_12617,N_12049);
nor U29774 (N_29774,N_18218,N_19131);
and U29775 (N_29775,N_12058,N_16178);
xor U29776 (N_29776,N_15289,N_17198);
and U29777 (N_29777,N_19420,N_13221);
or U29778 (N_29778,N_16233,N_11092);
or U29779 (N_29779,N_10960,N_19508);
nand U29780 (N_29780,N_17848,N_10460);
nand U29781 (N_29781,N_16960,N_16268);
or U29782 (N_29782,N_10965,N_19786);
or U29783 (N_29783,N_13411,N_19664);
xor U29784 (N_29784,N_18056,N_10338);
nand U29785 (N_29785,N_17580,N_15655);
and U29786 (N_29786,N_19404,N_14109);
nand U29787 (N_29787,N_12580,N_14017);
and U29788 (N_29788,N_12841,N_13894);
or U29789 (N_29789,N_10145,N_17281);
or U29790 (N_29790,N_17484,N_13865);
and U29791 (N_29791,N_15366,N_12258);
xnor U29792 (N_29792,N_17704,N_19121);
nor U29793 (N_29793,N_19773,N_10841);
or U29794 (N_29794,N_13670,N_12756);
xnor U29795 (N_29795,N_16706,N_18458);
nor U29796 (N_29796,N_15364,N_10572);
xnor U29797 (N_29797,N_16917,N_11923);
xnor U29798 (N_29798,N_15031,N_10458);
or U29799 (N_29799,N_12682,N_12313);
or U29800 (N_29800,N_17692,N_13651);
nand U29801 (N_29801,N_18295,N_15109);
nand U29802 (N_29802,N_15055,N_15879);
nand U29803 (N_29803,N_12482,N_19824);
or U29804 (N_29804,N_12724,N_15445);
or U29805 (N_29805,N_18849,N_15427);
nand U29806 (N_29806,N_19404,N_10046);
nor U29807 (N_29807,N_18815,N_15589);
xnor U29808 (N_29808,N_12217,N_15162);
nor U29809 (N_29809,N_19361,N_12878);
nor U29810 (N_29810,N_15771,N_15211);
or U29811 (N_29811,N_10291,N_13756);
or U29812 (N_29812,N_19890,N_17843);
or U29813 (N_29813,N_10831,N_16517);
and U29814 (N_29814,N_17146,N_13187);
xnor U29815 (N_29815,N_13144,N_15338);
nor U29816 (N_29816,N_12312,N_15960);
xnor U29817 (N_29817,N_17412,N_15902);
and U29818 (N_29818,N_13933,N_18751);
or U29819 (N_29819,N_13577,N_16896);
nor U29820 (N_29820,N_13391,N_18507);
nand U29821 (N_29821,N_13687,N_10274);
and U29822 (N_29822,N_13028,N_18926);
nor U29823 (N_29823,N_14707,N_15012);
and U29824 (N_29824,N_19933,N_10010);
nor U29825 (N_29825,N_13316,N_17560);
xor U29826 (N_29826,N_12039,N_17330);
nor U29827 (N_29827,N_16069,N_19702);
and U29828 (N_29828,N_14451,N_18083);
nor U29829 (N_29829,N_16313,N_12612);
nand U29830 (N_29830,N_19928,N_13896);
xor U29831 (N_29831,N_16747,N_12053);
and U29832 (N_29832,N_15782,N_12292);
xor U29833 (N_29833,N_13668,N_11180);
nor U29834 (N_29834,N_11119,N_15861);
and U29835 (N_29835,N_10540,N_11287);
xor U29836 (N_29836,N_16460,N_11209);
nand U29837 (N_29837,N_19463,N_17049);
xor U29838 (N_29838,N_19476,N_12892);
nor U29839 (N_29839,N_18464,N_13666);
and U29840 (N_29840,N_18648,N_10685);
or U29841 (N_29841,N_14796,N_17037);
and U29842 (N_29842,N_15371,N_15973);
and U29843 (N_29843,N_11794,N_12406);
or U29844 (N_29844,N_19726,N_15043);
nor U29845 (N_29845,N_18503,N_13506);
or U29846 (N_29846,N_13698,N_13853);
or U29847 (N_29847,N_15578,N_14039);
and U29848 (N_29848,N_15929,N_12664);
or U29849 (N_29849,N_16693,N_15321);
nor U29850 (N_29850,N_11841,N_12888);
or U29851 (N_29851,N_19253,N_14261);
and U29852 (N_29852,N_17748,N_11010);
nand U29853 (N_29853,N_13311,N_17405);
xnor U29854 (N_29854,N_12096,N_19425);
and U29855 (N_29855,N_18307,N_17065);
xor U29856 (N_29856,N_11405,N_14228);
and U29857 (N_29857,N_10530,N_12783);
xor U29858 (N_29858,N_11976,N_16811);
and U29859 (N_29859,N_15856,N_11471);
nor U29860 (N_29860,N_14010,N_10194);
nand U29861 (N_29861,N_13287,N_11788);
and U29862 (N_29862,N_11581,N_19699);
and U29863 (N_29863,N_16561,N_11399);
nand U29864 (N_29864,N_19004,N_19005);
nand U29865 (N_29865,N_17785,N_17621);
and U29866 (N_29866,N_16231,N_13807);
nand U29867 (N_29867,N_13811,N_17831);
or U29868 (N_29868,N_11420,N_14628);
and U29869 (N_29869,N_13170,N_17715);
and U29870 (N_29870,N_17280,N_15692);
or U29871 (N_29871,N_16927,N_16969);
nand U29872 (N_29872,N_14615,N_13212);
and U29873 (N_29873,N_15559,N_17637);
xor U29874 (N_29874,N_14812,N_11781);
and U29875 (N_29875,N_10309,N_14021);
and U29876 (N_29876,N_19229,N_10778);
nor U29877 (N_29877,N_10453,N_18930);
nor U29878 (N_29878,N_17676,N_12457);
xnor U29879 (N_29879,N_13874,N_13264);
or U29880 (N_29880,N_18831,N_19047);
or U29881 (N_29881,N_12522,N_12320);
or U29882 (N_29882,N_16034,N_12201);
and U29883 (N_29883,N_15102,N_16405);
nor U29884 (N_29884,N_19436,N_18957);
nand U29885 (N_29885,N_17186,N_17348);
nor U29886 (N_29886,N_16653,N_14778);
nor U29887 (N_29887,N_17649,N_11536);
nor U29888 (N_29888,N_12781,N_16252);
nor U29889 (N_29889,N_18779,N_19762);
or U29890 (N_29890,N_18479,N_17679);
and U29891 (N_29891,N_12473,N_12776);
nor U29892 (N_29892,N_12045,N_10401);
and U29893 (N_29893,N_10303,N_19796);
or U29894 (N_29894,N_11031,N_16519);
nand U29895 (N_29895,N_10785,N_16860);
or U29896 (N_29896,N_18740,N_15076);
or U29897 (N_29897,N_16591,N_12615);
nor U29898 (N_29898,N_18461,N_15540);
and U29899 (N_29899,N_14225,N_19141);
nor U29900 (N_29900,N_12866,N_19571);
nor U29901 (N_29901,N_15565,N_15154);
or U29902 (N_29902,N_14681,N_19843);
and U29903 (N_29903,N_19182,N_12300);
xor U29904 (N_29904,N_12196,N_19539);
xor U29905 (N_29905,N_17165,N_10893);
nand U29906 (N_29906,N_17221,N_19985);
or U29907 (N_29907,N_10311,N_16260);
or U29908 (N_29908,N_19405,N_15967);
xnor U29909 (N_29909,N_14719,N_13075);
and U29910 (N_29910,N_17284,N_15340);
and U29911 (N_29911,N_11133,N_12440);
and U29912 (N_29912,N_19385,N_10040);
nand U29913 (N_29913,N_17141,N_10610);
or U29914 (N_29914,N_13656,N_18625);
and U29915 (N_29915,N_18615,N_10653);
xnor U29916 (N_29916,N_15163,N_18662);
and U29917 (N_29917,N_11704,N_13839);
and U29918 (N_29918,N_16593,N_14168);
xnor U29919 (N_29919,N_12488,N_10489);
nand U29920 (N_29920,N_19316,N_10939);
nand U29921 (N_29921,N_15626,N_13054);
nor U29922 (N_29922,N_11364,N_12790);
nand U29923 (N_29923,N_18131,N_19893);
nor U29924 (N_29924,N_15808,N_15704);
or U29925 (N_29925,N_15752,N_11927);
nor U29926 (N_29926,N_14324,N_11497);
and U29927 (N_29927,N_16874,N_15715);
nand U29928 (N_29928,N_10848,N_15230);
xor U29929 (N_29929,N_10617,N_17074);
and U29930 (N_29930,N_13735,N_19398);
nand U29931 (N_29931,N_11006,N_15187);
nand U29932 (N_29932,N_16321,N_10194);
xor U29933 (N_29933,N_14148,N_12481);
and U29934 (N_29934,N_17471,N_16270);
nand U29935 (N_29935,N_11614,N_12061);
nor U29936 (N_29936,N_14691,N_10042);
nor U29937 (N_29937,N_18554,N_18566);
and U29938 (N_29938,N_14759,N_19396);
nor U29939 (N_29939,N_18248,N_17091);
nor U29940 (N_29940,N_18851,N_18752);
or U29941 (N_29941,N_14493,N_13550);
and U29942 (N_29942,N_18579,N_16710);
xnor U29943 (N_29943,N_19958,N_16792);
or U29944 (N_29944,N_17472,N_12424);
nand U29945 (N_29945,N_16962,N_19891);
or U29946 (N_29946,N_19570,N_19463);
xor U29947 (N_29947,N_19431,N_13931);
xor U29948 (N_29948,N_18747,N_19888);
or U29949 (N_29949,N_13535,N_13350);
nand U29950 (N_29950,N_19655,N_12129);
nand U29951 (N_29951,N_14438,N_18244);
and U29952 (N_29952,N_16983,N_14376);
nand U29953 (N_29953,N_17463,N_14993);
nor U29954 (N_29954,N_15840,N_10894);
nor U29955 (N_29955,N_18702,N_17607);
or U29956 (N_29956,N_18768,N_14761);
nand U29957 (N_29957,N_13508,N_13033);
nand U29958 (N_29958,N_18595,N_13340);
and U29959 (N_29959,N_10869,N_15174);
nand U29960 (N_29960,N_18243,N_12397);
or U29961 (N_29961,N_11407,N_19924);
nand U29962 (N_29962,N_14667,N_18262);
or U29963 (N_29963,N_18883,N_11812);
or U29964 (N_29964,N_18278,N_16954);
xor U29965 (N_29965,N_15804,N_11780);
and U29966 (N_29966,N_12200,N_17465);
nor U29967 (N_29967,N_14364,N_14028);
xnor U29968 (N_29968,N_19482,N_15763);
xnor U29969 (N_29969,N_18437,N_10364);
nand U29970 (N_29970,N_14760,N_18469);
or U29971 (N_29971,N_19338,N_17186);
and U29972 (N_29972,N_13740,N_19937);
or U29973 (N_29973,N_14565,N_16002);
or U29974 (N_29974,N_18495,N_13204);
nor U29975 (N_29975,N_13693,N_15255);
nand U29976 (N_29976,N_19449,N_13748);
or U29977 (N_29977,N_18684,N_17540);
or U29978 (N_29978,N_14150,N_11967);
or U29979 (N_29979,N_12202,N_12812);
or U29980 (N_29980,N_15448,N_15169);
xor U29981 (N_29981,N_15857,N_13490);
xnor U29982 (N_29982,N_11187,N_13678);
xnor U29983 (N_29983,N_12511,N_18529);
nor U29984 (N_29984,N_18681,N_10804);
xnor U29985 (N_29985,N_12437,N_10361);
and U29986 (N_29986,N_15896,N_10601);
xnor U29987 (N_29987,N_16240,N_13016);
and U29988 (N_29988,N_14301,N_11712);
nand U29989 (N_29989,N_18920,N_18566);
xnor U29990 (N_29990,N_11860,N_15814);
or U29991 (N_29991,N_12501,N_19922);
nor U29992 (N_29992,N_18087,N_18044);
or U29993 (N_29993,N_17057,N_18042);
or U29994 (N_29994,N_14832,N_13370);
xor U29995 (N_29995,N_12208,N_14857);
nor U29996 (N_29996,N_14971,N_15215);
nand U29997 (N_29997,N_10804,N_11439);
and U29998 (N_29998,N_14860,N_18240);
xor U29999 (N_29999,N_13804,N_13507);
or U30000 (N_30000,N_21736,N_29317);
nand U30001 (N_30001,N_29243,N_27737);
nor U30002 (N_30002,N_27694,N_20813);
nor U30003 (N_30003,N_25373,N_25948);
and U30004 (N_30004,N_21338,N_27819);
nor U30005 (N_30005,N_21911,N_26506);
or U30006 (N_30006,N_29244,N_27035);
nor U30007 (N_30007,N_29492,N_21704);
nand U30008 (N_30008,N_20859,N_25952);
or U30009 (N_30009,N_25688,N_22825);
nand U30010 (N_30010,N_25222,N_22436);
nand U30011 (N_30011,N_22195,N_24027);
xnor U30012 (N_30012,N_24625,N_21010);
or U30013 (N_30013,N_22801,N_26598);
nor U30014 (N_30014,N_29905,N_28378);
and U30015 (N_30015,N_25122,N_22311);
and U30016 (N_30016,N_20144,N_26920);
and U30017 (N_30017,N_23358,N_24634);
or U30018 (N_30018,N_25731,N_28329);
or U30019 (N_30019,N_26925,N_26395);
nand U30020 (N_30020,N_22315,N_27452);
or U30021 (N_30021,N_23916,N_29154);
nor U30022 (N_30022,N_29093,N_27173);
nand U30023 (N_30023,N_28614,N_27171);
or U30024 (N_30024,N_29202,N_23478);
or U30025 (N_30025,N_25247,N_20278);
and U30026 (N_30026,N_27266,N_29906);
or U30027 (N_30027,N_25142,N_25683);
or U30028 (N_30028,N_24401,N_28622);
xnor U30029 (N_30029,N_23785,N_29869);
nand U30030 (N_30030,N_21804,N_26803);
xnor U30031 (N_30031,N_27410,N_23963);
nand U30032 (N_30032,N_21958,N_24515);
or U30033 (N_30033,N_23042,N_25910);
nand U30034 (N_30034,N_24667,N_23806);
or U30035 (N_30035,N_28208,N_28305);
xnor U30036 (N_30036,N_20472,N_26829);
nand U30037 (N_30037,N_24534,N_26793);
and U30038 (N_30038,N_28279,N_25821);
or U30039 (N_30039,N_22251,N_21062);
nand U30040 (N_30040,N_27283,N_28187);
xnor U30041 (N_30041,N_23787,N_20412);
nand U30042 (N_30042,N_21087,N_23547);
or U30043 (N_30043,N_29249,N_21796);
xnor U30044 (N_30044,N_27041,N_27004);
xor U30045 (N_30045,N_29727,N_22782);
nand U30046 (N_30046,N_23775,N_29911);
and U30047 (N_30047,N_21583,N_22439);
or U30048 (N_30048,N_26146,N_29238);
nand U30049 (N_30049,N_24519,N_27952);
nor U30050 (N_30050,N_29004,N_22192);
or U30051 (N_30051,N_23540,N_24063);
nor U30052 (N_30052,N_26630,N_22144);
and U30053 (N_30053,N_28884,N_27495);
nor U30054 (N_30054,N_27780,N_26475);
and U30055 (N_30055,N_28625,N_24553);
and U30056 (N_30056,N_23935,N_24783);
and U30057 (N_30057,N_28004,N_21970);
nor U30058 (N_30058,N_27243,N_23119);
xor U30059 (N_30059,N_20673,N_25070);
or U30060 (N_30060,N_28910,N_26875);
nor U30061 (N_30061,N_25524,N_29099);
or U30062 (N_30062,N_27227,N_25543);
nor U30063 (N_30063,N_20799,N_21733);
xor U30064 (N_30064,N_29194,N_26227);
nor U30065 (N_30065,N_22664,N_29731);
nor U30066 (N_30066,N_23772,N_28021);
nor U30067 (N_30067,N_23603,N_25740);
nor U30068 (N_30068,N_21288,N_26125);
nor U30069 (N_30069,N_25190,N_24766);
xnor U30070 (N_30070,N_24296,N_22685);
or U30071 (N_30071,N_25227,N_29551);
nor U30072 (N_30072,N_20196,N_22725);
nor U30073 (N_30073,N_20002,N_27589);
nand U30074 (N_30074,N_24219,N_24500);
xor U30075 (N_30075,N_24838,N_20747);
nor U30076 (N_30076,N_28182,N_28957);
and U30077 (N_30077,N_23304,N_21459);
and U30078 (N_30078,N_21749,N_22169);
xor U30079 (N_30079,N_27645,N_29502);
nor U30080 (N_30080,N_23398,N_27509);
nor U30081 (N_30081,N_21500,N_24335);
xnor U30082 (N_30082,N_25351,N_21417);
and U30083 (N_30083,N_25497,N_24542);
and U30084 (N_30084,N_26690,N_25776);
nand U30085 (N_30085,N_24647,N_24740);
and U30086 (N_30086,N_20214,N_23660);
nor U30087 (N_30087,N_24489,N_21432);
xor U30088 (N_30088,N_20887,N_29797);
or U30089 (N_30089,N_26388,N_27080);
and U30090 (N_30090,N_26197,N_22682);
nand U30091 (N_30091,N_23382,N_28411);
or U30092 (N_30092,N_26709,N_29000);
xor U30093 (N_30093,N_26921,N_29732);
and U30094 (N_30094,N_23548,N_25499);
and U30095 (N_30095,N_26502,N_29356);
xnor U30096 (N_30096,N_21170,N_26302);
xor U30097 (N_30097,N_22493,N_29517);
xor U30098 (N_30098,N_23536,N_28508);
nor U30099 (N_30099,N_24950,N_28976);
xor U30100 (N_30100,N_24019,N_21108);
and U30101 (N_30101,N_27449,N_28521);
and U30102 (N_30102,N_21613,N_22078);
or U30103 (N_30103,N_23172,N_23363);
nor U30104 (N_30104,N_28686,N_29286);
xnor U30105 (N_30105,N_29603,N_25737);
and U30106 (N_30106,N_22843,N_26192);
xor U30107 (N_30107,N_26084,N_20063);
nand U30108 (N_30108,N_23108,N_27650);
and U30109 (N_30109,N_28262,N_22077);
nand U30110 (N_30110,N_21554,N_21348);
nand U30111 (N_30111,N_22827,N_26551);
xnor U30112 (N_30112,N_21446,N_22521);
or U30113 (N_30113,N_20425,N_24986);
xnor U30114 (N_30114,N_29833,N_26979);
and U30115 (N_30115,N_25449,N_29720);
or U30116 (N_30116,N_26474,N_20627);
xor U30117 (N_30117,N_26115,N_25355);
or U30118 (N_30118,N_22928,N_21060);
xnor U30119 (N_30119,N_22022,N_29707);
or U30120 (N_30120,N_25433,N_26618);
and U30121 (N_30121,N_24840,N_26657);
xnor U30122 (N_30122,N_27138,N_28184);
xor U30123 (N_30123,N_28924,N_29148);
or U30124 (N_30124,N_22499,N_24725);
or U30125 (N_30125,N_25513,N_24535);
and U30126 (N_30126,N_23873,N_22502);
or U30127 (N_30127,N_27859,N_21762);
nand U30128 (N_30128,N_24315,N_22866);
nand U30129 (N_30129,N_27318,N_25392);
and U30130 (N_30130,N_24244,N_25824);
nand U30131 (N_30131,N_23589,N_20894);
or U30132 (N_30132,N_24373,N_22904);
nor U30133 (N_30133,N_21548,N_29664);
or U30134 (N_30134,N_24139,N_25055);
or U30135 (N_30135,N_29121,N_24913);
nor U30136 (N_30136,N_28132,N_21519);
nor U30137 (N_30137,N_26007,N_21175);
nor U30138 (N_30138,N_20003,N_24116);
xnor U30139 (N_30139,N_24909,N_28885);
and U30140 (N_30140,N_27064,N_26738);
xor U30141 (N_30141,N_20606,N_26765);
xnor U30142 (N_30142,N_25091,N_20356);
nand U30143 (N_30143,N_20635,N_21824);
xor U30144 (N_30144,N_20619,N_29879);
xnor U30145 (N_30145,N_27541,N_24214);
and U30146 (N_30146,N_26027,N_20744);
xnor U30147 (N_30147,N_26678,N_22349);
or U30148 (N_30148,N_26180,N_25003);
nand U30149 (N_30149,N_28782,N_28531);
or U30150 (N_30150,N_29400,N_22329);
and U30151 (N_30151,N_24754,N_22445);
and U30152 (N_30152,N_21042,N_27553);
and U30153 (N_30153,N_20400,N_23483);
or U30154 (N_30154,N_24097,N_20118);
xnor U30155 (N_30155,N_22853,N_22520);
nand U30156 (N_30156,N_24583,N_28068);
and U30157 (N_30157,N_28160,N_21999);
or U30158 (N_30158,N_26574,N_20485);
or U30159 (N_30159,N_28699,N_28624);
xor U30160 (N_30160,N_26298,N_26129);
and U30161 (N_30161,N_26661,N_23355);
xnor U30162 (N_30162,N_23177,N_21747);
and U30163 (N_30163,N_27336,N_22231);
nor U30164 (N_30164,N_20961,N_21024);
xor U30165 (N_30165,N_27400,N_29451);
nand U30166 (N_30166,N_20071,N_23594);
nor U30167 (N_30167,N_23945,N_26977);
nor U30168 (N_30168,N_22990,N_26255);
or U30169 (N_30169,N_26648,N_24526);
nand U30170 (N_30170,N_25479,N_26567);
nand U30171 (N_30171,N_25897,N_20841);
and U30172 (N_30172,N_24906,N_29967);
nor U30173 (N_30173,N_22792,N_20181);
or U30174 (N_30174,N_26572,N_27195);
nor U30175 (N_30175,N_27028,N_25819);
xor U30176 (N_30176,N_28586,N_26672);
nor U30177 (N_30177,N_20505,N_21306);
nor U30178 (N_30178,N_28309,N_21649);
nor U30179 (N_30179,N_29776,N_28167);
and U30180 (N_30180,N_26570,N_24125);
or U30181 (N_30181,N_23032,N_22126);
and U30182 (N_30182,N_26120,N_27699);
nor U30183 (N_30183,N_21965,N_23324);
xnor U30184 (N_30184,N_28428,N_29354);
nor U30185 (N_30185,N_20678,N_29936);
nor U30186 (N_30186,N_26173,N_27305);
and U30187 (N_30187,N_26465,N_22629);
nand U30188 (N_30188,N_20880,N_26834);
and U30189 (N_30189,N_24105,N_25714);
nor U30190 (N_30190,N_28570,N_25577);
or U30191 (N_30191,N_20090,N_29966);
or U30192 (N_30192,N_21125,N_27657);
nor U30193 (N_30193,N_22809,N_26074);
xnor U30194 (N_30194,N_25949,N_25833);
xnor U30195 (N_30195,N_27221,N_29075);
or U30196 (N_30196,N_26892,N_23998);
nor U30197 (N_30197,N_29842,N_25464);
nand U30198 (N_30198,N_27574,N_23175);
nor U30199 (N_30199,N_24012,N_27775);
nand U30200 (N_30200,N_23939,N_27701);
xnor U30201 (N_30201,N_26396,N_22736);
nor U30202 (N_30202,N_26526,N_21391);
nor U30203 (N_30203,N_29804,N_24473);
nand U30204 (N_30204,N_20232,N_27098);
or U30205 (N_30205,N_27262,N_28331);
xnor U30206 (N_30206,N_26862,N_23724);
xor U30207 (N_30207,N_29634,N_27590);
and U30208 (N_30208,N_25839,N_20420);
nor U30209 (N_30209,N_23243,N_20160);
nand U30210 (N_30210,N_26401,N_20453);
xor U30211 (N_30211,N_24297,N_27597);
and U30212 (N_30212,N_24811,N_29163);
and U30213 (N_30213,N_20106,N_28405);
and U30214 (N_30214,N_24270,N_29239);
nor U30215 (N_30215,N_21028,N_28314);
nor U30216 (N_30216,N_27844,N_26004);
nor U30217 (N_30217,N_26859,N_29704);
and U30218 (N_30218,N_26792,N_28941);
xnor U30219 (N_30219,N_22277,N_20981);
or U30220 (N_30220,N_23327,N_27425);
nand U30221 (N_30221,N_29805,N_22261);
and U30222 (N_30222,N_20138,N_22396);
or U30223 (N_30223,N_21689,N_26922);
nand U30224 (N_30224,N_23598,N_27199);
or U30225 (N_30225,N_22187,N_26536);
xnor U30226 (N_30226,N_22376,N_22540);
and U30227 (N_30227,N_27365,N_29064);
xor U30228 (N_30228,N_21488,N_29612);
nand U30229 (N_30229,N_29611,N_24772);
xnor U30230 (N_30230,N_26616,N_24084);
or U30231 (N_30231,N_20336,N_21284);
nor U30232 (N_30232,N_26868,N_22253);
or U30233 (N_30233,N_28151,N_22858);
xnor U30234 (N_30234,N_20419,N_27571);
nand U30235 (N_30235,N_25257,N_26720);
nand U30236 (N_30236,N_21243,N_24470);
and U30237 (N_30237,N_22587,N_22369);
or U30238 (N_30238,N_23459,N_27334);
or U30239 (N_30239,N_28585,N_26756);
nor U30240 (N_30240,N_21846,N_24308);
xnor U30241 (N_30241,N_26402,N_21771);
xor U30242 (N_30242,N_27757,N_26663);
nand U30243 (N_30243,N_21674,N_22425);
or U30244 (N_30244,N_26256,N_23275);
or U30245 (N_30245,N_22119,N_24719);
nand U30246 (N_30246,N_25229,N_28636);
nor U30247 (N_30247,N_27211,N_21334);
nand U30248 (N_30248,N_28410,N_24452);
and U30249 (N_30249,N_24053,N_28365);
nor U30250 (N_30250,N_20337,N_23608);
nand U30251 (N_30251,N_21561,N_26202);
and U30252 (N_30252,N_29444,N_20967);
nand U30253 (N_30253,N_23303,N_26557);
nand U30254 (N_30254,N_27323,N_29373);
nand U30255 (N_30255,N_20751,N_21217);
nand U30256 (N_30256,N_28790,N_20237);
nand U30257 (N_30257,N_20397,N_26917);
or U30258 (N_30258,N_20818,N_22469);
nand U30259 (N_30259,N_23588,N_24806);
nor U30260 (N_30260,N_22008,N_27889);
or U30261 (N_30261,N_22748,N_27263);
xnor U30262 (N_30262,N_20948,N_28598);
or U30263 (N_30263,N_28210,N_24919);
xnor U30264 (N_30264,N_27248,N_22173);
and U30265 (N_30265,N_22756,N_21345);
xnor U30266 (N_30266,N_25427,N_25525);
and U30267 (N_30267,N_25841,N_22970);
nor U30268 (N_30268,N_29604,N_21027);
nand U30269 (N_30269,N_25000,N_26527);
and U30270 (N_30270,N_21317,N_22494);
or U30271 (N_30271,N_24467,N_28389);
nor U30272 (N_30272,N_24414,N_28883);
xnor U30273 (N_30273,N_21399,N_28766);
or U30274 (N_30274,N_26975,N_24856);
and U30275 (N_30275,N_26232,N_22006);
and U30276 (N_30276,N_26309,N_24355);
xor U30277 (N_30277,N_22863,N_21420);
and U30278 (N_30278,N_20631,N_24872);
nand U30279 (N_30279,N_27594,N_23635);
or U30280 (N_30280,N_20504,N_29207);
xor U30281 (N_30281,N_25377,N_23212);
or U30282 (N_30282,N_23720,N_21489);
nor U30283 (N_30283,N_26887,N_22010);
or U30284 (N_30284,N_28731,N_25183);
and U30285 (N_30285,N_26705,N_21408);
xnor U30286 (N_30286,N_25958,N_23912);
nand U30287 (N_30287,N_27261,N_21894);
or U30288 (N_30288,N_22818,N_23696);
xnor U30289 (N_30289,N_20441,N_28078);
nor U30290 (N_30290,N_24585,N_28089);
nor U30291 (N_30291,N_27569,N_26906);
xor U30292 (N_30292,N_23083,N_24372);
nand U30293 (N_30293,N_24817,N_26441);
xnor U30294 (N_30294,N_26942,N_20262);
and U30295 (N_30295,N_25665,N_20695);
nor U30296 (N_30296,N_27133,N_22754);
or U30297 (N_30297,N_26766,N_27249);
and U30298 (N_30298,N_24521,N_25586);
and U30299 (N_30299,N_29985,N_23490);
xnor U30300 (N_30300,N_23665,N_25324);
nor U30301 (N_30301,N_21422,N_20568);
and U30302 (N_30302,N_27577,N_20333);
or U30303 (N_30303,N_27386,N_23843);
and U30304 (N_30304,N_21695,N_24656);
nand U30305 (N_30305,N_21315,N_27142);
and U30306 (N_30306,N_29042,N_23493);
or U30307 (N_30307,N_21002,N_27457);
nand U30308 (N_30308,N_27743,N_21651);
and U30309 (N_30309,N_28606,N_29170);
and U30310 (N_30310,N_25342,N_26322);
nor U30311 (N_30311,N_26500,N_22992);
xnor U30312 (N_30312,N_28162,N_24700);
nand U30313 (N_30313,N_23612,N_28181);
xor U30314 (N_30314,N_20285,N_25837);
xnor U30315 (N_30315,N_29161,N_27114);
or U30316 (N_30316,N_24215,N_22908);
or U30317 (N_30317,N_24490,N_20559);
xor U30318 (N_30318,N_23114,N_27271);
nor U30319 (N_30319,N_28874,N_24112);
xnor U30320 (N_30320,N_20642,N_29224);
nand U30321 (N_30321,N_26050,N_25167);
or U30322 (N_30322,N_21298,N_23021);
nand U30323 (N_30323,N_23579,N_20884);
or U30324 (N_30324,N_29076,N_20348);
nand U30325 (N_30325,N_21957,N_29119);
xnor U30326 (N_30326,N_29717,N_20035);
nor U30327 (N_30327,N_26400,N_25307);
nor U30328 (N_30328,N_23826,N_25706);
nor U30329 (N_30329,N_25490,N_25083);
xor U30330 (N_30330,N_26193,N_28859);
nor U30331 (N_30331,N_22586,N_26196);
or U30332 (N_30332,N_27402,N_22063);
xor U30333 (N_30333,N_27084,N_21173);
and U30334 (N_30334,N_29234,N_25571);
nand U30335 (N_30335,N_21126,N_28308);
or U30336 (N_30336,N_21429,N_21910);
nor U30337 (N_30337,N_22117,N_26316);
xnor U30338 (N_30338,N_25096,N_28930);
and U30339 (N_30339,N_23088,N_25795);
or U30340 (N_30340,N_28943,N_29722);
or U30341 (N_30341,N_22563,N_21735);
and U30342 (N_30342,N_22501,N_25651);
xnor U30343 (N_30343,N_24374,N_28303);
nand U30344 (N_30344,N_24514,N_24967);
nand U30345 (N_30345,N_25446,N_27346);
xnor U30346 (N_30346,N_25905,N_21169);
nor U30347 (N_30347,N_29606,N_26848);
xnor U30348 (N_30348,N_24680,N_25878);
and U30349 (N_30349,N_25850,N_20726);
or U30350 (N_30350,N_24358,N_24261);
nor U30351 (N_30351,N_27347,N_28447);
nor U30352 (N_30352,N_20329,N_22532);
nor U30353 (N_30353,N_24032,N_28524);
nand U30354 (N_30354,N_29783,N_27315);
nand U30355 (N_30355,N_28295,N_25738);
nand U30356 (N_30356,N_23819,N_21642);
xnor U30357 (N_30357,N_28652,N_29706);
nand U30358 (N_30358,N_20561,N_25058);
or U30359 (N_30359,N_25644,N_23139);
xor U30360 (N_30360,N_21073,N_29149);
and U30361 (N_30361,N_27514,N_22097);
and U30362 (N_30362,N_21775,N_23052);
nor U30363 (N_30363,N_23049,N_22623);
nor U30364 (N_30364,N_20513,N_27893);
or U30365 (N_30365,N_25606,N_21692);
nand U30366 (N_30366,N_25283,N_27061);
xor U30367 (N_30367,N_23979,N_21938);
and U30368 (N_30368,N_29900,N_24092);
xor U30369 (N_30369,N_23118,N_27135);
nand U30370 (N_30370,N_20649,N_20815);
xor U30371 (N_30371,N_27710,N_25260);
nor U30372 (N_30372,N_23600,N_23408);
and U30373 (N_30373,N_22226,N_25434);
nor U30374 (N_30374,N_26121,N_21301);
xnor U30375 (N_30375,N_27825,N_23312);
and U30376 (N_30376,N_23499,N_22463);
nor U30377 (N_30377,N_20448,N_20620);
xnor U30378 (N_30378,N_23976,N_28933);
nor U30379 (N_30379,N_26505,N_29640);
nand U30380 (N_30380,N_28090,N_20896);
nand U30381 (N_30381,N_28115,N_25539);
nor U30382 (N_30382,N_26640,N_25541);
or U30383 (N_30383,N_24235,N_26960);
nand U30384 (N_30384,N_25855,N_20767);
or U30385 (N_30385,N_20738,N_29363);
xnor U30386 (N_30386,N_26362,N_29488);
nand U30387 (N_30387,N_27802,N_23271);
or U30388 (N_30388,N_29065,N_21133);
xor U30389 (N_30389,N_24283,N_24733);
or U30390 (N_30390,N_23410,N_21457);
xor U30391 (N_30391,N_22161,N_29445);
or U30392 (N_30392,N_29933,N_24353);
nor U30393 (N_30393,N_25925,N_22118);
nand U30394 (N_30394,N_23395,N_20427);
and U30395 (N_30395,N_29775,N_26160);
nand U30396 (N_30396,N_20811,N_24339);
nand U30397 (N_30397,N_26449,N_26753);
and U30398 (N_30398,N_25781,N_25242);
or U30399 (N_30399,N_22609,N_26870);
nand U30400 (N_30400,N_21978,N_22994);
nand U30401 (N_30401,N_25898,N_21037);
xor U30402 (N_30402,N_27647,N_27534);
or U30403 (N_30403,N_23313,N_20178);
nor U30404 (N_30404,N_27122,N_23448);
and U30405 (N_30405,N_22945,N_20770);
and U30406 (N_30406,N_21623,N_23704);
or U30407 (N_30407,N_20552,N_28207);
nor U30408 (N_30408,N_21964,N_23325);
or U30409 (N_30409,N_26021,N_25483);
or U30410 (N_30410,N_21951,N_21770);
nor U30411 (N_30411,N_21461,N_20509);
or U30412 (N_30412,N_22874,N_29029);
nand U30413 (N_30413,N_21293,N_20174);
nor U30414 (N_30414,N_28798,N_21874);
xor U30415 (N_30415,N_23283,N_27210);
nand U30416 (N_30416,N_21349,N_25405);
or U30417 (N_30417,N_28734,N_21249);
and U30418 (N_30418,N_28268,N_28890);
or U30419 (N_30419,N_22073,N_25144);
nand U30420 (N_30420,N_24759,N_20790);
xor U30421 (N_30421,N_29630,N_20360);
nand U30422 (N_30422,N_24411,N_22290);
nor U30423 (N_30423,N_24403,N_26123);
and U30424 (N_30424,N_29629,N_26980);
nor U30425 (N_30425,N_26175,N_23040);
and U30426 (N_30426,N_23809,N_24461);
nand U30427 (N_30427,N_25649,N_28043);
xor U30428 (N_30428,N_25224,N_28876);
or U30429 (N_30429,N_28176,N_29235);
and U30430 (N_30430,N_23747,N_20468);
xor U30431 (N_30431,N_23872,N_20184);
xnor U30432 (N_30432,N_25179,N_22316);
or U30433 (N_30433,N_24338,N_29068);
or U30434 (N_30434,N_23610,N_20394);
and U30435 (N_30435,N_26907,N_22106);
nor U30436 (N_30436,N_28178,N_26219);
nor U30437 (N_30437,N_27504,N_23035);
nand U30438 (N_30438,N_24047,N_25274);
and U30439 (N_30439,N_25961,N_22632);
and U30440 (N_30440,N_26546,N_23427);
nor U30441 (N_30441,N_23102,N_28581);
xnor U30442 (N_30442,N_20550,N_28947);
and U30443 (N_30443,N_25888,N_27515);
xor U30444 (N_30444,N_23260,N_24511);
or U30445 (N_30445,N_28364,N_24712);
nand U30446 (N_30446,N_29590,N_25895);
or U30447 (N_30447,N_23498,N_29114);
xnor U30448 (N_30448,N_28845,N_27938);
or U30449 (N_30449,N_28568,N_29398);
nor U30450 (N_30450,N_27911,N_29394);
or U30451 (N_30451,N_22602,N_28402);
and U30452 (N_30452,N_26884,N_24937);
nand U30453 (N_30453,N_20656,N_27726);
nor U30454 (N_30454,N_27126,N_29728);
xnor U30455 (N_30455,N_28227,N_22556);
and U30456 (N_30456,N_29292,N_27872);
nand U30457 (N_30457,N_27218,N_27115);
or U30458 (N_30458,N_21036,N_22003);
nand U30459 (N_30459,N_23160,N_21632);
and U30460 (N_30460,N_22570,N_28399);
or U30461 (N_30461,N_29272,N_29669);
or U30462 (N_30462,N_29493,N_27018);
and U30463 (N_30463,N_23778,N_20129);
nand U30464 (N_30464,N_25210,N_25472);
or U30465 (N_30465,N_26656,N_22759);
and U30466 (N_30466,N_29824,N_24073);
nand U30467 (N_30467,N_24697,N_27505);
xor U30468 (N_30468,N_25551,N_22619);
and U30469 (N_30469,N_28929,N_24138);
nor U30470 (N_30470,N_27936,N_21276);
and U30471 (N_30471,N_28903,N_25032);
nor U30472 (N_30472,N_20313,N_29041);
xnor U30473 (N_30473,N_24836,N_28339);
xnor U30474 (N_30474,N_25052,N_24660);
nor U30475 (N_30475,N_28058,N_25908);
nor U30476 (N_30476,N_27898,N_28315);
xor U30477 (N_30477,N_20795,N_20252);
xnor U30478 (N_30478,N_22597,N_28861);
or U30479 (N_30479,N_26966,N_20959);
nor U30480 (N_30480,N_27067,N_28471);
and U30481 (N_30481,N_24090,N_23482);
nand U30482 (N_30482,N_29079,N_21669);
and U30483 (N_30483,N_29694,N_24229);
or U30484 (N_30484,N_21636,N_26597);
nand U30485 (N_30485,N_20061,N_26547);
xnor U30486 (N_30486,N_20155,N_24342);
and U30487 (N_30487,N_23079,N_25362);
nor U30488 (N_30488,N_22893,N_29850);
or U30489 (N_30489,N_27517,N_26017);
xor U30490 (N_30490,N_20889,N_25994);
xor U30491 (N_30491,N_22631,N_20375);
nor U30492 (N_30492,N_23227,N_29387);
xnor U30493 (N_30493,N_27473,N_20351);
nor U30494 (N_30494,N_28671,N_26083);
nor U30495 (N_30495,N_29320,N_26646);
or U30496 (N_30496,N_20450,N_24234);
nor U30497 (N_30497,N_21843,N_29124);
nand U30498 (N_30498,N_21971,N_24321);
nor U30499 (N_30499,N_29744,N_20662);
xnor U30500 (N_30500,N_25486,N_20211);
and U30501 (N_30501,N_23928,N_25110);
xnor U30502 (N_30502,N_25605,N_23409);
or U30503 (N_30503,N_26103,N_21064);
or U30504 (N_30504,N_25106,N_20683);
or U30505 (N_30505,N_28747,N_20886);
nor U30506 (N_30506,N_29708,N_23567);
xnor U30507 (N_30507,N_29881,N_21681);
nand U30508 (N_30508,N_26850,N_23130);
or U30509 (N_30509,N_29179,N_27909);
xnor U30510 (N_30510,N_26321,N_28748);
xor U30511 (N_30511,N_27764,N_28513);
nand U30512 (N_30512,N_24650,N_20587);
nor U30513 (N_30513,N_26488,N_27464);
xnor U30514 (N_30514,N_23340,N_29530);
and U30515 (N_30515,N_23865,N_29131);
nand U30516 (N_30516,N_25914,N_27637);
or U30517 (N_30517,N_24434,N_29572);
nor U30518 (N_30518,N_27823,N_23165);
and U30519 (N_30519,N_20300,N_27241);
and U30520 (N_30520,N_23002,N_21476);
nand U30521 (N_30521,N_27016,N_28826);
nor U30522 (N_30522,N_22422,N_20681);
xnor U30523 (N_30523,N_22796,N_24230);
nor U30524 (N_30524,N_23520,N_21141);
and U30525 (N_30525,N_24791,N_29779);
nor U30526 (N_30526,N_27390,N_20526);
xor U30527 (N_30527,N_28523,N_25001);
nor U30528 (N_30528,N_22962,N_21291);
and U30529 (N_30529,N_22115,N_22282);
nor U30530 (N_30530,N_26609,N_23648);
or U30531 (N_30531,N_27989,N_25340);
nand U30532 (N_30532,N_26524,N_22956);
xnor U30533 (N_30533,N_28049,N_20978);
and U30534 (N_30534,N_23795,N_21946);
xor U30535 (N_30535,N_21480,N_27461);
and U30536 (N_30536,N_27443,N_24532);
and U30537 (N_30537,N_26170,N_28475);
xor U30538 (N_30538,N_22497,N_25366);
nor U30539 (N_30539,N_26295,N_21615);
xnor U30540 (N_30540,N_22338,N_23756);
nand U30541 (N_30541,N_24005,N_21553);
or U30542 (N_30542,N_29686,N_25113);
xor U30543 (N_30543,N_23031,N_22810);
nand U30544 (N_30544,N_21223,N_20204);
nor U30545 (N_30545,N_21437,N_29855);
xor U30546 (N_30546,N_26314,N_24023);
or U30547 (N_30547,N_22090,N_23670);
or U30548 (N_30548,N_26679,N_27667);
or U30549 (N_30549,N_26589,N_21586);
nand U30550 (N_30550,N_28050,N_20257);
nand U30551 (N_30551,N_28687,N_21352);
nand U30552 (N_30552,N_22636,N_21974);
and U30553 (N_30553,N_25005,N_20049);
nand U30554 (N_30554,N_22849,N_20931);
xor U30555 (N_30555,N_25099,N_26635);
or U30556 (N_30556,N_26446,N_28742);
or U30557 (N_30557,N_25053,N_27170);
or U30558 (N_30558,N_22356,N_22698);
and U30559 (N_30559,N_25769,N_27416);
xor U30560 (N_30560,N_28675,N_20392);
or U30561 (N_30561,N_20571,N_22660);
or U30562 (N_30562,N_27873,N_24510);
or U30563 (N_30563,N_28919,N_29447);
and U30564 (N_30564,N_21609,N_25172);
or U30565 (N_30565,N_21820,N_28376);
nand U30566 (N_30566,N_26918,N_27314);
nand U30567 (N_30567,N_27153,N_24495);
nor U30568 (N_30568,N_22049,N_26380);
or U30569 (N_30569,N_29274,N_26697);
and U30570 (N_30570,N_21584,N_24994);
nand U30571 (N_30571,N_25326,N_21097);
nand U30572 (N_30572,N_22362,N_22574);
and U30573 (N_30573,N_20920,N_24348);
nor U30574 (N_30574,N_29188,N_26250);
nor U30575 (N_30575,N_25754,N_20251);
and U30576 (N_30576,N_26665,N_24508);
and U30577 (N_30577,N_28579,N_28864);
nor U30578 (N_30578,N_29430,N_29162);
xor U30579 (N_30579,N_23474,N_25358);
xor U30580 (N_30580,N_23962,N_28904);
or U30581 (N_30581,N_29268,N_25923);
nand U30582 (N_30582,N_27982,N_21581);
nand U30583 (N_30583,N_29739,N_22232);
and U30584 (N_30584,N_22924,N_27556);
or U30585 (N_30585,N_26411,N_23877);
nor U30586 (N_30586,N_24100,N_29471);
nand U30587 (N_30587,N_22598,N_21044);
and U30588 (N_30588,N_26897,N_21833);
nand U30589 (N_30589,N_27620,N_28996);
nand U30590 (N_30590,N_24825,N_27176);
nand U30591 (N_30591,N_20669,N_20817);
or U30592 (N_30592,N_29329,N_26794);
nand U30593 (N_30593,N_28705,N_20218);
and U30594 (N_30594,N_29327,N_26049);
or U30595 (N_30595,N_27085,N_23571);
nor U30596 (N_30596,N_26016,N_24960);
or U30597 (N_30597,N_23242,N_29654);
nor U30598 (N_30598,N_27281,N_27997);
nor U30599 (N_30599,N_28567,N_23701);
and U30600 (N_30600,N_21535,N_26151);
nor U30601 (N_30601,N_26830,N_29877);
nor U30602 (N_30602,N_20027,N_20919);
nor U30603 (N_30603,N_21738,N_21921);
nand U30604 (N_30604,N_22974,N_22643);
nand U30605 (N_30605,N_23923,N_23551);
nor U30606 (N_30606,N_22139,N_20295);
nor U30607 (N_30607,N_29157,N_20021);
xnor U30608 (N_30608,N_27481,N_24915);
xnor U30609 (N_30609,N_22020,N_28164);
nand U30610 (N_30610,N_26726,N_22470);
xor U30611 (N_30611,N_20511,N_27867);
xor U30612 (N_30612,N_27850,N_25414);
or U30613 (N_30613,N_26499,N_23154);
nand U30614 (N_30614,N_25262,N_22246);
xnor U30615 (N_30615,N_22148,N_29535);
nand U30616 (N_30616,N_25012,N_26025);
xnor U30617 (N_30617,N_20685,N_29176);
nand U30618 (N_30618,N_22044,N_26419);
xnor U30619 (N_30619,N_27471,N_21536);
or U30620 (N_30620,N_24727,N_24284);
nor U30621 (N_30621,N_23698,N_22211);
and U30622 (N_30622,N_27213,N_21579);
nand U30623 (N_30623,N_21452,N_26903);
nand U30624 (N_30624,N_23103,N_20140);
nor U30625 (N_30625,N_20580,N_24696);
nand U30626 (N_30626,N_25020,N_25094);
nor U30627 (N_30627,N_23721,N_29864);
nor U30628 (N_30628,N_26459,N_26620);
nor U30629 (N_30629,N_26142,N_22324);
and U30630 (N_30630,N_28515,N_23309);
xor U30631 (N_30631,N_20169,N_29711);
or U30632 (N_30632,N_27357,N_23927);
or U30633 (N_30633,N_25940,N_25826);
and U30634 (N_30634,N_29407,N_27924);
or U30635 (N_30635,N_26073,N_27149);
or U30636 (N_30636,N_24491,N_26407);
or U30637 (N_30637,N_23677,N_20101);
nand U30638 (N_30638,N_23972,N_29050);
and U30639 (N_30639,N_27190,N_25039);
nand U30640 (N_30640,N_27580,N_20095);
xnor U30641 (N_30641,N_27027,N_20772);
nand U30642 (N_30642,N_20282,N_22190);
nand U30643 (N_30643,N_25250,N_28824);
and U30644 (N_30644,N_23213,N_20556);
and U30645 (N_30645,N_23281,N_25228);
xnor U30646 (N_30646,N_22518,N_29345);
nand U30647 (N_30647,N_26762,N_28322);
or U30648 (N_30648,N_24512,N_24428);
nor U30649 (N_30649,N_24089,N_28511);
or U30650 (N_30650,N_25121,N_23887);
nand U30651 (N_30651,N_21931,N_29273);
nand U30652 (N_30652,N_22207,N_20743);
nor U30653 (N_30653,N_29210,N_22707);
nand U30654 (N_30654,N_26463,N_25302);
nor U30655 (N_30655,N_28920,N_24885);
or U30656 (N_30656,N_21322,N_29497);
xnor U30657 (N_30657,N_29443,N_29795);
xnor U30658 (N_30658,N_28429,N_23808);
nand U30659 (N_30659,N_26778,N_22772);
and U30660 (N_30660,N_22285,N_24544);
nor U30661 (N_30661,N_21504,N_20791);
and U30662 (N_30662,N_27433,N_23494);
or U30663 (N_30663,N_21848,N_26386);
nor U30664 (N_30664,N_25018,N_26716);
or U30665 (N_30665,N_26246,N_23337);
nor U30666 (N_30666,N_26453,N_25438);
nand U30667 (N_30667,N_23273,N_24658);
or U30668 (N_30668,N_25212,N_21057);
nor U30669 (N_30669,N_26481,N_28103);
or U30670 (N_30670,N_28487,N_29172);
and U30671 (N_30671,N_29767,N_27290);
nor U30672 (N_30672,N_21728,N_25984);
and U30673 (N_30673,N_23936,N_21719);
nor U30674 (N_30674,N_24983,N_28044);
and U30675 (N_30675,N_23385,N_27278);
or U30676 (N_30676,N_21862,N_23138);
nor U30677 (N_30677,N_27466,N_23847);
nor U30678 (N_30678,N_29586,N_24035);
and U30679 (N_30679,N_20404,N_27447);
nor U30680 (N_30680,N_26688,N_29189);
or U30681 (N_30681,N_22840,N_23051);
or U30682 (N_30682,N_23993,N_24668);
nor U30683 (N_30683,N_23296,N_26086);
nand U30684 (N_30684,N_23107,N_24904);
xnor U30685 (N_30685,N_29026,N_25834);
nand U30686 (N_30686,N_21360,N_23584);
xnor U30687 (N_30687,N_25783,N_25995);
or U30688 (N_30688,N_26826,N_29355);
or U30689 (N_30689,N_25827,N_23413);
or U30690 (N_30690,N_29437,N_20043);
and U30691 (N_30691,N_26282,N_22746);
xor U30692 (N_30692,N_24203,N_29840);
and U30693 (N_30693,N_20500,N_26953);
and U30694 (N_30694,N_28473,N_29940);
or U30695 (N_30695,N_27236,N_21783);
or U30696 (N_30696,N_26333,N_26008);
xor U30697 (N_30697,N_29888,N_24134);
and U30698 (N_30698,N_22798,N_29044);
nor U30699 (N_30699,N_26294,N_28719);
xnor U30700 (N_30700,N_23817,N_23232);
or U30701 (N_30701,N_20494,N_27366);
or U30702 (N_30702,N_20946,N_23076);
or U30703 (N_30703,N_20059,N_24129);
nand U30704 (N_30704,N_23090,N_27407);
nor U30705 (N_30705,N_24445,N_25163);
or U30706 (N_30706,N_24880,N_24145);
and U30707 (N_30707,N_23466,N_22752);
nor U30708 (N_30708,N_20867,N_29063);
nor U30709 (N_30709,N_24404,N_24785);
nand U30710 (N_30710,N_27289,N_27923);
xnor U30711 (N_30711,N_21817,N_22846);
nand U30712 (N_30712,N_25768,N_20371);
or U30713 (N_30713,N_20629,N_27364);
and U30714 (N_30714,N_28257,N_20007);
nand U30715 (N_30715,N_27423,N_20121);
or U30716 (N_30716,N_27194,N_21838);
nor U30717 (N_30717,N_27550,N_25980);
nor U30718 (N_30718,N_26373,N_26237);
and U30719 (N_30719,N_21105,N_27626);
or U30720 (N_30720,N_27090,N_20266);
nand U30721 (N_30721,N_27049,N_22820);
nor U30722 (N_30722,N_26664,N_22228);
nand U30723 (N_30723,N_27742,N_29303);
and U30724 (N_30724,N_20528,N_22194);
nand U30725 (N_30725,N_29607,N_28759);
nor U30726 (N_30726,N_21424,N_26771);
or U30727 (N_30727,N_21549,N_25558);
nor U30728 (N_30728,N_21940,N_27507);
xor U30729 (N_30729,N_28901,N_27427);
nand U30730 (N_30730,N_29762,N_28583);
nand U30731 (N_30731,N_21633,N_28332);
nand U30732 (N_30732,N_20917,N_28739);
nand U30733 (N_30733,N_28944,N_28977);
nor U30734 (N_30734,N_24015,N_29259);
and U30735 (N_30735,N_22498,N_20701);
nor U30736 (N_30736,N_23797,N_22699);
nor U30737 (N_30737,N_26532,N_23085);
xnor U30738 (N_30738,N_28668,N_20794);
nand U30739 (N_30739,N_27394,N_25197);
or U30740 (N_30740,N_23379,N_28278);
or U30741 (N_30741,N_20876,N_25698);
nand U30742 (N_30742,N_22331,N_23011);
xnor U30743 (N_30743,N_22312,N_21502);
nand U30744 (N_30744,N_26458,N_24277);
nor U30745 (N_30745,N_22326,N_24078);
xnor U30746 (N_30746,N_28466,N_29331);
nor U30747 (N_30747,N_29165,N_28018);
xor U30748 (N_30748,N_29482,N_21413);
or U30749 (N_30749,N_21713,N_22953);
nand U30750 (N_30750,N_22405,N_20008);
or U30751 (N_30751,N_22136,N_21753);
and U30752 (N_30752,N_24924,N_27954);
or U30753 (N_30753,N_23505,N_27738);
and U30754 (N_30754,N_27540,N_26818);
nand U30755 (N_30755,N_25128,N_29883);
nand U30756 (N_30756,N_26938,N_22640);
nor U30757 (N_30757,N_24692,N_21319);
nand U30758 (N_30758,N_26356,N_22484);
nand U30759 (N_30759,N_23822,N_29684);
or U30760 (N_30760,N_22365,N_27301);
or U30761 (N_30761,N_23256,N_27188);
or U30762 (N_30762,N_25215,N_25359);
and U30763 (N_30763,N_26667,N_29683);
nand U30764 (N_30764,N_20975,N_22147);
or U30765 (N_30765,N_20127,N_23472);
xor U30766 (N_30766,N_28788,N_26530);
or U30767 (N_30767,N_28638,N_29700);
nor U30768 (N_30768,N_26320,N_26736);
nand U30769 (N_30769,N_29701,N_23224);
nand U30770 (N_30770,N_21780,N_20449);
nor U30771 (N_30771,N_27605,N_25777);
nand U30772 (N_30772,N_20719,N_27838);
or U30773 (N_30773,N_21813,N_28007);
nand U30774 (N_30774,N_20200,N_23850);
nand U30775 (N_30775,N_21109,N_26414);
nand U30776 (N_30776,N_26094,N_22758);
nand U30777 (N_30777,N_27575,N_28195);
nor U30778 (N_30778,N_28623,N_29389);
or U30779 (N_30779,N_29875,N_28255);
nand U30780 (N_30780,N_28472,N_29218);
nand U30781 (N_30781,N_26355,N_21449);
or U30782 (N_30782,N_26451,N_24365);
xnor U30783 (N_30783,N_24682,N_24953);
and U30784 (N_30784,N_23284,N_24384);
xnor U30785 (N_30785,N_27681,N_27920);
or U30786 (N_30786,N_28858,N_23893);
nor U30787 (N_30787,N_24828,N_23044);
and U30788 (N_30788,N_25267,N_24170);
nand U30789 (N_30789,N_27877,N_28776);
and U30790 (N_30790,N_25635,N_27732);
xor U30791 (N_30791,N_27886,N_21124);
or U30792 (N_30792,N_29383,N_20833);
xor U30793 (N_30793,N_25017,N_20439);
xnor U30794 (N_30794,N_22740,N_21296);
nand U30795 (N_30795,N_21656,N_28720);
and U30796 (N_30796,N_21680,N_25481);
or U30797 (N_30797,N_25098,N_24350);
nand U30798 (N_30798,N_29005,N_24142);
or U30799 (N_30799,N_26036,N_29178);
or U30800 (N_30800,N_29442,N_21631);
or U30801 (N_30801,N_25140,N_23113);
or U30802 (N_30802,N_29542,N_23683);
or U30803 (N_30803,N_28576,N_22056);
nor U30804 (N_30804,N_24549,N_23897);
nor U30805 (N_30805,N_29653,N_20780);
nand U30806 (N_30806,N_24807,N_25162);
or U30807 (N_30807,N_21255,N_25061);
or U30808 (N_30808,N_28820,N_21310);
nor U30809 (N_30809,N_22667,N_28359);
and U30810 (N_30810,N_24131,N_20788);
and U30811 (N_30811,N_21755,N_20892);
and U30812 (N_30812,N_27998,N_20442);
or U30813 (N_30813,N_28156,N_29823);
and U30814 (N_30814,N_26382,N_29213);
xnor U30815 (N_30815,N_29485,N_25387);
xnor U30816 (N_30816,N_26280,N_29483);
nor U30817 (N_30817,N_26523,N_25462);
nand U30818 (N_30818,N_21934,N_22714);
nand U30819 (N_30819,N_27895,N_28244);
and U30820 (N_30820,N_22553,N_28263);
and U30821 (N_30821,N_20991,N_26802);
nand U30822 (N_30822,N_22011,N_22122);
or U30823 (N_30823,N_26370,N_25956);
nor U30824 (N_30824,N_24750,N_24257);
nand U30825 (N_30825,N_24109,N_29229);
xor U30826 (N_30826,N_28633,N_29109);
nor U30827 (N_30827,N_27216,N_28841);
or U30828 (N_30828,N_27034,N_22958);
xor U30829 (N_30829,N_26271,N_21621);
or U30830 (N_30830,N_28067,N_24212);
and U30831 (N_30831,N_23813,N_23387);
and U30832 (N_30832,N_22371,N_24699);
or U30833 (N_30833,N_27468,N_29263);
nor U30834 (N_30834,N_29281,N_22217);
nand U30835 (N_30835,N_26819,N_20321);
xor U30836 (N_30836,N_20533,N_20615);
nor U30837 (N_30837,N_22048,N_20544);
nor U30838 (N_30838,N_26628,N_25973);
or U30839 (N_30839,N_29677,N_24842);
nor U30840 (N_30840,N_23384,N_25178);
xor U30841 (N_30841,N_23070,N_22569);
or U30842 (N_30842,N_21893,N_26484);
and U30843 (N_30843,N_20136,N_26674);
nand U30844 (N_30844,N_27455,N_23700);
nand U30845 (N_30845,N_24780,N_29086);
and U30846 (N_30846,N_25580,N_26081);
or U30847 (N_30847,N_27124,N_22679);
nor U30848 (N_30848,N_24624,N_28275);
xor U30849 (N_30849,N_21367,N_22717);
or U30850 (N_30850,N_28283,N_22548);
or U30851 (N_30851,N_29458,N_22367);
xor U30852 (N_30852,N_28834,N_24181);
nor U30853 (N_30853,N_22389,N_24482);
nor U30854 (N_30854,N_28343,N_21686);
and U30855 (N_30855,N_28037,N_28760);
xnor U30856 (N_30856,N_21159,N_28972);
and U30857 (N_30857,N_29040,N_23336);
or U30858 (N_30858,N_29045,N_28503);
xor U30859 (N_30859,N_22742,N_23006);
nand U30860 (N_30860,N_24366,N_25800);
nor U30861 (N_30861,N_28569,N_26392);
and U30862 (N_30862,N_24686,N_26095);
xnor U30863 (N_30863,N_20888,N_26058);
and U30864 (N_30864,N_23828,N_22304);
and U30865 (N_30865,N_25744,N_29928);
xor U30866 (N_30866,N_24390,N_27220);
or U30867 (N_30867,N_20322,N_24330);
and U30868 (N_30868,N_23094,N_24399);
nand U30869 (N_30869,N_27254,N_22345);
nor U30870 (N_30870,N_27653,N_22247);
nand U30871 (N_30871,N_22108,N_28481);
nand U30872 (N_30872,N_23602,N_20011);
and U30873 (N_30873,N_29538,N_23607);
xnor U30874 (N_30874,N_24882,N_28033);
nand U30875 (N_30875,N_24831,N_24260);
and U30876 (N_30876,N_28970,N_21503);
and U30877 (N_30877,N_21678,N_28430);
and U30878 (N_30878,N_25043,N_20871);
or U30879 (N_30879,N_27494,N_25581);
xnor U30880 (N_30880,N_22449,N_29074);
nor U30881 (N_30881,N_27885,N_22804);
and U30882 (N_30882,N_25046,N_28422);
nand U30883 (N_30883,N_20648,N_23761);
nand U30884 (N_30884,N_26413,N_26686);
xnor U30885 (N_30885,N_20997,N_25871);
nand U30886 (N_30886,N_23124,N_27795);
xnor U30887 (N_30887,N_22573,N_22838);
or U30888 (N_30888,N_23978,N_29341);
and U30889 (N_30889,N_21287,N_24091);
or U30890 (N_30890,N_20480,N_25196);
nor U30891 (N_30891,N_24313,N_27995);
nand U30892 (N_30892,N_22243,N_24616);
or U30893 (N_30893,N_21485,N_24652);
or U30894 (N_30894,N_22875,N_29539);
xnor U30895 (N_30895,N_20004,N_23010);
and U30896 (N_30896,N_20289,N_23020);
or U30897 (N_30897,N_22676,N_21278);
xor U30898 (N_30898,N_22728,N_24865);
and U30899 (N_30899,N_22220,N_29834);
nand U30900 (N_30900,N_23915,N_26457);
nor U30901 (N_30901,N_21202,N_28251);
nor U30902 (N_30902,N_20883,N_22039);
or U30903 (N_30903,N_25095,N_26470);
and U30904 (N_30904,N_28801,N_29749);
nor U30905 (N_30905,N_22596,N_23319);
nor U30906 (N_30906,N_27837,N_26269);
nor U30907 (N_30907,N_26087,N_25488);
nor U30908 (N_30908,N_21361,N_20482);
or U30909 (N_30909,N_25024,N_20022);
and U30910 (N_30910,N_23779,N_26445);
nand U30911 (N_30911,N_22092,N_25875);
xnor U30912 (N_30912,N_29448,N_29087);
nand U30913 (N_30913,N_24781,N_21041);
nand U30914 (N_30914,N_27480,N_27104);
xnor U30915 (N_30915,N_20812,N_29101);
nand U30916 (N_30916,N_24009,N_22157);
or U30917 (N_30917,N_27117,N_25755);
and U30918 (N_30918,N_23854,N_29104);
nand U30919 (N_30919,N_20398,N_29166);
xnor U30920 (N_30920,N_27865,N_20602);
or U30921 (N_30921,N_25133,N_29761);
and U30922 (N_30922,N_24566,N_24757);
nor U30923 (N_30923,N_25960,N_25181);
or U30924 (N_30924,N_29462,N_23290);
or U30925 (N_30925,N_22854,N_24834);
or U30926 (N_30926,N_27472,N_24784);
or U30927 (N_30927,N_26085,N_24250);
nand U30928 (N_30928,N_27313,N_28757);
nor U30929 (N_30929,N_29862,N_27387);
and U30930 (N_30930,N_24908,N_22076);
nand U30931 (N_30931,N_24143,N_26652);
or U30932 (N_30932,N_23206,N_23492);
nand U30933 (N_30933,N_27428,N_27264);
nor U30934 (N_30934,N_27560,N_28350);
xnor U30935 (N_30935,N_24322,N_27648);
nand U30936 (N_30936,N_20640,N_24779);
or U30937 (N_30937,N_27043,N_23964);
and U30938 (N_30938,N_25388,N_24628);
and U30939 (N_30939,N_21093,N_24739);
nor U30940 (N_30940,N_28869,N_25469);
xor U30941 (N_30941,N_22514,N_22421);
or U30942 (N_30942,N_26615,N_27434);
or U30943 (N_30943,N_28937,N_25982);
or U30944 (N_30944,N_22380,N_20560);
or U30945 (N_30945,N_20326,N_21685);
xnor U30946 (N_30946,N_21075,N_28562);
nand U30947 (N_30947,N_21643,N_29143);
nand U30948 (N_30948,N_22753,N_25666);
nor U30949 (N_30949,N_27450,N_21375);
nand U30950 (N_30950,N_20388,N_24396);
and U30951 (N_30951,N_23931,N_25346);
and U30952 (N_30952,N_21303,N_21939);
and U30953 (N_30953,N_26935,N_26673);
and U30954 (N_30954,N_29186,N_23125);
or U30955 (N_30955,N_23381,N_27816);
xnor U30956 (N_30956,N_27689,N_22830);
nand U30957 (N_30957,N_29296,N_24443);
and U30958 (N_30958,N_24165,N_25409);
nand U30959 (N_30959,N_24081,N_26060);
xor U30960 (N_30960,N_22889,N_24409);
nand U30961 (N_30961,N_21145,N_21407);
nor U30962 (N_30962,N_23736,N_23183);
or U30963 (N_30963,N_22434,N_29975);
nor U30964 (N_30964,N_24336,N_26586);
or U30965 (N_30965,N_23753,N_26432);
and U30966 (N_30966,N_29947,N_23933);
or U30967 (N_30967,N_20349,N_25139);
and U30968 (N_30968,N_21611,N_20347);
or U30969 (N_30969,N_24190,N_23842);
nor U30970 (N_30970,N_27368,N_24282);
and U30971 (N_30971,N_26313,N_26517);
nor U30972 (N_30972,N_21198,N_23692);
or U30973 (N_30973,N_20691,N_20031);
or U30974 (N_30974,N_20284,N_26364);
nand U30975 (N_30975,N_22146,N_23123);
and U30976 (N_30976,N_21456,N_27076);
nand U30977 (N_30977,N_28495,N_24619);
xnor U30978 (N_30978,N_24280,N_27852);
and U30979 (N_30979,N_21923,N_23241);
and U30980 (N_30980,N_23960,N_23711);
and U30981 (N_30981,N_29060,N_25013);
nand U30982 (N_30982,N_22341,N_24388);
nor U30983 (N_30983,N_23816,N_21998);
xor U30984 (N_30984,N_27948,N_28426);
nand U30985 (N_30985,N_26761,N_21808);
xnor U30986 (N_30986,N_28289,N_23055);
or U30987 (N_30987,N_26759,N_25779);
xor U30988 (N_30988,N_29811,N_28366);
and U30989 (N_30989,N_28146,N_25748);
nor U30990 (N_30990,N_28674,N_23840);
or U30991 (N_30991,N_25729,N_27788);
xnor U30992 (N_30992,N_29175,N_26682);
nand U30993 (N_30993,N_28336,N_25712);
and U30994 (N_30994,N_21389,N_23531);
xnor U30995 (N_30995,N_28435,N_29860);
nor U30996 (N_30996,N_28771,N_24337);
and U30997 (N_30997,N_23791,N_27736);
xnor U30998 (N_30998,N_27296,N_28536);
and U30999 (N_30999,N_28127,N_28588);
and U31000 (N_31000,N_23033,N_24262);
and U31001 (N_31001,N_21915,N_26276);
or U31002 (N_31002,N_21812,N_27052);
xor U31003 (N_31003,N_25725,N_23432);
or U31004 (N_31004,N_24984,N_23074);
nor U31005 (N_31005,N_29140,N_22175);
nand U31006 (N_31006,N_21696,N_25717);
nand U31007 (N_31007,N_23643,N_21725);
or U31008 (N_31008,N_25125,N_23529);
nor U31009 (N_31009,N_20083,N_21714);
nand U31010 (N_31010,N_22129,N_27883);
nor U31011 (N_31011,N_28221,N_21932);
nand U31012 (N_31012,N_26297,N_22868);
nor U31013 (N_31013,N_22516,N_29237);
nand U31014 (N_31014,N_20148,N_28584);
nand U31015 (N_31015,N_28219,N_24621);
or U31016 (N_31016,N_28627,N_29511);
xor U31017 (N_31017,N_21984,N_29789);
nor U31018 (N_31018,N_27813,N_22017);
or U31019 (N_31019,N_21516,N_28928);
and U31020 (N_31020,N_26172,N_27664);
xor U31021 (N_31021,N_26752,N_20197);
nand U31022 (N_31022,N_27251,N_26512);
xor U31023 (N_31023,N_29516,N_22021);
nand U31024 (N_31024,N_20183,N_22851);
and U31025 (N_31025,N_23347,N_28922);
nor U31026 (N_31026,N_27672,N_22673);
or U31027 (N_31027,N_25763,N_26218);
and U31028 (N_31028,N_23203,N_20895);
nand U31029 (N_31029,N_27984,N_23092);
xnor U31030 (N_31030,N_28334,N_21085);
xnor U31031 (N_31031,N_20176,N_20203);
or U31032 (N_31032,N_27411,N_23640);
nand U31033 (N_31033,N_20224,N_25810);
nand U31034 (N_31034,N_20039,N_25693);
and U31035 (N_31035,N_27787,N_20564);
nand U31036 (N_31036,N_29495,N_21094);
xnor U31037 (N_31037,N_28987,N_23560);
or U31038 (N_31038,N_20921,N_21684);
xnor U31039 (N_31039,N_27633,N_28385);
or U31040 (N_31040,N_20850,N_29573);
xor U31041 (N_31041,N_29512,N_22034);
and U31042 (N_31042,N_26377,N_23561);
or U31043 (N_31043,N_29164,N_21889);
or U31044 (N_31044,N_25368,N_24525);
and U31045 (N_31045,N_20259,N_28038);
nor U31046 (N_31046,N_29576,N_26741);
nand U31047 (N_31047,N_26015,N_28440);
or U31048 (N_31048,N_26636,N_22603);
and U31049 (N_31049,N_23799,N_29228);
nor U31050 (N_31050,N_25583,N_25516);
and U31051 (N_31051,N_23047,N_26997);
xnor U31052 (N_31052,N_28666,N_27491);
nor U31053 (N_31053,N_28911,N_20464);
xor U31054 (N_31054,N_21969,N_29199);
or U31055 (N_31055,N_20457,N_20341);
xor U31056 (N_31056,N_29069,N_22164);
or U31057 (N_31057,N_26833,N_28199);
or U31058 (N_31058,N_24191,N_25727);
and U31059 (N_31059,N_28467,N_29897);
or U31060 (N_31060,N_23246,N_20963);
or U31061 (N_31061,N_20458,N_29047);
nand U31062 (N_31062,N_24539,N_26948);
and U31063 (N_31063,N_26398,N_21559);
or U31064 (N_31064,N_28974,N_23771);
nand U31065 (N_31065,N_26035,N_24029);
nand U31066 (N_31066,N_23226,N_25269);
nor U31067 (N_31067,N_27977,N_24483);
nand U31068 (N_31068,N_24829,N_21879);
or U31069 (N_31069,N_22289,N_26135);
xnor U31070 (N_31070,N_20834,N_27554);
nor U31071 (N_31071,N_29464,N_23666);
and U31072 (N_31072,N_22711,N_22308);
nor U31073 (N_31073,N_27935,N_29334);
or U31074 (N_31074,N_29721,N_21630);
nand U31075 (N_31075,N_23524,N_20944);
xor U31076 (N_31076,N_22474,N_29513);
or U31077 (N_31077,N_25759,N_29358);
or U31078 (N_31078,N_20470,N_22604);
or U31079 (N_31079,N_22033,N_24479);
nand U31080 (N_31080,N_26118,N_22957);
nor U31081 (N_31081,N_20784,N_27396);
xor U31082 (N_31082,N_29111,N_21732);
xnor U31083 (N_31083,N_28517,N_21116);
or U31084 (N_31084,N_20708,N_29367);
or U31085 (N_31085,N_27144,N_28214);
and U31086 (N_31086,N_26012,N_26542);
xnor U31087 (N_31087,N_29651,N_21800);
or U31088 (N_31088,N_20925,N_25624);
or U31089 (N_31089,N_23231,N_27824);
xor U31090 (N_31090,N_29392,N_23414);
xor U31091 (N_31091,N_24218,N_22760);
and U31092 (N_31092,N_29845,N_23039);
or U31093 (N_31093,N_29764,N_29898);
nor U31094 (N_31094,N_25597,N_21212);
or U31095 (N_31095,N_21397,N_23576);
nand U31096 (N_31096,N_21152,N_28012);
nand U31097 (N_31097,N_28642,N_29467);
nand U31098 (N_31098,N_25413,N_21261);
nor U31099 (N_31099,N_21155,N_29153);
and U31100 (N_31100,N_20831,N_28486);
xor U31101 (N_31101,N_29382,N_24847);
and U31102 (N_31102,N_20217,N_25246);
nand U31103 (N_31103,N_22652,N_26866);
nand U31104 (N_31104,N_29934,N_21949);
and U31105 (N_31105,N_28157,N_23614);
xnor U31106 (N_31106,N_21274,N_20508);
and U31107 (N_31107,N_25854,N_27501);
nand U31108 (N_31108,N_27200,N_28992);
and U31109 (N_31109,N_23869,N_27009);
nand U31110 (N_31110,N_27968,N_22204);
xor U31111 (N_31111,N_26622,N_24069);
and U31112 (N_31112,N_22431,N_23653);
and U31113 (N_31113,N_22042,N_24654);
nor U31114 (N_31114,N_28042,N_29690);
or U31115 (N_31115,N_22590,N_29649);
nand U31116 (N_31116,N_26471,N_26068);
or U31117 (N_31117,N_20797,N_29525);
or U31118 (N_31118,N_27361,N_24475);
and U31119 (N_31119,N_28491,N_27881);
xor U31120 (N_31120,N_22417,N_24006);
or U31121 (N_31121,N_25650,N_29541);
and U31122 (N_31122,N_21439,N_27068);
nor U31123 (N_31123,N_20355,N_26490);
xor U31124 (N_31124,N_29342,N_20220);
and U31125 (N_31125,N_21727,N_22457);
nor U31126 (N_31126,N_27731,N_27389);
nor U31127 (N_31127,N_27342,N_20524);
or U31128 (N_31128,N_28641,N_24592);
or U31129 (N_31129,N_28230,N_25191);
nor U31130 (N_31130,N_20847,N_22199);
or U31131 (N_31131,N_24900,N_20694);
xnor U31132 (N_31132,N_23196,N_22052);
nor U31133 (N_31133,N_28787,N_29987);
xor U31134 (N_31134,N_26384,N_27209);
or U31135 (N_31135,N_20365,N_28862);
xor U31136 (N_31136,N_22954,N_25253);
nor U31137 (N_31137,N_26381,N_21994);
nand U31138 (N_31138,N_24793,N_20288);
or U31139 (N_31139,N_20599,N_22561);
nor U31140 (N_31140,N_22778,N_22240);
or U31141 (N_31141,N_28085,N_26226);
and U31142 (N_31142,N_28993,N_29699);
or U31143 (N_31143,N_20611,N_28953);
and U31144 (N_31144,N_24171,N_23316);
and U31145 (N_31145,N_20382,N_21767);
or U31146 (N_31146,N_28003,N_24347);
and U31147 (N_31147,N_28288,N_25318);
nor U31148 (N_31148,N_23356,N_23827);
nand U31149 (N_31149,N_25109,N_26780);
or U31150 (N_31150,N_21920,N_23814);
nor U31151 (N_31151,N_25171,N_25386);
or U31152 (N_31152,N_22113,N_23804);
xor U31153 (N_31153,N_25182,N_21604);
xnor U31154 (N_31154,N_24163,N_22419);
or U31155 (N_31155,N_21135,N_20652);
and U31156 (N_31156,N_20885,N_28379);
nor U31157 (N_31157,N_22468,N_23781);
xnor U31158 (N_31158,N_28403,N_25216);
nand U31159 (N_31159,N_21806,N_24436);
nor U31160 (N_31160,N_20984,N_21861);
or U31161 (N_31161,N_29846,N_28036);
and U31162 (N_31162,N_26350,N_26116);
and U31163 (N_31163,N_21564,N_29230);
nand U31164 (N_31164,N_27187,N_29012);
or U31165 (N_31165,N_22930,N_21836);
nand U31166 (N_31166,N_26529,N_27791);
nand U31167 (N_31167,N_20126,N_24615);
nand U31168 (N_31168,N_28749,N_20263);
or U31169 (N_31169,N_29280,N_28644);
or U31170 (N_31170,N_28387,N_25240);
or U31171 (N_31171,N_29903,N_24703);
and U31172 (N_31172,N_24917,N_20809);
nor U31173 (N_31173,N_28293,N_26303);
nor U31174 (N_31174,N_21272,N_21182);
xnor U31175 (N_31175,N_20248,N_23402);
and U31176 (N_31176,N_21794,N_23392);
xnor U31177 (N_31177,N_26947,N_21541);
or U31178 (N_31178,N_21162,N_27993);
nand U31179 (N_31179,N_25890,N_29125);
xor U31180 (N_31180,N_22471,N_20293);
nand U31181 (N_31181,N_23276,N_26361);
and U31182 (N_31182,N_22294,N_22351);
nor U31183 (N_31183,N_22099,N_25798);
or U31184 (N_31184,N_28660,N_22709);
nand U31185 (N_31185,N_23425,N_22125);
nand U31186 (N_31186,N_22466,N_23564);
and U31187 (N_31187,N_27953,N_29061);
or U31188 (N_31188,N_29055,N_26211);
xor U31189 (N_31189,N_27286,N_25814);
nor U31190 (N_31190,N_23752,N_25418);
or U31191 (N_31191,N_22835,N_20111);
nand U31192 (N_31192,N_25509,N_26216);
nand U31193 (N_31193,N_20114,N_28148);
and U31194 (N_31194,N_28958,N_26607);
nand U31195 (N_31195,N_25119,N_21708);
and U31196 (N_31196,N_22030,N_23061);
or U31197 (N_31197,N_22098,N_26127);
nand U31198 (N_31198,N_24246,N_21157);
xor U31199 (N_31199,N_21784,N_22657);
or U31200 (N_31200,N_23058,N_25522);
xnor U31201 (N_31201,N_24968,N_27448);
nor U31202 (N_31202,N_24642,N_27864);
or U31203 (N_31203,N_26957,N_29899);
or U31204 (N_31204,N_27148,N_25699);
nand U31205 (N_31205,N_27687,N_28064);
or U31206 (N_31206,N_27486,N_23453);
or U31207 (N_31207,N_27185,N_26565);
nand U31208 (N_31208,N_21702,N_28646);
xnor U31209 (N_31209,N_23004,N_26109);
nand U31210 (N_31210,N_24896,N_26696);
xnor U31211 (N_31211,N_21207,N_23871);
and U31212 (N_31212,N_20335,N_29550);
and U31213 (N_31213,N_25859,N_27962);
nand U31214 (N_31214,N_27215,N_27015);
xnor U31215 (N_31215,N_24753,N_21351);
and U31216 (N_31216,N_23521,N_29937);
or U31217 (N_31217,N_25188,N_24273);
and U31218 (N_31218,N_26604,N_26669);
or U31219 (N_31219,N_27371,N_27900);
or U31220 (N_31220,N_23475,N_20493);
or U31221 (N_31221,N_22867,N_22981);
or U31222 (N_31222,N_25447,N_25896);
and U31223 (N_31223,N_27944,N_28291);
or U31224 (N_31224,N_22392,N_26020);
xor U31225 (N_31225,N_25985,N_28392);
nor U31226 (N_31226,N_22672,N_23911);
and U31227 (N_31227,N_24184,N_23484);
or U31228 (N_31228,N_24751,N_20085);
and U31229 (N_31229,N_28081,N_20105);
or U31230 (N_31230,N_25652,N_28243);
or U31231 (N_31231,N_29745,N_27520);
and U31232 (N_31232,N_24061,N_20069);
or U31233 (N_31233,N_20246,N_27778);
and U31234 (N_31234,N_27781,N_29094);
nor U31235 (N_31235,N_21880,N_20410);
and U31236 (N_31236,N_29771,N_22340);
and U31237 (N_31237,N_27702,N_27551);
xor U31238 (N_31238,N_28927,N_22483);
or U31239 (N_31239,N_26569,N_24017);
nand U31240 (N_31240,N_27498,N_27806);
xor U31241 (N_31241,N_23550,N_23650);
xnor U31242 (N_31242,N_20934,N_29593);
xor U31243 (N_31243,N_20361,N_26797);
nand U31244 (N_31244,N_28954,N_29821);
nor U31245 (N_31245,N_28634,N_22622);
or U31246 (N_31246,N_29644,N_24198);
and U31247 (N_31247,N_23291,N_23645);
nand U31248 (N_31248,N_22229,N_24946);
xnor U31249 (N_31249,N_21878,N_26755);
or U31250 (N_31250,N_22062,N_26291);
or U31251 (N_31251,N_25743,N_23491);
or U31252 (N_31252,N_27379,N_26403);
and U31253 (N_31253,N_22920,N_21525);
or U31254 (N_31254,N_26014,N_24987);
or U31255 (N_31255,N_26994,N_25491);
nand U31256 (N_31256,N_26308,N_29479);
xor U31257 (N_31257,N_20205,N_25947);
nand U31258 (N_31258,N_27442,N_20250);
and U31259 (N_31259,N_29655,N_25654);
xnor U31260 (N_31260,N_24180,N_21761);
nand U31261 (N_31261,N_20860,N_29025);
xor U31262 (N_31262,N_29585,N_20712);
xor U31263 (N_31263,N_22826,N_23863);
and U31264 (N_31264,N_26779,N_29609);
xnor U31265 (N_31265,N_28716,N_27374);
xor U31266 (N_31266,N_28701,N_25015);
nor U31267 (N_31267,N_27947,N_21729);
or U31268 (N_31268,N_29405,N_21248);
xor U31269 (N_31269,N_20748,N_21873);
or U31270 (N_31270,N_22089,N_26629);
xnor U31271 (N_31271,N_27479,N_22131);
and U31272 (N_31272,N_25036,N_22903);
or U31273 (N_31273,N_22581,N_20868);
and U31274 (N_31274,N_29902,N_28526);
nor U31275 (N_31275,N_25054,N_21750);
xor U31276 (N_31276,N_20765,N_25813);
nor U31277 (N_31277,N_27746,N_26161);
or U31278 (N_31278,N_20655,N_25011);
or U31279 (N_31279,N_22907,N_24723);
nor U31280 (N_31280,N_24528,N_28280);
nor U31281 (N_31281,N_20527,N_26416);
nand U31282 (N_31282,N_20908,N_25175);
nor U31283 (N_31283,N_29036,N_28220);
and U31284 (N_31284,N_21852,N_21395);
and U31285 (N_31285,N_23726,N_28736);
or U31286 (N_31286,N_20459,N_29556);
nor U31287 (N_31287,N_21618,N_20238);
nor U31288 (N_31288,N_28878,N_24541);
xnor U31289 (N_31289,N_27939,N_20116);
nand U31290 (N_31290,N_21172,N_21046);
xnor U31291 (N_31291,N_23064,N_25595);
and U31292 (N_31292,N_23568,N_24086);
or U31293 (N_31293,N_25214,N_27925);
nor U31294 (N_31294,N_20177,N_24974);
or U31295 (N_31295,N_24030,N_27137);
or U31296 (N_31296,N_24824,N_25049);
and U31297 (N_31297,N_20545,N_25428);
nand U31298 (N_31298,N_24507,N_21547);
or U31299 (N_31299,N_24478,N_28872);
nand U31300 (N_31300,N_23424,N_24509);
or U31301 (N_31301,N_28211,N_20423);
nand U31302 (N_31302,N_23463,N_23443);
or U31303 (N_31303,N_22193,N_25401);
nand U31304 (N_31304,N_21316,N_24094);
or U31305 (N_31305,N_29730,N_25411);
xor U31306 (N_31306,N_21506,N_29017);
and U31307 (N_31307,N_24546,N_25230);
and U31308 (N_31308,N_21454,N_21444);
nand U31309 (N_31309,N_29838,N_22547);
nand U31310 (N_31310,N_29215,N_24777);
and U31311 (N_31311,N_20323,N_21558);
nor U31312 (N_31312,N_26089,N_24899);
nand U31313 (N_31313,N_29814,N_22831);
nor U31314 (N_31314,N_22950,N_23672);
nand U31315 (N_31315,N_20491,N_20195);
nand U31316 (N_31316,N_21299,N_20010);
and U31317 (N_31317,N_23394,N_29347);
nand U31318 (N_31318,N_22313,N_28212);
or U31319 (N_31319,N_29072,N_24651);
and U31320 (N_31320,N_21121,N_25614);
nor U31321 (N_31321,N_20913,N_26339);
nor U31322 (N_31322,N_28373,N_23445);
and U31323 (N_31323,N_23388,N_22151);
nor U31324 (N_31324,N_22882,N_27713);
nor U31325 (N_31325,N_24346,N_25452);
nor U31326 (N_31326,N_23940,N_28098);
and U31327 (N_31327,N_23684,N_28807);
or U31328 (N_31328,N_23104,N_23558);
xnor U31329 (N_31329,N_20849,N_23900);
nand U31330 (N_31330,N_27242,N_20698);
or U31331 (N_31331,N_29746,N_28702);
or U31332 (N_31332,N_23685,N_22461);
and U31333 (N_31333,N_25166,N_27237);
xor U31334 (N_31334,N_28573,N_27800);
nand U31335 (N_31335,N_23544,N_24440);
nor U31336 (N_31336,N_23938,N_21482);
and U31337 (N_31337,N_24465,N_25864);
and U31338 (N_31338,N_22593,N_26468);
nor U31339 (N_31339,N_22584,N_29120);
or U31340 (N_31340,N_28294,N_20534);
nand U31341 (N_31341,N_24238,N_28839);
nor U31342 (N_31342,N_23695,N_27753);
nor U31343 (N_31343,N_28506,N_23805);
and U31344 (N_31344,N_28131,N_23193);
nor U31345 (N_31345,N_20446,N_26064);
and U31346 (N_31346,N_26855,N_29961);
nand U31347 (N_31347,N_23539,N_26365);
xor U31348 (N_31348,N_25972,N_27419);
or U31349 (N_31349,N_23792,N_20447);
xor U31350 (N_31350,N_28296,N_22523);
nor U31351 (N_31351,N_23371,N_26344);
and U31352 (N_31352,N_29808,N_21768);
nor U31353 (N_31353,N_26131,N_20757);
or U31354 (N_31354,N_22877,N_25778);
nor U31355 (N_31355,N_27467,N_24770);
xnor U31356 (N_31356,N_22009,N_20146);
or U31357 (N_31357,N_28848,N_21019);
xor U31358 (N_31358,N_26976,N_28271);
nor U31359 (N_31359,N_27555,N_22803);
nor U31360 (N_31360,N_25487,N_24991);
nor U31361 (N_31361,N_28246,N_23983);
or U31362 (N_31362,N_21280,N_21321);
nor U31363 (N_31363,N_27820,N_22695);
xor U31364 (N_31364,N_20555,N_20771);
xor U31365 (N_31365,N_21464,N_21935);
and U31366 (N_31366,N_22541,N_29837);
nand U31367 (N_31367,N_21244,N_21897);
or U31368 (N_31368,N_23258,N_24979);
or U31369 (N_31369,N_23240,N_22669);
nor U31370 (N_31370,N_26592,N_28450);
xor U31371 (N_31371,N_23988,N_23029);
and U31372 (N_31372,N_26706,N_22948);
nand U31373 (N_31373,N_25992,N_21149);
nor U31374 (N_31374,N_21061,N_24221);
and U31375 (N_31375,N_27272,N_29051);
and U31376 (N_31376,N_26631,N_22167);
nand U31377 (N_31377,N_26108,N_21973);
nand U31378 (N_31378,N_20030,N_20633);
or U31379 (N_31379,N_26009,N_28697);
or U31380 (N_31380,N_29361,N_21835);
nand U31381 (N_31381,N_29977,N_20026);
nor U31382 (N_31382,N_21120,N_26582);
and U31383 (N_31383,N_27079,N_23914);
nand U31384 (N_31384,N_20857,N_24802);
nand U31385 (N_31385,N_25675,N_28549);
xnor U31386 (N_31386,N_26205,N_26951);
or U31387 (N_31387,N_28377,N_23950);
or U31388 (N_31388,N_24841,N_22168);
and U31389 (N_31389,N_24803,N_22887);
nand U31390 (N_31390,N_22143,N_29992);
xnor U31391 (N_31391,N_29236,N_28963);
nor U31392 (N_31392,N_29100,N_26072);
nor U31393 (N_31393,N_22677,N_25226);
nor U31394 (N_31394,N_21826,N_26723);
and U31395 (N_31395,N_28730,N_28643);
and U31396 (N_31396,N_22899,N_25753);
nor U31397 (N_31397,N_24274,N_28084);
or U31398 (N_31398,N_25844,N_25802);
xnor U31399 (N_31399,N_28163,N_22788);
nor U31400 (N_31400,N_27519,N_23205);
or U31401 (N_31401,N_21798,N_23717);
and U31402 (N_31402,N_20950,N_24530);
and U31403 (N_31403,N_27729,N_25422);
nor U31404 (N_31404,N_25981,N_22264);
xor U31405 (N_31405,N_23449,N_20413);
nand U31406 (N_31406,N_25425,N_20158);
xor U31407 (N_31407,N_28355,N_29737);
or U31408 (N_31408,N_22731,N_25263);
nor U31409 (N_31409,N_26149,N_25919);
xor U31410 (N_31410,N_20621,N_21859);
and U31411 (N_31411,N_20666,N_20435);
or U31412 (N_31412,N_29852,N_27125);
and U31413 (N_31413,N_20803,N_27307);
nor U31414 (N_31414,N_24160,N_27558);
nand U31415 (N_31415,N_20644,N_25863);
or U31416 (N_31416,N_28451,N_26872);
xor U31417 (N_31417,N_27961,N_22766);
or U31418 (N_31418,N_20070,N_20700);
and U31419 (N_31419,N_27383,N_28605);
nand U31420 (N_31420,N_21718,N_24506);
or U31421 (N_31421,N_22744,N_29391);
or U31422 (N_31422,N_25441,N_20821);
xnor U31423 (N_31423,N_25764,N_24095);
or U31424 (N_31424,N_26113,N_20741);
nand U31425 (N_31425,N_26195,N_27020);
nand U31426 (N_31426,N_22823,N_26786);
nand U31427 (N_31427,N_21841,N_25760);
nor U31428 (N_31428,N_28353,N_21805);
and U31429 (N_31429,N_21877,N_23638);
and U31430 (N_31430,N_24268,N_22651);
nand U31431 (N_31431,N_22037,N_25534);
and U31432 (N_31432,N_29085,N_24056);
xnor U31433 (N_31433,N_23322,N_28202);
or U31434 (N_31434,N_20832,N_29156);
or U31435 (N_31435,N_26133,N_25432);
nand U31436 (N_31436,N_21460,N_28978);
xor U31437 (N_31437,N_20040,N_21074);
and U31438 (N_31438,N_20091,N_27019);
nor U31439 (N_31439,N_20663,N_24394);
and U31440 (N_31440,N_20787,N_24318);
and U31441 (N_31441,N_28274,N_25185);
and U31442 (N_31442,N_21419,N_22975);
xor U31443 (N_31443,N_27349,N_28779);
xor U31444 (N_31444,N_23220,N_28683);
and U31445 (N_31445,N_23830,N_26936);
nor U31446 (N_31446,N_20769,N_29034);
or U31447 (N_31447,N_20992,N_29973);
or U31448 (N_31448,N_23966,N_26056);
and U31449 (N_31449,N_24167,N_21790);
nor U31450 (N_31450,N_24823,N_26543);
or U31451 (N_31451,N_20839,N_21189);
nand U31452 (N_31452,N_25926,N_20573);
and U31453 (N_31453,N_24240,N_29986);
or U31454 (N_31454,N_29531,N_20924);
nor U31455 (N_31455,N_27561,N_24630);
nor U31456 (N_31456,N_23556,N_28341);
or U31457 (N_31457,N_23292,N_27026);
nor U31458 (N_31458,N_28027,N_25955);
nor U31459 (N_31459,N_28276,N_21925);
nand U31460 (N_31460,N_26642,N_23430);
xor U31461 (N_31461,N_23164,N_24499);
or U31462 (N_31462,N_22292,N_23434);
xnor U31463 (N_31463,N_22344,N_20816);
xnor U31464 (N_31464,N_29205,N_26242);
xnor U31465 (N_31465,N_27578,N_25807);
nand U31466 (N_31466,N_20952,N_22562);
nand U31467 (N_31467,N_28000,N_25496);
and U31468 (N_31468,N_28073,N_28338);
and U31469 (N_31469,N_22265,N_29569);
or U31470 (N_31470,N_26801,N_20073);
and U31471 (N_31471,N_27714,N_20277);
nor U31472 (N_31472,N_26763,N_28170);
and U31473 (N_31473,N_22865,N_29110);
xor U31474 (N_31474,N_25198,N_28351);
or U31475 (N_31475,N_25041,N_25319);
nor U31476 (N_31476,N_22884,N_22355);
or U31477 (N_31477,N_21983,N_21161);
nand U31478 (N_31478,N_27531,N_21870);
xor U31479 (N_31479,N_22064,N_27437);
or U31480 (N_31480,N_21523,N_25612);
nand U31481 (N_31481,N_22739,N_28191);
and U31482 (N_31482,N_27169,N_28122);
nor U31483 (N_31483,N_29133,N_24571);
or U31484 (N_31484,N_23135,N_28902);
nand U31485 (N_31485,N_24608,N_24982);
xor U31486 (N_31486,N_26357,N_24496);
or U31487 (N_31487,N_21785,N_24156);
or U31488 (N_31488,N_22794,N_20161);
nand U31489 (N_31489,N_21034,N_25299);
and U31490 (N_31490,N_22715,N_28663);
nor U31491 (N_31491,N_29763,N_27352);
xnor U31492 (N_31492,N_22407,N_27640);
xor U31493 (N_31493,N_21134,N_20658);
or U31494 (N_31494,N_21641,N_23352);
nand U31495 (N_31495,N_25501,N_28342);
xnor U31496 (N_31496,N_29491,N_23314);
nor U31497 (N_31497,N_29766,N_28391);
nand U31498 (N_31498,N_23288,N_25588);
and U31499 (N_31499,N_27069,N_27053);
and U31500 (N_31500,N_23215,N_22805);
and U31501 (N_31501,N_23506,N_28738);
xnor U31502 (N_31502,N_27436,N_24459);
nand U31503 (N_31503,N_22872,N_28667);
xor U31504 (N_31504,N_27256,N_29314);
xnor U31505 (N_31505,N_25112,N_26963);
and U31506 (N_31506,N_27814,N_24787);
nor U31507 (N_31507,N_28438,N_20964);
nor U31508 (N_31508,N_27217,N_28011);
or U31509 (N_31509,N_20939,N_20484);
xor U31510 (N_31510,N_27421,N_27051);
or U31511 (N_31511,N_27320,N_23106);
or U31512 (N_31512,N_29487,N_26732);
or U31513 (N_31513,N_24843,N_25435);
and U31514 (N_31514,N_28048,N_27980);
or U31515 (N_31515,N_27700,N_27740);
or U31516 (N_31516,N_23400,N_26915);
and U31517 (N_31517,N_27718,N_22814);
or U31518 (N_31518,N_20402,N_27716);
and U31519 (N_31519,N_23501,N_20570);
nor U31520 (N_31520,N_25086,N_27930);
and U31521 (N_31521,N_22191,N_27058);
nand U31522 (N_31522,N_25883,N_27958);
or U31523 (N_31523,N_27112,N_26710);
nor U31524 (N_31524,N_28969,N_26886);
nand U31525 (N_31525,N_28710,N_28587);
xnor U31526 (N_31526,N_26804,N_28091);
xnor U31527 (N_31527,N_26473,N_29592);
and U31528 (N_31528,N_24629,N_29264);
nand U31529 (N_31529,N_23760,N_20677);
nor U31530 (N_31530,N_20387,N_29552);
nor U31531 (N_31531,N_21793,N_26438);
nand U31532 (N_31532,N_22057,N_22533);
nor U31533 (N_31533,N_28286,N_24210);
nand U31534 (N_31534,N_27380,N_20636);
xnor U31535 (N_31535,N_22165,N_26039);
and U31536 (N_31536,N_21722,N_20838);
xor U31537 (N_31537,N_28386,N_21807);
nand U31538 (N_31538,N_22334,N_27969);
and U31539 (N_31539,N_26832,N_24432);
and U31540 (N_31540,N_20641,N_25861);
or U31541 (N_31541,N_28896,N_29283);
nand U31542 (N_31542,N_24080,N_21697);
nand U31543 (N_31543,N_25537,N_20988);
and U31544 (N_31544,N_27929,N_28436);
xnor U31545 (N_31545,N_21111,N_23924);
xor U31546 (N_31546,N_26718,N_24513);
nor U31547 (N_31547,N_23405,N_21009);
xnor U31548 (N_31548,N_28298,N_20717);
and U31549 (N_31549,N_25004,N_25044);
nor U31550 (N_31550,N_24075,N_24976);
xor U31551 (N_31551,N_24289,N_27707);
nand U31552 (N_31552,N_28559,N_28589);
or U31553 (N_31553,N_29021,N_25369);
nor U31554 (N_31554,N_21510,N_27636);
xor U31555 (N_31555,N_27503,N_23071);
or U31556 (N_31556,N_25828,N_28547);
and U31557 (N_31557,N_28706,N_22279);
nor U31558 (N_31558,N_27649,N_21888);
or U31559 (N_31559,N_27758,N_26198);
or U31560 (N_31560,N_22999,N_22941);
nor U31561 (N_31561,N_26061,N_25647);
and U31562 (N_31562,N_23837,N_25634);
and U31563 (N_31563,N_21563,N_26244);
or U31564 (N_31564,N_23067,N_28828);
xnor U31565 (N_31565,N_25286,N_21945);
xor U31566 (N_31566,N_27634,N_24502);
or U31567 (N_31567,N_22123,N_29853);
xnor U31568 (N_31568,N_29858,N_25233);
nand U31569 (N_31569,N_29672,N_24944);
and U31570 (N_31570,N_21427,N_27552);
xor U31571 (N_31571,N_28065,N_29360);
xnor U31572 (N_31572,N_24176,N_26082);
nor U31573 (N_31573,N_24062,N_28850);
nand U31574 (N_31574,N_25593,N_29747);
and U31575 (N_31575,N_24004,N_29416);
nor U31576 (N_31576,N_24448,N_20198);
or U31577 (N_31577,N_28816,N_24077);
and U31578 (N_31578,N_27426,N_25220);
nand U31579 (N_31579,N_26814,N_28510);
xor U31580 (N_31580,N_28323,N_22786);
nor U31581 (N_31581,N_27646,N_26179);
xor U31582 (N_31582,N_25857,N_20930);
or U31583 (N_31583,N_24659,N_29158);
nand U31584 (N_31584,N_22055,N_23302);
and U31585 (N_31585,N_23992,N_29439);
nand U31586 (N_31586,N_26714,N_28106);
nor U31587 (N_31587,N_20664,N_25996);
and U31588 (N_31588,N_29679,N_22303);
nor U31589 (N_31589,N_20665,N_29115);
nand U31590 (N_31590,N_23406,N_29452);
xnor U31591 (N_31591,N_29526,N_23605);
nor U31592 (N_31592,N_25556,N_28397);
and U31593 (N_31593,N_22301,N_27306);
xnor U31594 (N_31594,N_26700,N_29105);
and U31595 (N_31595,N_29816,N_28577);
or U31596 (N_31596,N_23649,N_26257);
or U31597 (N_31597,N_21050,N_25082);
nor U31598 (N_31598,N_25937,N_29819);
nor U31599 (N_31599,N_27767,N_28613);
nand U31600 (N_31600,N_26034,N_21860);
or U31601 (N_31601,N_23163,N_27759);
xor U31602 (N_31602,N_20131,N_21596);
nor U31603 (N_31603,N_22690,N_25770);
or U31604 (N_31604,N_26823,N_29579);
xor U31605 (N_31605,N_22448,N_28076);
xnor U31606 (N_31606,N_28480,N_24977);
nor U31607 (N_31607,N_24306,N_24344);
or U31608 (N_31608,N_25572,N_26426);
xor U31609 (N_31609,N_21847,N_29626);
nor U31610 (N_31610,N_27277,N_22510);
or U31611 (N_31611,N_23277,N_27849);
or U31612 (N_31612,N_26336,N_28615);
nor U31613 (N_31613,N_29053,N_29865);
xor U31614 (N_31614,N_22177,N_21234);
xor U31615 (N_31615,N_25709,N_29289);
nand U31616 (N_31616,N_24329,N_24671);
nand U31617 (N_31617,N_26827,N_29972);
nor U31618 (N_31618,N_20153,N_27078);
nand U31619 (N_31619,N_27499,N_20722);
nor U31620 (N_31620,N_20330,N_27815);
or U31621 (N_31621,N_27782,N_20460);
nand U31622 (N_31622,N_23301,N_20589);
and U31623 (N_31623,N_23438,N_28539);
or U31624 (N_31624,N_26735,N_24096);
xor U31625 (N_31625,N_29152,N_21724);
or U31626 (N_31626,N_20103,N_24705);
xnor U31627 (N_31627,N_29399,N_22481);
nor U31628 (N_31628,N_25689,N_29574);
nand U31629 (N_31629,N_22906,N_29930);
xor U31630 (N_31630,N_27045,N_27696);
and U31631 (N_31631,N_21130,N_29501);
or U31632 (N_31632,N_23143,N_21928);
or U31633 (N_31633,N_24678,N_27120);
and U31634 (N_31634,N_26448,N_25168);
or U31635 (N_31635,N_25530,N_26838);
nand U31636 (N_31636,N_27094,N_20094);
and U31637 (N_31637,N_22300,N_28124);
nand U31638 (N_31638,N_25964,N_22712);
or U31639 (N_31639,N_22784,N_21382);
nor U31640 (N_31640,N_28025,N_23906);
xor U31641 (N_31641,N_27683,N_28768);
nand U31642 (N_31642,N_29039,N_23728);
xor U31643 (N_31643,N_27109,N_27395);
nor U31644 (N_31644,N_23637,N_24258);
or U31645 (N_31645,N_25030,N_21055);
xor U31646 (N_31646,N_26447,N_20845);
or U31647 (N_31647,N_22200,N_20171);
and U31648 (N_31648,N_25809,N_22832);
nor U31649 (N_31649,N_21063,N_29826);
and U31650 (N_31650,N_21140,N_20229);
nand U31651 (N_31651,N_28600,N_28529);
and U31652 (N_31652,N_24870,N_24093);
nor U31653 (N_31653,N_25108,N_25431);
nor U31654 (N_31654,N_21629,N_29078);
and U31655 (N_31655,N_22120,N_28321);
or U31656 (N_31656,N_22087,N_27295);
nand U31657 (N_31657,N_27599,N_24497);
nor U31658 (N_31658,N_24694,N_29856);
nor U31659 (N_31659,N_25579,N_25430);
xor U31660 (N_31660,N_29742,N_29698);
nand U31661 (N_31661,N_20074,N_29831);
and U31662 (N_31662,N_21021,N_21418);
nand U31663 (N_31663,N_21110,N_22074);
nor U31664 (N_31664,N_25638,N_26680);
xnor U31665 (N_31665,N_20009,N_29646);
and U31666 (N_31666,N_22659,N_20783);
nand U31667 (N_31667,N_23845,N_29689);
or U31668 (N_31668,N_23669,N_20029);
and U31669 (N_31669,N_25815,N_28761);
nor U31670 (N_31670,N_29923,N_26805);
xnor U31671 (N_31671,N_23268,N_20062);
xnor U31672 (N_31672,N_24269,N_22702);
nand U31673 (N_31673,N_29910,N_26888);
or U31674 (N_31674,N_23346,N_26286);
nand U31675 (N_31675,N_23631,N_29397);
nand U31676 (N_31676,N_23774,N_29313);
nand U31677 (N_31677,N_22844,N_20890);
and U31678 (N_31678,N_24421,N_26345);
nor U31679 (N_31679,N_29191,N_28206);
or U31680 (N_31680,N_22993,N_25150);
xor U31681 (N_31681,N_25376,N_26785);
and U31682 (N_31682,N_23511,N_22628);
and U31683 (N_31683,N_24552,N_22272);
and U31684 (N_31684,N_20525,N_23572);
and U31685 (N_31685,N_23378,N_25762);
xnor U31686 (N_31686,N_27684,N_23585);
nor U31687 (N_31687,N_28360,N_20162);
and U31688 (N_31688,N_26600,N_28942);
xnor U31689 (N_31689,N_23552,N_23578);
and U31690 (N_31690,N_21677,N_20310);
or U31691 (N_31691,N_26117,N_23233);
xor U31692 (N_31692,N_20639,N_24398);
nor U31693 (N_31693,N_28478,N_24923);
or U31694 (N_31694,N_20706,N_22687);
xnor U31695 (N_31695,N_23334,N_29330);
and U31696 (N_31696,N_26455,N_27377);
nand U31697 (N_31697,N_24789,N_23509);
or U31698 (N_31698,N_26806,N_25361);
and U31699 (N_31699,N_29959,N_25023);
nor U31700 (N_31700,N_27513,N_27269);
nand U31701 (N_31701,N_20179,N_21304);
or U31702 (N_31702,N_26208,N_29994);
nand U31703 (N_31703,N_26421,N_21025);
nand U31704 (N_31704,N_27907,N_20024);
or U31705 (N_31705,N_28873,N_20149);
xor U31706 (N_31706,N_25327,N_26687);
or U31707 (N_31707,N_27310,N_21039);
nor U31708 (N_31708,N_20098,N_24228);
or U31709 (N_31709,N_26023,N_23770);
xor U31710 (N_31710,N_27432,N_22322);
xnor U31711 (N_31711,N_24034,N_29787);
and U31712 (N_31712,N_28135,N_25758);
xnor U31713 (N_31713,N_28923,N_20674);
and U31714 (N_31714,N_25068,N_23777);
and U31715 (N_31715,N_20977,N_24407);
or U31716 (N_31716,N_20911,N_26865);
xor U31717 (N_31717,N_26552,N_20357);
or U31718 (N_31718,N_26051,N_22791);
and U31719 (N_31719,N_20081,N_21400);
and U31720 (N_31720,N_21676,N_26128);
nand U31721 (N_31721,N_22614,N_20709);
nor U31722 (N_31722,N_20440,N_24249);
xor U31723 (N_31723,N_21799,N_22096);
nor U31724 (N_31724,N_27239,N_29600);
and U31725 (N_31725,N_27807,N_28009);
or U31726 (N_31726,N_22837,N_27673);
nand U31727 (N_31727,N_21378,N_26168);
nor U31728 (N_31728,N_27691,N_24901);
and U31729 (N_31729,N_23116,N_22088);
nand U31730 (N_31730,N_27496,N_29200);
and U31731 (N_31731,N_20467,N_23673);
xor U31732 (N_31732,N_21387,N_27184);
and U31733 (N_31733,N_27165,N_29499);
nand U31734 (N_31734,N_21905,N_25998);
or U31735 (N_31735,N_28620,N_28118);
nor U31736 (N_31736,N_22616,N_27976);
or U31737 (N_31737,N_22896,N_24914);
or U31738 (N_31738,N_20363,N_27029);
nor U31739 (N_31739,N_23559,N_23134);
nand U31740 (N_31740,N_26689,N_22004);
nand U31741 (N_31741,N_24666,N_21470);
and U31742 (N_31742,N_26518,N_23091);
nand U31743 (N_31743,N_28431,N_24135);
nand U31744 (N_31744,N_21828,N_26052);
or U31745 (N_31745,N_24410,N_28062);
nor U31746 (N_31746,N_26881,N_26549);
or U31747 (N_31747,N_25546,N_28083);
or U31748 (N_31748,N_28072,N_27972);
xor U31749 (N_31749,N_29024,N_21803);
nand U31750 (N_31750,N_25818,N_26775);
and U31751 (N_31751,N_22662,N_26305);
and U31752 (N_31752,N_26914,N_29820);
and U31753 (N_31753,N_29909,N_26671);
or U31754 (N_31754,N_20735,N_27233);
nand U31755 (N_31755,N_28887,N_28396);
or U31756 (N_31756,N_24695,N_20466);
and U31757 (N_31757,N_23452,N_29559);
or U31758 (N_31758,N_25155,N_25904);
nor U31759 (N_31759,N_23741,N_23145);
or U31760 (N_31760,N_28628,N_26045);
and U31761 (N_31761,N_29310,N_27358);
or U31762 (N_31762,N_25915,N_26186);
nor U31763 (N_31763,N_28982,N_22916);
nand U31764 (N_31764,N_22260,N_24567);
and U31765 (N_31765,N_26878,N_28732);
xnor U31766 (N_31766,N_27183,N_22460);
and U31767 (N_31767,N_23060,N_24111);
and U31768 (N_31768,N_23611,N_20298);
nor U31769 (N_31769,N_21053,N_25275);
or U31770 (N_31770,N_25154,N_27523);
nor U31771 (N_31771,N_24254,N_23508);
nor U31772 (N_31772,N_24256,N_25829);
and U31773 (N_31773,N_21769,N_25161);
xnor U31774 (N_31774,N_28455,N_26774);
nor U31775 (N_31775,N_29136,N_24057);
and U31776 (N_31776,N_28247,N_23204);
xnor U31777 (N_31777,N_24397,N_24188);
nor U31778 (N_31778,N_25287,N_29490);
nor U31779 (N_31779,N_23068,N_26070);
xnor U31780 (N_31780,N_27754,N_21414);
xnor U31781 (N_31781,N_23832,N_24724);
and U31782 (N_31782,N_24102,N_20052);
nor U31783 (N_31783,N_28057,N_25521);
or U31784 (N_31784,N_27083,N_24216);
or U31785 (N_31785,N_26169,N_20186);
or U31786 (N_31786,N_27941,N_21467);
and U31787 (N_31787,N_28462,N_26496);
nor U31788 (N_31788,N_29676,N_29002);
and U31789 (N_31789,N_21230,N_23913);
or U31790 (N_31790,N_24778,N_20879);
or U31791 (N_31791,N_25204,N_26281);
nand U31792 (N_31792,N_20957,N_27846);
nand U31793 (N_31793,N_20739,N_26337);
nand U31794 (N_31794,N_29818,N_25174);
xor U31795 (N_31795,N_29807,N_23981);
xor U31796 (N_31796,N_21650,N_24903);
xor U31797 (N_31797,N_26770,N_24316);
nand U31798 (N_31798,N_25073,N_26038);
xnor U31799 (N_31799,N_22897,N_28052);
nor U31800 (N_31800,N_21816,N_24118);
xor U31801 (N_31801,N_24183,N_20354);
nand U31802 (N_31802,N_22416,N_25476);
xor U31803 (N_31803,N_24738,N_26156);
xnor U31804 (N_31804,N_22219,N_22472);
nor U31805 (N_31805,N_20032,N_29801);
nor U31806 (N_31806,N_24568,N_20434);
xor U31807 (N_31807,N_24955,N_29046);
nand U31808 (N_31808,N_23465,N_27105);
and U31809 (N_31809,N_23658,N_20983);
or U31810 (N_31810,N_21084,N_25485);
nor U31811 (N_31811,N_25103,N_22757);
or U31812 (N_31812,N_25587,N_20297);
nand U31813 (N_31813,N_29446,N_22206);
nor U31814 (N_31814,N_24957,N_23350);
xor U31815 (N_31815,N_22453,N_22675);
nand U31816 (N_31816,N_29489,N_23748);
nand U31817 (N_31817,N_26840,N_26858);
and U31818 (N_31818,N_28484,N_29738);
nand U31819 (N_31819,N_24604,N_27851);
nand U31820 (N_31820,N_28470,N_28330);
xnor U31821 (N_31821,N_29449,N_22065);
and U31822 (N_31822,N_29668,N_27453);
nand U31823 (N_31823,N_29514,N_28499);
or U31824 (N_31824,N_24292,N_20820);
xnor U31825 (N_31825,N_23100,N_29441);
nor U31826 (N_31826,N_22582,N_24159);
nand U31827 (N_31827,N_29786,N_23725);
nand U31828 (N_31828,N_24736,N_26776);
or U31829 (N_31829,N_29595,N_20455);
xnor U31830 (N_31830,N_21539,N_28751);
and U31831 (N_31831,N_28889,N_21171);
nand U31832 (N_31832,N_21766,N_20575);
xor U31833 (N_31833,N_26348,N_28653);
nand U31834 (N_31834,N_22564,N_25966);
or U31835 (N_31835,N_22869,N_25877);
and U31836 (N_31836,N_26893,N_21726);
xor U31837 (N_31837,N_20903,N_22218);
nand U31838 (N_31838,N_23627,N_25406);
nand U31839 (N_31839,N_24043,N_26444);
nor U31840 (N_31840,N_29932,N_25371);
nand U31841 (N_31841,N_25021,N_27157);
nand U31842 (N_31842,N_27799,N_21490);
nor U31843 (N_31843,N_25244,N_24124);
nor U31844 (N_31844,N_27511,N_20381);
and U31845 (N_31845,N_20082,N_24039);
and U31846 (N_31846,N_27160,N_27113);
and U31847 (N_31847,N_29591,N_23401);
and U31848 (N_31848,N_25963,N_23995);
nor U31849 (N_31849,N_25969,N_20339);
nor U31850 (N_31850,N_25983,N_22536);
nand U31851 (N_31851,N_28743,N_20592);
xnor U31852 (N_31852,N_22019,N_26905);
or U31853 (N_31853,N_24973,N_22186);
or U31854 (N_31854,N_25383,N_25970);
and U31855 (N_31855,N_29896,N_20104);
nand U31856 (N_31856,N_20367,N_25069);
and U31857 (N_31857,N_26062,N_23734);
nand U31858 (N_31858,N_21143,N_28190);
nor U31859 (N_31859,N_23870,N_26042);
nand U31860 (N_31860,N_28102,N_28596);
and U31861 (N_31861,N_26729,N_25505);
nand U31862 (N_31862,N_22828,N_28908);
nor U31863 (N_31863,N_27826,N_29583);
xnor U31864 (N_31864,N_29203,N_23022);
or U31865 (N_31865,N_27099,N_25389);
or U31866 (N_31866,N_20737,N_25787);
xnor U31867 (N_31867,N_29871,N_20954);
nand U31868 (N_31868,N_21834,N_29751);
xor U31869 (N_31869,N_28259,N_22109);
xnor U31870 (N_31870,N_20045,N_25848);
nand U31871 (N_31871,N_27785,N_29710);
nor U31872 (N_31872,N_20910,N_26742);
nor U31873 (N_31873,N_21963,N_29944);
or U31874 (N_31874,N_23274,N_26277);
nor U31875 (N_31875,N_22987,N_27884);
xor U31876 (N_31876,N_27235,N_21067);
and U31877 (N_31877,N_20192,N_21776);
nand U31878 (N_31878,N_24554,N_26647);
nand U31879 (N_31879,N_26929,N_22333);
nand U31880 (N_31880,N_25293,N_24890);
and U31881 (N_31881,N_20650,N_23991);
or U31882 (N_31882,N_24684,N_24429);
and U31883 (N_31883,N_28713,N_27960);
nand U31884 (N_31884,N_28655,N_22781);
xor U31885 (N_31885,N_20415,N_29190);
nor U31886 (N_31886,N_22213,N_22692);
or U31887 (N_31887,N_28362,N_23618);
and U31888 (N_31888,N_20659,N_22288);
nor U31889 (N_31889,N_22539,N_20716);
nor U31890 (N_31890,N_28142,N_28465);
nor U31891 (N_31891,N_23839,N_23045);
nand U31892 (N_31892,N_20965,N_22280);
and U31893 (N_31893,N_20048,N_21013);
and U31894 (N_31894,N_21381,N_25669);
nor U31895 (N_31895,N_22776,N_28093);
nor U31896 (N_31896,N_21199,N_24786);
nand U31897 (N_31897,N_25285,N_25412);
nor U31898 (N_31898,N_27593,N_21655);
or U31899 (N_31899,N_28175,N_20255);
nand U31900 (N_31900,N_25929,N_25626);
nor U31901 (N_31901,N_21390,N_25991);
and U31902 (N_31902,N_25902,N_23788);
xor U31903 (N_31903,N_22172,N_24602);
nand U31904 (N_31904,N_20626,N_26930);
nand U31905 (N_31905,N_22567,N_26347);
or U31906 (N_31906,N_23252,N_23230);
and U31907 (N_31907,N_29167,N_20914);
or U31908 (N_31908,N_29849,N_20807);
nor U31909 (N_31909,N_27617,N_20037);
or U31910 (N_31910,N_24626,N_25316);
and U31911 (N_31911,N_29204,N_26430);
nor U31912 (N_31912,N_28333,N_29565);
nor U31913 (N_31913,N_21782,N_25676);
nand U31914 (N_31914,N_26560,N_29980);
xor U31915 (N_31915,N_26699,N_20253);
xnor U31916 (N_31916,N_26501,N_20433);
and U31917 (N_31917,N_21854,N_22737);
and U31918 (N_31918,N_24503,N_22967);
xor U31919 (N_31919,N_21773,N_23458);
xnor U31920 (N_31920,N_22929,N_24618);
and U31921 (N_31921,N_27750,N_26404);
nand U31922 (N_31922,N_26995,N_21242);
nor U31923 (N_31923,N_24153,N_25078);
nand U31924 (N_31924,N_23075,N_23418);
xnor U31925 (N_31925,N_27093,N_25502);
nor U31926 (N_31926,N_27845,N_22447);
or U31927 (N_31927,N_28618,N_25892);
or U31928 (N_31928,N_28821,N_21177);
xor U31929 (N_31929,N_20166,N_21550);
nor U31930 (N_31930,N_28552,N_25467);
nor U31931 (N_31931,N_21950,N_21210);
nor U31932 (N_31932,N_29718,N_28001);
nand U31933 (N_31933,N_26067,N_25118);
nand U31934 (N_31934,N_23450,N_26713);
nand U31935 (N_31935,N_27355,N_22262);
and U31936 (N_31936,N_27676,N_20437);
nor U31937 (N_31937,N_21404,N_27524);
nand U31938 (N_31938,N_23996,N_20758);
nand U31939 (N_31939,N_28082,N_26114);
nand U31940 (N_31940,N_23513,N_21577);
nand U31941 (N_31941,N_22630,N_26578);
and U31942 (N_31942,N_28945,N_20750);
and U31943 (N_31943,N_28774,N_27036);
and U31944 (N_31944,N_21509,N_24596);
nor U31945 (N_31945,N_22508,N_25219);
and U31946 (N_31946,N_25202,N_26715);
nand U31947 (N_31947,N_28216,N_27518);
nor U31948 (N_31948,N_25695,N_27155);
xnor U31949 (N_31949,N_21398,N_22641);
nor U31950 (N_31950,N_26011,N_22424);
xnor U31951 (N_31951,N_29659,N_23294);
or U31952 (N_31952,N_22070,N_26989);
nand U31953 (N_31953,N_25255,N_23034);
and U31954 (N_31954,N_20543,N_25305);
nor U31955 (N_31955,N_22795,N_25107);
and U31956 (N_31956,N_27719,N_29788);
nand U31957 (N_31957,N_21358,N_24498);
and U31958 (N_31958,N_21904,N_21012);
and U31959 (N_31959,N_28723,N_20132);
xnor U31960 (N_31960,N_28400,N_23315);
xnor U31961 (N_31961,N_26399,N_28783);
or U31962 (N_31962,N_23228,N_24166);
or U31963 (N_31963,N_21228,N_26422);
nand U31964 (N_31964,N_25330,N_22330);
xor U31965 (N_31965,N_21279,N_24239);
xor U31966 (N_31966,N_20180,N_27698);
xnor U31967 (N_31967,N_26698,N_26326);
nand U31968 (N_31968,N_25790,N_20476);
nor U31969 (N_31969,N_25532,N_29543);
nor U31970 (N_31970,N_22100,N_27174);
nand U31971 (N_31971,N_27722,N_27705);
nand U31972 (N_31972,N_25710,N_29688);
and U31973 (N_31973,N_29866,N_29725);
xor U31974 (N_31974,N_22225,N_24993);
nor U31975 (N_31975,N_26666,N_25137);
nand U31976 (N_31976,N_28130,N_23901);
nand U31977 (N_31977,N_27928,N_25152);
xnor U31978 (N_31978,N_27635,N_25599);
xor U31979 (N_31979,N_29277,N_25265);
nor U31980 (N_31980,N_26769,N_20383);
nor U31981 (N_31981,N_22883,N_22130);
nor U31982 (N_31982,N_20785,N_23421);
nor U31983 (N_31983,N_20016,N_24715);
nor U31984 (N_31984,N_28421,N_29454);
and U31985 (N_31985,N_22027,N_21607);
nor U31986 (N_31986,N_21428,N_29379);
nor U31987 (N_31987,N_23286,N_20054);
nor U31988 (N_31988,N_29217,N_20331);
and U31989 (N_31989,N_24852,N_26708);
nand U31990 (N_31990,N_23956,N_21822);
nor U31991 (N_31991,N_25700,N_28934);
and U31992 (N_31992,N_25549,N_24468);
nor U31993 (N_31993,N_25243,N_28773);
nand U31994 (N_31994,N_28722,N_27641);
nor U31995 (N_31995,N_28490,N_28203);
and U31996 (N_31996,N_20646,N_29369);
and U31997 (N_31997,N_25860,N_22909);
and U31998 (N_31998,N_22180,N_23009);
or U31999 (N_31999,N_27332,N_20479);
nand U32000 (N_32000,N_23141,N_29141);
nand U32001 (N_32001,N_29796,N_29231);
and U32002 (N_32002,N_29851,N_28711);
and U32003 (N_32003,N_21144,N_24202);
nand U32004 (N_32004,N_24932,N_27529);
xor U32005 (N_32005,N_27460,N_27622);
nand U32006 (N_32006,N_25461,N_21138);
or U32007 (N_32007,N_21943,N_21392);
xor U32008 (N_32008,N_26292,N_29035);
or U32009 (N_32009,N_23456,N_26253);
nor U32010 (N_32010,N_22489,N_21379);
and U32011 (N_32011,N_24746,N_23169);
xnor U32012 (N_32012,N_26153,N_25564);
nor U32013 (N_32013,N_25237,N_28010);
xnor U32014 (N_32014,N_28670,N_22400);
nand U32015 (N_32015,N_28327,N_24758);
xnor U32016 (N_32016,N_24291,N_20733);
nand U32017 (N_32017,N_25390,N_27212);
nand U32018 (N_32018,N_24679,N_26354);
and U32019 (N_32019,N_27608,N_26817);
xnor U32020 (N_32020,N_27483,N_23802);
or U32021 (N_32021,N_26503,N_27735);
nand U32022 (N_32022,N_23661,N_24371);
nand U32023 (N_32023,N_28964,N_23620);
xnor U32024 (N_32024,N_20718,N_24107);
or U32025 (N_32025,N_28047,N_21129);
nor U32026 (N_32026,N_26331,N_21384);
nand U32027 (N_32027,N_23155,N_29663);
nor U32028 (N_32028,N_24423,N_21364);
or U32029 (N_32029,N_22174,N_24349);
xor U32030 (N_32030,N_29503,N_25156);
nor U32031 (N_32031,N_27134,N_29375);
or U32032 (N_32032,N_27110,N_20567);
nand U32033 (N_32033,N_22201,N_26307);
xnor U32034 (N_32034,N_21081,N_27378);
or U32035 (N_32035,N_27840,N_21122);
nor U32036 (N_32036,N_22550,N_21344);
or U32037 (N_32037,N_23644,N_23546);
nor U32038 (N_32038,N_24586,N_28707);
or U32039 (N_32039,N_23794,N_28192);
nor U32040 (N_32040,N_22694,N_28344);
xnor U32041 (N_32041,N_20900,N_28543);
nor U32042 (N_32042,N_23189,N_20623);
nor U32043 (N_32043,N_29386,N_29758);
xnor U32044 (N_32044,N_29628,N_29914);
xnor U32045 (N_32045,N_29570,N_28222);
xnor U32046 (N_32046,N_28717,N_29424);
xor U32047 (N_32047,N_20373,N_28468);
and U32048 (N_32048,N_27619,N_21312);
or U32049 (N_32049,N_24794,N_23829);
and U32050 (N_32050,N_21578,N_25602);
and U32051 (N_32051,N_28762,N_29836);
and U32052 (N_32052,N_28754,N_29848);
nor U32053 (N_32053,N_29477,N_28218);
nand U32054 (N_32054,N_22208,N_25097);
or U32055 (N_32055,N_20240,N_27159);
xnor U32056 (N_32056,N_26711,N_23516);
xor U32057 (N_32057,N_20529,N_27101);
nand U32058 (N_32058,N_29857,N_27150);
xor U32059 (N_32059,N_25494,N_25251);
nand U32060 (N_32060,N_28046,N_22612);
or U32061 (N_32061,N_29546,N_23321);
nand U32062 (N_32062,N_25935,N_20411);
or U32063 (N_32063,N_25974,N_29081);
and U32064 (N_32064,N_27228,N_29922);
or U32065 (N_32065,N_22427,N_27119);
nand U32066 (N_32066,N_20742,N_25079);
nor U32067 (N_32067,N_25613,N_25151);
nand U32068 (N_32068,N_25264,N_29333);
xor U32069 (N_32069,N_28066,N_23577);
or U32070 (N_32070,N_25900,N_24575);
and U32071 (N_32071,N_28383,N_24954);
xor U32072 (N_32072,N_24711,N_28981);
and U32073 (N_32073,N_26901,N_23755);
nand U32074 (N_32074,N_29362,N_24873);
nand U32075 (N_32075,N_23727,N_21995);
or U32076 (N_32076,N_23069,N_24916);
nor U32077 (N_32077,N_22696,N_29429);
or U32078 (N_32078,N_28802,N_20822);
or U32079 (N_32079,N_21494,N_24769);
xor U32080 (N_32080,N_20013,N_23554);
nand U32081 (N_32081,N_24205,N_25077);
and U32082 (N_32082,N_26368,N_23532);
nand U32083 (N_32083,N_23514,N_24074);
and U32084 (N_32084,N_20721,N_24951);
and U32085 (N_32085,N_28714,N_29211);
xor U32086 (N_32086,N_20776,N_26511);
or U32087 (N_32087,N_27834,N_24790);
nor U32088 (N_32088,N_29716,N_21233);
or U32089 (N_32089,N_27688,N_26946);
nor U32090 (N_32090,N_27964,N_20878);
or U32091 (N_32091,N_22988,N_25019);
xnor U32092 (N_32092,N_21648,N_26933);
nor U32093 (N_32093,N_23167,N_20319);
nor U32094 (N_32094,N_23959,N_27690);
nor U32095 (N_32095,N_29642,N_23574);
nand U32096 (N_32096,N_27201,N_27431);
and U32097 (N_32097,N_21628,N_21362);
xnor U32098 (N_32098,N_22599,N_24691);
nor U32099 (N_32099,N_21431,N_28715);
or U32100 (N_32100,N_26683,N_27832);
nand U32101 (N_32101,N_28388,N_25639);
and U32102 (N_32102,N_29469,N_22762);
nor U32103 (N_32103,N_23820,N_25632);
nor U32104 (N_32104,N_28948,N_21589);
and U32105 (N_32105,N_21855,N_28008);
and U32106 (N_32106,N_29080,N_22871);
nor U32107 (N_32107,N_22455,N_29048);
and U32108 (N_32108,N_26544,N_20766);
and U32109 (N_32109,N_20909,N_20806);
xnor U32110 (N_32110,N_25445,N_20102);
nand U32111 (N_32111,N_22864,N_20585);
xor U32112 (N_32112,N_29007,N_23451);
xnor U32113 (N_32113,N_21565,N_28054);
nor U32114 (N_32114,N_28575,N_28912);
and U32115 (N_32115,N_21425,N_25022);
nor U32116 (N_32116,N_24101,N_21047);
or U32117 (N_32117,N_28453,N_21267);
xor U32118 (N_32118,N_25547,N_27761);
nand U32119 (N_32119,N_21942,N_21007);
nor U32120 (N_32120,N_23156,N_27033);
xnor U32121 (N_32121,N_24538,N_21603);
nor U32122 (N_32122,N_28852,N_27508);
and U32123 (N_32123,N_24312,N_28926);
or U32124 (N_32124,N_22259,N_22663);
or U32125 (N_32125,N_20973,N_27585);
nor U32126 (N_32126,N_24441,N_20244);
nor U32127 (N_32127,N_28960,N_26462);
or U32128 (N_32128,N_21895,N_25440);
xnor U32129 (N_32129,N_21239,N_24584);
nor U32130 (N_32130,N_24300,N_26230);
and U32131 (N_32131,N_20827,N_21751);
and U32132 (N_32132,N_29555,N_20563);
xor U32133 (N_32133,N_26508,N_21737);
or U32134 (N_32134,N_29832,N_26940);
nor U32135 (N_32135,N_23140,N_24158);
nor U32136 (N_32136,N_25400,N_27915);
and U32137 (N_32137,N_29298,N_21347);
nor U32138 (N_32138,N_29500,N_28520);
nand U32139 (N_32139,N_28983,N_25946);
nand U32140 (N_32140,N_24850,N_20364);
xor U32141 (N_32141,N_28105,N_22283);
xnor U32142 (N_32142,N_24800,N_21723);
nor U32143 (N_32143,N_29294,N_28409);
nor U32144 (N_32144,N_28542,N_24935);
nand U32145 (N_32145,N_20163,N_23773);
and U32146 (N_32146,N_22777,N_25124);
xnor U32147 (N_32147,N_25303,N_20829);
xor U32148 (N_32148,N_23681,N_29433);
xnor U32149 (N_32149,N_29825,N_22138);
nand U32150 (N_32150,N_27161,N_23888);
xor U32151 (N_32151,N_28079,N_22538);
nand U32152 (N_32152,N_28607,N_22534);
or U32153 (N_32153,N_29540,N_25314);
nor U32154 (N_32154,N_27102,N_29197);
or U32155 (N_32155,N_20971,N_22529);
or U32156 (N_32156,N_26359,N_29792);
xnor U32157 (N_32157,N_29983,N_25134);
xor U32158 (N_32158,N_20874,N_26573);
xor U32159 (N_32159,N_24362,N_21101);
nand U32160 (N_32160,N_27238,N_20938);
and U32161 (N_32161,N_28522,N_28835);
nand U32162 (N_32162,N_28108,N_23715);
nand U32163 (N_32163,N_22635,N_28370);
or U32164 (N_32164,N_26283,N_26745);
nor U32165 (N_32165,N_26274,N_24363);
or U32166 (N_32166,N_23856,N_22648);
and U32167 (N_32167,N_25889,N_21266);
or U32168 (N_32168,N_27107,N_20275);
nand U32169 (N_32169,N_24593,N_29935);
nor U32170 (N_32170,N_22624,N_25851);
or U32171 (N_32171,N_23628,N_20539);
and U32172 (N_32172,N_25629,N_23377);
or U32173 (N_32173,N_23997,N_27888);
xnor U32174 (N_32174,N_21575,N_29192);
nor U32175 (N_32175,N_29867,N_25788);
or U32176 (N_32176,N_20574,N_20417);
and U32177 (N_32177,N_25279,N_28795);
nor U32178 (N_32178,N_23012,N_23357);
and U32179 (N_32179,N_20923,N_22544);
nand U32180 (N_32180,N_24474,N_21996);
nand U32181 (N_32181,N_28685,N_22005);
or U32182 (N_32182,N_27100,N_25301);
or U32183 (N_32183,N_28527,N_26371);
nor U32184 (N_32184,N_26535,N_25609);
nand U32185 (N_32185,N_22287,N_23048);
or U32186 (N_32186,N_28676,N_26104);
xnor U32187 (N_32187,N_25578,N_20690);
xor U32188 (N_32188,N_27793,N_29008);
or U32189 (N_32189,N_29054,N_24819);
or U32190 (N_32190,N_22325,N_24523);
xnor U32191 (N_32191,N_21142,N_24242);
nand U32192 (N_32192,N_24286,N_27975);
xnor U32193 (N_32193,N_21107,N_29692);
nand U32194 (N_32194,N_26851,N_21534);
xnor U32195 (N_32195,N_29554,N_25722);
nand U32196 (N_32196,N_23287,N_26889);
and U32197 (N_32197,N_23922,N_20734);
and U32198 (N_32198,N_22072,N_28031);
and U32199 (N_32199,N_28815,N_27932);
and U32200 (N_32200,N_29693,N_23266);
and U32201 (N_32201,N_27376,N_24548);
nand U32202 (N_32202,N_25999,N_24863);
nor U32203 (N_32203,N_22150,N_29639);
nand U32204 (N_32204,N_25442,N_25187);
and U32205 (N_32205,N_25804,N_21450);
or U32206 (N_32206,N_27572,N_22822);
nand U32207 (N_32207,N_28997,N_23951);
or U32208 (N_32208,N_21151,N_20287);
nand U32209 (N_32209,N_20369,N_26315);
or U32210 (N_32210,N_25470,N_23723);
xor U32211 (N_32211,N_26639,N_20165);
nand U32212 (N_32212,N_20391,N_25563);
nor U32213 (N_32213,N_22878,N_27300);
xnor U32214 (N_32214,N_21463,N_25276);
nor U32215 (N_32215,N_20226,N_22327);
xnor U32216 (N_32216,N_20998,N_20097);
or U32217 (N_32217,N_26591,N_29198);
nor U32218 (N_32218,N_25508,N_23128);
and U32219 (N_32219,N_26476,N_29687);
or U32220 (N_32220,N_26861,N_21546);
nor U32221 (N_32221,N_27204,N_29709);
or U32222 (N_32222,N_25749,N_23207);
and U32223 (N_32223,N_23267,N_25379);
nor U32224 (N_32224,N_21625,N_22184);
xor U32225 (N_32225,N_27769,N_25685);
and U32226 (N_32226,N_24653,N_20853);
xor U32227 (N_32227,N_29246,N_26633);
nor U32228 (N_32228,N_26076,N_28485);
and U32229 (N_32229,N_20842,N_21252);
and U32230 (N_32230,N_23835,N_23821);
or U32231 (N_32231,N_21309,N_28832);
nor U32232 (N_32232,N_27855,N_28855);
and U32233 (N_32233,N_22888,N_25557);
and U32234 (N_32234,N_24051,N_27226);
nand U32235 (N_32235,N_21662,N_22478);
nand U32236 (N_32236,N_26461,N_29385);
and U32237 (N_32237,N_28194,N_26909);
xor U32238 (N_32238,N_23238,N_25990);
and U32239 (N_32239,N_23025,N_21616);
or U32240 (N_32240,N_27803,N_25259);
xor U32241 (N_32241,N_27032,N_24582);
or U32242 (N_32242,N_25658,N_28168);
or U32243 (N_32243,N_20256,N_24855);
nand U32244 (N_32244,N_21745,N_25006);
xnor U32245 (N_32245,N_27926,N_29578);
xnor U32246 (N_32246,N_29931,N_20692);
nor U32247 (N_32247,N_27444,N_28554);
xor U32248 (N_32248,N_24613,N_26391);
and U32249 (N_32249,N_24605,N_28694);
nand U32250 (N_32250,N_29953,N_23545);
xor U32251 (N_32251,N_26835,N_21597);
or U32252 (N_32252,N_23905,N_20000);
xor U32253 (N_32253,N_23188,N_24154);
nand U32254 (N_32254,N_26939,N_29638);
xor U32255 (N_32255,N_23272,N_27129);
and U32256 (N_32256,N_24894,N_24442);
xnor U32257 (N_32257,N_22032,N_20607);
xnor U32258 (N_32258,N_23886,N_23894);
or U32259 (N_32259,N_21475,N_22726);
nand U32260 (N_32260,N_26387,N_21313);
nand U32261 (N_32261,N_23553,N_22978);
nor U32262 (N_32262,N_20588,N_29988);
and U32263 (N_32263,N_27292,N_21990);
or U32264 (N_32264,N_28639,N_26228);
xor U32265 (N_32265,N_27792,N_20515);
or U32266 (N_32266,N_25808,N_27584);
nor U32267 (N_32267,N_20051,N_27892);
and U32268 (N_32268,N_20840,N_29395);
nor U32269 (N_32269,N_22639,N_28174);
and U32270 (N_32270,N_24505,N_23368);
nand U32271 (N_32271,N_28116,N_25120);
and U32272 (N_32272,N_20966,N_24122);
or U32273 (N_32273,N_29678,N_23476);
and U32274 (N_32274,N_25348,N_20687);
and U32275 (N_32275,N_25064,N_23668);
xor U32276 (N_32276,N_27741,N_22504);
nand U32277 (N_32277,N_22420,N_27528);
nor U32278 (N_32278,N_26956,N_29473);
nor U32279 (N_32279,N_20242,N_27193);
xnor U32280 (N_32280,N_28560,N_23818);
nand U32281 (N_32281,N_20305,N_29242);
or U32282 (N_32282,N_22722,N_26750);
and U32283 (N_32283,N_27406,N_25645);
nand U32284 (N_32284,N_28432,N_25010);
xnor U32285 (N_32285,N_29374,N_27678);
nand U32286 (N_32286,N_28609,N_21222);
xor U32287 (N_32287,N_25027,N_29719);
nand U32288 (N_32288,N_26606,N_28061);
nor U32289 (N_32289,N_21595,N_22647);
nor U32290 (N_32290,N_20495,N_26876);
and U32291 (N_32291,N_23952,N_26625);
and U32292 (N_32292,N_22852,N_24389);
nand U32293 (N_32293,N_23712,N_24810);
or U32294 (N_32294,N_22745,N_20316);
and U32295 (N_32295,N_22700,N_23298);
xor U32296 (N_32296,N_24710,N_24597);
nor U32297 (N_32297,N_20137,N_29714);
or U32298 (N_32298,N_20897,N_24690);
or U32299 (N_32299,N_28418,N_28512);
nand U32300 (N_32300,N_28669,N_28401);
or U32301 (N_32301,N_23318,N_28433);
nand U32302 (N_32302,N_22517,N_29016);
or U32303 (N_32303,N_24895,N_26514);
and U32304 (N_32304,N_28860,N_24631);
or U32305 (N_32305,N_27023,N_26234);
nand U32306 (N_32306,N_25084,N_29913);
nand U32307 (N_32307,N_25705,N_23859);
xnor U32308 (N_32308,N_28456,N_25724);
and U32309 (N_32309,N_23709,N_27563);
and U32310 (N_32310,N_24718,N_26531);
nor U32311 (N_32311,N_27730,N_29841);
nand U32312 (N_32312,N_28060,N_29117);
or U32313 (N_32313,N_23597,N_24130);
and U32314 (N_32314,N_24226,N_20216);
xnor U32315 (N_32315,N_27469,N_21003);
nand U32316 (N_32316,N_22432,N_22375);
and U32317 (N_32317,N_22799,N_26964);
nor U32318 (N_32318,N_27922,N_27260);
and U32319 (N_32319,N_21869,N_27092);
nand U32320 (N_32320,N_28551,N_25331);
nor U32321 (N_32321,N_22565,N_20078);
and U32322 (N_32322,N_29290,N_29481);
or U32323 (N_32323,N_27362,N_27038);
nand U32324 (N_32324,N_21896,N_27401);
or U32325 (N_32325,N_27037,N_23537);
or U32326 (N_32326,N_28469,N_20856);
xnor U32327 (N_32327,N_24672,N_21487);
or U32328 (N_32328,N_26863,N_22482);
or U32329 (N_32329,N_25894,N_28892);
and U32330 (N_32330,N_24764,N_23121);
xnor U32331 (N_32331,N_24945,N_27403);
and U32332 (N_32332,N_20430,N_28424);
xnor U32333 (N_32333,N_24573,N_22505);
xnor U32334 (N_32334,N_25132,N_29222);
nand U32335 (N_32335,N_27070,N_21545);
nand U32336 (N_32336,N_22555,N_23096);
or U32337 (N_32337,N_25328,N_24049);
nand U32338 (N_32338,N_28020,N_25933);
nand U32339 (N_32339,N_20501,N_26747);
xor U32340 (N_32340,N_27874,N_25350);
xnor U32341 (N_32341,N_24859,N_25395);
nor U32342 (N_32342,N_27103,N_20866);
xor U32343 (N_32343,N_21526,N_29919);
and U32344 (N_32344,N_29981,N_21435);
xnor U32345 (N_32345,N_24065,N_29023);
and U32346 (N_32346,N_25456,N_28994);
nor U32347 (N_32347,N_26105,N_22686);
nand U32348 (N_32348,N_27252,N_24099);
nand U32349 (N_32349,N_23214,N_29580);
xnor U32350 (N_32350,N_21307,N_25684);
and U32351 (N_32351,N_20538,N_24633);
and U32352 (N_32352,N_26877,N_21185);
nor U32353 (N_32353,N_23586,N_29181);
and U32354 (N_32354,N_21588,N_25707);
or U32355 (N_32355,N_24887,N_25186);
nand U32356 (N_32356,N_29998,N_26590);
xor U32357 (N_32357,N_25660,N_25681);
and U32358 (N_32358,N_24204,N_29755);
nand U32359 (N_32359,N_26554,N_29209);
xor U32360 (N_32360,N_26949,N_23907);
and U32361 (N_32361,N_29652,N_29459);
xor U32362 (N_32362,N_27562,N_22337);
nand U32363 (N_32363,N_28104,N_20753);
or U32364 (N_32364,N_21331,N_27809);
nor U32365 (N_32365,N_20389,N_26033);
and U32366 (N_32366,N_25847,N_23765);
or U32367 (N_32367,N_20864,N_21430);
xnor U32368 (N_32368,N_28818,N_20033);
xor U32369 (N_32369,N_26924,N_24918);
and U32370 (N_32370,N_28185,N_24067);
or U32371 (N_32371,N_21569,N_29610);
xnor U32372 (N_32372,N_26393,N_23957);
xor U32373 (N_32373,N_27146,N_20877);
or U32374 (N_32374,N_23412,N_21899);
nor U32375 (N_32375,N_29844,N_29201);
and U32376 (N_32376,N_26599,N_23365);
and U32377 (N_32377,N_20990,N_27582);
nor U32378 (N_32378,N_25458,N_21712);
nor U32379 (N_32379,N_23557,N_24460);
or U32380 (N_32380,N_23200,N_26343);
nand U32381 (N_32381,N_22202,N_20535);
nor U32382 (N_32382,N_29066,N_27708);
and U32383 (N_32383,N_29504,N_28541);
or U32384 (N_32384,N_29344,N_22198);
nand U32385 (N_32385,N_24623,N_26748);
xor U32386 (N_32386,N_20905,N_26233);
and U32387 (N_32387,N_28317,N_20996);
and U32388 (N_32388,N_21000,N_29378);
and U32389 (N_32389,N_25708,N_28718);
and U32390 (N_32390,N_21214,N_21917);
xor U32391 (N_32391,N_25158,N_27916);
nor U32392 (N_32392,N_20705,N_26102);
xor U32393 (N_32393,N_22095,N_26394);
and U32394 (N_32394,N_22811,N_25625);
nand U32395 (N_32395,N_26982,N_23447);
and U32396 (N_32396,N_24961,N_22245);
or U32397 (N_32397,N_29371,N_24504);
or U32398 (N_32398,N_26456,N_24007);
xnor U32399 (N_32399,N_29321,N_20496);
xor U32400 (N_32400,N_29847,N_24486);
and U32401 (N_32401,N_29428,N_20362);
and U32402 (N_32402,N_28111,N_28416);
and U32403 (N_32403,N_22035,N_24255);
and U32404 (N_32404,N_26725,N_22492);
xnor U32405 (N_32405,N_28961,N_27002);
nor U32406 (N_32406,N_23173,N_22710);
nand U32407 (N_32407,N_26106,N_22479);
or U32408 (N_32408,N_23201,N_24406);
xor U32409 (N_32409,N_29253,N_23679);
and U32410 (N_32410,N_23170,N_25791);
nor U32411 (N_32411,N_28136,N_27409);
xnor U32412 (N_32412,N_24003,N_22787);
nand U32413 (N_32413,N_25978,N_26746);
and U32414 (N_32414,N_22638,N_21991);
or U32415 (N_32415,N_26869,N_23460);
nand U32416 (N_32416,N_23671,N_26849);
xnor U32417 (N_32417,N_21863,N_27459);
or U32418 (N_32418,N_27180,N_29038);
xnor U32419 (N_32419,N_22079,N_24193);
or U32420 (N_32420,N_21757,N_27056);
xnor U32421 (N_32421,N_22233,N_26171);
and U32422 (N_32422,N_28063,N_27250);
nor U32423 (N_32423,N_23399,N_29892);
xor U32424 (N_32424,N_29258,N_23833);
or U32425 (N_32425,N_20438,N_29921);
xnor U32426 (N_32426,N_25090,N_20521);
or U32427 (N_32427,N_23823,N_25381);
nor U32428 (N_32428,N_29735,N_27316);
and U32429 (N_32429,N_27544,N_27231);
xnor U32430 (N_32430,N_22205,N_28092);
xnor U32431 (N_32431,N_26157,N_26537);
xor U32432 (N_32432,N_21571,N_27328);
nor U32433 (N_32433,N_24345,N_21739);
nor U32434 (N_32434,N_29734,N_28561);
nand U32435 (N_32435,N_25836,N_29917);
or U32436 (N_32436,N_23330,N_27695);
nor U32437 (N_32437,N_21458,N_27965);
or U32438 (N_32438,N_26660,N_25976);
nor U32439 (N_32439,N_26088,N_26078);
nor U32440 (N_32440,N_28580,N_26847);
nand U32441 (N_32441,N_25415,N_21412);
xnor U32442 (N_32442,N_25603,N_26844);
nor U32443 (N_32443,N_29950,N_25747);
xnor U32444 (N_32444,N_21979,N_27706);
xor U32445 (N_32445,N_24930,N_28786);
nand U32446 (N_32446,N_23131,N_28840);
or U32447 (N_32447,N_29139,N_23656);
nor U32448 (N_32448,N_26443,N_21051);
xor U32449 (N_32449,N_23582,N_25659);
xor U32450 (N_32450,N_25436,N_24563);
nor U32451 (N_32451,N_27279,N_23095);
or U32452 (N_32452,N_21864,N_28493);
xnor U32453 (N_32453,N_26764,N_25728);
or U32454 (N_32454,N_24590,N_23533);
xor U32455 (N_32455,N_24767,N_29420);
or U32456 (N_32456,N_21501,N_26044);
nor U32457 (N_32457,N_24933,N_25975);
or U32458 (N_32458,N_23690,N_29071);
nor U32459 (N_32459,N_25225,N_23364);
nor U32460 (N_32460,N_29056,N_21763);
nand U32461 (N_32461,N_28316,N_26442);
nor U32462 (N_32462,N_27192,N_23264);
nor U32463 (N_32463,N_26740,N_24888);
and U32464 (N_32464,N_29251,N_27715);
nand U32465 (N_32465,N_27671,N_23678);
nand U32466 (N_32466,N_26450,N_25115);
and U32467 (N_32467,N_28236,N_27643);
nand U32468 (N_32468,N_23737,N_20870);
nand U32469 (N_32469,N_21016,N_23194);
xnor U32470 (N_32470,N_22053,N_29351);
xor U32471 (N_32471,N_28200,N_29974);
xor U32472 (N_32472,N_28595,N_28240);
xnor U32473 (N_32473,N_22433,N_27350);
xnor U32474 (N_32474,N_20819,N_24701);
nor U32475 (N_32475,N_22923,N_20537);
and U32476 (N_32476,N_21065,N_23523);
and U32477 (N_32477,N_23706,N_28504);
xor U32478 (N_32478,N_27625,N_26493);
or U32479 (N_32479,N_20906,N_23641);
and U32480 (N_32480,N_26568,N_23186);
and U32481 (N_32481,N_20647,N_28616);
or U32482 (N_32482,N_25872,N_23919);
or U32483 (N_32483,N_26520,N_29893);
and U32484 (N_32484,N_22528,N_27478);
nor U32485 (N_32485,N_26140,N_28474);
or U32486 (N_32486,N_29108,N_21119);
nor U32487 (N_32487,N_29942,N_23014);
nand U32488 (N_32488,N_26248,N_24975);
nor U32489 (N_32489,N_28851,N_27978);
and U32490 (N_32490,N_22522,N_27591);
nor U32491 (N_32491,N_22646,N_21797);
nand U32492 (N_32492,N_28772,N_20901);
xnor U32493 (N_32493,N_25466,N_23005);
nor U32494 (N_32494,N_28172,N_27621);
and U32495 (N_32495,N_27156,N_25582);
nor U32496 (N_32496,N_28637,N_27728);
or U32497 (N_32497,N_20473,N_23613);
nand U32498 (N_32498,N_25238,N_20617);
nand U32499 (N_32499,N_24152,N_28056);
nor U32500 (N_32500,N_24140,N_25424);
nand U32501 (N_32501,N_29365,N_28649);
nor U32502 (N_32502,N_26464,N_23732);
nand U32503 (N_32503,N_25555,N_22554);
and U32504 (N_32504,N_24377,N_29553);
xor U32505 (N_32505,N_22043,N_25289);
xor U32506 (N_32506,N_28729,N_27288);
xor U32507 (N_32507,N_28574,N_28654);
and U32508 (N_32508,N_25757,N_27821);
nor U32509 (N_32509,N_24393,N_28041);
xnor U32510 (N_32510,N_29208,N_22156);
xor U32511 (N_32511,N_22926,N_24940);
xor U32512 (N_32512,N_25404,N_29575);
or U32513 (N_32513,N_24762,N_25349);
xor U32514 (N_32514,N_27247,N_22162);
xnor U32515 (N_32515,N_29271,N_27429);
and U32516 (N_32516,N_24709,N_27000);
nand U32517 (N_32517,N_24052,N_28505);
and U32518 (N_32518,N_20881,N_28349);
nor U32519 (N_32519,N_29396,N_28797);
and U32520 (N_32520,N_26254,N_20503);
or U32521 (N_32521,N_24864,N_29404);
or U32522 (N_32522,N_24174,N_28267);
xnor U32523 (N_32523,N_21933,N_22859);
and U32524 (N_32524,N_29715,N_24620);
or U32525 (N_32525,N_24560,N_24303);
and U32526 (N_32526,N_28300,N_24851);
xnor U32527 (N_32527,N_25065,N_29348);
or U32528 (N_32528,N_28664,N_21014);
and U32529 (N_32529,N_22061,N_29943);
xnor U32530 (N_32530,N_26189,N_22197);
xor U32531 (N_32531,N_24681,N_26564);
or U32532 (N_32532,N_22965,N_25192);
and U32533 (N_32533,N_29813,N_24000);
and U32534 (N_32534,N_25364,N_29014);
nand U32535 (N_32535,N_22591,N_24381);
nor U32536 (N_32536,N_23591,N_24570);
nor U32537 (N_32537,N_28138,N_26290);
xor U32538 (N_32538,N_21913,N_26203);
or U32539 (N_32539,N_25071,N_20067);
or U32540 (N_32540,N_26820,N_26212);
or U32541 (N_32541,N_25527,N_22462);
or U32542 (N_32542,N_22681,N_22242);
and U32543 (N_32543,N_20596,N_22557);
nor U32544 (N_32544,N_20507,N_27797);
nor U32545 (N_32545,N_23697,N_23857);
nand U32546 (N_32546,N_21448,N_21698);
or U32547 (N_32547,N_20187,N_28537);
xor U32548 (N_32548,N_25993,N_29955);
nand U32549 (N_32549,N_22894,N_22142);
xor U32550 (N_32550,N_28284,N_21247);
or U32551 (N_32551,N_28171,N_27108);
nor U32552 (N_32552,N_25591,N_28340);
xor U32553 (N_32553,N_25399,N_29843);
and U32554 (N_32554,N_25295,N_29090);
and U32555 (N_32555,N_22627,N_25239);
or U32556 (N_32556,N_20108,N_26821);
nand U32557 (N_32557,N_24420,N_26602);
nor U32558 (N_32558,N_20684,N_24187);
xor U32559 (N_32559,N_24013,N_22951);
nor U32560 (N_32560,N_26583,N_29453);
and U32561 (N_32561,N_22703,N_20189);
nand U32562 (N_32562,N_23245,N_21801);
and U32563 (N_32563,N_20506,N_20053);
nand U32564 (N_32564,N_25034,N_25149);
nand U32565 (N_32565,N_27604,N_27847);
or U32566 (N_32566,N_21441,N_28114);
nand U32567 (N_32567,N_28014,N_26941);
nand U32568 (N_32568,N_26654,N_26229);
or U32569 (N_32569,N_29508,N_29740);
xor U32570 (N_32570,N_26231,N_24581);
or U32571 (N_32571,N_29384,N_21764);
xor U32572 (N_32572,N_23861,N_23159);
nor U32573 (N_32573,N_24220,N_29423);
nor U32574 (N_32574,N_27870,N_25849);
or U32575 (N_32575,N_25903,N_29817);
and U32576 (N_32576,N_26808,N_20219);
or U32577 (N_32577,N_26978,N_21514);
or U32578 (N_32578,N_20745,N_20969);
xor U32579 (N_32579,N_21181,N_22102);
nor U32580 (N_32580,N_22991,N_23397);
and U32581 (N_32581,N_27330,N_20590);
and U32582 (N_32582,N_24137,N_25736);
xnor U32583 (N_32583,N_22302,N_25868);
nor U32584 (N_32584,N_21077,N_22693);
nor U32585 (N_32585,N_23024,N_29839);
nand U32586 (N_32586,N_29096,N_22526);
and U32587 (N_32587,N_22771,N_23329);
nand U32588 (N_32588,N_20660,N_26791);
or U32589 (N_32589,N_24408,N_28117);
or U32590 (N_32590,N_28955,N_23244);
nor U32591 (N_32591,N_22495,N_25105);
nand U32592 (N_32592,N_29180,N_25723);
xnor U32593 (N_32593,N_23629,N_24182);
nor U32594 (N_32594,N_25775,N_22558);
and U32595 (N_32595,N_28080,N_22917);
or U32596 (N_32596,N_20143,N_22969);
xor U32597 (N_32597,N_20755,N_23297);
nand U32598 (N_32598,N_22931,N_23335);
xor U32599 (N_32599,N_21594,N_29425);
and U32600 (N_32600,N_26931,N_21825);
nand U32601 (N_32601,N_22658,N_21682);
nor U32602 (N_32602,N_29083,N_29147);
nor U32603 (N_32603,N_24942,N_24674);
or U32604 (N_32604,N_28534,N_22386);
and U32605 (N_32605,N_29059,N_24661);
nand U32606 (N_32606,N_26428,N_22942);
or U32607 (N_32607,N_28688,N_26139);
nor U32608 (N_32608,N_20172,N_28726);
or U32609 (N_32609,N_29089,N_27118);
and U32610 (N_32610,N_29368,N_22697);
or U32611 (N_32611,N_22221,N_27223);
or U32612 (N_32612,N_23464,N_22230);
xor U32613 (N_32613,N_21989,N_20128);
nand U32614 (N_32614,N_26703,N_26789);
nand U32615 (N_32615,N_20301,N_25329);
nand U32616 (N_32616,N_26891,N_22116);
nand U32617 (N_32617,N_29568,N_26712);
xnor U32618 (N_32618,N_26860,N_28335);
xor U32619 (N_32619,N_28755,N_21369);
nor U32620 (N_32620,N_20703,N_22841);
and U32621 (N_32621,N_23507,N_25498);
nor U32622 (N_32622,N_28931,N_20697);
and U32623 (N_32623,N_28921,N_20612);
nor U32624 (N_32624,N_26048,N_27587);
or U32625 (N_32625,N_21263,N_28857);
or U32626 (N_32626,N_29784,N_22626);
and U32627 (N_32627,N_21080,N_26751);
xnor U32628 (N_32628,N_28758,N_22412);
xnor U32629 (N_32629,N_21018,N_26904);
or U32630 (N_32630,N_25205,N_22968);
nand U32631 (N_32631,N_23735,N_20120);
nand U32632 (N_32632,N_24877,N_25322);
nand U32633 (N_32633,N_21530,N_24341);
nor U32634 (N_32634,N_21752,N_21232);
or U32635 (N_32635,N_21297,N_20325);
and U32636 (N_32636,N_21148,N_26515);
or U32637 (N_32637,N_21593,N_24113);
nand U32638 (N_32638,N_26272,N_28784);
nor U32639 (N_32639,N_21479,N_29520);
nor U32640 (N_32640,N_21082,N_23028);
nand U32641 (N_32641,N_21038,N_22515);
nand U32642 (N_32642,N_20350,N_24391);
or U32643 (N_32643,N_20805,N_23920);
xor U32644 (N_32644,N_24471,N_20514);
xor U32645 (N_32645,N_24241,N_22227);
nand U32646 (N_32646,N_24551,N_27456);
nand U32647 (N_32647,N_24172,N_22067);
nor U32648 (N_32648,N_21657,N_27008);
nor U32649 (N_32649,N_23417,N_29435);
nand U32650 (N_32650,N_29827,N_25317);
and U32651 (N_32651,N_22339,N_21383);
or U32652 (N_32652,N_24822,N_29885);
xor U32653 (N_32653,N_24845,N_29873);
or U32654 (N_32654,N_21302,N_20378);
and U32655 (N_32655,N_20264,N_27860);
xnor U32656 (N_32656,N_25842,N_27360);
and U32657 (N_32657,N_23269,N_20972);
xor U32658 (N_32658,N_26730,N_29113);
nand U32659 (N_32659,N_24717,N_23549);
or U32660 (N_32660,N_23345,N_28417);
nand U32661 (N_32661,N_21006,N_23825);
and U32662 (N_32662,N_24020,N_26874);
xor U32663 (N_32663,N_29118,N_23790);
xor U32664 (N_32664,N_28183,N_28459);
nor U32665 (N_32665,N_21186,N_29712);
or U32666 (N_32666,N_22216,N_26992);
xnor U32667 (N_32667,N_28367,N_28437);
and U32668 (N_32668,N_26871,N_20724);
or U32669 (N_32669,N_29982,N_25482);
and U32670 (N_32670,N_20173,N_25598);
xor U32671 (N_32671,N_25200,N_23967);
and U32672 (N_32672,N_27284,N_26030);
nor U32673 (N_32673,N_20974,N_20848);
and U32674 (N_32674,N_25468,N_20935);
nand U32675 (N_32675,N_29275,N_27868);
or U32676 (N_32676,N_23390,N_27304);
xnor U32677 (N_32677,N_29577,N_26843);
nand U32678 (N_32678,N_27106,N_20830);
xnor U32679 (N_32679,N_22084,N_28763);
or U32680 (N_32680,N_22373,N_25235);
xor U32681 (N_32681,N_27257,N_20962);
nor U32682 (N_32682,N_27843,N_20047);
nor U32683 (N_32683,N_27709,N_23150);
nand U32684 (N_32684,N_28558,N_29835);
nor U32685 (N_32685,N_22359,N_24609);
and U32686 (N_32686,N_29685,N_28272);
xnor U32687 (N_32687,N_28915,N_22655);
nand U32688 (N_32688,N_24104,N_22546);
nand U32689 (N_32689,N_22140,N_29527);
or U32690 (N_32690,N_29912,N_20107);
xor U32691 (N_32691,N_29417,N_29122);
or U32692 (N_32692,N_22881,N_22671);
xor U32693 (N_32693,N_23221,N_27424);
xor U32694 (N_32694,N_20699,N_24737);
nand U32695 (N_32695,N_20553,N_20779);
nor U32696 (N_32696,N_24458,N_29567);
nand U32697 (N_32697,N_20182,N_20157);
xnor U32698 (N_32698,N_24874,N_21203);
nor U32699 (N_32699,N_27805,N_24189);
nand U32700 (N_32700,N_21543,N_29782);
and U32701 (N_32701,N_25951,N_29006);
xnor U32702 (N_32702,N_24574,N_25333);
nor U32703 (N_32703,N_27751,N_25529);
xor U32704 (N_32704,N_21270,N_23054);
nand U32705 (N_32705,N_25072,N_26525);
and U32706 (N_32706,N_21608,N_22576);
or U32707 (N_32707,N_26143,N_21471);
and U32708 (N_32708,N_24632,N_27762);
nand U32709 (N_32709,N_23457,N_26492);
nor U32710 (N_32710,N_28865,N_25344);
nor U32711 (N_32711,N_26839,N_26207);
and U32712 (N_32712,N_21245,N_29256);
nor U32713 (N_32713,N_21259,N_26148);
xor U32714 (N_32714,N_21871,N_26101);
nand U32715 (N_32715,N_25745,N_22059);
nor U32716 (N_32716,N_26970,N_27097);
xor U32717 (N_32717,N_24400,N_21830);
or U32718 (N_32718,N_27568,N_21573);
or U32719 (N_32719,N_29529,N_23184);
or U32720 (N_32720,N_25321,N_20749);
xor U32721 (N_32721,N_24559,N_20376);
nor U32722 (N_32722,N_29276,N_23481);
xor U32723 (N_32723,N_25611,N_25474);
and U32724 (N_32724,N_27913,N_20147);
or U32725 (N_32725,N_29137,N_29142);
xor U32726 (N_32726,N_21246,N_29682);
nand U32727 (N_32727,N_28381,N_26174);
nor U32728 (N_32728,N_24952,N_29809);
or U32729 (N_32729,N_27303,N_25566);
or U32730 (N_32730,N_27388,N_29150);
or U32731 (N_32731,N_26954,N_22980);
nand U32732 (N_32732,N_22720,N_21098);
nor U32733 (N_32733,N_24343,N_27525);
xnor U32734 (N_32734,N_28995,N_20579);
nand U32735 (N_32735,N_24892,N_27222);
and U32736 (N_32736,N_21845,N_23740);
or U32737 (N_32737,N_26911,N_23575);
xor U32738 (N_32738,N_29661,N_22403);
nor U32739 (N_32739,N_20643,N_29588);
and U32740 (N_32740,N_21481,N_24577);
nand U32741 (N_32741,N_25664,N_24232);
and U32742 (N_32742,N_27878,N_29364);
and U32743 (N_32743,N_26621,N_27985);
nor U32744 (N_32744,N_29752,N_28973);
nand U32745 (N_32745,N_23479,N_20670);
nor U32746 (N_32746,N_28264,N_26659);
or U32747 (N_32747,N_28886,N_25045);
nor U32748 (N_32748,N_24730,N_26842);
or U32749 (N_32749,N_20426,N_27127);
xor U32750 (N_32750,N_22348,N_26985);
and U32751 (N_32751,N_21193,N_20249);
xor U32752 (N_32752,N_29997,N_28657);
and U32753 (N_32753,N_29410,N_24326);
xnor U32754 (N_32754,N_22305,N_20134);
xnor U32755 (N_32755,N_24060,N_21176);
or U32756 (N_32756,N_24451,N_26055);
and U32757 (N_32757,N_27234,N_25298);
nand U32758 (N_32758,N_27988,N_26926);
and U32759 (N_32759,N_25357,N_21924);
xnor U32760 (N_32760,N_28197,N_25281);
nand U32761 (N_32761,N_21872,N_25354);
and U32762 (N_32762,N_25636,N_24265);
or U32763 (N_32763,N_23986,N_28461);
nor U32764 (N_32764,N_23688,N_26539);
or U32765 (N_32765,N_29297,N_28916);
and U32766 (N_32766,N_28040,N_23373);
xor U32767 (N_32767,N_21469,N_27059);
xor U32768 (N_32768,N_21380,N_24227);
and U32769 (N_32769,N_26090,N_20566);
and U32770 (N_32770,N_20490,N_21538);
or U32771 (N_32771,N_29662,N_27259);
and U32772 (N_32772,N_26374,N_27808);
and U32773 (N_32773,N_23262,N_22299);
nor U32774 (N_32774,N_28871,N_27618);
nand U32775 (N_32775,N_20077,N_27145);
nand U32776 (N_32776,N_26952,N_24247);
and U32777 (N_32777,N_27339,N_22082);
or U32778 (N_32778,N_27986,N_20518);
nand U32779 (N_32779,N_25938,N_24359);
nor U32780 (N_32780,N_24117,N_27392);
nand U32781 (N_32781,N_22093,N_21610);
xor U32782 (N_32782,N_29697,N_29798);
or U32783 (N_32783,N_21497,N_23918);
nor U32784 (N_32784,N_27786,N_22487);
or U32785 (N_32785,N_29564,N_23285);
nand U32786 (N_32786,N_21661,N_22780);
xor U32787 (N_32787,N_21792,N_25831);
nand U32788 (N_32788,N_23308,N_29882);
nand U32789 (N_32789,N_25922,N_22735);
nor U32790 (N_32790,N_24357,N_23543);
nand U32791 (N_32791,N_25931,N_23750);
or U32792 (N_32792,N_24484,N_29665);
nor U32793 (N_32793,N_26209,N_25338);
nor U32794 (N_32794,N_23824,N_29403);
and U32795 (N_32795,N_23133,N_28427);
nand U32796 (N_32796,N_29736,N_27755);
nand U32797 (N_32797,N_23953,N_29062);
xor U32798 (N_32798,N_23093,N_21137);
and U32799 (N_32799,N_20041,N_25478);
and U32800 (N_32800,N_28656,N_23599);
or U32801 (N_32801,N_25245,N_26267);
nand U32802 (N_32802,N_25713,N_21744);
xnor U32803 (N_32803,N_22397,N_28870);
nor U32804 (N_32804,N_24714,N_22729);
or U32805 (N_32805,N_21876,N_29095);
or U32806 (N_32806,N_29357,N_29160);
nor U32807 (N_32807,N_20477,N_21829);
xor U32808 (N_32808,N_20510,N_23178);
nand U32809 (N_32809,N_21667,N_29058);
nand U32810 (N_32810,N_21164,N_22038);
nand U32811 (N_32811,N_20222,N_25033);
nor U32812 (N_32812,N_25437,N_28611);
nor U32813 (N_32813,N_27163,N_21346);
or U32814 (N_32814,N_25568,N_29318);
or U32815 (N_32815,N_20943,N_23943);
nand U32816 (N_32816,N_28071,N_29340);
nor U32817 (N_32817,N_22391,N_23982);
nand U32818 (N_32818,N_25042,N_23261);
nand U32819 (N_32819,N_24687,N_29533);
and U32820 (N_32820,N_26296,N_23713);
and U32821 (N_32821,N_28516,N_23082);
and U32822 (N_32822,N_21262,N_28173);
xor U32823 (N_32823,N_27408,N_24098);
and U32824 (N_32824,N_28393,N_28750);
and U32825 (N_32825,N_25271,N_22621);
nand U32826 (N_32826,N_20342,N_25703);
or U32827 (N_32827,N_27063,N_27345);
or U32828 (N_32828,N_26895,N_23890);
and U32829 (N_32829,N_29507,N_20279);
nor U32830 (N_32830,N_20359,N_20088);
nand U32831 (N_32831,N_22842,N_25843);
nand U32832 (N_32832,N_29182,N_23619);
nand U32833 (N_32833,N_24304,N_29599);
and U32834 (N_32834,N_28237,N_24380);
and U32835 (N_32835,N_22293,N_29413);
xnor U32836 (N_32836,N_27903,N_23745);
nand U32837 (N_32837,N_27828,N_26241);
and U32838 (N_32838,N_26158,N_24963);
nand U32839 (N_32839,N_23542,N_26577);
and U32840 (N_32840,N_27025,N_20372);
nand U32841 (N_32841,N_26558,N_29854);
xor U32842 (N_32842,N_26022,N_22588);
or U32843 (N_32843,N_21668,N_29171);
nor U32844 (N_32844,N_24001,N_23714);
and U32845 (N_32845,N_22278,N_25590);
xor U32846 (N_32846,N_24492,N_22189);
and U32847 (N_32847,N_20469,N_29295);
nand U32848 (N_32848,N_24449,N_27207);
nand U32849 (N_32849,N_22382,N_21528);
xnor U32850 (N_32850,N_29777,N_28853);
xor U32851 (N_32851,N_25766,N_20135);
xnor U32852 (N_32852,N_25901,N_20201);
nor U32853 (N_32853,N_24416,N_29627);
nand U32854 (N_32854,N_22719,N_25805);
nor U32855 (N_32855,N_21325,N_28877);
or U32856 (N_32856,N_21977,N_26285);
nor U32857 (N_32857,N_26562,N_27668);
or U32858 (N_32858,N_22224,N_25111);
xnor U32859 (N_32859,N_23639,N_20918);
nor U32860 (N_32860,N_20715,N_26757);
and U32861 (N_32861,N_22802,N_27652);
nor U32862 (N_32862,N_23780,N_22535);
and U32863 (N_32863,N_21405,N_27399);
xnor U32864 (N_32864,N_21590,N_20141);
nor U32865 (N_32865,N_24040,N_28120);
or U32866 (N_32866,N_28811,N_23903);
and U32867 (N_32867,N_20634,N_20936);
or U32868 (N_32868,N_22925,N_22910);
nand U32869 (N_32869,N_24194,N_26194);
or U32870 (N_32870,N_21777,N_27576);
nand U32871 (N_32871,N_22163,N_26943);
xor U32872 (N_32872,N_28533,N_20399);
and U32873 (N_32873,N_25170,N_27369);
and U32874 (N_32874,N_25280,N_28778);
and U32875 (N_32875,N_22789,N_27353);
nor U32876 (N_32876,N_23404,N_28110);
nor U32877 (N_32877,N_20862,N_28509);
nand U32878 (N_32878,N_24606,N_24920);
nand U32879 (N_32879,N_28161,N_22406);
and U32880 (N_32880,N_27861,N_20844);
or U32881 (N_32881,N_21865,N_27527);
nand U32882 (N_32882,N_24677,N_27974);
nor U32883 (N_32883,N_26053,N_26379);
nand U32884 (N_32884,N_28345,N_27178);
nand U32885 (N_32885,N_25375,N_28140);
or U32886 (N_32886,N_27182,N_22770);
and U32887 (N_32887,N_27966,N_22170);
nor U32888 (N_32888,N_24821,N_23270);
and U32889 (N_32889,N_21944,N_25391);
and U32890 (N_32890,N_26815,N_28846);
nand U32891 (N_32891,N_25382,N_20084);
nand U32892 (N_32892,N_23958,N_22024);
nor U32893 (N_32893,N_27258,N_21635);
nand U32894 (N_32894,N_20225,N_20167);
xnor U32895 (N_32895,N_20292,N_23926);
and U32896 (N_32896,N_23306,N_21574);
nand U32897 (N_32897,N_24999,N_23179);
xor U32898 (N_32898,N_27057,N_25987);
or U32899 (N_32899,N_28794,N_26311);
nand U32900 (N_32900,N_21614,N_25493);
nand U32901 (N_32901,N_29376,N_21209);
or U32902 (N_32902,N_21099,N_28141);
xnor U32903 (N_32903,N_24425,N_24997);
nor U32904 (N_32904,N_29003,N_29254);
nor U32905 (N_32905,N_27796,N_29582);
and U32906 (N_32906,N_28313,N_28556);
nand U32907 (N_32907,N_21308,N_25756);
xnor U32908 (N_32908,N_24934,N_22775);
xor U32909 (N_32909,N_20979,N_22000);
or U32910 (N_32910,N_28312,N_21956);
xnor U32911 (N_32911,N_27512,N_22656);
or U32912 (N_32912,N_28745,N_28420);
xor U32913 (N_32913,N_21927,N_20601);
and U32914 (N_32914,N_21721,N_25789);
xor U32915 (N_32915,N_27141,N_27232);
or U32916 (N_32916,N_24070,N_25840);
xor U32917 (N_32917,N_28099,N_27087);
and U32918 (N_32918,N_21997,N_22025);
and U32919 (N_32919,N_21058,N_26215);
nor U32920 (N_32920,N_20044,N_21652);
nor U32921 (N_32921,N_20406,N_24369);
nand U32922 (N_32922,N_24662,N_20454);
nor U32923 (N_32923,N_29750,N_20036);
nor U32924 (N_32924,N_22464,N_28810);
xnor U32925 (N_32925,N_22530,N_24907);
nor U32926 (N_32926,N_28571,N_21241);
or U32927 (N_32927,N_21102,N_29518);
xor U32928 (N_32928,N_21533,N_23566);
and U32929 (N_32929,N_21026,N_29010);
xor U32930 (N_32930,N_20499,N_28348);
and U32931 (N_32931,N_21968,N_26001);
and U32932 (N_32932,N_22733,N_24761);
nor U32933 (N_32933,N_21440,N_27908);
xnor U32934 (N_32934,N_20296,N_20532);
nor U32935 (N_32935,N_21587,N_29305);
nand U32936 (N_32936,N_20228,N_25489);
nor U32937 (N_32937,N_28015,N_22360);
or U32938 (N_32938,N_26047,N_29338);
nor U32939 (N_32939,N_20740,N_27557);
or U32940 (N_32940,N_22450,N_21372);
or U32941 (N_32941,N_24868,N_20937);
nand U32942 (N_32942,N_29335,N_28260);
or U32943 (N_32943,N_20324,N_24168);
or U32944 (N_32944,N_25194,N_25670);
nand U32945 (N_32945,N_27356,N_20720);
and U32946 (N_32946,N_21795,N_21226);
or U32947 (N_32947,N_23667,N_22971);
and U32948 (N_32948,N_24294,N_26923);
or U32949 (N_32949,N_22785,N_24664);
nand U32950 (N_32950,N_21542,N_25256);
nand U32951 (N_32951,N_26927,N_21936);
and U32952 (N_32952,N_27274,N_26183);
xnor U32953 (N_32953,N_20994,N_22185);
xnor U32954 (N_32954,N_27579,N_28740);
or U32955 (N_32955,N_21810,N_26691);
and U32956 (N_32956,N_22255,N_28234);
and U32957 (N_32957,N_28454,N_27072);
xnor U32958 (N_32958,N_24314,N_28324);
nand U32959 (N_32959,N_22922,N_24059);
nand U32960 (N_32960,N_23367,N_29778);
and U32961 (N_32961,N_27896,N_20152);
xnor U32962 (N_32962,N_29635,N_22239);
and U32963 (N_32963,N_27606,N_27405);
and U32964 (N_32964,N_28525,N_20645);
and U32965 (N_32965,N_28893,N_23716);
xnor U32966 (N_32966,N_22269,N_25822);
nor U32967 (N_32967,N_22727,N_24480);
nand U32968 (N_32968,N_24263,N_25480);
or U32969 (N_32969,N_27546,N_22320);
nand U32970 (N_32970,N_27311,N_28825);
and U32971 (N_32971,N_26122,N_25300);
or U32972 (N_32972,N_23622,N_20089);
and U32973 (N_32973,N_28097,N_28662);
xor U32974 (N_32974,N_20272,N_24378);
nor U32975 (N_32975,N_25101,N_22454);
or U32976 (N_32976,N_28169,N_24055);
nand U32977 (N_32977,N_20854,N_24233);
nor U32978 (N_32978,N_28193,N_26385);
and U32979 (N_32979,N_26091,N_21866);
nor U32980 (N_32980,N_20072,N_22595);
nand U32981 (N_32981,N_28186,N_28796);
nor U32982 (N_32982,N_21353,N_26611);
or U32983 (N_32983,N_26579,N_23999);
nor U32984 (N_32984,N_24437,N_27983);
nand U32985 (N_32985,N_23439,N_28617);
xor U32986 (N_32986,N_21001,N_24720);
nand U32987 (N_32987,N_22885,N_23435);
nand U32988 (N_32988,N_23386,N_21849);
and U32989 (N_32989,N_27367,N_20175);
nand U32990 (N_32990,N_20686,N_20531);
or U32991 (N_32991,N_29949,N_27477);
nand U32992 (N_32992,N_23764,N_26999);
or U32993 (N_32993,N_26111,N_24547);
xor U32994 (N_32994,N_27994,N_25008);
nand U32995 (N_32995,N_22440,N_21672);
and U32996 (N_32996,N_23433,N_22114);
xor U32997 (N_32997,N_27147,N_26594);
xnor U32998 (N_32998,N_25592,N_22601);
nand U32999 (N_32999,N_24927,N_29765);
and U33000 (N_33000,N_20583,N_20702);
nand U33001 (N_33001,N_22845,N_22346);
xor U33002 (N_33002,N_25648,N_26637);
or U33003 (N_33003,N_28984,N_23625);
and U33004 (N_33004,N_24045,N_23694);
xnor U33005 (N_33005,N_20680,N_29135);
nor U33006 (N_33006,N_26692,N_24941);
or U33007 (N_33007,N_24103,N_23630);
and U33008 (N_33008,N_25016,N_20344);
nand U33009 (N_33009,N_20613,N_27583);
nor U33010 (N_33010,N_25589,N_27322);
xor U33011 (N_33011,N_28273,N_28155);
nand U33012 (N_33012,N_21875,N_23968);
and U33013 (N_33013,N_25270,N_26890);
and U33014 (N_33014,N_29621,N_25655);
nor U33015 (N_33015,N_20823,N_25797);
and U33016 (N_33016,N_27463,N_22738);
xor U33017 (N_33017,N_21385,N_22222);
and U33018 (N_33018,N_26002,N_25512);
and U33019 (N_33019,N_29647,N_29768);
nor U33020 (N_33020,N_29614,N_23910);
or U33021 (N_33021,N_28703,N_23166);
xor U33022 (N_33022,N_20628,N_28780);
xnor U33023 (N_33023,N_23223,N_29450);
xnor U33024 (N_33024,N_22428,N_28320);
xnor U33025 (N_33025,N_20759,N_25173);
xor U33026 (N_33026,N_27734,N_28413);
and U33027 (N_33027,N_20215,N_25672);
xor U33028 (N_33028,N_20221,N_27801);
nor U33029 (N_33029,N_22870,N_22806);
or U33030 (N_33030,N_29794,N_22182);
xor U33031 (N_33031,N_28735,N_24305);
and U33032 (N_33032,N_21537,N_27887);
and U33033 (N_33033,N_29088,N_27030);
or U33034 (N_33034,N_27121,N_23674);
or U33035 (N_33035,N_24462,N_26494);
nor U33036 (N_33036,N_23353,N_21515);
xnor U33037 (N_33037,N_23380,N_22850);
and U33038 (N_33038,N_24962,N_22708);
nand U33039 (N_33039,N_25443,N_25816);
nor U33040 (N_33040,N_22075,N_27430);
or U33041 (N_33041,N_28261,N_28101);
or U33042 (N_33042,N_29225,N_21264);
nor U33043 (N_33043,N_23800,N_20327);
xor U33044 (N_33044,N_29402,N_23389);
nand U33045 (N_33045,N_23455,N_29332);
and U33046 (N_33046,N_29781,N_21178);
nor U33047 (N_33047,N_22307,N_26478);
xor U33048 (N_33048,N_27774,N_23636);
xnor U33049 (N_33049,N_27703,N_24301);
xnor U33050 (N_33050,N_22963,N_24516);
or U33051 (N_33051,N_24657,N_29082);
xor U33052 (N_33052,N_20985,N_26369);
xor U33053 (N_33053,N_29112,N_20066);
nor U33054 (N_33054,N_20403,N_23680);
nand U33055 (N_33055,N_23305,N_26435);
and U33056 (N_33056,N_21069,N_24148);
nor U33057 (N_33057,N_20593,N_27656);
xor U33058 (N_33058,N_25471,N_24665);
or U33059 (N_33059,N_26704,N_21617);
or U33060 (N_33060,N_26807,N_28126);
xor U33061 (N_33061,N_22408,N_26563);
xnor U33062 (N_33062,N_26367,N_23403);
xnor U33063 (N_33063,N_22724,N_29214);
xnor U33064 (N_33064,N_28949,N_27128);
xnor U33065 (N_33065,N_24958,N_20610);
xnor U33066 (N_33066,N_26340,N_23359);
nand U33067 (N_33067,N_20810,N_21011);
and U33068 (N_33068,N_29625,N_25913);
and U33069 (N_33069,N_22459,N_29184);
nand U33070 (N_33070,N_25007,N_25667);
nor U33071 (N_33071,N_27039,N_22480);
xnor U33072 (N_33072,N_29196,N_21127);
xor U33073 (N_33073,N_23396,N_22797);
or U33074 (N_33074,N_22955,N_24972);
xnor U33075 (N_33075,N_23504,N_28165);
nand U33076 (N_33076,N_20015,N_21823);
xor U33077 (N_33077,N_23110,N_23708);
xnor U33078 (N_33078,N_22071,N_22932);
xnor U33079 (N_33079,N_27660,N_29800);
xnor U33080 (N_33080,N_22124,N_26433);
nand U33081 (N_33081,N_25126,N_27197);
and U33082 (N_33082,N_28382,N_23515);
nand U33083 (N_33083,N_21772,N_20777);
nor U33084 (N_33084,N_28631,N_25977);
nand U33085 (N_33085,N_29422,N_25690);
xnor U33086 (N_33086,N_21273,N_23485);
nand U33087 (N_33087,N_21113,N_27638);
nor U33088 (N_33088,N_29613,N_20487);
nand U33089 (N_33089,N_21601,N_25419);
and U33090 (N_33090,N_26439,N_21690);
or U33091 (N_33091,N_24966,N_22314);
or U33092 (N_33092,N_29266,N_25628);
and U33093 (N_33093,N_20731,N_28113);
and U33094 (N_33094,N_24683,N_28328);
or U33095 (N_33095,N_24550,N_23063);
nand U33096 (N_33096,N_25223,N_25968);
and U33097 (N_33097,N_22855,N_22080);
or U33098 (N_33098,N_25730,N_25165);
and U33099 (N_33099,N_26971,N_22886);
xnor U33100 (N_33100,N_26853,N_28224);
xnor U33101 (N_33101,N_21333,N_28696);
or U33102 (N_33102,N_27082,N_22045);
and U33103 (N_33103,N_27393,N_26440);
and U33104 (N_33104,N_26154,N_27549);
nand U33105 (N_33105,N_26702,N_28709);
nor U33106 (N_33106,N_29257,N_27595);
xor U33107 (N_33107,N_28630,N_22815);
nand U33108 (N_33108,N_26614,N_22816);
or U33109 (N_33109,N_26670,N_22860);
and U33110 (N_33110,N_29328,N_20235);
xor U33111 (N_33111,N_26489,N_27475);
nor U33112 (N_33112,N_22214,N_20451);
xor U33113 (N_33113,N_21166,N_28095);
and U33114 (N_33114,N_28479,N_23867);
and U33115 (N_33115,N_20999,N_29524);
xnor U33116 (N_33116,N_23411,N_20396);
or U33117 (N_33117,N_21258,N_24132);
nor U33118 (N_33118,N_26772,N_27007);
or U33119 (N_33119,N_27022,N_20622);
and U33120 (N_33120,N_29636,N_27906);
or U33121 (N_33121,N_21283,N_25965);
and U33122 (N_33122,N_25870,N_21743);
nor U33123 (N_33123,N_22674,N_27040);
xor U33124 (N_33124,N_26685,N_29092);
nor U33125 (N_33125,N_25074,N_29769);
nand U33126 (N_33126,N_21040,N_25063);
or U33127 (N_33127,N_25484,N_22496);
nand U33128 (N_33128,N_26937,N_28906);
nor U33129 (N_33129,N_25794,N_27302);
and U33130 (N_33130,N_22933,N_21281);
nand U33131 (N_33131,N_20208,N_27335);
nor U33132 (N_33132,N_26773,N_28777);
nor U33133 (N_33133,N_28791,N_25562);
nor U33134 (N_33134,N_20899,N_20609);
nor U33135 (N_33135,N_21165,N_24022);
or U33136 (N_33136,N_20432,N_26397);
or U33137 (N_33137,N_21477,N_23216);
or U33138 (N_33138,N_24155,N_21976);
nand U33139 (N_33139,N_28843,N_28494);
nand U33140 (N_33140,N_29952,N_29968);
nand U33141 (N_33141,N_21842,N_21520);
or U33142 (N_33142,N_29696,N_29312);
and U33143 (N_33143,N_21647,N_21508);
nor U33144 (N_33144,N_29219,N_23925);
nand U33145 (N_33145,N_23428,N_23525);
nand U33146 (N_33146,N_20729,N_27435);
and U33147 (N_33147,N_23471,N_22374);
nor U33148 (N_33148,N_26167,N_27297);
nand U33149 (N_33149,N_20651,N_28965);
xor U33150 (N_33150,N_21211,N_28051);
or U33151 (N_33151,N_23973,N_26003);
or U33152 (N_33152,N_27420,N_27537);
and U33153 (N_33153,N_20393,N_20471);
nand U33154 (N_33154,N_25294,N_21730);
nand U33155 (N_33155,N_21337,N_28677);
and U33156 (N_33156,N_20902,N_22512);
nand U33157 (N_33157,N_28804,N_24641);
and U33158 (N_33158,N_21197,N_24830);
nand U33159 (N_33159,N_21986,N_27329);
and U33160 (N_33160,N_26845,N_20273);
or U33161 (N_33161,N_21220,N_24564);
and U33162 (N_33162,N_22166,N_23733);
and U33163 (N_33163,N_20150,N_27255);
xor U33164 (N_33164,N_26466,N_22040);
xnor U33165 (N_33165,N_29414,N_24741);
xor U33166 (N_33166,N_21560,N_24430);
and U33167 (N_33167,N_27848,N_21499);
nand U33168 (N_33168,N_26028,N_28612);
and U33169 (N_33169,N_24879,N_21049);
and U33170 (N_33170,N_23762,N_26744);
or U33171 (N_33171,N_27073,N_20714);
or U33172 (N_33172,N_21802,N_20416);
nor U33173 (N_33173,N_22976,N_21356);
and U33174 (N_33174,N_27175,N_26163);
or U33175 (N_33175,N_24529,N_20986);
nand U33176 (N_33176,N_21687,N_28831);
nor U33177 (N_33177,N_24164,N_28024);
nand U33178 (N_33178,N_21300,N_21716);
and U33179 (N_33179,N_21250,N_26266);
nand U33180 (N_33180,N_27623,N_21341);
xor U33181 (N_33181,N_24044,N_21221);
and U33182 (N_33182,N_22577,N_23229);
or U33183 (N_33183,N_26351,N_28458);
and U33184 (N_33184,N_23954,N_20481);
or U33185 (N_33185,N_23372,N_22411);
nand U33186 (N_33186,N_28700,N_23247);
or U33187 (N_33187,N_22506,N_29759);
or U33188 (N_33188,N_25221,N_28695);
and U33189 (N_33189,N_25862,N_24161);
or U33190 (N_33190,N_22176,N_24351);
and U33191 (N_33191,N_29976,N_23415);
xnor U33192 (N_33192,N_26701,N_25610);
nand U33193 (N_33193,N_26559,N_24998);
and U33194 (N_33194,N_27309,N_29617);
nor U33195 (N_33195,N_28281,N_20276);
nor U33196 (N_33196,N_27669,N_27839);
nand U33197 (N_33197,N_29656,N_23898);
xnor U33198 (N_33198,N_24669,N_28765);
nor U33199 (N_33199,N_27912,N_27905);
nand U33200 (N_33200,N_21215,N_24867);
xor U33201 (N_33201,N_20318,N_29352);
and U33202 (N_33202,N_28733,N_22476);
nand U33203 (N_33203,N_28769,N_22363);
nor U33204 (N_33204,N_20540,N_28661);
nand U33205 (N_33205,N_22001,N_24649);
or U33206 (N_33206,N_26424,N_22915);
nand U33207 (N_33207,N_25500,N_29615);
xnor U33208 (N_33208,N_28866,N_20947);
nand U33209 (N_33209,N_25835,N_28005);
xor U33210 (N_33210,N_22718,N_27340);
nor U33211 (N_33211,N_27268,N_23742);
and U33212 (N_33212,N_26330,N_21765);
nand U33213 (N_33213,N_23663,N_27899);
nand U33214 (N_33214,N_24293,N_24801);
and U33215 (N_33215,N_26378,N_23689);
or U33216 (N_33216,N_24771,N_29350);
xnor U33217 (N_33217,N_23099,N_24331);
nand U33218 (N_33218,N_23601,N_27829);
nor U33219 (N_33219,N_29970,N_29695);
nand U33220 (N_33220,N_26293,N_24426);
or U33221 (N_33221,N_20949,N_21496);
xnor U33222 (N_33222,N_29884,N_21916);
or U33223 (N_33223,N_25272,N_29308);
nor U33224 (N_33224,N_25750,N_26273);
and U33225 (N_33225,N_24768,N_22688);
or U33226 (N_33226,N_27902,N_22937);
nor U33227 (N_33227,N_26477,N_28069);
and U33228 (N_33228,N_23642,N_20421);
and U33229 (N_33229,N_28645,N_26259);
and U33230 (N_33230,N_24481,N_21156);
nor U33231 (N_33231,N_20368,N_27151);
and U33232 (N_33232,N_27321,N_20982);
and U33233 (N_33233,N_26358,N_26479);
and U33234 (N_33234,N_20443,N_27581);
nor U33235 (N_33235,N_27596,N_21544);
and U33236 (N_33236,N_27910,N_29380);
nand U33237 (N_33237,N_21646,N_20338);
xnor U33238 (N_33238,N_27485,N_21919);
xor U33239 (N_33239,N_24837,N_23168);
nor U33240 (N_33240,N_24083,N_26423);
nand U33241 (N_33241,N_20429,N_24209);
xor U33242 (N_33242,N_27048,N_27214);
xor U33243 (N_33243,N_25856,N_27811);
xnor U33244 (N_33244,N_27136,N_27191);
or U33245 (N_33245,N_20014,N_27692);
nand U33246 (N_33246,N_20034,N_26879);
nor U33247 (N_33247,N_27391,N_25249);
or U33248 (N_33248,N_21180,N_22212);
nand U33249 (N_33249,N_29084,N_29743);
and U33250 (N_33250,N_20117,N_25702);
xor U33251 (N_33251,N_21066,N_23570);
and U33252 (N_33252,N_26601,N_29757);
nor U33253 (N_33253,N_23782,N_26327);
and U33254 (N_33254,N_27693,N_22347);
nor U33255 (N_33255,N_21238,N_29929);
or U33256 (N_33256,N_21486,N_21966);
nand U33257 (N_33257,N_21257,N_23969);
and U33258 (N_33258,N_27489,N_23538);
xnor U33259 (N_33259,N_29460,N_24224);
xor U33260 (N_33260,N_21136,N_26516);
or U33261 (N_33261,N_22986,N_23569);
nand U33262 (N_33262,N_26675,N_29566);
or U33263 (N_33263,N_25085,N_21426);
nand U33264 (N_33264,N_28159,N_26341);
or U33265 (N_33265,N_23073,N_25515);
nand U33266 (N_33266,N_23751,N_25320);
xor U33267 (N_33267,N_22281,N_25029);
and U33268 (N_33268,N_28952,N_25918);
nand U33269 (N_33269,N_27679,N_28498);
nor U33270 (N_33270,N_29729,N_20115);
nor U33271 (N_33271,N_25252,N_21260);
nor U33272 (N_33272,N_22267,N_25620);
nand U33273 (N_33273,N_25761,N_22542);
nand U33274 (N_33274,N_24598,N_25177);
or U33275 (N_33275,N_24253,N_21787);
and U33276 (N_33276,N_28299,N_23858);
nor U33277 (N_33277,N_21290,N_22755);
xnor U33278 (N_33278,N_21644,N_27044);
xor U33279 (N_33279,N_21256,N_20343);
and U33280 (N_33280,N_22892,N_24493);
and U33281 (N_33281,N_28034,N_25884);
nor U33282 (N_33282,N_27326,N_26304);
nor U33283 (N_33283,N_25575,N_20461);
xor U33284 (N_33284,N_21582,N_25291);
nand U33285 (N_33285,N_25615,N_23431);
or U33286 (N_33286,N_24295,N_20312);
nor U33287 (N_33287,N_21505,N_29287);
nand U33288 (N_33288,N_24835,N_29960);
nand U33289 (N_33289,N_24195,N_23934);
or U33290 (N_33290,N_29279,N_25785);
nand U33291 (N_33291,N_21521,N_20657);
nor U33292 (N_33292,N_25962,N_29948);
nor U33293 (N_33293,N_25510,N_22112);
and U33294 (N_33294,N_29602,N_28137);
or U33295 (N_33295,N_22297,N_25465);
nand U33296 (N_33296,N_22134,N_22559);
xor U33297 (N_33297,N_24200,N_27779);
xor U33298 (N_33298,N_21438,N_22296);
nor U33299 (N_33299,N_25936,N_29412);
nor U33300 (N_33300,N_25523,N_29946);
nor U33301 (N_33301,N_28975,N_29667);
nand U33302 (N_33302,N_27497,N_26695);
nor U33303 (N_33303,N_27901,N_23949);
nand U33304 (N_33304,N_26916,N_20151);
xor U33305 (N_33305,N_28698,N_29876);
or U33306 (N_33306,N_27871,N_24601);
nand U33307 (N_33307,N_24021,N_26998);
nor U33308 (N_33308,N_21557,N_25916);
nor U33309 (N_33309,N_22946,N_28238);
or U33310 (N_33310,N_26150,N_28519);
or U33311 (N_33311,N_20055,N_23038);
xnor U33312 (N_33312,N_24947,N_20018);
xor U33313 (N_33313,N_26571,N_23255);
nor U33314 (N_33314,N_24588,N_26623);
nor U33315 (N_33315,N_26132,N_22813);
and U33316 (N_33316,N_21227,N_24676);
and U33317 (N_33317,N_25473,N_25463);
nand U33318 (N_33318,N_28894,N_22385);
xnor U33319 (N_33319,N_29261,N_25671);
or U33320 (N_33320,N_22880,N_22985);
and U33321 (N_33321,N_25199,N_29995);
nand U33322 (N_33322,N_29978,N_26983);
xnor U33323 (N_33323,N_22834,N_21903);
xnor U33324 (N_33324,N_26556,N_22665);
nand U33325 (N_33325,N_21484,N_27566);
nand U33326 (N_33326,N_20798,N_21071);
xor U33327 (N_33327,N_24978,N_21665);
or U33328 (N_33328,N_25241,N_20239);
nand U33329 (N_33329,N_20940,N_28833);
or U33330 (N_33330,N_21955,N_27439);
or U33331 (N_33331,N_21524,N_29436);
nor U33332 (N_33332,N_29632,N_23985);
and U33333 (N_33333,N_23880,N_27013);
xor U33334 (N_33334,N_29293,N_26221);
nand U33335 (N_33335,N_25048,N_26885);
xnor U33336 (N_33336,N_26013,N_23338);
nand U33337 (N_33337,N_23066,N_22442);
or U33338 (N_33338,N_23783,N_20548);
or U33339 (N_33339,N_21416,N_26899);
xor U33340 (N_33340,N_29785,N_24995);
xnor U33341 (N_33341,N_20209,N_25459);
or U33342 (N_33342,N_23796,N_25213);
xor U33343 (N_33343,N_21115,N_23659);
nand U33344 (N_33344,N_20824,N_27338);
and U33345 (N_33345,N_22485,N_27533);
xor U33346 (N_33346,N_24883,N_25087);
xnor U33347 (N_33347,N_28419,N_24797);
nand U33348 (N_33348,N_21146,N_26581);
and U33349 (N_33349,N_20064,N_23908);
or U33350 (N_33350,N_29455,N_25335);
xor U33351 (N_33351,N_27398,N_20618);
nor U33352 (N_33352,N_24655,N_26894);
xnor U33353 (N_33353,N_23510,N_28153);
or U33354 (N_33354,N_24713,N_21123);
or U33355 (N_33355,N_20774,N_29278);
and U33356 (N_33356,N_28800,N_24415);
nand U33357 (N_33357,N_21941,N_27422);
nand U33358 (N_33358,N_23120,N_28301);
and U33359 (N_33359,N_20851,N_27071);
or U33360 (N_33360,N_29506,N_26485);
nand U33361 (N_33361,N_27686,N_26145);
nor U33362 (N_33362,N_25548,N_24025);
or U33363 (N_33363,N_28483,N_22829);
nand U33364 (N_33364,N_20728,N_23148);
or U33365 (N_33365,N_20199,N_27219);
or U33366 (N_33366,N_26032,N_20025);
xnor U33367 (N_33367,N_25858,N_29924);
or U33368 (N_33368,N_25767,N_24721);
nand U33369 (N_33369,N_24114,N_20080);
nor U33370 (N_33370,N_22223,N_22152);
xor U33371 (N_33371,N_29282,N_27492);
or U33372 (N_33372,N_20309,N_21619);
nand U33373 (N_33373,N_20736,N_28712);
nor U33374 (N_33374,N_20340,N_26617);
nor U33375 (N_33375,N_28442,N_22388);
nor U33376 (N_33376,N_20386,N_20099);
and U33377 (N_33377,N_20142,N_20096);
or U33378 (N_33378,N_27765,N_21434);
nand U33379 (N_33379,N_27745,N_26813);
or U33380 (N_33380,N_20231,N_22592);
xnor U33381 (N_33381,N_28727,N_26632);
or U33382 (N_33382,N_25726,N_26836);
xnor U33383 (N_33383,N_28898,N_29650);
nor U33384 (N_33384,N_27628,N_27327);
nand U33385 (N_33385,N_23416,N_27588);
nand U33386 (N_33386,N_29116,N_22158);
nand U33387 (N_33387,N_22467,N_27077);
or U33388 (N_33388,N_20112,N_24494);
and U33389 (N_33389,N_25520,N_25080);
xor U33390 (N_33390,N_21017,N_22276);
nor U33391 (N_33391,N_25421,N_27629);
nand U33392 (N_33392,N_29346,N_27476);
and U33393 (N_33393,N_29753,N_25939);
and U33394 (N_33394,N_24884,N_21926);
xor U33395 (N_33395,N_20875,N_22617);
and U33396 (N_33396,N_28593,N_21436);
nor U33397 (N_33397,N_23407,N_29306);
nor U33398 (N_33398,N_24643,N_21005);
and U33399 (N_33399,N_23929,N_29494);
nor U33400 (N_33400,N_29601,N_27723);
xor U33401 (N_33401,N_21892,N_20486);
and U33402 (N_33402,N_24466,N_25117);
xnor U33403 (N_33403,N_21090,N_25184);
nand U33404 (N_33404,N_22107,N_22610);
nor U33405 (N_33405,N_25339,N_28799);
nand U33406 (N_33406,N_23328,N_21117);
and U33407 (N_33407,N_21746,N_25159);
xnor U33408 (N_33408,N_20065,N_20730);
or U33409 (N_33409,N_29726,N_21881);
xor U33410 (N_33410,N_23236,N_25911);
or U33411 (N_33411,N_25394,N_28302);
nor U33412 (N_33412,N_22973,N_26587);
nor U33413 (N_33413,N_29247,N_23754);
nor U33414 (N_33414,N_28544,N_27253);
and U33415 (N_33415,N_22634,N_23596);
nand U33416 (N_33416,N_25573,N_25453);
nand U33417 (N_33417,N_24354,N_25038);
or U33418 (N_33418,N_29723,N_22366);
xnor U33419 (N_33419,N_28936,N_20497);
nand U33420 (N_33420,N_21167,N_27654);
nor U33421 (N_33421,N_29388,N_28250);
xor U33422 (N_33422,N_20968,N_26811);
nand U33423 (N_33423,N_22398,N_28476);
or U33424 (N_33424,N_21474,N_26335);
nor U33425 (N_33425,N_21691,N_22203);
nor U33426 (N_33426,N_26210,N_29127);
nand U33427 (N_33427,N_24068,N_28492);
xor U33428 (N_33428,N_27763,N_23617);
nand U33429 (N_33429,N_29544,N_26973);
and U33430 (N_33430,N_20489,N_29013);
and U33431 (N_33431,N_27603,N_24450);
and U33432 (N_33432,N_24456,N_24046);
nor U33433 (N_33433,N_23436,N_26190);
nor U33434 (N_33434,N_25953,N_27927);
xor U33435 (N_33435,N_21703,N_27454);
and U33436 (N_33436,N_21670,N_28564);
xor U33437 (N_33437,N_29705,N_22133);
or U33438 (N_33438,N_29270,N_29326);
xor U33439 (N_33439,N_25296,N_23786);
or U33440 (N_33440,N_25114,N_26913);
or U33441 (N_33441,N_24281,N_23147);
nor U33442 (N_33442,N_26491,N_26243);
nand U33443 (N_33443,N_21154,N_22996);
or U33444 (N_33444,N_26366,N_21975);
xor U33445 (N_33445,N_21972,N_28875);
or U33446 (N_33446,N_28659,N_29918);
or U33447 (N_33447,N_24026,N_26743);
or U33448 (N_33448,N_20315,N_25806);
and U33449 (N_33449,N_21693,N_22633);
nor U33450 (N_33450,N_23971,N_23293);
xor U33451 (N_33451,N_21552,N_23555);
or U33452 (N_33452,N_20314,N_29138);
nand U33453 (N_33453,N_20835,N_26412);
xor U33454 (N_33454,N_20366,N_22111);
and U33455 (N_33455,N_27853,N_20436);
or U33456 (N_33456,N_26141,N_26596);
nand U33457 (N_33457,N_23977,N_22615);
or U33458 (N_33458,N_24243,N_26214);
xor U33459 (N_33459,N_27265,N_23127);
xor U33460 (N_33460,N_27474,N_21660);
and U33461 (N_33461,N_24732,N_29927);
and U33462 (N_33462,N_29019,N_27955);
or U33463 (N_33463,N_23299,N_29901);
or U33464 (N_33464,N_22128,N_27530);
or U33465 (N_33465,N_25873,N_26275);
nand U33466 (N_33466,N_27697,N_21742);
nor U33467 (N_33467,N_27712,N_28147);
nor U33468 (N_33468,N_20558,N_21421);
nor U33469 (N_33469,N_22394,N_27567);
and U33470 (N_33470,N_24251,N_28680);
nand U33471 (N_33471,N_21902,N_22947);
xor U33472 (N_33472,N_23098,N_21598);
nand U33473 (N_33473,N_27607,N_21411);
nand U33474 (N_33474,N_27665,N_28891);
nor U33475 (N_33475,N_23862,N_28112);
and U33476 (N_33476,N_22817,N_23375);
and U33477 (N_33477,N_20502,N_26684);
nand U33478 (N_33478,N_23801,N_21654);
or U33479 (N_33479,N_28563,N_23279);
xor U33480 (N_33480,N_21032,N_20260);
nand U33481 (N_33481,N_21401,N_21201);
xnor U33482 (N_33482,N_28129,N_28094);
xnor U33483 (N_33483,N_23710,N_20576);
nor U33484 (N_33484,N_23441,N_20907);
and U33485 (N_33485,N_22336,N_23036);
or U33486 (N_33486,N_27836,N_21701);
nand U33487 (N_33487,N_28988,N_24627);
nor U33488 (N_33488,N_24578,N_23176);
and U33489 (N_33489,N_29240,N_21254);
nand U33490 (N_33490,N_20778,N_28026);
xor U33491 (N_33491,N_25169,N_22857);
nand U33492 (N_33492,N_24860,N_23037);
nand U33493 (N_33493,N_22372,N_22524);
nand U33494 (N_33494,N_26553,N_28827);
nand U33495 (N_33495,N_25734,N_25631);
nand U33496 (N_33496,N_20428,N_25554);
and U33497 (N_33497,N_21128,N_29070);
nor U33498 (N_33498,N_29803,N_21850);
xnor U33499 (N_33499,N_26225,N_27894);
xnor U33500 (N_33500,N_28179,N_28756);
nor U33501 (N_33501,N_25037,N_24931);
nor U33502 (N_33502,N_22342,N_24948);
and U33503 (N_33503,N_22730,N_28354);
xor U33504 (N_33504,N_27858,N_27536);
nand U33505 (N_33505,N_28501,N_26077);
nor U33506 (N_33506,N_29802,N_26240);
nor U33507 (N_33507,N_21355,N_20754);
nor U33508 (N_33508,N_27240,N_25157);
and U33509 (N_33509,N_25308,N_27516);
xnor U33510 (N_33510,N_28290,N_22443);
xor U33511 (N_33511,N_29193,N_27502);
nor U33512 (N_33512,N_29102,N_27945);
or U33513 (N_33513,N_22323,N_25752);
xor U33514 (N_33514,N_25374,N_20793);
nor U33515 (N_33515,N_24925,N_22423);
xnor U33516 (N_33516,N_23654,N_26235);
and U33517 (N_33517,N_22642,N_28704);
or U33518 (N_33518,N_28287,N_25886);
xor U33519 (N_33519,N_22488,N_24439);
xor U33520 (N_33520,N_25559,N_24048);
and U33521 (N_33521,N_29561,N_24213);
or U33522 (N_33522,N_24795,N_25823);
and U33523 (N_33523,N_25604,N_22155);
nand U33524 (N_33524,N_27186,N_24225);
nor U33525 (N_33525,N_20993,N_21237);
and U33526 (N_33526,N_28394,N_27934);
xnor U33527 (N_33527,N_28239,N_26585);
and U33528 (N_33528,N_27522,N_29255);
nand U33529 (N_33529,N_27704,N_25711);
nand U33530 (N_33530,N_27344,N_20873);
xnor U33531 (N_33531,N_29366,N_23719);
and U33532 (N_33532,N_21423,N_29608);
and U33533 (N_33533,N_24455,N_27586);
nand U33534 (N_33534,N_25315,N_21531);
and U33535 (N_33535,N_20922,N_22069);
xor U33536 (N_33536,N_20547,N_24926);
and U33537 (N_33537,N_27547,N_27140);
and U33538 (N_33538,N_23362,N_28346);
nand U33539 (N_33539,N_23097,N_29536);
and U33540 (N_33540,N_26460,N_27598);
or U33541 (N_33541,N_28550,N_21373);
and U33542 (N_33542,N_21453,N_24760);
or U33543 (N_33543,N_28325,N_27065);
nor U33544 (N_33544,N_21988,N_26857);
and U33545 (N_33545,N_21208,N_25715);
nand U33546 (N_33546,N_20520,N_29032);
nor U33547 (N_33547,N_22578,N_22879);
and U33548 (N_33548,N_23947,N_27752);
xnor U33549 (N_33549,N_27050,N_20236);
nand U33550 (N_33550,N_28946,N_22807);
nor U33551 (N_33551,N_20100,N_25060);
xor U33552 (N_33552,N_20038,N_25403);
nand U33553 (N_33553,N_21679,N_22271);
nand U33554 (N_33554,N_25416,N_21329);
xnor U33555 (N_33555,N_25131,N_27950);
and U33556 (N_33556,N_28842,N_26739);
or U33557 (N_33557,N_29418,N_24639);
or U33558 (N_33558,N_28269,N_22890);
nand U33559 (N_33559,N_25880,N_27198);
or U33560 (N_33560,N_23080,N_24809);
or U33561 (N_33561,N_23941,N_29232);
nand U33562 (N_33562,N_23059,N_20516);
or U33563 (N_33563,N_26969,N_21555);
nor U33564 (N_33564,N_20223,N_23062);
or U33565 (N_33565,N_23209,N_21857);
nor U33566 (N_33566,N_26352,N_26126);
or U33567 (N_33567,N_22543,N_22475);
xnor U33568 (N_33568,N_21396,N_28829);
xnor U33569 (N_33569,N_26734,N_23026);
nor U33570 (N_33570,N_24206,N_20230);
and U33571 (N_33571,N_24898,N_20828);
or U33572 (N_33572,N_20808,N_26063);
nand U33573 (N_33573,N_22560,N_29311);
xor U33574 (N_33574,N_25945,N_21183);
xor U33575 (N_33575,N_26287,N_27831);
and U33576 (N_33576,N_29145,N_22002);
and U33577 (N_33577,N_22054,N_20270);
or U33578 (N_33578,N_22486,N_26498);
nor U33579 (N_33579,N_28837,N_29304);
xor U33580 (N_33580,N_28601,N_29177);
and U33581 (N_33581,N_29584,N_29022);
xor U33582 (N_33582,N_26854,N_25881);
nor U33583 (N_33583,N_23374,N_24076);
nor U33584 (N_33584,N_23699,N_27904);
and U33585 (N_33585,N_24121,N_28464);
nand U33586 (N_33586,N_24276,N_22379);
nor U33587 (N_33587,N_20792,N_24418);
and U33588 (N_33588,N_26024,N_20006);
xor U33589 (N_33589,N_27943,N_25201);
xnor U33590 (N_33590,N_29868,N_27451);
xor U33591 (N_33591,N_23191,N_27973);
nand U33592 (N_33592,N_28803,N_29954);
and U33593 (N_33593,N_29713,N_20953);
or U33594 (N_33594,N_23259,N_29733);
nor U33595 (N_33595,N_28380,N_28125);
or U33596 (N_33596,N_25682,N_20444);
and U33597 (N_33597,N_28913,N_29780);
nor U33598 (N_33598,N_26638,N_22473);
nand U33599 (N_33599,N_27592,N_20352);
and U33600 (N_33600,N_27612,N_22268);
nand U33601 (N_33601,N_24707,N_29941);
nor U33602 (N_33602,N_26758,N_22383);
nor U33603 (N_33603,N_25774,N_22645);
or U33604 (N_33604,N_23081,N_29822);
and U33605 (N_33605,N_28225,N_28604);
or U33606 (N_33606,N_25429,N_26467);
and U33607 (N_33607,N_25146,N_25360);
or U33608 (N_33608,N_28868,N_20598);
and U33609 (N_33609,N_20424,N_23185);
and U33610 (N_33610,N_23534,N_27060);
or U33611 (N_33611,N_25325,N_23348);
and U33612 (N_33612,N_29020,N_26300);
xor U33613 (N_33613,N_23065,N_25679);
nor U33614 (N_33614,N_20431,N_23848);
nand U33615 (N_33615,N_29528,N_20377);
xnor U33616 (N_33616,N_25618,N_21357);
nand U33617 (N_33617,N_27172,N_28806);
or U33618 (N_33618,N_26375,N_20764);
nand U33619 (N_33619,N_28838,N_20825);
nor U33620 (N_33620,N_23488,N_20492);
xor U33621 (N_33621,N_21906,N_26883);
nand U33622 (N_33622,N_29465,N_29891);
or U33623 (N_33623,N_29146,N_22914);
nor U33624 (N_33624,N_23027,N_24252);
or U33625 (N_33625,N_28310,N_21224);
nand U33626 (N_33626,N_20119,N_26480);
nand U33627 (N_33627,N_24157,N_22254);
nand U33628 (N_33628,N_26521,N_29195);
and U33629 (N_33629,N_28822,N_29159);
or U33630 (N_33630,N_24375,N_29558);
nor U33631 (N_33631,N_22012,N_28962);
or U33632 (N_33632,N_26497,N_22127);
or U33633 (N_33633,N_28956,N_21734);
and U33634 (N_33634,N_27789,N_29126);
and U33635 (N_33635,N_27282,N_20346);
and U33636 (N_33636,N_25887,N_20206);
nand U33637 (N_33637,N_24858,N_21831);
or U33638 (N_33638,N_20087,N_28452);
nand U33639 (N_33639,N_24716,N_24911);
xor U33640 (N_33640,N_28149,N_21612);
and U33641 (N_33641,N_24487,N_22836);
or U33642 (N_33642,N_23763,N_22058);
and U33643 (N_33643,N_26360,N_20929);
and U33644 (N_33644,N_26968,N_26987);
and U33645 (N_33645,N_22215,N_29547);
and U33646 (N_33646,N_28235,N_24447);
or U33647 (N_33647,N_20542,N_28347);
nor U33648 (N_33648,N_26427,N_25771);
nor U33649 (N_33649,N_26268,N_25811);
and U33650 (N_33650,N_25341,N_29221);
and U33651 (N_33651,N_27293,N_21088);
and U33652 (N_33652,N_29027,N_26418);
xnor U33653 (N_33653,N_26119,N_22905);
and U33654 (N_33654,N_21350,N_28444);
and U33655 (N_33655,N_24382,N_22437);
or U33656 (N_33656,N_24755,N_22153);
and U33657 (N_33657,N_20191,N_21840);
and U33658 (N_33658,N_29925,N_20463);
or U33659 (N_33659,N_20210,N_20826);
nor U33660 (N_33660,N_25193,N_25164);
and U33661 (N_33661,N_22178,N_22105);
or U33662 (N_33662,N_21741,N_23142);
or U33663 (N_33663,N_29548,N_26944);
or U33664 (N_33664,N_21268,N_25035);
xnor U33665 (N_33665,N_22060,N_24929);
nand U33666 (N_33666,N_20530,N_21754);
and U33667 (N_33667,N_29532,N_27055);
nand U33668 (N_33668,N_27440,N_25135);
nor U33669 (N_33669,N_23970,N_21705);
or U33670 (N_33670,N_27768,N_23495);
or U33671 (N_33671,N_26900,N_20762);
and U33672 (N_33672,N_22159,N_23853);
or U33673 (N_33673,N_25189,N_27465);
or U33674 (N_33674,N_24395,N_26454);
xor U33675 (N_33675,N_26719,N_25846);
or U33676 (N_33676,N_22839,N_22537);
or U33677 (N_33677,N_25009,N_24565);
nand U33678 (N_33678,N_24902,N_26534);
and U33679 (N_33679,N_26213,N_24989);
nor U33680 (N_33680,N_27298,N_27205);
xnor U33681 (N_33681,N_25627,N_21363);
and U33682 (N_33682,N_25879,N_20012);
and U33683 (N_33683,N_20498,N_28029);
or U33684 (N_33684,N_27602,N_26224);
or U33685 (N_33685,N_24556,N_21394);
xnor U33686 (N_33686,N_21814,N_21683);
xnor U33687 (N_33687,N_25934,N_29359);
xor U33688 (N_33688,N_25954,N_20536);
nor U33689 (N_33689,N_22335,N_25891);
nor U33690 (N_33690,N_28248,N_22160);
xnor U33691 (N_33691,N_22637,N_27325);
xnor U33692 (N_33692,N_27794,N_28809);
nand U33693 (N_33693,N_22701,N_23573);
xor U33694 (N_33694,N_25538,N_26318);
and U33695 (N_33695,N_27319,N_21327);
nand U33696 (N_33696,N_28895,N_21605);
xor U33697 (N_33697,N_20113,N_21960);
nand U33698 (N_33698,N_25310,N_23852);
xor U33699 (N_33699,N_23899,N_23190);
xor U33700 (N_33700,N_22384,N_24463);
and U33701 (N_33701,N_29643,N_25542);
nand U33702 (N_33702,N_28665,N_20418);
nor U33703 (N_33703,N_21639,N_20345);
and U33704 (N_33704,N_21106,N_23146);
nand U33705 (N_33705,N_20557,N_22353);
and U33706 (N_33706,N_20307,N_29594);
nor U33707 (N_33707,N_20637,N_27154);
or U33708 (N_33708,N_21781,N_23023);
nand U33709 (N_33709,N_21045,N_21709);
and U33710 (N_33710,N_29691,N_21786);
xor U33711 (N_33711,N_28986,N_27990);
or U33712 (N_33712,N_29597,N_24041);
nor U33713 (N_33713,N_24368,N_22381);
or U33714 (N_33714,N_24173,N_21447);
nor U33715 (N_33715,N_27270,N_25544);
or U33716 (N_33716,N_29674,N_29958);
and U33717 (N_33717,N_27417,N_27659);
or U33718 (N_33718,N_20267,N_25928);
nor U33719 (N_33719,N_23000,N_21200);
nand U33720 (N_33720,N_23758,N_21993);
nor U33721 (N_33721,N_25567,N_21374);
nor U33722 (N_33722,N_20630,N_27487);
or U33723 (N_33723,N_28423,N_28764);
nor U33724 (N_33724,N_23486,N_22911);
or U33725 (N_33725,N_23370,N_20517);
and U33726 (N_33726,N_24708,N_27548);
or U33727 (N_33727,N_20001,N_29660);
and U33728 (N_33728,N_24848,N_24637);
and U33729 (N_33729,N_28582,N_26908);
or U33730 (N_33730,N_22519,N_29260);
nand U33731 (N_33731,N_21710,N_23019);
and U33732 (N_33732,N_21634,N_23013);
nand U33733 (N_33733,N_22913,N_23517);
xnor U33734 (N_33734,N_20286,N_25944);
and U33735 (N_33735,N_27777,N_26576);
or U33736 (N_33736,N_20185,N_22774);
nor U33737 (N_33737,N_25290,N_25697);
nand U33738 (N_33738,N_22995,N_22310);
or U33739 (N_33739,N_23541,N_22763);
or U33740 (N_33740,N_27024,N_28553);
nand U33741 (N_33741,N_22743,N_23077);
xnor U33742 (N_33742,N_25160,N_25941);
nand U33743 (N_33743,N_27285,N_25180);
nor U33744 (N_33744,N_24307,N_28518);
or U33745 (N_33745,N_24248,N_29509);
nor U33746 (N_33746,N_22395,N_29316);
and U33747 (N_33747,N_23187,N_20852);
nand U33748 (N_33748,N_26288,N_27535);
nor U33749 (N_33749,N_28844,N_29748);
nor U33750 (N_33750,N_24555,N_24376);
nor U33751 (N_33751,N_24782,N_27333);
nand U33752 (N_33752,N_27343,N_22552);
and U33753 (N_33753,N_23768,N_29151);
or U33754 (N_33754,N_25454,N_22236);
nor U33755 (N_33755,N_23646,N_29440);
nor U33756 (N_33756,N_21359,N_23151);
xor U33757 (N_33757,N_27005,N_27012);
or U33758 (N_33758,N_25258,N_23948);
or U33759 (N_33759,N_29657,N_21532);
nand U33760 (N_33760,N_25457,N_24545);
or U33761 (N_33761,N_22589,N_25393);
xnor U33762 (N_33762,N_25646,N_25528);
or U33763 (N_33763,N_20893,N_20122);
and U33764 (N_33764,N_21513,N_24208);
and U33765 (N_33765,N_27244,N_29103);
nand U33766 (N_33766,N_28228,N_24477);
and U33767 (N_33767,N_26191,N_22531);
or U33768 (N_33768,N_27827,N_26054);
nand U33769 (N_33769,N_29623,N_27559);
and U33770 (N_33770,N_26717,N_25336);
and U33771 (N_33771,N_21311,N_21821);
xnor U33772 (N_33772,N_23253,N_22441);
nand U33773 (N_33773,N_29648,N_27677);
or U33774 (N_33774,N_24108,N_28398);
xnor U33775 (N_33775,N_28306,N_29478);
xnor U33776 (N_33776,N_27363,N_20569);
or U33777 (N_33777,N_29018,N_26693);
and U33778 (N_33778,N_21809,N_28496);
nor U33779 (N_33779,N_28817,N_21900);
xor U33780 (N_33780,N_24266,N_22983);
xnor U33781 (N_33781,N_28789,N_24236);
or U33782 (N_33782,N_22370,N_28121);
nand U33783 (N_33783,N_20075,N_29496);
nand U33784 (N_33784,N_22848,N_20271);
xnor U33785 (N_33785,N_25704,N_28006);
xor U33786 (N_33786,N_24969,N_28357);
nand U33787 (N_33787,N_23263,N_28985);
xnor U33788 (N_33788,N_27616,N_25218);
and U33789 (N_33789,N_28792,N_20385);
or U33790 (N_33790,N_22343,N_22041);
or U33791 (N_33791,N_23422,N_21320);
and U33792 (N_33792,N_24722,N_20761);
and U33793 (N_33793,N_25014,N_27937);
nand U33794 (N_33794,N_27744,N_24517);
and U33795 (N_33795,N_25266,N_28682);
or U33796 (N_33796,N_26137,N_28209);
nor U33797 (N_33797,N_26608,N_23282);
nand U33798 (N_33798,N_24222,N_26041);
or U33799 (N_33799,N_27291,N_24731);
or U33800 (N_33800,N_28189,N_21731);
nor U33801 (N_33801,N_21953,N_26018);
and U33802 (N_33802,N_27663,N_21907);
nand U33803 (N_33803,N_27611,N_21694);
nor U33804 (N_33804,N_24340,N_22390);
or U33805 (N_33805,N_24488,N_26561);
nand U33806 (N_33806,N_24992,N_27202);
nand U33807 (N_33807,N_23017,N_22465);
nand U33808 (N_33808,N_28249,N_27957);
nand U33809 (N_33809,N_25893,N_22773);
xnor U33810 (N_33810,N_26676,N_26784);
or U33811 (N_33811,N_22959,N_24352);
nor U33812 (N_33812,N_24897,N_29307);
xnor U33813 (N_33813,N_21468,N_21285);
and U33814 (N_33814,N_25536,N_28708);
or U33815 (N_33815,N_23587,N_20796);
nor U33816 (N_33816,N_23793,N_24524);
or U33817 (N_33817,N_28412,N_22856);
nand U33818 (N_33818,N_23604,N_26986);
or U33819 (N_33819,N_24648,N_24912);
nor U33820 (N_33820,N_28724,N_27158);
xor U33821 (N_33821,N_21600,N_26721);
nor U33822 (N_33822,N_22298,N_28968);
xnor U33823 (N_33823,N_26626,N_22783);
or U33824 (N_33824,N_26389,N_23237);
nor U33825 (N_33825,N_25601,N_29336);
nor U33826 (N_33826,N_26263,N_21982);
and U33827 (N_33827,N_20139,N_28565);
or U33828 (N_33828,N_28188,N_20554);
xnor U33829 (N_33829,N_26247,N_26299);
or U33830 (N_33830,N_27818,N_29562);
nand U33831 (N_33831,N_24815,N_22824);
xnor U33832 (N_33832,N_24832,N_22919);
nand U33833 (N_33833,N_28415,N_21740);
or U33834 (N_33834,N_25067,N_26124);
nor U33835 (N_33835,N_21717,N_25297);
nor U33836 (N_33836,N_24424,N_22600);
nand U33837 (N_33837,N_27348,N_20265);
nand U33838 (N_33838,N_26046,N_24014);
xor U33839 (N_33839,N_26201,N_24010);
nand U33840 (N_33840,N_27046,N_29522);
xor U33841 (N_33841,N_21206,N_23744);
and U33842 (N_33842,N_21930,N_26588);
nand U33843 (N_33843,N_28070,N_28959);
and U33844 (N_33844,N_22812,N_23239);
nor U33845 (N_33845,N_22458,N_26182);
xnor U33846 (N_33846,N_26919,N_24472);
xor U33847 (N_33847,N_21054,N_26279);
xor U33848 (N_33848,N_25596,N_23202);
xor U33849 (N_33849,N_27822,N_29173);
nand U33850 (N_33850,N_26238,N_24379);
xor U33851 (N_33851,N_22918,N_26405);
and U33852 (N_33852,N_29409,N_26864);
nor U33853 (N_33853,N_21160,N_27784);
nand U33854 (N_33854,N_20268,N_20653);
nand U33855 (N_33855,N_23144,N_23592);
nor U33856 (N_33856,N_24186,N_29658);
nor U33857 (N_33857,N_24356,N_23519);
nor U33858 (N_33858,N_22583,N_21711);
nand U33859 (N_33859,N_21253,N_27776);
or U33860 (N_33860,N_24417,N_24317);
nand U33861 (N_33861,N_29534,N_26824);
or U33862 (N_33862,N_25367,N_21072);
nor U33863 (N_33863,N_26651,N_20093);
or U33864 (N_33864,N_20976,N_29979);
nor U33865 (N_33865,N_23341,N_24444);
xnor U33866 (N_33866,N_24469,N_29223);
and U33867 (N_33867,N_26880,N_22414);
nand U33868 (N_33868,N_21043,N_25439);
xor U33869 (N_33869,N_21498,N_26486);
xor U33870 (N_33870,N_27918,N_29252);
nand U33871 (N_33871,N_21901,N_28909);
xor U33872 (N_33872,N_24302,N_25378);
nor U33873 (N_33873,N_26749,N_23841);
nor U33874 (N_33874,N_26262,N_24033);
or U33875 (N_33875,N_27267,N_21491);
and U33876 (N_33876,N_27111,N_29589);
nor U33877 (N_33877,N_21815,N_28548);
nor U33878 (N_33878,N_25799,N_28753);
xnor U33879 (N_33879,N_27224,N_24299);
or U33880 (N_33880,N_27670,N_23518);
or U33881 (N_33881,N_21179,N_24446);
and U33882 (N_33882,N_22036,N_25784);
nor U33883 (N_33883,N_25932,N_22808);
nor U33884 (N_33884,N_29098,N_20023);
and U33885 (N_33885,N_28229,N_27866);
and U33886 (N_33886,N_25531,N_28055);
and U33887 (N_33887,N_24128,N_21483);
xnor U33888 (N_33888,N_23730,N_23369);
nand U33889 (N_33889,N_26610,N_28905);
and U33890 (N_33890,N_21229,N_25311);
xor U33891 (N_33891,N_22545,N_21343);
and U33892 (N_33892,N_25622,N_24645);
nand U33893 (N_33893,N_23454,N_29463);
and U33894 (N_33894,N_28619,N_21188);
or U33895 (N_33895,N_24002,N_23583);
nor U33896 (N_33896,N_23738,N_22944);
nor U33897 (N_33897,N_27614,N_20213);
nor U33898 (N_33898,N_23171,N_27088);
xnor U33899 (N_33899,N_24066,N_24706);
xor U33900 (N_33900,N_29233,N_23391);
and U33901 (N_33901,N_22438,N_27095);
nor U33902 (N_33902,N_25195,N_26323);
xor U33903 (N_33903,N_24689,N_24612);
xor U33904 (N_33904,N_22137,N_22430);
xor U33905 (N_33905,N_23662,N_25741);
nand U33906 (N_33906,N_28002,N_26961);
xor U33907 (N_33907,N_21213,N_25906);
and U33908 (N_33908,N_23015,N_25141);
xor U33909 (N_33909,N_21473,N_23393);
and U33910 (N_33910,N_28938,N_21150);
nand U33911 (N_33911,N_23320,N_28650);
xor U33912 (N_33912,N_20675,N_26452);
xor U33913 (N_33913,N_28242,N_22749);
nand U33914 (N_33914,N_22964,N_20933);
nor U33915 (N_33915,N_24536,N_22014);
xnor U33916 (N_33916,N_24402,N_20019);
nor U33917 (N_33917,N_21240,N_25410);
or U33918 (N_33918,N_21386,N_21788);
or U33919 (N_33919,N_23624,N_25574);
nand U33920 (N_33920,N_29587,N_24037);
or U33921 (N_33921,N_21225,N_29324);
nor U33922 (N_33922,N_29498,N_20384);
or U33923 (N_33923,N_27003,N_21837);
nor U33924 (N_33924,N_29461,N_26783);
or U33925 (N_33925,N_28867,N_23278);
xor U33926 (N_33926,N_29810,N_26580);
or U33927 (N_33927,N_28907,N_23946);
nand U33928 (N_33928,N_23739,N_27130);
nand U33929 (N_33929,N_27510,N_28258);
nor U33930 (N_33930,N_24197,N_22068);
or U33931 (N_33931,N_20723,N_20836);
and U33932 (N_33932,N_26584,N_21030);
nand U33933 (N_33933,N_24812,N_21100);
or U33934 (N_33934,N_27382,N_29741);
nor U33935 (N_33935,N_25656,N_28728);
nor U33936 (N_33936,N_25062,N_25852);
nor U33937 (N_33937,N_25561,N_23265);
and U33938 (N_33938,N_20056,N_26415);
nand U33939 (N_33939,N_24267,N_24862);
nor U33940 (N_33940,N_23046,N_21666);
nand U33941 (N_33941,N_21015,N_25971);
xor U33942 (N_33942,N_29265,N_23199);
xnor U33943 (N_33943,N_20303,N_29015);
and U33944 (N_33944,N_28566,N_21779);
nor U33945 (N_33945,N_23682,N_28404);
nand U33946 (N_33946,N_25492,N_25560);
and U33947 (N_33947,N_28196,N_24561);
or U33948 (N_33948,N_28204,N_21194);
nand U33949 (N_33949,N_26080,N_28425);
and U33950 (N_33950,N_25460,N_25282);
and U33951 (N_33951,N_27921,N_25927);
and U33952 (N_33952,N_25786,N_24527);
or U33953 (N_33953,N_21292,N_20904);
or U33954 (N_33954,N_24050,N_23526);
nor U33955 (N_33955,N_21664,N_22415);
xnor U33956 (N_33956,N_24217,N_25720);
nor U33957 (N_33957,N_28888,N_24587);
or U33958 (N_33958,N_27446,N_25211);
nand U33959 (N_33959,N_29793,N_28678);
and U33960 (N_33960,N_21445,N_28177);
nor U33961 (N_33961,N_20932,N_23581);
xnor U33962 (N_33962,N_20773,N_28019);
xor U33963 (N_33963,N_26945,N_29097);
xnor U33964 (N_33964,N_27384,N_23503);
or U33965 (N_33965,N_24580,N_29563);
nor U33966 (N_33966,N_21131,N_23161);
or U33967 (N_33967,N_20858,N_26653);
nand U33968 (N_33968,N_29770,N_20926);
nor U33969 (N_33969,N_25420,N_22625);
nand U33970 (N_33970,N_20076,N_26406);
nor U33971 (N_33971,N_25989,N_20752);
nor U33972 (N_33972,N_24939,N_28658);
and U33973 (N_33973,N_23621,N_25637);
xnor U33974 (N_33974,N_21789,N_22250);
nand U33975 (N_33975,N_20283,N_26950);
xor U33976 (N_33976,N_21031,N_22404);
or U33977 (N_33977,N_22309,N_22585);
nand U33978 (N_33978,N_28074,N_22678);
and U33979 (N_33979,N_28814,N_24603);
nand U33980 (N_33980,N_28205,N_20970);
or U33981 (N_33981,N_28088,N_23851);
nor U33982 (N_33982,N_28372,N_25869);
nor U33983 (N_33983,N_24169,N_22352);
or U33984 (N_33984,N_20800,N_25407);
and U33985 (N_33985,N_28592,N_22575);
xor U33986 (N_33986,N_22960,N_25423);
or U33987 (N_33987,N_22650,N_26777);
xnor U33988 (N_33988,N_26312,N_22644);
nand U33989 (N_33989,N_21332,N_25674);
and U33990 (N_33990,N_26349,N_28603);
nand U33991 (N_33991,N_22490,N_25153);
nor U33992 (N_33992,N_29957,N_20632);
and U33993 (N_33993,N_24614,N_28725);
xor U33994 (N_33994,N_24663,N_23043);
nand U33995 (N_33995,N_20254,N_28143);
and U33996 (N_33996,N_20614,N_26575);
nor U33997 (N_33997,N_20604,N_28443);
nand U33998 (N_33998,N_26164,N_22862);
nor U33999 (N_33999,N_21637,N_27341);
and U34000 (N_34000,N_23811,N_27609);
and U34001 (N_34001,N_21163,N_21433);
nand U34002 (N_34002,N_24798,N_26566);
nand U34003 (N_34003,N_29052,N_26645);
nand U34004 (N_34004,N_28979,N_27610);
and U34005 (N_34005,N_26507,N_24433);
or U34006 (N_34006,N_25206,N_24196);
and U34007 (N_34007,N_20625,N_26538);
nand U34008 (N_34008,N_28406,N_21868);
or U34009 (N_34009,N_25506,N_21406);
nand U34010 (N_34010,N_24752,N_23122);
nand U34011 (N_34011,N_21570,N_28023);
nand U34012 (N_34012,N_25519,N_23647);
nor U34013 (N_34013,N_28407,N_28629);
or U34014 (N_34014,N_25059,N_29468);
xnor U34015 (N_34015,N_20786,N_26722);
or U34016 (N_34016,N_25363,N_26882);
or U34017 (N_34017,N_21451,N_24576);
and U34018 (N_34018,N_29624,N_23149);
and U34019 (N_34019,N_25208,N_20512);
or U34020 (N_34020,N_21556,N_28602);
xnor U34021 (N_34021,N_24476,N_27862);
or U34022 (N_34022,N_29681,N_21522);
nand U34023 (N_34023,N_21368,N_22252);
or U34024 (N_34024,N_29620,N_22935);
or U34025 (N_34025,N_24106,N_25278);
nor U34026 (N_34026,N_22734,N_26278);
and U34027 (N_34027,N_22368,N_20855);
and U34028 (N_34028,N_27835,N_27294);
and U34029 (N_34029,N_28980,N_26431);
nor U34030 (N_34030,N_27570,N_23687);
nor U34031 (N_34031,N_23676,N_28304);
nand U34032 (N_34032,N_22110,N_21340);
or U34033 (N_34033,N_28693,N_21403);
and U34034 (N_34034,N_23195,N_29724);
and U34035 (N_34035,N_22997,N_29284);
and U34036 (N_34036,N_26107,N_23467);
nand U34037 (N_34037,N_23180,N_24031);
or U34038 (N_34038,N_21715,N_25732);
xor U34039 (N_34039,N_29456,N_27711);
xor U34040 (N_34040,N_26065,N_26236);
or U34041 (N_34041,N_22527,N_26306);
xor U34042 (N_34042,N_22051,N_24875);
xnor U34043 (N_34043,N_29605,N_28371);
nor U34044 (N_34044,N_25444,N_23333);
nor U34045 (N_34045,N_20865,N_22141);
nand U34046 (N_34046,N_23634,N_25231);
or U34047 (N_34047,N_23339,N_24611);
nor U34048 (N_34048,N_28990,N_29168);
nand U34049 (N_34049,N_28215,N_24179);
nor U34050 (N_34050,N_24323,N_27956);
xor U34051 (N_34051,N_21947,N_26694);
nand U34052 (N_34052,N_29560,N_27841);
xnor U34053 (N_34053,N_27542,N_21759);
nor U34054 (N_34054,N_20294,N_25867);
and U34055 (N_34055,N_28775,N_24419);
nand U34056 (N_34056,N_25830,N_28384);
and U34057 (N_34057,N_27857,N_22732);
xnor U34058 (N_34058,N_20124,N_25268);
nand U34059 (N_34059,N_29011,N_22683);
nor U34060 (N_34060,N_27230,N_23562);
nand U34061 (N_34061,N_24054,N_26112);
and U34062 (N_34062,N_20474,N_28254);
nor U34063 (N_34063,N_29432,N_28277);
xnor U34064 (N_34064,N_21370,N_22768);
or U34065 (N_34065,N_27817,N_28231);
nor U34066 (N_34066,N_28626,N_24288);
or U34067 (N_34067,N_20960,N_23480);
or U34068 (N_34068,N_25838,N_25426);
and U34069 (N_34069,N_23219,N_22898);
nor U34070 (N_34070,N_29596,N_21818);
or U34071 (N_34071,N_20156,N_26873);
or U34072 (N_34072,N_29510,N_25607);
nand U34073 (N_34073,N_28746,N_21324);
or U34074 (N_34074,N_23896,N_24311);
or U34075 (N_34075,N_21890,N_22258);
nand U34076 (N_34076,N_27725,N_21295);
xnor U34077 (N_34077,N_25594,N_20522);
or U34078 (N_34078,N_27075,N_29894);
nor U34079 (N_34079,N_26984,N_29486);
xor U34080 (N_34080,N_25092,N_25504);
nor U34081 (N_34081,N_23593,N_22901);
or U34082 (N_34082,N_23606,N_27441);
nor U34083 (N_34083,N_21512,N_26603);
xnor U34084 (N_34084,N_29325,N_28737);
and U34085 (N_34085,N_25623,N_20679);
xor U34086 (N_34086,N_20958,N_26425);
and U34087 (N_34087,N_22446,N_25721);
or U34088 (N_34088,N_20863,N_29703);
or U34089 (N_34089,N_28966,N_20987);
and U34090 (N_34090,N_26383,N_22977);
and U34091 (N_34091,N_29870,N_21592);
nor U34092 (N_34092,N_27543,N_28256);
nand U34093 (N_34093,N_29323,N_26376);
xnor U34094 (N_34094,N_24192,N_24008);
nor U34095 (N_34095,N_29220,N_21305);
xor U34096 (N_34096,N_20727,N_27206);
and U34097 (N_34097,N_23535,N_20234);
or U34098 (N_34098,N_26641,N_23003);
xnor U34099 (N_34099,N_29267,N_29169);
or U34100 (N_34100,N_26353,N_22779);
and U34101 (N_34101,N_27404,N_29622);
xnor U34102 (N_34102,N_25742,N_23838);
and U34103 (N_34103,N_26782,N_27001);
or U34104 (N_34104,N_21908,N_23323);
nor U34105 (N_34105,N_23812,N_28640);
and U34106 (N_34106,N_22273,N_28879);
and U34107 (N_34107,N_26037,N_28823);
xnor U34108 (N_34108,N_27979,N_21511);
nand U34109 (N_34109,N_24071,N_21658);
nand U34110 (N_34110,N_26955,N_29129);
or U34111 (N_34111,N_27143,N_27011);
xnor U34112 (N_34112,N_25116,N_29666);
xnor U34113 (N_34113,N_21937,N_20395);
nor U34114 (N_34114,N_20775,N_29963);
and U34115 (N_34115,N_29859,N_29472);
nand U34116 (N_34116,N_28781,N_25845);
or U34117 (N_34117,N_26974,N_24970);
nand U34118 (N_34118,N_27856,N_23423);
nor U34119 (N_34119,N_28158,N_24141);
or U34120 (N_34120,N_23089,N_24808);
xnor U34121 (N_34121,N_23875,N_22013);
xor U34122 (N_34122,N_28477,N_26483);
nor U34123 (N_34123,N_26910,N_24617);
or U34124 (N_34124,N_23860,N_20756);
nand U34125 (N_34125,N_26006,N_20017);
and U34126 (N_34126,N_26166,N_29999);
xnor U34127 (N_34127,N_23932,N_21079);
xor U34128 (N_34128,N_24383,N_20746);
nor U34129 (N_34129,N_28489,N_24364);
nand U34130 (N_34130,N_23257,N_20212);
and U34131 (N_34131,N_23885,N_27770);
nand U34132 (N_34132,N_20380,N_20194);
and U34133 (N_34133,N_27351,N_25209);
and U34134 (N_34134,N_28292,N_22511);
or U34135 (N_34135,N_27869,N_25093);
or U34136 (N_34136,N_25921,N_22429);
nand U34137 (N_34137,N_22031,N_29890);
nor U34138 (N_34138,N_26019,N_28813);
nor U34139 (N_34139,N_25643,N_24072);
and U34140 (N_34140,N_21216,N_24018);
nor U34141 (N_34141,N_24996,N_20462);
or U34142 (N_34142,N_21819,N_25657);
nor U34143 (N_34143,N_25701,N_27229);
nand U34144 (N_34144,N_20523,N_26981);
nand U34145 (N_34145,N_25552,N_23468);
nand U34146 (N_34146,N_21020,N_20578);
nand U34147 (N_34147,N_25148,N_23878);
or U34148 (N_34148,N_24422,N_24640);
nand U34149 (N_34149,N_24773,N_27324);
and U34150 (N_34150,N_21048,N_22705);
or U34151 (N_34151,N_29812,N_26043);
nand U34152 (N_34152,N_27914,N_23053);
xor U34153 (N_34153,N_26165,N_26932);
and U34154 (N_34154,N_28998,N_25668);
nor U34155 (N_34155,N_24115,N_22979);
or U34156 (N_34156,N_28856,N_21004);
nor U34157 (N_34157,N_23109,N_23157);
nand U34158 (N_34158,N_28245,N_23864);
nor U34159 (N_34159,N_28374,N_23001);
or U34160 (N_34160,N_29990,N_25040);
nor U34161 (N_34161,N_23975,N_24820);
or U34162 (N_34162,N_28880,N_20311);
and U34163 (N_34163,N_28414,N_29991);
nor U34164 (N_34164,N_23158,N_27181);
xnor U34165 (N_34165,N_24959,N_27096);
nor U34166 (N_34166,N_27521,N_20638);
xnor U34167 (N_34167,N_22982,N_27642);
nand U34168 (N_34168,N_22741,N_20782);
or U34169 (N_34169,N_21922,N_28352);
nor U34170 (N_34170,N_27538,N_24310);
xor U34171 (N_34171,N_28672,N_29791);
xor U34172 (N_34172,N_22257,N_29880);
or U34173 (N_34173,N_24943,N_24735);
nand U34174 (N_34174,N_24936,N_22927);
nor U34175 (N_34175,N_25104,N_27897);
or U34176 (N_34176,N_21591,N_25450);
xnor U34177 (N_34177,N_23429,N_22605);
nor U34178 (N_34178,N_24876,N_24501);
nor U34179 (N_34179,N_29641,N_22188);
nand U34180 (N_34180,N_20353,N_23512);
nand U34181 (N_34181,N_23807,N_22572);
and U34182 (N_34182,N_24763,N_29091);
nand U34183 (N_34183,N_28270,N_26260);
xnor U34184 (N_34184,N_25820,N_27276);
and U34185 (N_34185,N_28591,N_28311);
xor U34186 (N_34186,N_20379,N_20159);
and U34187 (N_34187,N_23767,N_25075);
or U34188 (N_34188,N_23580,N_29920);
nor U34189 (N_34189,N_29926,N_23955);
or U34190 (N_34190,N_20374,N_25397);
and U34191 (N_34191,N_26217,N_25653);
and U34192 (N_34192,N_23016,N_26681);
and U34193 (N_34193,N_22940,N_24776);
and U34194 (N_34194,N_21980,N_21023);
or U34195 (N_34195,N_20541,N_20584);
xor U34196 (N_34196,N_24805,N_28368);
nor U34197 (N_34197,N_20042,N_24079);
and U34198 (N_34198,N_28991,N_29377);
xor U34199 (N_34199,N_20046,N_26619);
or U34200 (N_34200,N_20837,N_26409);
xor U34201 (N_34201,N_20320,N_23470);
nand U34202 (N_34202,N_26788,N_22413);
xor U34203 (N_34203,N_23743,N_24928);
or U34204 (N_34204,N_22608,N_25203);
nand U34205 (N_34205,N_20915,N_25526);
or U34206 (N_34206,N_28307,N_26650);
nand U34207 (N_34207,N_24693,N_24844);
and U34208 (N_34208,N_26059,N_28502);
and U34209 (N_34209,N_20079,N_24796);
xnor U34210 (N_34210,N_24085,N_28457);
or U34211 (N_34211,N_22354,N_24211);
and U34212 (N_34212,N_25288,N_24328);
and U34213 (N_34213,N_23280,N_25553);
or U34214 (N_34214,N_21335,N_28265);
nor U34215 (N_34215,N_24816,N_25694);
xor U34216 (N_34216,N_27717,N_23530);
or U34217 (N_34217,N_20682,N_29476);
nand U34218 (N_34218,N_24144,N_21410);
and U34219 (N_34219,N_28594,N_29123);
or U34220 (N_34220,N_21912,N_25025);
nand U34221 (N_34221,N_22713,N_25540);
and U34222 (N_34222,N_24199,N_22274);
xor U34223 (N_34223,N_21673,N_25002);
and U34224 (N_34224,N_22704,N_25370);
nor U34225 (N_34225,N_23078,N_25917);
nand U34226 (N_34226,N_22943,N_24127);
xnor U34227 (N_34227,N_28253,N_27337);
or U34228 (N_34228,N_24110,N_27086);
nand U34229 (N_34229,N_23008,N_27275);
nand U34230 (N_34230,N_29806,N_29028);
nand U34231 (N_34231,N_24427,N_26796);
nand U34232 (N_34232,N_22026,N_20551);
nand U34233 (N_34233,N_26800,N_26959);
and U34234 (N_34234,N_26902,N_29155);
xnor U34235 (N_34235,N_23496,N_25687);
or U34236 (N_34236,N_25874,N_29434);
xnor U34237 (N_34237,N_24988,N_21052);
nand U34238 (N_34238,N_25130,N_23849);
or U34239 (N_34239,N_25312,N_23803);
nor U34240 (N_34240,N_28785,N_23132);
or U34241 (N_34241,N_21068,N_22912);
xor U34242 (N_34242,N_24405,N_24599);
or U34243 (N_34243,N_25057,N_27412);
xor U34244 (N_34244,N_22104,N_21455);
nor U34245 (N_34245,N_25292,N_25518);
and U34246 (N_34246,N_21918,N_21402);
nor U34247 (N_34247,N_24438,N_28035);
or U34248 (N_34248,N_21083,N_29390);
xor U34249 (N_34249,N_26627,N_23990);
xnor U34250 (N_34250,N_24591,N_28045);
nand U34251 (N_34251,N_24849,N_23311);
or U34252 (N_34252,N_20846,N_27418);
and U34253 (N_34253,N_24178,N_24453);
and U34254 (N_34254,N_26509,N_24123);
xor U34255 (N_34255,N_20945,N_21114);
nor U34256 (N_34256,N_24788,N_29415);
xor U34257 (N_34257,N_29989,N_22029);
nand U34258 (N_34258,N_21442,N_27756);
or U34259 (N_34259,N_29227,N_27167);
nand U34260 (N_34260,N_27771,N_23473);
xnor U34261 (N_34261,N_20145,N_29637);
and U34262 (N_34262,N_27917,N_20247);
nor U34263 (N_34263,N_29965,N_28395);
nor U34264 (N_34264,N_29049,N_26809);
xnor U34265 (N_34265,N_28369,N_20951);
nor U34266 (N_34266,N_21330,N_26239);
nand U34267 (N_34267,N_23136,N_25979);
nand U34268 (N_34268,N_22921,N_23609);
nand U34269 (N_34269,N_21493,N_29438);
nand U34270 (N_34270,N_29618,N_20869);
nand U34271 (N_34271,N_28439,N_29426);
nand U34272 (N_34272,N_25691,N_21118);
nand U34273 (N_34273,N_23072,N_21147);
xnor U34274 (N_34274,N_23307,N_29938);
or U34275 (N_34275,N_28448,N_23310);
nor U34276 (N_34276,N_22723,N_24149);
or U34277 (N_34277,N_27971,N_24120);
nand U34278 (N_34278,N_28180,N_21462);
nor U34279 (N_34279,N_23440,N_25026);
or U34280 (N_34280,N_26162,N_24857);
nor U34281 (N_34281,N_24814,N_28882);
and U34282 (N_34282,N_25619,N_23731);
nor U34283 (N_34283,N_26988,N_22318);
nor U34284 (N_34284,N_22132,N_26781);
and U34285 (N_34285,N_23942,N_26519);
nor U34286 (N_34286,N_27359,N_20843);
xnor U34287 (N_34287,N_24921,N_20891);
xnor U34288 (N_34288,N_26972,N_28691);
xnor U34289 (N_34289,N_29030,N_21236);
nor U34290 (N_34290,N_22691,N_26261);
or U34291 (N_34291,N_20358,N_23331);
nor U34292 (N_34292,N_23527,N_28690);
xor U34293 (N_34293,N_26799,N_24147);
nand U34294 (N_34294,N_27949,N_23718);
nor U34295 (N_34295,N_27273,N_23351);
xor U34296 (N_34296,N_24646,N_20942);
nand U34297 (N_34297,N_24150,N_29130);
and U34298 (N_34298,N_21376,N_27959);
nand U34299 (N_34299,N_29680,N_24028);
nor U34300 (N_34300,N_26136,N_20020);
nand U34301 (N_34301,N_24272,N_27842);
nor U34302 (N_34302,N_29907,N_26550);
xnor U34303 (N_34303,N_23105,N_23249);
and U34304 (N_34304,N_24827,N_27166);
xnor U34305 (N_34305,N_25907,N_23810);
nand U34306 (N_34306,N_27876,N_29187);
nand U34307 (N_34307,N_25692,N_25661);
nor U34308 (N_34308,N_25284,N_24726);
xnor U34309 (N_34309,N_24644,N_21168);
nand U34310 (N_34310,N_22183,N_21891);
nand U34311 (N_34311,N_28679,N_24162);
nor U34312 (N_34312,N_22525,N_26958);
and U34313 (N_34313,N_20193,N_25207);
nand U34314 (N_34314,N_20546,N_22790);
nand U34315 (N_34315,N_20302,N_21231);
and U34316 (N_34316,N_29760,N_25511);
and U34317 (N_34317,N_28441,N_26837);
xnor U34318 (N_34318,N_26504,N_28793);
and U34319 (N_34319,N_24175,N_21954);
xnor U34320 (N_34320,N_25967,N_27116);
nand U34321 (N_34321,N_28940,N_28530);
or U34322 (N_34322,N_24320,N_27632);
xnor U34323 (N_34323,N_20465,N_27438);
and U34324 (N_34324,N_24826,N_24557);
or U34325 (N_34325,N_26760,N_22091);
and U34326 (N_34326,N_25899,N_29878);
xnor U34327 (N_34327,N_28016,N_25066);
or U34328 (N_34328,N_26325,N_24540);
xnor U34329 (N_34329,N_23729,N_22248);
and U34330 (N_34330,N_23326,N_28326);
or U34331 (N_34331,N_23844,N_29245);
and U34332 (N_34332,N_22179,N_27564);
nand U34333 (N_34333,N_22209,N_22618);
xnor U34334 (N_34334,N_25739,N_24275);
and U34335 (N_34335,N_23705,N_26528);
and U34336 (N_34336,N_21095,N_23921);
nor U34337 (N_34337,N_23944,N_28767);
nand U34338 (N_34338,N_27682,N_20661);
and U34339 (N_34339,N_23086,N_25765);
nand U34340 (N_34340,N_25217,N_25792);
nor U34341 (N_34341,N_26967,N_29799);
or U34342 (N_34342,N_26031,N_20050);
xnor U34343 (N_34343,N_25621,N_27760);
nand U34344 (N_34344,N_27245,N_29581);
nand U34345 (N_34345,N_23846,N_23874);
nand U34346 (N_34346,N_21112,N_21184);
xnor U34347 (N_34347,N_23961,N_27991);
nand U34348 (N_34348,N_26510,N_23590);
nand U34349 (N_34349,N_23487,N_20597);
nand U34350 (N_34350,N_28899,N_24818);
xor U34351 (N_34351,N_25076,N_27987);
nand U34352 (N_34352,N_25773,N_22066);
nand U34353 (N_34353,N_25585,N_22196);
xor U34354 (N_34354,N_21409,N_20202);
xnor U34355 (N_34355,N_23174,N_29886);
xor U34356 (N_34356,N_22620,N_26092);
nand U34357 (N_34357,N_28999,N_20164);
nand U34358 (N_34358,N_24775,N_21884);
and U34359 (N_34359,N_29863,N_20582);
nand U34360 (N_34360,N_21076,N_22418);
and U34361 (N_34361,N_21959,N_27662);
nand U34362 (N_34362,N_24327,N_25616);
nand U34363 (N_34363,N_26204,N_26541);
and U34364 (N_34364,N_28358,N_22377);
nor U34365 (N_34365,N_21653,N_22007);
xor U34366 (N_34366,N_21103,N_24905);
xor U34367 (N_34367,N_25232,N_26029);
nor U34368 (N_34368,N_27152,N_22238);
xnor U34369 (N_34369,N_28134,N_27062);
and U34370 (N_34370,N_26540,N_21518);
or U34371 (N_34371,N_22364,N_28538);
xnor U34372 (N_34372,N_24387,N_22154);
nand U34373 (N_34373,N_24278,N_23300);
nor U34374 (N_34374,N_27890,N_23749);
nor U34375 (N_34375,N_23366,N_21443);
nor U34376 (N_34376,N_28252,N_27951);
xor U34377 (N_34377,N_24878,N_22939);
xnor U34378 (N_34378,N_29037,N_26410);
and U34379 (N_34379,N_20549,N_20258);
or U34380 (N_34380,N_23248,N_24562);
nor U34381 (N_34381,N_22145,N_27066);
xnor U34382 (N_34382,N_25912,N_20760);
or U34383 (N_34383,N_26613,N_20028);
xor U34384 (N_34384,N_23087,N_24279);
and U34385 (N_34385,N_29861,N_20154);
nand U34386 (N_34386,N_21981,N_22409);
xor U34387 (N_34387,N_25081,N_23889);
nand U34388 (N_34388,N_26928,N_20789);
nand U34389 (N_34389,N_26155,N_28119);
nand U34390 (N_34390,N_22989,N_24869);
nor U34391 (N_34391,N_25100,N_27600);
xor U34392 (N_34392,N_23117,N_22961);
and U34393 (N_34393,N_23989,N_25876);
xor U34394 (N_34394,N_24891,N_25136);
nor U34395 (N_34395,N_25545,N_22387);
and U34396 (N_34396,N_21566,N_24231);
nand U34397 (N_34397,N_25372,N_21339);
or U34398 (N_34398,N_20781,N_22284);
xnor U34399 (N_34399,N_21318,N_27666);
and U34400 (N_34400,N_28932,N_21602);
xnor U34401 (N_34401,N_24334,N_27312);
xor U34402 (N_34402,N_20696,N_23693);
nand U34403 (N_34403,N_23446,N_29571);
nor U34404 (N_34404,N_26177,N_27081);
xor U34405 (N_34405,N_20243,N_25680);
nand U34406 (N_34406,N_20591,N_27089);
nor U34407 (N_34407,N_21562,N_22861);
nand U34408 (N_34408,N_26898,N_23208);
or U34409 (N_34409,N_22016,N_20281);
or U34410 (N_34410,N_26487,N_24332);
and U34411 (N_34411,N_21620,N_26662);
nor U34412 (N_34412,N_20802,N_22393);
xnor U34413 (N_34413,N_29956,N_26026);
nand U34414 (N_34414,N_26258,N_26737);
or U34415 (N_34415,N_26096,N_22121);
xor U34416 (N_34416,N_28918,N_29009);
and U34417 (N_34417,N_20713,N_26429);
and U34418 (N_34418,N_20407,N_23420);
and U34419 (N_34419,N_22286,N_25102);
and U34420 (N_34420,N_22571,N_26816);
xor U34421 (N_34421,N_28500,N_23974);
nor U34422 (N_34422,N_29829,N_28721);
xnor U34423 (N_34423,N_20241,N_26408);
nand U34424 (N_34424,N_28532,N_24749);
nor U34425 (N_34425,N_21089,N_24881);
xnor U34426 (N_34426,N_27674,N_27031);
nand U34427 (N_34427,N_22401,N_28375);
nor U34428 (N_34428,N_22306,N_27225);
nand U34429 (N_34429,N_22607,N_22086);
xnor U34430 (N_34430,N_23426,N_28232);
nor U34431 (N_34431,N_23879,N_26110);
xnor U34432 (N_34432,N_28849,N_27413);
nand U34433 (N_34433,N_26079,N_25345);
or U34434 (N_34434,N_26437,N_24985);
nor U34435 (N_34435,N_24861,N_20594);
and U34436 (N_34436,N_23675,N_29466);
nor U34437 (N_34437,N_28939,N_27532);
and U34438 (N_34438,N_25673,N_25514);
xor U34439 (N_34439,N_24673,N_24264);
or U34440 (N_34440,N_29183,N_25570);
nand U34441 (N_34441,N_24151,N_29702);
and U34442 (N_34442,N_25885,N_26707);
nor U34443 (N_34443,N_25313,N_21606);
nand U34444 (N_34444,N_24522,N_27500);
nand U34445 (N_34445,N_23563,N_24011);
or U34446 (N_34446,N_23883,N_21909);
and U34447 (N_34447,N_21314,N_22684);
xor U34448 (N_34448,N_24748,N_20328);
nand U34449 (N_34449,N_20572,N_27685);
nor U34450 (N_34450,N_27539,N_24367);
nor U34451 (N_34451,N_22321,N_29134);
and U34452 (N_34452,N_27651,N_26040);
or U34453 (N_34453,N_24600,N_22611);
or U34454 (N_34454,N_27940,N_27047);
nand U34455 (N_34455,N_21282,N_25920);
xor U34456 (N_34456,N_25832,N_22275);
or U34457 (N_34457,N_20725,N_27615);
or U34458 (N_34458,N_28935,N_24088);
nor U34459 (N_34459,N_26264,N_26896);
nor U34460 (N_34460,N_25882,N_26206);
xnor U34461 (N_34461,N_20603,N_21568);
or U34462 (N_34462,N_21056,N_22800);
nand U34463 (N_34463,N_20814,N_21365);
or U34464 (N_34464,N_22721,N_25943);
or U34465 (N_34465,N_25261,N_23444);
or U34466 (N_34466,N_20308,N_28075);
or U34467 (N_34467,N_27772,N_21033);
nand U34468 (N_34468,N_24636,N_28217);
and U34469 (N_34469,N_25959,N_25796);
or U34470 (N_34470,N_26991,N_28572);
nor U34471 (N_34471,N_24271,N_27854);
nor U34472 (N_34472,N_28017,N_23342);
xor U34473 (N_34473,N_21377,N_22435);
xnor U34474 (N_34474,N_20989,N_27727);
nor U34475 (N_34475,N_23884,N_21929);
xnor U34476 (N_34476,N_29984,N_29815);
xnor U34477 (N_34477,N_26795,N_28535);
and U34478 (N_34478,N_25617,N_29545);
nand U34479 (N_34479,N_21342,N_29315);
and U34480 (N_34480,N_27385,N_23855);
nor U34481 (N_34481,N_28836,N_23623);
nor U34482 (N_34482,N_22670,N_23084);
xor U34483 (N_34483,N_25176,N_29043);
nor U34484 (N_34484,N_26677,N_21858);
and U34485 (N_34485,N_25812,N_21204);
or U34486 (N_34486,N_26812,N_29673);
xnor U34487 (N_34487,N_24177,N_23652);
xnor U34488 (N_34488,N_23101,N_29206);
xor U34489 (N_34489,N_29889,N_26733);
or U34490 (N_34490,N_22507,N_28166);
nor U34491 (N_34491,N_21671,N_24370);
and U34492 (N_34492,N_25507,N_28597);
xor U34493 (N_34493,N_23442,N_22357);
nand U34494 (N_34494,N_20768,N_23930);
or U34495 (N_34495,N_28144,N_26270);
or U34496 (N_34496,N_20390,N_20624);
xnor U34497 (N_34497,N_22291,N_26790);
xor U34498 (N_34498,N_25751,N_25630);
nand U34499 (N_34499,N_27458,N_23030);
nor U34500 (N_34500,N_27655,N_24595);
nand U34501 (N_34501,N_23937,N_21517);
and U34502 (N_34502,N_24589,N_24744);
nor U34503 (N_34503,N_23210,N_28555);
and U34504 (N_34504,N_24207,N_24392);
or U34505 (N_34505,N_27999,N_23834);
nand U34506 (N_34506,N_25356,N_29073);
or U34507 (N_34507,N_22579,N_21760);
nand U34508 (N_34508,N_20005,N_27879);
or U34509 (N_34509,N_28599,N_27203);
nand U34510 (N_34510,N_28950,N_28241);
and U34511 (N_34511,N_28635,N_28578);
nand U34512 (N_34512,N_24259,N_22350);
and U34513 (N_34513,N_21059,N_27624);
nand U34514 (N_34514,N_23965,N_21961);
or U34515 (N_34515,N_25909,N_25332);
xor U34516 (N_34516,N_20882,N_25678);
nor U34517 (N_34517,N_24742,N_29945);
or U34518 (N_34518,N_24734,N_22402);
or U34519 (N_34519,N_23891,N_22410);
nand U34520 (N_34520,N_21388,N_24774);
or U34521 (N_34521,N_25942,N_27639);
or U34522 (N_34522,N_21827,N_24435);
or U34523 (N_34523,N_24813,N_29285);
nor U34524 (N_34524,N_20280,N_26912);
nor U34525 (N_34525,N_26658,N_20801);
and U34526 (N_34526,N_21070,N_22716);
nor U34527 (N_34527,N_28446,N_27891);
nor U34528 (N_34528,N_20130,N_21323);
and U34529 (N_34529,N_23383,N_24799);
and U34530 (N_34530,N_24747,N_21371);
xor U34531 (N_34531,N_23565,N_26728);
and U34532 (N_34532,N_29872,N_23691);
xnor U34533 (N_34533,N_22456,N_27308);
xnor U34534 (N_34534,N_23868,N_26495);
nor U34535 (N_34535,N_27963,N_24237);
or U34536 (N_34536,N_28032,N_22023);
nor U34537 (N_34537,N_29431,N_27810);
and U34538 (N_34538,N_27720,N_21139);
and U34539 (N_34539,N_29401,N_20676);
or U34540 (N_34540,N_23137,N_28139);
nor U34541 (N_34541,N_28337,N_23222);
xnor U34542 (N_34542,N_24024,N_22477);
nor U34543 (N_34543,N_26624,N_22689);
xnor U34544 (N_34544,N_20478,N_21104);
or U34545 (N_34545,N_26334,N_23354);
xnor U34546 (N_34546,N_20409,N_28621);
and U34547 (N_34547,N_26469,N_26310);
nor U34548 (N_34548,N_28545,N_24956);
nand U34549 (N_34549,N_21415,N_20057);
xor U34550 (N_34550,N_22984,N_23181);
xnor U34551 (N_34551,N_26472,N_27317);
and U34552 (N_34552,N_24133,N_27415);
xnor U34553 (N_34553,N_29411,N_28445);
nor U34554 (N_34554,N_25640,N_29370);
or U34555 (N_34555,N_20600,N_27196);
and U34556 (N_34556,N_21624,N_27493);
and U34557 (N_34557,N_28647,N_23111);
xnor U34558 (N_34558,N_26178,N_26199);
or U34559 (N_34559,N_23707,N_20109);
xor U34560 (N_34560,N_24729,N_24675);
nand U34561 (N_34561,N_22649,N_24485);
or U34562 (N_34562,N_27373,N_26482);
or U34563 (N_34563,N_29916,N_27812);
and U34564 (N_34564,N_25031,N_21851);
nand U34565 (N_34565,N_22047,N_29067);
nand U34566 (N_34566,N_24064,N_27381);
nand U34567 (N_34567,N_26731,N_21580);
and U34568 (N_34568,N_25988,N_23153);
nor U34569 (N_34569,N_23129,N_28460);
nor U34570 (N_34570,N_20861,N_29322);
xnor U34571 (N_34571,N_20898,N_26130);
xor U34572 (N_34572,N_21465,N_24245);
and U34573 (N_34573,N_28863,N_26144);
nand U34574 (N_34574,N_26593,N_27790);
nand U34575 (N_34575,N_26152,N_24309);
and U34576 (N_34576,N_27123,N_27733);
and U34577 (N_34577,N_29774,N_26522);
or U34578 (N_34578,N_26831,N_23616);
nor U34579 (N_34579,N_25782,N_26319);
or U34580 (N_34580,N_26867,N_26284);
or U34581 (N_34581,N_21962,N_21265);
and U34582 (N_34582,N_25853,N_25050);
and U34583 (N_34583,N_21086,N_21218);
and U34584 (N_34584,N_23041,N_23984);
or U34585 (N_34585,N_26934,N_29969);
nand U34586 (N_34586,N_22653,N_25236);
nand U34587 (N_34587,N_21774,N_23192);
nor U34588 (N_34588,N_20422,N_29475);
and U34589 (N_34589,N_26990,N_21472);
xnor U34590 (N_34590,N_23197,N_28059);
and U34591 (N_34591,N_28408,N_26555);
xor U34592 (N_34592,N_24607,N_24949);
nand U34593 (N_34593,N_26071,N_26649);
nor U34594 (N_34594,N_21914,N_22568);
or U34595 (N_34595,N_21153,N_22444);
or U34596 (N_34596,N_29993,N_25803);
nor U34597 (N_34597,N_21540,N_24385);
nand U34598 (N_34598,N_24804,N_25248);
nand U34599 (N_34599,N_22103,N_28363);
or U34600 (N_34600,N_20452,N_23497);
nand U34601 (N_34601,N_27880,N_24635);
or U34602 (N_34602,N_26138,N_24412);
or U34603 (N_34603,N_26420,N_27882);
or U34604 (N_34604,N_28223,N_22900);
xnor U34605 (N_34605,N_24833,N_23626);
xnor U34606 (N_34606,N_26390,N_21811);
or U34607 (N_34607,N_27724,N_27208);
or U34608 (N_34608,N_21856,N_21886);
xor U34609 (N_34609,N_21887,N_22566);
or U34610 (N_34610,N_24688,N_28770);
nor U34611 (N_34611,N_21599,N_28610);
or U34612 (N_34612,N_27942,N_25780);
nor U34613 (N_34613,N_20475,N_24533);
and U34614 (N_34614,N_29915,N_20086);
nand U34615 (N_34615,N_20916,N_21707);
nand U34616 (N_34616,N_27739,N_26372);
and U34617 (N_34617,N_28266,N_27162);
or U34618 (N_34618,N_21251,N_24893);
xor U34619 (N_34619,N_24558,N_27331);
nand U34620 (N_34620,N_27863,N_25277);
nand U34621 (N_34621,N_26841,N_24457);
and U34622 (N_34622,N_26289,N_25950);
and U34623 (N_34623,N_28546,N_23776);
xor U34624 (N_34624,N_23881,N_22270);
or U34625 (N_34625,N_28847,N_27631);
nor U34626 (N_34626,N_26249,N_28681);
xnor U34627 (N_34627,N_26000,N_26846);
xnor U34628 (N_34628,N_21328,N_27131);
xor U34629 (N_34629,N_22769,N_25455);
nand U34630 (N_34630,N_24622,N_28361);
and U34631 (N_34631,N_25254,N_25417);
or U34632 (N_34632,N_22317,N_25384);
and U34633 (N_34633,N_24866,N_20269);
nand U34634 (N_34634,N_29077,N_20711);
xor U34635 (N_34635,N_29216,N_27833);
xnor U34636 (N_34636,N_29557,N_26100);
xnor U34637 (N_34637,N_20245,N_24704);
nand U34638 (N_34638,N_24324,N_23344);
and U34639 (N_34639,N_26655,N_25334);
xor U34640 (N_34640,N_23018,N_22767);
and U34641 (N_34641,N_22244,N_26852);
nand U34642 (N_34642,N_26754,N_23419);
nand U34643 (N_34643,N_26787,N_24386);
nand U34644 (N_34644,N_24980,N_22135);
and U34645 (N_34645,N_29480,N_29515);
nand U34646 (N_34646,N_29519,N_25495);
xnor U34647 (N_34647,N_21507,N_23651);
nand U34648 (N_34648,N_22050,N_21832);
and U34649 (N_34649,N_26159,N_21235);
xor U34650 (N_34650,N_23349,N_22509);
xnor U34651 (N_34651,N_26097,N_28285);
or U34652 (N_34652,N_28925,N_21326);
nand U34653 (N_34653,N_24971,N_21294);
or U34654 (N_34654,N_23500,N_28109);
nor U34655 (N_34655,N_29951,N_29904);
and U34656 (N_34656,N_29962,N_23217);
nor U34657 (N_34657,N_24846,N_21867);
and U34658 (N_34658,N_26533,N_22668);
and U34659 (N_34659,N_27189,N_24454);
and U34660 (N_34660,N_24965,N_28100);
xor U34661 (N_34661,N_23437,N_29185);
nand U34662 (N_34662,N_24413,N_23007);
or U34663 (N_34663,N_26768,N_23343);
or U34664 (N_34664,N_29971,N_25398);
nor U34665 (N_34665,N_29474,N_23769);
xor U34666 (N_34666,N_29521,N_20995);
nand U34667 (N_34667,N_28540,N_28608);
or U34668 (N_34668,N_29616,N_23703);
xnor U34669 (N_34669,N_24670,N_24610);
nor U34670 (N_34670,N_23657,N_29381);
nor U34671 (N_34671,N_25147,N_27177);
nor U34672 (N_34672,N_27445,N_26223);
xor U34673 (N_34673,N_24146,N_24886);
nor U34674 (N_34674,N_21839,N_23655);
and U34675 (N_34675,N_26513,N_25385);
xnor U34676 (N_34676,N_26634,N_26644);
xnor U34677 (N_34677,N_26545,N_24543);
nand U34678 (N_34678,N_23987,N_27526);
and U34679 (N_34679,N_23904,N_22094);
and U34680 (N_34680,N_22891,N_21640);
nand U34681 (N_34681,N_21393,N_22580);
nand U34682 (N_34682,N_23836,N_24910);
nand U34683 (N_34683,N_23502,N_27933);
and U34684 (N_34684,N_26595,N_22551);
xor U34685 (N_34685,N_27287,N_27179);
nor U34686 (N_34686,N_29675,N_28812);
nor U34687 (N_34687,N_27017,N_29319);
or U34688 (N_34688,N_28488,N_20190);
nor U34689 (N_34689,N_24518,N_28692);
or U34690 (N_34690,N_21853,N_28145);
nand U34691 (N_34691,N_22241,N_22847);
nand U34692 (N_34692,N_20068,N_20693);
xor U34693 (N_34693,N_20370,N_24728);
or U34694 (N_34694,N_28390,N_25353);
xor U34695 (N_34695,N_29772,N_21277);
or U34696 (N_34696,N_20616,N_26328);
xnor U34697 (N_34697,N_26098,N_25380);
nand U34698 (N_34698,N_24201,N_29670);
nand U34699 (N_34699,N_26147,N_26548);
and U34700 (N_34700,N_24922,N_20334);
and U34701 (N_34701,N_25817,N_25337);
or U34702 (N_34702,N_20763,N_23902);
and U34703 (N_34703,N_22821,N_23182);
nor U34704 (N_34704,N_23980,N_29939);
nand U34705 (N_34705,N_23218,N_29537);
or U34706 (N_34706,N_27981,N_23057);
xor U34707 (N_34707,N_22895,N_28854);
and U34708 (N_34708,N_22015,N_20207);
and U34709 (N_34709,N_28077,N_24016);
xnor U34710 (N_34710,N_28741,N_20261);
nand U34711 (N_34711,N_22328,N_25957);
xor U34712 (N_34712,N_27372,N_22666);
nor U34713 (N_34713,N_24537,N_29631);
or U34714 (N_34714,N_29408,N_26099);
nor U34715 (N_34715,N_20060,N_23702);
nand U34716 (N_34716,N_24702,N_21627);
and U34717 (N_34717,N_26767,N_27006);
xor U34718 (N_34718,N_24889,N_29269);
and U34719 (N_34719,N_22938,N_26093);
and U34720 (N_34720,N_28497,N_28449);
nand U34721 (N_34721,N_23831,N_22952);
nor U34722 (N_34722,N_20488,N_24854);
or U34723 (N_34723,N_25825,N_25663);
nor U34724 (N_34724,N_27299,N_20605);
or U34725 (N_34725,N_24990,N_28805);
xnor U34726 (N_34726,N_21191,N_24287);
or U34727 (N_34727,N_28128,N_26436);
xnor U34728 (N_34728,N_29128,N_25352);
nor U34729 (N_34729,N_22661,N_20125);
nand U34730 (N_34730,N_26417,N_25801);
or U34731 (N_34731,N_23469,N_22500);
nor U34732 (N_34732,N_29887,N_27573);
xor U34733 (N_34733,N_24361,N_26332);
or U34734 (N_34734,N_26075,N_29523);
xnor U34735 (N_34735,N_20689,N_28133);
nand U34736 (N_34736,N_21700,N_21885);
xor U34737 (N_34737,N_21882,N_20710);
nand U34738 (N_34738,N_24569,N_23909);
and U34739 (N_34739,N_27766,N_27798);
xor U34740 (N_34740,N_20123,N_27091);
xor U34741 (N_34741,N_20955,N_23757);
and U34742 (N_34742,N_22966,N_22319);
nand U34743 (N_34743,N_21174,N_21158);
and U34744 (N_34744,N_27565,N_21622);
xor U34745 (N_34745,N_21638,N_23789);
xor U34746 (N_34746,N_24464,N_23766);
or U34747 (N_34747,N_23317,N_21205);
nand U34748 (N_34748,N_26965,N_29619);
xnor U34749 (N_34749,N_26962,N_26324);
and U34750 (N_34750,N_28013,N_26251);
nand U34751 (N_34751,N_23528,N_25234);
nand U34752 (N_34752,N_23876,N_29773);
xor U34753 (N_34753,N_20058,N_21022);
nand U34754 (N_34754,N_29031,N_27680);
nor U34755 (N_34755,N_29337,N_27168);
xnor U34756 (N_34756,N_28030,N_29633);
xor U34757 (N_34757,N_25503,N_22549);
and U34758 (N_34758,N_21585,N_29132);
nand U34759 (N_34759,N_27354,N_21289);
nand U34760 (N_34760,N_25273,N_21985);
and U34761 (N_34761,N_21336,N_29309);
nand U34762 (N_34762,N_21008,N_22747);
nand U34763 (N_34763,N_29754,N_24290);
nand U34764 (N_34764,N_26338,N_21466);
or U34765 (N_34765,N_22451,N_27164);
or U34766 (N_34766,N_27830,N_29421);
nor U34767 (N_34767,N_22426,N_22235);
or U34768 (N_34768,N_24839,N_22819);
xnor U34769 (N_34769,N_21663,N_25662);
and U34770 (N_34770,N_20732,N_25576);
nand U34771 (N_34771,N_27721,N_21576);
nand U34772 (N_34772,N_25733,N_22399);
nand U34773 (N_34773,N_21992,N_20291);
nor U34774 (N_34774,N_25056,N_28022);
and U34775 (N_34775,N_21758,N_28123);
and U34776 (N_34776,N_24981,N_24185);
xnor U34777 (N_34777,N_27021,N_28201);
and U34778 (N_34778,N_29226,N_25127);
nor U34779 (N_34779,N_20227,N_25865);
nor U34780 (N_34780,N_29144,N_20188);
nand U34781 (N_34781,N_23152,N_25306);
and U34782 (N_34782,N_22101,N_23198);
nor U34783 (N_34783,N_24756,N_25347);
nand U34784 (N_34784,N_28053,N_23759);
nor U34785 (N_34785,N_21778,N_27074);
nor U34786 (N_34786,N_20586,N_27675);
nand U34787 (N_34787,N_29756,N_25746);
nor U34788 (N_34788,N_23289,N_24698);
nand U34789 (N_34789,N_27630,N_25924);
xnor U34790 (N_34790,N_22081,N_21096);
nand U34791 (N_34791,N_28684,N_27783);
or U34792 (N_34792,N_21626,N_29248);
nand U34793 (N_34793,N_21645,N_20577);
nand U34794 (N_34794,N_29908,N_27462);
or U34795 (N_34795,N_20671,N_24333);
nor U34796 (N_34796,N_26363,N_23632);
and U34797 (N_34797,N_23798,N_27749);
xnor U34798 (N_34798,N_27967,N_25402);
nand U34799 (N_34799,N_27875,N_25584);
nand U34800 (N_34800,N_25600,N_26643);
nand U34801 (N_34801,N_29262,N_21529);
or U34802 (N_34802,N_20456,N_29343);
nor U34803 (N_34803,N_21495,N_26727);
and U34804 (N_34804,N_26605,N_27010);
and U34805 (N_34805,N_27658,N_25633);
nor U34806 (N_34806,N_24572,N_27773);
nand U34807 (N_34807,N_23295,N_29302);
or U34808 (N_34808,N_26798,N_22873);
xnor U34809 (N_34809,N_23746,N_26134);
nor U34810 (N_34810,N_27375,N_22764);
or U34811 (N_34811,N_23115,N_24792);
xor U34812 (N_34812,N_25930,N_23522);
nand U34813 (N_34813,N_23250,N_20608);
nand U34814 (N_34814,N_29349,N_25028);
and U34815 (N_34815,N_20928,N_28482);
nor U34816 (N_34816,N_29393,N_21967);
and U34817 (N_34817,N_23615,N_24745);
nand U34818 (N_34818,N_27488,N_25641);
nor U34819 (N_34819,N_27747,N_25696);
or U34820 (N_34820,N_24042,N_21035);
nor U34821 (N_34821,N_21952,N_23866);
or U34822 (N_34822,N_28226,N_22171);
xor U34823 (N_34823,N_27601,N_20290);
and U34824 (N_34824,N_28819,N_26434);
or U34825 (N_34825,N_23360,N_25304);
and U34826 (N_34826,N_28086,N_25047);
xor U34827 (N_34827,N_21883,N_23251);
nand U34828 (N_34828,N_20668,N_29419);
nand U34829 (N_34829,N_22210,N_24223);
and U34830 (N_34830,N_28900,N_23917);
or U34831 (N_34831,N_22249,N_25677);
or U34832 (N_34832,N_23056,N_28673);
nand U34833 (N_34833,N_28914,N_29250);
or U34834 (N_34834,N_22266,N_26668);
or U34835 (N_34835,N_23477,N_29107);
or U34836 (N_34836,N_28107,N_20707);
or U34837 (N_34837,N_23225,N_21286);
nor U34838 (N_34838,N_24087,N_20562);
or U34839 (N_34839,N_28282,N_25129);
nor U34840 (N_34840,N_26996,N_20667);
or U34841 (N_34841,N_25719,N_28356);
xnor U34842 (N_34842,N_27482,N_21354);
and U34843 (N_34843,N_28213,N_22606);
nor U34844 (N_34844,N_24765,N_20317);
nand U34845 (N_34845,N_25608,N_28744);
xnor U34846 (N_34846,N_21699,N_28198);
or U34847 (N_34847,N_23994,N_25323);
and U34848 (N_34848,N_20332,N_25565);
nor U34849 (N_34849,N_27996,N_29174);
nor U34850 (N_34850,N_21478,N_24638);
nor U34851 (N_34851,N_29372,N_29996);
or U34852 (N_34852,N_25143,N_25550);
nor U34853 (N_34853,N_24325,N_28154);
nand U34854 (N_34854,N_21844,N_25365);
xnor U34855 (N_34855,N_23332,N_22237);
nand U34856 (N_34856,N_22046,N_26828);
xnor U34857 (N_34857,N_29874,N_24579);
or U34858 (N_34858,N_23235,N_20401);
and U34859 (N_34859,N_27506,N_25718);
nor U34860 (N_34860,N_26822,N_27931);
nand U34861 (N_34861,N_25089,N_21132);
nand U34862 (N_34862,N_29033,N_28297);
or U34863 (N_34863,N_28514,N_28830);
and U34864 (N_34864,N_23664,N_20233);
and U34865 (N_34865,N_20304,N_25396);
and U34866 (N_34866,N_23211,N_20414);
xor U34867 (N_34867,N_20980,N_21187);
nor U34868 (N_34868,N_26346,N_20170);
and U34869 (N_34869,N_28590,N_26825);
xor U34870 (N_34870,N_29964,N_22765);
or U34871 (N_34871,N_20565,N_24520);
and U34872 (N_34872,N_23489,N_29549);
xor U34873 (N_34873,N_27484,N_24938);
and U34874 (N_34874,N_20306,N_29406);
and U34875 (N_34875,N_21196,N_23112);
or U34876 (N_34876,N_23162,N_23234);
xnor U34877 (N_34877,N_22028,N_20092);
and U34878 (N_34878,N_20672,N_24319);
nand U34879 (N_34879,N_24298,N_28096);
or U34880 (N_34880,N_25517,N_20110);
and U34881 (N_34881,N_20956,N_27946);
nor U34882 (N_34882,N_24082,N_20704);
and U34883 (N_34883,N_27804,N_27139);
or U34884 (N_34884,N_20941,N_26005);
xor U34885 (N_34885,N_28319,N_22491);
or U34886 (N_34886,N_29301,N_20912);
xnor U34887 (N_34887,N_27414,N_25145);
or U34888 (N_34888,N_22706,N_21492);
xor U34889 (N_34889,N_22513,N_28507);
nor U34890 (N_34890,N_21195,N_28463);
or U34891 (N_34891,N_22972,N_22085);
nor U34892 (N_34892,N_20299,N_29291);
nor U34893 (N_34893,N_29645,N_29505);
or U34894 (N_34894,N_25475,N_20408);
xnor U34895 (N_34895,N_29830,N_20688);
xor U34896 (N_34896,N_29470,N_22680);
xor U34897 (N_34897,N_24964,N_27042);
or U34898 (N_34898,N_23126,N_20654);
xor U34899 (N_34899,N_26329,N_22256);
nor U34900 (N_34900,N_23722,N_22949);
and U34901 (N_34901,N_21898,N_21659);
nor U34902 (N_34902,N_22452,N_21192);
and U34903 (N_34903,N_22934,N_29598);
and U34904 (N_34904,N_29288,N_21720);
xor U34905 (N_34905,N_21269,N_21791);
nand U34906 (N_34906,N_25448,N_23882);
nand U34907 (N_34907,N_20581,N_21688);
or U34908 (N_34908,N_29457,N_24136);
xnor U34909 (N_34909,N_24285,N_21092);
and U34910 (N_34910,N_23895,N_27470);
xnor U34911 (N_34911,N_22654,N_25772);
xor U34912 (N_34912,N_27970,N_25451);
or U34913 (N_34913,N_23376,N_28917);
or U34914 (N_34914,N_29001,N_21987);
xor U34915 (N_34915,N_24531,N_25477);
nor U34916 (N_34916,N_22751,N_26317);
or U34917 (N_34917,N_22358,N_29241);
or U34918 (N_34918,N_22833,N_26252);
and U34919 (N_34919,N_29212,N_27992);
nor U34920 (N_34920,N_20483,N_29484);
nor U34921 (N_34921,N_22761,N_28651);
xnor U34922 (N_34922,N_23361,N_21271);
xnor U34923 (N_34923,N_23784,N_25088);
nor U34924 (N_34924,N_28808,N_26245);
nor U34925 (N_34925,N_26342,N_27748);
nand U34926 (N_34926,N_23050,N_22361);
or U34927 (N_34927,N_21567,N_27919);
xor U34928 (N_34928,N_28318,N_22295);
xnor U34929 (N_34929,N_25051,N_20872);
nor U34930 (N_34930,N_27246,N_27644);
nor U34931 (N_34931,N_26187,N_26993);
xor U34932 (N_34932,N_22750,N_22936);
or U34933 (N_34933,N_27370,N_20519);
nand U34934 (N_34934,N_23815,N_23254);
nor U34935 (N_34935,N_25642,N_21948);
xor U34936 (N_34936,N_27613,N_26181);
or U34937 (N_34937,N_22263,N_20168);
nor U34938 (N_34938,N_21366,N_26184);
nand U34939 (N_34939,N_26188,N_28971);
xnor U34940 (N_34940,N_22234,N_26810);
or U34941 (N_34941,N_28752,N_26185);
or U34942 (N_34942,N_25997,N_23595);
xor U34943 (N_34943,N_21190,N_24126);
and U34944 (N_34944,N_25866,N_28951);
nand U34945 (N_34945,N_28648,N_21078);
nor U34946 (N_34946,N_21756,N_20595);
xor U34947 (N_34947,N_25735,N_24871);
and U34948 (N_34948,N_22378,N_26066);
nor U34949 (N_34949,N_28632,N_27397);
or U34950 (N_34950,N_29895,N_24743);
nand U34951 (N_34951,N_24036,N_20274);
xnor U34952 (N_34952,N_23462,N_27661);
nand U34953 (N_34953,N_22793,N_22503);
nor U34954 (N_34954,N_29299,N_22181);
nor U34955 (N_34955,N_26176,N_28233);
nor U34956 (N_34956,N_22876,N_25533);
and U34957 (N_34957,N_28689,N_21219);
nand U34958 (N_34958,N_28897,N_22332);
and U34959 (N_34959,N_27545,N_25793);
or U34960 (N_34960,N_21275,N_24038);
or U34961 (N_34961,N_29339,N_21551);
or U34962 (N_34962,N_26856,N_26724);
nand U34963 (N_34963,N_24058,N_20927);
or U34964 (N_34964,N_24594,N_21748);
nand U34965 (N_34965,N_25569,N_22018);
nor U34966 (N_34966,N_22594,N_29671);
and U34967 (N_34967,N_29300,N_26265);
nor U34968 (N_34968,N_25686,N_26301);
or U34969 (N_34969,N_29790,N_22998);
nand U34970 (N_34970,N_29828,N_25986);
xnor U34971 (N_34971,N_21029,N_21706);
and U34972 (N_34972,N_27490,N_24853);
or U34973 (N_34973,N_20133,N_21675);
and U34974 (N_34974,N_27627,N_28557);
nor U34975 (N_34975,N_28087,N_25138);
nand U34976 (N_34976,N_25408,N_25535);
nor U34977 (N_34977,N_27280,N_28028);
xnor U34978 (N_34978,N_26612,N_20405);
and U34979 (N_34979,N_28152,N_27014);
and U34980 (N_34980,N_24431,N_22149);
nand U34981 (N_34981,N_21572,N_24360);
or U34982 (N_34982,N_26010,N_23892);
or U34983 (N_34983,N_29057,N_26069);
xor U34984 (N_34984,N_22083,N_27132);
nor U34985 (N_34985,N_25343,N_26220);
or U34986 (N_34986,N_28881,N_20804);
nand U34987 (N_34987,N_22902,N_26057);
nor U34988 (N_34988,N_29353,N_29106);
nor U34989 (N_34989,N_23686,N_25309);
nor U34990 (N_34990,N_28967,N_29427);
or U34991 (N_34991,N_26222,N_21527);
nand U34992 (N_34992,N_21091,N_28150);
nor U34993 (N_34993,N_28434,N_25123);
xor U34994 (N_34994,N_23461,N_22613);
and U34995 (N_34995,N_28039,N_26200);
xnor U34996 (N_34996,N_24685,N_25716);
xor U34997 (N_34997,N_24119,N_28989);
or U34998 (N_34998,N_28528,N_20445);
nand U34999 (N_34999,N_27054,N_23633);
xor U35000 (N_35000,N_23060,N_29166);
nor U35001 (N_35001,N_29236,N_23303);
xnor U35002 (N_35002,N_22585,N_21847);
xor U35003 (N_35003,N_20701,N_27120);
or U35004 (N_35004,N_24308,N_23267);
xnor U35005 (N_35005,N_28190,N_26406);
or U35006 (N_35006,N_27419,N_28698);
nor U35007 (N_35007,N_24587,N_26527);
xor U35008 (N_35008,N_21217,N_26211);
xnor U35009 (N_35009,N_24297,N_27288);
nor U35010 (N_35010,N_25978,N_26334);
or U35011 (N_35011,N_25766,N_26986);
xor U35012 (N_35012,N_20162,N_24421);
or U35013 (N_35013,N_29574,N_20224);
xnor U35014 (N_35014,N_21628,N_27883);
and U35015 (N_35015,N_25173,N_29136);
xnor U35016 (N_35016,N_25904,N_22779);
xor U35017 (N_35017,N_23502,N_25481);
and U35018 (N_35018,N_21308,N_26406);
nor U35019 (N_35019,N_22983,N_29854);
xor U35020 (N_35020,N_28296,N_28521);
nand U35021 (N_35021,N_25700,N_23055);
nand U35022 (N_35022,N_28515,N_25807);
or U35023 (N_35023,N_25037,N_20436);
nand U35024 (N_35024,N_23994,N_21307);
nor U35025 (N_35025,N_20587,N_27971);
and U35026 (N_35026,N_22497,N_21832);
or U35027 (N_35027,N_26933,N_21920);
nand U35028 (N_35028,N_28272,N_22861);
nor U35029 (N_35029,N_29995,N_29721);
nor U35030 (N_35030,N_27351,N_25907);
nor U35031 (N_35031,N_26080,N_20890);
nand U35032 (N_35032,N_22853,N_28463);
xnor U35033 (N_35033,N_23180,N_25509);
or U35034 (N_35034,N_26816,N_28608);
xnor U35035 (N_35035,N_20387,N_28533);
xnor U35036 (N_35036,N_27181,N_24889);
xor U35037 (N_35037,N_20896,N_22565);
nor U35038 (N_35038,N_22810,N_24627);
or U35039 (N_35039,N_28215,N_27714);
nand U35040 (N_35040,N_22799,N_28897);
or U35041 (N_35041,N_23859,N_25013);
nor U35042 (N_35042,N_21918,N_28897);
nand U35043 (N_35043,N_20026,N_27257);
xnor U35044 (N_35044,N_26636,N_21278);
or U35045 (N_35045,N_23464,N_24829);
or U35046 (N_35046,N_23278,N_22954);
nor U35047 (N_35047,N_23782,N_22968);
and U35048 (N_35048,N_25008,N_23206);
nand U35049 (N_35049,N_27934,N_21716);
xor U35050 (N_35050,N_20795,N_22430);
nor U35051 (N_35051,N_28452,N_27246);
and U35052 (N_35052,N_29800,N_22948);
nand U35053 (N_35053,N_21214,N_21022);
or U35054 (N_35054,N_23518,N_25122);
and U35055 (N_35055,N_27735,N_20082);
or U35056 (N_35056,N_22251,N_29719);
or U35057 (N_35057,N_29998,N_28388);
or U35058 (N_35058,N_20859,N_23583);
nand U35059 (N_35059,N_23667,N_28193);
nor U35060 (N_35060,N_24767,N_28161);
xor U35061 (N_35061,N_21976,N_24117);
and U35062 (N_35062,N_21801,N_24298);
nor U35063 (N_35063,N_29169,N_28347);
xor U35064 (N_35064,N_22708,N_21071);
nand U35065 (N_35065,N_24739,N_28217);
xnor U35066 (N_35066,N_26934,N_23269);
nor U35067 (N_35067,N_23613,N_28715);
nor U35068 (N_35068,N_20272,N_25228);
nand U35069 (N_35069,N_24101,N_22428);
nor U35070 (N_35070,N_26895,N_20258);
nand U35071 (N_35071,N_25112,N_21283);
xor U35072 (N_35072,N_29463,N_21060);
nand U35073 (N_35073,N_25011,N_22095);
and U35074 (N_35074,N_26222,N_24005);
nor U35075 (N_35075,N_24248,N_29978);
nor U35076 (N_35076,N_28564,N_26289);
or U35077 (N_35077,N_28728,N_29670);
xnor U35078 (N_35078,N_28590,N_26398);
nor U35079 (N_35079,N_27587,N_28542);
xnor U35080 (N_35080,N_29537,N_27121);
or U35081 (N_35081,N_23284,N_24157);
and U35082 (N_35082,N_22678,N_27667);
and U35083 (N_35083,N_25468,N_27739);
or U35084 (N_35084,N_20810,N_28983);
nand U35085 (N_35085,N_24920,N_26545);
nor U35086 (N_35086,N_25310,N_25344);
xor U35087 (N_35087,N_26160,N_28066);
or U35088 (N_35088,N_21095,N_24898);
or U35089 (N_35089,N_29699,N_25232);
nor U35090 (N_35090,N_22110,N_27035);
nand U35091 (N_35091,N_26844,N_28834);
or U35092 (N_35092,N_28150,N_27171);
nor U35093 (N_35093,N_24389,N_22273);
nor U35094 (N_35094,N_27046,N_21851);
xnor U35095 (N_35095,N_25894,N_24646);
nor U35096 (N_35096,N_28323,N_23489);
and U35097 (N_35097,N_25517,N_24540);
xnor U35098 (N_35098,N_22237,N_24909);
xnor U35099 (N_35099,N_28625,N_25618);
or U35100 (N_35100,N_20068,N_21248);
or U35101 (N_35101,N_21521,N_20322);
nand U35102 (N_35102,N_25751,N_21915);
xor U35103 (N_35103,N_23055,N_20422);
xnor U35104 (N_35104,N_29192,N_20380);
and U35105 (N_35105,N_21043,N_29326);
nand U35106 (N_35106,N_23771,N_22571);
and U35107 (N_35107,N_23527,N_26463);
and U35108 (N_35108,N_21517,N_26556);
nor U35109 (N_35109,N_29162,N_27334);
nor U35110 (N_35110,N_21500,N_29530);
xnor U35111 (N_35111,N_24592,N_21379);
xor U35112 (N_35112,N_21725,N_20228);
nor U35113 (N_35113,N_28000,N_28793);
nand U35114 (N_35114,N_25860,N_21222);
xor U35115 (N_35115,N_28363,N_26185);
and U35116 (N_35116,N_23938,N_29358);
nand U35117 (N_35117,N_24041,N_28755);
or U35118 (N_35118,N_29269,N_20907);
xnor U35119 (N_35119,N_29720,N_24088);
and U35120 (N_35120,N_21783,N_22872);
and U35121 (N_35121,N_21553,N_27722);
and U35122 (N_35122,N_21286,N_26094);
or U35123 (N_35123,N_27042,N_26674);
nor U35124 (N_35124,N_29496,N_28505);
and U35125 (N_35125,N_20412,N_23577);
or U35126 (N_35126,N_21819,N_25864);
nand U35127 (N_35127,N_28111,N_28138);
nor U35128 (N_35128,N_25650,N_21928);
and U35129 (N_35129,N_25303,N_21370);
and U35130 (N_35130,N_21568,N_29364);
or U35131 (N_35131,N_20906,N_26321);
nand U35132 (N_35132,N_27529,N_21580);
and U35133 (N_35133,N_20594,N_28459);
and U35134 (N_35134,N_29808,N_22032);
xnor U35135 (N_35135,N_21317,N_24291);
xor U35136 (N_35136,N_27448,N_28639);
xnor U35137 (N_35137,N_28488,N_27276);
or U35138 (N_35138,N_27848,N_20391);
or U35139 (N_35139,N_22460,N_24231);
and U35140 (N_35140,N_22248,N_26484);
and U35141 (N_35141,N_27347,N_24011);
or U35142 (N_35142,N_23628,N_22518);
and U35143 (N_35143,N_26998,N_28592);
nor U35144 (N_35144,N_22590,N_28276);
nand U35145 (N_35145,N_28205,N_24222);
xor U35146 (N_35146,N_22057,N_22089);
or U35147 (N_35147,N_21105,N_26454);
nand U35148 (N_35148,N_24105,N_25710);
and U35149 (N_35149,N_27187,N_21799);
nor U35150 (N_35150,N_28442,N_26192);
xnor U35151 (N_35151,N_25919,N_26084);
nand U35152 (N_35152,N_20557,N_21362);
xor U35153 (N_35153,N_25028,N_23740);
xnor U35154 (N_35154,N_28926,N_28053);
and U35155 (N_35155,N_21987,N_27015);
and U35156 (N_35156,N_22898,N_22998);
or U35157 (N_35157,N_22720,N_21782);
xnor U35158 (N_35158,N_22342,N_29328);
nor U35159 (N_35159,N_27123,N_24012);
or U35160 (N_35160,N_27997,N_27912);
and U35161 (N_35161,N_26709,N_22143);
or U35162 (N_35162,N_25209,N_24639);
or U35163 (N_35163,N_22112,N_22613);
or U35164 (N_35164,N_20000,N_20672);
or U35165 (N_35165,N_23656,N_24000);
nand U35166 (N_35166,N_21093,N_24697);
nand U35167 (N_35167,N_23237,N_22645);
nor U35168 (N_35168,N_20817,N_29472);
nand U35169 (N_35169,N_25987,N_23997);
nand U35170 (N_35170,N_27808,N_21212);
xor U35171 (N_35171,N_23820,N_23500);
xnor U35172 (N_35172,N_22666,N_29857);
xor U35173 (N_35173,N_20442,N_23988);
xnor U35174 (N_35174,N_25680,N_23127);
and U35175 (N_35175,N_21910,N_27907);
and U35176 (N_35176,N_29647,N_29488);
and U35177 (N_35177,N_26301,N_28510);
and U35178 (N_35178,N_20473,N_23462);
nand U35179 (N_35179,N_24096,N_24399);
nor U35180 (N_35180,N_26667,N_20906);
nand U35181 (N_35181,N_21464,N_28247);
nor U35182 (N_35182,N_27392,N_29355);
and U35183 (N_35183,N_27990,N_27138);
xnor U35184 (N_35184,N_21895,N_22384);
nor U35185 (N_35185,N_22228,N_20350);
nor U35186 (N_35186,N_21543,N_23888);
and U35187 (N_35187,N_23644,N_25658);
nor U35188 (N_35188,N_24579,N_25226);
xor U35189 (N_35189,N_27251,N_27559);
or U35190 (N_35190,N_27300,N_25404);
nand U35191 (N_35191,N_27242,N_29251);
xor U35192 (N_35192,N_28668,N_21686);
xor U35193 (N_35193,N_22026,N_25451);
xnor U35194 (N_35194,N_22884,N_20192);
nand U35195 (N_35195,N_21014,N_26793);
or U35196 (N_35196,N_26793,N_22837);
nor U35197 (N_35197,N_22358,N_20493);
or U35198 (N_35198,N_29289,N_29989);
or U35199 (N_35199,N_25627,N_26586);
nand U35200 (N_35200,N_25669,N_29452);
or U35201 (N_35201,N_23609,N_24300);
and U35202 (N_35202,N_20759,N_25845);
and U35203 (N_35203,N_21658,N_25567);
or U35204 (N_35204,N_26526,N_26134);
or U35205 (N_35205,N_25672,N_25293);
xor U35206 (N_35206,N_20980,N_21031);
xnor U35207 (N_35207,N_27157,N_25560);
nor U35208 (N_35208,N_20092,N_24925);
and U35209 (N_35209,N_29074,N_22574);
nor U35210 (N_35210,N_26176,N_22294);
nor U35211 (N_35211,N_28570,N_28449);
and U35212 (N_35212,N_24245,N_26161);
or U35213 (N_35213,N_21350,N_27323);
or U35214 (N_35214,N_24107,N_22808);
nor U35215 (N_35215,N_23562,N_27514);
nor U35216 (N_35216,N_26856,N_23566);
or U35217 (N_35217,N_29008,N_27454);
nor U35218 (N_35218,N_27018,N_28261);
nand U35219 (N_35219,N_27206,N_29371);
xor U35220 (N_35220,N_22436,N_20651);
and U35221 (N_35221,N_26322,N_21309);
nor U35222 (N_35222,N_24603,N_28073);
nand U35223 (N_35223,N_21261,N_28498);
nand U35224 (N_35224,N_25095,N_25814);
nor U35225 (N_35225,N_26359,N_23177);
nand U35226 (N_35226,N_21154,N_29631);
or U35227 (N_35227,N_27690,N_28088);
or U35228 (N_35228,N_29721,N_21221);
nand U35229 (N_35229,N_29156,N_27483);
or U35230 (N_35230,N_20450,N_25250);
nor U35231 (N_35231,N_27970,N_20298);
nand U35232 (N_35232,N_28009,N_22335);
nor U35233 (N_35233,N_28807,N_24894);
nor U35234 (N_35234,N_24328,N_25364);
or U35235 (N_35235,N_24279,N_21367);
xor U35236 (N_35236,N_21882,N_21674);
nor U35237 (N_35237,N_23857,N_24287);
or U35238 (N_35238,N_26447,N_23075);
nand U35239 (N_35239,N_28135,N_22019);
or U35240 (N_35240,N_29139,N_27694);
nor U35241 (N_35241,N_29119,N_24718);
nor U35242 (N_35242,N_21253,N_28921);
nor U35243 (N_35243,N_22164,N_29485);
or U35244 (N_35244,N_29521,N_28038);
or U35245 (N_35245,N_25748,N_21058);
and U35246 (N_35246,N_23918,N_23429);
and U35247 (N_35247,N_29168,N_27809);
nor U35248 (N_35248,N_20735,N_20330);
nor U35249 (N_35249,N_21519,N_25575);
xor U35250 (N_35250,N_22007,N_21701);
nand U35251 (N_35251,N_28571,N_22446);
nor U35252 (N_35252,N_22081,N_29973);
or U35253 (N_35253,N_20250,N_27600);
xor U35254 (N_35254,N_24358,N_25969);
and U35255 (N_35255,N_24830,N_21438);
xor U35256 (N_35256,N_25109,N_22317);
and U35257 (N_35257,N_28972,N_22773);
nor U35258 (N_35258,N_27113,N_20237);
nand U35259 (N_35259,N_20173,N_20963);
nor U35260 (N_35260,N_22745,N_24190);
xnor U35261 (N_35261,N_26347,N_25051);
nor U35262 (N_35262,N_26826,N_22695);
xnor U35263 (N_35263,N_25744,N_27787);
xnor U35264 (N_35264,N_26425,N_20846);
nand U35265 (N_35265,N_27608,N_23805);
or U35266 (N_35266,N_24188,N_27327);
and U35267 (N_35267,N_27436,N_29782);
xor U35268 (N_35268,N_29023,N_24636);
nand U35269 (N_35269,N_24317,N_20215);
nor U35270 (N_35270,N_25852,N_21578);
nor U35271 (N_35271,N_28516,N_21122);
nor U35272 (N_35272,N_23855,N_23578);
and U35273 (N_35273,N_29939,N_24920);
and U35274 (N_35274,N_22908,N_24268);
and U35275 (N_35275,N_28041,N_24317);
nor U35276 (N_35276,N_21247,N_21378);
and U35277 (N_35277,N_24044,N_20494);
nand U35278 (N_35278,N_29464,N_25439);
or U35279 (N_35279,N_21486,N_23457);
or U35280 (N_35280,N_23447,N_26316);
nand U35281 (N_35281,N_20115,N_24989);
xnor U35282 (N_35282,N_28991,N_25651);
or U35283 (N_35283,N_20362,N_28827);
nor U35284 (N_35284,N_26336,N_29954);
xnor U35285 (N_35285,N_25817,N_23252);
xnor U35286 (N_35286,N_25988,N_23182);
and U35287 (N_35287,N_20164,N_25418);
or U35288 (N_35288,N_29316,N_24995);
and U35289 (N_35289,N_26956,N_26176);
and U35290 (N_35290,N_25941,N_22424);
and U35291 (N_35291,N_20748,N_28231);
nor U35292 (N_35292,N_25311,N_20028);
xnor U35293 (N_35293,N_23788,N_25444);
and U35294 (N_35294,N_28536,N_23287);
nand U35295 (N_35295,N_22329,N_21067);
nor U35296 (N_35296,N_22874,N_29960);
and U35297 (N_35297,N_26873,N_26863);
nor U35298 (N_35298,N_22473,N_27590);
nand U35299 (N_35299,N_26722,N_24513);
nor U35300 (N_35300,N_28148,N_21402);
nor U35301 (N_35301,N_24027,N_20887);
nand U35302 (N_35302,N_21404,N_28878);
nand U35303 (N_35303,N_24386,N_28090);
xnor U35304 (N_35304,N_29264,N_21919);
xor U35305 (N_35305,N_24862,N_20404);
nand U35306 (N_35306,N_21228,N_21148);
nor U35307 (N_35307,N_21114,N_25146);
nand U35308 (N_35308,N_29553,N_26839);
nor U35309 (N_35309,N_27686,N_25846);
nand U35310 (N_35310,N_28731,N_25263);
nand U35311 (N_35311,N_27642,N_28320);
nor U35312 (N_35312,N_28643,N_28909);
xnor U35313 (N_35313,N_26581,N_22081);
or U35314 (N_35314,N_26082,N_21017);
xor U35315 (N_35315,N_21478,N_22129);
xor U35316 (N_35316,N_27947,N_25866);
or U35317 (N_35317,N_27140,N_25913);
nand U35318 (N_35318,N_25745,N_28316);
or U35319 (N_35319,N_25514,N_23867);
xnor U35320 (N_35320,N_21242,N_28809);
xor U35321 (N_35321,N_26193,N_25039);
nand U35322 (N_35322,N_25606,N_27514);
or U35323 (N_35323,N_25686,N_27348);
nand U35324 (N_35324,N_24830,N_26825);
and U35325 (N_35325,N_24364,N_23327);
nor U35326 (N_35326,N_26024,N_27271);
xor U35327 (N_35327,N_29117,N_24313);
and U35328 (N_35328,N_23666,N_20540);
nor U35329 (N_35329,N_28017,N_21510);
xnor U35330 (N_35330,N_23893,N_22232);
or U35331 (N_35331,N_23231,N_29833);
nor U35332 (N_35332,N_23360,N_25626);
nor U35333 (N_35333,N_23768,N_24104);
and U35334 (N_35334,N_24813,N_29302);
xnor U35335 (N_35335,N_21077,N_25090);
and U35336 (N_35336,N_28341,N_24711);
nor U35337 (N_35337,N_25588,N_24769);
nand U35338 (N_35338,N_28079,N_21444);
and U35339 (N_35339,N_21752,N_29228);
nand U35340 (N_35340,N_22756,N_20115);
and U35341 (N_35341,N_22732,N_27137);
xor U35342 (N_35342,N_23215,N_26714);
nor U35343 (N_35343,N_29556,N_23122);
nand U35344 (N_35344,N_24678,N_29889);
and U35345 (N_35345,N_22184,N_20830);
nand U35346 (N_35346,N_23697,N_25803);
nor U35347 (N_35347,N_27688,N_25193);
nor U35348 (N_35348,N_23842,N_24777);
and U35349 (N_35349,N_22854,N_22013);
or U35350 (N_35350,N_27526,N_23281);
or U35351 (N_35351,N_21450,N_25875);
xor U35352 (N_35352,N_26341,N_20194);
or U35353 (N_35353,N_28812,N_20469);
and U35354 (N_35354,N_25599,N_26259);
or U35355 (N_35355,N_26136,N_25540);
and U35356 (N_35356,N_29884,N_24965);
and U35357 (N_35357,N_21570,N_24665);
xnor U35358 (N_35358,N_25720,N_21807);
nand U35359 (N_35359,N_21835,N_29189);
nor U35360 (N_35360,N_20505,N_22904);
nor U35361 (N_35361,N_26501,N_27433);
nand U35362 (N_35362,N_23759,N_25315);
or U35363 (N_35363,N_28905,N_26871);
nor U35364 (N_35364,N_29466,N_20426);
nor U35365 (N_35365,N_29497,N_21145);
xnor U35366 (N_35366,N_29897,N_21761);
nor U35367 (N_35367,N_27253,N_25769);
or U35368 (N_35368,N_21056,N_24095);
nor U35369 (N_35369,N_29342,N_28070);
nand U35370 (N_35370,N_29335,N_20019);
xor U35371 (N_35371,N_21740,N_24406);
nor U35372 (N_35372,N_28618,N_27652);
or U35373 (N_35373,N_25069,N_21090);
and U35374 (N_35374,N_24906,N_23361);
and U35375 (N_35375,N_20875,N_28482);
nand U35376 (N_35376,N_29118,N_27782);
and U35377 (N_35377,N_20634,N_27057);
and U35378 (N_35378,N_24853,N_24429);
nor U35379 (N_35379,N_28466,N_24099);
or U35380 (N_35380,N_29734,N_29429);
nor U35381 (N_35381,N_24465,N_23313);
nor U35382 (N_35382,N_20030,N_25204);
and U35383 (N_35383,N_23462,N_26964);
and U35384 (N_35384,N_22956,N_29397);
or U35385 (N_35385,N_27216,N_26152);
and U35386 (N_35386,N_23721,N_23672);
xnor U35387 (N_35387,N_23112,N_23926);
nand U35388 (N_35388,N_29192,N_21314);
nor U35389 (N_35389,N_25636,N_29314);
and U35390 (N_35390,N_28042,N_28684);
xnor U35391 (N_35391,N_27084,N_25184);
nor U35392 (N_35392,N_29707,N_26743);
and U35393 (N_35393,N_23729,N_22347);
and U35394 (N_35394,N_26264,N_23857);
xnor U35395 (N_35395,N_25039,N_23373);
or U35396 (N_35396,N_24391,N_23897);
nand U35397 (N_35397,N_27695,N_23551);
xor U35398 (N_35398,N_21978,N_26700);
or U35399 (N_35399,N_28530,N_26821);
nand U35400 (N_35400,N_23607,N_29400);
xnor U35401 (N_35401,N_28394,N_29645);
and U35402 (N_35402,N_21116,N_21786);
and U35403 (N_35403,N_27812,N_25665);
and U35404 (N_35404,N_25042,N_23251);
nand U35405 (N_35405,N_24024,N_28389);
or U35406 (N_35406,N_21524,N_27902);
or U35407 (N_35407,N_23886,N_27757);
nor U35408 (N_35408,N_21391,N_28487);
nand U35409 (N_35409,N_28058,N_21045);
and U35410 (N_35410,N_29240,N_29260);
nor U35411 (N_35411,N_21092,N_27927);
nand U35412 (N_35412,N_28127,N_29865);
and U35413 (N_35413,N_20031,N_21241);
or U35414 (N_35414,N_28959,N_29643);
or U35415 (N_35415,N_27172,N_20865);
or U35416 (N_35416,N_25900,N_29227);
or U35417 (N_35417,N_27181,N_20521);
nor U35418 (N_35418,N_25979,N_23248);
nor U35419 (N_35419,N_21521,N_21374);
or U35420 (N_35420,N_26779,N_27323);
nor U35421 (N_35421,N_20644,N_20667);
xor U35422 (N_35422,N_28078,N_23517);
nand U35423 (N_35423,N_20504,N_25384);
xor U35424 (N_35424,N_23217,N_21605);
nand U35425 (N_35425,N_29184,N_22000);
nand U35426 (N_35426,N_27334,N_23125);
or U35427 (N_35427,N_27308,N_28753);
xnor U35428 (N_35428,N_24760,N_20259);
and U35429 (N_35429,N_22728,N_27025);
or U35430 (N_35430,N_25021,N_24849);
nor U35431 (N_35431,N_29997,N_23150);
nand U35432 (N_35432,N_25772,N_23282);
and U35433 (N_35433,N_28862,N_22387);
nand U35434 (N_35434,N_27254,N_22430);
or U35435 (N_35435,N_23304,N_28351);
xnor U35436 (N_35436,N_21616,N_24752);
xnor U35437 (N_35437,N_24648,N_22685);
nor U35438 (N_35438,N_28098,N_21751);
nor U35439 (N_35439,N_27361,N_24548);
nor U35440 (N_35440,N_20452,N_21060);
nand U35441 (N_35441,N_20535,N_22906);
nor U35442 (N_35442,N_24303,N_21742);
nor U35443 (N_35443,N_25527,N_23405);
or U35444 (N_35444,N_28084,N_23618);
or U35445 (N_35445,N_29828,N_28928);
nand U35446 (N_35446,N_26420,N_20805);
and U35447 (N_35447,N_28905,N_25902);
and U35448 (N_35448,N_27577,N_21993);
nor U35449 (N_35449,N_22838,N_24609);
nor U35450 (N_35450,N_21111,N_28337);
nor U35451 (N_35451,N_29863,N_25338);
xor U35452 (N_35452,N_21926,N_25677);
nand U35453 (N_35453,N_24217,N_21521);
xor U35454 (N_35454,N_29863,N_20004);
xnor U35455 (N_35455,N_22432,N_24214);
nor U35456 (N_35456,N_28677,N_23686);
nor U35457 (N_35457,N_23941,N_25323);
xnor U35458 (N_35458,N_21775,N_20370);
xnor U35459 (N_35459,N_29367,N_21604);
or U35460 (N_35460,N_21700,N_25117);
nor U35461 (N_35461,N_26265,N_24068);
nor U35462 (N_35462,N_26191,N_29149);
nor U35463 (N_35463,N_22739,N_29841);
xor U35464 (N_35464,N_26447,N_27261);
nor U35465 (N_35465,N_29135,N_29669);
xor U35466 (N_35466,N_28821,N_28780);
nand U35467 (N_35467,N_23140,N_23942);
and U35468 (N_35468,N_27013,N_22760);
or U35469 (N_35469,N_21927,N_23359);
xor U35470 (N_35470,N_20426,N_23686);
and U35471 (N_35471,N_21858,N_24027);
xnor U35472 (N_35472,N_24618,N_27209);
xor U35473 (N_35473,N_26769,N_25166);
xnor U35474 (N_35474,N_22819,N_22735);
nor U35475 (N_35475,N_23779,N_29632);
or U35476 (N_35476,N_22873,N_25449);
nor U35477 (N_35477,N_28160,N_21017);
xnor U35478 (N_35478,N_29566,N_27109);
nor U35479 (N_35479,N_27051,N_20743);
nand U35480 (N_35480,N_24820,N_28914);
nor U35481 (N_35481,N_27445,N_28722);
xnor U35482 (N_35482,N_25934,N_24358);
or U35483 (N_35483,N_27809,N_22439);
nand U35484 (N_35484,N_26604,N_27523);
or U35485 (N_35485,N_24011,N_27664);
nand U35486 (N_35486,N_23069,N_21158);
or U35487 (N_35487,N_23260,N_23846);
and U35488 (N_35488,N_24793,N_28112);
xnor U35489 (N_35489,N_24539,N_23557);
and U35490 (N_35490,N_24186,N_25108);
or U35491 (N_35491,N_20848,N_20944);
and U35492 (N_35492,N_25423,N_27920);
nor U35493 (N_35493,N_23834,N_22582);
nand U35494 (N_35494,N_26453,N_25869);
nand U35495 (N_35495,N_20840,N_24908);
xnor U35496 (N_35496,N_20904,N_20108);
and U35497 (N_35497,N_20075,N_28494);
nor U35498 (N_35498,N_24267,N_27669);
and U35499 (N_35499,N_24693,N_21692);
and U35500 (N_35500,N_26631,N_21499);
nand U35501 (N_35501,N_22017,N_22127);
nand U35502 (N_35502,N_25783,N_27771);
nor U35503 (N_35503,N_26473,N_23442);
xor U35504 (N_35504,N_29063,N_22381);
nand U35505 (N_35505,N_22422,N_25686);
xnor U35506 (N_35506,N_27173,N_21357);
or U35507 (N_35507,N_25692,N_24803);
xnor U35508 (N_35508,N_21822,N_26574);
nand U35509 (N_35509,N_28018,N_20790);
and U35510 (N_35510,N_22771,N_27505);
and U35511 (N_35511,N_26919,N_24241);
nand U35512 (N_35512,N_28474,N_28765);
xnor U35513 (N_35513,N_29221,N_27658);
and U35514 (N_35514,N_21977,N_25878);
nor U35515 (N_35515,N_28399,N_29152);
and U35516 (N_35516,N_29414,N_27645);
and U35517 (N_35517,N_24479,N_24804);
nor U35518 (N_35518,N_20296,N_21134);
or U35519 (N_35519,N_23180,N_24321);
xor U35520 (N_35520,N_27589,N_25232);
and U35521 (N_35521,N_28678,N_20273);
and U35522 (N_35522,N_25618,N_27810);
xor U35523 (N_35523,N_21414,N_28576);
and U35524 (N_35524,N_25369,N_28289);
xor U35525 (N_35525,N_21715,N_28772);
nor U35526 (N_35526,N_29157,N_28529);
or U35527 (N_35527,N_24825,N_20457);
or U35528 (N_35528,N_29220,N_25142);
and U35529 (N_35529,N_25947,N_27978);
nor U35530 (N_35530,N_21496,N_23027);
xnor U35531 (N_35531,N_26457,N_22563);
and U35532 (N_35532,N_20531,N_25522);
nor U35533 (N_35533,N_28744,N_28153);
nor U35534 (N_35534,N_23775,N_23654);
nand U35535 (N_35535,N_24569,N_21560);
nor U35536 (N_35536,N_25643,N_23738);
nand U35537 (N_35537,N_27956,N_23890);
nand U35538 (N_35538,N_20642,N_23446);
nor U35539 (N_35539,N_29495,N_22875);
and U35540 (N_35540,N_24709,N_26428);
xor U35541 (N_35541,N_23233,N_26413);
xnor U35542 (N_35542,N_29119,N_28827);
nor U35543 (N_35543,N_22409,N_28794);
or U35544 (N_35544,N_26614,N_26863);
xor U35545 (N_35545,N_23727,N_21201);
nor U35546 (N_35546,N_21775,N_25828);
xor U35547 (N_35547,N_28648,N_28295);
xnor U35548 (N_35548,N_25222,N_23449);
xor U35549 (N_35549,N_27610,N_20709);
nor U35550 (N_35550,N_23372,N_22793);
nand U35551 (N_35551,N_26872,N_22844);
or U35552 (N_35552,N_21839,N_27466);
nand U35553 (N_35553,N_28111,N_20125);
or U35554 (N_35554,N_21309,N_28425);
nor U35555 (N_35555,N_23203,N_21570);
nand U35556 (N_35556,N_25336,N_25391);
nor U35557 (N_35557,N_24672,N_22878);
nand U35558 (N_35558,N_24475,N_29141);
nand U35559 (N_35559,N_20262,N_22147);
and U35560 (N_35560,N_20860,N_20413);
and U35561 (N_35561,N_27222,N_24984);
nand U35562 (N_35562,N_25547,N_22167);
xor U35563 (N_35563,N_21744,N_21871);
nor U35564 (N_35564,N_24333,N_26607);
xnor U35565 (N_35565,N_26887,N_20498);
nand U35566 (N_35566,N_22141,N_27019);
and U35567 (N_35567,N_27080,N_25327);
and U35568 (N_35568,N_23852,N_24499);
and U35569 (N_35569,N_22345,N_24044);
nor U35570 (N_35570,N_27711,N_22584);
nand U35571 (N_35571,N_20902,N_20778);
xnor U35572 (N_35572,N_24302,N_24960);
or U35573 (N_35573,N_28292,N_24634);
nand U35574 (N_35574,N_25231,N_26147);
xor U35575 (N_35575,N_20672,N_25384);
xnor U35576 (N_35576,N_29415,N_26325);
and U35577 (N_35577,N_28636,N_20414);
nand U35578 (N_35578,N_23446,N_23171);
nand U35579 (N_35579,N_29829,N_29709);
nand U35580 (N_35580,N_23362,N_29056);
nand U35581 (N_35581,N_21309,N_29915);
and U35582 (N_35582,N_27925,N_23812);
xor U35583 (N_35583,N_26225,N_29817);
xor U35584 (N_35584,N_25278,N_20234);
and U35585 (N_35585,N_29809,N_24447);
and U35586 (N_35586,N_22420,N_24170);
xor U35587 (N_35587,N_24145,N_20493);
and U35588 (N_35588,N_26169,N_22504);
and U35589 (N_35589,N_22275,N_22447);
xor U35590 (N_35590,N_24569,N_20017);
nor U35591 (N_35591,N_21478,N_25993);
or U35592 (N_35592,N_28934,N_20303);
nand U35593 (N_35593,N_20242,N_25604);
xor U35594 (N_35594,N_20805,N_28818);
or U35595 (N_35595,N_25094,N_29589);
xnor U35596 (N_35596,N_20115,N_24668);
nor U35597 (N_35597,N_23369,N_24048);
nor U35598 (N_35598,N_24083,N_22443);
and U35599 (N_35599,N_27122,N_24433);
or U35600 (N_35600,N_29154,N_21116);
nand U35601 (N_35601,N_26303,N_28805);
and U35602 (N_35602,N_27332,N_26725);
and U35603 (N_35603,N_24390,N_23895);
nor U35604 (N_35604,N_20340,N_24251);
or U35605 (N_35605,N_24037,N_20024);
xnor U35606 (N_35606,N_21587,N_20023);
nand U35607 (N_35607,N_25169,N_23295);
nor U35608 (N_35608,N_23811,N_24897);
xor U35609 (N_35609,N_29217,N_26965);
and U35610 (N_35610,N_24998,N_27509);
and U35611 (N_35611,N_20785,N_22726);
xor U35612 (N_35612,N_28098,N_21818);
nand U35613 (N_35613,N_24758,N_23326);
and U35614 (N_35614,N_21254,N_25911);
nor U35615 (N_35615,N_27375,N_28792);
and U35616 (N_35616,N_25171,N_23409);
nor U35617 (N_35617,N_29898,N_29805);
nor U35618 (N_35618,N_20456,N_21379);
xnor U35619 (N_35619,N_28274,N_29509);
xor U35620 (N_35620,N_26646,N_24703);
nand U35621 (N_35621,N_28150,N_27920);
and U35622 (N_35622,N_26582,N_20882);
nand U35623 (N_35623,N_28944,N_28501);
or U35624 (N_35624,N_24146,N_20794);
nand U35625 (N_35625,N_22137,N_23485);
nand U35626 (N_35626,N_21229,N_23768);
xnor U35627 (N_35627,N_27172,N_27569);
nor U35628 (N_35628,N_26908,N_21313);
or U35629 (N_35629,N_20759,N_23237);
nand U35630 (N_35630,N_28202,N_26596);
xor U35631 (N_35631,N_27411,N_22887);
nand U35632 (N_35632,N_21024,N_27773);
xor U35633 (N_35633,N_20924,N_28287);
or U35634 (N_35634,N_26061,N_28501);
xnor U35635 (N_35635,N_24573,N_25586);
xor U35636 (N_35636,N_29094,N_23423);
nand U35637 (N_35637,N_26028,N_29358);
and U35638 (N_35638,N_27987,N_22864);
nor U35639 (N_35639,N_20941,N_23315);
xnor U35640 (N_35640,N_28907,N_23541);
nand U35641 (N_35641,N_27684,N_27809);
and U35642 (N_35642,N_25363,N_27694);
or U35643 (N_35643,N_23804,N_27200);
or U35644 (N_35644,N_22197,N_22516);
xnor U35645 (N_35645,N_24410,N_21542);
nor U35646 (N_35646,N_23615,N_22125);
nor U35647 (N_35647,N_25091,N_26048);
nor U35648 (N_35648,N_28080,N_20602);
or U35649 (N_35649,N_28074,N_25754);
xnor U35650 (N_35650,N_21483,N_28992);
or U35651 (N_35651,N_21023,N_22921);
or U35652 (N_35652,N_28341,N_27068);
nor U35653 (N_35653,N_23723,N_23198);
nand U35654 (N_35654,N_22656,N_20519);
nand U35655 (N_35655,N_25900,N_28411);
xnor U35656 (N_35656,N_21165,N_21053);
or U35657 (N_35657,N_28573,N_26964);
nand U35658 (N_35658,N_27725,N_24194);
and U35659 (N_35659,N_28915,N_22741);
xnor U35660 (N_35660,N_22628,N_23686);
or U35661 (N_35661,N_21726,N_24888);
and U35662 (N_35662,N_20960,N_24507);
xnor U35663 (N_35663,N_24285,N_26761);
nand U35664 (N_35664,N_21083,N_20083);
nor U35665 (N_35665,N_24437,N_21736);
and U35666 (N_35666,N_29178,N_27417);
xor U35667 (N_35667,N_21297,N_29933);
nand U35668 (N_35668,N_23660,N_26584);
xor U35669 (N_35669,N_20257,N_29310);
nand U35670 (N_35670,N_27516,N_25101);
or U35671 (N_35671,N_23699,N_20372);
xnor U35672 (N_35672,N_27306,N_24233);
nand U35673 (N_35673,N_24861,N_25262);
nand U35674 (N_35674,N_20815,N_20535);
nor U35675 (N_35675,N_26013,N_21894);
xor U35676 (N_35676,N_24167,N_29644);
nand U35677 (N_35677,N_21498,N_22815);
xor U35678 (N_35678,N_27280,N_20231);
xnor U35679 (N_35679,N_24980,N_20784);
xnor U35680 (N_35680,N_21249,N_21778);
or U35681 (N_35681,N_24718,N_26301);
or U35682 (N_35682,N_28651,N_24304);
nand U35683 (N_35683,N_22261,N_26092);
or U35684 (N_35684,N_26605,N_22370);
nor U35685 (N_35685,N_22279,N_23456);
and U35686 (N_35686,N_28547,N_24610);
nand U35687 (N_35687,N_20536,N_24191);
xnor U35688 (N_35688,N_26489,N_24977);
xnor U35689 (N_35689,N_25382,N_29726);
xnor U35690 (N_35690,N_29297,N_27154);
nand U35691 (N_35691,N_28303,N_21395);
nand U35692 (N_35692,N_27559,N_23928);
or U35693 (N_35693,N_28291,N_22757);
xor U35694 (N_35694,N_27585,N_25314);
or U35695 (N_35695,N_22551,N_24748);
nand U35696 (N_35696,N_26905,N_21492);
or U35697 (N_35697,N_29764,N_25480);
nand U35698 (N_35698,N_24738,N_25763);
or U35699 (N_35699,N_28597,N_23798);
nand U35700 (N_35700,N_22100,N_22537);
or U35701 (N_35701,N_27741,N_29033);
nand U35702 (N_35702,N_27165,N_22022);
nor U35703 (N_35703,N_29504,N_24768);
and U35704 (N_35704,N_29291,N_21183);
nor U35705 (N_35705,N_23431,N_26687);
and U35706 (N_35706,N_22020,N_20524);
and U35707 (N_35707,N_23450,N_23242);
or U35708 (N_35708,N_24269,N_20792);
or U35709 (N_35709,N_22649,N_21736);
or U35710 (N_35710,N_22665,N_20922);
xnor U35711 (N_35711,N_23716,N_26006);
xor U35712 (N_35712,N_21634,N_25798);
nor U35713 (N_35713,N_24168,N_22889);
nand U35714 (N_35714,N_20532,N_28093);
and U35715 (N_35715,N_25384,N_21717);
nor U35716 (N_35716,N_23063,N_20314);
nor U35717 (N_35717,N_24056,N_27601);
nor U35718 (N_35718,N_27298,N_26804);
nor U35719 (N_35719,N_25969,N_23576);
xor U35720 (N_35720,N_23644,N_22969);
and U35721 (N_35721,N_29254,N_24335);
nand U35722 (N_35722,N_26989,N_22042);
xnor U35723 (N_35723,N_29719,N_22834);
nand U35724 (N_35724,N_24320,N_23939);
nor U35725 (N_35725,N_28050,N_24971);
xor U35726 (N_35726,N_23245,N_27467);
nand U35727 (N_35727,N_23676,N_28515);
and U35728 (N_35728,N_20904,N_23799);
xor U35729 (N_35729,N_25003,N_28460);
xnor U35730 (N_35730,N_29299,N_25177);
nor U35731 (N_35731,N_28602,N_22523);
or U35732 (N_35732,N_29369,N_26860);
and U35733 (N_35733,N_23758,N_21409);
or U35734 (N_35734,N_25653,N_27012);
nor U35735 (N_35735,N_26754,N_22437);
nor U35736 (N_35736,N_28399,N_28069);
and U35737 (N_35737,N_24700,N_27226);
xor U35738 (N_35738,N_21754,N_24619);
and U35739 (N_35739,N_21517,N_25751);
or U35740 (N_35740,N_26921,N_25485);
nor U35741 (N_35741,N_22729,N_22619);
nand U35742 (N_35742,N_20674,N_25969);
nor U35743 (N_35743,N_21450,N_25735);
xor U35744 (N_35744,N_20256,N_29480);
nor U35745 (N_35745,N_23514,N_29835);
and U35746 (N_35746,N_22044,N_26367);
and U35747 (N_35747,N_21142,N_29720);
nor U35748 (N_35748,N_25093,N_26761);
or U35749 (N_35749,N_26879,N_24211);
or U35750 (N_35750,N_29487,N_20353);
or U35751 (N_35751,N_27863,N_22026);
nor U35752 (N_35752,N_28715,N_28263);
and U35753 (N_35753,N_22925,N_24550);
and U35754 (N_35754,N_27037,N_28290);
nor U35755 (N_35755,N_26140,N_20051);
nand U35756 (N_35756,N_20793,N_29062);
nor U35757 (N_35757,N_28954,N_27300);
xnor U35758 (N_35758,N_25059,N_21099);
or U35759 (N_35759,N_28701,N_28442);
and U35760 (N_35760,N_21527,N_24018);
nor U35761 (N_35761,N_28866,N_21869);
xor U35762 (N_35762,N_21710,N_28092);
nor U35763 (N_35763,N_27687,N_26862);
nor U35764 (N_35764,N_29728,N_28147);
and U35765 (N_35765,N_26269,N_20862);
and U35766 (N_35766,N_20819,N_20379);
nand U35767 (N_35767,N_25402,N_29005);
or U35768 (N_35768,N_26192,N_27404);
or U35769 (N_35769,N_27299,N_23097);
nand U35770 (N_35770,N_20903,N_26913);
nor U35771 (N_35771,N_22092,N_22393);
nor U35772 (N_35772,N_23250,N_27327);
or U35773 (N_35773,N_23303,N_25660);
nand U35774 (N_35774,N_26840,N_29455);
nor U35775 (N_35775,N_21014,N_29140);
nand U35776 (N_35776,N_23628,N_25839);
or U35777 (N_35777,N_21003,N_28439);
and U35778 (N_35778,N_21183,N_28712);
nor U35779 (N_35779,N_22762,N_20968);
nand U35780 (N_35780,N_23242,N_21363);
nor U35781 (N_35781,N_29466,N_23901);
and U35782 (N_35782,N_26557,N_24488);
and U35783 (N_35783,N_22350,N_24908);
nor U35784 (N_35784,N_26692,N_23983);
xnor U35785 (N_35785,N_22824,N_29253);
nor U35786 (N_35786,N_26284,N_22208);
xnor U35787 (N_35787,N_23980,N_26184);
and U35788 (N_35788,N_23553,N_22261);
or U35789 (N_35789,N_23655,N_28626);
nand U35790 (N_35790,N_28585,N_27411);
nor U35791 (N_35791,N_25138,N_24141);
and U35792 (N_35792,N_20310,N_23966);
xor U35793 (N_35793,N_21593,N_24364);
nand U35794 (N_35794,N_21229,N_25116);
xor U35795 (N_35795,N_20490,N_22624);
and U35796 (N_35796,N_28685,N_28484);
xnor U35797 (N_35797,N_28857,N_29892);
and U35798 (N_35798,N_24636,N_24562);
xor U35799 (N_35799,N_27252,N_23438);
or U35800 (N_35800,N_20117,N_25150);
nand U35801 (N_35801,N_24879,N_26666);
nor U35802 (N_35802,N_26379,N_26852);
nor U35803 (N_35803,N_24342,N_28003);
nor U35804 (N_35804,N_29376,N_26324);
or U35805 (N_35805,N_24346,N_20809);
and U35806 (N_35806,N_24546,N_26265);
xnor U35807 (N_35807,N_20270,N_24387);
or U35808 (N_35808,N_22421,N_21168);
xnor U35809 (N_35809,N_24667,N_22092);
and U35810 (N_35810,N_28304,N_29948);
nand U35811 (N_35811,N_26446,N_26611);
nand U35812 (N_35812,N_23112,N_25129);
xnor U35813 (N_35813,N_23350,N_27953);
xnor U35814 (N_35814,N_24953,N_28923);
nand U35815 (N_35815,N_25415,N_26902);
and U35816 (N_35816,N_21583,N_29929);
xor U35817 (N_35817,N_29891,N_27476);
and U35818 (N_35818,N_24226,N_22567);
nand U35819 (N_35819,N_23047,N_20365);
nand U35820 (N_35820,N_26019,N_23828);
nand U35821 (N_35821,N_28573,N_25824);
nor U35822 (N_35822,N_29197,N_21881);
nand U35823 (N_35823,N_27546,N_25120);
nor U35824 (N_35824,N_27251,N_20776);
or U35825 (N_35825,N_27852,N_29647);
or U35826 (N_35826,N_21424,N_25593);
or U35827 (N_35827,N_28693,N_21816);
or U35828 (N_35828,N_24136,N_22074);
and U35829 (N_35829,N_20798,N_23759);
xnor U35830 (N_35830,N_23152,N_25532);
nor U35831 (N_35831,N_28384,N_29033);
nand U35832 (N_35832,N_20403,N_21403);
and U35833 (N_35833,N_28750,N_25877);
xor U35834 (N_35834,N_20214,N_26658);
or U35835 (N_35835,N_26799,N_20619);
and U35836 (N_35836,N_27130,N_24710);
and U35837 (N_35837,N_29297,N_20489);
xnor U35838 (N_35838,N_24442,N_29666);
xor U35839 (N_35839,N_20529,N_23775);
or U35840 (N_35840,N_26714,N_25220);
nand U35841 (N_35841,N_26592,N_29485);
or U35842 (N_35842,N_20919,N_25941);
and U35843 (N_35843,N_21954,N_27559);
nor U35844 (N_35844,N_24174,N_26261);
or U35845 (N_35845,N_26308,N_26355);
and U35846 (N_35846,N_23964,N_24658);
nand U35847 (N_35847,N_25345,N_24002);
or U35848 (N_35848,N_21479,N_28009);
nor U35849 (N_35849,N_26137,N_26150);
or U35850 (N_35850,N_26790,N_29611);
and U35851 (N_35851,N_27027,N_23755);
nor U35852 (N_35852,N_25356,N_22123);
nor U35853 (N_35853,N_21251,N_23864);
xnor U35854 (N_35854,N_22643,N_24963);
and U35855 (N_35855,N_26116,N_24378);
and U35856 (N_35856,N_24894,N_25955);
nand U35857 (N_35857,N_20012,N_27926);
nand U35858 (N_35858,N_26994,N_27307);
or U35859 (N_35859,N_28295,N_25863);
and U35860 (N_35860,N_23413,N_22047);
nand U35861 (N_35861,N_23765,N_26896);
and U35862 (N_35862,N_26901,N_23283);
nor U35863 (N_35863,N_26697,N_29394);
or U35864 (N_35864,N_29891,N_22004);
nand U35865 (N_35865,N_22731,N_23575);
xnor U35866 (N_35866,N_21645,N_27968);
xor U35867 (N_35867,N_29381,N_21180);
xnor U35868 (N_35868,N_27763,N_20759);
or U35869 (N_35869,N_20794,N_25471);
and U35870 (N_35870,N_23012,N_25871);
or U35871 (N_35871,N_25875,N_20924);
and U35872 (N_35872,N_23850,N_21904);
nor U35873 (N_35873,N_26091,N_23235);
nand U35874 (N_35874,N_22525,N_23568);
xnor U35875 (N_35875,N_29548,N_21081);
or U35876 (N_35876,N_20927,N_22134);
nor U35877 (N_35877,N_21481,N_28533);
and U35878 (N_35878,N_24179,N_27151);
nor U35879 (N_35879,N_28382,N_29910);
nand U35880 (N_35880,N_29214,N_24832);
nand U35881 (N_35881,N_29456,N_26221);
nand U35882 (N_35882,N_20953,N_29461);
nor U35883 (N_35883,N_26743,N_27752);
xnor U35884 (N_35884,N_20604,N_29656);
nand U35885 (N_35885,N_28238,N_21084);
and U35886 (N_35886,N_21224,N_22105);
nor U35887 (N_35887,N_21726,N_20687);
or U35888 (N_35888,N_29627,N_20502);
xor U35889 (N_35889,N_27181,N_26907);
or U35890 (N_35890,N_20547,N_27018);
and U35891 (N_35891,N_22565,N_26981);
and U35892 (N_35892,N_22874,N_22488);
nor U35893 (N_35893,N_27430,N_27532);
xor U35894 (N_35894,N_22271,N_23890);
and U35895 (N_35895,N_29253,N_29931);
and U35896 (N_35896,N_24997,N_26845);
nand U35897 (N_35897,N_29620,N_28249);
xnor U35898 (N_35898,N_26590,N_22623);
nor U35899 (N_35899,N_21022,N_23872);
nor U35900 (N_35900,N_25165,N_23308);
nor U35901 (N_35901,N_23245,N_26564);
nand U35902 (N_35902,N_27117,N_25769);
and U35903 (N_35903,N_25970,N_23630);
or U35904 (N_35904,N_21978,N_24504);
and U35905 (N_35905,N_20164,N_23397);
nor U35906 (N_35906,N_24952,N_25460);
nand U35907 (N_35907,N_23659,N_29822);
or U35908 (N_35908,N_21988,N_20105);
xor U35909 (N_35909,N_27609,N_29805);
nor U35910 (N_35910,N_21916,N_28987);
or U35911 (N_35911,N_21759,N_26343);
and U35912 (N_35912,N_27016,N_20360);
or U35913 (N_35913,N_27816,N_24365);
or U35914 (N_35914,N_28169,N_25467);
nand U35915 (N_35915,N_29537,N_25577);
and U35916 (N_35916,N_22420,N_26742);
nor U35917 (N_35917,N_28143,N_23211);
and U35918 (N_35918,N_20030,N_29278);
nor U35919 (N_35919,N_25741,N_27833);
and U35920 (N_35920,N_25620,N_23488);
or U35921 (N_35921,N_29325,N_20266);
or U35922 (N_35922,N_20101,N_22659);
nor U35923 (N_35923,N_24772,N_22204);
and U35924 (N_35924,N_20810,N_25698);
xnor U35925 (N_35925,N_23720,N_29110);
nor U35926 (N_35926,N_22349,N_21203);
nor U35927 (N_35927,N_28963,N_23430);
nor U35928 (N_35928,N_28852,N_29497);
or U35929 (N_35929,N_26683,N_28638);
xor U35930 (N_35930,N_28667,N_26402);
or U35931 (N_35931,N_29914,N_29143);
nor U35932 (N_35932,N_24148,N_29175);
or U35933 (N_35933,N_27619,N_20197);
xor U35934 (N_35934,N_20304,N_28121);
and U35935 (N_35935,N_20746,N_21622);
or U35936 (N_35936,N_21068,N_25006);
or U35937 (N_35937,N_24971,N_27873);
and U35938 (N_35938,N_20464,N_24965);
nand U35939 (N_35939,N_27658,N_27663);
and U35940 (N_35940,N_22030,N_22635);
nand U35941 (N_35941,N_22081,N_22514);
and U35942 (N_35942,N_25443,N_25588);
or U35943 (N_35943,N_21847,N_24160);
xor U35944 (N_35944,N_26699,N_21418);
and U35945 (N_35945,N_25063,N_21000);
or U35946 (N_35946,N_28384,N_29869);
nor U35947 (N_35947,N_24790,N_26470);
xnor U35948 (N_35948,N_23193,N_22130);
and U35949 (N_35949,N_24864,N_20854);
and U35950 (N_35950,N_20895,N_25926);
nand U35951 (N_35951,N_25627,N_26693);
xnor U35952 (N_35952,N_29408,N_27634);
and U35953 (N_35953,N_28715,N_21782);
or U35954 (N_35954,N_21457,N_25635);
xnor U35955 (N_35955,N_23809,N_23216);
nand U35956 (N_35956,N_29980,N_27197);
or U35957 (N_35957,N_24026,N_28681);
xnor U35958 (N_35958,N_25637,N_29028);
xor U35959 (N_35959,N_21603,N_22614);
and U35960 (N_35960,N_26644,N_21028);
nand U35961 (N_35961,N_22888,N_20357);
or U35962 (N_35962,N_27682,N_22095);
nor U35963 (N_35963,N_28039,N_22724);
and U35964 (N_35964,N_20059,N_20368);
nor U35965 (N_35965,N_28451,N_21845);
nand U35966 (N_35966,N_22566,N_27521);
and U35967 (N_35967,N_29472,N_22774);
nand U35968 (N_35968,N_24754,N_27066);
xnor U35969 (N_35969,N_28990,N_20129);
nand U35970 (N_35970,N_28506,N_24018);
nand U35971 (N_35971,N_25977,N_26221);
nand U35972 (N_35972,N_29276,N_27515);
xor U35973 (N_35973,N_20009,N_25251);
or U35974 (N_35974,N_24278,N_21217);
and U35975 (N_35975,N_27467,N_21948);
and U35976 (N_35976,N_25157,N_25115);
xor U35977 (N_35977,N_24461,N_21898);
xnor U35978 (N_35978,N_26528,N_26754);
nor U35979 (N_35979,N_20083,N_27357);
and U35980 (N_35980,N_23266,N_27361);
or U35981 (N_35981,N_22679,N_26327);
and U35982 (N_35982,N_29767,N_26938);
and U35983 (N_35983,N_25119,N_24829);
and U35984 (N_35984,N_24424,N_25682);
or U35985 (N_35985,N_25861,N_27911);
nand U35986 (N_35986,N_21543,N_27826);
nor U35987 (N_35987,N_28233,N_28525);
and U35988 (N_35988,N_21522,N_24479);
and U35989 (N_35989,N_26304,N_27495);
nand U35990 (N_35990,N_29989,N_20343);
nor U35991 (N_35991,N_22426,N_20865);
nand U35992 (N_35992,N_27210,N_26590);
or U35993 (N_35993,N_27311,N_20586);
and U35994 (N_35994,N_28348,N_23892);
nand U35995 (N_35995,N_27267,N_28214);
nand U35996 (N_35996,N_28645,N_21481);
or U35997 (N_35997,N_26201,N_26265);
or U35998 (N_35998,N_29827,N_20803);
and U35999 (N_35999,N_21950,N_27562);
nor U36000 (N_36000,N_21093,N_20812);
nand U36001 (N_36001,N_27327,N_23625);
nor U36002 (N_36002,N_25868,N_21331);
xnor U36003 (N_36003,N_24138,N_27121);
nand U36004 (N_36004,N_23767,N_21500);
xnor U36005 (N_36005,N_26551,N_21855);
nor U36006 (N_36006,N_21992,N_23680);
xnor U36007 (N_36007,N_23549,N_20593);
nor U36008 (N_36008,N_20516,N_28288);
or U36009 (N_36009,N_25164,N_29186);
nand U36010 (N_36010,N_22745,N_22695);
nor U36011 (N_36011,N_25083,N_22045);
or U36012 (N_36012,N_23793,N_27876);
nand U36013 (N_36013,N_22088,N_27308);
nand U36014 (N_36014,N_20088,N_28489);
nand U36015 (N_36015,N_29014,N_22957);
and U36016 (N_36016,N_23222,N_24735);
nor U36017 (N_36017,N_22388,N_26442);
nor U36018 (N_36018,N_24030,N_23963);
xor U36019 (N_36019,N_23934,N_24145);
and U36020 (N_36020,N_26893,N_23280);
xnor U36021 (N_36021,N_22447,N_23529);
nor U36022 (N_36022,N_20804,N_20506);
nand U36023 (N_36023,N_20007,N_28414);
nor U36024 (N_36024,N_28797,N_26457);
nand U36025 (N_36025,N_24532,N_28203);
nor U36026 (N_36026,N_22106,N_27942);
nand U36027 (N_36027,N_27120,N_25841);
nor U36028 (N_36028,N_29301,N_26066);
nand U36029 (N_36029,N_20053,N_28411);
nand U36030 (N_36030,N_27300,N_24672);
and U36031 (N_36031,N_26931,N_27996);
xnor U36032 (N_36032,N_28808,N_23238);
nand U36033 (N_36033,N_20521,N_20078);
xor U36034 (N_36034,N_22387,N_20228);
or U36035 (N_36035,N_21153,N_21919);
nor U36036 (N_36036,N_23423,N_27472);
xnor U36037 (N_36037,N_28214,N_23399);
nor U36038 (N_36038,N_28001,N_22971);
xor U36039 (N_36039,N_28385,N_24442);
and U36040 (N_36040,N_29503,N_21444);
nand U36041 (N_36041,N_26840,N_26553);
nand U36042 (N_36042,N_24988,N_27692);
and U36043 (N_36043,N_26551,N_21150);
nor U36044 (N_36044,N_26872,N_20066);
nor U36045 (N_36045,N_26228,N_29774);
xor U36046 (N_36046,N_23710,N_24661);
nor U36047 (N_36047,N_25069,N_29231);
xor U36048 (N_36048,N_29494,N_25108);
xor U36049 (N_36049,N_26925,N_23134);
and U36050 (N_36050,N_28426,N_29508);
nor U36051 (N_36051,N_26577,N_22799);
nand U36052 (N_36052,N_29425,N_29719);
nand U36053 (N_36053,N_28867,N_22262);
xnor U36054 (N_36054,N_28886,N_22157);
xor U36055 (N_36055,N_22915,N_21747);
nor U36056 (N_36056,N_26828,N_22538);
and U36057 (N_36057,N_26968,N_26640);
or U36058 (N_36058,N_25559,N_24428);
or U36059 (N_36059,N_28836,N_23164);
xnor U36060 (N_36060,N_20288,N_21106);
or U36061 (N_36061,N_20672,N_20281);
xor U36062 (N_36062,N_23591,N_28498);
xnor U36063 (N_36063,N_21108,N_27835);
nand U36064 (N_36064,N_24718,N_25489);
or U36065 (N_36065,N_22900,N_24533);
or U36066 (N_36066,N_22527,N_29507);
xor U36067 (N_36067,N_21013,N_26844);
nand U36068 (N_36068,N_22833,N_22767);
nor U36069 (N_36069,N_20942,N_27454);
and U36070 (N_36070,N_21783,N_26991);
xor U36071 (N_36071,N_21575,N_29921);
xor U36072 (N_36072,N_27850,N_24203);
or U36073 (N_36073,N_26181,N_27121);
and U36074 (N_36074,N_25624,N_23378);
xor U36075 (N_36075,N_24895,N_24022);
xnor U36076 (N_36076,N_24010,N_24540);
xnor U36077 (N_36077,N_29571,N_29374);
nand U36078 (N_36078,N_25714,N_25379);
or U36079 (N_36079,N_28952,N_22737);
nand U36080 (N_36080,N_25620,N_29092);
xor U36081 (N_36081,N_21126,N_23676);
nor U36082 (N_36082,N_29543,N_28193);
or U36083 (N_36083,N_29381,N_21923);
nor U36084 (N_36084,N_27049,N_25746);
or U36085 (N_36085,N_25931,N_26110);
or U36086 (N_36086,N_21303,N_21106);
or U36087 (N_36087,N_21661,N_24264);
xnor U36088 (N_36088,N_25572,N_22325);
and U36089 (N_36089,N_26234,N_21107);
or U36090 (N_36090,N_29165,N_28677);
and U36091 (N_36091,N_26916,N_26794);
xnor U36092 (N_36092,N_25010,N_23874);
and U36093 (N_36093,N_24103,N_29555);
xor U36094 (N_36094,N_20218,N_29075);
nand U36095 (N_36095,N_24562,N_24227);
nor U36096 (N_36096,N_28100,N_27775);
nand U36097 (N_36097,N_29872,N_23143);
nand U36098 (N_36098,N_25025,N_27727);
and U36099 (N_36099,N_27228,N_22765);
nor U36100 (N_36100,N_28817,N_25718);
nor U36101 (N_36101,N_21381,N_21423);
nand U36102 (N_36102,N_25248,N_28012);
xor U36103 (N_36103,N_27072,N_21570);
nand U36104 (N_36104,N_25355,N_27694);
nor U36105 (N_36105,N_20687,N_26501);
and U36106 (N_36106,N_23481,N_27492);
or U36107 (N_36107,N_29308,N_25204);
and U36108 (N_36108,N_26775,N_23486);
nor U36109 (N_36109,N_22871,N_26675);
or U36110 (N_36110,N_26788,N_26767);
nand U36111 (N_36111,N_21083,N_29164);
or U36112 (N_36112,N_26929,N_23058);
and U36113 (N_36113,N_24197,N_26629);
nand U36114 (N_36114,N_20522,N_21794);
and U36115 (N_36115,N_24111,N_23223);
nand U36116 (N_36116,N_23670,N_28071);
xor U36117 (N_36117,N_26212,N_24238);
and U36118 (N_36118,N_28391,N_28628);
nand U36119 (N_36119,N_25621,N_29757);
nand U36120 (N_36120,N_20112,N_29564);
xnor U36121 (N_36121,N_22182,N_24685);
or U36122 (N_36122,N_23943,N_25722);
xnor U36123 (N_36123,N_28743,N_22789);
nor U36124 (N_36124,N_25457,N_25594);
nand U36125 (N_36125,N_24538,N_29387);
nor U36126 (N_36126,N_20626,N_22321);
and U36127 (N_36127,N_28884,N_25358);
nand U36128 (N_36128,N_20080,N_21066);
nand U36129 (N_36129,N_29121,N_22159);
and U36130 (N_36130,N_20270,N_24235);
xnor U36131 (N_36131,N_27975,N_22604);
xor U36132 (N_36132,N_26814,N_22171);
or U36133 (N_36133,N_27607,N_28719);
or U36134 (N_36134,N_21639,N_20958);
or U36135 (N_36135,N_22686,N_27445);
nand U36136 (N_36136,N_27855,N_21105);
nand U36137 (N_36137,N_29171,N_28089);
xor U36138 (N_36138,N_26650,N_21515);
nand U36139 (N_36139,N_29162,N_26816);
nor U36140 (N_36140,N_25552,N_26106);
xnor U36141 (N_36141,N_20081,N_27484);
and U36142 (N_36142,N_21831,N_20921);
nor U36143 (N_36143,N_20321,N_21981);
and U36144 (N_36144,N_28027,N_25349);
nor U36145 (N_36145,N_22140,N_23491);
nand U36146 (N_36146,N_29978,N_28773);
nand U36147 (N_36147,N_29571,N_29304);
nand U36148 (N_36148,N_22337,N_27859);
xor U36149 (N_36149,N_22934,N_28731);
and U36150 (N_36150,N_21388,N_20971);
nor U36151 (N_36151,N_29904,N_28337);
and U36152 (N_36152,N_25345,N_29845);
xnor U36153 (N_36153,N_24375,N_29419);
nand U36154 (N_36154,N_27926,N_21023);
or U36155 (N_36155,N_29867,N_28905);
or U36156 (N_36156,N_23979,N_21580);
nor U36157 (N_36157,N_29016,N_25669);
nand U36158 (N_36158,N_27499,N_26979);
or U36159 (N_36159,N_25014,N_21192);
and U36160 (N_36160,N_25498,N_21924);
and U36161 (N_36161,N_23001,N_29931);
xor U36162 (N_36162,N_29243,N_23483);
xor U36163 (N_36163,N_21490,N_23875);
or U36164 (N_36164,N_27503,N_21402);
and U36165 (N_36165,N_20766,N_20574);
nand U36166 (N_36166,N_22095,N_24167);
xnor U36167 (N_36167,N_22647,N_22686);
or U36168 (N_36168,N_28437,N_21551);
and U36169 (N_36169,N_20109,N_29109);
nor U36170 (N_36170,N_25960,N_27632);
nor U36171 (N_36171,N_20841,N_28772);
xor U36172 (N_36172,N_25667,N_23709);
xor U36173 (N_36173,N_29746,N_21995);
nor U36174 (N_36174,N_26229,N_20561);
nor U36175 (N_36175,N_23056,N_27610);
or U36176 (N_36176,N_25299,N_20441);
nor U36177 (N_36177,N_24668,N_27885);
or U36178 (N_36178,N_22441,N_20521);
nor U36179 (N_36179,N_28432,N_24757);
or U36180 (N_36180,N_27027,N_20130);
or U36181 (N_36181,N_24246,N_24087);
nand U36182 (N_36182,N_29869,N_26906);
nor U36183 (N_36183,N_20876,N_22869);
nand U36184 (N_36184,N_22760,N_26524);
nand U36185 (N_36185,N_28710,N_21761);
xor U36186 (N_36186,N_20260,N_20258);
or U36187 (N_36187,N_23066,N_28016);
nor U36188 (N_36188,N_25734,N_24259);
nor U36189 (N_36189,N_26597,N_24031);
nand U36190 (N_36190,N_21135,N_23582);
nor U36191 (N_36191,N_26806,N_26528);
or U36192 (N_36192,N_21479,N_27824);
and U36193 (N_36193,N_26076,N_27257);
nand U36194 (N_36194,N_25466,N_23511);
xnor U36195 (N_36195,N_29386,N_21551);
and U36196 (N_36196,N_21580,N_22928);
nor U36197 (N_36197,N_20790,N_21010);
and U36198 (N_36198,N_29557,N_24385);
xor U36199 (N_36199,N_22193,N_22745);
nand U36200 (N_36200,N_24380,N_23903);
or U36201 (N_36201,N_27373,N_23579);
nor U36202 (N_36202,N_23829,N_26239);
or U36203 (N_36203,N_25356,N_22552);
nor U36204 (N_36204,N_25998,N_24828);
xnor U36205 (N_36205,N_21738,N_20411);
nor U36206 (N_36206,N_26140,N_26289);
or U36207 (N_36207,N_25045,N_22554);
and U36208 (N_36208,N_23187,N_20829);
xnor U36209 (N_36209,N_24189,N_21279);
xor U36210 (N_36210,N_26849,N_22136);
or U36211 (N_36211,N_28700,N_21505);
and U36212 (N_36212,N_29387,N_26813);
nand U36213 (N_36213,N_25032,N_23887);
and U36214 (N_36214,N_23312,N_20341);
and U36215 (N_36215,N_22113,N_23134);
or U36216 (N_36216,N_29657,N_28748);
nor U36217 (N_36217,N_24838,N_29559);
nand U36218 (N_36218,N_28953,N_24122);
or U36219 (N_36219,N_24456,N_22771);
nor U36220 (N_36220,N_25023,N_28357);
and U36221 (N_36221,N_22331,N_25606);
nor U36222 (N_36222,N_26546,N_27304);
xor U36223 (N_36223,N_25190,N_29511);
nor U36224 (N_36224,N_23317,N_21112);
nor U36225 (N_36225,N_24907,N_21515);
nor U36226 (N_36226,N_29961,N_26463);
xor U36227 (N_36227,N_26333,N_25317);
and U36228 (N_36228,N_27289,N_20576);
nand U36229 (N_36229,N_26530,N_27411);
nand U36230 (N_36230,N_25483,N_25672);
nor U36231 (N_36231,N_25408,N_26257);
xor U36232 (N_36232,N_20677,N_27954);
nor U36233 (N_36233,N_25513,N_24449);
or U36234 (N_36234,N_26448,N_26654);
nor U36235 (N_36235,N_26878,N_20504);
or U36236 (N_36236,N_20849,N_27361);
nand U36237 (N_36237,N_27772,N_27828);
nand U36238 (N_36238,N_23495,N_23460);
nand U36239 (N_36239,N_22418,N_25927);
or U36240 (N_36240,N_24522,N_22754);
xnor U36241 (N_36241,N_27580,N_20921);
nor U36242 (N_36242,N_28141,N_20260);
xnor U36243 (N_36243,N_27807,N_28154);
nor U36244 (N_36244,N_23627,N_27437);
nand U36245 (N_36245,N_27983,N_22711);
xor U36246 (N_36246,N_27282,N_21746);
xor U36247 (N_36247,N_29924,N_27855);
xnor U36248 (N_36248,N_28521,N_21246);
nand U36249 (N_36249,N_22746,N_29416);
nor U36250 (N_36250,N_23365,N_28187);
and U36251 (N_36251,N_20918,N_24466);
and U36252 (N_36252,N_23597,N_28461);
or U36253 (N_36253,N_23216,N_22660);
nor U36254 (N_36254,N_23537,N_28394);
or U36255 (N_36255,N_25891,N_25946);
and U36256 (N_36256,N_27343,N_21401);
and U36257 (N_36257,N_28039,N_24577);
nor U36258 (N_36258,N_23644,N_29854);
xnor U36259 (N_36259,N_21079,N_23783);
xnor U36260 (N_36260,N_25463,N_21646);
xor U36261 (N_36261,N_29672,N_29010);
xor U36262 (N_36262,N_28461,N_23050);
or U36263 (N_36263,N_22139,N_25199);
and U36264 (N_36264,N_29527,N_24476);
and U36265 (N_36265,N_28660,N_25562);
xnor U36266 (N_36266,N_22665,N_23662);
or U36267 (N_36267,N_20545,N_29281);
nand U36268 (N_36268,N_21521,N_21359);
nor U36269 (N_36269,N_20435,N_22693);
xnor U36270 (N_36270,N_21100,N_21761);
and U36271 (N_36271,N_29533,N_20998);
nor U36272 (N_36272,N_22637,N_24868);
or U36273 (N_36273,N_27193,N_22592);
and U36274 (N_36274,N_24061,N_21279);
and U36275 (N_36275,N_22415,N_29666);
nor U36276 (N_36276,N_20263,N_26126);
nand U36277 (N_36277,N_24900,N_23988);
and U36278 (N_36278,N_29591,N_24343);
or U36279 (N_36279,N_28399,N_25508);
nand U36280 (N_36280,N_23944,N_24525);
and U36281 (N_36281,N_24557,N_28763);
and U36282 (N_36282,N_22214,N_23218);
nor U36283 (N_36283,N_20123,N_27873);
xor U36284 (N_36284,N_29344,N_21367);
and U36285 (N_36285,N_29499,N_23460);
or U36286 (N_36286,N_22588,N_25016);
nand U36287 (N_36287,N_21605,N_26408);
nand U36288 (N_36288,N_21916,N_23087);
and U36289 (N_36289,N_21584,N_29127);
and U36290 (N_36290,N_24954,N_23813);
and U36291 (N_36291,N_23202,N_27011);
or U36292 (N_36292,N_28879,N_23853);
xor U36293 (N_36293,N_29629,N_24027);
or U36294 (N_36294,N_27475,N_23864);
nor U36295 (N_36295,N_28084,N_20603);
nor U36296 (N_36296,N_22647,N_22632);
and U36297 (N_36297,N_25593,N_20106);
xnor U36298 (N_36298,N_23612,N_22710);
nand U36299 (N_36299,N_27972,N_25658);
nand U36300 (N_36300,N_28728,N_24295);
or U36301 (N_36301,N_20790,N_20307);
or U36302 (N_36302,N_21331,N_28853);
or U36303 (N_36303,N_26787,N_25581);
and U36304 (N_36304,N_28039,N_20322);
and U36305 (N_36305,N_22287,N_26660);
xor U36306 (N_36306,N_29729,N_27953);
or U36307 (N_36307,N_28574,N_23064);
nand U36308 (N_36308,N_29843,N_26412);
nor U36309 (N_36309,N_23553,N_20963);
or U36310 (N_36310,N_20520,N_21909);
or U36311 (N_36311,N_26100,N_29542);
and U36312 (N_36312,N_23135,N_22121);
and U36313 (N_36313,N_20215,N_23510);
or U36314 (N_36314,N_21085,N_27241);
or U36315 (N_36315,N_24169,N_23605);
or U36316 (N_36316,N_23908,N_26548);
xor U36317 (N_36317,N_29610,N_27310);
nand U36318 (N_36318,N_23203,N_29310);
nand U36319 (N_36319,N_24218,N_24099);
nand U36320 (N_36320,N_26353,N_27799);
nand U36321 (N_36321,N_22538,N_23304);
nand U36322 (N_36322,N_28298,N_23960);
and U36323 (N_36323,N_22174,N_26526);
or U36324 (N_36324,N_24778,N_25484);
nand U36325 (N_36325,N_29589,N_22157);
nor U36326 (N_36326,N_22902,N_24474);
and U36327 (N_36327,N_28248,N_29237);
nand U36328 (N_36328,N_29320,N_25773);
xnor U36329 (N_36329,N_20587,N_23272);
or U36330 (N_36330,N_28555,N_29941);
and U36331 (N_36331,N_21378,N_26009);
or U36332 (N_36332,N_23318,N_20369);
nor U36333 (N_36333,N_29342,N_25938);
nand U36334 (N_36334,N_21454,N_20733);
nand U36335 (N_36335,N_22653,N_25729);
nand U36336 (N_36336,N_22979,N_27503);
or U36337 (N_36337,N_27652,N_24914);
nand U36338 (N_36338,N_20985,N_21523);
or U36339 (N_36339,N_25472,N_21201);
nor U36340 (N_36340,N_24761,N_26599);
or U36341 (N_36341,N_25054,N_23281);
nor U36342 (N_36342,N_28623,N_28913);
nand U36343 (N_36343,N_22869,N_21241);
and U36344 (N_36344,N_27359,N_27878);
xnor U36345 (N_36345,N_25527,N_24809);
nor U36346 (N_36346,N_29173,N_22833);
and U36347 (N_36347,N_26236,N_22768);
xnor U36348 (N_36348,N_24510,N_24777);
or U36349 (N_36349,N_23333,N_27140);
and U36350 (N_36350,N_24575,N_27202);
xnor U36351 (N_36351,N_23908,N_24628);
nor U36352 (N_36352,N_21913,N_21471);
or U36353 (N_36353,N_26049,N_28038);
nor U36354 (N_36354,N_29391,N_26594);
nor U36355 (N_36355,N_26709,N_20332);
and U36356 (N_36356,N_26372,N_25072);
or U36357 (N_36357,N_28681,N_28549);
nand U36358 (N_36358,N_25554,N_28127);
xor U36359 (N_36359,N_21047,N_24749);
nand U36360 (N_36360,N_23544,N_20944);
xor U36361 (N_36361,N_21703,N_21134);
nor U36362 (N_36362,N_20050,N_21012);
and U36363 (N_36363,N_23844,N_25549);
xor U36364 (N_36364,N_25064,N_27223);
nand U36365 (N_36365,N_22917,N_26739);
xor U36366 (N_36366,N_26652,N_22723);
and U36367 (N_36367,N_25593,N_24680);
and U36368 (N_36368,N_23317,N_21904);
and U36369 (N_36369,N_23498,N_21465);
xnor U36370 (N_36370,N_23051,N_28056);
or U36371 (N_36371,N_24050,N_24712);
nand U36372 (N_36372,N_22867,N_22372);
xnor U36373 (N_36373,N_25019,N_25520);
xnor U36374 (N_36374,N_25346,N_28721);
and U36375 (N_36375,N_24226,N_22248);
and U36376 (N_36376,N_20640,N_26559);
xor U36377 (N_36377,N_23144,N_21276);
nand U36378 (N_36378,N_22647,N_26581);
nand U36379 (N_36379,N_25359,N_21389);
or U36380 (N_36380,N_23512,N_25655);
or U36381 (N_36381,N_26118,N_22923);
and U36382 (N_36382,N_27022,N_20098);
nand U36383 (N_36383,N_27937,N_20058);
or U36384 (N_36384,N_24627,N_24551);
nand U36385 (N_36385,N_28055,N_26760);
and U36386 (N_36386,N_22170,N_22662);
and U36387 (N_36387,N_27366,N_27981);
and U36388 (N_36388,N_27734,N_27994);
xnor U36389 (N_36389,N_24023,N_29515);
xor U36390 (N_36390,N_29985,N_28551);
nand U36391 (N_36391,N_27285,N_27479);
nor U36392 (N_36392,N_27006,N_25366);
xor U36393 (N_36393,N_22339,N_28588);
nand U36394 (N_36394,N_27980,N_24525);
and U36395 (N_36395,N_28810,N_29471);
and U36396 (N_36396,N_26038,N_21509);
nand U36397 (N_36397,N_21547,N_21356);
nand U36398 (N_36398,N_27820,N_28205);
nand U36399 (N_36399,N_22212,N_25166);
nand U36400 (N_36400,N_22172,N_26703);
nor U36401 (N_36401,N_20172,N_25357);
xor U36402 (N_36402,N_25407,N_23304);
nor U36403 (N_36403,N_22918,N_27224);
or U36404 (N_36404,N_28741,N_23911);
or U36405 (N_36405,N_27341,N_20673);
nor U36406 (N_36406,N_28397,N_22795);
nor U36407 (N_36407,N_20070,N_25649);
xnor U36408 (N_36408,N_26408,N_26254);
nor U36409 (N_36409,N_20695,N_25339);
nor U36410 (N_36410,N_27922,N_29888);
or U36411 (N_36411,N_22252,N_24451);
and U36412 (N_36412,N_26082,N_28600);
or U36413 (N_36413,N_27446,N_25414);
xnor U36414 (N_36414,N_27495,N_22377);
or U36415 (N_36415,N_22283,N_22103);
nor U36416 (N_36416,N_28743,N_24819);
nor U36417 (N_36417,N_26387,N_23173);
xor U36418 (N_36418,N_29432,N_24702);
or U36419 (N_36419,N_24253,N_27486);
xor U36420 (N_36420,N_20229,N_29909);
or U36421 (N_36421,N_20430,N_25751);
xnor U36422 (N_36422,N_27187,N_27564);
nor U36423 (N_36423,N_29629,N_26506);
nand U36424 (N_36424,N_22574,N_26600);
and U36425 (N_36425,N_27849,N_25560);
nand U36426 (N_36426,N_25283,N_24681);
xor U36427 (N_36427,N_24482,N_27412);
nor U36428 (N_36428,N_29016,N_22444);
or U36429 (N_36429,N_21820,N_24064);
nand U36430 (N_36430,N_26018,N_24523);
xnor U36431 (N_36431,N_22808,N_22613);
xor U36432 (N_36432,N_22805,N_21571);
nor U36433 (N_36433,N_28703,N_23048);
nor U36434 (N_36434,N_25521,N_24889);
nor U36435 (N_36435,N_22747,N_24909);
nor U36436 (N_36436,N_21510,N_26552);
xor U36437 (N_36437,N_28208,N_20773);
nor U36438 (N_36438,N_23925,N_29409);
or U36439 (N_36439,N_21622,N_24677);
and U36440 (N_36440,N_21062,N_23918);
nor U36441 (N_36441,N_27388,N_28354);
nand U36442 (N_36442,N_28537,N_24628);
xnor U36443 (N_36443,N_25510,N_28103);
or U36444 (N_36444,N_28518,N_26350);
nor U36445 (N_36445,N_25685,N_20670);
nand U36446 (N_36446,N_21609,N_25518);
nor U36447 (N_36447,N_28637,N_22878);
nor U36448 (N_36448,N_25482,N_21083);
nor U36449 (N_36449,N_28217,N_27259);
nor U36450 (N_36450,N_25803,N_26883);
xnor U36451 (N_36451,N_24286,N_26910);
and U36452 (N_36452,N_28671,N_22741);
or U36453 (N_36453,N_28919,N_24634);
nor U36454 (N_36454,N_24644,N_21765);
or U36455 (N_36455,N_21649,N_24292);
and U36456 (N_36456,N_27443,N_24859);
nand U36457 (N_36457,N_22271,N_24028);
nand U36458 (N_36458,N_22448,N_27536);
nor U36459 (N_36459,N_23178,N_29962);
or U36460 (N_36460,N_24689,N_21414);
xor U36461 (N_36461,N_26439,N_20836);
nor U36462 (N_36462,N_28260,N_26233);
nand U36463 (N_36463,N_23759,N_27544);
or U36464 (N_36464,N_28568,N_29122);
nor U36465 (N_36465,N_23947,N_24017);
nand U36466 (N_36466,N_28523,N_21676);
and U36467 (N_36467,N_20945,N_21222);
or U36468 (N_36468,N_23487,N_26969);
or U36469 (N_36469,N_24131,N_24121);
nand U36470 (N_36470,N_23785,N_22849);
xor U36471 (N_36471,N_24391,N_21441);
nor U36472 (N_36472,N_23712,N_23274);
xor U36473 (N_36473,N_20198,N_28235);
xnor U36474 (N_36474,N_29862,N_20637);
or U36475 (N_36475,N_20399,N_21751);
nor U36476 (N_36476,N_24818,N_20000);
nor U36477 (N_36477,N_24121,N_27932);
and U36478 (N_36478,N_23640,N_26731);
and U36479 (N_36479,N_22282,N_20612);
or U36480 (N_36480,N_24024,N_24809);
xnor U36481 (N_36481,N_24482,N_27400);
and U36482 (N_36482,N_24014,N_25932);
or U36483 (N_36483,N_24884,N_21871);
xor U36484 (N_36484,N_26519,N_25076);
nand U36485 (N_36485,N_26034,N_25936);
xor U36486 (N_36486,N_21034,N_29201);
nor U36487 (N_36487,N_23686,N_24223);
nand U36488 (N_36488,N_25681,N_29313);
or U36489 (N_36489,N_24480,N_28142);
and U36490 (N_36490,N_24999,N_26873);
or U36491 (N_36491,N_26827,N_27472);
xnor U36492 (N_36492,N_29343,N_20168);
nand U36493 (N_36493,N_25064,N_20884);
nor U36494 (N_36494,N_24061,N_28610);
or U36495 (N_36495,N_24543,N_28728);
nand U36496 (N_36496,N_23102,N_26466);
nor U36497 (N_36497,N_29678,N_26572);
and U36498 (N_36498,N_23126,N_26164);
nand U36499 (N_36499,N_29792,N_23171);
nor U36500 (N_36500,N_21794,N_25523);
nor U36501 (N_36501,N_25101,N_25911);
nand U36502 (N_36502,N_23382,N_21852);
nor U36503 (N_36503,N_20335,N_23501);
xnor U36504 (N_36504,N_29032,N_22068);
or U36505 (N_36505,N_28566,N_25287);
nand U36506 (N_36506,N_21605,N_25502);
or U36507 (N_36507,N_24365,N_21558);
and U36508 (N_36508,N_29563,N_29071);
nor U36509 (N_36509,N_25662,N_25864);
xnor U36510 (N_36510,N_23147,N_27294);
and U36511 (N_36511,N_22103,N_25957);
and U36512 (N_36512,N_26153,N_25364);
nor U36513 (N_36513,N_23065,N_21703);
nand U36514 (N_36514,N_25399,N_27682);
nor U36515 (N_36515,N_29863,N_28018);
and U36516 (N_36516,N_26707,N_26355);
xnor U36517 (N_36517,N_20998,N_25834);
or U36518 (N_36518,N_22161,N_28031);
nand U36519 (N_36519,N_20081,N_26030);
xor U36520 (N_36520,N_22296,N_20332);
nand U36521 (N_36521,N_29810,N_27476);
and U36522 (N_36522,N_27721,N_21682);
nor U36523 (N_36523,N_23478,N_25246);
nand U36524 (N_36524,N_29105,N_28274);
nand U36525 (N_36525,N_26276,N_28149);
nand U36526 (N_36526,N_24879,N_21568);
or U36527 (N_36527,N_25979,N_23106);
nor U36528 (N_36528,N_25299,N_24647);
nand U36529 (N_36529,N_27215,N_25271);
or U36530 (N_36530,N_27788,N_20795);
and U36531 (N_36531,N_20976,N_25697);
and U36532 (N_36532,N_29668,N_27226);
nor U36533 (N_36533,N_24501,N_23811);
or U36534 (N_36534,N_27211,N_22368);
xnor U36535 (N_36535,N_27032,N_24083);
xor U36536 (N_36536,N_21078,N_22242);
xor U36537 (N_36537,N_21858,N_21119);
nor U36538 (N_36538,N_25062,N_23694);
nor U36539 (N_36539,N_25304,N_23581);
nand U36540 (N_36540,N_22123,N_26507);
nand U36541 (N_36541,N_20437,N_28081);
and U36542 (N_36542,N_29256,N_22908);
nand U36543 (N_36543,N_27578,N_24425);
nor U36544 (N_36544,N_25698,N_25419);
or U36545 (N_36545,N_22739,N_20846);
nor U36546 (N_36546,N_21631,N_27498);
xnor U36547 (N_36547,N_22094,N_27066);
nand U36548 (N_36548,N_24846,N_25582);
and U36549 (N_36549,N_28793,N_26785);
or U36550 (N_36550,N_25271,N_23270);
xnor U36551 (N_36551,N_26900,N_20271);
nor U36552 (N_36552,N_22404,N_26606);
or U36553 (N_36553,N_27088,N_29374);
xnor U36554 (N_36554,N_24062,N_29228);
and U36555 (N_36555,N_25236,N_26158);
or U36556 (N_36556,N_29324,N_24944);
xor U36557 (N_36557,N_21137,N_29481);
nor U36558 (N_36558,N_22069,N_23969);
xor U36559 (N_36559,N_24803,N_28542);
nor U36560 (N_36560,N_25126,N_20836);
nand U36561 (N_36561,N_24984,N_25846);
and U36562 (N_36562,N_27253,N_29887);
xnor U36563 (N_36563,N_21144,N_21339);
and U36564 (N_36564,N_28111,N_27618);
and U36565 (N_36565,N_20763,N_24658);
nor U36566 (N_36566,N_22421,N_23547);
or U36567 (N_36567,N_25806,N_20434);
or U36568 (N_36568,N_29083,N_29009);
nor U36569 (N_36569,N_27658,N_21561);
or U36570 (N_36570,N_27499,N_20252);
and U36571 (N_36571,N_20446,N_24161);
nand U36572 (N_36572,N_23652,N_23326);
xnor U36573 (N_36573,N_28724,N_24215);
or U36574 (N_36574,N_28121,N_28466);
and U36575 (N_36575,N_28637,N_25414);
xor U36576 (N_36576,N_27548,N_23554);
or U36577 (N_36577,N_24691,N_23258);
xor U36578 (N_36578,N_27462,N_20694);
or U36579 (N_36579,N_26571,N_23604);
nor U36580 (N_36580,N_20036,N_27376);
and U36581 (N_36581,N_28387,N_25420);
nor U36582 (N_36582,N_28836,N_20088);
or U36583 (N_36583,N_27123,N_22589);
nor U36584 (N_36584,N_29636,N_28865);
nor U36585 (N_36585,N_25599,N_29242);
nand U36586 (N_36586,N_27808,N_20355);
and U36587 (N_36587,N_27773,N_27755);
xnor U36588 (N_36588,N_24283,N_25581);
xor U36589 (N_36589,N_21862,N_26051);
nor U36590 (N_36590,N_26626,N_24588);
nand U36591 (N_36591,N_21307,N_20848);
xor U36592 (N_36592,N_29757,N_20913);
or U36593 (N_36593,N_21218,N_26133);
and U36594 (N_36594,N_25025,N_26156);
nor U36595 (N_36595,N_29551,N_29573);
or U36596 (N_36596,N_29182,N_23674);
nand U36597 (N_36597,N_20666,N_25439);
nand U36598 (N_36598,N_28412,N_29088);
xnor U36599 (N_36599,N_20026,N_25208);
xnor U36600 (N_36600,N_26027,N_28532);
xnor U36601 (N_36601,N_28165,N_21896);
and U36602 (N_36602,N_27390,N_23220);
xor U36603 (N_36603,N_23243,N_29264);
nor U36604 (N_36604,N_21806,N_25259);
or U36605 (N_36605,N_27962,N_21462);
or U36606 (N_36606,N_26038,N_20590);
xnor U36607 (N_36607,N_28010,N_25947);
and U36608 (N_36608,N_26177,N_24916);
nor U36609 (N_36609,N_24314,N_20760);
nand U36610 (N_36610,N_24910,N_25723);
nor U36611 (N_36611,N_28982,N_23833);
or U36612 (N_36612,N_27107,N_27841);
xor U36613 (N_36613,N_23438,N_29324);
nand U36614 (N_36614,N_21762,N_27726);
or U36615 (N_36615,N_22399,N_28832);
nor U36616 (N_36616,N_24131,N_29558);
nor U36617 (N_36617,N_28743,N_29024);
and U36618 (N_36618,N_23338,N_29347);
and U36619 (N_36619,N_20500,N_21095);
or U36620 (N_36620,N_20402,N_24102);
nor U36621 (N_36621,N_26309,N_20634);
nand U36622 (N_36622,N_26793,N_20150);
nand U36623 (N_36623,N_26087,N_27324);
and U36624 (N_36624,N_22059,N_21147);
nor U36625 (N_36625,N_22786,N_22011);
and U36626 (N_36626,N_27138,N_28753);
or U36627 (N_36627,N_23724,N_28327);
nor U36628 (N_36628,N_22286,N_21629);
xnor U36629 (N_36629,N_23225,N_20258);
xnor U36630 (N_36630,N_20136,N_28492);
or U36631 (N_36631,N_20073,N_28941);
xor U36632 (N_36632,N_26864,N_29170);
xor U36633 (N_36633,N_26733,N_21159);
xnor U36634 (N_36634,N_23513,N_25207);
or U36635 (N_36635,N_21544,N_26225);
and U36636 (N_36636,N_22550,N_22894);
and U36637 (N_36637,N_29851,N_27553);
and U36638 (N_36638,N_28268,N_24033);
or U36639 (N_36639,N_20954,N_21194);
xor U36640 (N_36640,N_25711,N_25211);
nand U36641 (N_36641,N_20867,N_24919);
nand U36642 (N_36642,N_25836,N_26095);
nor U36643 (N_36643,N_23271,N_27042);
nor U36644 (N_36644,N_26459,N_24488);
nand U36645 (N_36645,N_23732,N_28183);
nand U36646 (N_36646,N_24421,N_29491);
and U36647 (N_36647,N_23895,N_23505);
or U36648 (N_36648,N_21216,N_23079);
xor U36649 (N_36649,N_26571,N_20263);
or U36650 (N_36650,N_20256,N_29695);
xor U36651 (N_36651,N_21725,N_21929);
nor U36652 (N_36652,N_25455,N_29638);
or U36653 (N_36653,N_29828,N_21562);
nand U36654 (N_36654,N_26949,N_26718);
nand U36655 (N_36655,N_24976,N_25803);
nand U36656 (N_36656,N_29571,N_21524);
nor U36657 (N_36657,N_23057,N_24441);
nand U36658 (N_36658,N_23369,N_25576);
and U36659 (N_36659,N_29218,N_23597);
xor U36660 (N_36660,N_21719,N_21802);
nand U36661 (N_36661,N_28452,N_27805);
nand U36662 (N_36662,N_21446,N_20119);
xor U36663 (N_36663,N_25125,N_22932);
nor U36664 (N_36664,N_20001,N_27014);
nor U36665 (N_36665,N_26818,N_21995);
nor U36666 (N_36666,N_24009,N_26145);
nand U36667 (N_36667,N_27755,N_23064);
xor U36668 (N_36668,N_26017,N_22332);
nor U36669 (N_36669,N_21784,N_23838);
nor U36670 (N_36670,N_25483,N_26269);
and U36671 (N_36671,N_27706,N_23628);
nand U36672 (N_36672,N_21931,N_26607);
nor U36673 (N_36673,N_26388,N_23564);
xor U36674 (N_36674,N_20895,N_23324);
nand U36675 (N_36675,N_29969,N_22229);
nor U36676 (N_36676,N_25425,N_25998);
or U36677 (N_36677,N_29141,N_24768);
nand U36678 (N_36678,N_23760,N_22568);
xnor U36679 (N_36679,N_24929,N_24178);
or U36680 (N_36680,N_29009,N_29077);
or U36681 (N_36681,N_23582,N_20607);
nor U36682 (N_36682,N_24301,N_24938);
nand U36683 (N_36683,N_25462,N_20579);
or U36684 (N_36684,N_22716,N_24238);
or U36685 (N_36685,N_24770,N_27385);
or U36686 (N_36686,N_29096,N_26560);
or U36687 (N_36687,N_29571,N_25939);
nor U36688 (N_36688,N_28106,N_28099);
nand U36689 (N_36689,N_26317,N_21021);
and U36690 (N_36690,N_27112,N_28404);
or U36691 (N_36691,N_23648,N_21235);
nor U36692 (N_36692,N_27178,N_25708);
nor U36693 (N_36693,N_29191,N_21808);
xnor U36694 (N_36694,N_29085,N_24283);
nor U36695 (N_36695,N_20306,N_20226);
nand U36696 (N_36696,N_21163,N_27185);
nand U36697 (N_36697,N_29937,N_29029);
and U36698 (N_36698,N_21512,N_23284);
nand U36699 (N_36699,N_23442,N_25812);
nor U36700 (N_36700,N_22638,N_23740);
and U36701 (N_36701,N_29002,N_20490);
xnor U36702 (N_36702,N_22009,N_29954);
xor U36703 (N_36703,N_29329,N_24111);
nand U36704 (N_36704,N_22572,N_24887);
xor U36705 (N_36705,N_29765,N_25992);
nand U36706 (N_36706,N_23091,N_27307);
or U36707 (N_36707,N_22790,N_29719);
nor U36708 (N_36708,N_20440,N_29155);
or U36709 (N_36709,N_25923,N_27032);
xor U36710 (N_36710,N_24983,N_27977);
or U36711 (N_36711,N_29660,N_20748);
nand U36712 (N_36712,N_26049,N_24853);
nor U36713 (N_36713,N_20391,N_26035);
nor U36714 (N_36714,N_22810,N_22550);
nand U36715 (N_36715,N_28196,N_22918);
and U36716 (N_36716,N_24838,N_26060);
and U36717 (N_36717,N_28246,N_26479);
and U36718 (N_36718,N_29197,N_20476);
xor U36719 (N_36719,N_29873,N_23392);
and U36720 (N_36720,N_22255,N_27702);
nand U36721 (N_36721,N_25601,N_25901);
xnor U36722 (N_36722,N_27188,N_22456);
and U36723 (N_36723,N_27047,N_20122);
xor U36724 (N_36724,N_28824,N_25403);
and U36725 (N_36725,N_27314,N_20560);
xnor U36726 (N_36726,N_22146,N_20025);
nand U36727 (N_36727,N_27733,N_21319);
xor U36728 (N_36728,N_25968,N_20369);
xnor U36729 (N_36729,N_21221,N_20619);
nor U36730 (N_36730,N_29556,N_23264);
or U36731 (N_36731,N_28251,N_26889);
nor U36732 (N_36732,N_23345,N_22508);
nor U36733 (N_36733,N_28787,N_24672);
nor U36734 (N_36734,N_24728,N_23264);
nor U36735 (N_36735,N_24523,N_23550);
nand U36736 (N_36736,N_23670,N_28267);
xor U36737 (N_36737,N_23005,N_20353);
xor U36738 (N_36738,N_25021,N_28515);
nand U36739 (N_36739,N_20196,N_20254);
and U36740 (N_36740,N_22424,N_28183);
xor U36741 (N_36741,N_27739,N_21976);
nor U36742 (N_36742,N_25814,N_27525);
nor U36743 (N_36743,N_28990,N_21403);
xor U36744 (N_36744,N_23878,N_22124);
or U36745 (N_36745,N_20507,N_22947);
or U36746 (N_36746,N_26091,N_28639);
nand U36747 (N_36747,N_23995,N_24001);
nand U36748 (N_36748,N_22359,N_28070);
or U36749 (N_36749,N_25982,N_22595);
nor U36750 (N_36750,N_22543,N_24707);
xnor U36751 (N_36751,N_28191,N_27947);
or U36752 (N_36752,N_29347,N_28228);
xnor U36753 (N_36753,N_25585,N_21342);
or U36754 (N_36754,N_29736,N_20557);
or U36755 (N_36755,N_27313,N_26266);
or U36756 (N_36756,N_24992,N_28305);
or U36757 (N_36757,N_20217,N_21175);
nand U36758 (N_36758,N_23184,N_22611);
and U36759 (N_36759,N_28357,N_23535);
nand U36760 (N_36760,N_20484,N_27614);
nand U36761 (N_36761,N_28207,N_28769);
or U36762 (N_36762,N_26986,N_22542);
or U36763 (N_36763,N_29928,N_26151);
nor U36764 (N_36764,N_27410,N_26910);
xnor U36765 (N_36765,N_28046,N_20919);
and U36766 (N_36766,N_26287,N_24647);
nor U36767 (N_36767,N_28583,N_24741);
or U36768 (N_36768,N_20887,N_20727);
and U36769 (N_36769,N_28803,N_24688);
or U36770 (N_36770,N_25753,N_22576);
nor U36771 (N_36771,N_29590,N_22668);
and U36772 (N_36772,N_27254,N_22059);
nand U36773 (N_36773,N_25378,N_27960);
nor U36774 (N_36774,N_20863,N_23239);
nand U36775 (N_36775,N_23024,N_26771);
xnor U36776 (N_36776,N_25469,N_25290);
xor U36777 (N_36777,N_25311,N_22111);
or U36778 (N_36778,N_27867,N_28871);
nor U36779 (N_36779,N_24919,N_25664);
and U36780 (N_36780,N_24898,N_22818);
nand U36781 (N_36781,N_24126,N_22966);
or U36782 (N_36782,N_21684,N_25991);
or U36783 (N_36783,N_22818,N_25644);
nor U36784 (N_36784,N_26875,N_24096);
nor U36785 (N_36785,N_20886,N_26343);
and U36786 (N_36786,N_28371,N_22736);
nor U36787 (N_36787,N_25274,N_21409);
nand U36788 (N_36788,N_27383,N_21587);
or U36789 (N_36789,N_23867,N_27138);
and U36790 (N_36790,N_20021,N_28823);
and U36791 (N_36791,N_29556,N_23073);
and U36792 (N_36792,N_24170,N_26392);
or U36793 (N_36793,N_26287,N_26528);
nor U36794 (N_36794,N_23528,N_21360);
nand U36795 (N_36795,N_28734,N_22902);
and U36796 (N_36796,N_23561,N_25748);
and U36797 (N_36797,N_28188,N_22236);
and U36798 (N_36798,N_23256,N_23614);
xnor U36799 (N_36799,N_24611,N_21796);
nor U36800 (N_36800,N_20379,N_20948);
nand U36801 (N_36801,N_29520,N_26673);
nand U36802 (N_36802,N_21045,N_21189);
nand U36803 (N_36803,N_25424,N_22454);
or U36804 (N_36804,N_27751,N_20843);
nand U36805 (N_36805,N_22732,N_23027);
nor U36806 (N_36806,N_26707,N_21426);
or U36807 (N_36807,N_29254,N_25264);
nor U36808 (N_36808,N_29679,N_26678);
nand U36809 (N_36809,N_24963,N_22965);
or U36810 (N_36810,N_25591,N_25889);
nand U36811 (N_36811,N_24309,N_28356);
xnor U36812 (N_36812,N_29941,N_27657);
or U36813 (N_36813,N_27561,N_21115);
or U36814 (N_36814,N_24750,N_21006);
nor U36815 (N_36815,N_21800,N_22633);
and U36816 (N_36816,N_22170,N_22081);
nor U36817 (N_36817,N_29231,N_29390);
nand U36818 (N_36818,N_23617,N_21604);
nor U36819 (N_36819,N_22303,N_25297);
xnor U36820 (N_36820,N_29777,N_24311);
nand U36821 (N_36821,N_28961,N_24641);
or U36822 (N_36822,N_24974,N_24122);
nor U36823 (N_36823,N_22390,N_28645);
nor U36824 (N_36824,N_28854,N_20026);
nand U36825 (N_36825,N_27553,N_22225);
or U36826 (N_36826,N_21106,N_29512);
nor U36827 (N_36827,N_28994,N_25186);
nand U36828 (N_36828,N_28890,N_25381);
nand U36829 (N_36829,N_22526,N_29097);
nand U36830 (N_36830,N_22930,N_20968);
nand U36831 (N_36831,N_24588,N_22655);
xnor U36832 (N_36832,N_20659,N_20613);
nor U36833 (N_36833,N_23873,N_29332);
nand U36834 (N_36834,N_29509,N_23830);
xnor U36835 (N_36835,N_22423,N_27971);
and U36836 (N_36836,N_29031,N_28270);
and U36837 (N_36837,N_26733,N_22503);
nor U36838 (N_36838,N_22512,N_27958);
nor U36839 (N_36839,N_21751,N_20494);
xor U36840 (N_36840,N_20907,N_24492);
or U36841 (N_36841,N_24999,N_20318);
nand U36842 (N_36842,N_23322,N_27886);
or U36843 (N_36843,N_21800,N_26124);
nand U36844 (N_36844,N_28123,N_26028);
and U36845 (N_36845,N_22190,N_27828);
nand U36846 (N_36846,N_22770,N_27584);
nand U36847 (N_36847,N_22832,N_29362);
xor U36848 (N_36848,N_24954,N_29686);
and U36849 (N_36849,N_21236,N_26369);
nor U36850 (N_36850,N_28650,N_24776);
or U36851 (N_36851,N_27123,N_28009);
or U36852 (N_36852,N_20853,N_27815);
nand U36853 (N_36853,N_23728,N_25863);
and U36854 (N_36854,N_26352,N_27909);
nand U36855 (N_36855,N_24271,N_28143);
xor U36856 (N_36856,N_27346,N_27588);
nor U36857 (N_36857,N_20639,N_24946);
nand U36858 (N_36858,N_21130,N_22276);
or U36859 (N_36859,N_24229,N_20485);
or U36860 (N_36860,N_22039,N_28639);
or U36861 (N_36861,N_20934,N_25179);
xnor U36862 (N_36862,N_22774,N_20373);
nand U36863 (N_36863,N_29918,N_29542);
nor U36864 (N_36864,N_27465,N_25400);
nand U36865 (N_36865,N_28753,N_20026);
nor U36866 (N_36866,N_22432,N_25398);
xor U36867 (N_36867,N_20190,N_29649);
xor U36868 (N_36868,N_23036,N_21770);
or U36869 (N_36869,N_23998,N_25838);
nand U36870 (N_36870,N_21848,N_25800);
xnor U36871 (N_36871,N_24153,N_20894);
and U36872 (N_36872,N_28924,N_28862);
and U36873 (N_36873,N_27924,N_25260);
xnor U36874 (N_36874,N_27410,N_23964);
xnor U36875 (N_36875,N_26855,N_25362);
or U36876 (N_36876,N_21933,N_20290);
xnor U36877 (N_36877,N_29303,N_26332);
xnor U36878 (N_36878,N_29070,N_26246);
and U36879 (N_36879,N_21742,N_25945);
and U36880 (N_36880,N_20321,N_26427);
nand U36881 (N_36881,N_27210,N_20364);
and U36882 (N_36882,N_25035,N_23781);
xor U36883 (N_36883,N_20729,N_26668);
xor U36884 (N_36884,N_24026,N_21281);
and U36885 (N_36885,N_25954,N_23800);
nor U36886 (N_36886,N_29748,N_23888);
and U36887 (N_36887,N_26986,N_20873);
nand U36888 (N_36888,N_20698,N_26412);
or U36889 (N_36889,N_21275,N_22062);
nor U36890 (N_36890,N_29763,N_21101);
xnor U36891 (N_36891,N_22775,N_26797);
xor U36892 (N_36892,N_24038,N_22171);
and U36893 (N_36893,N_23184,N_21388);
or U36894 (N_36894,N_20991,N_23744);
xnor U36895 (N_36895,N_24589,N_20376);
and U36896 (N_36896,N_29972,N_29289);
or U36897 (N_36897,N_24455,N_26499);
nor U36898 (N_36898,N_25359,N_25278);
or U36899 (N_36899,N_20471,N_25496);
nand U36900 (N_36900,N_24682,N_22762);
and U36901 (N_36901,N_25046,N_24802);
nor U36902 (N_36902,N_26169,N_25583);
and U36903 (N_36903,N_29421,N_26808);
nor U36904 (N_36904,N_25865,N_28495);
nand U36905 (N_36905,N_29186,N_26818);
nor U36906 (N_36906,N_25933,N_25544);
xnor U36907 (N_36907,N_27932,N_21613);
xnor U36908 (N_36908,N_25053,N_28655);
nand U36909 (N_36909,N_21114,N_27572);
xor U36910 (N_36910,N_23788,N_29404);
xnor U36911 (N_36911,N_24277,N_25181);
xor U36912 (N_36912,N_22548,N_21727);
nor U36913 (N_36913,N_23156,N_28915);
and U36914 (N_36914,N_28954,N_27732);
nor U36915 (N_36915,N_22877,N_25034);
or U36916 (N_36916,N_22327,N_29114);
xnor U36917 (N_36917,N_23547,N_28208);
nor U36918 (N_36918,N_28638,N_25380);
nand U36919 (N_36919,N_25930,N_25767);
or U36920 (N_36920,N_28896,N_20751);
and U36921 (N_36921,N_23428,N_21758);
or U36922 (N_36922,N_27956,N_27830);
and U36923 (N_36923,N_27298,N_22377);
nand U36924 (N_36924,N_23621,N_20280);
nor U36925 (N_36925,N_24736,N_20438);
xor U36926 (N_36926,N_21848,N_26032);
nand U36927 (N_36927,N_20410,N_23348);
nor U36928 (N_36928,N_29232,N_22825);
xor U36929 (N_36929,N_21231,N_27978);
or U36930 (N_36930,N_28521,N_26529);
or U36931 (N_36931,N_23582,N_27008);
nor U36932 (N_36932,N_20872,N_20071);
and U36933 (N_36933,N_26068,N_27732);
xnor U36934 (N_36934,N_29886,N_20172);
nand U36935 (N_36935,N_21694,N_28176);
nor U36936 (N_36936,N_27431,N_20433);
nor U36937 (N_36937,N_22601,N_25165);
nand U36938 (N_36938,N_23880,N_29210);
nand U36939 (N_36939,N_20388,N_21871);
nand U36940 (N_36940,N_23880,N_20897);
nand U36941 (N_36941,N_25928,N_23010);
or U36942 (N_36942,N_23255,N_29911);
and U36943 (N_36943,N_23351,N_26140);
nor U36944 (N_36944,N_24024,N_25894);
xor U36945 (N_36945,N_27088,N_21195);
nor U36946 (N_36946,N_22313,N_25198);
or U36947 (N_36947,N_21556,N_23116);
or U36948 (N_36948,N_23022,N_26310);
and U36949 (N_36949,N_28612,N_29499);
xor U36950 (N_36950,N_26683,N_27328);
nor U36951 (N_36951,N_29742,N_24607);
nor U36952 (N_36952,N_21790,N_24275);
or U36953 (N_36953,N_27869,N_22408);
and U36954 (N_36954,N_28651,N_29978);
or U36955 (N_36955,N_23530,N_26541);
nor U36956 (N_36956,N_28104,N_20810);
nor U36957 (N_36957,N_25769,N_24712);
or U36958 (N_36958,N_22600,N_24637);
nor U36959 (N_36959,N_22442,N_22870);
nand U36960 (N_36960,N_25771,N_20020);
and U36961 (N_36961,N_25441,N_24706);
nor U36962 (N_36962,N_26721,N_20250);
xnor U36963 (N_36963,N_28329,N_26310);
nand U36964 (N_36964,N_24881,N_21999);
nor U36965 (N_36965,N_20810,N_28414);
and U36966 (N_36966,N_20281,N_23634);
or U36967 (N_36967,N_25043,N_23360);
and U36968 (N_36968,N_27790,N_22690);
nand U36969 (N_36969,N_27038,N_24691);
xnor U36970 (N_36970,N_21534,N_25276);
nor U36971 (N_36971,N_20993,N_20797);
and U36972 (N_36972,N_29684,N_24234);
xor U36973 (N_36973,N_24957,N_29789);
nand U36974 (N_36974,N_29844,N_26880);
nand U36975 (N_36975,N_20658,N_27135);
xor U36976 (N_36976,N_22698,N_23480);
nor U36977 (N_36977,N_28697,N_24791);
xnor U36978 (N_36978,N_26323,N_25445);
and U36979 (N_36979,N_24528,N_23132);
or U36980 (N_36980,N_20799,N_20849);
nand U36981 (N_36981,N_25648,N_23878);
and U36982 (N_36982,N_20605,N_29737);
nand U36983 (N_36983,N_20139,N_20160);
or U36984 (N_36984,N_26667,N_23452);
nor U36985 (N_36985,N_21393,N_26278);
and U36986 (N_36986,N_23961,N_20022);
or U36987 (N_36987,N_22718,N_22653);
xnor U36988 (N_36988,N_26846,N_29845);
xnor U36989 (N_36989,N_28223,N_21994);
and U36990 (N_36990,N_20829,N_20285);
and U36991 (N_36991,N_29706,N_23425);
or U36992 (N_36992,N_25660,N_23180);
nand U36993 (N_36993,N_24300,N_23101);
nand U36994 (N_36994,N_29775,N_29640);
and U36995 (N_36995,N_22555,N_22051);
and U36996 (N_36996,N_20174,N_23938);
xor U36997 (N_36997,N_23259,N_28980);
xor U36998 (N_36998,N_22187,N_20239);
nand U36999 (N_36999,N_23675,N_23362);
xnor U37000 (N_37000,N_25399,N_20458);
nand U37001 (N_37001,N_24860,N_27243);
nor U37002 (N_37002,N_29606,N_20384);
and U37003 (N_37003,N_27816,N_24971);
xor U37004 (N_37004,N_26944,N_24570);
and U37005 (N_37005,N_24649,N_24189);
nor U37006 (N_37006,N_25211,N_26904);
nor U37007 (N_37007,N_29526,N_22606);
or U37008 (N_37008,N_20731,N_27340);
and U37009 (N_37009,N_26576,N_23330);
nand U37010 (N_37010,N_22512,N_21264);
xor U37011 (N_37011,N_24867,N_26528);
and U37012 (N_37012,N_26337,N_21667);
nand U37013 (N_37013,N_28194,N_29934);
and U37014 (N_37014,N_20074,N_23921);
nor U37015 (N_37015,N_24465,N_21315);
and U37016 (N_37016,N_29968,N_23803);
xor U37017 (N_37017,N_20348,N_24430);
nand U37018 (N_37018,N_21506,N_21867);
nand U37019 (N_37019,N_25050,N_28622);
xor U37020 (N_37020,N_21386,N_26960);
nand U37021 (N_37021,N_23867,N_23405);
and U37022 (N_37022,N_26456,N_29734);
and U37023 (N_37023,N_24661,N_25160);
nand U37024 (N_37024,N_23746,N_26215);
xnor U37025 (N_37025,N_26910,N_28182);
nor U37026 (N_37026,N_24934,N_24313);
nand U37027 (N_37027,N_22019,N_20448);
nand U37028 (N_37028,N_26375,N_21075);
xor U37029 (N_37029,N_27697,N_21267);
and U37030 (N_37030,N_23046,N_23051);
nand U37031 (N_37031,N_29910,N_24414);
nand U37032 (N_37032,N_25204,N_23988);
or U37033 (N_37033,N_21654,N_22240);
nor U37034 (N_37034,N_21296,N_22431);
or U37035 (N_37035,N_26622,N_25611);
or U37036 (N_37036,N_24315,N_25837);
xnor U37037 (N_37037,N_29019,N_28978);
xnor U37038 (N_37038,N_25340,N_28166);
xor U37039 (N_37039,N_20208,N_25034);
nor U37040 (N_37040,N_21923,N_26635);
nor U37041 (N_37041,N_24647,N_25382);
nand U37042 (N_37042,N_27434,N_20367);
or U37043 (N_37043,N_29964,N_21449);
nor U37044 (N_37044,N_22976,N_29894);
or U37045 (N_37045,N_26680,N_29054);
nand U37046 (N_37046,N_28171,N_24450);
and U37047 (N_37047,N_24648,N_25844);
nor U37048 (N_37048,N_21635,N_23499);
nand U37049 (N_37049,N_25854,N_29938);
xor U37050 (N_37050,N_25665,N_29858);
or U37051 (N_37051,N_21051,N_29649);
and U37052 (N_37052,N_21855,N_20438);
nand U37053 (N_37053,N_29345,N_26442);
or U37054 (N_37054,N_28787,N_23871);
nor U37055 (N_37055,N_25385,N_25356);
and U37056 (N_37056,N_27132,N_24614);
nand U37057 (N_37057,N_24483,N_23533);
xnor U37058 (N_37058,N_23612,N_29038);
nand U37059 (N_37059,N_29907,N_23731);
xnor U37060 (N_37060,N_28382,N_29746);
nand U37061 (N_37061,N_22712,N_27243);
and U37062 (N_37062,N_26444,N_23199);
or U37063 (N_37063,N_25061,N_29245);
nor U37064 (N_37064,N_27105,N_21647);
and U37065 (N_37065,N_26896,N_26400);
nor U37066 (N_37066,N_21391,N_26084);
and U37067 (N_37067,N_22835,N_21345);
nor U37068 (N_37068,N_25414,N_20783);
nand U37069 (N_37069,N_28628,N_25738);
nand U37070 (N_37070,N_24294,N_20329);
and U37071 (N_37071,N_24708,N_29146);
nor U37072 (N_37072,N_23884,N_27712);
xnor U37073 (N_37073,N_26892,N_20701);
nand U37074 (N_37074,N_26934,N_23408);
xor U37075 (N_37075,N_22230,N_29037);
xor U37076 (N_37076,N_20313,N_22261);
and U37077 (N_37077,N_22158,N_26258);
nor U37078 (N_37078,N_21985,N_26611);
and U37079 (N_37079,N_20731,N_24201);
or U37080 (N_37080,N_22921,N_23445);
or U37081 (N_37081,N_26842,N_27467);
nand U37082 (N_37082,N_25481,N_29588);
and U37083 (N_37083,N_29211,N_28677);
or U37084 (N_37084,N_25201,N_26894);
or U37085 (N_37085,N_23723,N_20384);
nor U37086 (N_37086,N_24366,N_29277);
or U37087 (N_37087,N_28683,N_29884);
or U37088 (N_37088,N_28272,N_26893);
and U37089 (N_37089,N_22025,N_25174);
or U37090 (N_37090,N_23348,N_21357);
or U37091 (N_37091,N_29942,N_24608);
or U37092 (N_37092,N_21454,N_28525);
xor U37093 (N_37093,N_22522,N_21833);
nand U37094 (N_37094,N_25904,N_23436);
and U37095 (N_37095,N_27968,N_29989);
xor U37096 (N_37096,N_22387,N_22055);
or U37097 (N_37097,N_23886,N_27370);
xor U37098 (N_37098,N_27562,N_23734);
and U37099 (N_37099,N_23685,N_27452);
xnor U37100 (N_37100,N_21121,N_25225);
and U37101 (N_37101,N_23778,N_20381);
nand U37102 (N_37102,N_27264,N_29666);
xnor U37103 (N_37103,N_23617,N_25472);
and U37104 (N_37104,N_29408,N_27151);
nor U37105 (N_37105,N_26126,N_27676);
xnor U37106 (N_37106,N_20765,N_21770);
nand U37107 (N_37107,N_21763,N_27306);
xnor U37108 (N_37108,N_29409,N_23476);
nor U37109 (N_37109,N_21037,N_27339);
xor U37110 (N_37110,N_24859,N_29173);
xor U37111 (N_37111,N_24248,N_23939);
and U37112 (N_37112,N_28983,N_25292);
and U37113 (N_37113,N_27119,N_27726);
nor U37114 (N_37114,N_25835,N_25286);
nor U37115 (N_37115,N_20709,N_29105);
nand U37116 (N_37116,N_25113,N_26147);
nor U37117 (N_37117,N_25529,N_20997);
nand U37118 (N_37118,N_27279,N_26782);
and U37119 (N_37119,N_20097,N_20068);
and U37120 (N_37120,N_26981,N_25898);
or U37121 (N_37121,N_22482,N_20698);
xnor U37122 (N_37122,N_27162,N_20774);
and U37123 (N_37123,N_22633,N_23233);
or U37124 (N_37124,N_20002,N_25060);
or U37125 (N_37125,N_20788,N_29567);
and U37126 (N_37126,N_23628,N_22001);
nand U37127 (N_37127,N_25203,N_27548);
xnor U37128 (N_37128,N_20509,N_24513);
nor U37129 (N_37129,N_29317,N_24700);
or U37130 (N_37130,N_27099,N_29677);
or U37131 (N_37131,N_29695,N_27239);
xor U37132 (N_37132,N_25810,N_27954);
xor U37133 (N_37133,N_23240,N_28732);
xnor U37134 (N_37134,N_25406,N_26574);
xor U37135 (N_37135,N_24420,N_28959);
nand U37136 (N_37136,N_28928,N_22857);
or U37137 (N_37137,N_28355,N_22533);
or U37138 (N_37138,N_22336,N_29268);
or U37139 (N_37139,N_23713,N_26430);
nor U37140 (N_37140,N_22276,N_23201);
and U37141 (N_37141,N_25169,N_29318);
or U37142 (N_37142,N_24264,N_27253);
nor U37143 (N_37143,N_26268,N_22138);
nor U37144 (N_37144,N_26610,N_21597);
nand U37145 (N_37145,N_24589,N_22328);
or U37146 (N_37146,N_21102,N_28697);
nand U37147 (N_37147,N_22214,N_28321);
nand U37148 (N_37148,N_26085,N_28744);
xnor U37149 (N_37149,N_21258,N_25980);
or U37150 (N_37150,N_28056,N_21302);
nand U37151 (N_37151,N_27558,N_28094);
or U37152 (N_37152,N_27308,N_21338);
xnor U37153 (N_37153,N_26353,N_25296);
or U37154 (N_37154,N_22556,N_24797);
xnor U37155 (N_37155,N_22217,N_22751);
xnor U37156 (N_37156,N_22678,N_23732);
nor U37157 (N_37157,N_21836,N_25031);
and U37158 (N_37158,N_26327,N_26472);
or U37159 (N_37159,N_25877,N_21804);
nand U37160 (N_37160,N_25073,N_23303);
nor U37161 (N_37161,N_29142,N_26934);
or U37162 (N_37162,N_20666,N_24208);
or U37163 (N_37163,N_20218,N_22459);
nor U37164 (N_37164,N_21981,N_23526);
and U37165 (N_37165,N_21964,N_24744);
or U37166 (N_37166,N_20941,N_20371);
xnor U37167 (N_37167,N_27202,N_25011);
xor U37168 (N_37168,N_27562,N_28527);
nand U37169 (N_37169,N_23232,N_21779);
or U37170 (N_37170,N_27698,N_29558);
nand U37171 (N_37171,N_29014,N_24338);
nor U37172 (N_37172,N_22613,N_25745);
nor U37173 (N_37173,N_26321,N_29529);
nand U37174 (N_37174,N_29253,N_27046);
xnor U37175 (N_37175,N_20515,N_27878);
and U37176 (N_37176,N_28090,N_27536);
xor U37177 (N_37177,N_21119,N_21050);
nand U37178 (N_37178,N_24545,N_29106);
or U37179 (N_37179,N_21120,N_22480);
or U37180 (N_37180,N_20098,N_23653);
nor U37181 (N_37181,N_25338,N_25503);
and U37182 (N_37182,N_23056,N_24267);
or U37183 (N_37183,N_25398,N_26119);
nand U37184 (N_37184,N_26543,N_22267);
and U37185 (N_37185,N_20441,N_28321);
nor U37186 (N_37186,N_20398,N_29992);
nand U37187 (N_37187,N_25256,N_20844);
or U37188 (N_37188,N_20172,N_23737);
nand U37189 (N_37189,N_22890,N_26823);
nor U37190 (N_37190,N_25859,N_28330);
and U37191 (N_37191,N_23260,N_21115);
xnor U37192 (N_37192,N_26699,N_27840);
or U37193 (N_37193,N_28575,N_24681);
nand U37194 (N_37194,N_25441,N_22365);
xnor U37195 (N_37195,N_21678,N_26312);
nand U37196 (N_37196,N_24472,N_24300);
and U37197 (N_37197,N_27603,N_20494);
nand U37198 (N_37198,N_24548,N_26061);
nand U37199 (N_37199,N_25058,N_29243);
xor U37200 (N_37200,N_25442,N_20010);
xor U37201 (N_37201,N_22598,N_28977);
nand U37202 (N_37202,N_29612,N_22993);
nand U37203 (N_37203,N_26111,N_21389);
nor U37204 (N_37204,N_21124,N_22064);
and U37205 (N_37205,N_29478,N_23949);
nor U37206 (N_37206,N_21977,N_22951);
nor U37207 (N_37207,N_22865,N_27192);
nand U37208 (N_37208,N_24301,N_22901);
nand U37209 (N_37209,N_28432,N_29169);
xor U37210 (N_37210,N_22233,N_24731);
xor U37211 (N_37211,N_20108,N_24872);
xor U37212 (N_37212,N_26142,N_21762);
or U37213 (N_37213,N_22075,N_28105);
nand U37214 (N_37214,N_23061,N_29664);
or U37215 (N_37215,N_25650,N_21611);
nor U37216 (N_37216,N_29365,N_28502);
nand U37217 (N_37217,N_27558,N_27649);
nand U37218 (N_37218,N_24366,N_20202);
nor U37219 (N_37219,N_22738,N_26158);
nor U37220 (N_37220,N_28208,N_29394);
and U37221 (N_37221,N_22724,N_27338);
nand U37222 (N_37222,N_28899,N_28179);
and U37223 (N_37223,N_23827,N_25008);
xnor U37224 (N_37224,N_29046,N_23550);
and U37225 (N_37225,N_27826,N_24735);
nor U37226 (N_37226,N_26916,N_27323);
nand U37227 (N_37227,N_26577,N_26237);
and U37228 (N_37228,N_24546,N_25221);
or U37229 (N_37229,N_25929,N_23671);
and U37230 (N_37230,N_23384,N_25248);
nand U37231 (N_37231,N_21055,N_20014);
and U37232 (N_37232,N_20130,N_23881);
nand U37233 (N_37233,N_20767,N_28575);
nand U37234 (N_37234,N_27331,N_21309);
or U37235 (N_37235,N_20212,N_27429);
nand U37236 (N_37236,N_23590,N_29018);
xnor U37237 (N_37237,N_26501,N_20791);
and U37238 (N_37238,N_22255,N_24566);
and U37239 (N_37239,N_28892,N_28330);
and U37240 (N_37240,N_21332,N_20007);
nand U37241 (N_37241,N_22048,N_28411);
nor U37242 (N_37242,N_26297,N_25711);
and U37243 (N_37243,N_27132,N_22227);
nand U37244 (N_37244,N_26421,N_21653);
and U37245 (N_37245,N_29246,N_28034);
nor U37246 (N_37246,N_27335,N_22485);
nand U37247 (N_37247,N_25521,N_25929);
xor U37248 (N_37248,N_27019,N_23696);
nor U37249 (N_37249,N_22810,N_23703);
and U37250 (N_37250,N_29474,N_25249);
nand U37251 (N_37251,N_27598,N_29172);
nand U37252 (N_37252,N_23320,N_24116);
nor U37253 (N_37253,N_27766,N_29112);
and U37254 (N_37254,N_20816,N_27994);
nor U37255 (N_37255,N_21341,N_21566);
nand U37256 (N_37256,N_25714,N_23552);
and U37257 (N_37257,N_20546,N_29981);
nand U37258 (N_37258,N_25925,N_29901);
and U37259 (N_37259,N_23291,N_27235);
and U37260 (N_37260,N_24650,N_21170);
xor U37261 (N_37261,N_23249,N_21619);
xnor U37262 (N_37262,N_27088,N_26905);
or U37263 (N_37263,N_29714,N_26107);
nor U37264 (N_37264,N_29852,N_22099);
nand U37265 (N_37265,N_24235,N_28185);
or U37266 (N_37266,N_25943,N_23297);
nor U37267 (N_37267,N_23374,N_23861);
nand U37268 (N_37268,N_25631,N_26700);
nand U37269 (N_37269,N_28943,N_28875);
xnor U37270 (N_37270,N_24221,N_28504);
and U37271 (N_37271,N_28261,N_28112);
xnor U37272 (N_37272,N_29297,N_20634);
or U37273 (N_37273,N_25953,N_26134);
and U37274 (N_37274,N_22199,N_26012);
nand U37275 (N_37275,N_20193,N_29852);
and U37276 (N_37276,N_25517,N_21075);
nor U37277 (N_37277,N_22371,N_26021);
and U37278 (N_37278,N_21128,N_27982);
nor U37279 (N_37279,N_27622,N_28593);
nand U37280 (N_37280,N_26506,N_25768);
xnor U37281 (N_37281,N_26148,N_28534);
nand U37282 (N_37282,N_24265,N_24089);
nand U37283 (N_37283,N_21133,N_28781);
xor U37284 (N_37284,N_28252,N_29564);
or U37285 (N_37285,N_27982,N_28837);
or U37286 (N_37286,N_22735,N_20444);
or U37287 (N_37287,N_28341,N_20943);
or U37288 (N_37288,N_27789,N_25400);
nand U37289 (N_37289,N_27862,N_20086);
and U37290 (N_37290,N_22386,N_20448);
and U37291 (N_37291,N_29088,N_25333);
or U37292 (N_37292,N_28256,N_27376);
nand U37293 (N_37293,N_20957,N_22259);
or U37294 (N_37294,N_22521,N_22281);
xnor U37295 (N_37295,N_24687,N_28919);
nor U37296 (N_37296,N_21048,N_27137);
xor U37297 (N_37297,N_23775,N_20943);
or U37298 (N_37298,N_26892,N_25092);
nand U37299 (N_37299,N_28616,N_28556);
nor U37300 (N_37300,N_23663,N_22654);
nand U37301 (N_37301,N_28823,N_25704);
or U37302 (N_37302,N_24240,N_20371);
and U37303 (N_37303,N_23665,N_27689);
nand U37304 (N_37304,N_29366,N_29562);
or U37305 (N_37305,N_28010,N_20186);
or U37306 (N_37306,N_24613,N_21709);
xnor U37307 (N_37307,N_24035,N_29795);
and U37308 (N_37308,N_29075,N_29930);
nand U37309 (N_37309,N_21000,N_21405);
or U37310 (N_37310,N_21924,N_27235);
nor U37311 (N_37311,N_26288,N_28699);
xnor U37312 (N_37312,N_26501,N_21440);
nor U37313 (N_37313,N_21228,N_21408);
nor U37314 (N_37314,N_26043,N_24206);
or U37315 (N_37315,N_21826,N_22983);
xor U37316 (N_37316,N_28041,N_27025);
nor U37317 (N_37317,N_22016,N_22945);
nor U37318 (N_37318,N_29406,N_25648);
nand U37319 (N_37319,N_23432,N_26291);
and U37320 (N_37320,N_29995,N_22935);
nand U37321 (N_37321,N_25936,N_21672);
xnor U37322 (N_37322,N_28505,N_24349);
xnor U37323 (N_37323,N_29746,N_22307);
nand U37324 (N_37324,N_24131,N_24615);
or U37325 (N_37325,N_24685,N_28892);
or U37326 (N_37326,N_25202,N_26612);
xor U37327 (N_37327,N_20317,N_23536);
nor U37328 (N_37328,N_23900,N_29653);
and U37329 (N_37329,N_27582,N_29473);
xor U37330 (N_37330,N_24375,N_22665);
and U37331 (N_37331,N_25667,N_28724);
nand U37332 (N_37332,N_28836,N_29300);
nor U37333 (N_37333,N_21532,N_20012);
and U37334 (N_37334,N_26965,N_23170);
nor U37335 (N_37335,N_27876,N_21395);
or U37336 (N_37336,N_23297,N_22978);
xor U37337 (N_37337,N_27147,N_20016);
nand U37338 (N_37338,N_25245,N_21927);
nor U37339 (N_37339,N_23729,N_22512);
nand U37340 (N_37340,N_24965,N_24924);
and U37341 (N_37341,N_25825,N_27401);
nand U37342 (N_37342,N_25554,N_28649);
xor U37343 (N_37343,N_20732,N_26205);
nor U37344 (N_37344,N_27086,N_20875);
nor U37345 (N_37345,N_22826,N_22337);
or U37346 (N_37346,N_24543,N_29331);
nor U37347 (N_37347,N_25997,N_29794);
or U37348 (N_37348,N_21618,N_23550);
xor U37349 (N_37349,N_22845,N_24510);
or U37350 (N_37350,N_29302,N_26210);
and U37351 (N_37351,N_21067,N_20795);
and U37352 (N_37352,N_23178,N_27822);
and U37353 (N_37353,N_24202,N_22913);
nor U37354 (N_37354,N_29593,N_29750);
or U37355 (N_37355,N_22215,N_28471);
or U37356 (N_37356,N_29159,N_27565);
nand U37357 (N_37357,N_20708,N_20283);
or U37358 (N_37358,N_29490,N_21705);
nor U37359 (N_37359,N_23758,N_26010);
nand U37360 (N_37360,N_28567,N_28538);
nor U37361 (N_37361,N_20687,N_24642);
and U37362 (N_37362,N_25415,N_24883);
nor U37363 (N_37363,N_29882,N_26923);
or U37364 (N_37364,N_28089,N_27847);
and U37365 (N_37365,N_28638,N_22483);
xor U37366 (N_37366,N_20299,N_23762);
and U37367 (N_37367,N_28133,N_20533);
nor U37368 (N_37368,N_21633,N_21238);
nand U37369 (N_37369,N_24591,N_23798);
xor U37370 (N_37370,N_28323,N_29918);
xnor U37371 (N_37371,N_21120,N_28842);
nand U37372 (N_37372,N_29278,N_23475);
nand U37373 (N_37373,N_20061,N_20503);
xor U37374 (N_37374,N_25001,N_21947);
or U37375 (N_37375,N_21719,N_21432);
xor U37376 (N_37376,N_28344,N_25801);
or U37377 (N_37377,N_26806,N_24977);
or U37378 (N_37378,N_24462,N_29826);
nor U37379 (N_37379,N_26846,N_27811);
nor U37380 (N_37380,N_24921,N_22179);
or U37381 (N_37381,N_27296,N_28279);
nand U37382 (N_37382,N_28817,N_24488);
xnor U37383 (N_37383,N_20093,N_20324);
nor U37384 (N_37384,N_20341,N_26212);
and U37385 (N_37385,N_21322,N_24745);
and U37386 (N_37386,N_21453,N_22371);
or U37387 (N_37387,N_27259,N_28093);
nor U37388 (N_37388,N_22942,N_21465);
or U37389 (N_37389,N_23388,N_24867);
xor U37390 (N_37390,N_24478,N_21338);
nor U37391 (N_37391,N_23455,N_23870);
or U37392 (N_37392,N_24983,N_27127);
and U37393 (N_37393,N_20510,N_21491);
or U37394 (N_37394,N_24052,N_25029);
and U37395 (N_37395,N_27568,N_22460);
and U37396 (N_37396,N_25180,N_24322);
xnor U37397 (N_37397,N_26285,N_23693);
nand U37398 (N_37398,N_27279,N_24048);
xnor U37399 (N_37399,N_22559,N_24300);
nand U37400 (N_37400,N_27169,N_26164);
or U37401 (N_37401,N_24574,N_26870);
xor U37402 (N_37402,N_28463,N_29565);
nand U37403 (N_37403,N_21834,N_21797);
or U37404 (N_37404,N_22322,N_21293);
and U37405 (N_37405,N_20556,N_22140);
nor U37406 (N_37406,N_29074,N_28003);
and U37407 (N_37407,N_23415,N_26847);
and U37408 (N_37408,N_29739,N_21610);
and U37409 (N_37409,N_26014,N_25428);
or U37410 (N_37410,N_24530,N_27366);
and U37411 (N_37411,N_27521,N_26902);
nor U37412 (N_37412,N_25842,N_29534);
nand U37413 (N_37413,N_29470,N_29294);
nor U37414 (N_37414,N_24358,N_26982);
nor U37415 (N_37415,N_27479,N_25989);
nand U37416 (N_37416,N_24755,N_25713);
and U37417 (N_37417,N_22486,N_26976);
or U37418 (N_37418,N_21473,N_26874);
or U37419 (N_37419,N_23477,N_27844);
nor U37420 (N_37420,N_24550,N_23006);
xnor U37421 (N_37421,N_20669,N_21341);
or U37422 (N_37422,N_28692,N_26908);
and U37423 (N_37423,N_29385,N_28559);
and U37424 (N_37424,N_28242,N_26771);
xnor U37425 (N_37425,N_20698,N_26488);
nor U37426 (N_37426,N_27597,N_23471);
xnor U37427 (N_37427,N_24973,N_20136);
xnor U37428 (N_37428,N_23519,N_29735);
nand U37429 (N_37429,N_26667,N_24948);
nand U37430 (N_37430,N_28911,N_29917);
nor U37431 (N_37431,N_28043,N_27063);
and U37432 (N_37432,N_28294,N_21116);
xor U37433 (N_37433,N_25337,N_29014);
nor U37434 (N_37434,N_20277,N_24539);
nor U37435 (N_37435,N_29187,N_28465);
xor U37436 (N_37436,N_24044,N_22388);
nor U37437 (N_37437,N_23168,N_23974);
xor U37438 (N_37438,N_24751,N_23293);
xnor U37439 (N_37439,N_28020,N_24031);
and U37440 (N_37440,N_25143,N_29394);
and U37441 (N_37441,N_25050,N_24401);
xor U37442 (N_37442,N_21326,N_22336);
nor U37443 (N_37443,N_26021,N_26103);
nor U37444 (N_37444,N_25257,N_20770);
or U37445 (N_37445,N_20486,N_29525);
nor U37446 (N_37446,N_20629,N_20675);
or U37447 (N_37447,N_24296,N_23167);
nor U37448 (N_37448,N_23926,N_24370);
or U37449 (N_37449,N_29427,N_23077);
nor U37450 (N_37450,N_21130,N_26792);
nor U37451 (N_37451,N_28827,N_20647);
or U37452 (N_37452,N_26740,N_23789);
nand U37453 (N_37453,N_27685,N_27272);
nand U37454 (N_37454,N_24824,N_26493);
and U37455 (N_37455,N_29460,N_20484);
nor U37456 (N_37456,N_23386,N_24550);
xor U37457 (N_37457,N_24816,N_29439);
or U37458 (N_37458,N_26520,N_24145);
nor U37459 (N_37459,N_28495,N_29120);
and U37460 (N_37460,N_28885,N_24949);
and U37461 (N_37461,N_22321,N_25546);
xnor U37462 (N_37462,N_21501,N_27799);
or U37463 (N_37463,N_25032,N_25787);
or U37464 (N_37464,N_27695,N_27393);
nor U37465 (N_37465,N_26370,N_26201);
or U37466 (N_37466,N_27830,N_25523);
and U37467 (N_37467,N_20136,N_27490);
nor U37468 (N_37468,N_27037,N_28644);
nor U37469 (N_37469,N_21638,N_27832);
xnor U37470 (N_37470,N_21725,N_25384);
and U37471 (N_37471,N_24482,N_24578);
xor U37472 (N_37472,N_26986,N_21103);
nand U37473 (N_37473,N_21991,N_22908);
nand U37474 (N_37474,N_24824,N_25917);
and U37475 (N_37475,N_27835,N_24164);
nand U37476 (N_37476,N_20883,N_27266);
or U37477 (N_37477,N_29000,N_26334);
xor U37478 (N_37478,N_29717,N_21790);
nand U37479 (N_37479,N_20122,N_27158);
nor U37480 (N_37480,N_27822,N_23768);
or U37481 (N_37481,N_22556,N_23336);
and U37482 (N_37482,N_28368,N_21806);
nor U37483 (N_37483,N_24111,N_28264);
nand U37484 (N_37484,N_27446,N_21224);
nor U37485 (N_37485,N_28646,N_26761);
or U37486 (N_37486,N_29809,N_29253);
and U37487 (N_37487,N_21725,N_27206);
or U37488 (N_37488,N_27486,N_21877);
xor U37489 (N_37489,N_24808,N_23312);
and U37490 (N_37490,N_28633,N_25165);
and U37491 (N_37491,N_23330,N_28032);
nand U37492 (N_37492,N_21562,N_23688);
nand U37493 (N_37493,N_25892,N_29871);
or U37494 (N_37494,N_24746,N_20397);
xnor U37495 (N_37495,N_25410,N_25254);
nor U37496 (N_37496,N_23977,N_21881);
and U37497 (N_37497,N_24991,N_28795);
nand U37498 (N_37498,N_23748,N_20199);
xnor U37499 (N_37499,N_21117,N_25799);
nor U37500 (N_37500,N_22031,N_23675);
xnor U37501 (N_37501,N_28887,N_20881);
nor U37502 (N_37502,N_28026,N_28023);
nor U37503 (N_37503,N_22740,N_28225);
or U37504 (N_37504,N_25512,N_21295);
nor U37505 (N_37505,N_20172,N_29118);
xnor U37506 (N_37506,N_20031,N_28349);
xor U37507 (N_37507,N_25875,N_21863);
and U37508 (N_37508,N_25224,N_26471);
or U37509 (N_37509,N_29498,N_27994);
or U37510 (N_37510,N_21857,N_25350);
xnor U37511 (N_37511,N_22803,N_21461);
or U37512 (N_37512,N_26994,N_24885);
and U37513 (N_37513,N_27698,N_29087);
or U37514 (N_37514,N_21253,N_29457);
or U37515 (N_37515,N_29958,N_22766);
nor U37516 (N_37516,N_23436,N_24771);
nand U37517 (N_37517,N_25613,N_24751);
or U37518 (N_37518,N_21371,N_24153);
or U37519 (N_37519,N_29795,N_21391);
and U37520 (N_37520,N_22176,N_29928);
nor U37521 (N_37521,N_27506,N_22261);
nor U37522 (N_37522,N_25018,N_25506);
nand U37523 (N_37523,N_22573,N_29078);
and U37524 (N_37524,N_23206,N_24568);
nor U37525 (N_37525,N_27838,N_26178);
nand U37526 (N_37526,N_20065,N_27753);
nor U37527 (N_37527,N_25977,N_25587);
or U37528 (N_37528,N_24049,N_22459);
nor U37529 (N_37529,N_29774,N_28063);
xnor U37530 (N_37530,N_25965,N_20948);
nand U37531 (N_37531,N_20798,N_26518);
or U37532 (N_37532,N_27496,N_27728);
and U37533 (N_37533,N_27771,N_25185);
nand U37534 (N_37534,N_24069,N_22817);
nor U37535 (N_37535,N_29455,N_21649);
xor U37536 (N_37536,N_22979,N_23867);
nor U37537 (N_37537,N_22850,N_22551);
xnor U37538 (N_37538,N_25459,N_29074);
nor U37539 (N_37539,N_23925,N_29115);
nand U37540 (N_37540,N_21141,N_28219);
or U37541 (N_37541,N_25517,N_23664);
or U37542 (N_37542,N_20767,N_20456);
and U37543 (N_37543,N_23285,N_29896);
and U37544 (N_37544,N_27337,N_24685);
nand U37545 (N_37545,N_27743,N_25000);
xnor U37546 (N_37546,N_28610,N_25431);
nor U37547 (N_37547,N_21847,N_25628);
nor U37548 (N_37548,N_28140,N_27350);
xor U37549 (N_37549,N_26997,N_23396);
xnor U37550 (N_37550,N_22023,N_20167);
nand U37551 (N_37551,N_23073,N_29330);
nand U37552 (N_37552,N_27004,N_21532);
nand U37553 (N_37553,N_28051,N_27175);
nor U37554 (N_37554,N_28728,N_28939);
xor U37555 (N_37555,N_23117,N_21805);
and U37556 (N_37556,N_23696,N_28190);
and U37557 (N_37557,N_25427,N_21673);
or U37558 (N_37558,N_25202,N_22963);
or U37559 (N_37559,N_20092,N_24178);
or U37560 (N_37560,N_23718,N_26525);
xnor U37561 (N_37561,N_22272,N_22577);
or U37562 (N_37562,N_26152,N_29175);
and U37563 (N_37563,N_27593,N_20883);
and U37564 (N_37564,N_21814,N_27704);
nand U37565 (N_37565,N_23113,N_25648);
or U37566 (N_37566,N_26515,N_27444);
nor U37567 (N_37567,N_25526,N_20397);
nand U37568 (N_37568,N_25184,N_26152);
nand U37569 (N_37569,N_29353,N_26601);
nand U37570 (N_37570,N_26912,N_21837);
nand U37571 (N_37571,N_29122,N_24018);
nor U37572 (N_37572,N_29525,N_20039);
nand U37573 (N_37573,N_25174,N_25344);
xor U37574 (N_37574,N_23763,N_29535);
nand U37575 (N_37575,N_24236,N_24283);
nand U37576 (N_37576,N_24446,N_29380);
nor U37577 (N_37577,N_21401,N_22786);
xnor U37578 (N_37578,N_21016,N_25165);
or U37579 (N_37579,N_23022,N_23249);
nor U37580 (N_37580,N_23714,N_24831);
nand U37581 (N_37581,N_23616,N_29064);
or U37582 (N_37582,N_24943,N_23613);
xnor U37583 (N_37583,N_28938,N_22421);
nand U37584 (N_37584,N_20060,N_22446);
or U37585 (N_37585,N_21656,N_23080);
and U37586 (N_37586,N_20684,N_29205);
nand U37587 (N_37587,N_25297,N_26013);
xnor U37588 (N_37588,N_28895,N_23412);
and U37589 (N_37589,N_29562,N_20333);
nand U37590 (N_37590,N_28027,N_21490);
or U37591 (N_37591,N_28254,N_27343);
nand U37592 (N_37592,N_25197,N_20438);
and U37593 (N_37593,N_24798,N_20850);
xnor U37594 (N_37594,N_26315,N_20865);
nor U37595 (N_37595,N_23254,N_20082);
nand U37596 (N_37596,N_25807,N_25333);
and U37597 (N_37597,N_22750,N_22538);
xor U37598 (N_37598,N_22844,N_24315);
xnor U37599 (N_37599,N_24044,N_27922);
nor U37600 (N_37600,N_20610,N_26442);
xor U37601 (N_37601,N_27087,N_21649);
or U37602 (N_37602,N_29002,N_20281);
nand U37603 (N_37603,N_25971,N_20017);
xor U37604 (N_37604,N_29851,N_23456);
or U37605 (N_37605,N_26004,N_28260);
nor U37606 (N_37606,N_28036,N_28976);
or U37607 (N_37607,N_25386,N_22939);
or U37608 (N_37608,N_22139,N_22333);
nor U37609 (N_37609,N_22870,N_28995);
nand U37610 (N_37610,N_24226,N_24002);
nand U37611 (N_37611,N_22234,N_22745);
nand U37612 (N_37612,N_27428,N_20765);
or U37613 (N_37613,N_22507,N_22733);
and U37614 (N_37614,N_28514,N_24474);
xnor U37615 (N_37615,N_21614,N_21932);
nor U37616 (N_37616,N_27445,N_20457);
nor U37617 (N_37617,N_23261,N_22842);
and U37618 (N_37618,N_21016,N_25062);
and U37619 (N_37619,N_28323,N_23111);
xnor U37620 (N_37620,N_28468,N_25005);
or U37621 (N_37621,N_27601,N_25059);
nor U37622 (N_37622,N_23101,N_25111);
nor U37623 (N_37623,N_20038,N_24692);
nand U37624 (N_37624,N_29602,N_20903);
nand U37625 (N_37625,N_26779,N_26459);
nor U37626 (N_37626,N_28278,N_28089);
and U37627 (N_37627,N_22074,N_21652);
and U37628 (N_37628,N_22695,N_23764);
nor U37629 (N_37629,N_25868,N_22544);
or U37630 (N_37630,N_25416,N_28553);
xnor U37631 (N_37631,N_26500,N_29654);
nand U37632 (N_37632,N_28718,N_20977);
nor U37633 (N_37633,N_27893,N_20052);
and U37634 (N_37634,N_25718,N_28620);
nor U37635 (N_37635,N_21491,N_23679);
and U37636 (N_37636,N_26099,N_29251);
nor U37637 (N_37637,N_23785,N_26730);
and U37638 (N_37638,N_27135,N_23949);
nor U37639 (N_37639,N_24289,N_24377);
nor U37640 (N_37640,N_26044,N_20629);
nand U37641 (N_37641,N_23674,N_21282);
and U37642 (N_37642,N_28738,N_27096);
nand U37643 (N_37643,N_23693,N_20707);
and U37644 (N_37644,N_21411,N_21577);
xor U37645 (N_37645,N_28034,N_27279);
xor U37646 (N_37646,N_28493,N_26419);
nor U37647 (N_37647,N_20178,N_20869);
nand U37648 (N_37648,N_26965,N_23395);
nand U37649 (N_37649,N_25923,N_24352);
or U37650 (N_37650,N_26632,N_24591);
and U37651 (N_37651,N_20500,N_28882);
xor U37652 (N_37652,N_24836,N_28811);
or U37653 (N_37653,N_23964,N_26189);
nand U37654 (N_37654,N_25640,N_22494);
nand U37655 (N_37655,N_25249,N_23323);
xor U37656 (N_37656,N_22729,N_29694);
xnor U37657 (N_37657,N_28511,N_20658);
and U37658 (N_37658,N_24765,N_20537);
and U37659 (N_37659,N_21477,N_29611);
nand U37660 (N_37660,N_27287,N_28487);
xor U37661 (N_37661,N_27638,N_20436);
or U37662 (N_37662,N_25577,N_25399);
and U37663 (N_37663,N_28817,N_21150);
nor U37664 (N_37664,N_23249,N_24852);
and U37665 (N_37665,N_23562,N_25599);
nor U37666 (N_37666,N_27411,N_29474);
nor U37667 (N_37667,N_29811,N_23357);
or U37668 (N_37668,N_28232,N_25775);
and U37669 (N_37669,N_27066,N_26294);
nand U37670 (N_37670,N_23057,N_21618);
nor U37671 (N_37671,N_23493,N_29561);
xor U37672 (N_37672,N_21078,N_24132);
or U37673 (N_37673,N_22857,N_29168);
nand U37674 (N_37674,N_20691,N_25850);
nor U37675 (N_37675,N_25107,N_24032);
or U37676 (N_37676,N_22043,N_26203);
or U37677 (N_37677,N_21909,N_25649);
nand U37678 (N_37678,N_22343,N_22031);
nor U37679 (N_37679,N_25268,N_25808);
xor U37680 (N_37680,N_22947,N_28745);
or U37681 (N_37681,N_24354,N_21704);
xor U37682 (N_37682,N_20898,N_29439);
nand U37683 (N_37683,N_27931,N_23361);
or U37684 (N_37684,N_28324,N_25310);
xnor U37685 (N_37685,N_22792,N_29838);
xnor U37686 (N_37686,N_24796,N_28768);
nor U37687 (N_37687,N_20993,N_29936);
nor U37688 (N_37688,N_27179,N_23548);
and U37689 (N_37689,N_24142,N_27604);
or U37690 (N_37690,N_25243,N_24963);
xnor U37691 (N_37691,N_25260,N_27665);
nand U37692 (N_37692,N_24876,N_28463);
nor U37693 (N_37693,N_28434,N_28518);
and U37694 (N_37694,N_20179,N_22343);
xnor U37695 (N_37695,N_24598,N_23733);
nand U37696 (N_37696,N_27005,N_23846);
nand U37697 (N_37697,N_25260,N_28296);
nand U37698 (N_37698,N_23237,N_29833);
or U37699 (N_37699,N_28466,N_28620);
and U37700 (N_37700,N_28099,N_28390);
xnor U37701 (N_37701,N_22730,N_26892);
xor U37702 (N_37702,N_26155,N_27135);
xnor U37703 (N_37703,N_20479,N_25683);
or U37704 (N_37704,N_26589,N_20587);
or U37705 (N_37705,N_20080,N_20200);
or U37706 (N_37706,N_28929,N_21505);
or U37707 (N_37707,N_21603,N_29832);
nand U37708 (N_37708,N_26020,N_28545);
nand U37709 (N_37709,N_20689,N_26756);
and U37710 (N_37710,N_21157,N_23202);
or U37711 (N_37711,N_20821,N_22717);
nor U37712 (N_37712,N_28188,N_27281);
nor U37713 (N_37713,N_25283,N_22305);
xnor U37714 (N_37714,N_20509,N_27938);
xnor U37715 (N_37715,N_24745,N_24085);
nor U37716 (N_37716,N_21379,N_27446);
nand U37717 (N_37717,N_24575,N_21599);
nor U37718 (N_37718,N_25827,N_24666);
nand U37719 (N_37719,N_29781,N_20411);
or U37720 (N_37720,N_20754,N_23737);
nand U37721 (N_37721,N_21045,N_25942);
or U37722 (N_37722,N_28535,N_21126);
nand U37723 (N_37723,N_25801,N_27998);
or U37724 (N_37724,N_28308,N_27284);
xnor U37725 (N_37725,N_29502,N_25463);
or U37726 (N_37726,N_21138,N_25381);
nor U37727 (N_37727,N_21214,N_24519);
nor U37728 (N_37728,N_21214,N_28768);
or U37729 (N_37729,N_25972,N_22867);
nor U37730 (N_37730,N_21729,N_22903);
and U37731 (N_37731,N_27487,N_25097);
nor U37732 (N_37732,N_25383,N_21804);
xor U37733 (N_37733,N_28454,N_26166);
and U37734 (N_37734,N_25554,N_27834);
nand U37735 (N_37735,N_29759,N_28614);
and U37736 (N_37736,N_27304,N_20077);
xnor U37737 (N_37737,N_23209,N_22658);
xor U37738 (N_37738,N_23050,N_29230);
xor U37739 (N_37739,N_24127,N_25320);
or U37740 (N_37740,N_27749,N_21877);
nand U37741 (N_37741,N_23909,N_24516);
xor U37742 (N_37742,N_24165,N_24461);
nand U37743 (N_37743,N_28592,N_24709);
nor U37744 (N_37744,N_26512,N_27864);
or U37745 (N_37745,N_20579,N_27379);
nand U37746 (N_37746,N_25406,N_25207);
xnor U37747 (N_37747,N_20481,N_20641);
xnor U37748 (N_37748,N_28254,N_29284);
xor U37749 (N_37749,N_29334,N_26775);
and U37750 (N_37750,N_26794,N_26048);
nor U37751 (N_37751,N_24267,N_24815);
nor U37752 (N_37752,N_29267,N_28327);
and U37753 (N_37753,N_20507,N_20806);
xor U37754 (N_37754,N_27995,N_26190);
and U37755 (N_37755,N_24580,N_27276);
nand U37756 (N_37756,N_22710,N_25368);
nor U37757 (N_37757,N_22879,N_20011);
or U37758 (N_37758,N_22536,N_28118);
nand U37759 (N_37759,N_29586,N_26880);
nor U37760 (N_37760,N_21586,N_28722);
nor U37761 (N_37761,N_21665,N_24997);
xnor U37762 (N_37762,N_21578,N_25380);
and U37763 (N_37763,N_25028,N_27586);
xor U37764 (N_37764,N_28698,N_21415);
nor U37765 (N_37765,N_29601,N_20230);
xor U37766 (N_37766,N_24324,N_24711);
or U37767 (N_37767,N_27590,N_20027);
or U37768 (N_37768,N_25969,N_22389);
and U37769 (N_37769,N_22210,N_20499);
nor U37770 (N_37770,N_24091,N_22172);
nor U37771 (N_37771,N_21892,N_25876);
or U37772 (N_37772,N_26795,N_20375);
nand U37773 (N_37773,N_24762,N_26101);
xor U37774 (N_37774,N_26986,N_27699);
nor U37775 (N_37775,N_23746,N_29231);
nor U37776 (N_37776,N_22086,N_26300);
and U37777 (N_37777,N_29226,N_25069);
and U37778 (N_37778,N_25154,N_29460);
and U37779 (N_37779,N_27808,N_21363);
xor U37780 (N_37780,N_22392,N_29669);
nor U37781 (N_37781,N_29176,N_23768);
or U37782 (N_37782,N_21932,N_28809);
nand U37783 (N_37783,N_21410,N_20921);
or U37784 (N_37784,N_25679,N_29012);
xnor U37785 (N_37785,N_24083,N_28501);
nand U37786 (N_37786,N_23483,N_25552);
nor U37787 (N_37787,N_22319,N_22955);
or U37788 (N_37788,N_22541,N_27370);
and U37789 (N_37789,N_23481,N_23587);
or U37790 (N_37790,N_22829,N_20268);
nor U37791 (N_37791,N_25814,N_27931);
nor U37792 (N_37792,N_21811,N_20035);
or U37793 (N_37793,N_24389,N_20075);
xnor U37794 (N_37794,N_26449,N_21931);
xor U37795 (N_37795,N_24710,N_27927);
or U37796 (N_37796,N_27399,N_23253);
or U37797 (N_37797,N_28704,N_23956);
xor U37798 (N_37798,N_29930,N_24105);
nor U37799 (N_37799,N_25272,N_21447);
nor U37800 (N_37800,N_23343,N_24131);
xor U37801 (N_37801,N_26369,N_29440);
and U37802 (N_37802,N_27580,N_23828);
nand U37803 (N_37803,N_25936,N_20454);
and U37804 (N_37804,N_27496,N_23047);
and U37805 (N_37805,N_27207,N_25659);
nor U37806 (N_37806,N_21296,N_23201);
or U37807 (N_37807,N_21980,N_23641);
or U37808 (N_37808,N_24517,N_20111);
and U37809 (N_37809,N_25817,N_27204);
xnor U37810 (N_37810,N_26898,N_24824);
nand U37811 (N_37811,N_22244,N_25077);
nand U37812 (N_37812,N_20588,N_24924);
or U37813 (N_37813,N_21597,N_24468);
nor U37814 (N_37814,N_23451,N_29364);
xor U37815 (N_37815,N_26187,N_29858);
nand U37816 (N_37816,N_26419,N_26259);
and U37817 (N_37817,N_25659,N_21763);
or U37818 (N_37818,N_27880,N_28213);
xor U37819 (N_37819,N_20839,N_23413);
nand U37820 (N_37820,N_29944,N_26229);
and U37821 (N_37821,N_26959,N_29530);
nor U37822 (N_37822,N_24474,N_24021);
nand U37823 (N_37823,N_22853,N_29730);
and U37824 (N_37824,N_24395,N_24534);
xor U37825 (N_37825,N_22825,N_28027);
nand U37826 (N_37826,N_26568,N_25014);
nand U37827 (N_37827,N_25068,N_22364);
nor U37828 (N_37828,N_25262,N_22155);
xor U37829 (N_37829,N_21502,N_22292);
nor U37830 (N_37830,N_23224,N_22407);
nand U37831 (N_37831,N_28609,N_29940);
or U37832 (N_37832,N_23099,N_26665);
or U37833 (N_37833,N_23210,N_23939);
and U37834 (N_37834,N_23613,N_26733);
nand U37835 (N_37835,N_26100,N_24647);
nor U37836 (N_37836,N_21766,N_24788);
xnor U37837 (N_37837,N_22211,N_21468);
nor U37838 (N_37838,N_22922,N_25184);
nor U37839 (N_37839,N_27800,N_29285);
xor U37840 (N_37840,N_21918,N_23883);
or U37841 (N_37841,N_25076,N_25768);
xnor U37842 (N_37842,N_21853,N_25888);
and U37843 (N_37843,N_23516,N_27379);
and U37844 (N_37844,N_26256,N_29562);
nor U37845 (N_37845,N_22522,N_29904);
xor U37846 (N_37846,N_24045,N_29884);
or U37847 (N_37847,N_22522,N_22278);
nor U37848 (N_37848,N_23821,N_22450);
nor U37849 (N_37849,N_24430,N_29498);
and U37850 (N_37850,N_24153,N_24065);
nor U37851 (N_37851,N_24537,N_23848);
xnor U37852 (N_37852,N_28906,N_24752);
xor U37853 (N_37853,N_26864,N_25680);
and U37854 (N_37854,N_23176,N_21274);
or U37855 (N_37855,N_29183,N_24475);
or U37856 (N_37856,N_26994,N_29455);
and U37857 (N_37857,N_20141,N_23889);
nor U37858 (N_37858,N_24380,N_26238);
or U37859 (N_37859,N_20016,N_25700);
nand U37860 (N_37860,N_24815,N_28747);
and U37861 (N_37861,N_21717,N_22020);
and U37862 (N_37862,N_26584,N_27882);
or U37863 (N_37863,N_23676,N_29498);
nand U37864 (N_37864,N_20483,N_20039);
nand U37865 (N_37865,N_28326,N_29649);
nor U37866 (N_37866,N_25374,N_28322);
nand U37867 (N_37867,N_28360,N_29742);
and U37868 (N_37868,N_29932,N_28174);
nand U37869 (N_37869,N_21474,N_20136);
nand U37870 (N_37870,N_22069,N_21889);
nand U37871 (N_37871,N_25898,N_25281);
and U37872 (N_37872,N_29286,N_26698);
nand U37873 (N_37873,N_27795,N_29134);
or U37874 (N_37874,N_29055,N_28898);
or U37875 (N_37875,N_26927,N_21430);
nor U37876 (N_37876,N_21112,N_26682);
xnor U37877 (N_37877,N_24930,N_23963);
or U37878 (N_37878,N_26937,N_20437);
nand U37879 (N_37879,N_20457,N_23620);
nor U37880 (N_37880,N_25878,N_21747);
nand U37881 (N_37881,N_29477,N_29175);
nand U37882 (N_37882,N_22294,N_26811);
and U37883 (N_37883,N_22276,N_25433);
nand U37884 (N_37884,N_29196,N_24815);
nor U37885 (N_37885,N_26483,N_22965);
nand U37886 (N_37886,N_23782,N_29197);
nor U37887 (N_37887,N_21158,N_27105);
and U37888 (N_37888,N_27287,N_26627);
nand U37889 (N_37889,N_21135,N_23010);
nand U37890 (N_37890,N_22190,N_23729);
xor U37891 (N_37891,N_29042,N_28642);
nand U37892 (N_37892,N_29419,N_20272);
nand U37893 (N_37893,N_26751,N_24895);
nor U37894 (N_37894,N_22014,N_24214);
and U37895 (N_37895,N_28149,N_29992);
or U37896 (N_37896,N_22225,N_27910);
xor U37897 (N_37897,N_25074,N_28552);
and U37898 (N_37898,N_29509,N_21333);
nor U37899 (N_37899,N_29800,N_20695);
or U37900 (N_37900,N_27877,N_28467);
nor U37901 (N_37901,N_21899,N_27109);
and U37902 (N_37902,N_23762,N_29392);
nand U37903 (N_37903,N_26093,N_24348);
nand U37904 (N_37904,N_23103,N_29654);
or U37905 (N_37905,N_24686,N_21851);
nor U37906 (N_37906,N_27597,N_20651);
and U37907 (N_37907,N_22199,N_23987);
xor U37908 (N_37908,N_27876,N_26960);
nor U37909 (N_37909,N_29851,N_23965);
or U37910 (N_37910,N_23843,N_24780);
nor U37911 (N_37911,N_23768,N_27336);
and U37912 (N_37912,N_20425,N_20029);
and U37913 (N_37913,N_23069,N_22302);
and U37914 (N_37914,N_21468,N_28203);
and U37915 (N_37915,N_27224,N_25703);
nor U37916 (N_37916,N_21800,N_21882);
nand U37917 (N_37917,N_20669,N_27998);
xor U37918 (N_37918,N_23196,N_21393);
nor U37919 (N_37919,N_21734,N_28294);
xor U37920 (N_37920,N_25355,N_21891);
and U37921 (N_37921,N_28226,N_25291);
and U37922 (N_37922,N_23605,N_29864);
and U37923 (N_37923,N_21036,N_20927);
nor U37924 (N_37924,N_22364,N_21756);
or U37925 (N_37925,N_28475,N_24761);
nand U37926 (N_37926,N_27758,N_23209);
xnor U37927 (N_37927,N_24306,N_26064);
nand U37928 (N_37928,N_26285,N_24762);
and U37929 (N_37929,N_23786,N_22325);
xor U37930 (N_37930,N_22383,N_24343);
and U37931 (N_37931,N_27176,N_23789);
or U37932 (N_37932,N_28031,N_28570);
nor U37933 (N_37933,N_24758,N_21154);
and U37934 (N_37934,N_24412,N_26469);
nand U37935 (N_37935,N_29042,N_22817);
xor U37936 (N_37936,N_23801,N_20656);
nor U37937 (N_37937,N_24788,N_27572);
or U37938 (N_37938,N_22210,N_25235);
nor U37939 (N_37939,N_23879,N_26754);
xor U37940 (N_37940,N_23918,N_21034);
xnor U37941 (N_37941,N_26883,N_27002);
xnor U37942 (N_37942,N_26834,N_29509);
nand U37943 (N_37943,N_27665,N_21205);
or U37944 (N_37944,N_20052,N_28436);
xor U37945 (N_37945,N_28140,N_20319);
and U37946 (N_37946,N_22983,N_23023);
nor U37947 (N_37947,N_24415,N_28022);
or U37948 (N_37948,N_25797,N_23883);
nor U37949 (N_37949,N_26151,N_21483);
nor U37950 (N_37950,N_28967,N_26546);
xnor U37951 (N_37951,N_27611,N_23135);
nand U37952 (N_37952,N_24629,N_23532);
xor U37953 (N_37953,N_26036,N_27537);
nand U37954 (N_37954,N_28794,N_22535);
and U37955 (N_37955,N_28269,N_24890);
nor U37956 (N_37956,N_21574,N_20150);
or U37957 (N_37957,N_20153,N_20487);
and U37958 (N_37958,N_25689,N_25308);
xnor U37959 (N_37959,N_28613,N_22356);
or U37960 (N_37960,N_28724,N_26421);
xnor U37961 (N_37961,N_23101,N_22276);
xor U37962 (N_37962,N_27334,N_22053);
xnor U37963 (N_37963,N_27911,N_21001);
nor U37964 (N_37964,N_24390,N_26208);
or U37965 (N_37965,N_26287,N_20825);
or U37966 (N_37966,N_27212,N_21644);
nand U37967 (N_37967,N_25086,N_23966);
nor U37968 (N_37968,N_21049,N_21862);
nand U37969 (N_37969,N_24226,N_26489);
or U37970 (N_37970,N_28948,N_20197);
nor U37971 (N_37971,N_23114,N_29478);
and U37972 (N_37972,N_27677,N_20970);
or U37973 (N_37973,N_20517,N_29704);
nand U37974 (N_37974,N_23332,N_21533);
xnor U37975 (N_37975,N_27479,N_24462);
nor U37976 (N_37976,N_24051,N_22637);
nor U37977 (N_37977,N_23871,N_28553);
nand U37978 (N_37978,N_26874,N_28970);
xor U37979 (N_37979,N_26604,N_24101);
and U37980 (N_37980,N_28708,N_24595);
nand U37981 (N_37981,N_28341,N_21739);
nor U37982 (N_37982,N_24146,N_20086);
or U37983 (N_37983,N_29496,N_21640);
nor U37984 (N_37984,N_28260,N_25922);
or U37985 (N_37985,N_20272,N_29823);
nor U37986 (N_37986,N_22021,N_20719);
xor U37987 (N_37987,N_26828,N_21772);
nand U37988 (N_37988,N_25613,N_24359);
nand U37989 (N_37989,N_29682,N_20536);
nand U37990 (N_37990,N_29353,N_22430);
nor U37991 (N_37991,N_23949,N_26141);
and U37992 (N_37992,N_27496,N_25689);
and U37993 (N_37993,N_23480,N_24844);
and U37994 (N_37994,N_22612,N_25359);
and U37995 (N_37995,N_22615,N_20970);
or U37996 (N_37996,N_22882,N_24051);
and U37997 (N_37997,N_20810,N_20350);
or U37998 (N_37998,N_24945,N_24027);
nand U37999 (N_37999,N_23044,N_29085);
nor U38000 (N_38000,N_27939,N_20752);
nand U38001 (N_38001,N_24863,N_29796);
or U38002 (N_38002,N_28228,N_29882);
xnor U38003 (N_38003,N_27134,N_24884);
and U38004 (N_38004,N_28705,N_22292);
nor U38005 (N_38005,N_28063,N_24168);
or U38006 (N_38006,N_24547,N_22718);
nand U38007 (N_38007,N_22125,N_26606);
and U38008 (N_38008,N_23022,N_20288);
and U38009 (N_38009,N_22923,N_26855);
and U38010 (N_38010,N_24974,N_29358);
or U38011 (N_38011,N_26723,N_24161);
nand U38012 (N_38012,N_20635,N_21684);
or U38013 (N_38013,N_25750,N_23865);
nor U38014 (N_38014,N_27687,N_23961);
nor U38015 (N_38015,N_27797,N_25373);
nor U38016 (N_38016,N_28432,N_20167);
nor U38017 (N_38017,N_23300,N_26050);
or U38018 (N_38018,N_27741,N_26248);
nand U38019 (N_38019,N_27294,N_25781);
nand U38020 (N_38020,N_22874,N_29268);
xnor U38021 (N_38021,N_29837,N_26065);
xnor U38022 (N_38022,N_21191,N_21538);
nand U38023 (N_38023,N_23332,N_29339);
and U38024 (N_38024,N_21380,N_27301);
or U38025 (N_38025,N_21407,N_24952);
nor U38026 (N_38026,N_25041,N_22456);
and U38027 (N_38027,N_22692,N_26756);
xor U38028 (N_38028,N_20203,N_21828);
and U38029 (N_38029,N_26221,N_25773);
nand U38030 (N_38030,N_26648,N_22089);
nor U38031 (N_38031,N_27615,N_22567);
and U38032 (N_38032,N_21081,N_26552);
or U38033 (N_38033,N_28261,N_23200);
nand U38034 (N_38034,N_20840,N_26975);
xnor U38035 (N_38035,N_22843,N_29723);
and U38036 (N_38036,N_24232,N_28862);
nor U38037 (N_38037,N_25578,N_28992);
nand U38038 (N_38038,N_26112,N_23268);
or U38039 (N_38039,N_26121,N_24366);
or U38040 (N_38040,N_24937,N_29450);
and U38041 (N_38041,N_20791,N_22461);
xnor U38042 (N_38042,N_23939,N_21962);
nand U38043 (N_38043,N_21996,N_29614);
and U38044 (N_38044,N_26213,N_27063);
nand U38045 (N_38045,N_24744,N_20954);
xor U38046 (N_38046,N_24141,N_22950);
nor U38047 (N_38047,N_23660,N_21137);
nand U38048 (N_38048,N_23009,N_20793);
xor U38049 (N_38049,N_25504,N_25424);
xnor U38050 (N_38050,N_23916,N_27143);
and U38051 (N_38051,N_21288,N_28389);
xnor U38052 (N_38052,N_28338,N_20136);
nand U38053 (N_38053,N_28050,N_26268);
nand U38054 (N_38054,N_28598,N_20888);
and U38055 (N_38055,N_29761,N_22777);
and U38056 (N_38056,N_20814,N_27176);
or U38057 (N_38057,N_25362,N_27054);
nand U38058 (N_38058,N_23773,N_24557);
nand U38059 (N_38059,N_23420,N_29957);
nor U38060 (N_38060,N_22309,N_22542);
nor U38061 (N_38061,N_20695,N_22703);
nand U38062 (N_38062,N_20869,N_22886);
and U38063 (N_38063,N_24463,N_21392);
nor U38064 (N_38064,N_23102,N_28859);
or U38065 (N_38065,N_22973,N_28657);
nand U38066 (N_38066,N_27472,N_22514);
xnor U38067 (N_38067,N_22550,N_21997);
and U38068 (N_38068,N_25379,N_24747);
or U38069 (N_38069,N_28320,N_20169);
nor U38070 (N_38070,N_28507,N_22044);
and U38071 (N_38071,N_23914,N_20224);
or U38072 (N_38072,N_25331,N_21923);
or U38073 (N_38073,N_21897,N_22629);
xor U38074 (N_38074,N_20394,N_28508);
or U38075 (N_38075,N_23895,N_26661);
xor U38076 (N_38076,N_29868,N_24538);
nand U38077 (N_38077,N_23098,N_23837);
xnor U38078 (N_38078,N_27407,N_26311);
or U38079 (N_38079,N_22714,N_20352);
or U38080 (N_38080,N_26651,N_25874);
nor U38081 (N_38081,N_25083,N_24898);
and U38082 (N_38082,N_28113,N_29606);
and U38083 (N_38083,N_23751,N_24364);
and U38084 (N_38084,N_29238,N_25282);
nand U38085 (N_38085,N_28552,N_27151);
or U38086 (N_38086,N_21948,N_26756);
nor U38087 (N_38087,N_20387,N_28611);
nand U38088 (N_38088,N_24811,N_20552);
and U38089 (N_38089,N_23802,N_27321);
or U38090 (N_38090,N_20888,N_29657);
and U38091 (N_38091,N_28207,N_26103);
or U38092 (N_38092,N_26169,N_22437);
nand U38093 (N_38093,N_23842,N_21194);
and U38094 (N_38094,N_21642,N_27486);
or U38095 (N_38095,N_20833,N_27025);
nand U38096 (N_38096,N_28493,N_26274);
nor U38097 (N_38097,N_27339,N_25848);
and U38098 (N_38098,N_26799,N_25600);
xnor U38099 (N_38099,N_28587,N_21526);
xor U38100 (N_38100,N_24671,N_28858);
or U38101 (N_38101,N_24683,N_29463);
nand U38102 (N_38102,N_21195,N_21377);
or U38103 (N_38103,N_24701,N_20696);
nor U38104 (N_38104,N_25205,N_23248);
nand U38105 (N_38105,N_20772,N_26596);
xnor U38106 (N_38106,N_26389,N_23662);
nand U38107 (N_38107,N_20173,N_26928);
nand U38108 (N_38108,N_21830,N_28812);
nor U38109 (N_38109,N_28496,N_27131);
xnor U38110 (N_38110,N_23298,N_24186);
xor U38111 (N_38111,N_25263,N_24070);
xnor U38112 (N_38112,N_26659,N_26560);
or U38113 (N_38113,N_23139,N_29030);
and U38114 (N_38114,N_25110,N_26274);
nor U38115 (N_38115,N_22872,N_21188);
nor U38116 (N_38116,N_25231,N_27866);
xnor U38117 (N_38117,N_29948,N_27502);
or U38118 (N_38118,N_28993,N_27526);
nor U38119 (N_38119,N_23104,N_23458);
and U38120 (N_38120,N_23138,N_29591);
nor U38121 (N_38121,N_26680,N_25310);
nand U38122 (N_38122,N_29942,N_22674);
xor U38123 (N_38123,N_27933,N_25783);
xnor U38124 (N_38124,N_29499,N_23629);
or U38125 (N_38125,N_21901,N_26915);
or U38126 (N_38126,N_23950,N_29622);
or U38127 (N_38127,N_24089,N_26818);
and U38128 (N_38128,N_26443,N_22376);
or U38129 (N_38129,N_22547,N_25417);
nand U38130 (N_38130,N_25316,N_21678);
nand U38131 (N_38131,N_25942,N_25506);
xor U38132 (N_38132,N_22706,N_21556);
nand U38133 (N_38133,N_21672,N_29829);
and U38134 (N_38134,N_24167,N_28471);
nor U38135 (N_38135,N_28404,N_28255);
or U38136 (N_38136,N_29608,N_28835);
and U38137 (N_38137,N_26682,N_25269);
and U38138 (N_38138,N_22704,N_23784);
and U38139 (N_38139,N_24216,N_22140);
and U38140 (N_38140,N_28010,N_27442);
nand U38141 (N_38141,N_29859,N_21626);
nor U38142 (N_38142,N_23903,N_28894);
or U38143 (N_38143,N_23881,N_28902);
nand U38144 (N_38144,N_23242,N_20296);
xnor U38145 (N_38145,N_20163,N_29242);
nand U38146 (N_38146,N_27864,N_28836);
nand U38147 (N_38147,N_24505,N_22355);
and U38148 (N_38148,N_21639,N_26566);
nand U38149 (N_38149,N_28375,N_28950);
and U38150 (N_38150,N_22197,N_20910);
xnor U38151 (N_38151,N_23508,N_20922);
nor U38152 (N_38152,N_26139,N_27785);
nor U38153 (N_38153,N_29602,N_25955);
xnor U38154 (N_38154,N_22769,N_29223);
nand U38155 (N_38155,N_23300,N_27101);
and U38156 (N_38156,N_28542,N_28674);
nand U38157 (N_38157,N_25854,N_21169);
xor U38158 (N_38158,N_24863,N_23877);
nand U38159 (N_38159,N_23507,N_26465);
or U38160 (N_38160,N_23001,N_24976);
nor U38161 (N_38161,N_22782,N_23049);
xnor U38162 (N_38162,N_21969,N_26486);
or U38163 (N_38163,N_29589,N_28899);
nand U38164 (N_38164,N_28080,N_24861);
nand U38165 (N_38165,N_21766,N_25333);
nor U38166 (N_38166,N_24094,N_23633);
xnor U38167 (N_38167,N_27751,N_23868);
or U38168 (N_38168,N_27633,N_26114);
and U38169 (N_38169,N_21451,N_28381);
nand U38170 (N_38170,N_24165,N_29184);
nor U38171 (N_38171,N_28498,N_23883);
or U38172 (N_38172,N_27292,N_22453);
nor U38173 (N_38173,N_29314,N_21542);
nand U38174 (N_38174,N_26457,N_21067);
nand U38175 (N_38175,N_20928,N_22849);
nand U38176 (N_38176,N_28657,N_28743);
or U38177 (N_38177,N_23910,N_29194);
nor U38178 (N_38178,N_27640,N_20718);
or U38179 (N_38179,N_25947,N_25768);
nor U38180 (N_38180,N_25941,N_22737);
nor U38181 (N_38181,N_20793,N_25372);
and U38182 (N_38182,N_20134,N_28326);
nor U38183 (N_38183,N_20425,N_20025);
nand U38184 (N_38184,N_23272,N_28860);
xor U38185 (N_38185,N_23159,N_25203);
or U38186 (N_38186,N_25872,N_27850);
nor U38187 (N_38187,N_22095,N_25147);
nor U38188 (N_38188,N_25434,N_25447);
xnor U38189 (N_38189,N_28926,N_27767);
or U38190 (N_38190,N_20555,N_28516);
nor U38191 (N_38191,N_23669,N_22693);
nand U38192 (N_38192,N_21881,N_28282);
or U38193 (N_38193,N_28253,N_26280);
or U38194 (N_38194,N_24050,N_24097);
xnor U38195 (N_38195,N_25760,N_27068);
nor U38196 (N_38196,N_27771,N_29312);
xor U38197 (N_38197,N_28151,N_22928);
nor U38198 (N_38198,N_22545,N_24415);
nand U38199 (N_38199,N_29821,N_25101);
and U38200 (N_38200,N_27675,N_28000);
nor U38201 (N_38201,N_20142,N_27076);
xor U38202 (N_38202,N_27194,N_28130);
nor U38203 (N_38203,N_29394,N_23234);
or U38204 (N_38204,N_24652,N_27429);
xor U38205 (N_38205,N_27565,N_25655);
nor U38206 (N_38206,N_25274,N_25502);
nand U38207 (N_38207,N_22586,N_28720);
xnor U38208 (N_38208,N_24650,N_25460);
xor U38209 (N_38209,N_25116,N_27321);
nor U38210 (N_38210,N_28536,N_22789);
or U38211 (N_38211,N_24766,N_29481);
xor U38212 (N_38212,N_25786,N_28373);
and U38213 (N_38213,N_28218,N_23902);
or U38214 (N_38214,N_24156,N_23130);
nand U38215 (N_38215,N_22172,N_22229);
nor U38216 (N_38216,N_24909,N_25163);
xnor U38217 (N_38217,N_27259,N_25516);
nand U38218 (N_38218,N_24304,N_23517);
xor U38219 (N_38219,N_28802,N_27133);
xnor U38220 (N_38220,N_28404,N_29672);
nor U38221 (N_38221,N_22512,N_22684);
nor U38222 (N_38222,N_28440,N_22449);
or U38223 (N_38223,N_27814,N_28838);
nand U38224 (N_38224,N_20529,N_23711);
nor U38225 (N_38225,N_24500,N_27108);
or U38226 (N_38226,N_29977,N_27899);
nor U38227 (N_38227,N_27085,N_26765);
xor U38228 (N_38228,N_22218,N_28407);
and U38229 (N_38229,N_22688,N_23913);
nor U38230 (N_38230,N_23656,N_21723);
xor U38231 (N_38231,N_28782,N_25332);
nor U38232 (N_38232,N_21561,N_22231);
xnor U38233 (N_38233,N_27267,N_26694);
xnor U38234 (N_38234,N_22316,N_24771);
nand U38235 (N_38235,N_22847,N_20045);
or U38236 (N_38236,N_22505,N_25807);
or U38237 (N_38237,N_27185,N_24126);
nor U38238 (N_38238,N_29722,N_20706);
and U38239 (N_38239,N_22219,N_21709);
xor U38240 (N_38240,N_25521,N_21562);
and U38241 (N_38241,N_20370,N_25477);
or U38242 (N_38242,N_22558,N_26974);
nor U38243 (N_38243,N_20202,N_22297);
nor U38244 (N_38244,N_21835,N_24488);
and U38245 (N_38245,N_26364,N_24535);
xnor U38246 (N_38246,N_23424,N_29730);
xor U38247 (N_38247,N_21283,N_21394);
nor U38248 (N_38248,N_25039,N_21350);
or U38249 (N_38249,N_28019,N_26678);
xnor U38250 (N_38250,N_28286,N_24651);
nor U38251 (N_38251,N_21857,N_22977);
nand U38252 (N_38252,N_23621,N_20991);
nor U38253 (N_38253,N_28866,N_27885);
and U38254 (N_38254,N_29443,N_27340);
and U38255 (N_38255,N_23221,N_23370);
and U38256 (N_38256,N_23522,N_23624);
nand U38257 (N_38257,N_28916,N_27943);
and U38258 (N_38258,N_24411,N_20066);
or U38259 (N_38259,N_29890,N_26718);
or U38260 (N_38260,N_21476,N_23363);
or U38261 (N_38261,N_20949,N_20173);
nand U38262 (N_38262,N_29082,N_27067);
nor U38263 (N_38263,N_24939,N_27171);
xnor U38264 (N_38264,N_27669,N_21890);
nor U38265 (N_38265,N_22193,N_22643);
nor U38266 (N_38266,N_20923,N_24452);
and U38267 (N_38267,N_24943,N_25102);
nand U38268 (N_38268,N_29691,N_27145);
or U38269 (N_38269,N_23547,N_22836);
and U38270 (N_38270,N_29665,N_21766);
or U38271 (N_38271,N_23633,N_23952);
or U38272 (N_38272,N_22669,N_25910);
xor U38273 (N_38273,N_27522,N_29912);
xnor U38274 (N_38274,N_29640,N_21359);
or U38275 (N_38275,N_24184,N_20834);
xor U38276 (N_38276,N_23990,N_25089);
nor U38277 (N_38277,N_25071,N_26662);
nand U38278 (N_38278,N_20892,N_21854);
xor U38279 (N_38279,N_24270,N_24755);
nor U38280 (N_38280,N_21525,N_23432);
xnor U38281 (N_38281,N_26042,N_22058);
or U38282 (N_38282,N_25277,N_26465);
and U38283 (N_38283,N_28337,N_22674);
and U38284 (N_38284,N_20858,N_23121);
nor U38285 (N_38285,N_22771,N_25202);
xor U38286 (N_38286,N_25237,N_22746);
nand U38287 (N_38287,N_22680,N_22602);
or U38288 (N_38288,N_23583,N_21496);
nand U38289 (N_38289,N_23834,N_27624);
and U38290 (N_38290,N_25829,N_28901);
nor U38291 (N_38291,N_24192,N_24703);
nand U38292 (N_38292,N_22650,N_25243);
nand U38293 (N_38293,N_26119,N_26148);
nand U38294 (N_38294,N_29446,N_21738);
nor U38295 (N_38295,N_22376,N_23485);
nand U38296 (N_38296,N_25196,N_28421);
and U38297 (N_38297,N_20638,N_20405);
and U38298 (N_38298,N_29297,N_22204);
or U38299 (N_38299,N_24444,N_29770);
nor U38300 (N_38300,N_21497,N_23826);
xnor U38301 (N_38301,N_27526,N_22585);
and U38302 (N_38302,N_21318,N_26836);
and U38303 (N_38303,N_25819,N_29713);
and U38304 (N_38304,N_28987,N_28520);
xnor U38305 (N_38305,N_20772,N_27583);
nand U38306 (N_38306,N_24415,N_21171);
nor U38307 (N_38307,N_22047,N_25189);
xnor U38308 (N_38308,N_20255,N_23599);
nand U38309 (N_38309,N_27413,N_24741);
or U38310 (N_38310,N_27312,N_26306);
nor U38311 (N_38311,N_22193,N_26721);
nor U38312 (N_38312,N_20284,N_28217);
nand U38313 (N_38313,N_25512,N_26484);
nor U38314 (N_38314,N_24182,N_27732);
nor U38315 (N_38315,N_25696,N_22296);
nor U38316 (N_38316,N_29230,N_25785);
and U38317 (N_38317,N_22354,N_29227);
and U38318 (N_38318,N_27430,N_26207);
nand U38319 (N_38319,N_29027,N_21776);
nor U38320 (N_38320,N_23784,N_29642);
and U38321 (N_38321,N_24190,N_27859);
nor U38322 (N_38322,N_28146,N_24479);
xnor U38323 (N_38323,N_28418,N_25837);
nand U38324 (N_38324,N_25139,N_27330);
and U38325 (N_38325,N_28994,N_27521);
xor U38326 (N_38326,N_27825,N_25879);
nand U38327 (N_38327,N_24262,N_29496);
and U38328 (N_38328,N_26756,N_27556);
or U38329 (N_38329,N_28208,N_25228);
xor U38330 (N_38330,N_24204,N_22646);
or U38331 (N_38331,N_24135,N_27110);
nor U38332 (N_38332,N_22419,N_23306);
xnor U38333 (N_38333,N_25312,N_26640);
nor U38334 (N_38334,N_26268,N_21829);
nor U38335 (N_38335,N_24340,N_23803);
or U38336 (N_38336,N_20358,N_24420);
nor U38337 (N_38337,N_28153,N_22828);
nand U38338 (N_38338,N_28508,N_28627);
nand U38339 (N_38339,N_21673,N_23004);
xor U38340 (N_38340,N_25582,N_27327);
and U38341 (N_38341,N_25753,N_27712);
and U38342 (N_38342,N_29838,N_23919);
and U38343 (N_38343,N_20205,N_25408);
nand U38344 (N_38344,N_29841,N_21188);
nor U38345 (N_38345,N_26463,N_20140);
and U38346 (N_38346,N_24426,N_27271);
nand U38347 (N_38347,N_26053,N_20098);
nand U38348 (N_38348,N_25259,N_26030);
nor U38349 (N_38349,N_27664,N_24852);
xor U38350 (N_38350,N_20468,N_21016);
or U38351 (N_38351,N_28942,N_29585);
and U38352 (N_38352,N_29163,N_29334);
or U38353 (N_38353,N_28278,N_23487);
and U38354 (N_38354,N_20748,N_25996);
xnor U38355 (N_38355,N_26996,N_23712);
nand U38356 (N_38356,N_23681,N_29289);
nor U38357 (N_38357,N_29616,N_27212);
xor U38358 (N_38358,N_28094,N_28471);
nand U38359 (N_38359,N_22852,N_29014);
and U38360 (N_38360,N_24245,N_22712);
nor U38361 (N_38361,N_29899,N_27108);
xor U38362 (N_38362,N_29179,N_25486);
or U38363 (N_38363,N_20954,N_26223);
nor U38364 (N_38364,N_26740,N_22311);
xor U38365 (N_38365,N_25715,N_27249);
nor U38366 (N_38366,N_25144,N_24828);
nand U38367 (N_38367,N_27562,N_23483);
xnor U38368 (N_38368,N_20764,N_27180);
nand U38369 (N_38369,N_27040,N_20215);
xor U38370 (N_38370,N_25327,N_27434);
and U38371 (N_38371,N_22058,N_26018);
and U38372 (N_38372,N_21365,N_26683);
nor U38373 (N_38373,N_25675,N_26155);
xnor U38374 (N_38374,N_21850,N_25982);
and U38375 (N_38375,N_20153,N_21995);
xnor U38376 (N_38376,N_24219,N_21169);
or U38377 (N_38377,N_23736,N_22253);
nand U38378 (N_38378,N_29566,N_26951);
or U38379 (N_38379,N_21075,N_27168);
nor U38380 (N_38380,N_20708,N_20553);
and U38381 (N_38381,N_24068,N_28650);
nand U38382 (N_38382,N_23623,N_22011);
nor U38383 (N_38383,N_29333,N_26221);
xnor U38384 (N_38384,N_25248,N_21058);
or U38385 (N_38385,N_21833,N_25683);
nand U38386 (N_38386,N_23318,N_25836);
nand U38387 (N_38387,N_25006,N_29563);
and U38388 (N_38388,N_24271,N_20782);
nand U38389 (N_38389,N_27932,N_22093);
or U38390 (N_38390,N_24432,N_24981);
xor U38391 (N_38391,N_28280,N_26586);
or U38392 (N_38392,N_27682,N_25923);
nor U38393 (N_38393,N_20633,N_22174);
xnor U38394 (N_38394,N_28017,N_29458);
nand U38395 (N_38395,N_20956,N_25980);
and U38396 (N_38396,N_22933,N_28100);
or U38397 (N_38397,N_27420,N_26721);
and U38398 (N_38398,N_21209,N_21755);
nand U38399 (N_38399,N_25156,N_20289);
or U38400 (N_38400,N_25529,N_28347);
nand U38401 (N_38401,N_20805,N_23495);
or U38402 (N_38402,N_27860,N_23409);
nand U38403 (N_38403,N_21533,N_22072);
xor U38404 (N_38404,N_27782,N_29423);
xnor U38405 (N_38405,N_28982,N_20883);
nand U38406 (N_38406,N_28263,N_27626);
xnor U38407 (N_38407,N_27126,N_25238);
and U38408 (N_38408,N_27280,N_27548);
or U38409 (N_38409,N_23743,N_28492);
nand U38410 (N_38410,N_24627,N_28266);
or U38411 (N_38411,N_20909,N_23166);
xor U38412 (N_38412,N_22739,N_29666);
nand U38413 (N_38413,N_23140,N_20193);
or U38414 (N_38414,N_22435,N_22394);
xnor U38415 (N_38415,N_25222,N_26496);
or U38416 (N_38416,N_28303,N_26188);
nand U38417 (N_38417,N_26333,N_27037);
xnor U38418 (N_38418,N_26212,N_26539);
and U38419 (N_38419,N_26902,N_22104);
and U38420 (N_38420,N_23793,N_24381);
xor U38421 (N_38421,N_21209,N_20151);
or U38422 (N_38422,N_29144,N_25519);
nor U38423 (N_38423,N_20888,N_27349);
nand U38424 (N_38424,N_24820,N_20731);
or U38425 (N_38425,N_23344,N_28442);
nor U38426 (N_38426,N_21844,N_21339);
and U38427 (N_38427,N_29796,N_27883);
nor U38428 (N_38428,N_21306,N_26662);
nand U38429 (N_38429,N_23691,N_20394);
and U38430 (N_38430,N_27432,N_22067);
nor U38431 (N_38431,N_21509,N_21654);
xnor U38432 (N_38432,N_22501,N_26619);
xnor U38433 (N_38433,N_26082,N_29393);
nor U38434 (N_38434,N_21763,N_23034);
xor U38435 (N_38435,N_21824,N_27523);
nand U38436 (N_38436,N_21005,N_23589);
or U38437 (N_38437,N_27135,N_27643);
nor U38438 (N_38438,N_28165,N_28667);
and U38439 (N_38439,N_20287,N_21400);
nand U38440 (N_38440,N_28618,N_24789);
nor U38441 (N_38441,N_23693,N_29439);
xnor U38442 (N_38442,N_25929,N_22617);
or U38443 (N_38443,N_24795,N_22837);
nor U38444 (N_38444,N_27803,N_27009);
and U38445 (N_38445,N_25754,N_21129);
or U38446 (N_38446,N_22829,N_28157);
and U38447 (N_38447,N_21411,N_22914);
and U38448 (N_38448,N_26646,N_20336);
nand U38449 (N_38449,N_20082,N_24525);
or U38450 (N_38450,N_26922,N_29178);
xor U38451 (N_38451,N_24773,N_26854);
and U38452 (N_38452,N_26678,N_26420);
nor U38453 (N_38453,N_26623,N_28942);
nor U38454 (N_38454,N_29064,N_20912);
xor U38455 (N_38455,N_27102,N_25822);
nand U38456 (N_38456,N_22910,N_20385);
nand U38457 (N_38457,N_25721,N_26254);
or U38458 (N_38458,N_22279,N_20530);
nand U38459 (N_38459,N_26030,N_23887);
xor U38460 (N_38460,N_24740,N_21315);
nand U38461 (N_38461,N_20637,N_29423);
and U38462 (N_38462,N_21056,N_27639);
or U38463 (N_38463,N_20264,N_29066);
nand U38464 (N_38464,N_22073,N_29470);
or U38465 (N_38465,N_20791,N_28878);
xor U38466 (N_38466,N_25194,N_25990);
nor U38467 (N_38467,N_26525,N_27661);
xnor U38468 (N_38468,N_24814,N_20779);
and U38469 (N_38469,N_26281,N_21052);
nor U38470 (N_38470,N_21108,N_21594);
or U38471 (N_38471,N_27619,N_28901);
and U38472 (N_38472,N_23063,N_27468);
and U38473 (N_38473,N_25064,N_24656);
or U38474 (N_38474,N_29434,N_25354);
and U38475 (N_38475,N_25889,N_29193);
nand U38476 (N_38476,N_23173,N_21822);
xnor U38477 (N_38477,N_20235,N_28994);
nand U38478 (N_38478,N_20988,N_25649);
nand U38479 (N_38479,N_27679,N_24975);
xor U38480 (N_38480,N_29290,N_22269);
xor U38481 (N_38481,N_29290,N_21327);
and U38482 (N_38482,N_26403,N_23644);
and U38483 (N_38483,N_21774,N_24303);
and U38484 (N_38484,N_28245,N_28990);
nand U38485 (N_38485,N_20921,N_22509);
xor U38486 (N_38486,N_23956,N_22327);
or U38487 (N_38487,N_26333,N_22040);
nand U38488 (N_38488,N_26763,N_28935);
nand U38489 (N_38489,N_20409,N_25411);
nor U38490 (N_38490,N_23921,N_26016);
or U38491 (N_38491,N_20084,N_28291);
and U38492 (N_38492,N_26307,N_29126);
nor U38493 (N_38493,N_21701,N_25501);
nand U38494 (N_38494,N_21602,N_27241);
or U38495 (N_38495,N_27224,N_23019);
and U38496 (N_38496,N_26845,N_23887);
or U38497 (N_38497,N_24529,N_21870);
nand U38498 (N_38498,N_24527,N_28850);
and U38499 (N_38499,N_21114,N_25622);
nor U38500 (N_38500,N_24048,N_28101);
and U38501 (N_38501,N_28120,N_22220);
or U38502 (N_38502,N_21620,N_22299);
xor U38503 (N_38503,N_23629,N_26003);
nor U38504 (N_38504,N_25149,N_20681);
or U38505 (N_38505,N_28438,N_27228);
xnor U38506 (N_38506,N_27301,N_27776);
or U38507 (N_38507,N_29689,N_21107);
and U38508 (N_38508,N_21352,N_20802);
xor U38509 (N_38509,N_23819,N_22235);
xnor U38510 (N_38510,N_27746,N_23405);
and U38511 (N_38511,N_24306,N_23765);
or U38512 (N_38512,N_26389,N_26887);
nor U38513 (N_38513,N_23406,N_21397);
and U38514 (N_38514,N_26913,N_24734);
xor U38515 (N_38515,N_25485,N_20280);
nand U38516 (N_38516,N_28928,N_27574);
and U38517 (N_38517,N_29278,N_29384);
nand U38518 (N_38518,N_23901,N_24977);
xor U38519 (N_38519,N_21785,N_23669);
or U38520 (N_38520,N_27276,N_27003);
xnor U38521 (N_38521,N_25361,N_26107);
or U38522 (N_38522,N_28052,N_24023);
nor U38523 (N_38523,N_23259,N_20484);
and U38524 (N_38524,N_29097,N_22885);
nor U38525 (N_38525,N_20297,N_22344);
and U38526 (N_38526,N_27338,N_29308);
or U38527 (N_38527,N_26354,N_20145);
nor U38528 (N_38528,N_22902,N_24993);
nor U38529 (N_38529,N_22517,N_21911);
and U38530 (N_38530,N_26709,N_24795);
nor U38531 (N_38531,N_23211,N_24171);
nand U38532 (N_38532,N_25952,N_27915);
nor U38533 (N_38533,N_27113,N_23731);
and U38534 (N_38534,N_21911,N_22731);
nand U38535 (N_38535,N_23851,N_29469);
xor U38536 (N_38536,N_22896,N_29164);
nand U38537 (N_38537,N_27057,N_28390);
nand U38538 (N_38538,N_27998,N_25231);
nor U38539 (N_38539,N_23963,N_28782);
xnor U38540 (N_38540,N_28744,N_21696);
nor U38541 (N_38541,N_26612,N_20451);
nand U38542 (N_38542,N_22852,N_28547);
nand U38543 (N_38543,N_20269,N_27550);
or U38544 (N_38544,N_22845,N_28759);
and U38545 (N_38545,N_21035,N_21340);
and U38546 (N_38546,N_22848,N_27395);
or U38547 (N_38547,N_24894,N_23368);
xor U38548 (N_38548,N_27863,N_25908);
nor U38549 (N_38549,N_20215,N_27461);
and U38550 (N_38550,N_28261,N_21883);
and U38551 (N_38551,N_25097,N_20073);
nand U38552 (N_38552,N_28001,N_21817);
nand U38553 (N_38553,N_20776,N_21292);
xnor U38554 (N_38554,N_29008,N_27936);
nor U38555 (N_38555,N_25213,N_22689);
nand U38556 (N_38556,N_23614,N_25118);
xnor U38557 (N_38557,N_21175,N_24789);
or U38558 (N_38558,N_22714,N_20007);
xnor U38559 (N_38559,N_23229,N_21920);
and U38560 (N_38560,N_21890,N_21319);
and U38561 (N_38561,N_24676,N_21541);
xor U38562 (N_38562,N_20496,N_27446);
nand U38563 (N_38563,N_25116,N_28998);
xor U38564 (N_38564,N_25304,N_26555);
nand U38565 (N_38565,N_20945,N_21444);
nor U38566 (N_38566,N_29654,N_26859);
nand U38567 (N_38567,N_25796,N_23167);
or U38568 (N_38568,N_20954,N_27869);
nor U38569 (N_38569,N_28154,N_21988);
or U38570 (N_38570,N_23533,N_25245);
nand U38571 (N_38571,N_27288,N_25061);
nand U38572 (N_38572,N_22352,N_27731);
nand U38573 (N_38573,N_29886,N_23444);
xnor U38574 (N_38574,N_20953,N_25439);
nor U38575 (N_38575,N_20679,N_22897);
and U38576 (N_38576,N_26519,N_27600);
and U38577 (N_38577,N_22875,N_22630);
or U38578 (N_38578,N_29826,N_25198);
and U38579 (N_38579,N_25598,N_22564);
nand U38580 (N_38580,N_25460,N_21664);
xor U38581 (N_38581,N_20097,N_25928);
nor U38582 (N_38582,N_20303,N_25983);
nor U38583 (N_38583,N_22045,N_28027);
or U38584 (N_38584,N_25122,N_20990);
nand U38585 (N_38585,N_27098,N_27578);
nor U38586 (N_38586,N_27865,N_28628);
or U38587 (N_38587,N_25425,N_25925);
nor U38588 (N_38588,N_26899,N_29517);
nand U38589 (N_38589,N_29289,N_23323);
and U38590 (N_38590,N_22536,N_25760);
xor U38591 (N_38591,N_29633,N_22632);
nand U38592 (N_38592,N_20120,N_28472);
nand U38593 (N_38593,N_26824,N_25477);
or U38594 (N_38594,N_22321,N_28315);
nor U38595 (N_38595,N_22010,N_23916);
xnor U38596 (N_38596,N_23551,N_27463);
or U38597 (N_38597,N_23073,N_27461);
nand U38598 (N_38598,N_27520,N_29894);
nand U38599 (N_38599,N_25674,N_21790);
or U38600 (N_38600,N_20716,N_26928);
nand U38601 (N_38601,N_28772,N_29194);
xnor U38602 (N_38602,N_21248,N_28914);
xnor U38603 (N_38603,N_28257,N_28208);
and U38604 (N_38604,N_21753,N_24493);
nor U38605 (N_38605,N_27058,N_29310);
nor U38606 (N_38606,N_22929,N_28807);
and U38607 (N_38607,N_27411,N_26744);
xnor U38608 (N_38608,N_22557,N_28898);
or U38609 (N_38609,N_22698,N_24427);
or U38610 (N_38610,N_21871,N_27018);
xor U38611 (N_38611,N_24201,N_28402);
nand U38612 (N_38612,N_25182,N_28958);
or U38613 (N_38613,N_23629,N_24317);
and U38614 (N_38614,N_21770,N_27189);
nor U38615 (N_38615,N_24215,N_22187);
and U38616 (N_38616,N_25304,N_28239);
and U38617 (N_38617,N_23819,N_24025);
nor U38618 (N_38618,N_23904,N_28765);
nand U38619 (N_38619,N_24840,N_21871);
nor U38620 (N_38620,N_27881,N_27333);
nand U38621 (N_38621,N_29746,N_29832);
nor U38622 (N_38622,N_23919,N_24510);
nor U38623 (N_38623,N_22591,N_21571);
nand U38624 (N_38624,N_25237,N_28154);
or U38625 (N_38625,N_22108,N_29872);
and U38626 (N_38626,N_20182,N_26157);
and U38627 (N_38627,N_26237,N_28340);
xor U38628 (N_38628,N_26640,N_27113);
or U38629 (N_38629,N_25851,N_22784);
nand U38630 (N_38630,N_25220,N_26374);
nor U38631 (N_38631,N_28296,N_21890);
nand U38632 (N_38632,N_24655,N_24151);
nor U38633 (N_38633,N_26608,N_22233);
xor U38634 (N_38634,N_23417,N_29125);
and U38635 (N_38635,N_24526,N_21061);
or U38636 (N_38636,N_25899,N_22231);
xnor U38637 (N_38637,N_27576,N_24511);
or U38638 (N_38638,N_27197,N_29232);
or U38639 (N_38639,N_21028,N_28543);
or U38640 (N_38640,N_20741,N_24334);
xor U38641 (N_38641,N_23305,N_20739);
nand U38642 (N_38642,N_20211,N_23659);
xor U38643 (N_38643,N_26110,N_29887);
nor U38644 (N_38644,N_21913,N_25145);
nand U38645 (N_38645,N_27759,N_24479);
and U38646 (N_38646,N_20195,N_28888);
nor U38647 (N_38647,N_29114,N_29379);
nand U38648 (N_38648,N_28993,N_20720);
xor U38649 (N_38649,N_24261,N_25322);
xnor U38650 (N_38650,N_20060,N_23808);
or U38651 (N_38651,N_26910,N_25686);
nor U38652 (N_38652,N_27709,N_27285);
or U38653 (N_38653,N_23818,N_29209);
and U38654 (N_38654,N_24837,N_29853);
xor U38655 (N_38655,N_22404,N_22963);
and U38656 (N_38656,N_29897,N_20043);
and U38657 (N_38657,N_29202,N_20697);
or U38658 (N_38658,N_20303,N_28357);
xnor U38659 (N_38659,N_20154,N_28730);
nor U38660 (N_38660,N_29430,N_22059);
xor U38661 (N_38661,N_22351,N_27385);
nand U38662 (N_38662,N_27208,N_25136);
xnor U38663 (N_38663,N_25777,N_27696);
and U38664 (N_38664,N_22114,N_25212);
and U38665 (N_38665,N_28428,N_27953);
nand U38666 (N_38666,N_26027,N_28596);
nand U38667 (N_38667,N_21030,N_27801);
nand U38668 (N_38668,N_28045,N_29035);
nand U38669 (N_38669,N_20749,N_28875);
nand U38670 (N_38670,N_23548,N_26954);
and U38671 (N_38671,N_23618,N_20648);
and U38672 (N_38672,N_25308,N_29534);
nand U38673 (N_38673,N_20007,N_25770);
or U38674 (N_38674,N_28414,N_28115);
nor U38675 (N_38675,N_22985,N_20057);
nor U38676 (N_38676,N_23721,N_22272);
or U38677 (N_38677,N_28748,N_29236);
nand U38678 (N_38678,N_25497,N_29557);
and U38679 (N_38679,N_27707,N_24105);
xnor U38680 (N_38680,N_25548,N_25785);
or U38681 (N_38681,N_29618,N_28386);
or U38682 (N_38682,N_28106,N_24495);
nor U38683 (N_38683,N_23214,N_23044);
xor U38684 (N_38684,N_25764,N_20511);
and U38685 (N_38685,N_29515,N_21917);
nand U38686 (N_38686,N_20044,N_25403);
and U38687 (N_38687,N_23403,N_26767);
and U38688 (N_38688,N_24660,N_20961);
and U38689 (N_38689,N_22701,N_20282);
nor U38690 (N_38690,N_28456,N_24749);
or U38691 (N_38691,N_22066,N_29513);
nor U38692 (N_38692,N_24825,N_21269);
or U38693 (N_38693,N_29836,N_28807);
nor U38694 (N_38694,N_25629,N_27369);
or U38695 (N_38695,N_25192,N_25919);
xnor U38696 (N_38696,N_28821,N_20078);
and U38697 (N_38697,N_21456,N_26591);
nor U38698 (N_38698,N_29202,N_26513);
nor U38699 (N_38699,N_28067,N_20996);
and U38700 (N_38700,N_21769,N_25261);
and U38701 (N_38701,N_23123,N_21085);
and U38702 (N_38702,N_26897,N_25218);
and U38703 (N_38703,N_28122,N_24911);
or U38704 (N_38704,N_29321,N_20648);
xnor U38705 (N_38705,N_20587,N_23211);
and U38706 (N_38706,N_21102,N_23864);
nor U38707 (N_38707,N_25640,N_22684);
and U38708 (N_38708,N_20026,N_22778);
or U38709 (N_38709,N_21738,N_29638);
nor U38710 (N_38710,N_25408,N_25281);
nor U38711 (N_38711,N_25232,N_23233);
and U38712 (N_38712,N_26769,N_22816);
or U38713 (N_38713,N_22554,N_24264);
xor U38714 (N_38714,N_27897,N_28642);
xnor U38715 (N_38715,N_27879,N_29567);
and U38716 (N_38716,N_24624,N_29825);
xor U38717 (N_38717,N_21586,N_29495);
nand U38718 (N_38718,N_22430,N_26178);
and U38719 (N_38719,N_24655,N_27873);
xnor U38720 (N_38720,N_23400,N_27628);
or U38721 (N_38721,N_23540,N_23084);
xnor U38722 (N_38722,N_25724,N_26986);
nor U38723 (N_38723,N_26070,N_27810);
nand U38724 (N_38724,N_29436,N_22077);
and U38725 (N_38725,N_22761,N_21523);
xnor U38726 (N_38726,N_25195,N_20247);
nand U38727 (N_38727,N_20442,N_28751);
or U38728 (N_38728,N_27059,N_29858);
or U38729 (N_38729,N_25462,N_21161);
xnor U38730 (N_38730,N_21068,N_29068);
xnor U38731 (N_38731,N_28463,N_22356);
xnor U38732 (N_38732,N_27558,N_28088);
nor U38733 (N_38733,N_28368,N_27530);
nand U38734 (N_38734,N_24679,N_24751);
nand U38735 (N_38735,N_26541,N_22264);
nand U38736 (N_38736,N_21031,N_23383);
and U38737 (N_38737,N_22859,N_23459);
and U38738 (N_38738,N_22523,N_20585);
and U38739 (N_38739,N_28286,N_22990);
and U38740 (N_38740,N_29134,N_24666);
nand U38741 (N_38741,N_27066,N_22944);
nand U38742 (N_38742,N_24735,N_21976);
xor U38743 (N_38743,N_28773,N_23214);
nor U38744 (N_38744,N_26118,N_27385);
nor U38745 (N_38745,N_27993,N_23667);
or U38746 (N_38746,N_25819,N_22986);
nor U38747 (N_38747,N_28057,N_22597);
xnor U38748 (N_38748,N_27749,N_25480);
or U38749 (N_38749,N_29403,N_22309);
nand U38750 (N_38750,N_24646,N_21626);
nor U38751 (N_38751,N_27270,N_27661);
or U38752 (N_38752,N_20323,N_22258);
or U38753 (N_38753,N_28018,N_27394);
or U38754 (N_38754,N_27445,N_29333);
xor U38755 (N_38755,N_27057,N_26876);
xor U38756 (N_38756,N_22423,N_27490);
nor U38757 (N_38757,N_28641,N_24230);
xor U38758 (N_38758,N_24534,N_27346);
nor U38759 (N_38759,N_29339,N_26962);
xor U38760 (N_38760,N_21421,N_22168);
nand U38761 (N_38761,N_26933,N_24541);
xor U38762 (N_38762,N_29925,N_29490);
nand U38763 (N_38763,N_27410,N_27368);
nand U38764 (N_38764,N_23645,N_21512);
and U38765 (N_38765,N_23503,N_21525);
xnor U38766 (N_38766,N_20261,N_23434);
xor U38767 (N_38767,N_20568,N_27200);
and U38768 (N_38768,N_26584,N_27959);
nand U38769 (N_38769,N_21537,N_26640);
and U38770 (N_38770,N_21709,N_25822);
or U38771 (N_38771,N_23252,N_23056);
nand U38772 (N_38772,N_27981,N_27810);
or U38773 (N_38773,N_25860,N_26571);
xnor U38774 (N_38774,N_27035,N_20870);
or U38775 (N_38775,N_22145,N_28587);
or U38776 (N_38776,N_29349,N_21106);
and U38777 (N_38777,N_22640,N_22347);
xor U38778 (N_38778,N_23042,N_25158);
nand U38779 (N_38779,N_27956,N_21610);
nand U38780 (N_38780,N_29629,N_25129);
or U38781 (N_38781,N_26550,N_29965);
and U38782 (N_38782,N_21947,N_25950);
and U38783 (N_38783,N_22085,N_26120);
and U38784 (N_38784,N_24899,N_24633);
nor U38785 (N_38785,N_21456,N_25136);
or U38786 (N_38786,N_27888,N_24204);
nand U38787 (N_38787,N_28858,N_23165);
nand U38788 (N_38788,N_21694,N_21162);
and U38789 (N_38789,N_28704,N_28643);
and U38790 (N_38790,N_29258,N_24799);
nand U38791 (N_38791,N_27213,N_27334);
and U38792 (N_38792,N_23261,N_21580);
or U38793 (N_38793,N_26926,N_28258);
nand U38794 (N_38794,N_26188,N_25945);
and U38795 (N_38795,N_20904,N_20312);
nor U38796 (N_38796,N_27500,N_20550);
nand U38797 (N_38797,N_22974,N_24043);
xnor U38798 (N_38798,N_21972,N_22986);
nand U38799 (N_38799,N_21732,N_24312);
and U38800 (N_38800,N_28620,N_27495);
and U38801 (N_38801,N_27560,N_26546);
nand U38802 (N_38802,N_22358,N_24183);
and U38803 (N_38803,N_24301,N_24128);
nor U38804 (N_38804,N_22882,N_22768);
xor U38805 (N_38805,N_23490,N_26891);
or U38806 (N_38806,N_29551,N_29308);
and U38807 (N_38807,N_24865,N_23981);
or U38808 (N_38808,N_25021,N_23681);
nand U38809 (N_38809,N_22045,N_24929);
or U38810 (N_38810,N_28727,N_27874);
nand U38811 (N_38811,N_27445,N_24062);
nor U38812 (N_38812,N_21313,N_23324);
xor U38813 (N_38813,N_22254,N_28119);
nand U38814 (N_38814,N_24364,N_23491);
nand U38815 (N_38815,N_24162,N_20732);
xnor U38816 (N_38816,N_22079,N_26640);
nand U38817 (N_38817,N_22088,N_22784);
nor U38818 (N_38818,N_27629,N_25709);
nor U38819 (N_38819,N_26971,N_26276);
or U38820 (N_38820,N_21337,N_24801);
nor U38821 (N_38821,N_28469,N_22967);
or U38822 (N_38822,N_29650,N_28950);
and U38823 (N_38823,N_23307,N_22267);
nor U38824 (N_38824,N_28655,N_25993);
xor U38825 (N_38825,N_28972,N_21669);
nand U38826 (N_38826,N_28520,N_29335);
xor U38827 (N_38827,N_29016,N_27928);
nor U38828 (N_38828,N_24134,N_26926);
nand U38829 (N_38829,N_24243,N_29914);
and U38830 (N_38830,N_28563,N_23531);
and U38831 (N_38831,N_29466,N_26479);
and U38832 (N_38832,N_20608,N_28719);
xor U38833 (N_38833,N_28236,N_23806);
or U38834 (N_38834,N_24790,N_26217);
and U38835 (N_38835,N_24606,N_22161);
nor U38836 (N_38836,N_22634,N_21218);
and U38837 (N_38837,N_28124,N_23734);
or U38838 (N_38838,N_28497,N_26131);
xnor U38839 (N_38839,N_21089,N_21000);
and U38840 (N_38840,N_20694,N_29015);
xor U38841 (N_38841,N_21884,N_20810);
or U38842 (N_38842,N_24878,N_22317);
nor U38843 (N_38843,N_25405,N_20424);
nand U38844 (N_38844,N_22247,N_23461);
and U38845 (N_38845,N_25254,N_24789);
nor U38846 (N_38846,N_24093,N_24275);
nand U38847 (N_38847,N_20756,N_24597);
and U38848 (N_38848,N_24326,N_27744);
nand U38849 (N_38849,N_24856,N_27304);
and U38850 (N_38850,N_29417,N_21996);
nand U38851 (N_38851,N_23205,N_25622);
nor U38852 (N_38852,N_25853,N_27485);
and U38853 (N_38853,N_23452,N_28764);
nor U38854 (N_38854,N_20741,N_25880);
nor U38855 (N_38855,N_26169,N_22889);
nand U38856 (N_38856,N_22105,N_23693);
and U38857 (N_38857,N_22805,N_20868);
or U38858 (N_38858,N_20223,N_26909);
xor U38859 (N_38859,N_23294,N_29195);
nand U38860 (N_38860,N_27323,N_29338);
nor U38861 (N_38861,N_29580,N_29585);
nor U38862 (N_38862,N_21615,N_26734);
nand U38863 (N_38863,N_22682,N_23462);
nor U38864 (N_38864,N_25245,N_24995);
and U38865 (N_38865,N_23610,N_25294);
or U38866 (N_38866,N_20817,N_22482);
nand U38867 (N_38867,N_22582,N_23747);
nand U38868 (N_38868,N_21140,N_22230);
or U38869 (N_38869,N_28488,N_23128);
nand U38870 (N_38870,N_21026,N_20182);
nor U38871 (N_38871,N_25989,N_28804);
xor U38872 (N_38872,N_22514,N_22029);
nand U38873 (N_38873,N_23256,N_25559);
xor U38874 (N_38874,N_27985,N_23145);
and U38875 (N_38875,N_23561,N_26790);
nor U38876 (N_38876,N_26257,N_24895);
nand U38877 (N_38877,N_24711,N_20834);
xnor U38878 (N_38878,N_25063,N_26549);
xnor U38879 (N_38879,N_26039,N_22882);
or U38880 (N_38880,N_27553,N_29461);
xnor U38881 (N_38881,N_23017,N_27935);
xnor U38882 (N_38882,N_29126,N_27987);
or U38883 (N_38883,N_28879,N_22154);
or U38884 (N_38884,N_21000,N_26045);
xor U38885 (N_38885,N_23840,N_23593);
and U38886 (N_38886,N_21142,N_22627);
or U38887 (N_38887,N_23336,N_26330);
or U38888 (N_38888,N_28399,N_22789);
nand U38889 (N_38889,N_20186,N_20527);
nand U38890 (N_38890,N_20565,N_20271);
nand U38891 (N_38891,N_25841,N_25126);
nand U38892 (N_38892,N_23951,N_27346);
xnor U38893 (N_38893,N_21978,N_27376);
nor U38894 (N_38894,N_21086,N_27154);
nand U38895 (N_38895,N_24474,N_21739);
nand U38896 (N_38896,N_28844,N_20981);
nand U38897 (N_38897,N_24999,N_25412);
nand U38898 (N_38898,N_20410,N_26234);
nor U38899 (N_38899,N_29981,N_21629);
or U38900 (N_38900,N_21979,N_25958);
nand U38901 (N_38901,N_26915,N_24838);
xnor U38902 (N_38902,N_21173,N_25262);
nand U38903 (N_38903,N_25327,N_22477);
xnor U38904 (N_38904,N_29919,N_24654);
and U38905 (N_38905,N_27301,N_20451);
nand U38906 (N_38906,N_27840,N_26974);
xor U38907 (N_38907,N_24511,N_21641);
nor U38908 (N_38908,N_24240,N_25880);
nor U38909 (N_38909,N_21279,N_21702);
nor U38910 (N_38910,N_28658,N_21467);
or U38911 (N_38911,N_28468,N_23250);
nand U38912 (N_38912,N_25726,N_28673);
nor U38913 (N_38913,N_28764,N_22852);
or U38914 (N_38914,N_25681,N_29823);
and U38915 (N_38915,N_21483,N_22021);
and U38916 (N_38916,N_26123,N_23332);
or U38917 (N_38917,N_22836,N_29853);
xor U38918 (N_38918,N_27460,N_21307);
nand U38919 (N_38919,N_23924,N_24099);
nand U38920 (N_38920,N_20158,N_24037);
xnor U38921 (N_38921,N_22964,N_24340);
nor U38922 (N_38922,N_23957,N_21062);
and U38923 (N_38923,N_23054,N_23062);
or U38924 (N_38924,N_25725,N_25763);
nor U38925 (N_38925,N_28558,N_27825);
xor U38926 (N_38926,N_25158,N_26158);
nand U38927 (N_38927,N_27186,N_23354);
nor U38928 (N_38928,N_29710,N_20045);
and U38929 (N_38929,N_21594,N_27416);
or U38930 (N_38930,N_26035,N_20651);
nor U38931 (N_38931,N_22408,N_24990);
nor U38932 (N_38932,N_26303,N_27211);
nand U38933 (N_38933,N_25820,N_27522);
or U38934 (N_38934,N_28586,N_24978);
xnor U38935 (N_38935,N_22133,N_27115);
xor U38936 (N_38936,N_24562,N_21764);
nor U38937 (N_38937,N_26034,N_25299);
or U38938 (N_38938,N_23488,N_29012);
and U38939 (N_38939,N_26723,N_25920);
and U38940 (N_38940,N_20761,N_24050);
and U38941 (N_38941,N_24183,N_27391);
nor U38942 (N_38942,N_21005,N_26647);
nor U38943 (N_38943,N_20851,N_25578);
nor U38944 (N_38944,N_27401,N_24004);
or U38945 (N_38945,N_21480,N_26784);
xor U38946 (N_38946,N_29761,N_22178);
and U38947 (N_38947,N_27305,N_21079);
or U38948 (N_38948,N_23627,N_27439);
and U38949 (N_38949,N_28301,N_24304);
xnor U38950 (N_38950,N_28466,N_23475);
and U38951 (N_38951,N_24624,N_26655);
xnor U38952 (N_38952,N_26483,N_25068);
and U38953 (N_38953,N_21306,N_28528);
xor U38954 (N_38954,N_29645,N_20731);
xnor U38955 (N_38955,N_25996,N_27385);
or U38956 (N_38956,N_20773,N_29318);
nor U38957 (N_38957,N_20052,N_27895);
nor U38958 (N_38958,N_23300,N_21666);
nor U38959 (N_38959,N_29160,N_26674);
xnor U38960 (N_38960,N_24744,N_27178);
nor U38961 (N_38961,N_24620,N_22739);
xnor U38962 (N_38962,N_27157,N_21715);
xor U38963 (N_38963,N_20958,N_29008);
or U38964 (N_38964,N_28114,N_25758);
nand U38965 (N_38965,N_28040,N_29798);
or U38966 (N_38966,N_25725,N_25840);
nor U38967 (N_38967,N_20915,N_26639);
nor U38968 (N_38968,N_26880,N_26614);
nor U38969 (N_38969,N_29773,N_23198);
and U38970 (N_38970,N_20532,N_28767);
xnor U38971 (N_38971,N_29748,N_24753);
or U38972 (N_38972,N_26597,N_29764);
and U38973 (N_38973,N_22144,N_28929);
and U38974 (N_38974,N_20953,N_22155);
nand U38975 (N_38975,N_23098,N_27186);
and U38976 (N_38976,N_27790,N_21062);
nor U38977 (N_38977,N_27812,N_23833);
and U38978 (N_38978,N_24696,N_21366);
nor U38979 (N_38979,N_26069,N_23073);
nor U38980 (N_38980,N_20221,N_29751);
xnor U38981 (N_38981,N_20081,N_29963);
xor U38982 (N_38982,N_26390,N_27030);
and U38983 (N_38983,N_21607,N_24436);
nor U38984 (N_38984,N_23298,N_21896);
and U38985 (N_38985,N_28874,N_29891);
nor U38986 (N_38986,N_26750,N_20089);
and U38987 (N_38987,N_28583,N_20917);
xnor U38988 (N_38988,N_29966,N_27261);
and U38989 (N_38989,N_26700,N_26112);
nand U38990 (N_38990,N_21813,N_23296);
or U38991 (N_38991,N_21344,N_29979);
nand U38992 (N_38992,N_22661,N_20072);
xor U38993 (N_38993,N_26374,N_29266);
nand U38994 (N_38994,N_22135,N_24722);
or U38995 (N_38995,N_21079,N_22480);
nor U38996 (N_38996,N_20326,N_29066);
or U38997 (N_38997,N_20794,N_28607);
nand U38998 (N_38998,N_22238,N_21167);
nand U38999 (N_38999,N_23634,N_28680);
or U39000 (N_39000,N_27815,N_25274);
or U39001 (N_39001,N_25604,N_28346);
and U39002 (N_39002,N_23964,N_27471);
nand U39003 (N_39003,N_20375,N_22481);
or U39004 (N_39004,N_21604,N_28696);
and U39005 (N_39005,N_27420,N_25423);
nand U39006 (N_39006,N_23735,N_26234);
xor U39007 (N_39007,N_29129,N_25499);
xnor U39008 (N_39008,N_26653,N_21206);
nand U39009 (N_39009,N_20544,N_20793);
and U39010 (N_39010,N_24634,N_24663);
xor U39011 (N_39011,N_22557,N_26447);
and U39012 (N_39012,N_27381,N_25348);
nor U39013 (N_39013,N_27797,N_24083);
and U39014 (N_39014,N_24255,N_26039);
or U39015 (N_39015,N_21831,N_29299);
xnor U39016 (N_39016,N_28112,N_26546);
nor U39017 (N_39017,N_28338,N_20904);
nand U39018 (N_39018,N_22446,N_23121);
xnor U39019 (N_39019,N_29265,N_23830);
nand U39020 (N_39020,N_22549,N_21815);
and U39021 (N_39021,N_22046,N_20415);
xnor U39022 (N_39022,N_29582,N_27750);
or U39023 (N_39023,N_25685,N_26166);
or U39024 (N_39024,N_22708,N_24327);
nand U39025 (N_39025,N_28969,N_27518);
and U39026 (N_39026,N_25262,N_27470);
xnor U39027 (N_39027,N_27488,N_29100);
nor U39028 (N_39028,N_22902,N_27864);
nand U39029 (N_39029,N_23391,N_24478);
and U39030 (N_39030,N_29149,N_20504);
xor U39031 (N_39031,N_22990,N_25593);
xnor U39032 (N_39032,N_25527,N_27792);
or U39033 (N_39033,N_24333,N_25468);
and U39034 (N_39034,N_22263,N_24179);
xnor U39035 (N_39035,N_24249,N_23698);
and U39036 (N_39036,N_28111,N_24349);
and U39037 (N_39037,N_20457,N_27166);
nor U39038 (N_39038,N_20753,N_25913);
nand U39039 (N_39039,N_29011,N_28629);
and U39040 (N_39040,N_22308,N_20976);
xor U39041 (N_39041,N_26431,N_20650);
and U39042 (N_39042,N_25784,N_24449);
or U39043 (N_39043,N_27776,N_24972);
and U39044 (N_39044,N_26392,N_26302);
nor U39045 (N_39045,N_29331,N_21111);
nand U39046 (N_39046,N_20239,N_28550);
or U39047 (N_39047,N_26501,N_29833);
or U39048 (N_39048,N_21009,N_29103);
xor U39049 (N_39049,N_26930,N_21609);
or U39050 (N_39050,N_24084,N_27637);
xnor U39051 (N_39051,N_22808,N_26140);
xor U39052 (N_39052,N_21260,N_29737);
and U39053 (N_39053,N_27211,N_22958);
and U39054 (N_39054,N_20345,N_28052);
xor U39055 (N_39055,N_27214,N_29905);
nand U39056 (N_39056,N_22455,N_22454);
nand U39057 (N_39057,N_29568,N_21033);
and U39058 (N_39058,N_29890,N_26294);
nor U39059 (N_39059,N_20991,N_23388);
or U39060 (N_39060,N_29460,N_21460);
or U39061 (N_39061,N_22282,N_28482);
or U39062 (N_39062,N_25353,N_25529);
nor U39063 (N_39063,N_29070,N_21742);
or U39064 (N_39064,N_27868,N_20604);
nor U39065 (N_39065,N_28641,N_26475);
xor U39066 (N_39066,N_20070,N_21070);
nand U39067 (N_39067,N_22621,N_29578);
nand U39068 (N_39068,N_22505,N_26826);
xnor U39069 (N_39069,N_25696,N_26927);
nand U39070 (N_39070,N_23985,N_27807);
nor U39071 (N_39071,N_26165,N_20024);
xnor U39072 (N_39072,N_23849,N_27500);
nand U39073 (N_39073,N_27409,N_23555);
nand U39074 (N_39074,N_27896,N_25542);
or U39075 (N_39075,N_25911,N_21347);
nor U39076 (N_39076,N_20468,N_21759);
nor U39077 (N_39077,N_25744,N_28592);
nor U39078 (N_39078,N_20142,N_22637);
xor U39079 (N_39079,N_28308,N_20144);
nand U39080 (N_39080,N_22987,N_29545);
xnor U39081 (N_39081,N_29102,N_22811);
nor U39082 (N_39082,N_22158,N_23981);
nor U39083 (N_39083,N_26186,N_22624);
xnor U39084 (N_39084,N_21931,N_21031);
nand U39085 (N_39085,N_29722,N_21505);
xor U39086 (N_39086,N_27160,N_23967);
or U39087 (N_39087,N_26808,N_23789);
xnor U39088 (N_39088,N_24731,N_21446);
xor U39089 (N_39089,N_26205,N_25751);
nand U39090 (N_39090,N_27101,N_20033);
nor U39091 (N_39091,N_20052,N_25553);
nand U39092 (N_39092,N_24495,N_27306);
xor U39093 (N_39093,N_21779,N_25978);
and U39094 (N_39094,N_20529,N_22178);
or U39095 (N_39095,N_27318,N_26779);
and U39096 (N_39096,N_26746,N_28504);
nand U39097 (N_39097,N_27212,N_28101);
nand U39098 (N_39098,N_20976,N_24133);
xnor U39099 (N_39099,N_21054,N_24833);
and U39100 (N_39100,N_20796,N_29482);
nor U39101 (N_39101,N_22137,N_27440);
xor U39102 (N_39102,N_28079,N_27996);
nor U39103 (N_39103,N_23731,N_26385);
nor U39104 (N_39104,N_26903,N_27447);
nand U39105 (N_39105,N_24715,N_20822);
nor U39106 (N_39106,N_28771,N_23407);
or U39107 (N_39107,N_24950,N_25694);
xnor U39108 (N_39108,N_24689,N_27040);
nand U39109 (N_39109,N_23622,N_27585);
or U39110 (N_39110,N_23710,N_28064);
nand U39111 (N_39111,N_24099,N_27847);
nor U39112 (N_39112,N_21096,N_24698);
nand U39113 (N_39113,N_28963,N_28158);
nor U39114 (N_39114,N_28264,N_29550);
xnor U39115 (N_39115,N_24466,N_21817);
and U39116 (N_39116,N_26545,N_26726);
or U39117 (N_39117,N_21363,N_26178);
nand U39118 (N_39118,N_25074,N_29816);
or U39119 (N_39119,N_25281,N_22580);
or U39120 (N_39120,N_23765,N_22763);
xnor U39121 (N_39121,N_28509,N_27046);
or U39122 (N_39122,N_21545,N_23492);
nand U39123 (N_39123,N_25132,N_27644);
nor U39124 (N_39124,N_23748,N_22682);
nand U39125 (N_39125,N_26925,N_26172);
and U39126 (N_39126,N_21079,N_22993);
and U39127 (N_39127,N_24117,N_29847);
nor U39128 (N_39128,N_24821,N_22391);
or U39129 (N_39129,N_25361,N_26415);
nand U39130 (N_39130,N_22423,N_20773);
and U39131 (N_39131,N_28673,N_24449);
nand U39132 (N_39132,N_26402,N_26318);
and U39133 (N_39133,N_23200,N_23860);
nor U39134 (N_39134,N_24603,N_23404);
xor U39135 (N_39135,N_29424,N_29960);
nand U39136 (N_39136,N_22420,N_29917);
and U39137 (N_39137,N_24982,N_21351);
nand U39138 (N_39138,N_25889,N_24302);
and U39139 (N_39139,N_29772,N_20138);
nand U39140 (N_39140,N_21403,N_29632);
xnor U39141 (N_39141,N_28101,N_28742);
nand U39142 (N_39142,N_22489,N_29505);
and U39143 (N_39143,N_20854,N_24497);
and U39144 (N_39144,N_21913,N_20339);
nor U39145 (N_39145,N_25022,N_21752);
xor U39146 (N_39146,N_20164,N_27621);
nor U39147 (N_39147,N_20867,N_26121);
nand U39148 (N_39148,N_23884,N_27409);
and U39149 (N_39149,N_29816,N_20937);
and U39150 (N_39150,N_24070,N_21840);
xnor U39151 (N_39151,N_23530,N_20521);
xor U39152 (N_39152,N_20027,N_20346);
nor U39153 (N_39153,N_25381,N_28163);
and U39154 (N_39154,N_28440,N_23227);
nor U39155 (N_39155,N_28423,N_25453);
nand U39156 (N_39156,N_25123,N_20420);
or U39157 (N_39157,N_26314,N_25727);
or U39158 (N_39158,N_29725,N_26828);
xor U39159 (N_39159,N_28191,N_20021);
or U39160 (N_39160,N_27462,N_23576);
and U39161 (N_39161,N_27203,N_23491);
or U39162 (N_39162,N_24009,N_28455);
xor U39163 (N_39163,N_22115,N_21070);
xnor U39164 (N_39164,N_24603,N_21736);
and U39165 (N_39165,N_23120,N_25225);
and U39166 (N_39166,N_27660,N_29509);
nor U39167 (N_39167,N_29120,N_23202);
xnor U39168 (N_39168,N_26787,N_20326);
nand U39169 (N_39169,N_24590,N_24561);
nor U39170 (N_39170,N_27122,N_28328);
xor U39171 (N_39171,N_24732,N_26676);
nor U39172 (N_39172,N_26617,N_29521);
and U39173 (N_39173,N_29344,N_21714);
and U39174 (N_39174,N_27733,N_21276);
and U39175 (N_39175,N_28358,N_29490);
xnor U39176 (N_39176,N_23486,N_21984);
nor U39177 (N_39177,N_22798,N_21332);
xnor U39178 (N_39178,N_28837,N_26210);
or U39179 (N_39179,N_23853,N_26538);
and U39180 (N_39180,N_21620,N_23605);
nor U39181 (N_39181,N_25691,N_21269);
xnor U39182 (N_39182,N_22107,N_24278);
nand U39183 (N_39183,N_28737,N_21209);
nor U39184 (N_39184,N_27571,N_20403);
and U39185 (N_39185,N_29645,N_28723);
nand U39186 (N_39186,N_29710,N_20391);
nor U39187 (N_39187,N_25626,N_25389);
xor U39188 (N_39188,N_26844,N_25763);
and U39189 (N_39189,N_25267,N_27148);
or U39190 (N_39190,N_22889,N_20856);
or U39191 (N_39191,N_29468,N_23567);
or U39192 (N_39192,N_23348,N_20032);
xor U39193 (N_39193,N_25356,N_23013);
nor U39194 (N_39194,N_20543,N_20659);
or U39195 (N_39195,N_21369,N_26029);
and U39196 (N_39196,N_26886,N_28778);
and U39197 (N_39197,N_25573,N_24604);
xnor U39198 (N_39198,N_28410,N_20548);
xor U39199 (N_39199,N_29146,N_25623);
nand U39200 (N_39200,N_26517,N_29476);
or U39201 (N_39201,N_25531,N_24513);
and U39202 (N_39202,N_21819,N_28292);
nand U39203 (N_39203,N_26561,N_26714);
or U39204 (N_39204,N_27124,N_25103);
and U39205 (N_39205,N_29719,N_28649);
and U39206 (N_39206,N_27670,N_24025);
nor U39207 (N_39207,N_20055,N_24305);
or U39208 (N_39208,N_23090,N_21148);
nand U39209 (N_39209,N_20463,N_24683);
xor U39210 (N_39210,N_21954,N_24242);
xor U39211 (N_39211,N_20468,N_23209);
nor U39212 (N_39212,N_24446,N_21563);
nor U39213 (N_39213,N_27495,N_28469);
or U39214 (N_39214,N_27499,N_25085);
nand U39215 (N_39215,N_23669,N_25256);
and U39216 (N_39216,N_20193,N_26083);
xnor U39217 (N_39217,N_27863,N_23938);
or U39218 (N_39218,N_28156,N_27315);
or U39219 (N_39219,N_24011,N_22313);
nand U39220 (N_39220,N_22582,N_25213);
xor U39221 (N_39221,N_22417,N_22503);
nand U39222 (N_39222,N_25791,N_27799);
nand U39223 (N_39223,N_27067,N_21819);
xor U39224 (N_39224,N_21250,N_29653);
xnor U39225 (N_39225,N_25647,N_27475);
or U39226 (N_39226,N_24414,N_29076);
and U39227 (N_39227,N_27430,N_28053);
and U39228 (N_39228,N_29858,N_29195);
or U39229 (N_39229,N_24645,N_23447);
nor U39230 (N_39230,N_25445,N_28443);
or U39231 (N_39231,N_29479,N_26082);
nand U39232 (N_39232,N_29043,N_20257);
nand U39233 (N_39233,N_23385,N_21768);
xnor U39234 (N_39234,N_26967,N_26558);
and U39235 (N_39235,N_24833,N_25720);
nor U39236 (N_39236,N_27732,N_28843);
xor U39237 (N_39237,N_25140,N_26591);
xor U39238 (N_39238,N_29885,N_29205);
and U39239 (N_39239,N_24307,N_21614);
nand U39240 (N_39240,N_24093,N_20098);
xor U39241 (N_39241,N_24155,N_28127);
nand U39242 (N_39242,N_24660,N_22772);
nor U39243 (N_39243,N_29551,N_23254);
nand U39244 (N_39244,N_29539,N_26336);
and U39245 (N_39245,N_25201,N_23715);
or U39246 (N_39246,N_20224,N_28992);
nor U39247 (N_39247,N_20108,N_28888);
nand U39248 (N_39248,N_24723,N_25239);
or U39249 (N_39249,N_27067,N_26702);
nand U39250 (N_39250,N_21039,N_21786);
nor U39251 (N_39251,N_26685,N_23389);
nor U39252 (N_39252,N_26742,N_20559);
and U39253 (N_39253,N_26031,N_28731);
and U39254 (N_39254,N_26073,N_21955);
or U39255 (N_39255,N_22522,N_20297);
and U39256 (N_39256,N_29639,N_26619);
or U39257 (N_39257,N_28226,N_23332);
xor U39258 (N_39258,N_22986,N_25825);
or U39259 (N_39259,N_25142,N_21531);
and U39260 (N_39260,N_22027,N_28717);
nor U39261 (N_39261,N_28265,N_28540);
or U39262 (N_39262,N_20046,N_28918);
or U39263 (N_39263,N_20304,N_21567);
nor U39264 (N_39264,N_28476,N_29945);
nor U39265 (N_39265,N_26027,N_25950);
and U39266 (N_39266,N_20980,N_21010);
nor U39267 (N_39267,N_25515,N_29202);
xor U39268 (N_39268,N_26051,N_22090);
nor U39269 (N_39269,N_25226,N_29521);
xor U39270 (N_39270,N_29823,N_24971);
xor U39271 (N_39271,N_21849,N_25257);
nand U39272 (N_39272,N_26087,N_26707);
and U39273 (N_39273,N_25147,N_20307);
nand U39274 (N_39274,N_21529,N_25632);
xnor U39275 (N_39275,N_25360,N_25088);
and U39276 (N_39276,N_22283,N_20044);
or U39277 (N_39277,N_21982,N_24079);
and U39278 (N_39278,N_28916,N_20824);
nand U39279 (N_39279,N_24657,N_20969);
or U39280 (N_39280,N_28411,N_27567);
nand U39281 (N_39281,N_29826,N_29904);
nand U39282 (N_39282,N_29643,N_21691);
nand U39283 (N_39283,N_24196,N_24590);
and U39284 (N_39284,N_20065,N_23824);
or U39285 (N_39285,N_26239,N_21182);
nand U39286 (N_39286,N_23942,N_22426);
nand U39287 (N_39287,N_24754,N_26719);
xnor U39288 (N_39288,N_27494,N_28216);
or U39289 (N_39289,N_25855,N_20558);
nor U39290 (N_39290,N_28569,N_23743);
nor U39291 (N_39291,N_23908,N_20721);
and U39292 (N_39292,N_20819,N_25585);
xor U39293 (N_39293,N_29073,N_24587);
or U39294 (N_39294,N_23089,N_22468);
xnor U39295 (N_39295,N_23747,N_27330);
and U39296 (N_39296,N_29376,N_25022);
and U39297 (N_39297,N_28880,N_23011);
nand U39298 (N_39298,N_27244,N_28307);
or U39299 (N_39299,N_24255,N_28683);
nor U39300 (N_39300,N_27736,N_20248);
or U39301 (N_39301,N_27751,N_22941);
xor U39302 (N_39302,N_25035,N_24744);
nand U39303 (N_39303,N_23377,N_24876);
nand U39304 (N_39304,N_28952,N_27877);
xnor U39305 (N_39305,N_25101,N_22760);
nand U39306 (N_39306,N_20569,N_20798);
xor U39307 (N_39307,N_27584,N_27970);
xor U39308 (N_39308,N_23541,N_27406);
or U39309 (N_39309,N_28340,N_27965);
or U39310 (N_39310,N_20522,N_28102);
and U39311 (N_39311,N_27226,N_24345);
xnor U39312 (N_39312,N_24106,N_24393);
or U39313 (N_39313,N_23223,N_20748);
nand U39314 (N_39314,N_27873,N_28131);
and U39315 (N_39315,N_27324,N_26069);
xnor U39316 (N_39316,N_22163,N_21789);
nand U39317 (N_39317,N_27476,N_20580);
and U39318 (N_39318,N_26289,N_23731);
or U39319 (N_39319,N_26897,N_20828);
nor U39320 (N_39320,N_24594,N_24566);
xor U39321 (N_39321,N_29881,N_25799);
nand U39322 (N_39322,N_28729,N_27671);
xnor U39323 (N_39323,N_27334,N_29545);
nor U39324 (N_39324,N_28771,N_24683);
nand U39325 (N_39325,N_23017,N_20564);
and U39326 (N_39326,N_23261,N_25752);
or U39327 (N_39327,N_25343,N_22431);
or U39328 (N_39328,N_27494,N_25222);
or U39329 (N_39329,N_29666,N_23189);
and U39330 (N_39330,N_23317,N_23868);
xnor U39331 (N_39331,N_21096,N_24679);
xnor U39332 (N_39332,N_22435,N_21534);
xor U39333 (N_39333,N_27816,N_24679);
and U39334 (N_39334,N_28491,N_27015);
and U39335 (N_39335,N_27719,N_23739);
and U39336 (N_39336,N_24623,N_27667);
nor U39337 (N_39337,N_24285,N_24891);
nand U39338 (N_39338,N_24681,N_25737);
or U39339 (N_39339,N_20512,N_29665);
and U39340 (N_39340,N_27515,N_23543);
or U39341 (N_39341,N_28159,N_20783);
xor U39342 (N_39342,N_28372,N_21816);
nand U39343 (N_39343,N_23084,N_24908);
xnor U39344 (N_39344,N_28388,N_23753);
nor U39345 (N_39345,N_28125,N_24432);
nand U39346 (N_39346,N_23331,N_22915);
and U39347 (N_39347,N_28652,N_22487);
xor U39348 (N_39348,N_24564,N_29974);
nand U39349 (N_39349,N_29431,N_24161);
xor U39350 (N_39350,N_29221,N_23951);
nor U39351 (N_39351,N_22736,N_28850);
and U39352 (N_39352,N_28507,N_22951);
nand U39353 (N_39353,N_27401,N_28397);
and U39354 (N_39354,N_26745,N_22985);
or U39355 (N_39355,N_26038,N_23426);
and U39356 (N_39356,N_21982,N_28783);
and U39357 (N_39357,N_28459,N_21587);
and U39358 (N_39358,N_28275,N_28473);
or U39359 (N_39359,N_20818,N_24741);
or U39360 (N_39360,N_22957,N_24733);
nor U39361 (N_39361,N_28081,N_23376);
nor U39362 (N_39362,N_24114,N_28104);
nor U39363 (N_39363,N_27268,N_23716);
or U39364 (N_39364,N_24982,N_25350);
nand U39365 (N_39365,N_20655,N_29582);
and U39366 (N_39366,N_29735,N_28761);
and U39367 (N_39367,N_24503,N_25224);
and U39368 (N_39368,N_28272,N_26747);
and U39369 (N_39369,N_20218,N_25857);
nand U39370 (N_39370,N_29037,N_20295);
xnor U39371 (N_39371,N_22373,N_23402);
nor U39372 (N_39372,N_27227,N_25615);
nor U39373 (N_39373,N_23102,N_20866);
nor U39374 (N_39374,N_23468,N_24560);
and U39375 (N_39375,N_28598,N_25943);
or U39376 (N_39376,N_23957,N_23587);
xor U39377 (N_39377,N_24740,N_28582);
and U39378 (N_39378,N_23749,N_29330);
nor U39379 (N_39379,N_29011,N_29395);
nor U39380 (N_39380,N_29692,N_26112);
nand U39381 (N_39381,N_25290,N_29502);
xnor U39382 (N_39382,N_28069,N_24251);
xnor U39383 (N_39383,N_23588,N_23405);
xor U39384 (N_39384,N_26817,N_23952);
nor U39385 (N_39385,N_21852,N_24464);
nor U39386 (N_39386,N_23239,N_24968);
nor U39387 (N_39387,N_26253,N_29377);
nor U39388 (N_39388,N_22880,N_28383);
nand U39389 (N_39389,N_26999,N_25021);
nand U39390 (N_39390,N_21742,N_28913);
or U39391 (N_39391,N_24017,N_25830);
and U39392 (N_39392,N_27342,N_29934);
xor U39393 (N_39393,N_25192,N_29193);
and U39394 (N_39394,N_21570,N_26162);
nor U39395 (N_39395,N_25948,N_26790);
nand U39396 (N_39396,N_22010,N_27613);
nand U39397 (N_39397,N_26100,N_20666);
nor U39398 (N_39398,N_22742,N_25710);
or U39399 (N_39399,N_24506,N_27867);
and U39400 (N_39400,N_26704,N_21383);
xor U39401 (N_39401,N_27335,N_21332);
or U39402 (N_39402,N_23411,N_26530);
nor U39403 (N_39403,N_20096,N_27652);
xnor U39404 (N_39404,N_25605,N_26874);
nor U39405 (N_39405,N_24312,N_24617);
nor U39406 (N_39406,N_26395,N_22677);
xnor U39407 (N_39407,N_22474,N_20537);
nor U39408 (N_39408,N_26175,N_26615);
nor U39409 (N_39409,N_29371,N_26801);
and U39410 (N_39410,N_26220,N_26094);
nand U39411 (N_39411,N_27739,N_24714);
nand U39412 (N_39412,N_28818,N_21798);
and U39413 (N_39413,N_26433,N_22145);
or U39414 (N_39414,N_29352,N_29705);
nand U39415 (N_39415,N_23896,N_24224);
or U39416 (N_39416,N_24233,N_23390);
nand U39417 (N_39417,N_25157,N_27189);
xor U39418 (N_39418,N_26783,N_25656);
xnor U39419 (N_39419,N_21195,N_29648);
nor U39420 (N_39420,N_24348,N_26801);
nor U39421 (N_39421,N_23900,N_24752);
nand U39422 (N_39422,N_28088,N_23959);
or U39423 (N_39423,N_25107,N_20341);
nand U39424 (N_39424,N_22667,N_29005);
nand U39425 (N_39425,N_21971,N_28353);
xnor U39426 (N_39426,N_27094,N_28851);
xnor U39427 (N_39427,N_28348,N_24461);
xor U39428 (N_39428,N_29724,N_27288);
xnor U39429 (N_39429,N_21842,N_25709);
nand U39430 (N_39430,N_24633,N_20402);
nand U39431 (N_39431,N_21009,N_20953);
or U39432 (N_39432,N_28672,N_29249);
and U39433 (N_39433,N_26885,N_26759);
and U39434 (N_39434,N_25094,N_22500);
nand U39435 (N_39435,N_20648,N_20807);
xnor U39436 (N_39436,N_28229,N_23957);
or U39437 (N_39437,N_23188,N_22258);
or U39438 (N_39438,N_22400,N_26068);
nor U39439 (N_39439,N_22089,N_26054);
or U39440 (N_39440,N_21990,N_28520);
and U39441 (N_39441,N_23793,N_24180);
nand U39442 (N_39442,N_24269,N_24953);
xnor U39443 (N_39443,N_27561,N_22059);
nor U39444 (N_39444,N_23696,N_22549);
and U39445 (N_39445,N_23081,N_29323);
or U39446 (N_39446,N_22100,N_29707);
nor U39447 (N_39447,N_24661,N_27759);
xnor U39448 (N_39448,N_21156,N_20781);
nor U39449 (N_39449,N_22946,N_29670);
nand U39450 (N_39450,N_23637,N_28106);
nor U39451 (N_39451,N_25879,N_27488);
xnor U39452 (N_39452,N_27786,N_22697);
nor U39453 (N_39453,N_21833,N_23102);
or U39454 (N_39454,N_21030,N_21844);
and U39455 (N_39455,N_27905,N_26156);
and U39456 (N_39456,N_29513,N_29019);
xor U39457 (N_39457,N_26843,N_29294);
nor U39458 (N_39458,N_25007,N_23835);
nor U39459 (N_39459,N_21912,N_27591);
xor U39460 (N_39460,N_29930,N_26023);
nor U39461 (N_39461,N_27851,N_21844);
nor U39462 (N_39462,N_28153,N_26412);
xnor U39463 (N_39463,N_25828,N_24506);
or U39464 (N_39464,N_29754,N_23064);
nor U39465 (N_39465,N_29854,N_25145);
nor U39466 (N_39466,N_25389,N_21596);
or U39467 (N_39467,N_21937,N_27640);
nor U39468 (N_39468,N_21070,N_23632);
xor U39469 (N_39469,N_26784,N_28823);
nor U39470 (N_39470,N_22190,N_28238);
or U39471 (N_39471,N_24971,N_26475);
nand U39472 (N_39472,N_24627,N_21756);
and U39473 (N_39473,N_28526,N_25262);
nor U39474 (N_39474,N_26389,N_22534);
nor U39475 (N_39475,N_28164,N_26283);
or U39476 (N_39476,N_29524,N_22056);
or U39477 (N_39477,N_23308,N_29372);
or U39478 (N_39478,N_29365,N_29888);
xor U39479 (N_39479,N_28160,N_20819);
and U39480 (N_39480,N_26648,N_27668);
and U39481 (N_39481,N_29359,N_22339);
xnor U39482 (N_39482,N_20080,N_23818);
xnor U39483 (N_39483,N_21795,N_21683);
nor U39484 (N_39484,N_27583,N_29481);
xnor U39485 (N_39485,N_28941,N_25673);
and U39486 (N_39486,N_29885,N_29175);
nor U39487 (N_39487,N_28014,N_20361);
xor U39488 (N_39488,N_27930,N_23859);
xor U39489 (N_39489,N_24508,N_27117);
xor U39490 (N_39490,N_22106,N_24922);
or U39491 (N_39491,N_22693,N_29957);
nand U39492 (N_39492,N_21964,N_21054);
and U39493 (N_39493,N_22566,N_27621);
or U39494 (N_39494,N_25077,N_21365);
and U39495 (N_39495,N_29040,N_26645);
or U39496 (N_39496,N_25946,N_26032);
nand U39497 (N_39497,N_27832,N_27870);
nand U39498 (N_39498,N_24475,N_23396);
or U39499 (N_39499,N_24779,N_25930);
and U39500 (N_39500,N_25855,N_24967);
nand U39501 (N_39501,N_26734,N_28558);
and U39502 (N_39502,N_28219,N_21898);
and U39503 (N_39503,N_22366,N_26465);
nor U39504 (N_39504,N_28558,N_22427);
and U39505 (N_39505,N_22740,N_27056);
xor U39506 (N_39506,N_21570,N_22291);
nor U39507 (N_39507,N_21757,N_24702);
or U39508 (N_39508,N_27889,N_27663);
and U39509 (N_39509,N_20372,N_28177);
nand U39510 (N_39510,N_29237,N_20205);
nand U39511 (N_39511,N_29709,N_25593);
and U39512 (N_39512,N_25941,N_24489);
or U39513 (N_39513,N_22488,N_29783);
nor U39514 (N_39514,N_27544,N_29498);
or U39515 (N_39515,N_20472,N_28315);
nor U39516 (N_39516,N_24104,N_27115);
and U39517 (N_39517,N_26220,N_22407);
and U39518 (N_39518,N_28309,N_24521);
nand U39519 (N_39519,N_22120,N_29346);
xnor U39520 (N_39520,N_28320,N_24600);
and U39521 (N_39521,N_24595,N_23816);
and U39522 (N_39522,N_23702,N_29966);
nor U39523 (N_39523,N_28125,N_21730);
nand U39524 (N_39524,N_21575,N_26127);
or U39525 (N_39525,N_20631,N_21900);
nor U39526 (N_39526,N_24471,N_24295);
nand U39527 (N_39527,N_20617,N_27873);
xnor U39528 (N_39528,N_26844,N_22563);
xnor U39529 (N_39529,N_21697,N_22556);
or U39530 (N_39530,N_22138,N_20009);
and U39531 (N_39531,N_27643,N_22126);
nand U39532 (N_39532,N_29611,N_22714);
xnor U39533 (N_39533,N_20741,N_26447);
and U39534 (N_39534,N_20683,N_25385);
xnor U39535 (N_39535,N_29035,N_23293);
or U39536 (N_39536,N_21973,N_21430);
xnor U39537 (N_39537,N_24009,N_27592);
or U39538 (N_39538,N_28933,N_24053);
xor U39539 (N_39539,N_21672,N_25556);
and U39540 (N_39540,N_29754,N_21998);
xor U39541 (N_39541,N_28290,N_26837);
and U39542 (N_39542,N_20462,N_28591);
nor U39543 (N_39543,N_27169,N_23460);
and U39544 (N_39544,N_25663,N_27219);
or U39545 (N_39545,N_27511,N_26863);
nor U39546 (N_39546,N_29663,N_26211);
or U39547 (N_39547,N_26292,N_20138);
and U39548 (N_39548,N_29180,N_26438);
or U39549 (N_39549,N_28998,N_27307);
nand U39550 (N_39550,N_21138,N_23720);
xor U39551 (N_39551,N_25425,N_25095);
and U39552 (N_39552,N_22493,N_20070);
and U39553 (N_39553,N_20181,N_29348);
and U39554 (N_39554,N_27185,N_20546);
xnor U39555 (N_39555,N_22277,N_20585);
or U39556 (N_39556,N_28341,N_22806);
nand U39557 (N_39557,N_27620,N_21652);
and U39558 (N_39558,N_25804,N_20943);
nand U39559 (N_39559,N_29715,N_21203);
and U39560 (N_39560,N_26232,N_21411);
and U39561 (N_39561,N_22241,N_22353);
nand U39562 (N_39562,N_21689,N_22707);
or U39563 (N_39563,N_21985,N_26668);
nor U39564 (N_39564,N_23939,N_24386);
nor U39565 (N_39565,N_24468,N_21612);
or U39566 (N_39566,N_25869,N_25270);
or U39567 (N_39567,N_24042,N_28399);
nand U39568 (N_39568,N_26007,N_22161);
xnor U39569 (N_39569,N_26805,N_26712);
nor U39570 (N_39570,N_24702,N_28936);
and U39571 (N_39571,N_21959,N_24827);
xor U39572 (N_39572,N_24999,N_21943);
nand U39573 (N_39573,N_23726,N_29730);
or U39574 (N_39574,N_23827,N_20621);
nand U39575 (N_39575,N_23813,N_23197);
and U39576 (N_39576,N_29554,N_25436);
and U39577 (N_39577,N_20875,N_28131);
nor U39578 (N_39578,N_24949,N_23798);
nand U39579 (N_39579,N_20452,N_29939);
or U39580 (N_39580,N_27939,N_29500);
xor U39581 (N_39581,N_29113,N_22779);
nand U39582 (N_39582,N_24411,N_21993);
nand U39583 (N_39583,N_20392,N_22109);
or U39584 (N_39584,N_24431,N_27136);
and U39585 (N_39585,N_25331,N_20690);
and U39586 (N_39586,N_28970,N_21739);
and U39587 (N_39587,N_28569,N_20139);
or U39588 (N_39588,N_26925,N_24811);
and U39589 (N_39589,N_21979,N_27244);
and U39590 (N_39590,N_21047,N_22739);
nor U39591 (N_39591,N_23261,N_28993);
nor U39592 (N_39592,N_20620,N_28225);
nor U39593 (N_39593,N_21974,N_27703);
xnor U39594 (N_39594,N_27642,N_26803);
nand U39595 (N_39595,N_23394,N_28513);
and U39596 (N_39596,N_23290,N_29674);
xnor U39597 (N_39597,N_22182,N_29883);
xor U39598 (N_39598,N_29997,N_24393);
nand U39599 (N_39599,N_25556,N_22773);
nand U39600 (N_39600,N_23217,N_20567);
xnor U39601 (N_39601,N_28324,N_27171);
nand U39602 (N_39602,N_26585,N_26242);
and U39603 (N_39603,N_22752,N_21595);
and U39604 (N_39604,N_29046,N_29444);
nand U39605 (N_39605,N_22953,N_24645);
xnor U39606 (N_39606,N_27292,N_22468);
xnor U39607 (N_39607,N_26825,N_20370);
xor U39608 (N_39608,N_28053,N_26030);
nand U39609 (N_39609,N_26150,N_29215);
nor U39610 (N_39610,N_29514,N_27869);
nor U39611 (N_39611,N_20555,N_20916);
nor U39612 (N_39612,N_24431,N_21854);
xor U39613 (N_39613,N_26803,N_29944);
xnor U39614 (N_39614,N_28136,N_21380);
xor U39615 (N_39615,N_28527,N_27287);
nor U39616 (N_39616,N_23373,N_21916);
and U39617 (N_39617,N_21943,N_21324);
and U39618 (N_39618,N_25377,N_25412);
nand U39619 (N_39619,N_24125,N_23228);
nor U39620 (N_39620,N_25104,N_20639);
xor U39621 (N_39621,N_26918,N_24111);
or U39622 (N_39622,N_22084,N_21835);
or U39623 (N_39623,N_20375,N_25456);
nor U39624 (N_39624,N_22202,N_27792);
and U39625 (N_39625,N_27126,N_23957);
and U39626 (N_39626,N_26398,N_22606);
xor U39627 (N_39627,N_20093,N_21879);
nand U39628 (N_39628,N_29046,N_28900);
nor U39629 (N_39629,N_20811,N_26806);
or U39630 (N_39630,N_22185,N_29918);
nor U39631 (N_39631,N_29653,N_21200);
nand U39632 (N_39632,N_25196,N_25046);
and U39633 (N_39633,N_24361,N_26748);
nor U39634 (N_39634,N_22763,N_20199);
or U39635 (N_39635,N_29792,N_23995);
nor U39636 (N_39636,N_22565,N_28181);
or U39637 (N_39637,N_24501,N_28315);
and U39638 (N_39638,N_24314,N_24988);
nor U39639 (N_39639,N_27664,N_23808);
nand U39640 (N_39640,N_22564,N_22973);
nand U39641 (N_39641,N_27616,N_20588);
xor U39642 (N_39642,N_22712,N_20113);
or U39643 (N_39643,N_20297,N_28641);
nand U39644 (N_39644,N_26063,N_24841);
xor U39645 (N_39645,N_23090,N_25147);
nor U39646 (N_39646,N_25364,N_21389);
nand U39647 (N_39647,N_21874,N_28967);
nand U39648 (N_39648,N_23984,N_23634);
or U39649 (N_39649,N_24788,N_23197);
xnor U39650 (N_39650,N_27033,N_23690);
and U39651 (N_39651,N_20595,N_24347);
and U39652 (N_39652,N_20434,N_21316);
nand U39653 (N_39653,N_22185,N_23027);
or U39654 (N_39654,N_22466,N_22019);
nand U39655 (N_39655,N_22126,N_27924);
nand U39656 (N_39656,N_20456,N_20776);
and U39657 (N_39657,N_20071,N_25498);
nor U39658 (N_39658,N_22869,N_29474);
or U39659 (N_39659,N_20596,N_28444);
and U39660 (N_39660,N_24725,N_20890);
nand U39661 (N_39661,N_22019,N_27230);
or U39662 (N_39662,N_28030,N_25644);
or U39663 (N_39663,N_23976,N_22122);
or U39664 (N_39664,N_23617,N_25104);
xor U39665 (N_39665,N_26459,N_25597);
nor U39666 (N_39666,N_24343,N_29174);
nand U39667 (N_39667,N_25187,N_23234);
or U39668 (N_39668,N_29618,N_26841);
xnor U39669 (N_39669,N_29230,N_25350);
or U39670 (N_39670,N_25155,N_25527);
nor U39671 (N_39671,N_20472,N_26985);
xor U39672 (N_39672,N_26354,N_29354);
and U39673 (N_39673,N_26710,N_23942);
or U39674 (N_39674,N_25093,N_20246);
nor U39675 (N_39675,N_29596,N_28350);
or U39676 (N_39676,N_21848,N_22020);
nor U39677 (N_39677,N_23052,N_25841);
nand U39678 (N_39678,N_20893,N_21901);
xor U39679 (N_39679,N_28128,N_20934);
nand U39680 (N_39680,N_22180,N_27078);
xnor U39681 (N_39681,N_23747,N_21727);
xor U39682 (N_39682,N_24966,N_23212);
nand U39683 (N_39683,N_26609,N_26531);
nand U39684 (N_39684,N_29639,N_29120);
or U39685 (N_39685,N_24909,N_25259);
xnor U39686 (N_39686,N_22575,N_21071);
or U39687 (N_39687,N_28780,N_22225);
xnor U39688 (N_39688,N_28288,N_20974);
xnor U39689 (N_39689,N_24013,N_21262);
or U39690 (N_39690,N_26895,N_20514);
nand U39691 (N_39691,N_29393,N_22921);
xor U39692 (N_39692,N_27766,N_23195);
nor U39693 (N_39693,N_27857,N_24855);
nor U39694 (N_39694,N_21534,N_25722);
xnor U39695 (N_39695,N_26304,N_26089);
or U39696 (N_39696,N_26306,N_22347);
nand U39697 (N_39697,N_21395,N_28053);
xor U39698 (N_39698,N_20685,N_20882);
nand U39699 (N_39699,N_28096,N_23317);
and U39700 (N_39700,N_20842,N_21082);
or U39701 (N_39701,N_23508,N_26981);
nand U39702 (N_39702,N_23311,N_28807);
and U39703 (N_39703,N_25151,N_27064);
nor U39704 (N_39704,N_25026,N_26090);
or U39705 (N_39705,N_21281,N_20802);
or U39706 (N_39706,N_26750,N_29444);
and U39707 (N_39707,N_29663,N_25793);
or U39708 (N_39708,N_26503,N_20719);
and U39709 (N_39709,N_24572,N_27877);
nor U39710 (N_39710,N_27535,N_24225);
nor U39711 (N_39711,N_27310,N_23265);
nand U39712 (N_39712,N_20510,N_24272);
or U39713 (N_39713,N_21421,N_27482);
and U39714 (N_39714,N_20036,N_20871);
nor U39715 (N_39715,N_24102,N_23209);
and U39716 (N_39716,N_27444,N_22579);
and U39717 (N_39717,N_20740,N_25995);
nand U39718 (N_39718,N_21554,N_29398);
or U39719 (N_39719,N_25889,N_23141);
xor U39720 (N_39720,N_23257,N_26577);
xor U39721 (N_39721,N_29347,N_26861);
nand U39722 (N_39722,N_23963,N_20763);
nor U39723 (N_39723,N_26639,N_24833);
or U39724 (N_39724,N_26561,N_23138);
and U39725 (N_39725,N_21403,N_22982);
or U39726 (N_39726,N_24491,N_21489);
and U39727 (N_39727,N_22092,N_25701);
nand U39728 (N_39728,N_20982,N_25731);
and U39729 (N_39729,N_22647,N_26915);
nor U39730 (N_39730,N_24184,N_28785);
or U39731 (N_39731,N_29412,N_20998);
and U39732 (N_39732,N_20224,N_23009);
nor U39733 (N_39733,N_21797,N_23046);
and U39734 (N_39734,N_22398,N_29539);
nor U39735 (N_39735,N_27052,N_24892);
nor U39736 (N_39736,N_25267,N_20780);
xnor U39737 (N_39737,N_26794,N_29984);
or U39738 (N_39738,N_25635,N_23354);
xor U39739 (N_39739,N_20242,N_26767);
nand U39740 (N_39740,N_20624,N_23776);
nand U39741 (N_39741,N_25178,N_22967);
xnor U39742 (N_39742,N_26318,N_21466);
or U39743 (N_39743,N_21484,N_24964);
or U39744 (N_39744,N_23549,N_20265);
nor U39745 (N_39745,N_27295,N_24764);
or U39746 (N_39746,N_22118,N_28417);
or U39747 (N_39747,N_20960,N_25626);
and U39748 (N_39748,N_23360,N_26910);
or U39749 (N_39749,N_27762,N_23875);
xor U39750 (N_39750,N_22560,N_29182);
and U39751 (N_39751,N_24101,N_22944);
nand U39752 (N_39752,N_21009,N_24828);
nor U39753 (N_39753,N_25677,N_20794);
xnor U39754 (N_39754,N_22229,N_26268);
and U39755 (N_39755,N_25415,N_24997);
nand U39756 (N_39756,N_20929,N_27444);
and U39757 (N_39757,N_27611,N_29707);
nand U39758 (N_39758,N_28211,N_25721);
nor U39759 (N_39759,N_29172,N_23844);
and U39760 (N_39760,N_20135,N_29861);
xor U39761 (N_39761,N_24173,N_26315);
or U39762 (N_39762,N_29332,N_23403);
nand U39763 (N_39763,N_22046,N_27753);
and U39764 (N_39764,N_21170,N_28207);
and U39765 (N_39765,N_29402,N_29696);
nand U39766 (N_39766,N_22821,N_26453);
or U39767 (N_39767,N_24335,N_25075);
nand U39768 (N_39768,N_29401,N_25790);
xor U39769 (N_39769,N_24899,N_21420);
xor U39770 (N_39770,N_28629,N_26890);
nand U39771 (N_39771,N_20401,N_22776);
nand U39772 (N_39772,N_27195,N_27272);
xnor U39773 (N_39773,N_24231,N_24187);
nor U39774 (N_39774,N_27950,N_21419);
nor U39775 (N_39775,N_20839,N_28546);
and U39776 (N_39776,N_25780,N_27882);
nor U39777 (N_39777,N_23082,N_21132);
nor U39778 (N_39778,N_27380,N_20630);
and U39779 (N_39779,N_29303,N_24847);
or U39780 (N_39780,N_28208,N_27698);
nand U39781 (N_39781,N_28604,N_26529);
or U39782 (N_39782,N_27227,N_20285);
xor U39783 (N_39783,N_24452,N_21131);
xor U39784 (N_39784,N_26447,N_29521);
nand U39785 (N_39785,N_28211,N_21137);
and U39786 (N_39786,N_20830,N_26646);
or U39787 (N_39787,N_24689,N_26878);
and U39788 (N_39788,N_26118,N_21825);
or U39789 (N_39789,N_27994,N_23397);
and U39790 (N_39790,N_24084,N_27182);
or U39791 (N_39791,N_20854,N_26911);
nand U39792 (N_39792,N_26167,N_28999);
nor U39793 (N_39793,N_26264,N_20819);
nand U39794 (N_39794,N_23445,N_24142);
and U39795 (N_39795,N_27107,N_24657);
nand U39796 (N_39796,N_29400,N_29155);
and U39797 (N_39797,N_29108,N_23110);
or U39798 (N_39798,N_25478,N_26776);
xnor U39799 (N_39799,N_25511,N_27525);
and U39800 (N_39800,N_26800,N_29560);
or U39801 (N_39801,N_29351,N_25293);
or U39802 (N_39802,N_22382,N_24849);
nand U39803 (N_39803,N_27570,N_24460);
nor U39804 (N_39804,N_29996,N_28285);
or U39805 (N_39805,N_24771,N_26719);
nand U39806 (N_39806,N_28328,N_20192);
nand U39807 (N_39807,N_24309,N_27692);
and U39808 (N_39808,N_23911,N_28403);
nor U39809 (N_39809,N_22208,N_29940);
or U39810 (N_39810,N_28567,N_28366);
xor U39811 (N_39811,N_24743,N_21348);
or U39812 (N_39812,N_24054,N_20512);
nand U39813 (N_39813,N_22396,N_22128);
nor U39814 (N_39814,N_21941,N_23532);
and U39815 (N_39815,N_29813,N_29715);
xor U39816 (N_39816,N_23755,N_28578);
nor U39817 (N_39817,N_24862,N_22667);
or U39818 (N_39818,N_25565,N_22297);
or U39819 (N_39819,N_27492,N_22812);
and U39820 (N_39820,N_24581,N_29368);
and U39821 (N_39821,N_22557,N_22001);
nand U39822 (N_39822,N_28759,N_21946);
xnor U39823 (N_39823,N_27379,N_22012);
and U39824 (N_39824,N_28325,N_25339);
nand U39825 (N_39825,N_22488,N_29251);
xor U39826 (N_39826,N_26982,N_25158);
nand U39827 (N_39827,N_27722,N_21100);
nand U39828 (N_39828,N_25045,N_27477);
xnor U39829 (N_39829,N_26017,N_26639);
nor U39830 (N_39830,N_22679,N_26765);
or U39831 (N_39831,N_23958,N_26120);
and U39832 (N_39832,N_24076,N_27015);
or U39833 (N_39833,N_23264,N_29640);
nor U39834 (N_39834,N_23514,N_21749);
and U39835 (N_39835,N_22265,N_24691);
nand U39836 (N_39836,N_28093,N_24494);
and U39837 (N_39837,N_23861,N_25787);
nor U39838 (N_39838,N_24245,N_25975);
xor U39839 (N_39839,N_26599,N_21979);
nor U39840 (N_39840,N_28695,N_21672);
and U39841 (N_39841,N_25431,N_27802);
nor U39842 (N_39842,N_26272,N_23572);
xor U39843 (N_39843,N_20701,N_26671);
nand U39844 (N_39844,N_28713,N_22202);
nor U39845 (N_39845,N_27513,N_22257);
xnor U39846 (N_39846,N_25017,N_23234);
nand U39847 (N_39847,N_26325,N_27126);
or U39848 (N_39848,N_20319,N_27467);
nand U39849 (N_39849,N_28973,N_20284);
and U39850 (N_39850,N_26859,N_25108);
nor U39851 (N_39851,N_28335,N_22247);
xor U39852 (N_39852,N_26501,N_28438);
or U39853 (N_39853,N_27348,N_20334);
and U39854 (N_39854,N_25208,N_22460);
and U39855 (N_39855,N_28656,N_25503);
nor U39856 (N_39856,N_27197,N_26488);
nand U39857 (N_39857,N_27576,N_26445);
xor U39858 (N_39858,N_28780,N_26052);
and U39859 (N_39859,N_29621,N_29523);
nand U39860 (N_39860,N_27726,N_23777);
xor U39861 (N_39861,N_25814,N_22953);
or U39862 (N_39862,N_25984,N_27939);
or U39863 (N_39863,N_22651,N_29589);
nand U39864 (N_39864,N_24049,N_28000);
or U39865 (N_39865,N_28036,N_26892);
nand U39866 (N_39866,N_23427,N_22143);
nor U39867 (N_39867,N_21632,N_27564);
nor U39868 (N_39868,N_29932,N_23048);
or U39869 (N_39869,N_22971,N_20467);
nor U39870 (N_39870,N_23794,N_29808);
or U39871 (N_39871,N_28121,N_25484);
or U39872 (N_39872,N_25215,N_22600);
xnor U39873 (N_39873,N_28933,N_20535);
nand U39874 (N_39874,N_21145,N_23216);
nor U39875 (N_39875,N_21144,N_22731);
and U39876 (N_39876,N_20464,N_29898);
nand U39877 (N_39877,N_29566,N_29034);
or U39878 (N_39878,N_23004,N_22929);
nand U39879 (N_39879,N_24876,N_21848);
xnor U39880 (N_39880,N_20641,N_29864);
nand U39881 (N_39881,N_29436,N_24412);
nor U39882 (N_39882,N_22800,N_27937);
or U39883 (N_39883,N_20950,N_21249);
nand U39884 (N_39884,N_23585,N_22461);
nand U39885 (N_39885,N_21924,N_27810);
xnor U39886 (N_39886,N_23752,N_27567);
nand U39887 (N_39887,N_28282,N_23252);
and U39888 (N_39888,N_20410,N_20441);
or U39889 (N_39889,N_27990,N_25630);
and U39890 (N_39890,N_26077,N_20077);
xnor U39891 (N_39891,N_29012,N_27242);
nand U39892 (N_39892,N_26400,N_22007);
nand U39893 (N_39893,N_20635,N_24041);
nor U39894 (N_39894,N_29428,N_26172);
and U39895 (N_39895,N_25013,N_20708);
and U39896 (N_39896,N_21980,N_28826);
or U39897 (N_39897,N_27259,N_24268);
nor U39898 (N_39898,N_29210,N_20252);
and U39899 (N_39899,N_24074,N_27907);
xor U39900 (N_39900,N_28824,N_22263);
nand U39901 (N_39901,N_28637,N_25473);
xor U39902 (N_39902,N_28484,N_28458);
xor U39903 (N_39903,N_27666,N_27490);
nor U39904 (N_39904,N_24716,N_22763);
and U39905 (N_39905,N_27250,N_22040);
nor U39906 (N_39906,N_23638,N_20643);
xnor U39907 (N_39907,N_27585,N_26706);
xnor U39908 (N_39908,N_25685,N_28976);
nor U39909 (N_39909,N_23365,N_27340);
nor U39910 (N_39910,N_23361,N_23076);
nor U39911 (N_39911,N_22796,N_29475);
nor U39912 (N_39912,N_26943,N_29158);
nand U39913 (N_39913,N_28443,N_23530);
xnor U39914 (N_39914,N_22443,N_26709);
nand U39915 (N_39915,N_21867,N_20226);
and U39916 (N_39916,N_22739,N_23238);
nand U39917 (N_39917,N_25525,N_24538);
xor U39918 (N_39918,N_23380,N_22585);
xor U39919 (N_39919,N_29288,N_29584);
nor U39920 (N_39920,N_22082,N_29030);
nand U39921 (N_39921,N_29761,N_20696);
xnor U39922 (N_39922,N_26200,N_24312);
or U39923 (N_39923,N_29769,N_21297);
nand U39924 (N_39924,N_28864,N_25133);
nand U39925 (N_39925,N_26522,N_24711);
nor U39926 (N_39926,N_28367,N_26713);
nand U39927 (N_39927,N_25255,N_24401);
or U39928 (N_39928,N_25486,N_23707);
xor U39929 (N_39929,N_20514,N_26944);
nor U39930 (N_39930,N_25230,N_20376);
xnor U39931 (N_39931,N_29091,N_22298);
and U39932 (N_39932,N_28382,N_24764);
xor U39933 (N_39933,N_24837,N_29627);
nand U39934 (N_39934,N_28387,N_25561);
and U39935 (N_39935,N_23607,N_21094);
nand U39936 (N_39936,N_29341,N_28149);
and U39937 (N_39937,N_25789,N_22251);
xor U39938 (N_39938,N_26426,N_24469);
nor U39939 (N_39939,N_21523,N_21735);
nor U39940 (N_39940,N_22099,N_20319);
and U39941 (N_39941,N_29719,N_25470);
nand U39942 (N_39942,N_21930,N_27260);
or U39943 (N_39943,N_21624,N_27717);
and U39944 (N_39944,N_26610,N_26145);
xor U39945 (N_39945,N_20460,N_23789);
or U39946 (N_39946,N_22141,N_28374);
or U39947 (N_39947,N_22827,N_29974);
nand U39948 (N_39948,N_23870,N_23387);
nor U39949 (N_39949,N_29124,N_29712);
xor U39950 (N_39950,N_23939,N_27651);
or U39951 (N_39951,N_25927,N_23268);
xnor U39952 (N_39952,N_27095,N_21679);
nor U39953 (N_39953,N_29521,N_22317);
nand U39954 (N_39954,N_23708,N_21272);
nor U39955 (N_39955,N_24954,N_21719);
nor U39956 (N_39956,N_27714,N_23697);
nor U39957 (N_39957,N_27142,N_22991);
and U39958 (N_39958,N_25574,N_27775);
and U39959 (N_39959,N_20995,N_22794);
xor U39960 (N_39960,N_25315,N_25183);
xnor U39961 (N_39961,N_23902,N_21247);
nor U39962 (N_39962,N_26607,N_29520);
or U39963 (N_39963,N_26943,N_28090);
and U39964 (N_39964,N_20794,N_22955);
nand U39965 (N_39965,N_26704,N_20321);
nand U39966 (N_39966,N_29600,N_20066);
nand U39967 (N_39967,N_28370,N_20532);
nor U39968 (N_39968,N_23715,N_20011);
nand U39969 (N_39969,N_25581,N_29780);
or U39970 (N_39970,N_25900,N_23579);
and U39971 (N_39971,N_27699,N_29651);
nand U39972 (N_39972,N_25669,N_23000);
nor U39973 (N_39973,N_20062,N_22124);
nor U39974 (N_39974,N_28426,N_24494);
nand U39975 (N_39975,N_29555,N_26669);
or U39976 (N_39976,N_26409,N_26615);
nor U39977 (N_39977,N_28891,N_26055);
or U39978 (N_39978,N_25707,N_27662);
nand U39979 (N_39979,N_22186,N_23008);
nor U39980 (N_39980,N_25542,N_21328);
xor U39981 (N_39981,N_28277,N_23081);
or U39982 (N_39982,N_29923,N_24916);
or U39983 (N_39983,N_21562,N_20003);
nor U39984 (N_39984,N_29723,N_27150);
or U39985 (N_39985,N_21678,N_20875);
or U39986 (N_39986,N_24602,N_22784);
nand U39987 (N_39987,N_22716,N_24018);
or U39988 (N_39988,N_29851,N_20992);
and U39989 (N_39989,N_23012,N_23152);
xnor U39990 (N_39990,N_25483,N_25162);
or U39991 (N_39991,N_27830,N_20705);
or U39992 (N_39992,N_26438,N_27134);
xnor U39993 (N_39993,N_20434,N_28959);
xnor U39994 (N_39994,N_26415,N_26501);
and U39995 (N_39995,N_23204,N_21313);
nand U39996 (N_39996,N_20902,N_24113);
xor U39997 (N_39997,N_26204,N_23763);
nor U39998 (N_39998,N_21552,N_20043);
xor U39999 (N_39999,N_23151,N_24699);
nor U40000 (N_40000,N_37217,N_34655);
nand U40001 (N_40001,N_37639,N_35896);
and U40002 (N_40002,N_32367,N_38905);
nor U40003 (N_40003,N_36584,N_30780);
nand U40004 (N_40004,N_37935,N_39725);
nand U40005 (N_40005,N_32719,N_37010);
and U40006 (N_40006,N_37230,N_33840);
and U40007 (N_40007,N_38335,N_39743);
or U40008 (N_40008,N_32754,N_37906);
xor U40009 (N_40009,N_30464,N_33912);
and U40010 (N_40010,N_34746,N_30539);
or U40011 (N_40011,N_30666,N_38555);
xnor U40012 (N_40012,N_31218,N_34649);
xnor U40013 (N_40013,N_37018,N_34749);
and U40014 (N_40014,N_39051,N_37489);
or U40015 (N_40015,N_31197,N_39888);
nor U40016 (N_40016,N_37396,N_30579);
or U40017 (N_40017,N_38969,N_39169);
or U40018 (N_40018,N_35143,N_34105);
or U40019 (N_40019,N_32368,N_38250);
and U40020 (N_40020,N_35408,N_39625);
and U40021 (N_40021,N_37290,N_36336);
nand U40022 (N_40022,N_38971,N_31789);
xor U40023 (N_40023,N_33195,N_39635);
xor U40024 (N_40024,N_32912,N_31834);
xor U40025 (N_40025,N_38168,N_34834);
nor U40026 (N_40026,N_39052,N_38289);
or U40027 (N_40027,N_35085,N_38554);
nor U40028 (N_40028,N_37667,N_30167);
nand U40029 (N_40029,N_37644,N_30014);
nand U40030 (N_40030,N_37839,N_31132);
and U40031 (N_40031,N_33859,N_34221);
nand U40032 (N_40032,N_30067,N_37674);
nor U40033 (N_40033,N_34621,N_34230);
nand U40034 (N_40034,N_32493,N_31100);
and U40035 (N_40035,N_34522,N_37712);
nand U40036 (N_40036,N_39742,N_34499);
and U40037 (N_40037,N_30542,N_37573);
or U40038 (N_40038,N_33801,N_34155);
nand U40039 (N_40039,N_39066,N_30981);
and U40040 (N_40040,N_36847,N_36359);
nor U40041 (N_40041,N_33678,N_32560);
nand U40042 (N_40042,N_36196,N_30081);
and U40043 (N_40043,N_36451,N_31252);
or U40044 (N_40044,N_34757,N_38410);
nor U40045 (N_40045,N_38677,N_39445);
nand U40046 (N_40046,N_31783,N_37410);
nor U40047 (N_40047,N_37778,N_35199);
or U40048 (N_40048,N_37232,N_30468);
xor U40049 (N_40049,N_30752,N_36758);
nand U40050 (N_40050,N_38286,N_31026);
nand U40051 (N_40051,N_30737,N_39688);
or U40052 (N_40052,N_30144,N_34139);
and U40053 (N_40053,N_36787,N_37685);
or U40054 (N_40054,N_34058,N_34466);
nor U40055 (N_40055,N_36820,N_37451);
nor U40056 (N_40056,N_35994,N_32242);
and U40057 (N_40057,N_33651,N_31155);
nor U40058 (N_40058,N_31045,N_34001);
or U40059 (N_40059,N_37274,N_34955);
and U40060 (N_40060,N_34212,N_39538);
xor U40061 (N_40061,N_31751,N_37769);
nand U40062 (N_40062,N_33622,N_38644);
nand U40063 (N_40063,N_34358,N_38029);
xor U40064 (N_40064,N_31950,N_33380);
nor U40065 (N_40065,N_35126,N_33969);
and U40066 (N_40066,N_31562,N_35490);
and U40067 (N_40067,N_33100,N_39557);
nor U40068 (N_40068,N_38017,N_37606);
nor U40069 (N_40069,N_31978,N_35277);
nor U40070 (N_40070,N_38489,N_31015);
nor U40071 (N_40071,N_33992,N_36323);
nand U40072 (N_40072,N_35236,N_38453);
nor U40073 (N_40073,N_34280,N_33728);
and U40074 (N_40074,N_36025,N_33844);
xor U40075 (N_40075,N_30746,N_35892);
nor U40076 (N_40076,N_31047,N_35501);
xnor U40077 (N_40077,N_37428,N_35843);
nand U40078 (N_40078,N_36339,N_32557);
nand U40079 (N_40079,N_32096,N_33021);
and U40080 (N_40080,N_31354,N_39010);
or U40081 (N_40081,N_35433,N_38692);
nand U40082 (N_40082,N_30732,N_34100);
nand U40083 (N_40083,N_36666,N_33817);
nor U40084 (N_40084,N_35938,N_38902);
nand U40085 (N_40085,N_34448,N_38237);
xor U40086 (N_40086,N_39457,N_32530);
nand U40087 (N_40087,N_38239,N_38573);
nor U40088 (N_40088,N_30553,N_35806);
xnor U40089 (N_40089,N_30215,N_34332);
or U40090 (N_40090,N_30300,N_38257);
and U40091 (N_40091,N_37122,N_38356);
nand U40092 (N_40092,N_35731,N_33299);
nor U40093 (N_40093,N_35178,N_36059);
and U40094 (N_40094,N_32948,N_31678);
nor U40095 (N_40095,N_33115,N_33846);
or U40096 (N_40096,N_35937,N_32720);
and U40097 (N_40097,N_35627,N_37137);
or U40098 (N_40098,N_38024,N_31305);
nand U40099 (N_40099,N_34079,N_36718);
nor U40100 (N_40100,N_35726,N_39816);
or U40101 (N_40101,N_33883,N_32108);
and U40102 (N_40102,N_34496,N_33691);
nor U40103 (N_40103,N_33194,N_37724);
xnor U40104 (N_40104,N_34939,N_37790);
nor U40105 (N_40105,N_37206,N_39166);
nand U40106 (N_40106,N_39153,N_30816);
and U40107 (N_40107,N_38996,N_39098);
and U40108 (N_40108,N_39988,N_31530);
or U40109 (N_40109,N_31752,N_39879);
nand U40110 (N_40110,N_36511,N_35593);
nand U40111 (N_40111,N_30622,N_36976);
nand U40112 (N_40112,N_33874,N_34441);
or U40113 (N_40113,N_38082,N_35405);
nand U40114 (N_40114,N_32224,N_31502);
xor U40115 (N_40115,N_32992,N_32799);
nand U40116 (N_40116,N_31692,N_31193);
nand U40117 (N_40117,N_36414,N_38044);
xnor U40118 (N_40118,N_31005,N_31478);
or U40119 (N_40119,N_33759,N_30690);
and U40120 (N_40120,N_34866,N_38426);
or U40121 (N_40121,N_39399,N_36089);
nand U40122 (N_40122,N_36002,N_34098);
nand U40123 (N_40123,N_32322,N_36320);
and U40124 (N_40124,N_38772,N_35132);
xor U40125 (N_40125,N_32478,N_38682);
nor U40126 (N_40126,N_38213,N_33825);
and U40127 (N_40127,N_31027,N_39017);
or U40128 (N_40128,N_31420,N_33960);
and U40129 (N_40129,N_35929,N_37710);
or U40130 (N_40130,N_39281,N_39152);
and U40131 (N_40131,N_30580,N_33008);
nand U40132 (N_40132,N_35309,N_34384);
xnor U40133 (N_40133,N_38469,N_31779);
xnor U40134 (N_40134,N_31724,N_38538);
or U40135 (N_40135,N_34899,N_39055);
and U40136 (N_40136,N_39383,N_35391);
nor U40137 (N_40137,N_39817,N_32731);
or U40138 (N_40138,N_38976,N_38652);
nor U40139 (N_40139,N_39220,N_39539);
or U40140 (N_40140,N_34524,N_37093);
nand U40141 (N_40141,N_36113,N_33548);
and U40142 (N_40142,N_38157,N_36613);
nor U40143 (N_40143,N_30552,N_37417);
or U40144 (N_40144,N_38032,N_34375);
or U40145 (N_40145,N_36472,N_32612);
or U40146 (N_40146,N_37676,N_39218);
xnor U40147 (N_40147,N_34322,N_39854);
nand U40148 (N_40148,N_32737,N_35990);
or U40149 (N_40149,N_39221,N_33579);
and U40150 (N_40150,N_36244,N_30110);
nand U40151 (N_40151,N_32095,N_32578);
or U40152 (N_40152,N_32684,N_38020);
nor U40153 (N_40153,N_34137,N_31224);
nor U40154 (N_40154,N_33716,N_35007);
nor U40155 (N_40155,N_38717,N_30848);
nor U40156 (N_40156,N_31150,N_34238);
or U40157 (N_40157,N_36645,N_39384);
and U40158 (N_40158,N_30615,N_37821);
or U40159 (N_40159,N_30164,N_32247);
xor U40160 (N_40160,N_30751,N_39896);
nor U40161 (N_40161,N_37793,N_37576);
nor U40162 (N_40162,N_30920,N_30435);
and U40163 (N_40163,N_34924,N_38431);
and U40164 (N_40164,N_34640,N_39837);
or U40165 (N_40165,N_37182,N_35609);
nor U40166 (N_40166,N_33744,N_33701);
nand U40167 (N_40167,N_35859,N_30073);
or U40168 (N_40168,N_32820,N_32567);
xor U40169 (N_40169,N_33689,N_37243);
nand U40170 (N_40170,N_31659,N_30256);
xnor U40171 (N_40171,N_30318,N_34002);
or U40172 (N_40172,N_32909,N_32803);
and U40173 (N_40173,N_38264,N_38109);
or U40174 (N_40174,N_32654,N_35654);
nor U40175 (N_40175,N_30826,N_33899);
nand U40176 (N_40176,N_30336,N_36950);
and U40177 (N_40177,N_35350,N_35402);
xor U40178 (N_40178,N_33302,N_32791);
xor U40179 (N_40179,N_39600,N_33746);
nand U40180 (N_40180,N_30538,N_37782);
nor U40181 (N_40181,N_31068,N_36886);
nand U40182 (N_40182,N_33629,N_30398);
and U40183 (N_40183,N_32090,N_38986);
and U40184 (N_40184,N_33411,N_34437);
xor U40185 (N_40185,N_36245,N_30242);
xor U40186 (N_40186,N_32970,N_37160);
or U40187 (N_40187,N_31663,N_34304);
and U40188 (N_40188,N_32623,N_31187);
nor U40189 (N_40189,N_32550,N_35091);
and U40190 (N_40190,N_35807,N_30343);
nor U40191 (N_40191,N_31567,N_32352);
nor U40192 (N_40192,N_36227,N_32779);
nand U40193 (N_40193,N_33901,N_39892);
nor U40194 (N_40194,N_31759,N_38353);
nand U40195 (N_40195,N_36420,N_37306);
and U40196 (N_40196,N_33614,N_38982);
or U40197 (N_40197,N_34801,N_32818);
nor U40198 (N_40198,N_36770,N_35906);
and U40199 (N_40199,N_39130,N_34919);
nand U40200 (N_40200,N_30418,N_38057);
or U40201 (N_40201,N_39612,N_34403);
nand U40202 (N_40202,N_33949,N_33711);
or U40203 (N_40203,N_38146,N_34535);
and U40204 (N_40204,N_32703,N_30719);
or U40205 (N_40205,N_38299,N_37513);
or U40206 (N_40206,N_34878,N_39189);
xnor U40207 (N_40207,N_31716,N_31948);
or U40208 (N_40208,N_36671,N_33659);
or U40209 (N_40209,N_32042,N_33200);
nand U40210 (N_40210,N_33502,N_37805);
nand U40211 (N_40211,N_31559,N_39591);
nand U40212 (N_40212,N_39316,N_39437);
nand U40213 (N_40213,N_31351,N_38879);
nand U40214 (N_40214,N_39950,N_39155);
nand U40215 (N_40215,N_33534,N_30223);
nor U40216 (N_40216,N_31851,N_38136);
nand U40217 (N_40217,N_35748,N_34512);
or U40218 (N_40218,N_34550,N_32726);
nand U40219 (N_40219,N_33146,N_36794);
and U40220 (N_40220,N_37270,N_34637);
nand U40221 (N_40221,N_36468,N_31830);
nand U40222 (N_40222,N_31741,N_32705);
or U40223 (N_40223,N_36917,N_37740);
xnor U40224 (N_40224,N_37599,N_32158);
nand U40225 (N_40225,N_33414,N_39820);
nand U40226 (N_40226,N_31967,N_33887);
xnor U40227 (N_40227,N_39008,N_33886);
xnor U40228 (N_40228,N_37394,N_39570);
or U40229 (N_40229,N_34085,N_39451);
nand U40230 (N_40230,N_33601,N_35681);
nand U40231 (N_40231,N_33693,N_37110);
nor U40232 (N_40232,N_32311,N_31996);
nand U40233 (N_40233,N_32511,N_38149);
and U40234 (N_40234,N_35772,N_32525);
nor U40235 (N_40235,N_33860,N_37001);
xor U40236 (N_40236,N_37989,N_39195);
and U40237 (N_40237,N_37815,N_31903);
and U40238 (N_40238,N_33351,N_39035);
nor U40239 (N_40239,N_37746,N_33163);
nor U40240 (N_40240,N_31636,N_38002);
nor U40241 (N_40241,N_32023,N_35729);
nand U40242 (N_40242,N_32925,N_35644);
nor U40243 (N_40243,N_39842,N_35173);
nor U40244 (N_40244,N_34049,N_37469);
and U40245 (N_40245,N_35298,N_33583);
nor U40246 (N_40246,N_39069,N_32348);
xor U40247 (N_40247,N_37201,N_37012);
nand U40248 (N_40248,N_36231,N_31093);
xnor U40249 (N_40249,N_39546,N_33531);
or U40250 (N_40250,N_38627,N_32725);
nand U40251 (N_40251,N_33125,N_32866);
or U40252 (N_40252,N_34454,N_36772);
or U40253 (N_40253,N_33261,N_30049);
and U40254 (N_40254,N_31337,N_31376);
nor U40255 (N_40255,N_39589,N_36557);
or U40256 (N_40256,N_35365,N_36277);
xnor U40257 (N_40257,N_35914,N_37941);
nor U40258 (N_40258,N_33363,N_33246);
or U40259 (N_40259,N_34563,N_33309);
and U40260 (N_40260,N_31078,N_32824);
nor U40261 (N_40261,N_38139,N_34985);
or U40262 (N_40262,N_34928,N_34818);
or U40263 (N_40263,N_30740,N_34799);
xor U40264 (N_40264,N_36806,N_33813);
nand U40265 (N_40265,N_31002,N_39109);
or U40266 (N_40266,N_35233,N_33507);
nor U40267 (N_40267,N_34990,N_34824);
or U40268 (N_40268,N_32651,N_34915);
or U40269 (N_40269,N_30490,N_38176);
nand U40270 (N_40270,N_32995,N_33219);
nand U40271 (N_40271,N_32743,N_37499);
and U40272 (N_40272,N_32152,N_32298);
nand U40273 (N_40273,N_36525,N_35472);
or U40274 (N_40274,N_36792,N_30610);
xor U40275 (N_40275,N_35125,N_37249);
xnor U40276 (N_40276,N_34427,N_30240);
nor U40277 (N_40277,N_32362,N_33567);
nand U40278 (N_40278,N_34908,N_32113);
or U40279 (N_40279,N_36824,N_31826);
or U40280 (N_40280,N_32807,N_39951);
nor U40281 (N_40281,N_31297,N_32973);
nor U40282 (N_40282,N_39804,N_38786);
and U40283 (N_40283,N_35357,N_37351);
and U40284 (N_40284,N_30139,N_34172);
nand U40285 (N_40285,N_37794,N_38854);
or U40286 (N_40286,N_38781,N_39041);
and U40287 (N_40287,N_38634,N_34213);
xor U40288 (N_40288,N_32739,N_32517);
and U40289 (N_40289,N_36657,N_39039);
xor U40290 (N_40290,N_34672,N_33952);
or U40291 (N_40291,N_39320,N_35193);
and U40292 (N_40292,N_35884,N_37424);
xor U40293 (N_40293,N_33155,N_33478);
xor U40294 (N_40294,N_37826,N_34540);
nand U40295 (N_40295,N_35586,N_33438);
and U40296 (N_40296,N_35791,N_39826);
nor U40297 (N_40297,N_36432,N_35767);
or U40298 (N_40298,N_39885,N_37619);
or U40299 (N_40299,N_30374,N_34000);
or U40300 (N_40300,N_30488,N_33661);
nor U40301 (N_40301,N_34671,N_35219);
and U40302 (N_40302,N_34101,N_39328);
nor U40303 (N_40303,N_39860,N_39969);
nor U40304 (N_40304,N_35636,N_33066);
or U40305 (N_40305,N_33885,N_35614);
or U40306 (N_40306,N_32691,N_37730);
and U40307 (N_40307,N_31748,N_30939);
or U40308 (N_40308,N_39337,N_38273);
and U40309 (N_40309,N_30359,N_32016);
nor U40310 (N_40310,N_35668,N_37985);
xnor U40311 (N_40311,N_32827,N_37528);
nor U40312 (N_40312,N_35564,N_30152);
and U40313 (N_40313,N_36983,N_30113);
or U40314 (N_40314,N_31523,N_39535);
or U40315 (N_40315,N_32938,N_36480);
and U40316 (N_40316,N_35273,N_30052);
xnor U40317 (N_40317,N_37771,N_35555);
and U40318 (N_40318,N_38429,N_37621);
nand U40319 (N_40319,N_39596,N_37671);
and U40320 (N_40320,N_35226,N_35287);
nand U40321 (N_40321,N_30412,N_31853);
and U40322 (N_40322,N_32086,N_38797);
nand U40323 (N_40323,N_37708,N_35856);
nor U40324 (N_40324,N_37990,N_30799);
nor U40325 (N_40325,N_36170,N_36519);
nand U40326 (N_40326,N_39681,N_37388);
nor U40327 (N_40327,N_36836,N_36121);
and U40328 (N_40328,N_38315,N_30157);
nand U40329 (N_40329,N_35381,N_32950);
nand U40330 (N_40330,N_33740,N_39615);
xnor U40331 (N_40331,N_31966,N_39144);
xnor U40332 (N_40332,N_32307,N_38890);
and U40333 (N_40333,N_39653,N_34461);
xnor U40334 (N_40334,N_35670,N_32678);
nor U40335 (N_40335,N_34074,N_36808);
xnor U40336 (N_40336,N_34117,N_31407);
or U40337 (N_40337,N_36830,N_32130);
nand U40338 (N_40338,N_34313,N_37439);
xnor U40339 (N_40339,N_33552,N_32409);
and U40340 (N_40340,N_32747,N_34944);
xor U40341 (N_40341,N_38795,N_37519);
nand U40342 (N_40342,N_33004,N_34645);
nand U40343 (N_40343,N_39145,N_37476);
nor U40344 (N_40344,N_32723,N_37898);
or U40345 (N_40345,N_33437,N_39002);
xor U40346 (N_40346,N_30503,N_33143);
nor U40347 (N_40347,N_35290,N_32315);
and U40348 (N_40348,N_39419,N_37509);
nand U40349 (N_40349,N_35886,N_30898);
and U40350 (N_40350,N_36814,N_36075);
xor U40351 (N_40351,N_39724,N_31889);
xnor U40352 (N_40352,N_31225,N_35230);
or U40353 (N_40353,N_30984,N_31378);
or U40354 (N_40354,N_31831,N_35587);
xnor U40355 (N_40355,N_30403,N_39562);
or U40356 (N_40356,N_31323,N_32563);
or U40357 (N_40357,N_31051,N_34475);
or U40358 (N_40358,N_33165,N_36775);
nand U40359 (N_40359,N_33170,N_31681);
or U40360 (N_40360,N_30395,N_30676);
or U40361 (N_40361,N_35743,N_34426);
xor U40362 (N_40362,N_33816,N_32599);
nand U40363 (N_40363,N_31149,N_38098);
and U40364 (N_40364,N_32302,N_35499);
and U40365 (N_40365,N_36107,N_31960);
nand U40366 (N_40366,N_34064,N_34613);
nor U40367 (N_40367,N_31069,N_36255);
xor U40368 (N_40368,N_37059,N_38756);
nand U40369 (N_40369,N_30220,N_36745);
xor U40370 (N_40370,N_36291,N_34847);
nor U40371 (N_40371,N_35607,N_33154);
xnor U40372 (N_40372,N_38025,N_34107);
or U40373 (N_40373,N_36831,N_36407);
nor U40374 (N_40374,N_31884,N_34580);
xor U40375 (N_40375,N_30502,N_35559);
nor U40376 (N_40376,N_37026,N_31665);
xor U40377 (N_40377,N_30957,N_35596);
xnor U40378 (N_40378,N_34408,N_32122);
xnor U40379 (N_40379,N_31385,N_35918);
nor U40380 (N_40380,N_33439,N_32343);
nand U40381 (N_40381,N_30390,N_33172);
xor U40382 (N_40382,N_37204,N_32625);
nor U40383 (N_40383,N_37510,N_35005);
or U40384 (N_40384,N_31028,N_35372);
or U40385 (N_40385,N_30895,N_33410);
or U40386 (N_40386,N_36240,N_35455);
and U40387 (N_40387,N_31391,N_36651);
nor U40388 (N_40388,N_31575,N_34021);
or U40389 (N_40389,N_33365,N_38345);
nand U40390 (N_40390,N_33048,N_32460);
or U40391 (N_40391,N_32250,N_31139);
xor U40392 (N_40392,N_31894,N_39580);
nand U40393 (N_40393,N_32234,N_35049);
nand U40394 (N_40394,N_38015,N_38642);
and U40395 (N_40395,N_39735,N_33075);
or U40396 (N_40396,N_34873,N_32038);
and U40397 (N_40397,N_32055,N_39102);
xor U40398 (N_40398,N_34854,N_34065);
or U40399 (N_40399,N_31703,N_31500);
xnor U40400 (N_40400,N_38481,N_32890);
nor U40401 (N_40401,N_36605,N_31651);
xor U40402 (N_40402,N_30087,N_39730);
or U40403 (N_40403,N_37811,N_34651);
nand U40404 (N_40404,N_37765,N_35138);
xor U40405 (N_40405,N_31596,N_39167);
xor U40406 (N_40406,N_37134,N_37580);
and U40407 (N_40407,N_31288,N_30184);
nor U40408 (N_40408,N_33649,N_33533);
nor U40409 (N_40409,N_33749,N_38078);
and U40410 (N_40410,N_32554,N_30739);
nor U40411 (N_40411,N_36216,N_35849);
nand U40412 (N_40412,N_31480,N_32132);
nor U40413 (N_40413,N_37209,N_38590);
or U40414 (N_40414,N_37668,N_31684);
nor U40415 (N_40415,N_36331,N_32437);
xnor U40416 (N_40416,N_39699,N_38626);
or U40417 (N_40417,N_36991,N_37091);
and U40418 (N_40418,N_35953,N_31970);
nor U40419 (N_40419,N_35911,N_38200);
and U40420 (N_40420,N_39788,N_32410);
xnor U40421 (N_40421,N_38771,N_30168);
nor U40422 (N_40422,N_30536,N_35492);
xnor U40423 (N_40423,N_36145,N_33958);
nor U40424 (N_40424,N_38678,N_33079);
nor U40425 (N_40425,N_38870,N_36484);
and U40426 (N_40426,N_36801,N_37753);
or U40427 (N_40427,N_32127,N_37834);
nand U40428 (N_40428,N_36767,N_33287);
xor U40429 (N_40429,N_38591,N_36421);
nor U40430 (N_40430,N_38207,N_39894);
and U40431 (N_40431,N_38092,N_33779);
nand U40432 (N_40432,N_37508,N_38189);
nor U40433 (N_40433,N_35387,N_32497);
or U40434 (N_40434,N_35512,N_38514);
xnor U40435 (N_40435,N_39412,N_36592);
nand U40436 (N_40436,N_31148,N_34828);
and U40437 (N_40437,N_39924,N_32920);
xnor U40438 (N_40438,N_34954,N_39795);
and U40439 (N_40439,N_37322,N_36654);
nand U40440 (N_40440,N_39240,N_37867);
or U40441 (N_40441,N_39193,N_34495);
nor U40442 (N_40442,N_38341,N_38741);
nand U40443 (N_40443,N_30124,N_32642);
nand U40444 (N_40444,N_38903,N_32655);
nand U40445 (N_40445,N_36030,N_33795);
nand U40446 (N_40446,N_31459,N_35760);
and U40447 (N_40447,N_39658,N_39201);
and U40448 (N_40448,N_36928,N_32555);
or U40449 (N_40449,N_33926,N_33058);
or U40450 (N_40450,N_36713,N_31827);
or U40451 (N_40451,N_37473,N_32792);
and U40452 (N_40452,N_31731,N_36312);
or U40453 (N_40453,N_36788,N_38425);
or U40454 (N_40454,N_36805,N_37084);
and U40455 (N_40455,N_31079,N_38851);
xor U40456 (N_40456,N_33417,N_37039);
xnor U40457 (N_40457,N_37025,N_35984);
nand U40458 (N_40458,N_31605,N_38278);
and U40459 (N_40459,N_39272,N_39564);
nand U40460 (N_40460,N_36091,N_39468);
or U40461 (N_40461,N_30801,N_38269);
nor U40462 (N_40462,N_37009,N_30236);
nor U40463 (N_40463,N_39223,N_31279);
xor U40464 (N_40464,N_39769,N_37535);
xor U40465 (N_40465,N_34656,N_34451);
nor U40466 (N_40466,N_38133,N_38036);
and U40467 (N_40467,N_39284,N_33514);
and U40468 (N_40468,N_33254,N_30039);
or U40469 (N_40469,N_36232,N_34521);
and U40470 (N_40470,N_33944,N_33637);
xnor U40471 (N_40471,N_38849,N_37768);
xor U40472 (N_40472,N_33520,N_39282);
or U40473 (N_40473,N_33012,N_33033);
nand U40474 (N_40474,N_38377,N_34244);
or U40475 (N_40475,N_39243,N_35342);
xnor U40476 (N_40476,N_36222,N_36722);
or U40477 (N_40477,N_38871,N_35187);
xnor U40478 (N_40478,N_30238,N_35908);
or U40479 (N_40479,N_39222,N_35015);
xnor U40480 (N_40480,N_38165,N_33510);
or U40481 (N_40481,N_35053,N_32178);
nand U40482 (N_40482,N_33319,N_31604);
nand U40483 (N_40483,N_31617,N_38650);
nor U40484 (N_40484,N_38758,N_39181);
xnor U40485 (N_40485,N_33780,N_35176);
or U40486 (N_40486,N_34841,N_35105);
xnor U40487 (N_40487,N_37133,N_30896);
xor U40488 (N_40488,N_35592,N_39952);
nor U40489 (N_40489,N_30376,N_39433);
nor U40490 (N_40490,N_33845,N_38291);
and U40491 (N_40491,N_30279,N_31506);
and U40492 (N_40492,N_34532,N_37307);
nor U40493 (N_40493,N_39923,N_33289);
nand U40494 (N_40494,N_35653,N_33485);
or U40495 (N_40495,N_34949,N_33613);
and U40496 (N_40496,N_31533,N_35575);
and U40497 (N_40497,N_34407,N_37884);
or U40498 (N_40498,N_30341,N_39487);
nand U40499 (N_40499,N_36488,N_39526);
or U40500 (N_40500,N_34170,N_35597);
nor U40501 (N_40501,N_36644,N_33386);
nor U40502 (N_40502,N_32697,N_31095);
xnor U40503 (N_40503,N_38440,N_37261);
xor U40504 (N_40504,N_35329,N_35569);
nor U40505 (N_40505,N_32600,N_30672);
and U40506 (N_40506,N_31838,N_36153);
nand U40507 (N_40507,N_37830,N_38038);
or U40508 (N_40508,N_33072,N_39162);
xor U40509 (N_40509,N_39774,N_31504);
or U40510 (N_40510,N_31471,N_31843);
and U40511 (N_40511,N_30375,N_32819);
nand U40512 (N_40512,N_37774,N_37624);
and U40513 (N_40513,N_31188,N_30103);
nor U40514 (N_40514,N_30805,N_37933);
xnor U40515 (N_40515,N_34920,N_31906);
or U40516 (N_40516,N_34469,N_34906);
xnor U40517 (N_40517,N_30221,N_35640);
or U40518 (N_40518,N_39849,N_38958);
xor U40519 (N_40519,N_30397,N_34043);
nor U40520 (N_40520,N_37905,N_39374);
nand U40521 (N_40521,N_37144,N_33426);
and U40522 (N_40522,N_30339,N_35227);
xor U40523 (N_40523,N_33267,N_31885);
nand U40524 (N_40524,N_39147,N_31512);
nor U40525 (N_40525,N_37645,N_34470);
nor U40526 (N_40526,N_38907,N_37211);
or U40527 (N_40527,N_33080,N_36390);
or U40528 (N_40528,N_38305,N_38151);
xor U40529 (N_40529,N_33995,N_31673);
or U40530 (N_40530,N_31468,N_30294);
nand U40531 (N_40531,N_32264,N_32789);
nand U40532 (N_40532,N_38980,N_32239);
nand U40533 (N_40533,N_35314,N_34783);
nor U40534 (N_40534,N_37341,N_37496);
and U40535 (N_40535,N_30024,N_35921);
and U40536 (N_40536,N_35808,N_38733);
and U40537 (N_40537,N_38532,N_30530);
xor U40538 (N_40538,N_33399,N_32392);
nand U40539 (N_40539,N_34320,N_30881);
xnor U40540 (N_40540,N_36356,N_36946);
or U40541 (N_40541,N_30725,N_31040);
or U40542 (N_40542,N_35749,N_35599);
xnor U40543 (N_40543,N_30921,N_31536);
xor U40544 (N_40544,N_32117,N_37892);
and U40545 (N_40545,N_37744,N_32430);
or U40546 (N_40546,N_36308,N_30155);
nand U40547 (N_40547,N_39018,N_30394);
nor U40548 (N_40548,N_36148,N_39170);
nor U40549 (N_40549,N_33049,N_39308);
nor U40550 (N_40550,N_35446,N_39420);
and U40551 (N_40551,N_33406,N_39687);
nand U40552 (N_40552,N_37789,N_37086);
and U40553 (N_40553,N_33269,N_36575);
xor U40554 (N_40554,N_33781,N_34662);
or U40555 (N_40555,N_36281,N_32499);
nor U40556 (N_40556,N_36223,N_31278);
or U40557 (N_40557,N_39073,N_33419);
nand U40558 (N_40558,N_33674,N_33599);
xor U40559 (N_40559,N_33936,N_37996);
nor U40560 (N_40560,N_31243,N_33965);
nand U40561 (N_40561,N_39264,N_37156);
and U40562 (N_40562,N_38224,N_32468);
nor U40563 (N_40563,N_31497,N_32219);
nand U40564 (N_40564,N_33101,N_34256);
and U40565 (N_40565,N_35771,N_36463);
and U40566 (N_40566,N_35521,N_33334);
xor U40567 (N_40567,N_30176,N_33109);
nand U40568 (N_40568,N_39755,N_39205);
and U40569 (N_40569,N_31790,N_34216);
and U40570 (N_40570,N_31408,N_32476);
nand U40571 (N_40571,N_32645,N_38062);
and U40572 (N_40572,N_33941,N_31642);
xnor U40573 (N_40573,N_36550,N_39467);
or U40574 (N_40574,N_38814,N_38122);
and U40575 (N_40575,N_38855,N_32787);
xor U40576 (N_40576,N_38583,N_39219);
xnor U40577 (N_40577,N_36921,N_33168);
nor U40578 (N_40578,N_39173,N_39873);
nand U40579 (N_40579,N_31927,N_35546);
xor U40580 (N_40580,N_32369,N_32858);
nor U40581 (N_40581,N_32911,N_38318);
xnor U40582 (N_40582,N_30263,N_35106);
or U40583 (N_40583,N_39707,N_31557);
nand U40584 (N_40584,N_35028,N_30884);
nand U40585 (N_40585,N_35376,N_37637);
or U40586 (N_40586,N_32346,N_38656);
or U40587 (N_40587,N_32326,N_34060);
nor U40588 (N_40588,N_37092,N_34118);
or U40589 (N_40589,N_34700,N_39542);
nor U40590 (N_40590,N_34945,N_36627);
or U40591 (N_40591,N_35228,N_31313);
nand U40592 (N_40592,N_38248,N_38304);
and U40593 (N_40593,N_33570,N_33796);
or U40594 (N_40594,N_31130,N_34660);
nor U40595 (N_40595,N_32713,N_37956);
and U40596 (N_40596,N_30027,N_35537);
nand U40597 (N_40597,N_38941,N_32861);
xor U40598 (N_40598,N_34017,N_33354);
xor U40599 (N_40599,N_30405,N_36839);
and U40600 (N_40600,N_31119,N_36565);
nor U40601 (N_40601,N_30922,N_36620);
nor U40602 (N_40602,N_39094,N_36935);
nor U40603 (N_40603,N_32776,N_31720);
nor U40604 (N_40604,N_33090,N_33105);
or U40605 (N_40605,N_35059,N_36924);
nand U40606 (N_40606,N_30188,N_31620);
xnor U40607 (N_40607,N_39161,N_33785);
xnor U40608 (N_40608,N_36461,N_32533);
nor U40609 (N_40609,N_37893,N_36907);
or U40610 (N_40610,N_37615,N_36536);
nand U40611 (N_40611,N_32741,N_31165);
and U40612 (N_40612,N_35251,N_31511);
nor U40613 (N_40613,N_36074,N_31754);
xnor U40614 (N_40614,N_30949,N_33738);
xnor U40615 (N_40615,N_37924,N_36556);
and U40616 (N_40616,N_37596,N_31722);
and U40617 (N_40617,N_39369,N_33758);
and U40618 (N_40618,N_32138,N_36672);
or U40619 (N_40619,N_32847,N_38229);
nor U40620 (N_40620,N_30253,N_35779);
or U40621 (N_40621,N_31209,N_30335);
or U40622 (N_40622,N_33238,N_31195);
and U40623 (N_40623,N_35813,N_30248);
xnor U40624 (N_40624,N_34378,N_39289);
nor U40625 (N_40625,N_37463,N_30862);
nor U40626 (N_40626,N_30153,N_31346);
nand U40627 (N_40627,N_33123,N_30009);
or U40628 (N_40628,N_38325,N_35524);
and U40629 (N_40629,N_32797,N_34453);
xnor U40630 (N_40630,N_38880,N_34361);
xnor U40631 (N_40631,N_34381,N_39273);
and U40632 (N_40632,N_30150,N_31951);
nand U40633 (N_40633,N_37297,N_38588);
or U40634 (N_40634,N_39565,N_37876);
or U40635 (N_40635,N_36430,N_35827);
nand U40636 (N_40636,N_36553,N_39827);
nand U40637 (N_40637,N_32203,N_36132);
and U40638 (N_40638,N_33129,N_32375);
nand U40639 (N_40639,N_35988,N_34056);
or U40640 (N_40640,N_34509,N_31850);
nor U40641 (N_40641,N_33245,N_33896);
nor U40642 (N_40642,N_38534,N_35412);
nand U40643 (N_40643,N_33288,N_31707);
nand U40644 (N_40644,N_31153,N_36702);
or U40645 (N_40645,N_32899,N_35245);
xor U40646 (N_40646,N_36717,N_38053);
nand U40647 (N_40647,N_39907,N_30640);
nand U40648 (N_40648,N_34545,N_39016);
nor U40649 (N_40649,N_31984,N_32029);
or U40650 (N_40650,N_32991,N_37116);
nor U40651 (N_40651,N_34849,N_39787);
nor U40652 (N_40652,N_38087,N_37854);
or U40653 (N_40653,N_35244,N_31240);
and U40654 (N_40654,N_38270,N_34129);
and U40655 (N_40655,N_35780,N_34264);
xnor U40656 (N_40656,N_35811,N_37344);
or U40657 (N_40657,N_39480,N_34193);
or U40658 (N_40658,N_32160,N_37927);
nand U40659 (N_40659,N_36058,N_34881);
nand U40660 (N_40660,N_32323,N_36402);
nor U40661 (N_40661,N_34811,N_33489);
nor U40662 (N_40662,N_38177,N_33897);
or U40663 (N_40663,N_31321,N_31999);
and U40664 (N_40664,N_37043,N_34165);
or U40665 (N_40665,N_35383,N_35840);
nor U40666 (N_40666,N_35190,N_36481);
xnor U40667 (N_40667,N_37850,N_38672);
nor U40668 (N_40668,N_36048,N_39417);
xnor U40669 (N_40669,N_34409,N_34104);
xor U40670 (N_40670,N_36985,N_35481);
nor U40671 (N_40671,N_32853,N_35983);
nand U40672 (N_40672,N_31007,N_36043);
xnor U40673 (N_40673,N_35425,N_34609);
nand U40674 (N_40674,N_33496,N_38836);
nand U40675 (N_40675,N_36299,N_33980);
nor U40676 (N_40676,N_32394,N_31529);
and U40677 (N_40677,N_38774,N_38222);
nand U40678 (N_40678,N_32458,N_34391);
nor U40679 (N_40679,N_32305,N_37085);
nand U40680 (N_40680,N_30601,N_38753);
xnor U40681 (N_40681,N_30772,N_39389);
or U40682 (N_40682,N_33617,N_36719);
or U40683 (N_40683,N_30682,N_34389);
nand U40684 (N_40684,N_30338,N_39622);
or U40685 (N_40685,N_33057,N_31053);
nor U40686 (N_40686,N_35256,N_39823);
or U40687 (N_40687,N_32030,N_37004);
xor U40688 (N_40688,N_30097,N_39568);
nor U40689 (N_40689,N_38662,N_36741);
nand U40690 (N_40690,N_36547,N_38633);
nor U40691 (N_40691,N_31433,N_34589);
nor U40692 (N_40692,N_38399,N_38178);
or U40693 (N_40693,N_36067,N_36520);
xor U40694 (N_40694,N_30416,N_32683);
or U40695 (N_40695,N_34569,N_36124);
and U40696 (N_40696,N_30966,N_35038);
xnor U40697 (N_40697,N_32908,N_38234);
or U40698 (N_40698,N_35651,N_36674);
or U40699 (N_40699,N_38058,N_38895);
xor U40700 (N_40700,N_34484,N_30947);
and U40701 (N_40701,N_35514,N_30802);
nor U40702 (N_40702,N_31615,N_30636);
nand U40703 (N_40703,N_33568,N_30227);
and U40704 (N_40704,N_39814,N_36785);
nand U40705 (N_40705,N_39004,N_38625);
and U40706 (N_40706,N_33925,N_39700);
or U40707 (N_40707,N_32740,N_36630);
nor U40708 (N_40708,N_35800,N_30612);
xnor U40709 (N_40709,N_35191,N_37062);
and U40710 (N_40710,N_31016,N_31055);
nand U40711 (N_40711,N_32639,N_33643);
nand U40712 (N_40712,N_38158,N_39696);
xor U40713 (N_40713,N_39561,N_39662);
xnor U40714 (N_40714,N_34946,N_36817);
nand U40715 (N_40715,N_39819,N_31509);
xnor U40716 (N_40716,N_36524,N_34740);
nor U40717 (N_40717,N_31226,N_39598);
nand U40718 (N_40718,N_37558,N_37370);
nor U40719 (N_40719,N_37803,N_38080);
nand U40720 (N_40720,N_31001,N_32258);
nor U40721 (N_40721,N_31949,N_38458);
or U40722 (N_40722,N_34603,N_39404);
and U40723 (N_40723,N_36708,N_33041);
or U40724 (N_40724,N_34460,N_32648);
nor U40725 (N_40725,N_34054,N_37406);
xor U40726 (N_40726,N_36682,N_30836);
and U40727 (N_40727,N_34223,N_39721);
nor U40728 (N_40728,N_39948,N_33681);
xnor U40729 (N_40729,N_36916,N_33854);
nor U40730 (N_40730,N_32559,N_32157);
nor U40731 (N_40731,N_35540,N_30960);
or U40732 (N_40732,N_33920,N_32495);
and U40733 (N_40733,N_39897,N_30060);
and U40734 (N_40734,N_32749,N_32020);
xor U40735 (N_40735,N_30032,N_30001);
and U40736 (N_40736,N_31000,N_39778);
nor U40737 (N_40737,N_32411,N_32761);
and U40738 (N_40738,N_36016,N_38253);
or U40739 (N_40739,N_31070,N_36000);
nand U40740 (N_40740,N_31953,N_35691);
nor U40741 (N_40741,N_35266,N_35449);
and U40742 (N_40742,N_33937,N_36364);
nand U40743 (N_40743,N_35413,N_36085);
nor U40744 (N_40744,N_33382,N_32209);
nand U40745 (N_40745,N_37115,N_38367);
and U40746 (N_40746,N_30245,N_35826);
nand U40747 (N_40747,N_31758,N_36517);
or U40748 (N_40748,N_39460,N_37919);
xnor U40749 (N_40749,N_37371,N_36726);
xor U40750 (N_40750,N_31763,N_34438);
nor U40751 (N_40751,N_39928,N_39300);
nand U40752 (N_40752,N_38385,N_35682);
nor U40753 (N_40753,N_34781,N_30275);
xor U40754 (N_40754,N_33264,N_32384);
nor U40755 (N_40755,N_33451,N_39507);
nor U40756 (N_40756,N_36400,N_39825);
nand U40757 (N_40757,N_30761,N_36022);
nor U40758 (N_40758,N_34724,N_35831);
nand U40759 (N_40759,N_37484,N_31897);
xor U40760 (N_40760,N_37416,N_31576);
or U40761 (N_40761,N_36493,N_32194);
nor U40762 (N_40762,N_32006,N_39532);
xor U40763 (N_40763,N_31330,N_36021);
and U40764 (N_40764,N_32700,N_32971);
nor U40765 (N_40765,N_36168,N_36780);
nand U40766 (N_40766,N_34479,N_32288);
nand U40767 (N_40767,N_38388,N_39110);
xnor U40768 (N_40768,N_36088,N_32123);
nand U40769 (N_40769,N_39719,N_38560);
and U40770 (N_40770,N_31739,N_33429);
nor U40771 (N_40771,N_35496,N_30854);
xnor U40772 (N_40772,N_37714,N_30147);
or U40773 (N_40773,N_33089,N_38671);
xnor U40774 (N_40774,N_30996,N_39085);
xnor U40775 (N_40775,N_31386,N_31103);
or U40776 (N_40776,N_38292,N_37240);
nor U40777 (N_40777,N_36816,N_30423);
nand U40778 (N_40778,N_34728,N_38004);
or U40779 (N_40779,N_34341,N_35930);
nor U40780 (N_40780,N_31802,N_33635);
or U40781 (N_40781,N_35917,N_38479);
and U40782 (N_40782,N_33831,N_38166);
nor U40783 (N_40783,N_39172,N_32534);
xnor U40784 (N_40784,N_35171,N_30633);
xnor U40785 (N_40785,N_38936,N_38536);
nand U40786 (N_40786,N_38040,N_34447);
xor U40787 (N_40787,N_36603,N_35487);
xnor U40788 (N_40788,N_34751,N_31272);
xor U40789 (N_40789,N_33826,N_33082);
nor U40790 (N_40790,N_30877,N_36530);
nand U40791 (N_40791,N_38384,N_31056);
nand U40792 (N_40792,N_32014,N_35845);
or U40793 (N_40793,N_33685,N_35910);
nand U40794 (N_40794,N_32812,N_30965);
or U40795 (N_40795,N_36362,N_37272);
nand U40796 (N_40796,N_35829,N_32084);
xnor U40797 (N_40797,N_39863,N_35355);
and U40798 (N_40798,N_34232,N_39587);
nand U40799 (N_40799,N_33486,N_34596);
nor U40800 (N_40800,N_35104,N_38646);
or U40801 (N_40801,N_32832,N_35137);
nand U40802 (N_40802,N_38552,N_36369);
and U40803 (N_40803,N_32721,N_39059);
xor U40804 (N_40804,N_39278,N_38791);
nand U40805 (N_40805,N_36346,N_34301);
nand U40806 (N_40806,N_30356,N_37728);
and U40807 (N_40807,N_33543,N_38203);
nand U40808 (N_40808,N_38360,N_39695);
or U40809 (N_40809,N_30575,N_35048);
nand U40810 (N_40810,N_37414,N_38528);
nor U40811 (N_40811,N_37970,N_38621);
xor U40812 (N_40812,N_39684,N_35684);
nand U40813 (N_40813,N_31972,N_39644);
or U40814 (N_40814,N_36662,N_38891);
and U40815 (N_40815,N_35877,N_39453);
or U40816 (N_40816,N_39926,N_38000);
nand U40817 (N_40817,N_34154,N_36643);
and U40818 (N_40818,N_32826,N_36646);
or U40819 (N_40819,N_32526,N_38043);
xor U40820 (N_40820,N_34182,N_34843);
xor U40821 (N_40821,N_39182,N_38406);
and U40822 (N_40822,N_36204,N_31017);
nor U40823 (N_40823,N_31092,N_39309);
and U40824 (N_40824,N_32752,N_37368);
nor U40825 (N_40825,N_37662,N_31974);
xnor U40826 (N_40826,N_33490,N_33561);
nand U40827 (N_40827,N_33766,N_34744);
or U40828 (N_40828,N_33812,N_33206);
xor U40829 (N_40829,N_38359,N_30283);
and U40830 (N_40830,N_33658,N_32653);
nor U40831 (N_40831,N_39821,N_36185);
or U40832 (N_40832,N_31762,N_36659);
and U40833 (N_40833,N_30476,N_34791);
or U40834 (N_40834,N_39551,N_39253);
nor U40835 (N_40835,N_37572,N_39665);
nor U40836 (N_40836,N_38438,N_37138);
and U40837 (N_40837,N_35454,N_38857);
nor U40838 (N_40838,N_39310,N_30345);
xor U40839 (N_40839,N_38471,N_37837);
xnor U40840 (N_40840,N_30134,N_37772);
and U40841 (N_40841,N_30537,N_32610);
xor U40842 (N_40842,N_32252,N_36199);
xnor U40843 (N_40843,N_35021,N_36840);
xnor U40844 (N_40844,N_31551,N_30489);
nand U40845 (N_40845,N_31931,N_32518);
nor U40846 (N_40846,N_35377,N_35474);
and U40847 (N_40847,N_34584,N_34636);
and U40848 (N_40848,N_39876,N_31141);
and U40849 (N_40849,N_34111,N_37786);
nand U40850 (N_40850,N_37316,N_36126);
or U40851 (N_40851,N_32289,N_34392);
xnor U40852 (N_40852,N_36259,N_39732);
nor U40853 (N_40853,N_38470,N_33364);
nand U40854 (N_40854,N_34122,N_30379);
nor U40855 (N_40855,N_31898,N_36205);
nand U40856 (N_40856,N_33321,N_32467);
xor U40857 (N_40857,N_36845,N_38358);
or U40858 (N_40858,N_37157,N_36264);
xnor U40859 (N_40859,N_37105,N_39697);
xor U40860 (N_40860,N_32953,N_37063);
nor U40861 (N_40861,N_34935,N_37797);
nor U40862 (N_40862,N_32823,N_33005);
and U40863 (N_40863,N_38210,N_38943);
or U40864 (N_40864,N_39124,N_32414);
and U40865 (N_40865,N_35246,N_38076);
xor U40866 (N_40866,N_34995,N_31367);
or U40867 (N_40867,N_34202,N_34635);
nand U40868 (N_40868,N_39342,N_33468);
xnor U40869 (N_40869,N_39552,N_36640);
or U40870 (N_40870,N_37813,N_30621);
nor U40871 (N_40871,N_33822,N_34502);
xnor U40872 (N_40872,N_35638,N_32900);
or U40873 (N_40873,N_35774,N_35828);
nand U40874 (N_40874,N_38894,N_35323);
and U40875 (N_40875,N_38640,N_32333);
nand U40876 (N_40876,N_35356,N_32266);
and U40877 (N_40877,N_30317,N_36270);
nor U40878 (N_40878,N_37889,N_38437);
and U40879 (N_40879,N_31127,N_39933);
xnor U40880 (N_40880,N_30963,N_36800);
or U40881 (N_40881,N_31464,N_35590);
nand U40882 (N_40882,N_37804,N_39159);
xnor U40883 (N_40883,N_39541,N_35237);
or U40884 (N_40884,N_32043,N_39459);
nor U40885 (N_40885,N_32865,N_32261);
nor U40886 (N_40886,N_31034,N_38736);
or U40887 (N_40887,N_36580,N_39694);
xnor U40888 (N_40888,N_37704,N_30191);
nor U40889 (N_40889,N_37785,N_39639);
nor U40890 (N_40890,N_35578,N_38867);
xnor U40891 (N_40891,N_34628,N_37809);
or U40892 (N_40892,N_35166,N_30589);
nand U40893 (N_40893,N_32406,N_37612);
nand U40894 (N_40894,N_32917,N_37814);
or U40895 (N_40895,N_33310,N_34071);
xnor U40896 (N_40896,N_38517,N_37659);
and U40897 (N_40897,N_30905,N_33344);
nor U40898 (N_40898,N_35542,N_39773);
and U40899 (N_40899,N_35709,N_34308);
and U40900 (N_40900,N_34709,N_35285);
and U40901 (N_40901,N_36842,N_36165);
nor U40902 (N_40902,N_33193,N_31769);
nand U40903 (N_40903,N_32193,N_36625);
nand U40904 (N_40904,N_36428,N_35275);
nor U40905 (N_40905,N_34631,N_36956);
nand U40906 (N_40906,N_35121,N_30129);
nor U40907 (N_40907,N_35820,N_36954);
and U40908 (N_40908,N_37507,N_39626);
nand U40909 (N_40909,N_32334,N_30500);
or U40910 (N_40910,N_33412,N_32510);
xnor U40911 (N_40911,N_38968,N_34877);
and U40912 (N_40912,N_37550,N_33210);
nand U40913 (N_40913,N_30766,N_35404);
nand U40914 (N_40914,N_33176,N_32945);
or U40915 (N_40915,N_38948,N_36466);
or U40916 (N_40916,N_38267,N_33300);
xor U40917 (N_40917,N_30808,N_32036);
xnor U40918 (N_40918,N_30940,N_30664);
nor U40919 (N_40919,N_33435,N_36329);
and U40920 (N_40920,N_32279,N_31483);
nand U40921 (N_40921,N_34250,N_32514);
nand U40922 (N_40922,N_33625,N_38018);
or U40923 (N_40923,N_39651,N_33522);
or U40924 (N_40924,N_38067,N_38687);
nor U40925 (N_40925,N_34638,N_31699);
and U40926 (N_40926,N_38813,N_34703);
or U40927 (N_40927,N_33787,N_36397);
xnor U40928 (N_40928,N_37433,N_35184);
xor U40929 (N_40929,N_36812,N_34627);
nor U40930 (N_40930,N_38979,N_39444);
xor U40931 (N_40931,N_32922,N_33265);
xnor U40932 (N_40932,N_36198,N_33190);
nand U40933 (N_40933,N_33482,N_34942);
nand U40934 (N_40934,N_37321,N_36663);
and U40935 (N_40935,N_33818,N_33244);
xnor U40936 (N_40936,N_39346,N_32568);
or U40937 (N_40937,N_31492,N_30415);
nand U40938 (N_40938,N_32431,N_37432);
xor U40939 (N_40939,N_35081,N_30487);
nor U40940 (N_40940,N_30189,N_32666);
nand U40941 (N_40941,N_39869,N_34921);
nand U40942 (N_40942,N_39656,N_39401);
and U40943 (N_40943,N_36026,N_33723);
nand U40944 (N_40944,N_34969,N_32928);
or U40945 (N_40945,N_38853,N_39466);
nor U40946 (N_40946,N_39640,N_31008);
xnor U40947 (N_40947,N_30630,N_34979);
nand U40948 (N_40948,N_38754,N_37918);
and U40949 (N_40949,N_35200,N_36049);
and U40950 (N_40950,N_36864,N_37005);
nor U40951 (N_40951,N_38309,N_38990);
nor U40952 (N_40952,N_38459,N_33792);
or U40953 (N_40953,N_39753,N_39932);
xor U40954 (N_40954,N_34368,N_31339);
nor U40955 (N_40955,N_32303,N_35650);
and U40956 (N_40956,N_33042,N_36908);
and U40957 (N_40957,N_33110,N_32491);
or U40958 (N_40958,N_30018,N_37597);
xor U40959 (N_40959,N_36833,N_35207);
nor U40960 (N_40960,N_30424,N_34883);
xor U40961 (N_40961,N_34554,N_33688);
xnor U40962 (N_40962,N_31662,N_31574);
nor U40963 (N_40963,N_30606,N_36567);
or U40964 (N_40964,N_32051,N_34983);
and U40965 (N_40965,N_39027,N_37219);
and U40966 (N_40966,N_34667,N_36306);
xor U40967 (N_40967,N_32453,N_33322);
or U40968 (N_40968,N_34704,N_33710);
or U40969 (N_40969,N_37863,N_30505);
nor U40970 (N_40970,N_31076,N_38190);
or U40971 (N_40971,N_31106,N_37871);
and U40972 (N_40972,N_34087,N_39269);
or U40973 (N_40973,N_30022,N_39479);
and U40974 (N_40974,N_35439,N_37340);
xor U40975 (N_40975,N_38023,N_35955);
and U40976 (N_40976,N_31756,N_34510);
nand U40977 (N_40977,N_34747,N_31143);
xor U40978 (N_40978,N_34556,N_37118);
nor U40979 (N_40979,N_33849,N_38126);
xor U40980 (N_40980,N_36479,N_37969);
and U40981 (N_40981,N_36500,N_31012);
xor U40982 (N_40982,N_38048,N_33878);
xor U40983 (N_40983,N_35294,N_34792);
nor U40984 (N_40984,N_39241,N_38245);
nand U40985 (N_40985,N_39225,N_31686);
or U40986 (N_40986,N_39543,N_36217);
or U40987 (N_40987,N_31177,N_30219);
and U40988 (N_40988,N_38021,N_34601);
and U40989 (N_40989,N_33922,N_30249);
and U40990 (N_40990,N_39301,N_31945);
and U40991 (N_40991,N_39913,N_34615);
or U40992 (N_40992,N_36704,N_30402);
and U40993 (N_40993,N_39508,N_37506);
and U40994 (N_40994,N_33518,N_35630);
xnor U40995 (N_40995,N_35677,N_33387);
nand U40996 (N_40996,N_37928,N_30008);
and U40997 (N_40997,N_39375,N_33951);
nor U40998 (N_40998,N_38501,N_37787);
and U40999 (N_40999,N_39544,N_37549);
or U41000 (N_41000,N_32521,N_31979);
nor U41001 (N_41001,N_32934,N_30233);
nand U41002 (N_41002,N_37167,N_35210);
nand U41003 (N_41003,N_35531,N_31817);
nor U41004 (N_41004,N_34359,N_34248);
and U41005 (N_41005,N_33409,N_39136);
and U41006 (N_41006,N_30437,N_38793);
and U41007 (N_41007,N_35934,N_39636);
or U41008 (N_41008,N_32852,N_33504);
nand U41009 (N_41009,N_35563,N_33815);
or U41010 (N_41010,N_33516,N_35385);
nand U41011 (N_41011,N_31260,N_34204);
nand U41012 (N_41012,N_34681,N_33620);
or U41013 (N_41013,N_32583,N_36822);
or U41014 (N_41014,N_36601,N_35538);
and U41015 (N_41015,N_35034,N_30809);
nand U41016 (N_41016,N_36927,N_39079);
nor U41017 (N_41017,N_37947,N_31656);
and U41018 (N_41018,N_39012,N_36730);
or U41019 (N_41019,N_31267,N_34997);
xnor U41020 (N_41020,N_32507,N_35763);
and U41021 (N_41021,N_36122,N_38187);
nand U41022 (N_41022,N_39554,N_36716);
or U41023 (N_41023,N_38731,N_33943);
and U41024 (N_41024,N_33515,N_30948);
nor U41025 (N_41025,N_35738,N_36005);
xnor U41026 (N_41026,N_32736,N_32786);
and U41027 (N_41027,N_33456,N_30827);
and U41028 (N_41028,N_30463,N_37462);
nand U41029 (N_41029,N_30426,N_35272);
and U41030 (N_41030,N_32636,N_34669);
xor U41031 (N_41031,N_37075,N_38599);
or U41032 (N_41032,N_37901,N_35397);
nand U41033 (N_41033,N_37532,N_38428);
and U41034 (N_41034,N_34518,N_35453);
nand U41035 (N_41035,N_35291,N_31168);
nand U41036 (N_41036,N_31682,N_34882);
nor U41037 (N_41037,N_34723,N_30132);
or U41038 (N_41038,N_30924,N_39691);
and U41039 (N_41039,N_31033,N_32153);
and U41040 (N_41040,N_30387,N_34838);
xor U41041 (N_41041,N_30154,N_32366);
or U41042 (N_41042,N_35664,N_37438);
nor U41043 (N_41043,N_39115,N_36429);
xor U41044 (N_41044,N_31704,N_32998);
or U41045 (N_41045,N_34413,N_35987);
or U41046 (N_41046,N_31124,N_38077);
nand U41047 (N_41047,N_37625,N_38840);
and U41048 (N_41048,N_39045,N_38316);
nand U41049 (N_41049,N_38411,N_38605);
nand U41050 (N_41050,N_31377,N_30756);
nor U41051 (N_41051,N_35089,N_33113);
xnor U41052 (N_41052,N_38320,N_36720);
and U41053 (N_41053,N_33349,N_34034);
nand U41054 (N_41054,N_39305,N_38832);
and U41055 (N_41055,N_37033,N_38086);
or U41056 (N_41056,N_35315,N_33656);
or U41057 (N_41057,N_35017,N_39593);
nand U41058 (N_41058,N_38218,N_31282);
and U41059 (N_41059,N_37556,N_37628);
xnor U41060 (N_41060,N_30093,N_34337);
xnor U41061 (N_41061,N_36265,N_34848);
xnor U41062 (N_41062,N_32904,N_38931);
nand U41063 (N_41063,N_33594,N_30118);
nor U41064 (N_41064,N_31228,N_30715);
or U41065 (N_41065,N_30455,N_31191);
nor U41066 (N_41066,N_30649,N_31369);
nor U41067 (N_41067,N_39750,N_37074);
nand U41068 (N_41068,N_39126,N_32146);
nor U41069 (N_41069,N_32441,N_39338);
and U41070 (N_41070,N_33619,N_33403);
nor U41071 (N_41071,N_39637,N_30373);
nor U41072 (N_41072,N_31475,N_38403);
and U41073 (N_41073,N_32898,N_31232);
or U41074 (N_41074,N_31541,N_33784);
xor U41075 (N_41075,N_35662,N_37028);
or U41076 (N_41076,N_37592,N_30608);
and U41077 (N_41077,N_37309,N_37915);
or U41078 (N_41078,N_31324,N_36906);
nand U41079 (N_41079,N_34428,N_33361);
or U41080 (N_41080,N_31108,N_38790);
nand U41081 (N_41081,N_32433,N_31553);
or U41082 (N_41082,N_39216,N_31976);
xnor U41083 (N_41083,N_37191,N_32698);
nor U41084 (N_41084,N_33962,N_33778);
nand U41085 (N_41085,N_34493,N_33742);
or U41086 (N_41086,N_33655,N_33590);
or U41087 (N_41087,N_31277,N_33205);
nand U41088 (N_41088,N_36118,N_39646);
xnor U41089 (N_41089,N_36441,N_35465);
nor U41090 (N_41090,N_38763,N_37594);
or U41091 (N_41091,N_32216,N_39105);
and U41092 (N_41092,N_34784,N_39495);
or U41093 (N_41093,N_32982,N_30131);
nor U41094 (N_41094,N_30474,N_35139);
xnor U41095 (N_41095,N_33540,N_37094);
xnor U41096 (N_41096,N_35013,N_36009);
and U41097 (N_41097,N_37584,N_39157);
and U41098 (N_41098,N_31061,N_34996);
nor U41099 (N_41099,N_30684,N_37899);
nand U41100 (N_41100,N_35047,N_39270);
or U41101 (N_41101,N_33902,N_35676);
xnor U41102 (N_41102,N_35724,N_36936);
xnor U41103 (N_41103,N_39802,N_33028);
and U41104 (N_41104,N_31326,N_30316);
and U41105 (N_41105,N_32457,N_34145);
nand U41106 (N_41106,N_35753,N_36250);
and U41107 (N_41107,N_31049,N_36978);
nor U41108 (N_41108,N_30547,N_31757);
xnor U41109 (N_41109,N_32862,N_31908);
or U41110 (N_41110,N_34483,N_37702);
and U41111 (N_41111,N_30041,N_36194);
nor U41112 (N_41112,N_32699,N_33638);
xor U41113 (N_41113,N_33672,N_38268);
or U41114 (N_41114,N_37660,N_37586);
nor U41115 (N_41115,N_33017,N_37920);
nor U41116 (N_41116,N_36297,N_30094);
and U41117 (N_41117,N_35944,N_35986);
and U41118 (N_41118,N_33772,N_33400);
xnor U41119 (N_41119,N_33348,N_39123);
nor U41120 (N_41120,N_36294,N_37245);
xnor U41121 (N_41121,N_32144,N_38408);
and U41122 (N_41122,N_38681,N_36321);
nand U41123 (N_41123,N_32751,N_39371);
xnor U41124 (N_41124,N_34696,N_32054);
or U41125 (N_41125,N_39777,N_37687);
nand U41126 (N_41126,N_31611,N_39245);
xnor U41127 (N_41127,N_30211,N_36609);
nor U41128 (N_41128,N_38725,N_38156);
and U41129 (N_41129,N_35352,N_37524);
xnor U41130 (N_41130,N_35307,N_34070);
and U41131 (N_41131,N_39044,N_36852);
or U41132 (N_41132,N_37139,N_36544);
nor U41133 (N_41133,N_38064,N_32189);
or U41134 (N_41134,N_36827,N_36509);
nand U41135 (N_41135,N_32131,N_37657);
and U41136 (N_41136,N_39512,N_34754);
xnor U41137 (N_41137,N_35418,N_33059);
nand U41138 (N_41138,N_34120,N_35362);
nor U41139 (N_41139,N_39432,N_30815);
and U41140 (N_41140,N_32828,N_31309);
and U41141 (N_41141,N_30869,N_33034);
nor U41142 (N_41142,N_33580,N_33204);
and U41143 (N_41143,N_31577,N_31544);
and U41144 (N_41144,N_38142,N_34543);
or U41145 (N_41145,N_33765,N_34310);
and U41146 (N_41146,N_33471,N_38868);
xor U41147 (N_41147,N_33802,N_36380);
and U41148 (N_41148,N_37697,N_35466);
or U41149 (N_41149,N_38307,N_37102);
or U41150 (N_41150,N_33654,N_38987);
or U41151 (N_41151,N_32383,N_32793);
and U41152 (N_41152,N_35675,N_39829);
and U41153 (N_41153,N_36538,N_30368);
xor U41154 (N_41154,N_36969,N_37574);
xnor U41155 (N_41155,N_33633,N_32482);
nand U41156 (N_41156,N_36037,N_32200);
xor U41157 (N_41157,N_39973,N_36623);
or U41158 (N_41158,N_32377,N_35879);
and U41159 (N_41159,N_30839,N_38419);
xor U41160 (N_41160,N_33128,N_36633);
and U41161 (N_41161,N_39737,N_39421);
or U41162 (N_41162,N_37169,N_39603);
nor U41163 (N_41163,N_32318,N_32674);
xnor U41164 (N_41164,N_34722,N_34914);
and U41165 (N_41165,N_31419,N_37124);
nand U41166 (N_41166,N_34424,N_35183);
nand U41167 (N_41167,N_33355,N_30477);
nand U41168 (N_41168,N_34689,N_38884);
and U41169 (N_41169,N_36055,N_32770);
or U41170 (N_41170,N_31238,N_35620);
nor U41171 (N_41171,N_37773,N_32312);
xor U41172 (N_41172,N_37227,N_32641);
nand U41173 (N_41173,N_32783,N_37570);
nor U41174 (N_41174,N_39472,N_38539);
xnor U41175 (N_41175,N_31020,N_30807);
nand U41176 (N_41176,N_33203,N_38510);
and U41177 (N_41177,N_36241,N_31446);
xnor U41178 (N_41178,N_34958,N_37658);
xnor U41179 (N_41179,N_32968,N_32755);
nand U41180 (N_41180,N_34229,N_39757);
nand U41181 (N_41181,N_33431,N_36911);
nand U41182 (N_41182,N_34690,N_32407);
xor U41183 (N_41183,N_39114,N_36317);
and U41184 (N_41184,N_31690,N_38794);
nor U41185 (N_41185,N_33408,N_37117);
xor U41186 (N_41186,N_36876,N_34233);
xnor U41187 (N_41187,N_35602,N_32769);
and U41188 (N_41188,N_36454,N_35457);
nand U41189 (N_41189,N_31186,N_38997);
xor U41190 (N_41190,N_30728,N_39652);
nand U41191 (N_41191,N_34842,N_33220);
nand U41192 (N_41192,N_32155,N_35346);
or U41193 (N_41193,N_30758,N_37273);
nand U41194 (N_41194,N_38994,N_37993);
xnor U41195 (N_41195,N_34019,N_32941);
or U41196 (N_41196,N_31413,N_35460);
xor U41197 (N_41197,N_35769,N_39003);
and U41198 (N_41198,N_37427,N_30890);
nor U41199 (N_41199,N_33116,N_34570);
xnor U41200 (N_41200,N_35812,N_37859);
xor U41201 (N_41201,N_36626,N_35014);
and U41202 (N_41202,N_35360,N_33415);
and U41203 (N_41203,N_30461,N_31039);
and U41204 (N_41204,N_31689,N_37908);
or U41205 (N_41205,N_32175,N_34287);
xnor U41206 (N_41206,N_32523,N_31510);
xnor U41207 (N_41207,N_35027,N_39037);
xnor U41208 (N_41208,N_33517,N_31669);
or U41209 (N_41209,N_30101,N_31258);
and U41210 (N_41210,N_32906,N_32868);
nor U41211 (N_41211,N_38829,N_35164);
xor U41212 (N_41212,N_31705,N_35316);
and U41213 (N_41213,N_39327,N_32855);
xnor U41214 (N_41214,N_32088,N_34684);
and U41215 (N_41215,N_37385,N_34730);
nor U41216 (N_41216,N_39422,N_38447);
or U41217 (N_41217,N_35642,N_39175);
nand U41218 (N_41218,N_30226,N_33535);
and U41219 (N_41219,N_32474,N_35862);
or U41220 (N_41220,N_39992,N_34385);
nand U41221 (N_41221,N_39822,N_36279);
nor U41222 (N_41222,N_36558,N_35421);
nor U41223 (N_41223,N_35043,N_32675);
nor U41224 (N_41224,N_31735,N_30258);
or U41225 (N_41225,N_36433,N_35023);
and U41226 (N_41226,N_39549,N_32841);
nor U41227 (N_41227,N_35062,N_30524);
nand U41228 (N_41228,N_39028,N_39797);
and U41229 (N_41229,N_36880,N_38919);
xnor U41230 (N_41230,N_34547,N_32549);
or U41231 (N_41231,N_33473,N_39135);
or U41232 (N_41232,N_30116,N_38778);
xnor U41233 (N_41233,N_31940,N_31467);
nor U41234 (N_41234,N_32696,N_39491);
and U41235 (N_41235,N_33327,N_37605);
xnor U41236 (N_41236,N_39011,N_35361);
xor U41237 (N_41237,N_31788,N_34994);
or U41238 (N_41238,N_33527,N_37751);
nor U41239 (N_41239,N_32300,N_31421);
nand U41240 (N_41240,N_31854,N_38435);
nor U41241 (N_41241,N_30348,N_31366);
nand U41242 (N_41242,N_32843,N_38488);
xnor U41243 (N_41243,N_31543,N_34176);
and U41244 (N_41244,N_30306,N_31785);
nor U41245 (N_41245,N_37409,N_37498);
nand U41246 (N_41246,N_38323,N_31268);
nor U41247 (N_41247,N_32924,N_31461);
xor U41248 (N_41248,N_37638,N_34284);
nor U41249 (N_41249,N_34224,N_38845);
xnor U41250 (N_41250,N_39584,N_35130);
nor U41251 (N_41251,N_35527,N_36569);
xnor U41252 (N_41252,N_34925,N_34894);
nor U41253 (N_41253,N_31144,N_33421);
nor U41254 (N_41254,N_30372,N_31245);
and U41255 (N_41255,N_34500,N_33981);
and U41256 (N_41256,N_36377,N_32143);
nand U41257 (N_41257,N_35223,N_36769);
nor U41258 (N_41258,N_34416,N_38293);
nor U41259 (N_41259,N_32984,N_35867);
and U41260 (N_41260,N_37617,N_39744);
nand U41261 (N_41261,N_37752,N_31444);
nor U41262 (N_41262,N_37083,N_30859);
or U41263 (N_41263,N_37932,N_36436);
and U41264 (N_41264,N_38223,N_38603);
and U41265 (N_41265,N_30026,N_34490);
nor U41266 (N_41266,N_38295,N_37913);
nor U41267 (N_41267,N_39438,N_34511);
nand U41268 (N_41268,N_39183,N_30617);
or U41269 (N_41269,N_39607,N_37517);
and U41270 (N_41270,N_31862,N_33051);
nor U41271 (N_41271,N_39902,N_39809);
and U41272 (N_41272,N_35598,N_39025);
nor U41273 (N_41273,N_33684,N_39356);
nand U41274 (N_41274,N_34938,N_35063);
nor U41275 (N_41275,N_37421,N_30588);
xnor U41276 (N_41276,N_33954,N_31584);
nor U41277 (N_41277,N_32877,N_39548);
or U41278 (N_41278,N_35041,N_38660);
xor U41279 (N_41279,N_39499,N_30903);
or U41280 (N_41280,N_33307,N_35409);
and U41281 (N_41281,N_38095,N_38362);
xnor U41282 (N_41282,N_35388,N_34045);
xnor U41283 (N_41283,N_33448,N_32753);
nand U41284 (N_41284,N_34305,N_37031);
nor U41285 (N_41285,N_39889,N_37756);
or U41286 (N_41286,N_32733,N_32488);
nand U41287 (N_41287,N_35606,N_37068);
nor U41288 (N_41288,N_37065,N_31436);
xnor U41289 (N_41289,N_38992,N_31558);
xnor U41290 (N_41290,N_39986,N_39752);
and U41291 (N_41291,N_30047,N_35942);
xor U41292 (N_41292,N_38506,N_30170);
nand U41293 (N_41293,N_34741,N_35337);
nand U41294 (N_41294,N_30978,N_34984);
nor U41295 (N_41295,N_30228,N_39254);
nor U41296 (N_41296,N_31392,N_39381);
nand U41297 (N_41297,N_36504,N_35058);
nand U41298 (N_41298,N_33603,N_39711);
nand U41299 (N_41299,N_37653,N_36709);
xor U41300 (N_41300,N_32620,N_31310);
xor U41301 (N_41301,N_31814,N_38897);
nor U41302 (N_41302,N_39439,N_34620);
xnor U41303 (N_41303,N_30286,N_32259);
xnor U41304 (N_41304,N_33392,N_32324);
xor U41305 (N_41305,N_31071,N_37301);
nor U41306 (N_41306,N_34346,N_39746);
xor U41307 (N_41307,N_39352,N_38236);
nand U41308 (N_41308,N_32463,N_37719);
xor U41309 (N_41309,N_32989,N_37054);
and U41310 (N_41310,N_37354,N_38995);
xor U41311 (N_41311,N_34959,N_30213);
nand U41312 (N_41312,N_31194,N_31549);
or U41313 (N_41313,N_35020,N_39271);
or U41314 (N_41314,N_30112,N_39838);
and U41315 (N_41315,N_31435,N_30096);
xor U41316 (N_41316,N_33492,N_35870);
and U41317 (N_41317,N_33402,N_35946);
nor U41318 (N_41318,N_30853,N_39745);
or U41319 (N_41319,N_31099,N_32919);
nand U41320 (N_41320,N_34654,N_33118);
nand U41321 (N_41321,N_34362,N_35962);
nand U41322 (N_41322,N_30868,N_30619);
xor U41323 (N_41323,N_36283,N_31271);
and U41324 (N_41324,N_39190,N_33166);
xor U41325 (N_41325,N_31110,N_31649);
and U41326 (N_41326,N_30942,N_34195);
nand U41327 (N_41327,N_38010,N_35428);
nor U41328 (N_41328,N_37802,N_30529);
xor U41329 (N_41329,N_38297,N_36686);
or U41330 (N_41330,N_32363,N_37983);
xnor U41331 (N_41331,N_32082,N_38478);
or U41332 (N_41332,N_30092,N_31257);
nand U41333 (N_41333,N_34610,N_38242);
nor U41334 (N_41334,N_31042,N_31586);
and U41335 (N_41335,N_31560,N_39464);
nand U41336 (N_41336,N_32328,N_32340);
xor U41337 (N_41337,N_33855,N_37468);
and U41338 (N_41338,N_34463,N_37237);
xor U41339 (N_41339,N_36883,N_34168);
xor U41340 (N_41340,N_39847,N_37551);
nand U41341 (N_41341,N_38858,N_36328);
and U41342 (N_41342,N_33959,N_30020);
or U41343 (N_41343,N_36866,N_30558);
or U41344 (N_41344,N_33752,N_35704);
or U41345 (N_41345,N_34393,N_31532);
nor U41346 (N_41346,N_39925,N_30894);
and U41347 (N_41347,N_39799,N_39828);
nand U41348 (N_41348,N_35566,N_35837);
and U41349 (N_41349,N_35648,N_35789);
nor U41350 (N_41350,N_35111,N_39832);
or U41351 (N_41351,N_34004,N_30574);
nand U41352 (N_41352,N_39588,N_33371);
nor U41353 (N_41353,N_34765,N_39128);
xor U41354 (N_41354,N_35234,N_35135);
or U41355 (N_41355,N_35284,N_34024);
xnor U41356 (N_41356,N_37922,N_35725);
xor U41357 (N_41357,N_36590,N_39862);
nor U41358 (N_41358,N_36442,N_38266);
nor U41359 (N_41359,N_30845,N_30822);
nor U41360 (N_41360,N_35816,N_31540);
xor U41361 (N_41361,N_34685,N_36802);
or U41362 (N_41362,N_33186,N_39556);
xnor U41363 (N_41363,N_31939,N_33039);
and U41364 (N_41364,N_35351,N_31566);
nor U41365 (N_41365,N_30272,N_30142);
xnor U41366 (N_41366,N_34388,N_36161);
and U41367 (N_41367,N_37976,N_30856);
nor U41368 (N_41368,N_35554,N_31437);
nor U41369 (N_41369,N_33762,N_32888);
and U41370 (N_41370,N_34595,N_34143);
nand U41371 (N_41371,N_31126,N_31781);
nand U41372 (N_41372,N_34857,N_32427);
or U41373 (N_41373,N_38825,N_30177);
nand U41374 (N_41374,N_39178,N_37994);
and U41375 (N_41375,N_37684,N_33632);
nand U41376 (N_41376,N_34227,N_37533);
nand U41377 (N_41377,N_34960,N_38302);
or U41378 (N_41378,N_32220,N_35304);
and U41379 (N_41379,N_38988,N_33258);
or U41380 (N_41380,N_32228,N_35094);
or U41381 (N_41381,N_38219,N_31687);
or U41382 (N_41382,N_31585,N_30255);
and U41383 (N_41383,N_39754,N_36278);
nand U41384 (N_41384,N_30720,N_36764);
xnor U41385 (N_41385,N_36189,N_33713);
nand U41386 (N_41386,N_39119,N_37192);
nor U41387 (N_41387,N_31590,N_31166);
nand U41388 (N_41388,N_35792,N_38962);
nor U41389 (N_41389,N_37732,N_31926);
or U41390 (N_41390,N_34964,N_35196);
xor U41391 (N_41391,N_36578,N_31513);
and U41392 (N_41392,N_39810,N_31122);
nor U41393 (N_41393,N_35920,N_39785);
xor U41394 (N_41394,N_38769,N_30391);
nand U41395 (N_41395,N_38159,N_39000);
nand U41396 (N_41396,N_35120,N_30234);
xor U41397 (N_41397,N_34657,N_32335);
nand U41398 (N_41398,N_31563,N_30344);
xnor U41399 (N_41399,N_34336,N_35271);
nor U41400 (N_41400,N_33644,N_33315);
nand U41401 (N_41401,N_32680,N_30535);
nor U41402 (N_41402,N_30282,N_36598);
xor U41403 (N_41403,N_30838,N_30119);
nor U41404 (N_41404,N_34133,N_31441);
nor U41405 (N_41405,N_32355,N_39872);
and U41406 (N_41406,N_31674,N_31806);
xnor U41407 (N_41407,N_38680,N_34953);
xnor U41408 (N_41408,N_30568,N_32825);
or U41409 (N_41409,N_38143,N_35517);
or U41410 (N_41410,N_35582,N_33305);
nand U41411 (N_41411,N_31805,N_35263);
and U41412 (N_41412,N_33277,N_35880);
and U41413 (N_41413,N_30161,N_38935);
nand U41414 (N_41414,N_35061,N_37014);
nor U41415 (N_41415,N_32822,N_30085);
nor U41416 (N_41416,N_31215,N_32594);
and U41417 (N_41417,N_31773,N_39559);
or U41418 (N_41418,N_36391,N_32764);
and U41419 (N_41419,N_36846,N_30989);
nor U41420 (N_41420,N_34068,N_33433);
xor U41421 (N_41421,N_39511,N_30964);
and U41422 (N_41422,N_30763,N_37849);
xor U41423 (N_41423,N_36371,N_31625);
or U41424 (N_41424,N_33820,N_38779);
and U41425 (N_41425,N_36841,N_32918);
or U41426 (N_41426,N_38930,N_32718);
or U41427 (N_41427,N_33199,N_31066);
xnor U41428 (N_41428,N_31074,N_37984);
nand U41429 (N_41429,N_37268,N_39918);
or U41430 (N_41430,N_31998,N_32644);
nor U41431 (N_41431,N_32607,N_31303);
and U41432 (N_41432,N_36077,N_39946);
or U41433 (N_41433,N_33991,N_38262);
xor U41434 (N_41434,N_37208,N_36095);
xor U41435 (N_41435,N_30723,N_35124);
and U41436 (N_41436,N_32079,N_35520);
or U41437 (N_41437,N_32443,N_31780);
xnor U41438 (N_41438,N_34766,N_39968);
and U41439 (N_41439,N_39857,N_39563);
or U41440 (N_41440,N_36352,N_33157);
nand U41441 (N_41441,N_35869,N_31329);
nor U41442 (N_41442,N_30645,N_38559);
or U41443 (N_41443,N_35757,N_31588);
nand U41444 (N_41444,N_38085,N_30591);
nand U41445 (N_41445,N_39496,N_31338);
nand U41446 (N_41446,N_37718,N_38841);
nand U41447 (N_41447,N_39961,N_37345);
nand U41448 (N_41448,N_30613,N_30360);
or U41449 (N_41449,N_30927,N_34080);
or U41450 (N_41450,N_35400,N_37250);
nand U41451 (N_41451,N_31250,N_34274);
and U41452 (N_41452,N_36964,N_37381);
nand U41453 (N_41453,N_39210,N_38872);
or U41454 (N_41454,N_37602,N_34805);
and U41455 (N_41455,N_35504,N_38743);
nand U41456 (N_41456,N_35754,N_38760);
nand U41457 (N_41457,N_38424,N_37067);
or U41458 (N_41458,N_34717,N_39391);
xor U41459 (N_41459,N_37155,N_31140);
and U41460 (N_41460,N_36865,N_32357);
or U41461 (N_41461,N_36478,N_32221);
and U41462 (N_41462,N_31472,N_31849);
nor U41463 (N_41463,N_31723,N_36056);
nor U41464 (N_41464,N_38796,N_30311);
nand U41465 (N_41465,N_30675,N_38726);
or U41466 (N_41466,N_31685,N_34650);
and U41467 (N_41467,N_36086,N_38480);
xnor U41468 (N_41468,N_34073,N_32388);
nand U41469 (N_41469,N_31014,N_33141);
or U41470 (N_41470,N_39304,N_32416);
and U41471 (N_41471,N_39945,N_39722);
or U41472 (N_41472,N_39448,N_37492);
nor U41473 (N_41473,N_38643,N_38720);
and U41474 (N_41474,N_34557,N_34396);
or U41475 (N_41475,N_38972,N_37386);
and U41476 (N_41476,N_37024,N_32894);
or U41477 (N_41477,N_39649,N_39904);
or U41478 (N_41478,N_32887,N_34152);
nand U41479 (N_41479,N_30071,N_33278);
nor U41480 (N_41480,N_32990,N_30328);
and U41481 (N_41481,N_31729,N_36326);
or U41482 (N_41482,N_30266,N_33001);
xor U41483 (N_41483,N_39132,N_32017);
nor U41484 (N_41484,N_37376,N_30202);
or U41485 (N_41485,N_30785,N_33454);
xnor U41486 (N_41486,N_31449,N_31024);
nor U41487 (N_41487,N_37497,N_31183);
xor U41488 (N_41488,N_30704,N_32356);
or U41489 (N_41489,N_31650,N_34587);
nor U41490 (N_41490,N_30287,N_32231);
nor U41491 (N_41491,N_33718,N_37348);
xnor U41492 (N_41492,N_32652,N_31294);
nand U41493 (N_41493,N_32756,N_39935);
nor U41494 (N_41494,N_34863,N_32522);
xor U41495 (N_41495,N_32494,N_34468);
nor U41496 (N_41496,N_34665,N_34965);
nor U41497 (N_41497,N_34415,N_32104);
nand U41498 (N_41498,N_36378,N_33745);
and U41499 (N_41499,N_30334,N_32993);
nor U41500 (N_41500,N_34200,N_34574);
and U41501 (N_41501,N_31325,N_35494);
and U41502 (N_41502,N_32881,N_30046);
nand U41503 (N_41503,N_35663,N_39279);
or U41504 (N_41504,N_36152,N_37946);
nand U41505 (N_41505,N_36844,N_30994);
nand U41506 (N_41506,N_36896,N_35761);
and U41507 (N_41507,N_38614,N_32587);
nand U41508 (N_41508,N_36027,N_35364);
nand U41509 (N_41509,N_36691,N_33029);
nand U41510 (N_41510,N_36910,N_39141);
nor U41511 (N_41511,N_38182,N_35152);
or U41512 (N_41512,N_31430,N_38909);
nand U41513 (N_41513,N_36470,N_39996);
nor U41514 (N_41514,N_31648,N_34041);
and U41515 (N_41515,N_38414,N_31606);
or U41516 (N_41516,N_37758,N_33539);
or U41517 (N_41517,N_34729,N_35715);
and U41518 (N_41518,N_39302,N_33929);
nor U41519 (N_41519,N_35720,N_37077);
nor U41520 (N_41520,N_30932,N_36897);
nor U41521 (N_41521,N_31632,N_36734);
and U41522 (N_41522,N_38838,N_37176);
xnor U41523 (N_41523,N_38019,N_37791);
or U41524 (N_41524,N_35604,N_36774);
xor U41525 (N_41525,N_31304,N_31131);
and U41526 (N_41526,N_36608,N_35605);
and U41527 (N_41527,N_32685,N_35621);
xor U41528 (N_41528,N_34923,N_39575);
or U41529 (N_41529,N_31113,N_35483);
and U41530 (N_41530,N_33293,N_30624);
nand U41531 (N_41531,N_30532,N_31766);
and U41532 (N_41532,N_39617,N_37446);
or U41533 (N_41533,N_35699,N_35343);
or U41534 (N_41534,N_34478,N_37554);
and U41535 (N_41535,N_31402,N_30876);
or U41536 (N_41536,N_33440,N_33188);
nand U41537 (N_41537,N_31709,N_36116);
and U41538 (N_41538,N_36343,N_31169);
and U41539 (N_41539,N_37505,N_34314);
or U41540 (N_41540,N_33687,N_32021);
and U41541 (N_41541,N_34861,N_37516);
nand U41542 (N_41542,N_33771,N_32592);
nand U41543 (N_41543,N_35103,N_35122);
nor U41544 (N_41544,N_36112,N_30322);
nor U41545 (N_41545,N_34727,N_30753);
or U41546 (N_41546,N_36347,N_39734);
nor U41547 (N_41547,N_36635,N_37835);
nor U41548 (N_41548,N_30559,N_32849);
xnor U41549 (N_41549,N_31820,N_30261);
nand U41550 (N_41550,N_33236,N_30926);
xnor U41551 (N_41551,N_33595,N_30637);
and U41552 (N_41552,N_32901,N_30695);
nor U41553 (N_41553,N_34577,N_36221);
or U41554 (N_41554,N_38593,N_30082);
or U41555 (N_41555,N_34462,N_34832);
and U41556 (N_41556,N_38240,N_32905);
xnor U41557 (N_41557,N_35721,N_36560);
or U41558 (N_41558,N_38401,N_30726);
or U41559 (N_41559,N_34548,N_33164);
nand U41560 (N_41560,N_39692,N_38703);
nor U41561 (N_41561,N_37944,N_36571);
nor U41562 (N_41562,N_36776,N_33798);
or U41563 (N_41563,N_31772,N_31594);
nor U41564 (N_41564,N_31242,N_33223);
and U41565 (N_41565,N_31035,N_34236);
nor U41566 (N_41566,N_33495,N_35758);
and U41567 (N_41567,N_32944,N_38776);
nor U41568 (N_41568,N_38163,N_30478);
nand U41569 (N_41569,N_30199,N_34505);
nand U41570 (N_41570,N_31921,N_35624);
nor U41571 (N_41571,N_37831,N_35985);
and U41572 (N_41572,N_31878,N_30698);
nor U41573 (N_41573,N_33911,N_33640);
nor U41574 (N_41574,N_34148,N_32614);
and U41575 (N_41575,N_39177,N_37407);
xor U41576 (N_41576,N_31787,N_30871);
xnor U41577 (N_41577,N_33777,N_38246);
xor U41578 (N_41578,N_37448,N_36119);
and U41579 (N_41579,N_35526,N_31448);
nor U41580 (N_41580,N_31811,N_36658);
or U41581 (N_41581,N_38587,N_38108);
xor U41582 (N_41582,N_39165,N_35714);
nor U41583 (N_41583,N_39536,N_35095);
xor U41584 (N_41584,N_34714,N_35551);
or U41585 (N_41585,N_37495,N_37121);
and U41586 (N_41586,N_30860,N_36301);
nand U41587 (N_41587,N_30526,N_34189);
xor U41588 (N_41588,N_38787,N_31796);
or U41589 (N_41589,N_35051,N_36629);
nand U41590 (N_41590,N_38287,N_30543);
nor U41591 (N_41591,N_30450,N_34614);
nor U41592 (N_41592,N_32188,N_36518);
nor U41593 (N_41593,N_35855,N_39091);
xor U41594 (N_41594,N_36102,N_34178);
nor U41595 (N_41595,N_31121,N_33764);
and U41596 (N_41596,N_38699,N_34885);
and U41597 (N_41597,N_31994,N_35802);
and U41598 (N_41598,N_38940,N_37349);
and U41599 (N_41599,N_32223,N_33881);
xor U41600 (N_41600,N_38523,N_32466);
xnor U41601 (N_41601,N_39613,N_32374);
or U41602 (N_41602,N_33253,N_39628);
or U41603 (N_41603,N_36235,N_34440);
xor U41604 (N_41604,N_30548,N_36410);
or U41605 (N_41605,N_33546,N_34600);
nor U41606 (N_41606,N_34853,N_39344);
nand U41607 (N_41607,N_30583,N_35727);
nor U41608 (N_41608,N_36871,N_37363);
or U41609 (N_41609,N_30593,N_31481);
xor U41610 (N_41610,N_37696,N_31556);
and U41611 (N_41611,N_38684,N_36013);
nand U41612 (N_41612,N_33707,N_37523);
nand U41613 (N_41613,N_32767,N_34715);
or U41614 (N_41614,N_30840,N_37286);
nand U41615 (N_41615,N_32551,N_31643);
nor U41616 (N_41616,N_36994,N_35215);
nand U41617 (N_41617,N_32140,N_33990);
nor U41618 (N_41618,N_33462,N_37578);
or U41619 (N_41619,N_34592,N_37650);
or U41620 (N_41620,N_31524,N_34014);
xor U41621 (N_41621,N_30823,N_39292);
nand U41622 (N_41622,N_32107,N_30508);
nand U41623 (N_41623,N_34780,N_30632);
and U41624 (N_41624,N_32668,N_35435);
and U41625 (N_41625,N_33383,N_35750);
nor U41626 (N_41626,N_32574,N_32049);
or U41627 (N_41627,N_38999,N_30651);
nand U41628 (N_41628,N_36587,N_30392);
or U41629 (N_41629,N_30406,N_36271);
xnor U41630 (N_41630,N_30447,N_30705);
xor U41631 (N_41631,N_36815,N_39789);
xor U41632 (N_41632,N_38709,N_35198);
or U41633 (N_41633,N_33677,N_31164);
or U41634 (N_41634,N_32762,N_37225);
or U41635 (N_41635,N_38306,N_37734);
nand U41636 (N_41636,N_34758,N_31997);
nand U41637 (N_41637,N_37781,N_36992);
xor U41638 (N_41638,N_30846,N_36032);
nor U41639 (N_41639,N_32381,N_33218);
xor U41640 (N_41640,N_33803,N_32400);
nor U41641 (N_41641,N_31990,N_36541);
or U41642 (N_41642,N_37512,N_37975);
xor U41643 (N_41643,N_37013,N_34736);
nor U41644 (N_41644,N_37544,N_38111);
or U41645 (N_41645,N_34147,N_34697);
or U41646 (N_41646,N_34488,N_35079);
and U41647 (N_41647,N_35516,N_37474);
xnor U41648 (N_41648,N_30444,N_35046);
nor U41649 (N_41649,N_35824,N_37458);
nand U41650 (N_41650,N_30480,N_31137);
xnor U41651 (N_41651,N_39142,N_39720);
and U41652 (N_41652,N_31438,N_35333);
nor U41653 (N_41653,N_39796,N_30074);
xnor U41654 (N_41654,N_31863,N_30677);
and U41655 (N_41655,N_31227,N_33927);
nor U41656 (N_41656,N_31561,N_34380);
and U41657 (N_41657,N_37183,N_39713);
xnor U41658 (N_41658,N_35086,N_30638);
and U41659 (N_41659,N_30671,N_32880);
or U41660 (N_41660,N_34386,N_32605);
nand U41661 (N_41661,N_33657,N_37757);
nor U41662 (N_41662,N_36551,N_35153);
nand U41663 (N_41663,N_33715,N_35359);
nand U41664 (N_41664,N_33741,N_36854);
or U41665 (N_41665,N_34095,N_35557);
or U41666 (N_41666,N_30370,N_36932);
nor U41667 (N_41667,N_39803,N_39232);
nor U41668 (N_41668,N_38578,N_30691);
or U41669 (N_41669,N_32470,N_37525);
nor U41670 (N_41670,N_39712,N_37588);
nor U41671 (N_41671,N_38404,N_38721);
nand U41672 (N_41672,N_37205,N_37845);
xnor U41673 (N_41673,N_32634,N_39571);
nand U41674 (N_41674,N_32454,N_31036);
nor U41675 (N_41675,N_32262,N_33358);
or U41676 (N_41676,N_34077,N_35635);
nand U41677 (N_41677,N_33664,N_36450);
or U41678 (N_41678,N_36054,N_38623);
nor U41679 (N_41679,N_34816,N_30804);
and U41680 (N_41680,N_38113,N_34948);
or U41681 (N_41681,N_39929,N_38691);
or U41682 (N_41682,N_39048,N_36809);
nor U41683 (N_41683,N_37142,N_32018);
or U41684 (N_41684,N_36310,N_39019);
nand U41685 (N_41685,N_37447,N_36006);
nor U41686 (N_41686,N_31609,N_39909);
xnor U41687 (N_41687,N_37856,N_38611);
or U41688 (N_41688,N_34999,N_32850);
or U41689 (N_41689,N_33606,N_36707);
or U41690 (N_41690,N_33862,N_35665);
and U41691 (N_41691,N_36210,N_37555);
nand U41692 (N_41692,N_39620,N_32508);
or U41693 (N_41693,N_33366,N_36960);
nand U41694 (N_41694,N_32732,N_36431);
nor U41695 (N_41695,N_34982,N_31515);
xnor U41696 (N_41696,N_38864,N_35390);
xor U41697 (N_41697,N_30222,N_37399);
xor U41698 (N_41698,N_37842,N_33074);
or U41699 (N_41699,N_30789,N_38619);
nand U41700 (N_41700,N_38859,N_38407);
and U41701 (N_41701,N_31249,N_30495);
xor U41702 (N_41702,N_36071,N_33224);
and U41703 (N_41703,N_33997,N_39362);
xnor U41704 (N_41704,N_32816,N_33950);
and U41705 (N_41705,N_34184,N_38928);
and U41706 (N_41706,N_32398,N_30744);
nor U41707 (N_41707,N_30059,N_30494);
and U41708 (N_41708,N_36875,N_37825);
xor U41709 (N_41709,N_35623,N_38332);
and U41710 (N_41710,N_38380,N_35894);
nor U41711 (N_41711,N_31343,N_34476);
or U41712 (N_41712,N_30037,N_39443);
xor U41713 (N_41713,N_33137,N_34329);
nor U41714 (N_41714,N_33775,N_34864);
or U41715 (N_41715,N_37064,N_38770);
nand U41716 (N_41716,N_36942,N_35784);
nor U41717 (N_41717,N_39683,N_35004);
or U41718 (N_41718,N_37634,N_31440);
and U41719 (N_41719,N_38675,N_30700);
and U41720 (N_41720,N_34726,N_34282);
and U41721 (N_41721,N_34516,N_30982);
nand U41722 (N_41722,N_36923,N_38296);
and U41723 (N_41723,N_31114,N_34991);
nor U41724 (N_41724,N_36358,N_38147);
xor U41725 (N_41725,N_39670,N_37403);
or U41726 (N_41726,N_35974,N_35690);
xor U41727 (N_41727,N_37909,N_39678);
xnor U41728 (N_41728,N_37254,N_33352);
or U41729 (N_41729,N_35370,N_36023);
nand U41730 (N_41730,N_33946,N_31011);
nor U41731 (N_41731,N_31985,N_30369);
nor U41732 (N_41732,N_32543,N_32048);
nand U41733 (N_41733,N_39887,N_39673);
or U41734 (N_41734,N_33312,N_31619);
xor U41735 (N_41735,N_36593,N_39818);
nand U41736 (N_41736,N_33465,N_30735);
and U41737 (N_41737,N_39614,N_39361);
and U41738 (N_41738,N_38130,N_37504);
xor U41739 (N_41739,N_39370,N_33967);
and U41740 (N_41740,N_34759,N_30551);
nor U41741 (N_41741,N_37431,N_37123);
and U41742 (N_41742,N_33416,N_34477);
nand U41743 (N_41743,N_38059,N_32844);
nor U41744 (N_41744,N_38500,N_33957);
or U41745 (N_41745,N_37729,N_33463);
or U41746 (N_41746,N_33248,N_30724);
and U41747 (N_41747,N_33768,N_33102);
nand U41748 (N_41748,N_33797,N_30709);
and U41749 (N_41749,N_38628,N_37319);
and U41750 (N_41750,N_37731,N_37917);
nand U41751 (N_41751,N_30268,N_30325);
xnor U41752 (N_41752,N_39266,N_32633);
nand U41753 (N_41753,N_38767,N_38226);
or U41754 (N_41754,N_31120,N_33699);
nand U41755 (N_41755,N_32576,N_37971);
xnor U41756 (N_41756,N_38331,N_36186);
nor U41757 (N_41757,N_31905,N_35912);
nor U41758 (N_41758,N_34208,N_31462);
or U41759 (N_41759,N_30109,N_32192);
or U41760 (N_41760,N_35186,N_38324);
nand U41761 (N_41761,N_35865,N_36337);
xor U41762 (N_41762,N_39475,N_32402);
and U41763 (N_41763,N_31571,N_33610);
nor U41764 (N_41764,N_31334,N_30790);
nand U41765 (N_41765,N_30058,N_34710);
xnor U41766 (N_41766,N_31683,N_30206);
and U41767 (N_41767,N_36799,N_34374);
xor U41768 (N_41768,N_37661,N_33350);
and U41769 (N_41769,N_33774,N_31087);
or U41770 (N_41770,N_37181,N_30288);
nand U41771 (N_41771,N_39473,N_34802);
xnor U41772 (N_41772,N_33301,N_30451);
and U41773 (N_41773,N_36703,N_39377);
or U41774 (N_41774,N_34860,N_34775);
and U41775 (N_41775,N_33837,N_35728);
or U41776 (N_41776,N_36409,N_36303);
or U41777 (N_41777,N_34880,N_39731);
xor U41778 (N_41778,N_30609,N_38303);
nand U41779 (N_41779,N_35616,N_36821);
and U41780 (N_41780,N_34612,N_36934);
nand U41781 (N_41781,N_35206,N_34177);
xnor U41782 (N_41782,N_38638,N_35825);
and U41783 (N_41783,N_36212,N_36684);
nor U41784 (N_41784,N_30906,N_38261);
and U41785 (N_41785,N_30764,N_32361);
xnor U41786 (N_41786,N_36427,N_34538);
and U41787 (N_41787,N_33367,N_30169);
xnor U41788 (N_41788,N_30235,N_30834);
xor U41789 (N_41789,N_36322,N_39474);
nor U41790 (N_41790,N_37539,N_30021);
xor U41791 (N_41791,N_39657,N_33306);
nor U41792 (N_41792,N_34315,N_36733);
or U41793 (N_41793,N_31426,N_39610);
nand U41794 (N_41794,N_35335,N_32706);
xor U41795 (N_41795,N_33121,N_37678);
nand U41796 (N_41796,N_31048,N_37877);
xor U41797 (N_41797,N_34967,N_31345);
nor U41798 (N_41798,N_33597,N_39117);
or U41799 (N_41799,N_39465,N_34207);
nor U41800 (N_41800,N_36621,N_35556);
or U41801 (N_41801,N_30749,N_38137);
nor U41802 (N_41802,N_36533,N_30569);
nor U41803 (N_41803,N_34260,N_38953);
or U41804 (N_41804,N_38498,N_30835);
xor U41805 (N_41805,N_37310,N_33227);
or U41806 (N_41806,N_35380,N_38651);
and U41807 (N_41807,N_36018,N_33556);
or U41808 (N_41808,N_32243,N_37832);
nand U41809 (N_41809,N_32923,N_33078);
xor U41810 (N_41810,N_35764,N_35317);
and U41811 (N_41811,N_39641,N_33939);
nor U41812 (N_41812,N_31388,N_30308);
xnor U41813 (N_41813,N_30686,N_30000);
or U41814 (N_41814,N_30196,N_33679);
xor U41815 (N_41815,N_31535,N_33313);
nor U41816 (N_41816,N_38171,N_34755);
xor U41817 (N_41817,N_38254,N_33835);
and U41818 (N_41818,N_30331,N_38742);
or U41819 (N_41819,N_36060,N_31469);
nand U41820 (N_41820,N_34436,N_30481);
xnor U41821 (N_41821,N_30003,N_35536);
and U41822 (N_41822,N_31947,N_36688);
and U41823 (N_41823,N_35580,N_31263);
or U41824 (N_41824,N_31733,N_38798);
xnor U41825 (N_41825,N_36863,N_36669);
nor U41826 (N_41826,N_34030,N_31344);
nand U41827 (N_41827,N_35847,N_30386);
and U41828 (N_41828,N_38204,N_31447);
or U41829 (N_41829,N_39502,N_30626);
nand U41830 (N_41830,N_37537,N_33395);
xor U41831 (N_41831,N_30186,N_38003);
xor U41832 (N_41832,N_31200,N_35573);
and U41833 (N_41833,N_36007,N_36987);
nand U41834 (N_41834,N_32173,N_32798);
nand U41835 (N_41835,N_34099,N_33870);
or U41836 (N_41836,N_30911,N_37938);
nor U41837 (N_41837,N_36092,N_39831);
nand U41838 (N_41838,N_39521,N_37135);
nand U41839 (N_41839,N_32087,N_37171);
and U41840 (N_41840,N_36628,N_38863);
nor U41841 (N_41841,N_38196,N_38946);
or U41842 (N_41842,N_32851,N_33602);
xnor U41843 (N_41843,N_39585,N_32848);
nor U41844 (N_41844,N_39022,N_32609);
nand U41845 (N_41845,N_34225,N_38107);
nand U41846 (N_41846,N_37412,N_31808);
or U41847 (N_41847,N_34290,N_39938);
xnor U41848 (N_41848,N_32760,N_39120);
nand U41849 (N_41849,N_39985,N_32141);
nand U41850 (N_41850,N_35268,N_30301);
or U41851 (N_41851,N_33373,N_32562);
xnor U41852 (N_41852,N_38012,N_30570);
nand U41853 (N_41853,N_34125,N_34786);
or U41854 (N_41854,N_30443,N_35117);
nand U41855 (N_41855,N_35888,N_31081);
nand U41856 (N_41856,N_37480,N_33642);
xor U41857 (N_41857,N_37788,N_31911);
nand U41858 (N_41858,N_34582,N_34611);
nor U41859 (N_41859,N_36177,N_38280);
xnor U41860 (N_41860,N_36920,N_35872);
or U41861 (N_41861,N_34151,N_39784);
nor U41862 (N_41862,N_38865,N_38610);
or U41863 (N_41863,N_33627,N_31503);
or U41864 (N_41864,N_36677,N_32854);
xor U41865 (N_41865,N_39065,N_38959);
nor U41866 (N_41866,N_30941,N_37963);
nand U41867 (N_41867,N_37672,N_32276);
and U41868 (N_41868,N_33935,N_37355);
xnor U41869 (N_41869,N_37242,N_34387);
and U41870 (N_41870,N_31159,N_32359);
xnor U41871 (N_41871,N_37299,N_35835);
and U41872 (N_41872,N_33240,N_31170);
nand U41873 (N_41873,N_32635,N_34683);
nor U41874 (N_41874,N_30509,N_39927);
nor U41875 (N_41875,N_35745,N_35710);
and U41876 (N_41876,N_34762,N_35801);
or U41877 (N_41877,N_31357,N_37430);
nand U41878 (N_41878,N_38387,N_33036);
xor U41879 (N_41879,N_33235,N_30669);
and U41880 (N_41880,N_34131,N_39740);
and U41881 (N_41881,N_34012,N_36130);
or U41882 (N_41882,N_33061,N_34737);
xor U41883 (N_41883,N_30786,N_33737);
and U41884 (N_41884,N_31943,N_36004);
and U41885 (N_41885,N_34771,N_35260);
and U41886 (N_41886,N_39783,N_32707);
xor U41887 (N_41887,N_32490,N_34201);
nor U41888 (N_41888,N_34312,N_37196);
nor U41889 (N_41889,N_39668,N_36392);
nor U41890 (N_41890,N_38915,N_39898);
nand U41891 (N_41891,N_33388,N_33052);
or U41892 (N_41892,N_38615,N_34940);
and U41893 (N_41893,N_37895,N_39642);
nor U41894 (N_41894,N_33686,N_39624);
nor U41895 (N_41895,N_34066,N_39858);
and U41896 (N_41896,N_32615,N_35300);
nand U41897 (N_41897,N_32277,N_39775);
xnor U41898 (N_41898,N_36766,N_33932);
and U41899 (N_41899,N_31037,N_34788);
nand U41900 (N_41900,N_31335,N_37652);
or U41901 (N_41901,N_39318,N_39330);
xnor U41902 (N_41902,N_37561,N_35462);
nor U41903 (N_41903,N_30959,N_31891);
xnor U41904 (N_41904,N_31812,N_37478);
and U41905 (N_41905,N_30595,N_39609);
nand U41906 (N_41906,N_35786,N_33441);
nor U41907 (N_41907,N_39285,N_38537);
and U41908 (N_41908,N_39325,N_31956);
xor U41909 (N_41909,N_35280,N_38788);
xor U41910 (N_41910,N_37470,N_30365);
and U41911 (N_41911,N_35434,N_34750);
or U41912 (N_41912,N_39400,N_33853);
nand U41913 (N_41913,N_38397,N_36408);
nand U41914 (N_41914,N_38382,N_35010);
and U41915 (N_41915,N_32763,N_38734);
xor U41916 (N_41916,N_38738,N_32137);
nor U41917 (N_41917,N_31924,N_31234);
or U41918 (N_41918,N_34752,N_39484);
or U41919 (N_41919,N_30891,N_34623);
and U41920 (N_41920,N_38631,N_35185);
nor U41921 (N_41921,N_37833,N_35448);
xor U41922 (N_41922,N_38516,N_32916);
xor U41923 (N_41923,N_37383,N_39121);
or U41924 (N_41924,N_30673,N_33096);
nand U41925 (N_41925,N_31445,N_35179);
nand U41926 (N_41926,N_30528,N_30937);
or U41927 (N_41927,N_34377,N_38243);
nor U41928 (N_41928,N_38679,N_33148);
nor U41929 (N_41929,N_34410,N_31747);
and U41930 (N_41930,N_33142,N_31286);
nand U41931 (N_41931,N_38134,N_34951);
nor U41932 (N_41932,N_34713,N_31059);
nand U41933 (N_41933,N_37303,N_39893);
and U41934 (N_41934,N_37979,N_30875);
xor U41935 (N_41935,N_39395,N_37048);
and U41936 (N_41936,N_31382,N_37180);
nand U41937 (N_41937,N_34773,N_37212);
nor U41938 (N_41938,N_37426,N_32285);
and U41939 (N_41939,N_30038,N_34481);
nand U41940 (N_41940,N_37792,N_36273);
nor U41941 (N_41941,N_39682,N_38124);
nand U41942 (N_41942,N_32485,N_39675);
nand U41943 (N_41943,N_37861,N_30817);
nand U41944 (N_41944,N_32000,N_38433);
nor U41945 (N_41945,N_32293,N_33972);
nand U41946 (N_41946,N_35238,N_33250);
xor U41947 (N_41947,N_35345,N_34008);
nor U41948 (N_41948,N_36219,N_30794);
xor U41949 (N_41949,N_35009,N_32204);
nand U41950 (N_41950,N_35692,N_36545);
or U41951 (N_41951,N_38993,N_35115);
xor U41952 (N_41952,N_38547,N_37248);
or U41953 (N_41953,N_38911,N_39176);
and U41954 (N_41954,N_36239,N_38049);
nand U41955 (N_41955,N_36894,N_39062);
or U41956 (N_41956,N_36110,N_32712);
nand U41957 (N_41957,N_39942,N_32547);
xnor U41958 (N_41958,N_36097,N_30912);
xnor U41959 (N_41959,N_32831,N_38443);
nand U41960 (N_41960,N_30976,N_34083);
nand U41961 (N_41961,N_36610,N_35844);
or U41962 (N_41962,N_34968,N_37334);
nand U41963 (N_41963,N_36851,N_34720);
nor U41964 (N_41964,N_37195,N_31977);
nand U41965 (N_41965,N_30120,N_33266);
or U41966 (N_41966,N_39911,N_39295);
and U41967 (N_41967,N_38586,N_34978);
nor U41968 (N_41968,N_36981,N_32201);
and U41969 (N_41969,N_38169,N_34323);
and U41970 (N_41970,N_32423,N_39966);
nand U41971 (N_41971,N_36903,N_39096);
nor U41972 (N_41972,N_38112,N_32582);
nand U41973 (N_41973,N_35735,N_31710);
and U41974 (N_41974,N_39940,N_34491);
nor U41975 (N_41975,N_39749,N_33071);
or U41976 (N_41976,N_36870,N_35072);
nand U41977 (N_41977,N_30923,N_34166);
nand U41978 (N_41978,N_36318,N_39388);
nor U41979 (N_41979,N_38716,N_33457);
nand U41980 (N_41980,N_35570,N_37168);
or U41981 (N_41981,N_33975,N_33325);
xor U41982 (N_41982,N_38288,N_34226);
or U41983 (N_41983,N_31880,N_31298);
xor U41984 (N_41984,N_38071,N_38337);
nand U41985 (N_41985,N_33903,N_32081);
nand U41986 (N_41986,N_31522,N_37003);
xor U41987 (N_41987,N_39246,N_37313);
or U41988 (N_41988,N_37035,N_38034);
xnor U41989 (N_41989,N_36849,N_38475);
and U41990 (N_41990,N_31117,N_37130);
nor U41991 (N_41991,N_32344,N_34544);
xnor U41992 (N_41992,N_33790,N_38585);
or U41993 (N_41993,N_30546,N_33712);
xnor U41994 (N_41994,N_34013,N_32418);
nor U41995 (N_41995,N_32304,N_33618);
nand U41996 (N_41996,N_38550,N_31975);
and U41997 (N_41997,N_30667,N_32628);
xor U41998 (N_41998,N_36673,N_38563);
and U41999 (N_41999,N_33360,N_32710);
nor U42000 (N_42000,N_36374,N_30681);
or U42001 (N_42001,N_33499,N_39148);
nor U42002 (N_42002,N_37397,N_38238);
or U42003 (N_42003,N_36188,N_38766);
and U42004 (N_42004,N_32774,N_39960);
nor U42005 (N_42005,N_34961,N_39867);
and U42006 (N_42006,N_35254,N_34507);
and U42007 (N_42007,N_30171,N_38975);
xor U42008 (N_42008,N_36202,N_34819);
nand U42009 (N_42009,N_34745,N_31765);
or U42010 (N_42010,N_34897,N_30246);
nand U42011 (N_42011,N_38115,N_32103);
or U42012 (N_42012,N_37269,N_35168);
nand U42013 (N_42013,N_30358,N_35694);
nand U42014 (N_42014,N_37887,N_32101);
xor U42015 (N_42015,N_38465,N_33508);
nor U42016 (N_42016,N_35655,N_30954);
or U42017 (N_42017,N_32501,N_36393);
xnor U42018 (N_42018,N_32278,N_36098);
nand U42019 (N_42019,N_36417,N_32519);
and U42020 (N_42020,N_38007,N_36274);
nor U42021 (N_42021,N_34334,N_35145);
xor U42022 (N_42022,N_36269,N_37607);
nor U42023 (N_42023,N_30482,N_30095);
nand U42024 (N_42024,N_34203,N_38820);
or U42025 (N_42025,N_36586,N_38432);
nand U42026 (N_42026,N_35217,N_31208);
xnor U42027 (N_42027,N_35311,N_31216);
nor U42028 (N_42028,N_35871,N_33868);
or U42029 (N_42029,N_36855,N_39184);
nor U42030 (N_42030,N_37398,N_32512);
or U42031 (N_42031,N_35232,N_33393);
nand U42032 (N_42032,N_36293,N_31247);
and U42033 (N_42033,N_39255,N_36361);
nand U42034 (N_42034,N_36195,N_39449);
and U42035 (N_42035,N_32667,N_30706);
or U42036 (N_42036,N_33509,N_36791);
or U42037 (N_42037,N_34038,N_33645);
and U42038 (N_42038,N_38511,N_36263);
or U42039 (N_42039,N_31184,N_33119);
nand U42040 (N_42040,N_30616,N_33791);
or U42041 (N_42041,N_33064,N_32450);
nand U42042 (N_42042,N_37302,N_34988);
nor U42043 (N_42043,N_31318,N_34011);
nor U42044 (N_42044,N_37300,N_34401);
xor U42045 (N_42045,N_37651,N_34706);
nand U42046 (N_42046,N_35318,N_31573);
or U42047 (N_42047,N_32959,N_30408);
and U42048 (N_42048,N_37215,N_32611);
xnor U42049 (N_42049,N_33030,N_38837);
and U42050 (N_42050,N_31695,N_32118);
nor U42051 (N_42051,N_35441,N_35936);
or U42052 (N_42052,N_34159,N_33466);
xnor U42053 (N_42053,N_37284,N_38194);
xor U42054 (N_42054,N_30928,N_32596);
and U42055 (N_42055,N_38311,N_37271);
xor U42056 (N_42056,N_31688,N_34146);
xor U42057 (N_42057,N_35074,N_39275);
xnor U42058 (N_42058,N_37707,N_30600);
or U42059 (N_42059,N_34769,N_39531);
nand U42060 (N_42060,N_37514,N_30793);
or U42061 (N_42061,N_37910,N_38114);
nand U42062 (N_42062,N_36749,N_36721);
or U42063 (N_42063,N_38202,N_38831);
nand U42064 (N_42064,N_39454,N_34566);
or U42065 (N_42065,N_30668,N_34590);
and U42066 (N_42066,N_33930,N_33124);
nor U42067 (N_42067,N_38951,N_38460);
or U42068 (N_42068,N_34774,N_36375);
nand U42069 (N_42069,N_34498,N_38802);
nand U42070 (N_42070,N_39063,N_31505);
and U42071 (N_42071,N_35645,N_33799);
nor U42072 (N_42072,N_30065,N_36949);
xor U42073 (N_42073,N_37980,N_32447);
xor U42074 (N_42074,N_38757,N_31173);
and U42075 (N_42075,N_37390,N_31254);
nand U42076 (N_42076,N_30983,N_34594);
xor U42077 (N_42077,N_31083,N_38490);
xnor U42078 (N_42078,N_38228,N_34856);
xor U42079 (N_42079,N_38366,N_33483);
and U42080 (N_42080,N_38916,N_30057);
xor U42081 (N_42081,N_36832,N_32878);
or U42082 (N_42082,N_30050,N_38889);
or U42083 (N_42083,N_31913,N_38548);
nor U42084 (N_42084,N_36335,N_37860);
nor U42085 (N_42085,N_33337,N_38482);
nand U42086 (N_42086,N_32566,N_31080);
nor U42087 (N_42087,N_35502,N_35548);
nand U42088 (N_42088,N_38348,N_35419);
nand U42089 (N_42089,N_36253,N_30951);
nor U42090 (N_42090,N_35992,N_39727);
nor U42091 (N_42091,N_30130,N_31866);
or U42092 (N_42092,N_36735,N_33636);
or U42093 (N_42093,N_39425,N_34144);
nor U42094 (N_42094,N_37294,N_30992);
and U42095 (N_42095,N_35873,N_32455);
and U42096 (N_42096,N_35747,N_36699);
and U42097 (N_42097,N_32102,N_34103);
xor U42098 (N_42098,N_39333,N_36348);
or U42099 (N_42099,N_35156,N_30554);
nand U42100 (N_42100,N_30354,N_31128);
nor U42101 (N_42101,N_30747,N_34761);
xor U42102 (N_42102,N_38445,N_31308);
xor U42103 (N_42103,N_36031,N_31859);
nand U42104 (N_42104,N_35118,N_34907);
or U42105 (N_42105,N_37609,N_30962);
or U42106 (N_42106,N_30013,N_37838);
or U42107 (N_42107,N_39505,N_33145);
nor U42108 (N_42108,N_38561,N_32604);
or U42109 (N_42109,N_36701,N_38241);
nor U42110 (N_42110,N_36914,N_35157);
xnor U42111 (N_42111,N_36438,N_39602);
and U42112 (N_42112,N_34205,N_36158);
nand U42113 (N_42113,N_30943,N_38715);
nand U42114 (N_42114,N_39314,N_32595);
or U42115 (N_42115,N_31708,N_31406);
or U42116 (N_42116,N_33909,N_38711);
xnor U42117 (N_42117,N_37688,N_36404);
and U42118 (N_42118,N_34297,N_34124);
or U42119 (N_42119,N_37081,N_34352);
or U42120 (N_42120,N_35006,N_32254);
nand U42121 (N_42121,N_37613,N_35982);
nand U42122 (N_42122,N_32903,N_30381);
nor U42123 (N_42123,N_36881,N_38833);
xnor U42124 (N_42124,N_35488,N_37857);
nand U42125 (N_42125,N_37521,N_38592);
and U42126 (N_42126,N_36552,N_36760);
nand U42127 (N_42127,N_35161,N_35032);
xor U42128 (N_42128,N_33152,N_39086);
or U42129 (N_42129,N_31082,N_37483);
xnor U42130 (N_42130,N_31219,N_34778);
nor U42131 (N_42131,N_39807,N_30813);
nand U42132 (N_42132,N_35656,N_31484);
or U42133 (N_42133,N_33727,N_36176);
and U42134 (N_42134,N_34135,N_32105);
and U42135 (N_42135,N_33986,N_38051);
and U42136 (N_42136,N_36967,N_33910);
or U42137 (N_42137,N_32287,N_30448);
or U42138 (N_42138,N_39770,N_39890);
nand U42139 (N_42139,N_30915,N_31582);
nand U42140 (N_42140,N_37543,N_39237);
or U42141 (N_42141,N_30084,N_32569);
nor U42142 (N_42142,N_33598,N_30596);
or U42143 (N_42143,N_35861,N_37369);
nor U42144 (N_42144,N_37044,N_38199);
xor U42145 (N_42145,N_36051,N_37914);
and U42146 (N_42146,N_38497,N_35429);
nor U42147 (N_42147,N_31262,N_33872);
xor U42148 (N_42148,N_33444,N_36262);
nand U42149 (N_42149,N_39606,N_37113);
xor U42150 (N_42150,N_33544,N_39522);
xnor U42151 (N_42151,N_33324,N_34699);
or U42152 (N_42152,N_35174,N_38285);
and U42153 (N_42153,N_38035,N_30866);
and U42154 (N_42154,N_35995,N_32428);
xnor U42155 (N_42155,N_33729,N_38016);
xor U42156 (N_42156,N_31473,N_31499);
nand U42157 (N_42157,N_36576,N_37103);
nor U42158 (N_42158,N_35083,N_31645);
and U42159 (N_42159,N_37277,N_38618);
nor U42160 (N_42160,N_35054,N_31601);
and U42161 (N_42161,N_34277,N_36993);
and U42162 (N_42162,N_33839,N_39137);
and U42163 (N_42163,N_39366,N_30409);
xnor U42164 (N_42164,N_31349,N_38233);
nand U42165 (N_42165,N_39877,N_32662);
nor U42166 (N_42166,N_38702,N_36612);
nand U42167 (N_42167,N_38564,N_31694);
or U42168 (N_42168,N_36061,N_36169);
nor U42169 (N_42169,N_31860,N_32573);
xor U42170 (N_42170,N_32806,N_36499);
nand U42171 (N_42171,N_35941,N_36829);
or U42172 (N_42172,N_31336,N_39160);
and U42173 (N_42173,N_38954,N_36384);
nand U42174 (N_42174,N_39230,N_37631);
xnor U42175 (N_42175,N_33290,N_33160);
or U42176 (N_42176,N_33477,N_36705);
and U42177 (N_42177,N_32376,N_33308);
and U42178 (N_42178,N_34793,N_38066);
xnor U42179 (N_42179,N_32089,N_39125);
nor U42180 (N_42180,N_32165,N_31410);
xor U42181 (N_42181,N_35242,N_39971);
nor U42182 (N_42182,N_38745,N_34186);
xnor U42183 (N_42183,N_37641,N_31063);
and U42184 (N_42184,N_37545,N_38806);
nand U42185 (N_42185,N_37186,N_34158);
xnor U42186 (N_42186,N_32364,N_34188);
nor U42187 (N_42187,N_32879,N_33806);
xnor U42188 (N_42188,N_35841,N_35022);
xnor U42189 (N_42189,N_37060,N_35610);
nor U42190 (N_42190,N_35241,N_33099);
xor U42191 (N_42191,N_37163,N_37327);
and U42192 (N_42192,N_38256,N_39020);
nor U42193 (N_42193,N_32997,N_36247);
and U42194 (N_42194,N_37136,N_33616);
nand U42195 (N_42195,N_38138,N_34006);
nand U42196 (N_42196,N_37358,N_36988);
and U42197 (N_42197,N_31840,N_38689);
xor U42198 (N_42198,N_34564,N_32342);
or U42199 (N_42199,N_35895,N_36939);
xor U42200 (N_42200,N_35281,N_37455);
xor U42201 (N_42201,N_30066,N_31886);
nor U42202 (N_42202,N_30956,N_31332);
xnor U42203 (N_42203,N_35424,N_31628);
xnor U42204 (N_42204,N_32814,N_32829);
and U42205 (N_42205,N_32676,N_38572);
and U42206 (N_42206,N_33564,N_37777);
nor U42207 (N_42207,N_30688,N_36958);
or U42208 (N_42208,N_36650,N_30880);
and U42209 (N_42209,N_36641,N_39247);
nand U42210 (N_42210,N_37798,N_31794);
and U42211 (N_42211,N_30257,N_32063);
nor U42212 (N_42212,N_36452,N_38966);
and U42213 (N_42213,N_36069,N_38551);
or U42214 (N_42214,N_31818,N_39844);
nand U42215 (N_42215,N_39026,N_32119);
and U42216 (N_42216,N_33458,N_34063);
nor U42217 (N_42217,N_37698,N_32481);
or U42218 (N_42218,N_37552,N_32777);
xnor U42219 (N_42219,N_37400,N_35550);
nand U42220 (N_42220,N_36035,N_32780);
and U42221 (N_42221,N_31634,N_31201);
xor U42222 (N_42222,N_35253,N_38349);
nor U42223 (N_42223,N_37630,N_34622);
nand U42224 (N_42224,N_33924,N_34005);
nand U42225 (N_42225,N_36756,N_36041);
and U42226 (N_42226,N_33793,N_38504);
or U42227 (N_42227,N_35255,N_38850);
nand U42228 (N_42228,N_35858,N_38464);
xnor U42229 (N_42229,N_32066,N_30054);
or U42230 (N_42230,N_38730,N_38180);
nor U42231 (N_42231,N_39311,N_37623);
nand U42232 (N_42232,N_36017,N_32135);
nand U42233 (N_42233,N_38155,N_37441);
nor U42234 (N_42234,N_39348,N_39547);
or U42235 (N_42235,N_30140,N_37686);
and U42236 (N_42236,N_34708,N_31253);
or U42237 (N_42237,N_31182,N_35882);
or U42238 (N_42238,N_34738,N_35528);
xnor U42239 (N_42239,N_39340,N_36416);
xor U42240 (N_42240,N_35903,N_33397);
and U42241 (N_42241,N_39577,N_32218);
xor U42242 (N_42242,N_30899,N_36174);
nor U42243 (N_42243,N_34317,N_35773);
xor U42244 (N_42244,N_31740,N_36162);
or U42245 (N_42245,N_35301,N_35797);
or U42246 (N_42246,N_32327,N_37491);
nor U42247 (N_42247,N_31236,N_35395);
or U42248 (N_42248,N_35012,N_38011);
or U42249 (N_42249,N_35595,N_38543);
nor U42250 (N_42250,N_35533,N_30544);
nor U42251 (N_42251,N_39599,N_38054);
xor U42252 (N_42252,N_34059,N_31661);
nor U42253 (N_42253,N_39029,N_38922);
nand U42254 (N_42254,N_31727,N_35363);
and U42255 (N_42255,N_37560,N_30901);
or U42256 (N_42256,N_34214,N_32897);
nand U42257 (N_42257,N_33893,N_35403);
nand U42258 (N_42258,N_33671,N_35389);
xor U42259 (N_42259,N_30972,N_37643);
and U42260 (N_42260,N_33045,N_38391);
or U42261 (N_42261,N_37951,N_33877);
or U42262 (N_42262,N_32627,N_30028);
and U42263 (N_42263,N_38164,N_33376);
or U42264 (N_42264,N_36154,N_33211);
xor U42265 (N_42265,N_36938,N_34339);
nor U42266 (N_42266,N_30855,N_37050);
nand U42267 (N_42267,N_33682,N_30149);
or U42268 (N_42268,N_39866,N_32977);
and U42269 (N_42269,N_34795,N_36068);
and U42270 (N_42270,N_32889,N_39525);
or U42271 (N_42271,N_37140,N_37958);
or U42272 (N_42272,N_33875,N_32616);
xor U42273 (N_42273,N_35469,N_34705);
and U42274 (N_42274,N_31161,N_30878);
xnor U42275 (N_42275,N_39666,N_38313);
and U42276 (N_42276,N_37807,N_34607);
nand U42277 (N_42277,N_30207,N_33335);
or U42278 (N_42278,N_35374,N_34347);
or U42279 (N_42279,N_32722,N_32378);
nand U42280 (N_42280,N_38653,N_38582);
xor U42281 (N_42281,N_37601,N_35876);
and U42282 (N_42282,N_31167,N_39463);
and U42283 (N_42283,N_34331,N_31285);
or U42284 (N_42284,N_30663,N_36786);
nand U42285 (N_42285,N_30507,N_35951);
xnor U42286 (N_42286,N_36711,N_31373);
or U42287 (N_42287,N_37372,N_31782);
or U42288 (N_42288,N_34069,N_33694);
and U42289 (N_42289,N_33381,N_34647);
nand U42290 (N_42290,N_37305,N_33639);
or U42291 (N_42291,N_31548,N_38205);
nor U42292 (N_42292,N_35998,N_30122);
or U42293 (N_42293,N_33866,N_38926);
nor U42294 (N_42294,N_39097,N_33582);
and U42295 (N_42295,N_35375,N_36327);
and U42296 (N_42296,N_33907,N_34373);
and U42297 (N_42297,N_34909,N_39627);
or U42298 (N_42298,N_31528,N_38608);
and U42299 (N_42299,N_30573,N_30173);
nand U42300 (N_42300,N_39262,N_39122);
xnor U42301 (N_42301,N_37699,N_31760);
nor U42302 (N_42302,N_39093,N_39578);
xor U42303 (N_42303,N_31791,N_37057);
xor U42304 (N_42304,N_38649,N_36295);
nor U42305 (N_42305,N_31428,N_34136);
nand U42306 (N_42306,N_38249,N_32182);
xnor U42307 (N_42307,N_36183,N_32191);
nand U42308 (N_42308,N_36149,N_35269);
and U42309 (N_42309,N_30787,N_35991);
nor U42310 (N_42310,N_37820,N_35848);
and U42311 (N_42311,N_33717,N_31865);
and U42312 (N_42312,N_34175,N_30458);
nor U42313 (N_42313,N_35932,N_34876);
and U42314 (N_42314,N_34859,N_38502);
nand U42315 (N_42315,N_32308,N_39513);
nand U42316 (N_42316,N_31235,N_37691);
and U42317 (N_42317,N_36434,N_35172);
or U42318 (N_42318,N_32072,N_39501);
nand U42319 (N_42319,N_36548,N_30239);
and U42320 (N_42320,N_36473,N_33467);
nand U42321 (N_42321,N_38901,N_35529);
or U42322 (N_42322,N_38927,N_38028);
xnor U42323 (N_42323,N_38265,N_36968);
nand U42324 (N_42324,N_38338,N_30557);
and U42325 (N_42325,N_34418,N_37213);
or U42326 (N_42326,N_38135,N_32598);
nor U42327 (N_42327,N_33405,N_35897);
xor U42328 (N_42328,N_33169,N_32444);
xor U42329 (N_42329,N_34619,N_35952);
nor U42330 (N_42330,N_30319,N_31412);
nor U42331 (N_42331,N_33634,N_39267);
xor U42332 (N_42332,N_38088,N_32988);
nor U42333 (N_42333,N_30993,N_33221);
nor U42334 (N_42334,N_32110,N_34090);
nand U42335 (N_42335,N_31030,N_37626);
nand U42336 (N_42336,N_30872,N_35846);
and U42337 (N_42337,N_30146,N_32590);
and U42338 (N_42338,N_30718,N_31495);
or U42339 (N_42339,N_34397,N_30755);
xnor U42340 (N_42340,N_37346,N_38519);
nand U42341 (N_42341,N_38835,N_32817);
and U42342 (N_42342,N_38533,N_31909);
and U42343 (N_42343,N_36146,N_37088);
xor U42344 (N_42344,N_32434,N_33974);
or U42345 (N_42345,N_33735,N_35702);
xnor U42346 (N_42346,N_32804,N_36242);
and U42347 (N_42347,N_36996,N_38206);
and U42348 (N_42348,N_39072,N_33020);
nand U42349 (N_42349,N_36372,N_34061);
or U42350 (N_42350,N_35707,N_34836);
nor U42351 (N_42351,N_33612,N_32085);
nor U42352 (N_42352,N_30885,N_34156);
nor U42353 (N_42353,N_37335,N_32248);
xor U42354 (N_42354,N_33092,N_30230);
xnor U42355 (N_42355,N_35973,N_38924);
xnor U42356 (N_42356,N_36953,N_38694);
xnor U42357 (N_42357,N_33377,N_38804);
or U42358 (N_42358,N_36783,N_39703);
and U42359 (N_42359,N_37858,N_36138);
nor U42360 (N_42360,N_35019,N_37743);
xnor U42361 (N_42361,N_30364,N_32657);
xnor U42362 (N_42362,N_35146,N_36200);
nand U42363 (N_42363,N_33576,N_31348);
and U42364 (N_42364,N_38357,N_37308);
xor U42365 (N_42365,N_35756,N_33481);
or U42366 (N_42366,N_30670,N_35887);
or U42367 (N_42367,N_36632,N_31118);
nor U42368 (N_42368,N_30217,N_35470);
and U42369 (N_42369,N_32872,N_39714);
xor U42370 (N_42370,N_37868,N_32057);
xnor U42371 (N_42371,N_35568,N_32413);
and U42372 (N_42372,N_35647,N_38084);
nor U42373 (N_42373,N_30462,N_30106);
xor U42374 (N_42374,N_35819,N_32869);
xnor U42375 (N_42375,N_37632,N_36582);
nand U42376 (N_42376,N_33434,N_31825);
nand U42377 (N_42377,N_36106,N_36505);
and U42378 (N_42378,N_32026,N_34237);
nor U42379 (N_42379,N_38456,N_30629);
or U42380 (N_42380,N_35945,N_36225);
nand U42381 (N_42381,N_37008,N_39349);
or U42382 (N_42382,N_36458,N_36843);
xnor U42383 (N_42383,N_38487,N_33994);
or U42384 (N_42384,N_31210,N_30701);
and U42385 (N_42385,N_33755,N_33217);
or U42386 (N_42386,N_39717,N_32211);
nor U42387 (N_42387,N_33751,N_30776);
nor U42388 (N_42388,N_30759,N_36771);
or U42389 (N_42389,N_30800,N_37120);
xor U42390 (N_42390,N_37292,N_34140);
and U42391 (N_42391,N_31888,N_34355);
nand U42392 (N_42392,N_32294,N_38698);
and U42393 (N_42393,N_39813,N_33339);
nor U42394 (N_42394,N_36382,N_31813);
xnor U42395 (N_42395,N_37282,N_30607);
and U42396 (N_42396,N_36892,N_39164);
or U42397 (N_42397,N_34575,N_36902);
and U42398 (N_42398,N_30175,N_34130);
nor U42399 (N_42399,N_37175,N_31485);
and U42400 (N_42400,N_30382,N_31657);
and U42401 (N_42401,N_30174,N_33879);
nand U42402 (N_42402,N_38545,N_33472);
xor U42403 (N_42403,N_33867,N_34072);
and U42404 (N_42404,N_37350,N_36990);
nor U42405 (N_42405,N_30798,N_32932);
or U42406 (N_42406,N_39648,N_37812);
xor U42407 (N_42407,N_38179,N_34872);
xnor U42408 (N_42408,N_37150,N_32169);
xnor U42409 (N_42409,N_33577,N_36103);
or U42410 (N_42410,N_32464,N_30843);
or U42411 (N_42411,N_39790,N_30702);
xor U42412 (N_42412,N_32477,N_34251);
nand U42413 (N_42413,N_38690,N_38052);
or U42414 (N_42414,N_33669,N_36948);
or U42415 (N_42415,N_39861,N_37107);
xor U42416 (N_42416,N_39363,N_34501);
or U42417 (N_42417,N_35003,N_33260);
xor U42418 (N_42418,N_32267,N_30064);
nand U42419 (N_42419,N_38148,N_37943);
xor U42420 (N_42420,N_39111,N_30577);
xnor U42421 (N_42421,N_34187,N_33934);
or U42422 (N_42422,N_35069,N_39953);
nand U42423 (N_42423,N_30783,N_32571);
or U42424 (N_42424,N_33719,N_35310);
nand U42425 (N_42425,N_38141,N_37429);
xnor U42426 (N_42426,N_34541,N_31116);
xnor U42427 (N_42427,N_39604,N_33031);
xnor U42428 (N_42428,N_37666,N_35961);
nor U42429 (N_42429,N_39672,N_31717);
nor U42430 (N_42430,N_37759,N_38764);
and U42431 (N_42431,N_37047,N_36114);
nand U42432 (N_42432,N_32253,N_35486);
nand U42433 (N_42433,N_35076,N_33225);
xor U42434 (N_42434,N_39064,N_34163);
or U42435 (N_42435,N_38103,N_37827);
and U42436 (N_42436,N_32942,N_30133);
or U42437 (N_42437,N_35011,N_33374);
nand U42438 (N_42438,N_39339,N_34777);
nand U42439 (N_42439,N_37749,N_31350);
and U42440 (N_42440,N_36529,N_38580);
xnor U42441 (N_42441,N_30115,N_34989);
and U42442 (N_42442,N_31442,N_36877);
and U42443 (N_42443,N_31112,N_31525);
xor U42444 (N_42444,N_37325,N_35868);
or U42445 (N_42445,N_39980,N_38509);
or U42446 (N_42446,N_39034,N_39053);
nand U42447 (N_42447,N_33156,N_35631);
and U42448 (N_42448,N_37373,N_37968);
or U42449 (N_42449,N_38938,N_35860);
or U42450 (N_42450,N_32426,N_36078);
nor U42451 (N_42451,N_33731,N_33549);
nor U42452 (N_42452,N_33683,N_37146);
nand U42453 (N_42453,N_35214,N_36052);
nand U42454 (N_42454,N_37764,N_32019);
nor U42455 (N_42455,N_35591,N_30031);
and U42456 (N_42456,N_37378,N_33575);
or U42457 (N_42457,N_36725,N_36354);
nand U42458 (N_42458,N_38121,N_31152);
and U42459 (N_42459,N_38881,N_30893);
and U42460 (N_42460,N_30795,N_35116);
nand U42461 (N_42461,N_39353,N_35981);
nor U42462 (N_42462,N_38448,N_39227);
xor U42463 (N_42463,N_38596,N_31482);
nor U42464 (N_42464,N_38350,N_36508);
nor U42465 (N_42465,N_34686,N_35979);
nand U42466 (N_42466,N_35799,N_36687);
and U42467 (N_42467,N_36014,N_32265);
or U42468 (N_42468,N_37125,N_31487);
and U42469 (N_42469,N_33328,N_37819);
xnor U42470 (N_42470,N_30280,N_33900);
nand U42471 (N_42471,N_30452,N_36680);
xnor U42472 (N_42472,N_33977,N_37415);
or U42473 (N_42473,N_32230,N_33241);
nor U42474 (N_42474,N_36755,N_39233);
nand U42475 (N_42475,N_38847,N_39212);
nand U42476 (N_42476,N_37912,N_36445);
and U42477 (N_42477,N_30523,N_32417);
and U42478 (N_42478,N_32332,N_39504);
xor U42479 (N_42479,N_32186,N_35154);
nand U42480 (N_42480,N_31744,N_36341);
or U42481 (N_42481,N_39998,N_36487);
nand U42482 (N_42482,N_30005,N_32331);
nand U42483 (N_42483,N_30510,N_35883);
nand U42484 (N_42484,N_34926,N_38503);
and U42485 (N_42485,N_35093,N_35583);
nand U42486 (N_42486,N_35259,N_34067);
and U42487 (N_42487,N_33273,N_38718);
nand U42488 (N_42488,N_36955,N_35970);
xnor U42489 (N_42489,N_33984,N_33763);
xnor U42490 (N_42490,N_38160,N_38364);
nand U42491 (N_42491,N_30867,N_34902);
nor U42492 (N_42492,N_39908,N_32810);
nand U42493 (N_42493,N_38904,N_39032);
nand U42494 (N_42494,N_31932,N_32076);
or U42495 (N_42495,N_36793,N_31371);
and U42496 (N_42496,N_39922,N_34624);
or U42497 (N_42497,N_30713,N_37066);
nor U42498 (N_42498,N_36412,N_36123);
and U42499 (N_42499,N_31057,N_34886);
and U42500 (N_42500,N_37293,N_39406);
nand U42501 (N_42501,N_31084,N_30974);
xor U42502 (N_42502,N_36104,N_32282);
or U42503 (N_42503,N_36066,N_35878);
and U42504 (N_42504,N_37882,N_31580);
and U42505 (N_42505,N_38436,N_35489);
or U42506 (N_42506,N_33908,N_35001);
nand U42507 (N_42507,N_33453,N_38792);
nand U42508 (N_42508,N_30063,N_30299);
xor U42509 (N_42509,N_37252,N_31721);
xnor U42510 (N_42510,N_32093,N_37159);
nand U42511 (N_42511,N_32575,N_34423);
and U42512 (N_42512,N_32784,N_37479);
nand U42513 (N_42513,N_30178,N_39056);
xnor U42514 (N_42514,N_37716,N_39999);
xor U42515 (N_42515,N_36287,N_35141);
and U42516 (N_42516,N_35956,N_37610);
and U42517 (N_42517,N_33996,N_30102);
xor U42518 (N_42518,N_33880,N_36542);
nor U42519 (N_42519,N_32320,N_32273);
nor U42520 (N_42520,N_39140,N_32857);
or U42521 (N_42521,N_38181,N_35450);
xor U42522 (N_42522,N_39084,N_36929);
or U42523 (N_42523,N_35427,N_31730);
and U42524 (N_42524,N_39704,N_32268);
nor U42525 (N_42525,N_31969,N_31612);
nor U42526 (N_42526,N_38531,N_30121);
nor U42527 (N_42527,N_31882,N_30662);
nand U42528 (N_42528,N_30025,N_32440);
xor U42529 (N_42529,N_30858,N_33628);
xor U42530 (N_42530,N_35075,N_38336);
and U42531 (N_42531,N_30914,N_38221);
or U42532 (N_42532,N_33692,N_33016);
nor U42533 (N_42533,N_35064,N_33819);
or U42534 (N_42534,N_32643,N_36307);
nor U42535 (N_42535,N_32527,N_34711);
nand U42536 (N_42536,N_30506,N_30647);
and U42537 (N_42537,N_32775,N_32765);
xnor U42538 (N_42538,N_39995,N_32915);
nor U42539 (N_42539,N_36909,N_34296);
or U42540 (N_42540,N_36045,N_37571);
and U42541 (N_42541,N_30467,N_31465);
nor U42542 (N_42542,N_37418,N_33865);
or U42543 (N_42543,N_30512,N_38193);
nor U42544 (N_42544,N_36385,N_30162);
nor U42545 (N_42545,N_37408,N_39088);
and U42546 (N_42546,N_39874,N_34194);
nor U42547 (N_42547,N_30703,N_35417);
xnor U42548 (N_42548,N_38310,N_36752);
nor U42549 (N_42549,N_30434,N_30165);
xor U42550 (N_42550,N_38061,N_36647);
nand U42551 (N_42551,N_34701,N_32338);
and U42552 (N_42552,N_37317,N_35451);
nand U42553 (N_42553,N_34318,N_31046);
nor U42554 (N_42554,N_30970,N_30730);
and U42555 (N_42555,N_31358,N_30252);
and U42556 (N_42556,N_37852,N_31846);
nand U42557 (N_42557,N_39835,N_30422);
and U42558 (N_42558,N_38811,N_38515);
xnor U42559 (N_42559,N_38418,N_37342);
xor U42560 (N_42560,N_33805,N_38322);
nand U42561 (N_42561,N_33239,N_33054);
nor U42562 (N_42562,N_31728,N_39259);
nand U42563 (N_42563,N_36038,N_32985);
nor U42564 (N_42564,N_35667,N_39149);
or U42565 (N_42565,N_32545,N_39920);
and U42566 (N_42566,N_33469,N_36986);
xnor U42567 (N_42567,N_32353,N_39187);
or U42568 (N_42568,N_30051,N_39848);
or U42569 (N_42569,N_37620,N_38110);
nor U42570 (N_42570,N_30897,N_38527);
xor U42571 (N_42571,N_37974,N_32292);
and U42572 (N_42572,N_30576,N_36298);
and U42573 (N_42573,N_30944,N_30781);
xor U42574 (N_42574,N_38785,N_30346);
xor U42575 (N_42575,N_30201,N_35534);
nor U42576 (N_42576,N_33111,N_39322);
xnor U42577 (N_42577,N_31333,N_31463);
nor U42578 (N_42578,N_35444,N_32694);
nand U42579 (N_42579,N_32893,N_37391);
xor U42580 (N_42580,N_32179,N_39601);
nand U42581 (N_42581,N_39815,N_35891);
and U42582 (N_42582,N_39686,N_32432);
nand U42583 (N_42583,N_37709,N_33923);
nand U42584 (N_42584,N_30055,N_37897);
xnor U42585 (N_42585,N_32702,N_31712);
xnor U42586 (N_42586,N_37808,N_39376);
xnor U42587 (N_42587,N_35530,N_39763);
and U42588 (N_42588,N_33891,N_31869);
or U42589 (N_42589,N_39228,N_33551);
xor U42590 (N_42590,N_35182,N_35958);
xor U42591 (N_42591,N_36229,N_38606);
and U42592 (N_42592,N_34725,N_32075);
xnor U42593 (N_42593,N_34787,N_37799);
nand U42594 (N_42594,N_35068,N_37493);
xor U42595 (N_42595,N_32589,N_35445);
xor U42596 (N_42596,N_31618,N_38423);
nand U42597 (N_42597,N_34585,N_36825);
and U42598 (N_42598,N_34295,N_37890);
nand U42599 (N_42599,N_32263,N_36465);
and U42600 (N_42600,N_35565,N_30218);
and U42601 (N_42601,N_38329,N_38461);
or U42602 (N_42602,N_30492,N_31010);
nor U42603 (N_42603,N_31833,N_37402);
and U42604 (N_42604,N_33292,N_32134);
xor U42605 (N_42605,N_33573,N_32681);
or U42606 (N_42606,N_32341,N_36492);
xor U42607 (N_42607,N_37339,N_36724);
nand U42608 (N_42608,N_39840,N_38921);
and U42609 (N_42609,N_33884,N_38326);
nand U42610 (N_42610,N_35438,N_35415);
or U42611 (N_42611,N_30314,N_36024);
nor U42612 (N_42612,N_33528,N_31832);
nand U42613 (N_42613,N_31363,N_36689);
nand U42614 (N_42614,N_34562,N_33384);
nor U42615 (N_42615,N_31206,N_33259);
nor U42616 (N_42616,N_30302,N_37333);
nand U42617 (N_42617,N_34929,N_34539);
nor U42618 (N_42618,N_38869,N_33557);
or U42619 (N_42619,N_31038,N_36933);
and U42620 (N_42620,N_36020,N_30594);
or U42621 (N_42621,N_34443,N_34531);
xnor U42622 (N_42622,N_30527,N_34767);
or U42623 (N_42623,N_36349,N_39560);
nand U42624 (N_42624,N_35167,N_33942);
and U42625 (N_42625,N_33459,N_38783);
nand U42626 (N_42626,N_35781,N_38132);
xnor U42627 (N_42627,N_33209,N_30998);
nor U42628 (N_42628,N_35576,N_30614);
xor U42629 (N_42629,N_35902,N_30305);
and U42630 (N_42630,N_36406,N_32473);
or U42631 (N_42631,N_37454,N_35080);
or U42632 (N_42632,N_30562,N_33394);
and U42633 (N_42633,N_35632,N_30518);
xnor U42634 (N_42634,N_37711,N_34652);
xor U42635 (N_42635,N_38707,N_34648);
nor U42636 (N_42636,N_37998,N_35239);
nand U42637 (N_42637,N_32436,N_30143);
nand U42638 (N_42638,N_36305,N_39057);
or U42639 (N_42639,N_31738,N_32994);
nand U42640 (N_42640,N_39481,N_32213);
or U42641 (N_42641,N_30499,N_35177);
nand U42642 (N_42642,N_34183,N_31418);
nor U42643 (N_42643,N_31700,N_32531);
xor U42644 (N_42644,N_38014,N_36449);
or U42645 (N_42645,N_34559,N_33663);
xnor U42646 (N_42646,N_34829,N_38728);
nor U42647 (N_42647,N_32249,N_34546);
nand U42648 (N_42648,N_34561,N_31641);
and U42649 (N_42649,N_30470,N_35112);
nand U42650 (N_42650,N_35788,N_37485);
or U42651 (N_42651,N_38574,N_31006);
xor U42652 (N_42652,N_39242,N_31322);
nand U42653 (N_42653,N_38899,N_35482);
nor U42654 (N_42654,N_30748,N_30053);
nor U42655 (N_42655,N_32515,N_37872);
nor U42656 (N_42656,N_30882,N_36413);
xor U42657 (N_42657,N_37147,N_33025);
or U42658 (N_42658,N_33976,N_30520);
nor U42659 (N_42659,N_37997,N_31637);
nor U42660 (N_42660,N_30889,N_35866);
or U42661 (N_42661,N_36951,N_38800);
xnor U42662 (N_42662,N_38368,N_38378);
or U42663 (N_42663,N_36784,N_39680);
and U42664 (N_42664,N_33525,N_32781);
xnor U42665 (N_42665,N_31988,N_35248);
and U42666 (N_42666,N_35523,N_35552);
nor U42667 (N_42667,N_31239,N_32459);
xnor U42668 (N_42668,N_34760,N_39478);
nor U42669 (N_42669,N_39408,N_38704);
and U42670 (N_42670,N_37700,N_31054);
xnor U42671 (N_42671,N_32449,N_33010);
nand U42672 (N_42672,N_35368,N_32003);
xnor U42673 (N_42673,N_35686,N_32420);
and U42674 (N_42674,N_35851,N_39726);
or U42675 (N_42675,N_33372,N_38279);
and U42676 (N_42676,N_34492,N_32325);
xnor U42677 (N_42677,N_35078,N_35127);
nand U42678 (N_42678,N_38571,N_31767);
or U42679 (N_42679,N_35601,N_39718);
nand U42680 (N_42680,N_39510,N_36919);
nand U42681 (N_42681,N_36622,N_37488);
and U42682 (N_42682,N_39989,N_30736);
or U42683 (N_42683,N_37457,N_31486);
nand U42684 (N_42684,N_32570,N_37464);
xnor U42685 (N_42685,N_38363,N_32397);
nand U42686 (N_42686,N_33876,N_30930);
or U42687 (N_42687,N_36945,N_36739);
and U42688 (N_42688,N_37162,N_33120);
or U42689 (N_42689,N_39263,N_30986);
nor U42690 (N_42690,N_30953,N_31050);
and U42691 (N_42691,N_34862,N_36422);
nand U42692 (N_42692,N_33592,N_34093);
xor U42693 (N_42693,N_38777,N_31244);
xor U42694 (N_42694,N_35109,N_39661);
nor U42695 (N_42695,N_34039,N_31507);
xnor U42696 (N_42696,N_37581,N_30685);
xor U42697 (N_42697,N_31837,N_38917);
nor U42698 (N_42698,N_32552,N_34106);
nor U42699 (N_42699,N_33611,N_31736);
xor U42700 (N_42700,N_38073,N_30491);
nor U42701 (N_42701,N_35401,N_39655);
or U42702 (N_42702,N_36302,N_34519);
and U42703 (N_42703,N_33280,N_36209);
and U42704 (N_42704,N_39213,N_35971);
nor U42705 (N_42705,N_32080,N_35160);
nor U42706 (N_42706,N_38967,N_33985);
or U42707 (N_42707,N_36491,N_34956);
or U42708 (N_42708,N_32516,N_30315);
and U42709 (N_42709,N_34020,N_32504);
xnor U42710 (N_42710,N_32949,N_32883);
or U42711 (N_42711,N_38544,N_35821);
and U42712 (N_42712,N_34057,N_39288);
and U42713 (N_42713,N_31409,N_33425);
xnor U42714 (N_42714,N_36710,N_31776);
nor U42715 (N_42715,N_34891,N_38817);
nor U42716 (N_42716,N_36889,N_30831);
or U42717 (N_42717,N_33559,N_34536);
nor U42718 (N_42718,N_32867,N_36090);
or U42719 (N_42719,N_35202,N_34814);
nor U42720 (N_42720,N_37962,N_34123);
nor U42721 (N_42721,N_32801,N_36543);
nand U42722 (N_42722,N_31088,N_34382);
nor U42723 (N_42723,N_39462,N_30955);
or U42724 (N_42724,N_30833,N_33018);
xor U42725 (N_42725,N_33263,N_30040);
and U42726 (N_42726,N_33918,N_31624);
and U42727 (N_42727,N_33700,N_30135);
or U42728 (N_42728,N_37961,N_38670);
nand U42729 (N_42729,N_30812,N_38102);
nand U42730 (N_42730,N_38006,N_35922);
xor U42731 (N_42731,N_31775,N_30618);
nor U42732 (N_42732,N_35452,N_30917);
xnor U42733 (N_42733,N_33122,N_34265);
nand U42734 (N_42734,N_39070,N_34243);
nor U42735 (N_42735,N_34048,N_37475);
nor U42736 (N_42736,N_35158,N_33571);
or U42737 (N_42737,N_38104,N_30361);
xnor U42738 (N_42738,N_30821,N_39083);
nor U42739 (N_42739,N_34215,N_33730);
or U42740 (N_42740,N_39455,N_31319);
and U42741 (N_42741,N_34826,N_33898);
nand U42742 (N_42742,N_31520,N_39954);
xor U42743 (N_42743,N_34053,N_34306);
and U42744 (N_42744,N_35437,N_36884);
nor U42745 (N_42745,N_32842,N_31138);
nand U42746 (N_42746,N_38746,N_33000);
and U42747 (N_42747,N_36498,N_30521);
and U42748 (N_42748,N_33563,N_37715);
xnor U42749 (N_42749,N_35205,N_35830);
xnor U42750 (N_42750,N_30679,N_35371);
xnor U42751 (N_42751,N_31179,N_37173);
and U42752 (N_42752,N_36893,N_36015);
nand U42753 (N_42753,N_35646,N_30298);
xnor U42754 (N_42754,N_34218,N_34261);
nand U42755 (N_42755,N_34342,N_39006);
and U42756 (N_42756,N_30971,N_35498);
xor U42757 (N_42757,N_38613,N_35008);
nand U42758 (N_42758,N_32183,N_30377);
and U42759 (N_42759,N_39852,N_37598);
xor U42760 (N_42760,N_32581,N_39503);
xor U42761 (N_42761,N_31353,N_34644);
and U42762 (N_42762,N_34599,N_32821);
nand U42763 (N_42763,N_35889,N_34820);
nand U42764 (N_42764,N_33314,N_36512);
xnor U42765 (N_42765,N_39962,N_36044);
and U42766 (N_42766,N_38648,N_39917);
and U42767 (N_42767,N_30410,N_38762);
nor U42768 (N_42768,N_30934,N_32022);
and U42769 (N_42769,N_30128,N_36743);
or U42770 (N_42770,N_37016,N_35461);
nand U42771 (N_42771,N_37569,N_35626);
or U42772 (N_42772,N_35265,N_34632);
and U42773 (N_42773,N_39895,N_31534);
or U42774 (N_42774,N_37640,N_32062);
nor U42775 (N_42775,N_36155,N_39359);
nand U42776 (N_42776,N_32077,N_39597);
xnor U42777 (N_42777,N_35798,N_39899);
xor U42778 (N_42778,N_37007,N_32120);
and U42779 (N_42779,N_30126,N_33420);
and U42780 (N_42780,N_32572,N_37482);
nor U42781 (N_42781,N_37246,N_39156);
or U42782 (N_42782,N_39365,N_31778);
or U42783 (N_42783,N_38866,N_33320);
xnor U42784 (N_42784,N_31892,N_38294);
nand U42785 (N_42785,N_35695,N_38944);
nor U42786 (N_42786,N_38005,N_34333);
and U42787 (N_42787,N_30699,N_36125);
and U42788 (N_42788,N_36319,N_34527);
or U42789 (N_42789,N_35289,N_33283);
xor U42790 (N_42790,N_34219,N_32281);
xnor U42791 (N_42791,N_38821,N_36457);
nand U42792 (N_42792,N_36523,N_38370);
nor U42793 (N_42793,N_34376,N_36879);
nand U42794 (N_42794,N_30501,N_36373);
xnor U42795 (N_42795,N_35088,N_33138);
or U42796 (N_42796,N_34679,N_38556);
and U42797 (N_42797,N_31340,N_36072);
nand U42798 (N_42798,N_32986,N_32472);
or U42799 (N_42799,N_38208,N_34035);
and U42800 (N_42800,N_38765,N_30999);
or U42801 (N_42801,N_37288,N_31041);
and U42802 (N_42802,N_37725,N_32187);
or U42803 (N_42803,N_32202,N_38444);
or U42804 (N_42804,N_38442,N_38161);
or U42805 (N_42805,N_31904,N_32687);
xor U42806 (N_42806,N_31800,N_35539);
xnor U42807 (N_42807,N_31671,N_33356);
or U42808 (N_42808,N_33198,N_33670);
xor U42809 (N_42809,N_35964,N_37486);
xnor U42810 (N_42810,N_39009,N_38637);
and U42811 (N_42811,N_36642,N_36220);
nand U42812 (N_42812,N_34267,N_32227);
nor U42813 (N_42813,N_39082,N_33297);
xor U42814 (N_42814,N_33604,N_31174);
nand U42815 (N_42815,N_32025,N_37166);
nand U42816 (N_42816,N_31658,N_34366);
xnor U42817 (N_42817,N_35976,N_36947);
or U42818 (N_42818,N_38361,N_33945);
xor U42819 (N_42819,N_35705,N_39964);
and U42820 (N_42820,N_37568,N_38463);
and U42821 (N_42821,N_37337,N_39113);
xor U42822 (N_42822,N_36975,N_33243);
nor U42823 (N_42823,N_37965,N_35066);
nand U42824 (N_42824,N_39297,N_38153);
and U42825 (N_42825,N_38834,N_35641);
nand U42826 (N_42826,N_39283,N_37745);
and U42827 (N_42827,N_36399,N_31361);
nand U42828 (N_42828,N_32465,N_36965);
nor U42829 (N_42829,N_31429,N_31374);
nand U42830 (N_42830,N_39900,N_32730);
and U42831 (N_42831,N_39723,N_31077);
xnor U42832 (N_42832,N_31220,N_30549);
nor U42833 (N_42833,N_37445,N_31021);
xnor U42834 (N_42834,N_33704,N_34957);
and U42835 (N_42835,N_33725,N_31123);
nand U42836 (N_42836,N_33375,N_35541);
nor U42837 (N_42837,N_31025,N_31466);
nand U42838 (N_42838,N_30141,N_34015);
nor U42839 (N_42839,N_31086,N_32196);
and U42840 (N_42840,N_37049,N_30192);
xnor U42841 (N_42841,N_37972,N_31986);
xor U42842 (N_42842,N_38373,N_34910);
nor U42843 (N_42843,N_39705,N_31470);
nand U42844 (N_42844,N_39067,N_34529);
nor U42845 (N_42845,N_37128,N_30660);
nand U42846 (N_42846,N_35778,N_38041);
nand U42847 (N_42847,N_37129,N_34693);
nand U42848 (N_42848,N_30486,N_38346);
and U42849 (N_42849,N_31962,N_31289);
or U42850 (N_42850,N_36455,N_37727);
nand U42851 (N_42851,N_36163,N_32207);
and U42852 (N_42852,N_32618,N_34088);
and U42853 (N_42853,N_39782,N_30033);
nor U42854 (N_42854,N_33011,N_34831);
or U42855 (N_42855,N_35221,N_35966);
nor U42856 (N_42856,N_39976,N_39435);
nand U42857 (N_42857,N_37680,N_37164);
xor U42858 (N_42858,N_39250,N_34029);
and U42859 (N_42859,N_34565,N_31608);
nor U42860 (N_42860,N_36496,N_34164);
xor U42861 (N_42861,N_38775,N_35414);
and U42862 (N_42862,N_35319,N_35706);
or U42863 (N_42863,N_31599,N_36190);
or U42864 (N_42864,N_31803,N_37151);
and U42865 (N_42865,N_36661,N_35535);
nor U42866 (N_42866,N_32351,N_33103);
and U42867 (N_42867,N_39494,N_38055);
or U42868 (N_42868,N_34803,N_30229);
nor U42869 (N_42869,N_37733,N_36201);
or U42870 (N_42870,N_37862,N_39527);
nand U42871 (N_42871,N_37393,N_36655);
nand U42872 (N_42872,N_30918,N_35113);
or U42873 (N_42873,N_36197,N_36777);
and U42874 (N_42874,N_38861,N_36425);
and U42875 (N_42875,N_38505,N_36695);
nand U42876 (N_42876,N_32885,N_34199);
or U42877 (N_42877,N_39794,N_33983);
or U42878 (N_42878,N_34245,N_32502);
xnor U42879 (N_42879,N_39901,N_39553);
nand U42880 (N_42880,N_35392,N_36046);
and U42881 (N_42881,N_34269,N_37888);
nor U42882 (N_42882,N_34291,N_36797);
xnor U42883 (N_42883,N_35477,N_35852);
xnor U42884 (N_42884,N_39709,N_37494);
and U42885 (N_42885,N_31479,N_35577);
nor U42886 (N_42886,N_30111,N_34400);
and U42887 (N_42887,N_38042,N_36599);
or U42888 (N_42888,N_32682,N_36810);
nor U42889 (N_42889,N_35396,N_32106);
xnor U42890 (N_42890,N_38312,N_30657);
xnor U42891 (N_42891,N_31989,N_32926);
nor U42892 (N_42892,N_35386,N_30312);
nor U42893 (N_42893,N_38117,N_31935);
nand U42894 (N_42894,N_30516,N_37111);
xnor U42895 (N_42895,N_33347,N_36564);
nor U42896 (N_42896,N_30465,N_36230);
nor U42897 (N_42897,N_30205,N_36280);
xor U42898 (N_42898,N_34246,N_37000);
xor U42899 (N_42899,N_30773,N_33159);
and U42900 (N_42900,N_30396,N_37096);
xnor U42901 (N_42901,N_30216,N_34363);
nor U42902 (N_42902,N_31743,N_33323);
and U42903 (N_42903,N_39224,N_38598);
nor U42904 (N_42904,N_38620,N_35393);
or U42905 (N_42905,N_35746,N_38255);
nor U42906 (N_42906,N_37518,N_34810);
nand U42907 (N_42907,N_38416,N_37950);
or U42908 (N_42908,N_34661,N_35293);
and U42909 (N_42909,N_37082,N_34879);
nor U42910 (N_42910,N_33214,N_32147);
xor U42911 (N_42911,N_34288,N_35084);
nor U42912 (N_42912,N_37419,N_38037);
nand U42913 (N_42913,N_31356,N_31845);
nand U42914 (N_42914,N_37032,N_32067);
nand U42915 (N_42915,N_35257,N_34270);
xor U42916 (N_42916,N_32032,N_35136);
or U42917 (N_42917,N_34293,N_31142);
or U42918 (N_42918,N_37253,N_32967);
nor U42919 (N_42919,N_37766,N_36489);
nand U42920 (N_42920,N_37689,N_34972);
or U42921 (N_42921,N_32936,N_34815);
and U42922 (N_42922,N_31795,N_35464);
xor U42923 (N_42923,N_39239,N_31861);
nand U42924 (N_42924,N_39194,N_36925);
xnor U42925 (N_42925,N_33015,N_36595);
nor U42926 (N_42926,N_30254,N_34356);
nor U42927 (N_42927,N_31052,N_35790);
or U42928 (N_42928,N_31396,N_34753);
or U42929 (N_42929,N_32624,N_35678);
nand U42930 (N_42930,N_38334,N_36211);
and U42931 (N_42931,N_33566,N_36656);
nor U42932 (N_42932,N_32505,N_31610);
and U42933 (N_42933,N_36166,N_31701);
nand U42934 (N_42934,N_35734,N_33407);
or U42935 (N_42935,N_37220,N_34504);
nor U42936 (N_42936,N_39447,N_33562);
xnor U42937 (N_42937,N_34768,N_37109);
xor U42938 (N_42938,N_38144,N_35718);
nand U42939 (N_42939,N_35306,N_31900);
nor U42940 (N_42940,N_38394,N_34335);
and U42941 (N_42941,N_37198,N_31264);
or U42942 (N_42942,N_37434,N_31380);
or U42943 (N_42943,N_39335,N_35475);
nand U42944 (N_42944,N_34353,N_34653);
or U42945 (N_42945,N_38923,N_33095);
and U42946 (N_42946,N_38695,N_37076);
or U42947 (N_42947,N_30774,N_36649);
nor U42948 (N_42948,N_38579,N_31163);
xor U42949 (N_42949,N_38752,N_32546);
nand U42950 (N_42950,N_35508,N_30342);
nand U42951 (N_42951,N_39116,N_37600);
xor U42952 (N_42952,N_34092,N_30333);
nand U42953 (N_42953,N_36460,N_36167);
nand U42954 (N_42954,N_35960,N_36568);
xnor U42955 (N_42955,N_32412,N_36528);
and U42956 (N_42956,N_35099,N_37423);
nand U42957 (N_42957,N_37235,N_37226);
nand U42958 (N_42958,N_30197,N_32009);
nor U42959 (N_42959,N_37929,N_38846);
nor U42960 (N_42960,N_30083,N_36330);
nor U42961 (N_42961,N_37603,N_35901);
and U42962 (N_42962,N_34668,N_36737);
nor U42963 (N_42963,N_30997,N_30075);
xnor U42964 (N_42964,N_37069,N_38476);
and U42965 (N_42965,N_30803,N_35119);
or U42966 (N_42966,N_31075,N_31434);
or U42967 (N_42967,N_34324,N_33732);
nor U42968 (N_42968,N_37239,N_30484);
xor U42969 (N_42969,N_37583,N_30541);
xnor U42970 (N_42970,N_37401,N_37058);
nand U42971 (N_42971,N_33286,N_35500);
nor U42972 (N_42972,N_36637,N_32910);
nand U42973 (N_42973,N_32952,N_33303);
xor U42974 (N_42974,N_35765,N_36835);
xnor U42975 (N_42975,N_39252,N_30012);
xor U42976 (N_42976,N_36207,N_30190);
nor U42977 (N_42977,N_36439,N_37015);
or U42978 (N_42978,N_33754,N_39573);
xor U42979 (N_42979,N_32981,N_35589);
or U42980 (N_42980,N_31427,N_32536);
or U42981 (N_42981,N_35344,N_39416);
nand U42982 (N_42982,N_37503,N_34892);
xor U42983 (N_42983,N_37755,N_30151);
or U42984 (N_42984,N_34452,N_35796);
and U42985 (N_42985,N_34162,N_33179);
xnor U42986 (N_42986,N_30829,N_37405);
and U42987 (N_42987,N_39186,N_38803);
nand U42988 (N_42988,N_36187,N_33230);
xnor U42989 (N_42989,N_36234,N_37936);
nand U42990 (N_42990,N_30471,N_39806);
nand U42991 (N_42991,N_36617,N_33085);
nand U42992 (N_42992,N_36944,N_36215);
nor U42993 (N_42993,N_31715,N_30712);
nand U42994 (N_42994,N_36602,N_39387);
xnor U42995 (N_42995,N_32215,N_32033);
xor U42996 (N_42996,N_39493,N_32053);
xnor U42997 (N_42997,N_33871,N_34425);
nand U42998 (N_42998,N_30436,N_32701);
nand U42999 (N_42999,N_35286,N_34695);
nor U43000 (N_43000,N_30429,N_36514);
nand U43001 (N_43001,N_36534,N_34739);
xnor U43002 (N_43002,N_31009,N_37853);
nor U43003 (N_43003,N_34307,N_30863);
xor U43004 (N_43004,N_39231,N_33841);
nand U43005 (N_43005,N_37101,N_31718);
nor U43006 (N_43006,N_36137,N_37145);
and U43007 (N_43007,N_34974,N_32874);
nand U43008 (N_43008,N_33251,N_37056);
or U43009 (N_43009,N_37141,N_39458);
or U43010 (N_43010,N_33177,N_34126);
nand U43011 (N_43011,N_33130,N_34357);
nand U43012 (N_43012,N_36573,N_32438);
nor U43013 (N_43013,N_33596,N_36010);
xor U43014 (N_43014,N_30295,N_39390);
nand U43015 (N_43015,N_38609,N_30830);
nor U43016 (N_43016,N_35252,N_39779);
nor U43017 (N_43017,N_30163,N_30183);
or U43018 (N_43018,N_31312,N_31639);
nand U43019 (N_43019,N_37377,N_39047);
nor U43020 (N_43020,N_33675,N_38748);
nand U43021 (N_43021,N_31370,N_36172);
xnor U43022 (N_43022,N_33019,N_35142);
nand U43023 (N_43023,N_35905,N_32864);
nor U43024 (N_43024,N_36561,N_38365);
and U43025 (N_43025,N_33888,N_34257);
or U43026 (N_43026,N_30847,N_31887);
nor U43027 (N_43027,N_35671,N_34160);
and U43028 (N_43028,N_31185,N_30195);
xor U43029 (N_43029,N_31635,N_35305);
or U43030 (N_43030,N_37090,N_38330);
nand U43031 (N_43031,N_34268,N_34779);
xor U43032 (N_43032,N_35881,N_32379);
xor U43033 (N_43033,N_38474,N_32212);
and U43034 (N_43034,N_39334,N_33237);
or U43035 (N_43035,N_31360,N_30479);
and U43036 (N_43036,N_32024,N_30565);
and U43037 (N_43037,N_33646,N_37389);
or U43038 (N_43038,N_37565,N_39080);
or U43039 (N_43039,N_31914,N_37690);
nand U43040 (N_43040,N_30023,N_35793);
and U43041 (N_43041,N_39981,N_39733);
and U43042 (N_43042,N_39411,N_37750);
xor U43043 (N_43043,N_31824,N_36435);
and U43044 (N_43044,N_39179,N_31151);
or U43045 (N_43045,N_33368,N_32794);
and U43046 (N_43046,N_37311,N_33519);
xor U43047 (N_43047,N_33890,N_30769);
or U43048 (N_43048,N_38383,N_37870);
xor U43049 (N_43049,N_33560,N_34719);
or U43050 (N_43050,N_35334,N_35411);
nand U43051 (N_43051,N_39112,N_36696);
and U43052 (N_43052,N_39076,N_39741);
or U43053 (N_43053,N_30513,N_33035);
or U43054 (N_43054,N_30592,N_35639);
or U43055 (N_43055,N_39623,N_32115);
nor U43056 (N_43056,N_35270,N_38812);
nor U43057 (N_43057,N_31222,N_35669);
nor U43058 (N_43058,N_35192,N_32133);
or U43059 (N_43059,N_35037,N_30625);
or U43060 (N_43060,N_34806,N_39586);
and U43061 (N_43061,N_36469,N_35783);
nand U43062 (N_43062,N_31981,N_31231);
and U43063 (N_43063,N_33680,N_32935);
nand U43064 (N_43064,N_34970,N_33127);
nor U43065 (N_43065,N_33970,N_37681);
or U43066 (N_43066,N_30349,N_33341);
nand U43067 (N_43067,N_33449,N_35090);
nand U43068 (N_43068,N_32150,N_33748);
nor U43069 (N_43069,N_34402,N_38347);
xnor U43070 (N_43070,N_32309,N_30958);
nand U43071 (N_43071,N_35618,N_37608);
nand U43072 (N_43072,N_34421,N_35697);
nor U43073 (N_43073,N_33487,N_34398);
and U43074 (N_43074,N_37177,N_33187);
and U43075 (N_43075,N_38477,N_35204);
nand U43076 (N_43076,N_38317,N_36748);
nor U43077 (N_43077,N_30550,N_39492);
nor U43078 (N_43078,N_36999,N_34255);
xor U43079 (N_43079,N_33222,N_35288);
and U43080 (N_43080,N_35379,N_39930);
or U43081 (N_43081,N_31764,N_38283);
nand U43082 (N_43082,N_33213,N_35123);
nor U43083 (N_43083,N_38145,N_38186);
and U43084 (N_43084,N_31316,N_36363);
nor U43085 (N_43085,N_38009,N_37904);
nand U43086 (N_43086,N_33181,N_34379);
nand U43087 (N_43087,N_30564,N_32070);
nor U43088 (N_43088,N_31062,N_31816);
or U43089 (N_43089,N_34351,N_33276);
or U43090 (N_43090,N_35999,N_32040);
nand U43091 (N_43091,N_36913,N_32181);
nor U43092 (N_43092,N_31109,N_39312);
and U43093 (N_43093,N_34279,N_33274);
nor U43094 (N_43094,N_39590,N_34285);
nand U43095 (N_43095,N_38843,N_31302);
nand U43096 (N_43096,N_35426,N_32716);
xnor U43097 (N_43097,N_30916,N_37375);
and U43098 (N_43098,N_38352,N_36668);
xnor U43099 (N_43099,N_35509,N_33284);
or U43100 (N_43100,N_30811,N_38727);
and U43101 (N_43101,N_34231,N_33207);
xor U43102 (N_43102,N_31147,N_33955);
and U43103 (N_43103,N_35719,N_34890);
nor U43104 (N_43104,N_31375,N_31094);
nand U43105 (N_43105,N_34086,N_38685);
or U43106 (N_43106,N_39631,N_31922);
nand U43107 (N_43107,N_38072,N_39798);
nor U43108 (N_43108,N_32047,N_34367);
or U43109 (N_43109,N_32071,N_39881);
or U43110 (N_43110,N_30099,N_34798);
xor U43111 (N_43111,N_31680,N_36915);
nand U43112 (N_43112,N_30887,N_32078);
nor U43113 (N_43113,N_32251,N_39870);
and U43114 (N_43114,N_36099,N_31564);
or U43115 (N_43115,N_32015,N_38491);
nor U43116 (N_43116,N_30250,N_37735);
or U43117 (N_43117,N_33829,N_34851);
nand U43118 (N_43118,N_33734,N_35874);
and U43119 (N_43119,N_32380,N_32013);
and U43120 (N_43120,N_35077,N_39191);
nor U43121 (N_43121,N_32946,N_30555);
or U43122 (N_43122,N_32815,N_30384);
nor U43123 (N_43123,N_39676,N_30842);
and U43124 (N_43124,N_32766,N_31198);
and U43125 (N_43125,N_30030,N_35225);
and U43126 (N_43126,N_32588,N_37846);
xnor U43127 (N_43127,N_35312,N_31456);
or U43128 (N_43128,N_38409,N_38657);
and U43129 (N_43129,N_38597,N_38700);
or U43130 (N_43130,N_30900,N_39197);
nor U43131 (N_43131,N_34553,N_31836);
or U43132 (N_43132,N_36070,N_35201);
nand U43133 (N_43133,N_36675,N_36345);
nor U43134 (N_43134,N_31490,N_32452);
and U43135 (N_43135,N_35893,N_39372);
or U43136 (N_43136,N_38033,N_30166);
or U43137 (N_43137,N_35340,N_36191);
nor U43138 (N_43138,N_37264,N_36796);
xnor U43139 (N_43139,N_34837,N_33978);
xor U43140 (N_43140,N_37784,N_38852);
xnor U43141 (N_43141,N_30466,N_35927);
nor U43142 (N_43142,N_31725,N_34330);
or U43143 (N_43143,N_39367,N_38557);
nand U43144 (N_43144,N_32930,N_30076);
nor U43145 (N_43145,N_35733,N_35803);
nor U43146 (N_43146,N_34023,N_35947);
and U43147 (N_43147,N_37562,N_39379);
or U43148 (N_43148,N_39324,N_39660);
and U43149 (N_43149,N_38512,N_31493);
nand U43150 (N_43150,N_38192,N_31961);
nand U43151 (N_43151,N_37443,N_39530);
or U43152 (N_43152,N_35321,N_39049);
xnor U43153 (N_43153,N_38759,N_32475);
xnor U43154 (N_43154,N_34211,N_34114);
xor U43155 (N_43155,N_34404,N_36998);
nand U43156 (N_43156,N_36754,N_38127);
or U43157 (N_43157,N_38396,N_36490);
nor U43158 (N_43158,N_34629,N_32177);
and U43159 (N_43159,N_34809,N_37978);
nand U43160 (N_43160,N_35864,N_34542);
and U43161 (N_43161,N_39944,N_31555);
nor U43162 (N_43162,N_39277,N_30850);
or U43163 (N_43163,N_31653,N_36712);
nand U43164 (N_43164,N_32714,N_38046);
or U43165 (N_43165,N_34586,N_36143);
nand U43166 (N_43166,N_33162,N_37490);
and U43167 (N_43167,N_34639,N_31067);
and U43168 (N_43168,N_39188,N_39249);
nor U43169 (N_43169,N_35711,N_32382);
or U43170 (N_43170,N_37179,N_38030);
nand U43171 (N_43171,N_36501,N_36549);
or U43172 (N_43172,N_35547,N_31032);
nand U43173 (N_43173,N_36763,N_39423);
and U43174 (N_43174,N_34712,N_38641);
and U43175 (N_43175,N_39108,N_34992);
nor U43176 (N_43176,N_38739,N_33800);
nand U43177 (N_43177,N_36076,N_33511);
nand U43178 (N_43178,N_37779,N_34789);
nor U43179 (N_43179,N_32750,N_31857);
nand U43180 (N_43180,N_30643,N_31589);
xnor U43181 (N_43181,N_31496,N_32068);
and U43182 (N_43182,N_39200,N_31125);
nor U43183 (N_43183,N_38906,N_34489);
or U43184 (N_43184,N_36535,N_30533);
xnor U43185 (N_43185,N_39229,N_34010);
or U43186 (N_43186,N_30212,N_32164);
nand U43187 (N_43187,N_35035,N_36173);
nand U43188 (N_43188,N_31255,N_31457);
nor U43189 (N_43189,N_37945,N_30722);
nor U43190 (N_43190,N_31677,N_39244);
or U43191 (N_43191,N_38655,N_36611);
or U43192 (N_43192,N_30534,N_38074);
nand U43193 (N_43193,N_36583,N_37055);
nor U43194 (N_43194,N_30200,N_32272);
nor U43195 (N_43195,N_35220,N_37221);
xnor U43196 (N_43196,N_35349,N_35222);
or U43197 (N_43197,N_37046,N_39290);
and U43198 (N_43198,N_38390,N_34169);
and U43199 (N_43199,N_38981,N_39936);
or U43200 (N_43200,N_36019,N_33864);
nor U43201 (N_43201,N_36342,N_38420);
nand U43202 (N_43202,N_35968,N_35611);
nor U43203 (N_43203,N_30457,N_32529);
xor U43204 (N_43204,N_36868,N_32271);
nor U43205 (N_43205,N_37413,N_31203);
or U43206 (N_43206,N_34127,N_36171);
nand U43207 (N_43207,N_37530,N_37318);
and U43208 (N_43208,N_34390,N_38290);
and U43209 (N_43209,N_39095,N_32709);
nand U43210 (N_43210,N_36862,N_30243);
xnor U43211 (N_43211,N_35030,N_32638);
and U43212 (N_43212,N_38970,N_34442);
or U43213 (N_43213,N_32002,N_39997);
nand U43214 (N_43214,N_38277,N_38212);
nor U43215 (N_43215,N_34435,N_33398);
or U43216 (N_43216,N_31395,N_37881);
or U43217 (N_43217,N_35097,N_30987);
xnor U43218 (N_43218,N_35997,N_33578);
nor U43219 (N_43219,N_34591,N_38594);
nand U43220 (N_43220,N_35320,N_37655);
nand U43221 (N_43221,N_37957,N_39621);
nand U43222 (N_43222,N_38472,N_30779);
nor U43223 (N_43223,N_36333,N_30980);
and U43224 (N_43224,N_30367,N_33521);
nor U43225 (N_43225,N_33436,N_39321);
nand U43226 (N_43226,N_38819,N_30646);
nand U43227 (N_43227,N_38827,N_37767);
nor U43228 (N_43228,N_30585,N_36537);
or U43229 (N_43229,N_35149,N_32092);
and U43230 (N_43230,N_32180,N_36581);
or U43231 (N_43231,N_37379,N_36811);
nand U43232 (N_43232,N_30936,N_32214);
nand U43233 (N_43233,N_32148,N_39456);
xor U43234 (N_43234,N_32593,N_34963);
nand U43235 (N_43235,N_37126,N_38455);
nand U43236 (N_43236,N_38328,N_38392);
and U43237 (N_43237,N_36351,N_36206);
xor U43238 (N_43238,N_39298,N_36136);
nand U43239 (N_43239,N_33298,N_33180);
nor U43240 (N_43240,N_39791,N_34009);
and U43241 (N_43241,N_31920,N_34658);
nand U43242 (N_43242,N_34901,N_33047);
nand U43243 (N_43243,N_32524,N_32321);
nor U43244 (N_43244,N_33247,N_33389);
xnor U43245 (N_43245,N_31539,N_36706);
xor U43246 (N_43246,N_36079,N_35755);
or U43247 (N_43247,N_30145,N_32785);
or U43248 (N_43248,N_32479,N_34930);
nand U43249 (N_43249,N_38232,N_34161);
xnor U43250 (N_43250,N_36634,N_37108);
and U43251 (N_43251,N_32856,N_34796);
nor U43252 (N_43252,N_32270,N_35993);
or U43253 (N_43253,N_39500,N_39313);
and U43254 (N_43254,N_35052,N_32540);
nor U43255 (N_43255,N_38524,N_36778);
nor U43256 (N_43256,N_30919,N_32724);
nand U43257 (N_43257,N_34076,N_39209);
xor U43258 (N_43258,N_39386,N_39024);
nand U43259 (N_43259,N_33586,N_36370);
nand U43260 (N_43260,N_32126,N_37891);
nand U43261 (N_43261,N_33641,N_39206);
xor U43262 (N_43262,N_39355,N_38562);
xor U43263 (N_43263,N_32840,N_36746);
and U43264 (N_43264,N_37614,N_32659);
xnor U43265 (N_43265,N_38875,N_34112);
or U43266 (N_43266,N_38258,N_37930);
xor U43267 (N_43267,N_30967,N_35140);
and U43268 (N_43268,N_32004,N_34371);
nor U43269 (N_43269,N_35703,N_38259);
nor U43270 (N_43270,N_34807,N_31597);
xnor U43271 (N_43271,N_35919,N_33966);
and U43272 (N_43272,N_30366,N_30070);
nand U43273 (N_43273,N_35398,N_35777);
nor U43274 (N_43274,N_39013,N_39955);
nor U43275 (N_43275,N_39350,N_38722);
nand U43276 (N_43276,N_37187,N_30733);
or U43277 (N_43277,N_35471,N_37629);
or U43278 (N_43278,N_36762,N_37073);
xor U43279 (N_43279,N_37682,N_30631);
and U43280 (N_43280,N_37907,N_31915);
or U43281 (N_43281,N_33226,N_30586);
or U43282 (N_43282,N_37801,N_34678);
xor U43283 (N_43283,N_32782,N_34782);
xor U43284 (N_43284,N_39398,N_33750);
or U43285 (N_43285,N_35354,N_38244);
xnor U43286 (N_43286,N_33014,N_32313);
nor U43287 (N_43287,N_38197,N_38191);
nor U43288 (N_43288,N_31991,N_39851);
nor U43289 (N_43289,N_36180,N_32210);
nand U43290 (N_43290,N_30459,N_35795);
nand U43291 (N_43291,N_30313,N_32859);
xnor U43292 (N_43292,N_33279,N_33624);
xnor U43293 (N_43293,N_36252,N_32979);
xor U43294 (N_43294,N_38706,N_32940);
nor U43295 (N_43295,N_30873,N_36781);
nor U43296 (N_43296,N_30290,N_37332);
or U43297 (N_43297,N_34031,N_36761);
or U43298 (N_43298,N_33702,N_37722);
and U43299 (N_43299,N_35680,N_37864);
or U43300 (N_43300,N_30504,N_36368);
nor U43301 (N_43301,N_36819,N_36476);
or U43302 (N_43302,N_35150,N_32229);
or U43303 (N_43303,N_36728,N_33882);
nor U43304 (N_43304,N_38374,N_39418);
xnor U43305 (N_43305,N_36522,N_32679);
nor U43306 (N_43306,N_38282,N_33086);
xor U43307 (N_43307,N_31023,N_30453);
xnor U43308 (N_43308,N_39643,N_36141);
and U43309 (N_43309,N_37002,N_37461);
and U43310 (N_43310,N_38493,N_35195);
nor U43311 (N_43311,N_38636,N_37780);
or U43312 (N_43312,N_35240,N_34278);
or U43313 (N_43313,N_34142,N_33889);
nand U43314 (N_43314,N_33842,N_34228);
nor U43315 (N_43315,N_39987,N_31401);
xor U43316 (N_43316,N_37440,N_30324);
xor U43317 (N_43317,N_34328,N_36597);
xnor U43318 (N_43318,N_32154,N_38119);
nor U43319 (N_43319,N_36653,N_31572);
nand U43320 (N_43320,N_34817,N_35278);
xnor U43321 (N_43321,N_37029,N_38558);
nor U43322 (N_43322,N_37761,N_38710);
nand U43323 (N_43323,N_38492,N_34677);
and U43324 (N_43324,N_36029,N_37883);
xor U43325 (N_43325,N_30419,N_30439);
or U43326 (N_43326,N_39354,N_39659);
nor U43327 (N_43327,N_38667,N_37241);
and U43328 (N_43328,N_30582,N_37080);
or U43329 (N_43329,N_38673,N_30089);
or U43330 (N_43330,N_38932,N_30193);
nor U43331 (N_43331,N_35264,N_30043);
and U43332 (N_43332,N_36134,N_32245);
and U43333 (N_43333,N_36606,N_35339);
nor U43334 (N_43334,N_34047,N_37444);
or U43335 (N_43335,N_30729,N_30525);
nand U43336 (N_43336,N_30975,N_34414);
and U43337 (N_43337,N_31579,N_38630);
or U43338 (N_43338,N_34497,N_34444);
nand U43339 (N_43339,N_37036,N_33804);
and U43340 (N_43340,N_33404,N_38314);
nor U43341 (N_43341,N_30469,N_33553);
and U43342 (N_43342,N_38887,N_39276);
nor U43343 (N_43343,N_32136,N_35972);
xnor U43344 (N_43344,N_33450,N_37878);
or U43345 (N_43345,N_35044,N_31196);
xor U43346 (N_43346,N_34691,N_32520);
or U43347 (N_43347,N_34528,N_32419);
xnor U43348 (N_43348,N_37161,N_38026);
nand U43349 (N_43349,N_39343,N_36246);
and U43350 (N_43350,N_37817,N_30578);
and U43351 (N_43351,N_34977,N_30968);
nand U43352 (N_43352,N_39294,N_34800);
or U43353 (N_43353,N_31518,N_38263);
and U43354 (N_43354,N_34487,N_32951);
or U43355 (N_43355,N_38724,N_32500);
nor U43356 (N_43356,N_33108,N_37106);
nand U43357 (N_43357,N_36131,N_32892);
nor U43358 (N_43358,N_34299,N_38740);
and U43359 (N_43359,N_37663,N_32001);
or U43360 (N_43360,N_35832,N_37228);
nand U43361 (N_43361,N_39698,N_34458);
xnor U43362 (N_43362,N_34917,N_36237);
nand U43363 (N_43363,N_32813,N_36521);
nor U43364 (N_43364,N_30098,N_34141);
nor U43365 (N_43365,N_32290,N_31875);
xor U43366 (N_43366,N_37627,N_36411);
nor U43367 (N_43367,N_38957,N_35637);
nand U43368 (N_43368,N_36570,N_34763);
xnor U43369 (N_43369,N_32166,N_38913);
nor U43370 (N_43370,N_32422,N_35175);
xor U43371 (N_43371,N_39633,N_32670);
and U43372 (N_43372,N_31893,N_39450);
nor U43373 (N_43373,N_38719,N_38862);
or U43374 (N_43374,N_33569,N_39033);
nand U43375 (N_43375,N_39286,N_37131);
nor U43376 (N_43376,N_34567,N_30865);
nand U43377 (N_43377,N_38918,N_37900);
nor U43378 (N_43378,N_37520,N_36367);
nor U43379 (N_43379,N_33369,N_36379);
or U43380 (N_43380,N_32301,N_39265);
xnor U43381 (N_43381,N_32050,N_36773);
and U43382 (N_43382,N_38877,N_33856);
nor U43383 (N_43383,N_34450,N_37366);
nor U43384 (N_43384,N_34247,N_36289);
nand U43385 (N_43385,N_32037,N_31676);
and U43386 (N_43386,N_38658,N_37189);
and U43387 (N_43387,N_35249,N_32403);
xnor U43388 (N_43388,N_39574,N_36464);
and U43389 (N_43389,N_33062,N_38576);
nor U43390 (N_43390,N_39414,N_38321);
xnor U43391 (N_43391,N_39545,N_37589);
or U43392 (N_43392,N_37312,N_38632);
and U43393 (N_43393,N_38089,N_33968);
and U43394 (N_43394,N_31390,N_38154);
nand U43395 (N_43395,N_38584,N_37304);
nand U43396 (N_43396,N_38530,N_35151);
nand U43397 (N_43397,N_32283,N_30566);
xnor U43398 (N_43398,N_35658,N_33184);
xor U43399 (N_43399,N_32537,N_33088);
and U43400 (N_43400,N_39756,N_39315);
and U43401 (N_43401,N_35717,N_35581);
nor U43402 (N_43402,N_30330,N_32060);
and U43403 (N_43403,N_35619,N_33232);
nand U43404 (N_43404,N_35770,N_36952);
nor U43405 (N_43405,N_35752,N_30438);
or U43406 (N_43406,N_39919,N_34593);
nor U43407 (N_43407,N_31982,N_39430);
nand U43408 (N_43408,N_37677,N_39260);
or U43409 (N_43409,N_33648,N_30738);
and U43410 (N_43410,N_38801,N_31546);
and U43411 (N_43411,N_33268,N_38128);
or U43412 (N_43412,N_36120,N_32838);
nor U43413 (N_43413,N_31364,N_39747);
nand U43414 (N_43414,N_37564,N_37541);
nor U43415 (N_43415,N_36890,N_33068);
nand U43416 (N_43416,N_36779,N_31952);
xor U43417 (N_43417,N_39594,N_32336);
nand U43418 (N_43418,N_39781,N_37822);
nand U43419 (N_43419,N_32564,N_39846);
or U43420 (N_43420,N_33006,N_36443);
xor U43421 (N_43421,N_37642,N_34898);
nor U43422 (N_43422,N_36282,N_39865);
nor U43423 (N_43423,N_38105,N_38100);
nand U43424 (N_43424,N_35423,N_31403);
nand U43425 (N_43425,N_34032,N_30563);
or U43426 (N_43426,N_32415,N_37023);
and U43427 (N_43427,N_32773,N_36750);
and U43428 (N_43428,N_33652,N_39477);
nand U43429 (N_43429,N_37577,N_30977);
and U43430 (N_43430,N_32622,N_32114);
nand U43431 (N_43431,N_35744,N_35147);
xor U43432 (N_43432,N_33653,N_35899);
and U43433 (N_43433,N_31955,N_34473);
and U43434 (N_43434,N_37579,N_38209);
xor U43435 (N_43435,N_38096,N_35025);
nand U43436 (N_43436,N_34558,N_33318);
xnor U43437 (N_43437,N_31647,N_32297);
and U43438 (N_43438,N_38998,N_39702);
xnor U43439 (N_43439,N_36747,N_30114);
xor U43440 (N_43440,N_34383,N_36594);
nor U43441 (N_43441,N_32226,N_34551);
or U43442 (N_43442,N_30045,N_34369);
xnor U43443 (N_43443,N_35170,N_34943);
or U43444 (N_43444,N_34549,N_35430);
nand U43445 (N_43445,N_31111,N_34480);
nor U43446 (N_43446,N_38065,N_32535);
or U43447 (N_43447,N_38495,N_38565);
xnor U43448 (N_43448,N_35493,N_31266);
and U43449 (N_43449,N_39434,N_37233);
and U43450 (N_43450,N_35507,N_37851);
xnor U43451 (N_43451,N_31399,N_33171);
nor U43452 (N_43452,N_36828,N_33329);
and U43453 (N_43453,N_38247,N_34192);
xor U43454 (N_43454,N_34666,N_39583);
xnor U43455 (N_43455,N_34936,N_31453);
and U43456 (N_43456,N_35163,N_34311);
or U43457 (N_43457,N_31211,N_35485);
and U43458 (N_43458,N_38856,N_32291);
or U43459 (N_43459,N_31531,N_31180);
and U43460 (N_43460,N_37112,N_34075);
nand U43461 (N_43461,N_33827,N_39257);
nor U43462 (N_43462,N_30080,N_32788);
and U43463 (N_43463,N_35553,N_36860);
nor U43464 (N_43464,N_35545,N_33722);
and U43465 (N_43465,N_39663,N_30371);
xor U43466 (N_43466,N_33982,N_36736);
nand U43467 (N_43467,N_38965,N_39483);
or U43468 (N_43468,N_32542,N_36243);
nor U43469 (N_43469,N_37925,N_38942);
and U43470 (N_43470,N_37165,N_33743);
and U43471 (N_43471,N_35518,N_31477);
xnor U43472 (N_43472,N_32913,N_33446);
xnor U43473 (N_43473,N_38398,N_32704);
nand U43474 (N_43474,N_35689,N_38693);
nand U43475 (N_43475,N_39830,N_35224);
xnor U43476 (N_43476,N_36963,N_38486);
and U43477 (N_43477,N_39871,N_38661);
nor U43478 (N_43478,N_30069,N_36012);
xor U43479 (N_43479,N_35026,N_39685);
nor U43480 (N_43480,N_34721,N_37534);
nor U43481 (N_43481,N_37320,N_30757);
or U43482 (N_43482,N_35701,N_36213);
nor U43483 (N_43483,N_30148,N_38735);
xnor U43484 (N_43484,N_31928,N_34465);
and U43485 (N_43485,N_33726,N_30707);
nor U43486 (N_43486,N_38984,N_34016);
nor U43487 (N_43487,N_33002,N_30767);
or U43488 (N_43488,N_32073,N_37775);
nand U43489 (N_43489,N_36624,N_32748);
nor U43490 (N_43490,N_34171,N_39373);
xor U43491 (N_43491,N_32811,N_33588);
nand U43492 (N_43492,N_30442,N_38668);
and U43493 (N_43493,N_37367,N_36325);
and U43494 (N_43494,N_38231,N_39007);
nor U43495 (N_43495,N_31287,N_31895);
xor U43496 (N_43496,N_37595,N_32745);
and U43497 (N_43497,N_30788,N_35660);
nor U43498 (N_43498,N_34735,N_38844);
and U43499 (N_43499,N_31176,N_37717);
and U43500 (N_43500,N_34840,N_33631);
xor U43501 (N_43501,N_31792,N_39030);
nor U43502 (N_43502,N_36150,N_36111);
nor U43503 (N_43503,N_37538,N_32027);
xor U43504 (N_43504,N_34344,N_32235);
or U43505 (N_43505,N_32370,N_30925);
nand U43506 (N_43506,N_34197,N_31652);
and U43507 (N_43507,N_34869,N_39211);
and U43508 (N_43508,N_36181,N_35794);
nor U43509 (N_43509,N_33480,N_31431);
nor U43510 (N_43510,N_30768,N_31265);
xnor U43511 (N_43511,N_35863,N_33362);
and U43512 (N_43512,N_39645,N_31937);
xor U43513 (N_43513,N_37194,N_30571);
and U43514 (N_43514,N_34904,N_35189);
nor U43515 (N_43515,N_34625,N_31874);
nand U43516 (N_43516,N_33252,N_39994);
or U43517 (N_43517,N_37006,N_37257);
xor U43518 (N_43518,N_39959,N_39528);
xnor U43519 (N_43519,N_34253,N_32483);
xnor U43520 (N_43520,N_31091,N_38712);
xnor U43521 (N_43521,N_34515,N_35924);
or U43522 (N_43522,N_37279,N_39090);
and U43523 (N_43523,N_34692,N_33971);
or U43524 (N_43524,N_36759,N_35336);
or U43525 (N_43525,N_32983,N_32349);
xnor U43526 (N_43526,N_32802,N_30611);
nand U43527 (N_43527,N_33956,N_34517);
xnor U43528 (N_43528,N_35766,N_36685);
xor U43529 (N_43529,N_32198,N_39905);
nand U43530 (N_43530,N_30818,N_33572);
nor U43531 (N_43531,N_32800,N_36905);
nor U43532 (N_43532,N_30969,N_38466);
nand U43533 (N_43533,N_35394,N_35890);
or U43534 (N_43534,N_34456,N_39690);
xor U43535 (N_43535,N_30019,N_30209);
nor U43536 (N_43536,N_38376,N_39023);
xnor U43537 (N_43537,N_37939,N_38549);
xor U43538 (N_43538,N_31770,N_32690);
or U43539 (N_43539,N_34089,N_34833);
and U43540 (N_43540,N_30277,N_33257);
or U43541 (N_43541,N_38546,N_33094);
nand U43542 (N_43542,N_34674,N_32961);
nand U43543 (N_43543,N_39407,N_38339);
or U43544 (N_43544,N_39506,N_35209);
nor U43545 (N_43545,N_37089,N_34893);
xor U43546 (N_43546,N_34572,N_36765);
nand U43547 (N_43547,N_32577,N_35247);
or U43548 (N_43548,N_37823,N_38068);
or U43549 (N_43549,N_35571,N_30291);
xnor U43550 (N_43550,N_33993,N_30765);
and U43551 (N_43551,N_34259,N_38768);
nor U43552 (N_43552,N_31273,N_37231);
xnor U43553 (N_43553,N_39566,N_32372);
xnor U43554 (N_43554,N_39619,N_38581);
and U43555 (N_43555,N_30179,N_32876);
xnor U43556 (N_43556,N_39833,N_31311);
nand U43557 (N_43557,N_30810,N_38526);
nand U43558 (N_43558,N_36184,N_37153);
and U43559 (N_43559,N_37654,N_31501);
xnor U43560 (N_43560,N_38281,N_34604);
and U43561 (N_43561,N_34962,N_31458);
or U43562 (N_43562,N_33584,N_36315);
or U43563 (N_43563,N_30278,N_30104);
or U43564 (N_43564,N_31342,N_36837);
xnor U43565 (N_43565,N_39106,N_33998);
and U43566 (N_43566,N_30362,N_31160);
nor U43567 (N_43567,N_33401,N_31902);
or U43568 (N_43568,N_36100,N_36084);
nand U43569 (N_43569,N_37190,N_30068);
xor U43570 (N_43570,N_39768,N_30727);
or U43571 (N_43571,N_39174,N_33167);
or U43572 (N_43572,N_32329,N_30929);
xor U43573 (N_43573,N_38566,N_39061);
and U43574 (N_43574,N_30383,N_38090);
nor U43575 (N_43575,N_36693,N_35732);
nor U43576 (N_43576,N_39693,N_34987);
and U43577 (N_43577,N_34670,N_34365);
and U43578 (N_43578,N_31933,N_37911);
xor U43579 (N_43579,N_37546,N_38198);
or U43580 (N_43580,N_36151,N_31307);
or U43581 (N_43581,N_32424,N_31019);
and U43582 (N_43582,N_34110,N_37587);
nand U43583 (N_43583,N_32255,N_30642);
and U43584 (N_43584,N_39452,N_36272);
nor U43585 (N_43585,N_38427,N_38612);
nand U43586 (N_43586,N_36324,N_38008);
xnor U43587 (N_43587,N_36970,N_30902);
xnor U43588 (N_43588,N_36506,N_35436);
and U43589 (N_43589,N_31732,N_30187);
and U43590 (N_43590,N_33359,N_33056);
nor U43591 (N_43591,N_34191,N_31306);
nor U43592 (N_43592,N_37987,N_36676);
nor U43593 (N_43593,N_38230,N_34523);
nand U43594 (N_43594,N_38167,N_36389);
or U43595 (N_43595,N_33662,N_34526);
or U43596 (N_43596,N_33149,N_37222);
nand U43597 (N_43597,N_31290,N_36516);
or U43598 (N_43598,N_30441,N_31819);
or U43599 (N_43599,N_36160,N_32371);
nand U43600 (N_43600,N_31793,N_39729);
xnor U43601 (N_43601,N_31003,N_34537);
nor U43602 (N_43602,N_38070,N_34770);
nand U43603 (N_43603,N_32686,N_32978);
nand U43604 (N_43604,N_32695,N_33231);
or U43605 (N_43605,N_30870,N_33338);
xnor U43606 (N_43606,N_36804,N_30208);
nor U43607 (N_43607,N_30380,N_37042);
and U43608 (N_43608,N_37099,N_37347);
and U43609 (N_43609,N_33201,N_34281);
nor U43610 (N_43610,N_37154,N_36080);
nand U43611 (N_43611,N_34514,N_37027);
nor U43612 (N_43612,N_30721,N_36034);
xnor U43613 (N_43613,N_38647,N_32845);
and U43614 (N_43614,N_30952,N_34084);
nor U43615 (N_43615,N_38520,N_31102);
nand U43616 (N_43616,N_35148,N_30420);
xor U43617 (N_43617,N_34412,N_38983);
nand U43618 (N_43618,N_35629,N_34345);
nand U43619 (N_43619,N_33605,N_39875);
nor U43620 (N_43620,N_35716,N_37964);
or U43621 (N_43621,N_34242,N_37770);
xor U43622 (N_43622,N_38892,N_31664);
or U43623 (N_43623,N_35810,N_35957);
nand U43624 (N_43624,N_32584,N_35649);
and U43625 (N_43625,N_30029,N_39811);
nand U43626 (N_43626,N_37207,N_31450);
nor U43627 (N_43627,N_39748,N_32284);
or U43628 (N_43628,N_32100,N_38402);
nor U43629 (N_43629,N_31864,N_37244);
or U43630 (N_43630,N_37030,N_30791);
xnor U43631 (N_43631,N_30475,N_32446);
nor U43632 (N_43632,N_32873,N_33418);
nand U43633 (N_43633,N_36248,N_37959);
and U43634 (N_43634,N_33479,N_38417);
nand U43635 (N_43635,N_37188,N_32139);
xnor U43636 (N_43636,N_39647,N_32541);
or U43637 (N_43637,N_35016,N_32830);
nor U43638 (N_43638,N_30011,N_32528);
nand U43639 (N_43639,N_37079,N_30545);
and U43640 (N_43640,N_35468,N_39208);
or U43641 (N_43641,N_31476,N_39207);
nand U43642 (N_43642,N_33060,N_31104);
xor U43643 (N_43643,N_32591,N_36353);
or U43644 (N_43644,N_38513,N_35723);
and U43645 (N_43645,N_32886,N_31172);
nor U43646 (N_43646,N_30603,N_31592);
or U43647 (N_43647,N_35741,N_32360);
nand U43648 (N_43648,N_31488,N_31362);
and U43649 (N_43649,N_35759,N_34173);
and U43650 (N_43650,N_39882,N_36296);
and U43651 (N_43651,N_30497,N_31591);
and U43652 (N_43652,N_37104,N_34927);
and U43653 (N_43653,N_36813,N_38882);
nand U43654 (N_43654,N_30203,N_38663);
nor U43655 (N_43655,N_37693,N_31873);
nand U43656 (N_43656,N_34830,N_36503);
and U43657 (N_43657,N_30237,N_34494);
nor U43658 (N_43658,N_31964,N_31417);
nor U43659 (N_43659,N_37995,N_37593);
xnor U43660 (N_43660,N_33836,N_31828);
nor U43661 (N_43661,N_33196,N_32579);
and U43662 (N_43662,N_32975,N_33530);
xor U43663 (N_43663,N_34733,N_39163);
nand U43664 (N_43664,N_33761,N_36898);
nor U43665 (N_43665,N_37529,N_31411);
xnor U43666 (N_43666,N_34094,N_39199);
nor U43667 (N_43667,N_37960,N_31841);
nor U43668 (N_43668,N_37991,N_33782);
or U43669 (N_43669,N_35332,N_39307);
nor U43670 (N_43670,N_31537,N_32833);
xor U43671 (N_43671,N_38701,N_32041);
or U43672 (N_43672,N_34234,N_36753);
nand U43673 (N_43673,N_36973,N_38327);
and U43674 (N_43674,N_36931,N_34474);
xor U43675 (N_43675,N_39764,N_37465);
and U43676 (N_43676,N_32257,N_38575);
or U43677 (N_43677,N_32729,N_30674);
nand U43678 (N_43678,N_35511,N_32337);
and U43679 (N_43679,N_37132,N_31085);
or U43680 (N_43680,N_33271,N_36982);
and U43681 (N_43681,N_31394,N_35328);
and U43682 (N_43682,N_30892,N_33545);
nor U43683 (N_43683,N_34420,N_33703);
nand U43684 (N_43684,N_30653,N_31550);
nor U43685 (N_43685,N_39217,N_31992);
xnor U43686 (N_43686,N_34419,N_31627);
xor U43687 (N_43687,N_39555,N_36386);
xnor U43688 (N_43688,N_39760,N_33046);
nor U43689 (N_43689,N_39761,N_31706);
nor U43690 (N_43690,N_39958,N_39442);
or U43691 (N_43691,N_34871,N_38131);
nor U43692 (N_43692,N_31784,N_39347);
and U43693 (N_43693,N_33536,N_38860);
nor U43694 (N_43694,N_30904,N_30247);
and U43695 (N_43695,N_35915,N_34718);
or U43696 (N_43696,N_36885,N_34734);
and U43697 (N_43697,N_39906,N_33370);
nand U43698 (N_43698,N_37501,N_37296);
or U43699 (N_43699,N_36971,N_34641);
and U43700 (N_43700,N_30292,N_33475);
nand U43701 (N_43701,N_32142,N_39706);
nand U43702 (N_43702,N_32121,N_37880);
nand U43703 (N_43703,N_31799,N_33961);
xnor U43704 (N_43704,N_39558,N_32007);
nor U43705 (N_43705,N_36311,N_31489);
nand U43706 (N_43706,N_36128,N_36444);
and U43707 (N_43707,N_31568,N_36218);
or U43708 (N_43708,N_34618,N_31942);
or U43709 (N_43709,N_30743,N_35331);
nand U43710 (N_43710,N_33665,N_39903);
and U43711 (N_43711,N_34439,N_35406);
nand U43712 (N_43712,N_39800,N_34275);
nor U43713 (N_43713,N_34875,N_37114);
nand U43714 (N_43714,N_31229,N_39891);
xor U43715 (N_43715,N_30888,N_31753);
nand U43716 (N_43716,N_35980,N_36467);
or U43717 (N_43717,N_39476,N_34082);
or U43718 (N_43718,N_39765,N_31072);
and U43719 (N_43719,N_30814,N_34433);
nor U43720 (N_43720,N_37384,N_33794);
xor U43721 (N_43721,N_31514,N_35975);
and U43722 (N_43722,N_31105,N_32669);
and U43723 (N_43723,N_36977,N_34808);
or U43724 (N_43724,N_35231,N_38518);
xor U43725 (N_43725,N_33173,N_32163);
nand U43726 (N_43726,N_35713,N_33667);
and U43727 (N_43727,N_36731,N_38075);
or U43728 (N_43728,N_31424,N_37224);
nand U43729 (N_43729,N_32456,N_31508);
or U43730 (N_43730,N_37360,N_37992);
nand U43731 (N_43731,N_34303,N_35065);
nor U43732 (N_43732,N_37330,N_34222);
and U43733 (N_43733,N_35039,N_37953);
nand U43734 (N_43734,N_36937,N_33333);
or U43735 (N_43735,N_37011,N_33851);
xor U43736 (N_43736,N_37937,N_33191);
nor U43737 (N_43737,N_38097,N_36115);
nand U43738 (N_43738,N_37921,N_34289);
xnor U43739 (N_43739,N_39427,N_37178);
and U43740 (N_43740,N_35875,N_30428);
nor U43741 (N_43741,N_31622,N_33216);
xnor U43742 (N_43742,N_33783,N_34471);
and U43743 (N_43743,N_37754,N_31768);
nand U43744 (N_43744,N_32171,N_32907);
nand U43745 (N_43745,N_36867,N_36918);
nor U43746 (N_43746,N_37679,N_38457);
or U43747 (N_43747,N_33009,N_32206);
nor U43748 (N_43748,N_38886,N_31134);
and U43749 (N_43749,N_36683,N_36604);
xnor U43750 (N_43750,N_34174,N_39523);
xor U43751 (N_43751,N_36474,N_36853);
nor U43752 (N_43752,N_30297,N_37502);
nor U43753 (N_43753,N_30879,N_38342);
and U43754 (N_43754,N_31213,N_36826);
xor U43755 (N_43755,N_35588,N_34097);
xor U43756 (N_43756,N_32197,N_36887);
and U43757 (N_43757,N_39235,N_36614);
nor U43758 (N_43758,N_39293,N_34889);
nand U43759 (N_43759,N_32028,N_31202);
or U43760 (N_43760,N_31314,N_39081);
xnor U43761 (N_43761,N_33696,N_31439);
xor U43762 (N_43762,N_37692,N_39429);
and U43763 (N_43763,N_32688,N_31526);
nand U43764 (N_43764,N_38344,N_35348);
nand U43765 (N_43765,N_35261,N_35913);
nand U43766 (N_43766,N_37266,N_36290);
or U43767 (N_43767,N_32947,N_38123);
and U43768 (N_43768,N_33721,N_38747);
or U43769 (N_43769,N_34598,N_39710);
nor U43770 (N_43770,N_32613,N_37382);
xnor U43771 (N_43771,N_37200,N_31910);
or U43772 (N_43772,N_34271,N_36314);
nand U43773 (N_43773,N_38116,N_39143);
nor U43774 (N_43774,N_36175,N_30460);
xor U43775 (N_43775,N_35476,N_36559);
nand U43776 (N_43776,N_36094,N_31629);
or U43777 (N_43777,N_33037,N_33067);
and U43778 (N_43778,N_30694,N_32399);
and U43779 (N_43779,N_32758,N_35258);
nand U43780 (N_43780,N_36681,N_35341);
nand U43781 (N_43781,N_38964,N_32805);
or U43782 (N_43782,N_30908,N_39579);
or U43783 (N_43783,N_36140,N_36093);
and U43784 (N_43784,N_34581,N_30105);
xnor U43785 (N_43785,N_36147,N_34912);
or U43786 (N_43786,N_30123,N_34525);
nor U43787 (N_43787,N_32306,N_36873);
or U43788 (N_43788,N_35657,N_33852);
nand U43789 (N_43789,N_35853,N_38340);
nand U43790 (N_43790,N_39979,N_32664);
nor U43791 (N_43791,N_30156,N_33500);
nand U43792 (N_43792,N_33607,N_36028);
nor U43793 (N_43793,N_38939,N_31749);
xnor U43794 (N_43794,N_34588,N_31089);
and U43795 (N_43795,N_37559,N_31043);
or U43796 (N_43796,N_39078,N_30483);
nor U43797 (N_43797,N_31178,N_39296);
xnor U43798 (N_43798,N_32461,N_37275);
xnor U43799 (N_43799,N_37982,N_37776);
nand U43800 (N_43800,N_30627,N_34134);
nand U43801 (N_43801,N_30473,N_37675);
or U43802 (N_43802,N_37902,N_37540);
or U43803 (N_43803,N_37694,N_37061);
or U43804 (N_43804,N_34434,N_39129);
nor U43805 (N_43805,N_30413,N_34571);
and U43806 (N_43806,N_37547,N_35633);
nor U43807 (N_43807,N_30440,N_34149);
and U43808 (N_43808,N_35600,N_34343);
nand U43809 (N_43809,N_34823,N_32365);
or U43810 (N_43810,N_31852,N_37280);
and U43811 (N_43811,N_30407,N_31901);
xor U43812 (N_43812,N_39345,N_34360);
or U43813 (N_43813,N_30599,N_36292);
nand U43814 (N_43814,N_32052,N_37828);
xor U43815 (N_43815,N_32074,N_33621);
xnor U43816 (N_43816,N_32260,N_31876);
nor U43817 (N_43817,N_35907,N_38449);
nand U43818 (N_43818,N_30241,N_33295);
xnor U43819 (N_43819,N_32621,N_38508);
or U43820 (N_43820,N_34326,N_31777);
nand U43821 (N_43821,N_32972,N_31786);
or U43822 (N_43822,N_38354,N_36878);
and U43823 (N_43823,N_35505,N_35515);
nor U43824 (N_43824,N_31954,N_31199);
xor U43825 (N_43825,N_33650,N_38050);
and U43826 (N_43826,N_31809,N_30185);
nor U43827 (N_43827,N_31398,N_31934);
and U43828 (N_43828,N_31801,N_35965);
nor U43829 (N_43829,N_37281,N_38162);
xnor U43830 (N_43830,N_36631,N_31090);
and U43831 (N_43831,N_37380,N_32649);
xor U43832 (N_43832,N_32626,N_31578);
or U43833 (N_43833,N_33931,N_38371);
nand U43834 (N_43834,N_35814,N_30072);
nand U43835 (N_43835,N_30825,N_31822);
nor U43836 (N_43836,N_37095,N_38816);
nor U43837 (N_43837,N_36959,N_37879);
and U43838 (N_43838,N_38629,N_31925);
or U43839 (N_43839,N_31384,N_38174);
xor U43840 (N_43840,N_39131,N_37218);
nor U43841 (N_43841,N_39569,N_31291);
or U43842 (N_43842,N_35679,N_38173);
nand U43843 (N_43843,N_35613,N_34321);
nand U43844 (N_43844,N_39956,N_36652);
and U43845 (N_43845,N_35000,N_38842);
or U43846 (N_43846,N_37442,N_35295);
xor U43847 (N_43847,N_32738,N_35250);
nor U43848 (N_43848,N_30909,N_38496);
and U43849 (N_43849,N_37158,N_38093);
and U43850 (N_43850,N_39485,N_32059);
or U43851 (N_43851,N_35128,N_36665);
xnor U43852 (N_43852,N_31614,N_32768);
and U43853 (N_43853,N_30950,N_38952);
nor U43854 (N_43854,N_39751,N_39664);
nand U43855 (N_43855,N_34756,N_38183);
nand U43856 (N_43856,N_33769,N_31973);
xor U43857 (N_43857,N_30108,N_37829);
nor U43858 (N_43858,N_39886,N_35169);
xor U43859 (N_43859,N_37487,N_31993);
nand U43860 (N_43860,N_39582,N_33626);
nor U43861 (N_43861,N_35688,N_33913);
nor U43862 (N_43862,N_31365,N_32663);
xnor U43863 (N_43863,N_34096,N_30002);
nand U43864 (N_43864,N_39991,N_38991);
nand U43865 (N_43865,N_31745,N_34903);
xnor U43866 (N_43866,N_38914,N_33809);
or U43867 (N_43867,N_33423,N_37706);
and U43868 (N_43868,N_35782,N_38789);
nor U43869 (N_43869,N_34300,N_34319);
and U43870 (N_43870,N_39261,N_34896);
and U43871 (N_43871,N_36588,N_33272);
and U43872 (N_43872,N_39100,N_31414);
or U43873 (N_43873,N_30276,N_32339);
nor U43874 (N_43874,N_35978,N_33838);
nor U43875 (N_43875,N_35969,N_39967);
and U43876 (N_43876,N_36660,N_31810);
xor U43877 (N_43877,N_32044,N_36667);
and U43878 (N_43878,N_38381,N_30714);
xnor U43879 (N_43879,N_39941,N_31542);
and U43880 (N_43880,N_30485,N_35736);
or U43881 (N_43881,N_32629,N_31423);
or U43882 (N_43882,N_36515,N_31352);
nor U43883 (N_43883,N_34062,N_32927);
xnor U43884 (N_43884,N_34870,N_32715);
or U43885 (N_43885,N_38713,N_35634);
nand U43886 (N_43886,N_39099,N_37736);
and U43887 (N_43887,N_34467,N_36572);
nand U43888 (N_43888,N_38468,N_34116);
xnor U43889 (N_43889,N_33848,N_34113);
xnor U43890 (N_43890,N_36997,N_32396);
and U43891 (N_43891,N_34078,N_32098);
xnor U43892 (N_43892,N_36418,N_30293);
xor U43893 (N_43893,N_39880,N_36757);
nand U43894 (N_43894,N_30561,N_37466);
xnor U43895 (N_43895,N_32778,N_31848);
nand U43896 (N_43896,N_32405,N_35216);
or U43897 (N_43897,N_39843,N_34446);
xnor U43898 (N_43898,N_36532,N_34934);
and U43899 (N_43899,N_36388,N_39299);
nand U43900 (N_43900,N_37763,N_35458);
xnor U43901 (N_43901,N_32671,N_30260);
xnor U43902 (N_43902,N_36834,N_33850);
and U43903 (N_43903,N_35442,N_31270);
xnor U43904 (N_43904,N_34052,N_39133);
xor U43905 (N_43905,N_39766,N_33776);
nor U43906 (N_43906,N_34108,N_36507);
nand U43907 (N_43907,N_34663,N_31936);
nor U43908 (N_43908,N_36789,N_33690);
and U43909 (N_43909,N_33933,N_39291);
xnor U43910 (N_43910,N_32008,N_35737);
xnor U43911 (N_43911,N_37214,N_31623);
and U43912 (N_43912,N_38665,N_35218);
nand U43913 (N_43913,N_30289,N_30404);
or U43914 (N_43914,N_30754,N_34354);
xor U43915 (N_43915,N_32672,N_35473);
nand U43916 (N_43916,N_30016,N_31968);
nor U43917 (N_43917,N_33724,N_35165);
and U43918 (N_43918,N_34432,N_35815);
nor U43919 (N_43919,N_30820,N_32963);
and U43920 (N_43920,N_37364,N_39949);
or U43921 (N_43921,N_33698,N_37783);
xnor U43922 (N_43922,N_35042,N_31829);
nor U43923 (N_43923,N_37855,N_33963);
xor U43924 (N_43924,N_35229,N_36562);
nor U43925 (N_43925,N_30378,N_37942);
and U43926 (N_43926,N_30762,N_39101);
nor U43927 (N_43927,N_31136,N_35420);
or U43928 (N_43928,N_30048,N_30620);
or U43929 (N_43929,N_38828,N_38540);
or U43930 (N_43930,N_32693,N_35057);
xor U43931 (N_43931,N_36526,N_36300);
xnor U43932 (N_43932,N_30332,N_33470);
and U43933 (N_43933,N_34119,N_30323);
or U43934 (N_43934,N_39520,N_38616);
xor U43935 (N_43935,N_30304,N_33574);
and U43936 (N_43936,N_33053,N_30017);
nand U43937 (N_43937,N_30270,N_39836);
xor U43938 (N_43938,N_34748,N_38215);
or U43939 (N_43939,N_34743,N_34844);
xnor U43940 (N_43940,N_32162,N_39567);
nor U43941 (N_43941,N_33311,N_37748);
nand U43942 (N_43942,N_35131,N_36974);
and U43943 (N_43943,N_39040,N_30652);
nor U43944 (N_43944,N_31422,N_34472);
xor U43945 (N_43945,N_37836,N_31607);
nor U43946 (N_43946,N_35431,N_31204);
nor U43947 (N_43947,N_39771,N_38876);
xor U43948 (N_43948,N_30454,N_38809);
xnor U43949 (N_43949,N_30515,N_33357);
nand U43950 (N_43950,N_35203,N_32757);
and U43951 (N_43951,N_32217,N_39378);
nor U43952 (N_43952,N_39380,N_33043);
or U43953 (N_43953,N_37646,N_37669);
nand U43954 (N_43954,N_35243,N_33600);
nand U43955 (N_43955,N_32665,N_34132);
and U43956 (N_43956,N_32532,N_32393);
nand U43957 (N_43957,N_39616,N_33529);
or U43958 (N_43958,N_32601,N_32553);
and U43959 (N_43959,N_38873,N_39939);
and U43960 (N_43960,N_35367,N_34688);
and U43961 (N_43961,N_35503,N_37098);
nand U43962 (N_43962,N_32728,N_38214);
xnor U43963 (N_43963,N_30945,N_35898);
nor U43964 (N_43964,N_37323,N_34790);
xor U43965 (N_43965,N_31248,N_39618);
or U43966 (N_43966,N_31907,N_33081);
xnor U43967 (N_43967,N_37435,N_31115);
xnor U43968 (N_43968,N_38522,N_35742);
or U43969 (N_43969,N_31726,N_39482);
or U43970 (N_43970,N_35327,N_31696);
or U43971 (N_43971,N_36922,N_33317);
xnor U43972 (N_43972,N_31742,N_39947);
nand U43973 (N_43973,N_31261,N_32145);
nor U43974 (N_43974,N_38319,N_31569);
nor U43975 (N_43975,N_34888,N_37848);
and U43976 (N_43976,N_37966,N_32966);
xnor U43977 (N_43977,N_36101,N_31552);
nand U43978 (N_43978,N_35162,N_32005);
xor U43979 (N_43979,N_34022,N_32539);
xnor U43980 (N_43980,N_35561,N_30605);
or U43981 (N_43981,N_36483,N_35325);
xnor U43982 (N_43982,N_31022,N_31655);
xnor U43983 (N_43983,N_32034,N_35683);
or U43984 (N_43984,N_30775,N_35491);
xnor U43985 (N_43985,N_30090,N_31842);
xnor U43986 (N_43986,N_31646,N_35330);
and U43987 (N_43987,N_31698,N_32891);
xnor U43988 (N_43988,N_30522,N_38654);
or U43989 (N_43989,N_35197,N_35060);
xor U43990 (N_43990,N_33304,N_30446);
or U43991 (N_43991,N_33585,N_32656);
and U43992 (N_43992,N_35073,N_35071);
nand U43993 (N_43993,N_32809,N_39198);
xor U43994 (N_43994,N_34406,N_39982);
xor U43995 (N_43995,N_31397,N_35834);
xor U43996 (N_43996,N_35931,N_36962);
nand U43997 (N_43997,N_30004,N_33554);
xnor U43998 (N_43998,N_33714,N_38386);
and U43999 (N_43999,N_36073,N_31912);
or U44000 (N_44000,N_30661,N_38013);
or U44001 (N_44001,N_36366,N_35560);
xor U44002 (N_44002,N_37739,N_38600);
or U44003 (N_44003,N_30496,N_39855);
or U44004 (N_44004,N_38570,N_33442);
or U44005 (N_44005,N_38708,N_36486);
xnor U44006 (N_44006,N_38507,N_31603);
nor U44007 (N_44007,N_34422,N_35925);
xnor U44008 (N_44008,N_36164,N_39671);
or U44009 (N_44009,N_38412,N_31714);
xnor U44010 (N_44010,N_33390,N_31073);
or U44011 (N_44011,N_31598,N_37673);
or U44012 (N_44012,N_38001,N_33003);
or U44013 (N_44013,N_32914,N_33623);
nor U44014 (N_44014,N_39405,N_30180);
nand U44015 (N_44015,N_34128,N_39471);
nor U44016 (N_44016,N_35950,N_37315);
xor U44017 (N_44017,N_35928,N_36258);
xnor U44018 (N_44018,N_34263,N_33547);
nor U44019 (N_44019,N_36096,N_31175);
or U44020 (N_44020,N_33760,N_36087);
nor U44021 (N_44021,N_31881,N_31654);
nand U44022 (N_44022,N_32345,N_37404);
nor U44023 (N_44023,N_33705,N_34617);
nor U44024 (N_44024,N_33104,N_39975);
nor U44025 (N_44025,N_39674,N_37563);
and U44026 (N_44026,N_35672,N_35739);
and U44027 (N_44027,N_33786,N_34675);
nand U44028 (N_44028,N_36900,N_35098);
or U44029 (N_44029,N_34046,N_32509);
xor U44030 (N_44030,N_32286,N_39014);
nor U44031 (N_44031,N_39151,N_38251);
and U44032 (N_44032,N_33234,N_39514);
nand U44033 (N_44033,N_36387,N_39845);
nand U44034 (N_44034,N_36740,N_35522);
nand U44035 (N_44035,N_33202,N_32896);
nor U44036 (N_44036,N_39074,N_37331);
nor U44037 (N_44037,N_34578,N_32808);
and U44038 (N_44038,N_39498,N_35722);
or U44039 (N_44039,N_35303,N_33070);
nand U44040 (N_44040,N_37251,N_32429);
and U44041 (N_44041,N_30514,N_37747);
nand U44042 (N_44042,N_31300,N_31554);
or U44043 (N_44043,N_30310,N_39068);
xnor U44044 (N_44044,N_38729,N_31214);
or U44045 (N_44045,N_38271,N_36236);
or U44046 (N_44046,N_34918,N_32237);
nor U44047 (N_44047,N_34457,N_39934);
nand U44048 (N_44048,N_31315,N_31602);
and U44049 (N_44049,N_38810,N_33589);
xnor U44050 (N_44050,N_33494,N_37604);
xnor U44051 (N_44051,N_36790,N_39043);
nand U44052 (N_44052,N_37295,N_34868);
nand U44053 (N_44053,N_34338,N_39446);
and U44054 (N_44054,N_33948,N_38308);
and U44055 (N_44055,N_39931,N_30309);
xor U44056 (N_44056,N_32795,N_36510);
nor U44057 (N_44057,N_33185,N_37670);
and U44058 (N_44058,N_39634,N_38473);
nor U44059 (N_44059,N_35378,N_39834);
nor U44060 (N_44060,N_37713,N_31146);
and U44061 (N_44061,N_35622,N_32314);
nor U44062 (N_44062,N_30792,N_39440);
or U44063 (N_44063,N_33938,N_37618);
nand U44064 (N_44064,N_39268,N_37526);
xor U44065 (N_44065,N_38298,N_35114);
and U44066 (N_44066,N_34579,N_36256);
xnor U44067 (N_44067,N_30388,N_36033);
and U44068 (N_44068,N_30680,N_30851);
and U44069 (N_44069,N_34764,N_39415);
nand U44070 (N_44070,N_31129,N_31029);
nand U44071 (N_44071,N_38529,N_31241);
or U44072 (N_44072,N_37278,N_33050);
and U44073 (N_44073,N_37726,N_35282);
nand U44074 (N_44074,N_34534,N_31734);
or U44075 (N_44075,N_31711,N_32128);
and U44076 (N_44076,N_32742,N_30285);
nor U44077 (N_44077,N_33055,N_34993);
and U44078 (N_44078,N_39358,N_39071);
or U44079 (N_44079,N_32882,N_31638);
nor U44080 (N_44080,N_31491,N_31296);
nand U44081 (N_44081,N_32462,N_31631);
and U44082 (N_44082,N_38784,N_37721);
and U44083 (N_44083,N_34520,N_33091);
xor U44084 (N_44084,N_34794,N_35585);
or U44085 (N_44085,N_34254,N_31097);
and U44086 (N_44086,N_33422,N_36403);
nor U44087 (N_44087,N_31600,N_39762);
nand U44088 (N_44088,N_31918,N_31871);
and U44089 (N_44089,N_39943,N_38129);
or U44090 (N_44090,N_38413,N_33032);
nand U44091 (N_44091,N_32834,N_32484);
nor U44092 (N_44092,N_36966,N_35963);
and U44093 (N_44093,N_31916,N_31839);
or U44094 (N_44094,N_30210,N_30417);
xnor U44095 (N_44095,N_31761,N_38602);
nand U44096 (N_44096,N_39042,N_34911);
and U44097 (N_44097,N_39853,N_37841);
nor U44098 (N_44098,N_32129,N_32011);
xnor U44099 (N_44099,N_39103,N_31545);
and U44100 (N_44100,N_39965,N_33491);
nand U44101 (N_44101,N_31896,N_39236);
nor U44102 (N_44102,N_32933,N_39776);
and U44103 (N_44103,N_37796,N_35525);
xnor U44104 (N_44104,N_37197,N_30007);
nor U44105 (N_44105,N_31675,N_35024);
and U44106 (N_44106,N_32199,N_37986);
or U44107 (N_44107,N_38824,N_37353);
and U44108 (N_44108,N_36050,N_30320);
and U44109 (N_44109,N_31171,N_35943);
xnor U44110 (N_44110,N_34530,N_36995);
xnor U44111 (N_44111,N_33027,N_36456);
nor U44112 (N_44112,N_33906,N_30517);
xnor U44113 (N_44113,N_38635,N_33733);
nor U44114 (N_44114,N_30710,N_34973);
or U44115 (N_44115,N_35102,N_31259);
xnor U44116 (N_44116,N_33505,N_35996);
xor U44117 (N_44117,N_31256,N_33183);
nor U44118 (N_44118,N_31301,N_32846);
or U44119 (N_44119,N_34732,N_31383);
or U44120 (N_44120,N_34273,N_35809);
nand U44121 (N_44121,N_36513,N_38910);
and U44122 (N_44122,N_30864,N_31135);
or U44123 (N_44123,N_33346,N_32205);
nand U44124 (N_44124,N_32310,N_33915);
nand U44125 (N_44125,N_30995,N_33770);
xor U44126 (N_44126,N_36396,N_37021);
xor U44127 (N_44127,N_35532,N_35399);
or U44128 (N_44128,N_33788,N_38818);
and U44129 (N_44129,N_38723,N_36471);
xnor U44130 (N_44130,N_39326,N_38252);
nor U44131 (N_44131,N_30091,N_36226);
or U44132 (N_44132,N_32929,N_35659);
nand U44133 (N_44133,N_34449,N_34235);
nor U44134 (N_44134,N_30658,N_38674);
nor U44135 (N_44135,N_36596,N_31971);
xnor U44136 (N_44136,N_30648,N_38415);
and U44137 (N_44137,N_31957,N_31527);
nand U44138 (N_44138,N_35822,N_33555);
and U44139 (N_44139,N_31581,N_33609);
nand U44140 (N_44140,N_36257,N_32875);
nor U44141 (N_44141,N_31452,N_34845);
and U44142 (N_44142,N_36238,N_32965);
xor U44143 (N_44143,N_37374,N_39317);
and U44144 (N_44144,N_38912,N_34846);
xor U44145 (N_44145,N_32969,N_31691);
xor U44146 (N_44146,N_32208,N_36984);
and U44147 (N_44147,N_38393,N_37229);
and U44148 (N_44148,N_32045,N_33811);
xor U44149 (N_44149,N_34241,N_37223);
and U44150 (N_44150,N_35283,N_37017);
nor U44151 (N_44151,N_30931,N_35612);
nand U44152 (N_44152,N_32391,N_36332);
xnor U44153 (N_44153,N_35628,N_35775);
nor U44154 (N_44154,N_39716,N_33873);
and U44155 (N_44155,N_30326,N_30689);
nor U44156 (N_44156,N_32451,N_33117);
nor U44157 (N_44157,N_32061,N_37255);
and U44158 (N_44158,N_33591,N_33914);
and U44159 (N_44159,N_34309,N_30224);
and U44160 (N_44160,N_31281,N_39332);
nor U44161 (N_44161,N_30296,N_30716);
or U44162 (N_44162,N_36426,N_30231);
and U44163 (N_44163,N_35836,N_34646);
nand U44164 (N_44164,N_37387,N_30540);
nor U44165 (N_44165,N_37357,N_31798);
or U44166 (N_44166,N_33073,N_35708);
nand U44167 (N_44167,N_32222,N_30411);
or U44168 (N_44168,N_33294,N_39256);
nand U44169 (N_44169,N_38697,N_30567);
nor U44170 (N_44170,N_35101,N_34395);
nor U44171 (N_44171,N_39214,N_34952);
nand U44172 (N_44172,N_32486,N_37847);
xnor U44173 (N_44173,N_33391,N_32299);
or U44174 (N_44174,N_34459,N_35785);
and U44175 (N_44175,N_35625,N_39118);
nor U44176 (N_44176,N_32561,N_39171);
nand U44177 (N_44177,N_30597,N_39630);
nand U44178 (N_44178,N_31877,N_30158);
xor U44179 (N_44179,N_30693,N_32487);
nor U44180 (N_44180,N_38083,N_31368);
and U44181 (N_44181,N_36135,N_34702);
and U44182 (N_44182,N_37336,N_33767);
xor U44183 (N_44183,N_36591,N_37329);
nand U44184 (N_44184,N_37148,N_36670);
or U44185 (N_44185,N_32354,N_38822);
nand U44186 (N_44186,N_31189,N_32974);
xor U44187 (N_44187,N_39154,N_31251);
nor U44188 (N_44188,N_30259,N_35353);
and U44189 (N_44189,N_32236,N_31274);
or U44190 (N_44190,N_35422,N_37260);
or U44191 (N_44191,N_30796,N_33270);
xnor U44192 (N_44192,N_34167,N_37314);
nand U44193 (N_44193,N_30560,N_38683);
and U44194 (N_44194,N_34680,N_37720);
nor U44195 (N_44195,N_31963,N_36003);
nor U44196 (N_44196,N_39824,N_32442);
and U44197 (N_44197,N_35373,N_31400);
or U44198 (N_44198,N_31702,N_39509);
nor U44199 (N_44199,N_36284,N_37045);
nand U44200 (N_44200,N_35055,N_34933);
nor U44201 (N_44201,N_34947,N_37695);
or U44202 (N_44202,N_38284,N_37343);
or U44203 (N_44203,N_38659,N_35480);
or U44204 (N_44204,N_39403,N_30056);
xnor U44205 (N_44205,N_38462,N_33526);
xor U44206 (N_44206,N_30214,N_33340);
or U44207 (N_44207,N_32585,N_38422);
xnor U44208 (N_44208,N_34858,N_31890);
nor U44209 (N_44209,N_32445,N_38925);
xnor U44210 (N_44210,N_34626,N_37040);
xor U44211 (N_44211,N_30232,N_35661);
xnor U44212 (N_44212,N_32058,N_38056);
nor U44213 (N_44213,N_30225,N_35776);
xor U44214 (N_44214,N_35297,N_36980);
nand U44215 (N_44215,N_36276,N_30042);
nor U44216 (N_44216,N_31946,N_30844);
xor U44217 (N_44217,N_39215,N_34676);
nand U44218 (N_44218,N_30034,N_37500);
nor U44219 (N_44219,N_35322,N_32496);
and U44220 (N_44220,N_33541,N_32640);
nor U44221 (N_44221,N_32151,N_36214);
nor U44222 (N_44222,N_39738,N_32650);
and U44223 (N_44223,N_31133,N_32836);
nor U44224 (N_44224,N_31959,N_31679);
xor U44225 (N_44225,N_38617,N_31018);
xor U44226 (N_44226,N_34813,N_37967);
or U44227 (N_44227,N_35926,N_37411);
xnor U44228 (N_44228,N_33242,N_31154);
and U44229 (N_44229,N_36856,N_38389);
or U44230 (N_44230,N_32099,N_31443);
nand U44231 (N_44231,N_30010,N_37258);
and U44232 (N_44232,N_35818,N_33843);
xor U44233 (N_44233,N_34327,N_30432);
and U44234 (N_44234,N_34239,N_34276);
nor U44235 (N_44235,N_36001,N_30172);
nor U44236 (N_44236,N_32225,N_34839);
and U44237 (N_44237,N_39916,N_31317);
or U44238 (N_44238,N_35045,N_34364);
nor U44239 (N_44239,N_39134,N_37800);
xnor U44240 (N_44240,N_32184,N_30697);
and U44241 (N_44241,N_39238,N_35823);
or U44242 (N_44242,N_32149,N_34007);
xor U44243 (N_44243,N_35096,N_37952);
nor U44244 (N_44244,N_38499,N_33498);
nand U44245 (N_44245,N_36192,N_31670);
nand U44246 (N_44246,N_37810,N_36437);
xnor U44247 (N_44247,N_34486,N_37267);
nor U44248 (N_44248,N_32387,N_30656);
or U44249 (N_44249,N_33083,N_34033);
xnor U44250 (N_44250,N_36768,N_32962);
and U44251 (N_44251,N_38874,N_34206);
nand U44252 (N_44252,N_39519,N_39859);
or U44253 (N_44253,N_39203,N_32884);
xor U44254 (N_44254,N_36316,N_30852);
or U44255 (N_44255,N_38120,N_38755);
nor U44256 (N_44256,N_35584,N_37234);
nor U44257 (N_44257,N_38589,N_37436);
nand U44258 (N_44258,N_33833,N_36446);
nand U44259 (N_44259,N_34181,N_33114);
or U44260 (N_44260,N_32544,N_33353);
nand U44261 (N_44261,N_34630,N_31807);
xnor U44262 (N_44262,N_32921,N_30946);
xor U44263 (N_44263,N_38920,N_32233);
nor U44264 (N_44264,N_39839,N_30857);
xor U44265 (N_44265,N_33133,N_34180);
nand U44266 (N_44266,N_38888,N_32330);
and U44267 (N_44267,N_39489,N_36979);
nor U44268 (N_44268,N_38737,N_39274);
nor U44269 (N_44269,N_33131,N_31328);
or U44270 (N_44270,N_34249,N_36142);
and U44271 (N_44271,N_32347,N_31516);
xor U44272 (N_44272,N_39138,N_36475);
xor U44273 (N_44273,N_38188,N_32039);
nand U44274 (N_44274,N_30933,N_37481);
or U44275 (N_44275,N_31823,N_37611);
and U44276 (N_44276,N_33330,N_33443);
and U44277 (N_44277,N_37705,N_33999);
and U44278 (N_44278,N_32275,N_37437);
nand U44279 (N_44279,N_30741,N_39050);
nor U44280 (N_44280,N_37981,N_31737);
nand U44281 (N_44281,N_33174,N_33542);
or U44282 (N_44282,N_37701,N_36108);
xnor U44283 (N_44283,N_31212,N_35181);
nand U44284 (N_44284,N_37038,N_30711);
nand U44285 (N_44285,N_36727,N_37977);
nor U44286 (N_44286,N_32174,N_30355);
nand U44287 (N_44287,N_32646,N_38960);
nor U44288 (N_44288,N_30511,N_33892);
and U44289 (N_44289,N_30271,N_33940);
and U44290 (N_44290,N_38705,N_31044);
and U44291 (N_44291,N_33989,N_39533);
nor U44292 (N_44292,N_37903,N_34827);
xnor U44293 (N_44293,N_39139,N_33255);
xor U44294 (N_44294,N_36636,N_36823);
nor U44295 (N_44295,N_38235,N_39883);
nand U44296 (N_44296,N_31958,N_38175);
nor U44297 (N_44297,N_38099,N_33132);
nand U44298 (N_44298,N_32661,N_36286);
nor U44299 (N_44299,N_38172,N_36742);
or U44300 (N_44300,N_30819,N_37143);
xor U44301 (N_44301,N_35989,N_30587);
or U44302 (N_44302,N_36648,N_33460);
nand U44303 (N_44303,N_34966,N_39185);
and U44304 (N_44304,N_34028,N_37511);
and U44305 (N_44305,N_32863,N_33905);
nor U44306 (N_44306,N_32280,N_39984);
nor U44307 (N_44307,N_35033,N_35100);
nand U44308 (N_44308,N_33134,N_35495);
and U44309 (N_44309,N_32046,N_38799);
and U44310 (N_44310,N_36233,N_38908);
or U44311 (N_44311,N_36861,N_36036);
xnor U44312 (N_44312,N_33447,N_36249);
xnor U44313 (N_44313,N_36057,N_34986);
xnor U44314 (N_44314,N_37236,N_33208);
nor U44315 (N_44315,N_37818,N_32109);
xnor U44316 (N_44316,N_30590,N_32159);
nand U44317 (N_44317,N_38947,N_34411);
or U44318 (N_44318,N_39921,N_33808);
xnor U44319 (N_44319,N_31181,N_37037);
and U44320 (N_44320,N_30138,N_37875);
and U44321 (N_44321,N_37170,N_39515);
nor U44322 (N_44322,N_39516,N_37931);
and U44323 (N_44323,N_30832,N_33069);
xor U44324 (N_44324,N_34430,N_31771);
or U44325 (N_44325,N_32317,N_36502);
nand U44326 (N_44326,N_38276,N_38761);
xor U44327 (N_44327,N_37616,N_36539);
xor U44328 (N_44328,N_36961,N_32064);
xnor U44329 (N_44329,N_34050,N_39689);
nand U44330 (N_44330,N_31276,N_31930);
and U44331 (N_44331,N_37193,N_36941);
xnor U44332 (N_44332,N_39469,N_30665);
or U44333 (N_44333,N_39701,N_33953);
or U44334 (N_44334,N_37633,N_36208);
or U44335 (N_44335,N_32425,N_31517);
nor U44336 (N_44336,N_30117,N_32448);
nor U44337 (N_44337,N_33158,N_37338);
nor U44338 (N_44338,N_36895,N_32677);
xnor U44339 (N_44339,N_38439,N_37283);
or U44340 (N_44340,N_39306,N_39424);
xnor U44341 (N_44341,N_39632,N_38830);
nor U44342 (N_44342,N_31096,N_32435);
xor U44343 (N_44343,N_31327,N_31899);
and U44344 (N_44344,N_32954,N_30655);
or U44345 (N_44345,N_31565,N_37649);
nand U44346 (N_44346,N_37590,N_34931);
nand U44347 (N_44347,N_31299,N_31595);
xnor U44348 (N_44348,N_37459,N_33697);
nand U44349 (N_44349,N_36698,N_34198);
nor U44350 (N_44350,N_35939,N_37265);
nor U44351 (N_44351,N_36376,N_38669);
and U44352 (N_44352,N_32232,N_36082);
nand U44353 (N_44353,N_33332,N_39336);
xnor U44354 (N_44354,N_33189,N_39428);
and U44355 (N_44355,N_35308,N_35674);
xor U44356 (N_44356,N_33834,N_35549);
nor U44357 (N_44357,N_35804,N_32647);
nor U44358 (N_44358,N_34115,N_39486);
and U44359 (N_44359,N_30531,N_34025);
and U44360 (N_44360,N_39517,N_35155);
and U44361 (N_44361,N_35070,N_31031);
xnor U44362 (N_44362,N_33928,N_35180);
xor U44363 (N_44363,N_30262,N_33497);
and U44364 (N_44364,N_31498,N_37916);
xor U44365 (N_44365,N_36267,N_32492);
xor U44366 (N_44366,N_31668,N_31965);
xor U44367 (N_44367,N_39608,N_32960);
nand U44368 (N_44368,N_36926,N_30745);
or U44369 (N_44369,N_30204,N_36690);
xor U44370 (N_44370,N_31640,N_31013);
and U44371 (N_44371,N_37326,N_39341);
nand U44372 (N_44372,N_36423,N_30828);
or U44373 (N_44373,N_33379,N_36729);
nor U44374 (N_44374,N_38047,N_33706);
or U44375 (N_44375,N_37948,N_32580);
or U44376 (N_44376,N_36566,N_39736);
xnor U44377 (N_44377,N_38949,N_39005);
and U44378 (N_44378,N_33512,N_37172);
nand U44379 (N_44379,N_33979,N_30430);
and U44380 (N_44380,N_33947,N_33747);
xor U44381 (N_44381,N_34797,N_37527);
and U44382 (N_44382,N_38272,N_39168);
xnor U44383 (N_44383,N_36261,N_37723);
xnor U44384 (N_44384,N_35687,N_38101);
and U44385 (N_44385,N_32771,N_36803);
xnor U44386 (N_44386,N_30433,N_37806);
or U44387 (N_44387,N_32759,N_39107);
or U44388 (N_44388,N_30194,N_31230);
nand U44389 (N_44389,N_34190,N_37070);
xnor U44390 (N_44390,N_39104,N_35279);
and U44391 (N_44391,N_39202,N_37287);
nand U44392 (N_44392,N_34220,N_37622);
nor U44393 (N_44393,N_38140,N_38961);
nor U44394 (N_44394,N_34153,N_30086);
and U44395 (N_44395,N_33823,N_37656);
nand U44396 (N_44396,N_30399,N_31320);
xnor U44397 (N_44397,N_32256,N_33022);
nor U44398 (N_44398,N_34026,N_33282);
nor U44399 (N_44399,N_33789,N_30708);
xnor U44400 (N_44400,N_35292,N_36109);
nand U44401 (N_44401,N_32065,N_37477);
nand U44402 (N_44402,N_34349,N_30327);
nor U44403 (N_44403,N_34937,N_36285);
nand U44404 (N_44404,N_36869,N_35940);
xnor U44405 (N_44405,N_36105,N_38955);
and U44406 (N_44406,N_38091,N_31538);
nor U44407 (N_44407,N_33814,N_39426);
or U44408 (N_44408,N_32408,N_36577);
and U44409 (N_44409,N_38604,N_31158);
nor U44410 (N_44410,N_36874,N_39092);
xnor U44411 (N_44411,N_31923,N_31405);
nand U44412 (N_44412,N_30777,N_37844);
nor U44413 (N_44413,N_39441,N_33144);
xnor U44414 (N_44414,N_30849,N_37874);
and U44415 (N_44415,N_33824,N_33830);
or U44416 (N_44416,N_39780,N_34027);
nand U44417 (N_44417,N_33501,N_33537);
nor U44418 (N_44418,N_31205,N_34394);
nor U44419 (N_44419,N_32156,N_31995);
and U44420 (N_44420,N_39046,N_30182);
nand U44421 (N_44421,N_38686,N_37460);
xor U44422 (N_44422,N_36083,N_35762);
nand U44423 (N_44423,N_31246,N_32931);
xnor U44424 (N_44424,N_31389,N_38521);
nand U44425 (N_44425,N_32939,N_34325);
and U44426 (N_44426,N_34867,N_38195);
nor U44427 (N_44427,N_38688,N_37020);
nand U44428 (N_44428,N_33863,N_30347);
xnor U44429 (N_44429,N_32469,N_31162);
xor U44430 (N_44430,N_30678,N_34694);
nand U44431 (N_44431,N_38607,N_32269);
nor U44432 (N_44432,N_38060,N_33432);
and U44433 (N_44433,N_33987,N_32658);
or U44434 (N_44434,N_36203,N_35347);
nor U44435 (N_44435,N_35463,N_37926);
and U44436 (N_44436,N_39397,N_34731);
or U44437 (N_44437,N_30572,N_35740);
and U44438 (N_44438,N_30556,N_30650);
nand U44439 (N_44439,N_38081,N_37276);
or U44440 (N_44440,N_38225,N_31587);
nand U44441 (N_44441,N_33857,N_39396);
nor U44442 (N_44442,N_34506,N_35382);
nor U44443 (N_44443,N_34185,N_32513);
xor U44444 (N_44444,N_38933,N_39679);
and U44445 (N_44445,N_38978,N_36334);
nor U44446 (N_44446,N_36527,N_32083);
or U44447 (N_44447,N_37361,N_32630);
xnor U44448 (N_44448,N_30445,N_32161);
or U44449 (N_44449,N_32295,N_38749);
xnor U44450 (N_44450,N_39805,N_32390);
nor U44451 (N_44451,N_33424,N_35519);
or U44452 (N_44452,N_36288,N_38568);
nand U44453 (N_44453,N_32111,N_30337);
or U44454 (N_44454,N_30414,N_39758);
nand U44455 (N_44455,N_34643,N_32660);
or U44456 (N_44456,N_31416,N_38751);
nand U44457 (N_44457,N_31157,N_37955);
nand U44458 (N_44458,N_34266,N_35213);
and U44459 (N_44459,N_32031,N_37425);
nor U44460 (N_44460,N_37324,N_39303);
nor U44461 (N_44461,N_36157,N_39402);
nand U44462 (N_44462,N_30385,N_30935);
or U44463 (N_44463,N_38977,N_36424);
xor U44464 (N_44464,N_39963,N_34051);
xor U44465 (N_44465,N_39058,N_36482);
or U44466 (N_44466,N_36818,N_32124);
nand U44467 (N_44467,N_35384,N_32608);
and U44468 (N_44468,N_35040,N_38945);
xor U44469 (N_44469,N_30159,N_38485);
xor U44470 (N_44470,N_34606,N_33233);
or U44471 (N_44471,N_35194,N_38118);
nor U44472 (N_44472,N_36040,N_30623);
xor U44473 (N_44473,N_39497,N_34003);
and U44474 (N_44474,N_30519,N_37866);
nor U44475 (N_44475,N_34445,N_31719);
nand U44476 (N_44476,N_32274,N_31987);
and U44477 (N_44477,N_32603,N_31750);
or U44478 (N_44478,N_34998,N_38937);
nor U44479 (N_44479,N_34370,N_33097);
and U44480 (N_44480,N_34884,N_30731);
nand U44481 (N_44481,N_31593,N_36600);
or U44482 (N_44482,N_34976,N_39089);
and U44483 (N_44483,N_30353,N_36563);
xor U44484 (N_44484,N_38260,N_36859);
or U44485 (N_44485,N_37923,N_32069);
xor U44486 (N_44486,N_33445,N_32835);
xor U44487 (N_44487,N_38622,N_34707);
nand U44488 (N_44488,N_30641,N_33858);
xnor U44489 (N_44489,N_32389,N_33474);
nand U44490 (N_44490,N_35208,N_33192);
nor U44491 (N_44491,N_35087,N_34040);
nor U44492 (N_44492,N_35959,N_37362);
and U44493 (N_44493,N_39739,N_30961);
nand U44494 (N_44494,N_32241,N_34503);
xnor U44495 (N_44495,N_34210,N_32548);
nor U44496 (N_44496,N_33488,N_39054);
nor U44497 (N_44497,N_32673,N_35274);
nand U44498 (N_44498,N_31107,N_39385);
nor U44499 (N_44499,N_37359,N_30015);
xor U44500 (N_44500,N_33178,N_36585);
nand U44501 (N_44501,N_33044,N_33832);
or U44502 (N_44502,N_32094,N_38541);
or U44503 (N_44503,N_37635,N_37949);
nor U44504 (N_44504,N_34874,N_37522);
or U44505 (N_44505,N_38898,N_36619);
nand U44506 (N_44506,N_31804,N_32586);
nor U44507 (N_44507,N_33895,N_33917);
nor U44508 (N_44508,N_30077,N_32976);
xor U44509 (N_44509,N_35262,N_33695);
nor U44510 (N_44510,N_39914,N_36313);
or U44511 (N_44511,N_33215,N_38170);
nor U44512 (N_44512,N_32637,N_36360);
and U44513 (N_44513,N_35416,N_39972);
nor U44514 (N_44514,N_37760,N_33093);
or U44515 (N_44515,N_37636,N_39912);
and U44516 (N_44516,N_35479,N_37467);
and U44517 (N_44517,N_32964,N_32172);
xor U44518 (N_44518,N_32937,N_39667);
or U44519 (N_44519,N_33427,N_35603);
xnor U44520 (N_44520,N_34822,N_36228);
nand U44521 (N_44521,N_33343,N_30634);
nand U44522 (N_44522,N_35544,N_36700);
nor U44523 (N_44523,N_39021,N_34455);
or U44524 (N_44524,N_36062,N_38152);
nand U44525 (N_44525,N_33506,N_35933);
nor U44526 (N_44526,N_39392,N_38542);
xor U44527 (N_44527,N_30329,N_33275);
nand U44528 (N_44528,N_35513,N_36795);
nand U44529 (N_44529,N_37869,N_33484);
xnor U44530 (N_44530,N_33736,N_37566);
or U44531 (N_44531,N_36159,N_36448);
nor U44532 (N_44532,N_39075,N_30717);
nand U44533 (N_44533,N_33461,N_37019);
nor U44534 (N_44534,N_34576,N_31223);
nor U44535 (N_44535,N_39001,N_38395);
or U44536 (N_44536,N_34109,N_39801);
nor U44537 (N_44537,N_32386,N_32902);
nor U44538 (N_44538,N_35067,N_33919);
and U44539 (N_44539,N_35456,N_30078);
nor U44540 (N_44540,N_31283,N_31929);
and U44541 (N_44541,N_37262,N_30907);
and U44542 (N_44542,N_36365,N_38400);
and U44543 (N_44543,N_33084,N_33847);
or U44544 (N_44544,N_34372,N_33326);
and U44545 (N_44545,N_33212,N_36398);
or U44546 (N_44546,N_39850,N_36405);
xnor U44547 (N_44547,N_31583,N_30400);
or U44548 (N_44548,N_31292,N_35211);
nand U44549 (N_44549,N_38989,N_32746);
nand U44550 (N_44550,N_37553,N_34825);
xnor U44551 (N_44551,N_30472,N_37127);
xnor U44552 (N_44552,N_36144,N_36401);
or U44553 (N_44553,N_33291,N_36579);
and U44554 (N_44554,N_34887,N_38639);
and U44555 (N_44555,N_32404,N_30988);
nand U44556 (N_44556,N_30079,N_34157);
xnor U44557 (N_44557,N_32632,N_39915);
and U44558 (N_44558,N_31755,N_39978);
nand U44559 (N_44559,N_31858,N_35302);
nor U44560 (N_44560,N_30340,N_37557);
nand U44561 (N_44561,N_37456,N_30837);
or U44562 (N_44562,N_39884,N_38369);
xor U44563 (N_44563,N_33182,N_37210);
nor U44564 (N_44564,N_32943,N_38430);
or U44565 (N_44565,N_35144,N_39524);
nand U44566 (N_44566,N_37816,N_34042);
nor U44567 (N_44567,N_34240,N_36042);
nor U44568 (N_44568,N_38184,N_31644);
or U44569 (N_44569,N_35358,N_39015);
nand U44570 (N_44570,N_35133,N_38595);
and U44571 (N_44571,N_33396,N_37185);
nor U44572 (N_44572,N_36081,N_30797);
or U44573 (N_44573,N_38185,N_31381);
nor U44574 (N_44574,N_33063,N_31372);
and U44575 (N_44575,N_30251,N_36714);
and U44576 (N_44576,N_36607,N_36848);
xnor U44577 (N_44577,N_33281,N_34568);
or U44578 (N_44578,N_31359,N_34950);
nand U44579 (N_44579,N_32956,N_36858);
or U44580 (N_44580,N_36732,N_34583);
xor U44581 (N_44581,N_39196,N_35839);
or U44582 (N_44582,N_39251,N_35002);
nor U44583 (N_44583,N_35036,N_33139);
xor U44584 (N_44584,N_33430,N_32734);
nand U44585 (N_44585,N_31847,N_31451);
or U44586 (N_44586,N_36440,N_30274);
xnor U44587 (N_44587,N_33345,N_31821);
and U44588 (N_44588,N_38211,N_33428);
or U44589 (N_44589,N_39087,N_39413);
nand U44590 (N_44590,N_36692,N_33464);
nand U44591 (N_44591,N_32565,N_35276);
nand U44592 (N_44592,N_37149,N_30639);
nand U44593 (N_44593,N_30273,N_37152);
and U44594 (N_44594,N_35567,N_38569);
nand U44595 (N_44595,N_33476,N_34262);
or U44596 (N_44596,N_35904,N_38045);
nor U44597 (N_44597,N_30770,N_38379);
or U44598 (N_44598,N_34975,N_39792);
and U44599 (N_44599,N_30449,N_38343);
or U44600 (N_44600,N_38483,N_32556);
xnor U44601 (N_44601,N_30886,N_33262);
or U44602 (N_44602,N_32617,N_38351);
or U44603 (N_44603,N_37072,N_37097);
nand U44604 (N_44604,N_30598,N_32244);
nor U44605 (N_44605,N_32319,N_38434);
or U44606 (N_44606,N_31060,N_36664);
xor U44607 (N_44607,N_36807,N_33630);
xnor U44608 (N_44608,N_38985,N_30389);
xor U44609 (N_44609,N_32190,N_38125);
or U44610 (N_44610,N_34150,N_34555);
and U44611 (N_44611,N_36574,N_30910);
xnor U44612 (N_44612,N_37041,N_37548);
and U44613 (N_44613,N_38216,N_39357);
nor U44614 (N_44614,N_34865,N_38031);
and U44615 (N_44615,N_34852,N_37392);
and U44616 (N_44616,N_32350,N_37238);
xor U44617 (N_44617,N_33378,N_33720);
nand U44618 (N_44618,N_34350,N_39280);
nor U44619 (N_44619,N_35107,N_32597);
nand U44620 (N_44620,N_35698,N_34772);
nand U44621 (N_44621,N_38934,N_33821);
or U44622 (N_44622,N_38883,N_37174);
and U44623 (N_44623,N_31065,N_35954);
nor U44624 (N_44624,N_39808,N_38732);
and U44625 (N_44625,N_35484,N_36338);
nor U44626 (N_44626,N_36340,N_32480);
xnor U44627 (N_44627,N_38063,N_39287);
or U44628 (N_44628,N_30692,N_33147);
xor U44629 (N_44629,N_34716,N_38664);
xnor U44630 (N_44630,N_30696,N_31415);
or U44631 (N_44631,N_39518,N_33256);
and U44632 (N_44632,N_32711,N_33112);
xor U44633 (N_44633,N_37954,N_34804);
nor U44634 (N_44634,N_37471,N_30778);
nand U44635 (N_44635,N_33161,N_32421);
xor U44636 (N_44636,N_30493,N_36268);
xnor U44637 (N_44637,N_33150,N_31844);
and U44638 (N_44638,N_31221,N_36063);
and U44639 (N_44639,N_39540,N_39534);
nor U44640 (N_44640,N_30281,N_36546);
nand U44641 (N_44641,N_37052,N_35673);
and U44642 (N_44642,N_34258,N_36872);
and U44643 (N_44643,N_32619,N_39319);
nor U44644 (N_44644,N_31633,N_36053);
or U44645 (N_44645,N_31295,N_36381);
nand U44646 (N_44646,N_37395,N_30784);
or U44647 (N_44647,N_30350,N_33228);
nand U44648 (N_44648,N_38441,N_31454);
or U44649 (N_44649,N_35092,N_39368);
nand U44650 (N_44650,N_39977,N_38450);
nand U44651 (N_44651,N_39192,N_33452);
or U44652 (N_44652,N_35854,N_36344);
nor U44653 (N_44653,N_35700,N_34560);
nand U44654 (N_44654,N_37515,N_38452);
nand U44655 (N_44655,N_34673,N_38780);
or U44656 (N_44656,N_30874,N_38300);
xor U44657 (N_44657,N_38666,N_33007);
nor U44658 (N_44658,N_38227,N_35615);
nor U44659 (N_44659,N_31667,N_31355);
or U44660 (N_44660,N_37034,N_39970);
and U44661 (N_44661,N_39611,N_38375);
or U44662 (N_44662,N_39812,N_31237);
or U44663 (N_44663,N_34081,N_31815);
nand U44664 (N_44664,N_31269,N_36888);
and U44665 (N_44665,N_32772,N_31432);
and U44666 (N_44666,N_31879,N_31393);
xor U44667 (N_44667,N_36065,N_38274);
or U44668 (N_44668,N_30363,N_35652);
and U44669 (N_44669,N_38535,N_32240);
xor U44670 (N_44670,N_34179,N_33098);
nor U44671 (N_44671,N_37647,N_34286);
and U44672 (N_44672,N_39728,N_33076);
or U44673 (N_44673,N_34742,N_33513);
or U44674 (N_44674,N_34513,N_30841);
nor U44675 (N_44675,N_35685,N_35447);
nor U44676 (N_44676,N_35510,N_38405);
nor U44677 (N_44677,N_33904,N_30913);
nor U44678 (N_44678,N_31672,N_31660);
xor U44679 (N_44679,N_32689,N_31331);
and U44680 (N_44680,N_39036,N_39360);
nor U44681 (N_44681,N_39394,N_36477);
nor U44682 (N_44682,N_31621,N_36182);
or U44683 (N_44683,N_31293,N_33126);
or U44684 (N_44684,N_38839,N_31192);
nand U44685 (N_44685,N_31455,N_35787);
or U44686 (N_44686,N_39974,N_32503);
nand U44687 (N_44687,N_33296,N_36723);
xor U44688 (N_44688,N_36224,N_32385);
xnor U44689 (N_44689,N_36540,N_35497);
and U44690 (N_44690,N_33538,N_33558);
or U44691 (N_44691,N_38696,N_37100);
or U44692 (N_44692,N_37988,N_35267);
nand U44693 (N_44693,N_36251,N_31379);
nand U44694 (N_44694,N_38355,N_32195);
xnor U44695 (N_44695,N_34294,N_34916);
xor U44696 (N_44696,N_38094,N_35159);
or U44697 (N_44697,N_33524,N_39331);
and U44698 (N_44698,N_33135,N_34616);
xnor U44699 (N_44699,N_32035,N_34687);
or U44700 (N_44700,N_33894,N_31883);
nand U44701 (N_44701,N_35467,N_35558);
or U44702 (N_44702,N_30427,N_33964);
xor U44703 (N_44703,N_32170,N_30267);
or U44704 (N_44704,N_36129,N_32168);
nand U44705 (N_44705,N_37567,N_36555);
and U44706 (N_44706,N_33087,N_38929);
nand U44707 (N_44707,N_31570,N_38494);
xor U44708 (N_44708,N_36838,N_36064);
xnor U44709 (N_44709,N_36462,N_35459);
nand U44710 (N_44710,N_30883,N_33810);
and U44711 (N_44711,N_39158,N_31519);
nand U44712 (N_44712,N_35432,N_33413);
or U44713 (N_44713,N_38484,N_37022);
nand U44714 (N_44714,N_37840,N_34298);
nand U44715 (N_44715,N_33151,N_39410);
nor U44716 (N_44716,N_35900,N_34971);
or U44717 (N_44717,N_36039,N_33666);
nor U44718 (N_44718,N_30035,N_32602);
nand U44719 (N_44719,N_31280,N_34664);
nand U44720 (N_44720,N_36350,N_32708);
and U44721 (N_44721,N_34634,N_36394);
nand U44722 (N_44722,N_37285,N_38150);
nor U44723 (N_44723,N_30100,N_34196);
or U44724 (N_44724,N_31626,N_38823);
and U44725 (N_44725,N_38974,N_35407);
nor U44726 (N_44726,N_32471,N_39329);
xnor U44727 (N_44727,N_35338,N_32125);
or U44728 (N_44728,N_38220,N_33869);
or U44729 (N_44729,N_31746,N_38950);
nor U44730 (N_44730,N_32790,N_39772);
nor U44731 (N_44731,N_31872,N_39382);
nand U44732 (N_44732,N_38525,N_35838);
xor U44733 (N_44733,N_32439,N_30584);
or U44734 (N_44734,N_32606,N_30357);
and U44735 (N_44735,N_33136,N_30644);
or U44736 (N_44736,N_37202,N_38956);
and U44737 (N_44737,N_30604,N_31919);
xnor U44738 (N_44738,N_34209,N_36357);
nor U44739 (N_44739,N_37824,N_33608);
or U44740 (N_44740,N_33753,N_33773);
nand U44741 (N_44741,N_36008,N_36615);
nand U44742 (N_44742,N_36383,N_31870);
xor U44743 (N_44743,N_30401,N_32735);
or U44744 (N_44744,N_34217,N_38805);
nor U44745 (N_44745,N_30264,N_37531);
xor U44746 (N_44746,N_30938,N_36857);
nor U44747 (N_44747,N_34508,N_36179);
nor U44748 (N_44748,N_37422,N_35129);
and U44749 (N_44749,N_31944,N_30742);
and U44750 (N_44750,N_35134,N_34037);
xnor U44751 (N_44751,N_38217,N_30393);
xor U44752 (N_44752,N_37795,N_37078);
xor U44753 (N_44753,N_33615,N_32870);
or U44754 (N_44754,N_37973,N_36694);
nand U44755 (N_44755,N_39529,N_30782);
xor U44756 (N_44756,N_35296,N_30760);
xnor U44757 (N_44757,N_32238,N_30062);
nor U44758 (N_44758,N_30683,N_30088);
nand U44759 (N_44759,N_33593,N_35909);
or U44760 (N_44760,N_31983,N_39248);
xor U44761 (N_44761,N_37119,N_36453);
or U44762 (N_44762,N_30421,N_36395);
nor U44763 (N_44763,N_36047,N_34121);
nand U44764 (N_44764,N_37053,N_32692);
nor U44765 (N_44765,N_31856,N_30498);
xor U44766 (N_44766,N_39868,N_37352);
xnor U44767 (N_44767,N_33385,N_33175);
and U44768 (N_44768,N_38601,N_38106);
nor U44769 (N_44769,N_30973,N_34602);
nor U44770 (N_44770,N_34605,N_30303);
nand U44771 (N_44771,N_39060,N_34482);
and U44772 (N_44772,N_35369,N_39650);
or U44773 (N_44773,N_38022,N_38744);
xor U44774 (N_44774,N_39581,N_39364);
or U44775 (N_44775,N_36697,N_33676);
xnor U44776 (N_44776,N_35050,N_32796);
and U44777 (N_44777,N_34464,N_35916);
and U44778 (N_44778,N_39654,N_37737);
and U44779 (N_44779,N_38567,N_33316);
nand U44780 (N_44780,N_36943,N_36266);
or U44781 (N_44781,N_34431,N_30687);
nand U44782 (N_44782,N_39490,N_32010);
nor U44783 (N_44783,N_30824,N_38421);
xor U44784 (N_44784,N_38896,N_32401);
xor U44785 (N_44785,N_38553,N_36178);
nor U44786 (N_44786,N_33861,N_35935);
xnor U44787 (N_44787,N_34850,N_34429);
xor U44788 (N_44788,N_39759,N_37940);
xnor U44789 (N_44789,N_38878,N_34399);
nand U44790 (N_44790,N_30198,N_30127);
nand U44791 (N_44791,N_36899,N_38815);
xor U44792 (N_44792,N_34044,N_31058);
and U44793 (N_44793,N_39715,N_30771);
xnor U44794 (N_44794,N_33973,N_35842);
or U44795 (N_44795,N_35574,N_30425);
or U44796 (N_44796,N_38963,N_35326);
xor U44797 (N_44797,N_34932,N_35805);
and U44798 (N_44798,N_34905,N_30979);
nand U44799 (N_44799,N_32395,N_30734);
and U44800 (N_44800,N_37356,N_39669);
and U44801 (N_44801,N_33493,N_37741);
xor U44802 (N_44802,N_30581,N_38885);
and U44803 (N_44803,N_34941,N_32538);
nor U44804 (N_44804,N_35617,N_39629);
xnor U44805 (N_44805,N_34659,N_30321);
or U44806 (N_44806,N_30635,N_37263);
xor U44807 (N_44807,N_36304,N_37582);
nor U44808 (N_44808,N_37365,N_30125);
xnor U44809 (N_44809,N_35029,N_30456);
and U44810 (N_44810,N_32987,N_39431);
nor U44811 (N_44811,N_34091,N_38773);
or U44812 (N_44812,N_35850,N_39576);
or U44813 (N_44813,N_37256,N_36798);
or U44814 (N_44814,N_35443,N_38826);
nor U44815 (N_44815,N_32837,N_39150);
xor U44816 (N_44816,N_34597,N_37298);
or U44817 (N_44817,N_30352,N_37291);
nor U44818 (N_44818,N_30265,N_30659);
and U44819 (N_44819,N_32373,N_31425);
and U44820 (N_44820,N_37665,N_33285);
nand U44821 (N_44821,N_36485,N_31797);
or U44822 (N_44822,N_39550,N_35579);
and U44823 (N_44823,N_38676,N_39461);
nand U44824 (N_44824,N_32980,N_30244);
nor U44825 (N_44825,N_35666,N_37742);
nand U44826 (N_44826,N_36678,N_37449);
nand U44827 (N_44827,N_31774,N_34608);
nand U44828 (N_44828,N_37542,N_36415);
xor U44829 (N_44829,N_36193,N_36901);
xnor U44830 (N_44830,N_36127,N_30269);
and U44831 (N_44831,N_37420,N_35923);
or U44832 (N_44832,N_39031,N_37216);
xnor U44833 (N_44833,N_32996,N_30628);
nand U44834 (N_44834,N_30985,N_30654);
xor U44835 (N_44835,N_38973,N_33916);
nor U44836 (N_44836,N_39572,N_39937);
and U44837 (N_44837,N_32489,N_37873);
nand U44838 (N_44838,N_39786,N_36891);
nand U44839 (N_44839,N_31941,N_32895);
xor U44840 (N_44840,N_32167,N_31867);
xnor U44841 (N_44841,N_39957,N_38454);
and U44842 (N_44842,N_34922,N_39864);
and U44843 (N_44843,N_38451,N_30160);
nor U44844 (N_44844,N_32631,N_35949);
nor U44845 (N_44845,N_37071,N_32185);
or U44846 (N_44846,N_34895,N_39767);
or U44847 (N_44847,N_30806,N_34138);
or U44848 (N_44848,N_33532,N_39038);
nor U44849 (N_44849,N_38027,N_30036);
nand U44850 (N_44850,N_37762,N_33106);
nor U44851 (N_44851,N_37843,N_31868);
nand U44852 (N_44852,N_35562,N_37664);
or U44853 (N_44853,N_34821,N_38900);
nor U44854 (N_44854,N_37894,N_35885);
nor U44855 (N_44855,N_31713,N_39393);
and U44856 (N_44856,N_34102,N_35506);
nand U44857 (N_44857,N_35478,N_34316);
and U44858 (N_44858,N_39537,N_35751);
nor U44859 (N_44859,N_37453,N_33342);
or U44860 (N_44860,N_35299,N_36715);
xnor U44861 (N_44861,N_38301,N_32176);
or U44862 (N_44862,N_39488,N_34036);
or U44863 (N_44863,N_38446,N_33023);
xnor U44864 (N_44864,N_36260,N_36447);
or U44865 (N_44865,N_38333,N_35110);
nand U44866 (N_44866,N_31347,N_36133);
xor U44867 (N_44867,N_37865,N_36972);
nor U44868 (N_44868,N_36957,N_33336);
or U44869 (N_44869,N_39146,N_36904);
or U44870 (N_44870,N_33807,N_31156);
xor U44871 (N_44871,N_30431,N_36639);
xnor U44872 (N_44872,N_31547,N_31613);
nor U44873 (N_44873,N_37247,N_30351);
xnor U44874 (N_44874,N_32316,N_35235);
and U44875 (N_44875,N_32296,N_30044);
nand U44876 (N_44876,N_32958,N_34533);
and U44877 (N_44877,N_38893,N_37585);
and U44878 (N_44878,N_37885,N_33988);
or U44879 (N_44879,N_30061,N_37738);
nand U44880 (N_44880,N_37703,N_33550);
or U44881 (N_44881,N_37450,N_38848);
or U44882 (N_44882,N_33153,N_34272);
nand U44883 (N_44883,N_34682,N_39856);
nor U44884 (N_44884,N_37575,N_39226);
xnor U44885 (N_44885,N_31404,N_36738);
xnor U44886 (N_44886,N_31387,N_31064);
or U44887 (N_44887,N_35572,N_34785);
nand U44888 (N_44888,N_34340,N_37536);
and U44889 (N_44889,N_36912,N_37999);
or U44890 (N_44890,N_33587,N_32957);
xor U44891 (N_44891,N_33024,N_35324);
xor U44892 (N_44892,N_32871,N_32498);
xnor U44893 (N_44893,N_33503,N_31341);
nand U44894 (N_44894,N_34302,N_37289);
xor U44895 (N_44895,N_38645,N_31666);
xor U44896 (N_44896,N_37184,N_35108);
nand U44897 (N_44897,N_37591,N_30990);
and U44898 (N_44898,N_36275,N_30006);
nand U44899 (N_44899,N_35440,N_33660);
or U44900 (N_44900,N_35696,N_36751);
or U44901 (N_44901,N_37051,N_37259);
and U44902 (N_44902,N_37452,N_36679);
nand U44903 (N_44903,N_35693,N_31004);
xor U44904 (N_44904,N_31474,N_33065);
nor U44905 (N_44905,N_35082,N_35031);
or U44906 (N_44906,N_39677,N_32358);
xor U44907 (N_44907,N_36554,N_30602);
nor U44908 (N_44908,N_32717,N_36355);
nand U44909 (N_44909,N_35857,N_32116);
nor U44910 (N_44910,N_39841,N_34633);
and U44911 (N_44911,N_34698,N_34642);
nor U44912 (N_44912,N_39436,N_31630);
nand U44913 (N_44913,N_34283,N_36616);
nor U44914 (N_44914,N_39204,N_37896);
xnor U44915 (N_44915,N_39793,N_30136);
xnor U44916 (N_44916,N_32012,N_38275);
xor U44917 (N_44917,N_39605,N_36495);
and U44918 (N_44918,N_35056,N_36618);
nand U44919 (N_44919,N_34552,N_37648);
xnor U44920 (N_44920,N_35212,N_33828);
or U44921 (N_44921,N_33107,N_33647);
nand U44922 (N_44922,N_36459,N_37934);
and U44923 (N_44923,N_39234,N_31190);
nor U44924 (N_44924,N_34900,N_38750);
nand U44925 (N_44925,N_31101,N_35313);
xor U44926 (N_44926,N_33921,N_38039);
nand U44927 (N_44927,N_38372,N_39409);
or U44928 (N_44928,N_33668,N_36139);
xor U44929 (N_44929,N_34018,N_34252);
xor U44930 (N_44930,N_33038,N_35594);
nand U44931 (N_44931,N_31284,N_36254);
and U44932 (N_44932,N_39077,N_39323);
xnor U44933 (N_44933,N_36882,N_38782);
xnor U44934 (N_44934,N_35643,N_34980);
nor U44935 (N_44935,N_36494,N_31494);
nand U44936 (N_44936,N_37472,N_30284);
and U44937 (N_44937,N_32112,N_34405);
nor U44938 (N_44938,N_39708,N_31275);
nand U44939 (N_44939,N_30861,N_34981);
nand U44940 (N_44940,N_31917,N_30750);
nor U44941 (N_44941,N_31616,N_32246);
xor U44942 (N_44942,N_35833,N_31098);
and U44943 (N_44943,N_34055,N_36589);
and U44944 (N_44944,N_33739,N_36419);
nor U44945 (N_44945,N_33708,N_34417);
or U44946 (N_44946,N_30181,N_37683);
xnor U44947 (N_44947,N_36850,N_36638);
nor U44948 (N_44948,N_37328,N_31835);
nand U44949 (N_44949,N_33026,N_32839);
and U44950 (N_44950,N_37886,N_36117);
nor U44951 (N_44951,N_35608,N_34776);
nand U44952 (N_44952,N_33756,N_33229);
xnor U44953 (N_44953,N_39470,N_34348);
xnor U44954 (N_44954,N_33140,N_35817);
or U44955 (N_44955,N_32558,N_38577);
xor U44956 (N_44956,N_31697,N_32727);
xnor U44957 (N_44957,N_32744,N_36744);
or U44958 (N_44958,N_31938,N_35410);
or U44959 (N_44959,N_31521,N_38201);
nor U44960 (N_44960,N_39592,N_38467);
and U44961 (N_44961,N_35712,N_33673);
nor U44962 (N_44962,N_31980,N_33709);
nand U44963 (N_44963,N_31233,N_39910);
nor U44964 (N_44964,N_36782,N_36156);
and U44965 (N_44965,N_30107,N_35730);
xnor U44966 (N_44966,N_35768,N_30307);
xnor U44967 (N_44967,N_37087,N_33523);
and U44968 (N_44968,N_39258,N_38624);
or U44969 (N_44969,N_39127,N_31145);
nand U44970 (N_44970,N_38714,N_36531);
and U44971 (N_44971,N_32056,N_39638);
nand U44972 (N_44972,N_36011,N_36940);
or U44973 (N_44973,N_33565,N_38808);
or U44974 (N_44974,N_33077,N_34485);
nor U44975 (N_44975,N_32955,N_34855);
nand U44976 (N_44976,N_33757,N_38069);
or U44977 (N_44977,N_35977,N_36309);
nor U44978 (N_44978,N_33197,N_31207);
xnor U44979 (N_44979,N_39180,N_39983);
or U44980 (N_44980,N_32091,N_35543);
and U44981 (N_44981,N_33455,N_39878);
nor U44982 (N_44982,N_35948,N_30991);
nand U44983 (N_44983,N_36497,N_39993);
nand U44984 (N_44984,N_35967,N_36930);
nand U44985 (N_44985,N_32097,N_32506);
or U44986 (N_44986,N_32860,N_39990);
and U44987 (N_44987,N_36989,N_33040);
xor U44988 (N_44988,N_34913,N_34812);
and U44989 (N_44989,N_39595,N_31460);
and U44990 (N_44990,N_33249,N_31855);
or U44991 (N_44991,N_37199,N_32999);
and U44992 (N_44992,N_35018,N_38807);
or U44993 (N_44993,N_38079,N_30137);
nor U44994 (N_44994,N_34835,N_33581);
and U44995 (N_44995,N_34573,N_37203);
xor U44996 (N_44996,N_34292,N_35188);
nor U44997 (N_44997,N_33013,N_39351);
and U44998 (N_44998,N_31217,N_31693);
nor U44999 (N_44999,N_35366,N_33331);
and U45000 (N_45000,N_34509,N_30621);
xnor U45001 (N_45001,N_31257,N_39281);
xnor U45002 (N_45002,N_30633,N_35366);
xor U45003 (N_45003,N_36714,N_30773);
nand U45004 (N_45004,N_31734,N_38974);
xnor U45005 (N_45005,N_35990,N_32128);
nand U45006 (N_45006,N_33084,N_35384);
nor U45007 (N_45007,N_34965,N_30257);
nor U45008 (N_45008,N_39134,N_38621);
nor U45009 (N_45009,N_34048,N_39181);
or U45010 (N_45010,N_36249,N_35935);
and U45011 (N_45011,N_36691,N_38568);
nand U45012 (N_45012,N_34910,N_39798);
xnor U45013 (N_45013,N_31274,N_35941);
nand U45014 (N_45014,N_31417,N_34309);
and U45015 (N_45015,N_33263,N_35529);
xor U45016 (N_45016,N_38780,N_39686);
nand U45017 (N_45017,N_35300,N_31755);
and U45018 (N_45018,N_36027,N_31244);
xor U45019 (N_45019,N_38595,N_32445);
nand U45020 (N_45020,N_34694,N_30455);
nand U45021 (N_45021,N_31954,N_39339);
or U45022 (N_45022,N_37901,N_33552);
nor U45023 (N_45023,N_36135,N_33805);
xor U45024 (N_45024,N_30441,N_36029);
and U45025 (N_45025,N_31103,N_30847);
xnor U45026 (N_45026,N_35879,N_35963);
or U45027 (N_45027,N_31404,N_38722);
nand U45028 (N_45028,N_30890,N_32291);
xnor U45029 (N_45029,N_32574,N_30156);
nor U45030 (N_45030,N_34132,N_38443);
or U45031 (N_45031,N_39318,N_34349);
nand U45032 (N_45032,N_31045,N_37961);
nor U45033 (N_45033,N_38370,N_37052);
or U45034 (N_45034,N_39657,N_30331);
nor U45035 (N_45035,N_30327,N_32473);
nand U45036 (N_45036,N_31724,N_34939);
xnor U45037 (N_45037,N_33730,N_33937);
nor U45038 (N_45038,N_39411,N_33657);
nand U45039 (N_45039,N_36936,N_36939);
nand U45040 (N_45040,N_39506,N_39089);
nor U45041 (N_45041,N_35130,N_39207);
nor U45042 (N_45042,N_31924,N_36531);
or U45043 (N_45043,N_32776,N_39201);
nor U45044 (N_45044,N_39488,N_32237);
nand U45045 (N_45045,N_33291,N_36527);
xor U45046 (N_45046,N_37561,N_33523);
xnor U45047 (N_45047,N_37721,N_38505);
nand U45048 (N_45048,N_38990,N_33406);
xor U45049 (N_45049,N_39654,N_34123);
nor U45050 (N_45050,N_35573,N_37228);
or U45051 (N_45051,N_36482,N_38688);
or U45052 (N_45052,N_34194,N_37403);
or U45053 (N_45053,N_38708,N_30202);
nor U45054 (N_45054,N_39579,N_38462);
or U45055 (N_45055,N_32534,N_37212);
and U45056 (N_45056,N_37566,N_38232);
and U45057 (N_45057,N_34427,N_31271);
or U45058 (N_45058,N_32579,N_32603);
nand U45059 (N_45059,N_31734,N_31583);
or U45060 (N_45060,N_36455,N_33148);
and U45061 (N_45061,N_39925,N_35238);
or U45062 (N_45062,N_32182,N_37352);
xnor U45063 (N_45063,N_33419,N_34026);
and U45064 (N_45064,N_33961,N_36217);
nor U45065 (N_45065,N_32558,N_34674);
nand U45066 (N_45066,N_37046,N_37055);
nor U45067 (N_45067,N_38531,N_34949);
or U45068 (N_45068,N_32372,N_30281);
and U45069 (N_45069,N_36084,N_33075);
and U45070 (N_45070,N_34128,N_30914);
nand U45071 (N_45071,N_37667,N_38087);
and U45072 (N_45072,N_35596,N_32670);
and U45073 (N_45073,N_38941,N_39081);
nand U45074 (N_45074,N_35396,N_34832);
nor U45075 (N_45075,N_34331,N_37143);
or U45076 (N_45076,N_37115,N_33415);
and U45077 (N_45077,N_34878,N_35589);
and U45078 (N_45078,N_39203,N_38166);
nor U45079 (N_45079,N_32449,N_35440);
and U45080 (N_45080,N_34508,N_37732);
and U45081 (N_45081,N_34562,N_34969);
nor U45082 (N_45082,N_31383,N_39696);
or U45083 (N_45083,N_35200,N_33962);
or U45084 (N_45084,N_35512,N_36433);
xor U45085 (N_45085,N_36978,N_37893);
or U45086 (N_45086,N_31116,N_38532);
or U45087 (N_45087,N_39431,N_38407);
xor U45088 (N_45088,N_35299,N_30871);
or U45089 (N_45089,N_30055,N_33378);
and U45090 (N_45090,N_31275,N_35301);
and U45091 (N_45091,N_38129,N_33564);
nor U45092 (N_45092,N_30759,N_36318);
nor U45093 (N_45093,N_37811,N_39502);
or U45094 (N_45094,N_34162,N_38355);
or U45095 (N_45095,N_35662,N_30932);
nand U45096 (N_45096,N_35338,N_34324);
or U45097 (N_45097,N_31060,N_38832);
or U45098 (N_45098,N_36983,N_35999);
nand U45099 (N_45099,N_37638,N_35693);
and U45100 (N_45100,N_32229,N_32355);
nand U45101 (N_45101,N_32183,N_34360);
nor U45102 (N_45102,N_31464,N_34283);
nor U45103 (N_45103,N_37702,N_35581);
xnor U45104 (N_45104,N_34463,N_36957);
or U45105 (N_45105,N_33989,N_37779);
nand U45106 (N_45106,N_34468,N_32338);
xnor U45107 (N_45107,N_31668,N_37545);
xor U45108 (N_45108,N_34362,N_31263);
nand U45109 (N_45109,N_33144,N_39427);
or U45110 (N_45110,N_32485,N_32931);
or U45111 (N_45111,N_30542,N_36575);
nor U45112 (N_45112,N_31362,N_34623);
nand U45113 (N_45113,N_39388,N_30690);
xnor U45114 (N_45114,N_39437,N_34067);
nor U45115 (N_45115,N_30145,N_39441);
and U45116 (N_45116,N_31666,N_31966);
nor U45117 (N_45117,N_39286,N_38293);
and U45118 (N_45118,N_30543,N_34934);
or U45119 (N_45119,N_34530,N_36848);
and U45120 (N_45120,N_32984,N_35208);
nor U45121 (N_45121,N_36089,N_37590);
and U45122 (N_45122,N_31493,N_30034);
and U45123 (N_45123,N_34752,N_35825);
xnor U45124 (N_45124,N_35096,N_32694);
or U45125 (N_45125,N_31681,N_30085);
nor U45126 (N_45126,N_37596,N_38344);
or U45127 (N_45127,N_35229,N_31037);
nor U45128 (N_45128,N_38547,N_35607);
or U45129 (N_45129,N_38321,N_33508);
nand U45130 (N_45130,N_34620,N_34251);
nand U45131 (N_45131,N_38090,N_39226);
xnor U45132 (N_45132,N_35762,N_32996);
nand U45133 (N_45133,N_36978,N_35564);
and U45134 (N_45134,N_34712,N_35322);
nand U45135 (N_45135,N_35621,N_35077);
or U45136 (N_45136,N_39894,N_31257);
xnor U45137 (N_45137,N_38867,N_33520);
or U45138 (N_45138,N_33637,N_37292);
nor U45139 (N_45139,N_39531,N_31339);
and U45140 (N_45140,N_32762,N_34113);
nor U45141 (N_45141,N_30871,N_39502);
or U45142 (N_45142,N_38223,N_32108);
xor U45143 (N_45143,N_30755,N_31687);
nor U45144 (N_45144,N_39639,N_38725);
nand U45145 (N_45145,N_30853,N_32921);
nand U45146 (N_45146,N_36488,N_32616);
and U45147 (N_45147,N_32942,N_33555);
and U45148 (N_45148,N_32180,N_31708);
or U45149 (N_45149,N_30318,N_35464);
nand U45150 (N_45150,N_39875,N_31227);
xor U45151 (N_45151,N_30652,N_31485);
nor U45152 (N_45152,N_36251,N_36828);
nand U45153 (N_45153,N_38773,N_35294);
and U45154 (N_45154,N_37170,N_34779);
and U45155 (N_45155,N_39003,N_36346);
nand U45156 (N_45156,N_39635,N_37842);
nand U45157 (N_45157,N_33105,N_37883);
or U45158 (N_45158,N_32183,N_38214);
nand U45159 (N_45159,N_30072,N_31489);
nand U45160 (N_45160,N_30670,N_32276);
nor U45161 (N_45161,N_35467,N_38968);
xnor U45162 (N_45162,N_36596,N_33205);
nand U45163 (N_45163,N_39375,N_38974);
nand U45164 (N_45164,N_39584,N_38198);
nand U45165 (N_45165,N_34283,N_38557);
and U45166 (N_45166,N_32154,N_37528);
nand U45167 (N_45167,N_38661,N_32535);
xnor U45168 (N_45168,N_35142,N_32573);
nor U45169 (N_45169,N_37705,N_31578);
nor U45170 (N_45170,N_36709,N_32247);
or U45171 (N_45171,N_34141,N_33998);
or U45172 (N_45172,N_32547,N_39031);
xnor U45173 (N_45173,N_33348,N_30597);
xor U45174 (N_45174,N_34020,N_39583);
xor U45175 (N_45175,N_36403,N_36728);
nor U45176 (N_45176,N_34267,N_35984);
or U45177 (N_45177,N_32964,N_34199);
nand U45178 (N_45178,N_33433,N_37469);
nand U45179 (N_45179,N_30931,N_35938);
nor U45180 (N_45180,N_36521,N_37064);
xnor U45181 (N_45181,N_33623,N_35433);
xor U45182 (N_45182,N_32775,N_32406);
nand U45183 (N_45183,N_39673,N_31610);
nand U45184 (N_45184,N_35368,N_34017);
and U45185 (N_45185,N_38886,N_36721);
xor U45186 (N_45186,N_38283,N_38396);
or U45187 (N_45187,N_39500,N_36633);
or U45188 (N_45188,N_36151,N_36087);
or U45189 (N_45189,N_33511,N_37553);
and U45190 (N_45190,N_30429,N_37926);
nand U45191 (N_45191,N_30712,N_36264);
nor U45192 (N_45192,N_30347,N_33221);
nor U45193 (N_45193,N_33927,N_34187);
nand U45194 (N_45194,N_32368,N_31769);
nand U45195 (N_45195,N_37550,N_32567);
xor U45196 (N_45196,N_37546,N_33092);
xnor U45197 (N_45197,N_30080,N_33816);
nor U45198 (N_45198,N_31263,N_39855);
and U45199 (N_45199,N_37539,N_33144);
nor U45200 (N_45200,N_33485,N_30665);
or U45201 (N_45201,N_34503,N_38248);
or U45202 (N_45202,N_36382,N_39561);
nand U45203 (N_45203,N_39142,N_32943);
and U45204 (N_45204,N_35851,N_35561);
or U45205 (N_45205,N_32313,N_31883);
nor U45206 (N_45206,N_39332,N_34206);
nor U45207 (N_45207,N_30332,N_30283);
xor U45208 (N_45208,N_30299,N_36674);
xnor U45209 (N_45209,N_39830,N_32591);
or U45210 (N_45210,N_33898,N_32413);
xor U45211 (N_45211,N_33809,N_32003);
nand U45212 (N_45212,N_33801,N_32319);
xnor U45213 (N_45213,N_32680,N_30011);
xnor U45214 (N_45214,N_33069,N_36000);
nand U45215 (N_45215,N_36202,N_36511);
or U45216 (N_45216,N_36156,N_33209);
or U45217 (N_45217,N_34348,N_36176);
xnor U45218 (N_45218,N_32546,N_38918);
or U45219 (N_45219,N_33114,N_38741);
nand U45220 (N_45220,N_34489,N_32720);
or U45221 (N_45221,N_37276,N_39570);
nor U45222 (N_45222,N_31434,N_31417);
nand U45223 (N_45223,N_30621,N_39210);
and U45224 (N_45224,N_33526,N_38457);
and U45225 (N_45225,N_30313,N_34650);
nor U45226 (N_45226,N_39379,N_31305);
and U45227 (N_45227,N_31038,N_37157);
or U45228 (N_45228,N_30035,N_38829);
or U45229 (N_45229,N_30610,N_38899);
nand U45230 (N_45230,N_35353,N_33443);
nand U45231 (N_45231,N_38796,N_30741);
nor U45232 (N_45232,N_35957,N_34613);
and U45233 (N_45233,N_38127,N_32156);
and U45234 (N_45234,N_36814,N_37590);
xor U45235 (N_45235,N_31009,N_35586);
and U45236 (N_45236,N_34797,N_38144);
and U45237 (N_45237,N_31228,N_38978);
nor U45238 (N_45238,N_38979,N_36706);
and U45239 (N_45239,N_30257,N_36931);
or U45240 (N_45240,N_35233,N_33912);
and U45241 (N_45241,N_39116,N_35703);
nand U45242 (N_45242,N_34189,N_34823);
nand U45243 (N_45243,N_36023,N_39733);
and U45244 (N_45244,N_32356,N_36287);
and U45245 (N_45245,N_30801,N_34323);
or U45246 (N_45246,N_30529,N_36141);
or U45247 (N_45247,N_33288,N_38089);
and U45248 (N_45248,N_39334,N_31476);
and U45249 (N_45249,N_36214,N_37932);
xor U45250 (N_45250,N_33198,N_38683);
xor U45251 (N_45251,N_38612,N_30898);
and U45252 (N_45252,N_36602,N_34536);
xnor U45253 (N_45253,N_34791,N_36267);
and U45254 (N_45254,N_38660,N_38692);
or U45255 (N_45255,N_30917,N_37966);
or U45256 (N_45256,N_32828,N_38676);
nor U45257 (N_45257,N_36512,N_35764);
nor U45258 (N_45258,N_39865,N_32369);
nor U45259 (N_45259,N_35804,N_31833);
nor U45260 (N_45260,N_31299,N_36628);
xor U45261 (N_45261,N_37794,N_37041);
xor U45262 (N_45262,N_38682,N_36090);
or U45263 (N_45263,N_37186,N_34826);
and U45264 (N_45264,N_31061,N_33396);
nor U45265 (N_45265,N_35987,N_35359);
nand U45266 (N_45266,N_35316,N_38974);
nand U45267 (N_45267,N_37755,N_31817);
xnor U45268 (N_45268,N_36069,N_32466);
or U45269 (N_45269,N_34594,N_30636);
nand U45270 (N_45270,N_31141,N_31854);
nand U45271 (N_45271,N_32665,N_34237);
or U45272 (N_45272,N_36760,N_36624);
nand U45273 (N_45273,N_36070,N_32700);
and U45274 (N_45274,N_39815,N_39595);
xor U45275 (N_45275,N_37129,N_34809);
nand U45276 (N_45276,N_39200,N_31795);
xnor U45277 (N_45277,N_31150,N_30342);
xor U45278 (N_45278,N_38750,N_37071);
nor U45279 (N_45279,N_35848,N_39508);
and U45280 (N_45280,N_33305,N_30995);
and U45281 (N_45281,N_34027,N_34159);
and U45282 (N_45282,N_36482,N_32200);
or U45283 (N_45283,N_33571,N_39048);
or U45284 (N_45284,N_38211,N_34582);
and U45285 (N_45285,N_33435,N_34473);
xor U45286 (N_45286,N_34183,N_33162);
xnor U45287 (N_45287,N_36106,N_34284);
nand U45288 (N_45288,N_37947,N_32251);
xor U45289 (N_45289,N_33852,N_35419);
or U45290 (N_45290,N_31148,N_33100);
xor U45291 (N_45291,N_31957,N_34705);
nor U45292 (N_45292,N_33284,N_34439);
nand U45293 (N_45293,N_30274,N_39210);
or U45294 (N_45294,N_39920,N_31256);
or U45295 (N_45295,N_33591,N_37765);
nand U45296 (N_45296,N_35429,N_34594);
and U45297 (N_45297,N_37166,N_33322);
xor U45298 (N_45298,N_35984,N_37363);
xor U45299 (N_45299,N_35091,N_38732);
and U45300 (N_45300,N_34729,N_32471);
nand U45301 (N_45301,N_37768,N_32041);
nand U45302 (N_45302,N_39617,N_39294);
nand U45303 (N_45303,N_37463,N_34614);
and U45304 (N_45304,N_31200,N_30780);
or U45305 (N_45305,N_32666,N_31858);
nor U45306 (N_45306,N_31089,N_37722);
or U45307 (N_45307,N_33931,N_34693);
and U45308 (N_45308,N_31128,N_34190);
or U45309 (N_45309,N_31170,N_38869);
nand U45310 (N_45310,N_30299,N_30515);
and U45311 (N_45311,N_33195,N_32716);
xnor U45312 (N_45312,N_39123,N_38457);
nor U45313 (N_45313,N_35911,N_34901);
nand U45314 (N_45314,N_36508,N_38388);
xnor U45315 (N_45315,N_38109,N_38290);
or U45316 (N_45316,N_34680,N_33305);
nor U45317 (N_45317,N_31730,N_33586);
or U45318 (N_45318,N_35434,N_35538);
xor U45319 (N_45319,N_32408,N_36290);
xnor U45320 (N_45320,N_35565,N_38219);
nor U45321 (N_45321,N_30999,N_34609);
xnor U45322 (N_45322,N_32299,N_33108);
and U45323 (N_45323,N_31536,N_38237);
nor U45324 (N_45324,N_36121,N_39037);
and U45325 (N_45325,N_32080,N_30756);
or U45326 (N_45326,N_37378,N_30159);
nor U45327 (N_45327,N_32702,N_34211);
or U45328 (N_45328,N_35996,N_34971);
nand U45329 (N_45329,N_35358,N_31121);
and U45330 (N_45330,N_34959,N_39183);
or U45331 (N_45331,N_31152,N_31235);
nor U45332 (N_45332,N_34186,N_39652);
nor U45333 (N_45333,N_30393,N_32919);
xor U45334 (N_45334,N_35363,N_37814);
and U45335 (N_45335,N_31421,N_36065);
and U45336 (N_45336,N_36872,N_32748);
nor U45337 (N_45337,N_39962,N_31356);
nand U45338 (N_45338,N_35696,N_39120);
or U45339 (N_45339,N_37352,N_34951);
nor U45340 (N_45340,N_30774,N_32072);
and U45341 (N_45341,N_35175,N_32199);
nor U45342 (N_45342,N_32815,N_30181);
and U45343 (N_45343,N_39768,N_37906);
or U45344 (N_45344,N_34495,N_32297);
nand U45345 (N_45345,N_35660,N_39192);
or U45346 (N_45346,N_34865,N_30805);
xnor U45347 (N_45347,N_39768,N_39623);
xnor U45348 (N_45348,N_39875,N_34155);
nand U45349 (N_45349,N_33183,N_35511);
or U45350 (N_45350,N_31796,N_31739);
nand U45351 (N_45351,N_35791,N_32780);
and U45352 (N_45352,N_33345,N_38817);
nand U45353 (N_45353,N_36869,N_30108);
or U45354 (N_45354,N_31701,N_36444);
nand U45355 (N_45355,N_39632,N_32580);
nor U45356 (N_45356,N_32866,N_32400);
nand U45357 (N_45357,N_33379,N_37692);
nor U45358 (N_45358,N_30711,N_32682);
nor U45359 (N_45359,N_38895,N_33131);
nand U45360 (N_45360,N_34400,N_35355);
nand U45361 (N_45361,N_32202,N_33320);
nand U45362 (N_45362,N_37727,N_37873);
xnor U45363 (N_45363,N_31382,N_39787);
nor U45364 (N_45364,N_33311,N_31383);
nand U45365 (N_45365,N_30389,N_35443);
nor U45366 (N_45366,N_38503,N_35218);
nand U45367 (N_45367,N_37672,N_39552);
and U45368 (N_45368,N_30322,N_30747);
and U45369 (N_45369,N_35894,N_34520);
xor U45370 (N_45370,N_37385,N_34222);
xnor U45371 (N_45371,N_39843,N_35651);
nand U45372 (N_45372,N_32787,N_33926);
and U45373 (N_45373,N_35853,N_39377);
or U45374 (N_45374,N_31116,N_34439);
nand U45375 (N_45375,N_39554,N_36210);
and U45376 (N_45376,N_37634,N_34651);
nor U45377 (N_45377,N_32412,N_34610);
nand U45378 (N_45378,N_36250,N_36287);
xor U45379 (N_45379,N_30582,N_37379);
or U45380 (N_45380,N_39126,N_33728);
and U45381 (N_45381,N_36729,N_37784);
and U45382 (N_45382,N_34677,N_30057);
and U45383 (N_45383,N_33112,N_38539);
xor U45384 (N_45384,N_31858,N_39203);
or U45385 (N_45385,N_30406,N_35357);
xnor U45386 (N_45386,N_38329,N_31053);
xnor U45387 (N_45387,N_32430,N_39008);
and U45388 (N_45388,N_30234,N_31286);
nor U45389 (N_45389,N_37148,N_39768);
or U45390 (N_45390,N_32494,N_39942);
nand U45391 (N_45391,N_32409,N_39068);
or U45392 (N_45392,N_30723,N_38459);
nor U45393 (N_45393,N_36602,N_30476);
or U45394 (N_45394,N_34436,N_38300);
xnor U45395 (N_45395,N_31898,N_30911);
xnor U45396 (N_45396,N_33953,N_31981);
nand U45397 (N_45397,N_33996,N_39378);
and U45398 (N_45398,N_36615,N_32948);
nor U45399 (N_45399,N_31614,N_32903);
xnor U45400 (N_45400,N_33803,N_38090);
and U45401 (N_45401,N_30783,N_32935);
xnor U45402 (N_45402,N_31035,N_39301);
nor U45403 (N_45403,N_31900,N_39264);
nor U45404 (N_45404,N_32492,N_31278);
nor U45405 (N_45405,N_31351,N_32637);
or U45406 (N_45406,N_33591,N_31728);
or U45407 (N_45407,N_37142,N_31038);
nand U45408 (N_45408,N_39352,N_35832);
nor U45409 (N_45409,N_30096,N_32739);
xor U45410 (N_45410,N_38492,N_34289);
or U45411 (N_45411,N_32877,N_37301);
nand U45412 (N_45412,N_34488,N_34763);
nand U45413 (N_45413,N_30231,N_39108);
and U45414 (N_45414,N_37331,N_37892);
and U45415 (N_45415,N_33320,N_37681);
nor U45416 (N_45416,N_38624,N_33210);
xor U45417 (N_45417,N_39569,N_31386);
nand U45418 (N_45418,N_32270,N_35281);
nor U45419 (N_45419,N_33976,N_38748);
xor U45420 (N_45420,N_38804,N_36181);
nor U45421 (N_45421,N_33103,N_33441);
nor U45422 (N_45422,N_34914,N_37401);
nand U45423 (N_45423,N_38335,N_35577);
or U45424 (N_45424,N_39523,N_39842);
nor U45425 (N_45425,N_36959,N_32190);
nor U45426 (N_45426,N_32361,N_32969);
or U45427 (N_45427,N_37772,N_39918);
or U45428 (N_45428,N_37214,N_37969);
xnor U45429 (N_45429,N_37743,N_35431);
and U45430 (N_45430,N_32086,N_33350);
nor U45431 (N_45431,N_34938,N_39020);
nor U45432 (N_45432,N_37990,N_39244);
and U45433 (N_45433,N_34420,N_31227);
nand U45434 (N_45434,N_35655,N_35892);
xnor U45435 (N_45435,N_32565,N_34039);
and U45436 (N_45436,N_35744,N_35905);
nor U45437 (N_45437,N_38778,N_30151);
or U45438 (N_45438,N_35789,N_38445);
and U45439 (N_45439,N_34909,N_33654);
xor U45440 (N_45440,N_35155,N_38544);
nand U45441 (N_45441,N_39303,N_36895);
and U45442 (N_45442,N_31029,N_37659);
or U45443 (N_45443,N_34792,N_39619);
and U45444 (N_45444,N_30429,N_35894);
nor U45445 (N_45445,N_32926,N_39939);
nand U45446 (N_45446,N_30819,N_31369);
or U45447 (N_45447,N_37893,N_32980);
xnor U45448 (N_45448,N_37391,N_32097);
nand U45449 (N_45449,N_34884,N_31029);
or U45450 (N_45450,N_34838,N_38200);
xor U45451 (N_45451,N_38041,N_36463);
or U45452 (N_45452,N_31173,N_38063);
and U45453 (N_45453,N_34515,N_34850);
nand U45454 (N_45454,N_38028,N_31637);
xnor U45455 (N_45455,N_39984,N_38216);
and U45456 (N_45456,N_30846,N_32784);
or U45457 (N_45457,N_32055,N_30468);
nand U45458 (N_45458,N_37150,N_31239);
nand U45459 (N_45459,N_33336,N_37565);
nand U45460 (N_45460,N_37699,N_35676);
nand U45461 (N_45461,N_35794,N_39159);
and U45462 (N_45462,N_34862,N_33715);
or U45463 (N_45463,N_31222,N_36463);
nor U45464 (N_45464,N_32899,N_39835);
nand U45465 (N_45465,N_39383,N_38633);
nand U45466 (N_45466,N_33495,N_34692);
xnor U45467 (N_45467,N_39274,N_31479);
or U45468 (N_45468,N_36748,N_34573);
nand U45469 (N_45469,N_37045,N_35192);
or U45470 (N_45470,N_32874,N_36689);
nor U45471 (N_45471,N_32339,N_30988);
nor U45472 (N_45472,N_38609,N_34214);
xnor U45473 (N_45473,N_31750,N_33501);
or U45474 (N_45474,N_30515,N_38445);
xor U45475 (N_45475,N_34486,N_36859);
nand U45476 (N_45476,N_33196,N_33182);
xnor U45477 (N_45477,N_39698,N_31308);
or U45478 (N_45478,N_33765,N_30468);
and U45479 (N_45479,N_32439,N_35278);
nand U45480 (N_45480,N_36637,N_32317);
or U45481 (N_45481,N_39022,N_30322);
xor U45482 (N_45482,N_34703,N_34844);
and U45483 (N_45483,N_32937,N_39720);
nand U45484 (N_45484,N_31729,N_36849);
and U45485 (N_45485,N_32235,N_30985);
nand U45486 (N_45486,N_32629,N_33145);
nand U45487 (N_45487,N_39930,N_32728);
and U45488 (N_45488,N_31266,N_35732);
nor U45489 (N_45489,N_30673,N_37142);
or U45490 (N_45490,N_36697,N_35412);
and U45491 (N_45491,N_37549,N_36540);
nor U45492 (N_45492,N_38094,N_30863);
xor U45493 (N_45493,N_31227,N_37790);
and U45494 (N_45494,N_39540,N_30177);
xnor U45495 (N_45495,N_38265,N_36656);
or U45496 (N_45496,N_32254,N_37832);
or U45497 (N_45497,N_32853,N_34945);
or U45498 (N_45498,N_36575,N_39804);
nor U45499 (N_45499,N_37131,N_33866);
nand U45500 (N_45500,N_31712,N_35283);
nand U45501 (N_45501,N_36431,N_32706);
xnor U45502 (N_45502,N_36438,N_35334);
nand U45503 (N_45503,N_37610,N_38098);
xnor U45504 (N_45504,N_35305,N_32536);
nand U45505 (N_45505,N_39595,N_37758);
xnor U45506 (N_45506,N_32994,N_36583);
nand U45507 (N_45507,N_30389,N_33609);
nor U45508 (N_45508,N_36871,N_33353);
and U45509 (N_45509,N_35477,N_36979);
nand U45510 (N_45510,N_33126,N_34277);
nor U45511 (N_45511,N_39908,N_35059);
nand U45512 (N_45512,N_33795,N_34574);
nor U45513 (N_45513,N_33079,N_39658);
or U45514 (N_45514,N_36999,N_36686);
xnor U45515 (N_45515,N_32441,N_31379);
and U45516 (N_45516,N_39829,N_37185);
xnor U45517 (N_45517,N_33346,N_30593);
or U45518 (N_45518,N_32539,N_36646);
and U45519 (N_45519,N_35109,N_31298);
xor U45520 (N_45520,N_30906,N_32951);
and U45521 (N_45521,N_30443,N_38015);
or U45522 (N_45522,N_33546,N_36300);
and U45523 (N_45523,N_35661,N_36195);
and U45524 (N_45524,N_38278,N_33530);
xor U45525 (N_45525,N_33039,N_38676);
and U45526 (N_45526,N_36042,N_35364);
and U45527 (N_45527,N_36850,N_35331);
nand U45528 (N_45528,N_36479,N_35336);
nand U45529 (N_45529,N_39974,N_33462);
and U45530 (N_45530,N_37695,N_39106);
and U45531 (N_45531,N_33226,N_35441);
xor U45532 (N_45532,N_39957,N_37862);
nor U45533 (N_45533,N_34128,N_35672);
nor U45534 (N_45534,N_32732,N_33996);
nand U45535 (N_45535,N_37713,N_39985);
or U45536 (N_45536,N_33786,N_35742);
and U45537 (N_45537,N_31033,N_35711);
and U45538 (N_45538,N_38468,N_37779);
or U45539 (N_45539,N_32477,N_34009);
and U45540 (N_45540,N_39814,N_31877);
nand U45541 (N_45541,N_34018,N_30039);
and U45542 (N_45542,N_30833,N_38601);
nand U45543 (N_45543,N_30814,N_39212);
nand U45544 (N_45544,N_30735,N_31037);
nand U45545 (N_45545,N_38012,N_31298);
nand U45546 (N_45546,N_30353,N_37667);
nand U45547 (N_45547,N_38107,N_30297);
xor U45548 (N_45548,N_37969,N_30801);
nand U45549 (N_45549,N_37261,N_32818);
xor U45550 (N_45550,N_34482,N_34948);
and U45551 (N_45551,N_34718,N_31760);
and U45552 (N_45552,N_37880,N_33479);
and U45553 (N_45553,N_32742,N_38064);
and U45554 (N_45554,N_37497,N_30087);
or U45555 (N_45555,N_35189,N_36502);
nand U45556 (N_45556,N_34469,N_33092);
or U45557 (N_45557,N_35165,N_33369);
or U45558 (N_45558,N_30685,N_31547);
nor U45559 (N_45559,N_32260,N_30428);
nor U45560 (N_45560,N_30032,N_39857);
nor U45561 (N_45561,N_39084,N_33839);
and U45562 (N_45562,N_34397,N_30829);
nor U45563 (N_45563,N_32702,N_38137);
nor U45564 (N_45564,N_32227,N_39687);
nor U45565 (N_45565,N_31594,N_38447);
and U45566 (N_45566,N_35951,N_31813);
or U45567 (N_45567,N_37441,N_35935);
nor U45568 (N_45568,N_35876,N_31508);
and U45569 (N_45569,N_32481,N_36985);
and U45570 (N_45570,N_31213,N_34613);
and U45571 (N_45571,N_30681,N_39860);
or U45572 (N_45572,N_37951,N_39600);
or U45573 (N_45573,N_38467,N_30430);
or U45574 (N_45574,N_32632,N_33799);
xor U45575 (N_45575,N_35774,N_30644);
nand U45576 (N_45576,N_39921,N_37216);
nor U45577 (N_45577,N_31240,N_32210);
xnor U45578 (N_45578,N_33312,N_33115);
nor U45579 (N_45579,N_38932,N_37337);
or U45580 (N_45580,N_35176,N_38428);
or U45581 (N_45581,N_32555,N_33096);
and U45582 (N_45582,N_33277,N_34379);
and U45583 (N_45583,N_38693,N_37812);
xnor U45584 (N_45584,N_33652,N_30906);
nor U45585 (N_45585,N_35834,N_32795);
xnor U45586 (N_45586,N_36455,N_33394);
nand U45587 (N_45587,N_39823,N_31512);
nand U45588 (N_45588,N_39786,N_38741);
nand U45589 (N_45589,N_32525,N_39381);
or U45590 (N_45590,N_38898,N_33319);
and U45591 (N_45591,N_31825,N_31029);
nor U45592 (N_45592,N_32125,N_34564);
or U45593 (N_45593,N_38472,N_35969);
and U45594 (N_45594,N_33531,N_33216);
xor U45595 (N_45595,N_30673,N_35208);
nor U45596 (N_45596,N_35959,N_38103);
xnor U45597 (N_45597,N_33817,N_35019);
or U45598 (N_45598,N_38646,N_30536);
nand U45599 (N_45599,N_31573,N_33638);
or U45600 (N_45600,N_39282,N_33232);
and U45601 (N_45601,N_39772,N_34340);
nand U45602 (N_45602,N_37528,N_35831);
xnor U45603 (N_45603,N_39532,N_38393);
nor U45604 (N_45604,N_33865,N_37874);
or U45605 (N_45605,N_31650,N_30823);
and U45606 (N_45606,N_37424,N_32270);
and U45607 (N_45607,N_30386,N_38952);
xnor U45608 (N_45608,N_36506,N_32908);
xnor U45609 (N_45609,N_30769,N_33578);
xnor U45610 (N_45610,N_35020,N_38062);
and U45611 (N_45611,N_38835,N_32016);
xnor U45612 (N_45612,N_38773,N_30733);
nand U45613 (N_45613,N_38481,N_31685);
xor U45614 (N_45614,N_34582,N_32261);
xnor U45615 (N_45615,N_38595,N_32847);
nand U45616 (N_45616,N_37513,N_30938);
and U45617 (N_45617,N_32780,N_32985);
or U45618 (N_45618,N_35250,N_35523);
nand U45619 (N_45619,N_31279,N_36572);
nand U45620 (N_45620,N_38445,N_30830);
nand U45621 (N_45621,N_38189,N_33329);
xnor U45622 (N_45622,N_35228,N_39101);
and U45623 (N_45623,N_31756,N_37587);
nand U45624 (N_45624,N_33936,N_35396);
xnor U45625 (N_45625,N_30822,N_34361);
or U45626 (N_45626,N_37748,N_33486);
nor U45627 (N_45627,N_31199,N_37126);
or U45628 (N_45628,N_30629,N_30831);
and U45629 (N_45629,N_39746,N_38880);
and U45630 (N_45630,N_34107,N_39598);
or U45631 (N_45631,N_39836,N_33625);
nor U45632 (N_45632,N_35647,N_38679);
xor U45633 (N_45633,N_38403,N_36509);
nand U45634 (N_45634,N_37475,N_31646);
nor U45635 (N_45635,N_36844,N_33008);
nor U45636 (N_45636,N_30247,N_34685);
nand U45637 (N_45637,N_30743,N_32407);
or U45638 (N_45638,N_32761,N_32233);
or U45639 (N_45639,N_31016,N_39348);
or U45640 (N_45640,N_37828,N_39599);
and U45641 (N_45641,N_31257,N_32318);
xor U45642 (N_45642,N_35360,N_36655);
and U45643 (N_45643,N_31070,N_38083);
nand U45644 (N_45644,N_34846,N_36545);
or U45645 (N_45645,N_32300,N_33820);
nand U45646 (N_45646,N_33363,N_34675);
or U45647 (N_45647,N_36536,N_39129);
or U45648 (N_45648,N_31460,N_39363);
nand U45649 (N_45649,N_30280,N_32008);
and U45650 (N_45650,N_34718,N_32202);
nand U45651 (N_45651,N_31771,N_31725);
nand U45652 (N_45652,N_37768,N_31832);
xor U45653 (N_45653,N_33111,N_34325);
and U45654 (N_45654,N_31307,N_30208);
or U45655 (N_45655,N_38839,N_37889);
nand U45656 (N_45656,N_39293,N_37713);
or U45657 (N_45657,N_34486,N_33936);
nor U45658 (N_45658,N_36331,N_39643);
and U45659 (N_45659,N_33362,N_31828);
nor U45660 (N_45660,N_34811,N_37451);
and U45661 (N_45661,N_37813,N_31352);
or U45662 (N_45662,N_38163,N_31879);
nor U45663 (N_45663,N_36188,N_34819);
xor U45664 (N_45664,N_39374,N_37845);
nor U45665 (N_45665,N_35676,N_34178);
nor U45666 (N_45666,N_39200,N_34334);
xor U45667 (N_45667,N_30359,N_32349);
nor U45668 (N_45668,N_39458,N_38803);
and U45669 (N_45669,N_36862,N_30964);
xnor U45670 (N_45670,N_31709,N_31285);
and U45671 (N_45671,N_35379,N_33285);
nand U45672 (N_45672,N_36158,N_32199);
nor U45673 (N_45673,N_38917,N_38448);
nor U45674 (N_45674,N_38922,N_30280);
nand U45675 (N_45675,N_31923,N_35997);
nor U45676 (N_45676,N_37559,N_34749);
nand U45677 (N_45677,N_31918,N_33696);
and U45678 (N_45678,N_31162,N_35870);
nand U45679 (N_45679,N_39664,N_34475);
nor U45680 (N_45680,N_35629,N_35774);
nor U45681 (N_45681,N_37219,N_37879);
nor U45682 (N_45682,N_36140,N_36993);
and U45683 (N_45683,N_33371,N_30474);
nand U45684 (N_45684,N_38131,N_34746);
xor U45685 (N_45685,N_31411,N_31086);
and U45686 (N_45686,N_39475,N_32129);
nor U45687 (N_45687,N_31110,N_38796);
nand U45688 (N_45688,N_38401,N_37490);
xor U45689 (N_45689,N_30557,N_36443);
nand U45690 (N_45690,N_38374,N_33298);
nand U45691 (N_45691,N_38866,N_30195);
or U45692 (N_45692,N_36904,N_31892);
xnor U45693 (N_45693,N_31204,N_35160);
nand U45694 (N_45694,N_33139,N_38286);
nor U45695 (N_45695,N_30799,N_30489);
nand U45696 (N_45696,N_32676,N_34436);
xnor U45697 (N_45697,N_36007,N_36473);
or U45698 (N_45698,N_33585,N_31727);
nor U45699 (N_45699,N_39514,N_35345);
and U45700 (N_45700,N_38133,N_39791);
xnor U45701 (N_45701,N_34679,N_31127);
or U45702 (N_45702,N_38056,N_32257);
nand U45703 (N_45703,N_32950,N_36146);
nand U45704 (N_45704,N_31211,N_33850);
or U45705 (N_45705,N_37183,N_30407);
and U45706 (N_45706,N_31618,N_32046);
nand U45707 (N_45707,N_36702,N_31770);
or U45708 (N_45708,N_37195,N_34551);
or U45709 (N_45709,N_39290,N_32698);
xor U45710 (N_45710,N_36210,N_38784);
or U45711 (N_45711,N_32875,N_30253);
or U45712 (N_45712,N_33606,N_37194);
nand U45713 (N_45713,N_37113,N_34717);
or U45714 (N_45714,N_36238,N_31392);
or U45715 (N_45715,N_32355,N_38708);
or U45716 (N_45716,N_35086,N_35012);
or U45717 (N_45717,N_32169,N_35577);
and U45718 (N_45718,N_31297,N_35760);
and U45719 (N_45719,N_39530,N_31245);
nor U45720 (N_45720,N_31807,N_39569);
nor U45721 (N_45721,N_31372,N_38727);
and U45722 (N_45722,N_32829,N_38658);
or U45723 (N_45723,N_31410,N_35780);
or U45724 (N_45724,N_39076,N_39954);
and U45725 (N_45725,N_36073,N_31047);
xnor U45726 (N_45726,N_39134,N_32827);
and U45727 (N_45727,N_37998,N_39947);
nand U45728 (N_45728,N_36095,N_34201);
xor U45729 (N_45729,N_38495,N_30104);
nand U45730 (N_45730,N_33546,N_32643);
and U45731 (N_45731,N_38860,N_31870);
and U45732 (N_45732,N_32167,N_39455);
nand U45733 (N_45733,N_31362,N_31942);
or U45734 (N_45734,N_34776,N_31235);
or U45735 (N_45735,N_36457,N_34931);
xnor U45736 (N_45736,N_32766,N_35484);
and U45737 (N_45737,N_30850,N_34642);
or U45738 (N_45738,N_36743,N_36957);
nor U45739 (N_45739,N_36625,N_33775);
nand U45740 (N_45740,N_31648,N_37953);
xor U45741 (N_45741,N_31471,N_38339);
nor U45742 (N_45742,N_38665,N_31210);
and U45743 (N_45743,N_35575,N_31759);
and U45744 (N_45744,N_32114,N_37225);
nand U45745 (N_45745,N_32584,N_34884);
and U45746 (N_45746,N_33911,N_38972);
nor U45747 (N_45747,N_32817,N_39596);
nand U45748 (N_45748,N_35029,N_31758);
nand U45749 (N_45749,N_32752,N_35847);
and U45750 (N_45750,N_37049,N_34986);
or U45751 (N_45751,N_37359,N_36168);
nand U45752 (N_45752,N_34332,N_31924);
xor U45753 (N_45753,N_31502,N_35741);
or U45754 (N_45754,N_36835,N_36821);
nor U45755 (N_45755,N_30009,N_35679);
or U45756 (N_45756,N_33661,N_34259);
and U45757 (N_45757,N_33243,N_36854);
nor U45758 (N_45758,N_35359,N_34530);
or U45759 (N_45759,N_34466,N_39503);
xor U45760 (N_45760,N_36375,N_38025);
or U45761 (N_45761,N_33001,N_30310);
xnor U45762 (N_45762,N_37784,N_39014);
xnor U45763 (N_45763,N_33973,N_38551);
nand U45764 (N_45764,N_31695,N_33102);
nand U45765 (N_45765,N_37071,N_38874);
xor U45766 (N_45766,N_36760,N_32405);
or U45767 (N_45767,N_34040,N_39317);
or U45768 (N_45768,N_35588,N_35813);
xnor U45769 (N_45769,N_31125,N_34067);
nor U45770 (N_45770,N_36108,N_36187);
and U45771 (N_45771,N_38125,N_38186);
and U45772 (N_45772,N_39168,N_33556);
and U45773 (N_45773,N_33183,N_33699);
xor U45774 (N_45774,N_33880,N_36090);
xnor U45775 (N_45775,N_33935,N_32781);
nor U45776 (N_45776,N_31125,N_35054);
and U45777 (N_45777,N_34565,N_37283);
or U45778 (N_45778,N_31479,N_36900);
nor U45779 (N_45779,N_32009,N_34509);
xor U45780 (N_45780,N_31872,N_33525);
xnor U45781 (N_45781,N_36091,N_36909);
or U45782 (N_45782,N_34425,N_38591);
xor U45783 (N_45783,N_39541,N_30600);
xnor U45784 (N_45784,N_30174,N_35161);
nor U45785 (N_45785,N_36704,N_34351);
and U45786 (N_45786,N_33013,N_39112);
nand U45787 (N_45787,N_35641,N_33843);
or U45788 (N_45788,N_31038,N_30709);
nor U45789 (N_45789,N_37526,N_32800);
or U45790 (N_45790,N_35118,N_37948);
nor U45791 (N_45791,N_31940,N_35438);
xnor U45792 (N_45792,N_30514,N_32486);
xor U45793 (N_45793,N_30960,N_30854);
or U45794 (N_45794,N_39974,N_35481);
or U45795 (N_45795,N_37664,N_34719);
and U45796 (N_45796,N_33367,N_36238);
xnor U45797 (N_45797,N_30026,N_36072);
nor U45798 (N_45798,N_32409,N_38865);
and U45799 (N_45799,N_33988,N_33499);
nor U45800 (N_45800,N_36799,N_38537);
xnor U45801 (N_45801,N_34382,N_39969);
nand U45802 (N_45802,N_36829,N_38206);
nor U45803 (N_45803,N_38489,N_34368);
or U45804 (N_45804,N_34708,N_39056);
nand U45805 (N_45805,N_38556,N_30613);
xor U45806 (N_45806,N_35824,N_32982);
xor U45807 (N_45807,N_37168,N_33595);
or U45808 (N_45808,N_33995,N_38840);
nor U45809 (N_45809,N_38955,N_30478);
nor U45810 (N_45810,N_34472,N_36938);
nor U45811 (N_45811,N_30625,N_34309);
and U45812 (N_45812,N_30074,N_31580);
nor U45813 (N_45813,N_34464,N_30875);
nand U45814 (N_45814,N_38953,N_30791);
nand U45815 (N_45815,N_33452,N_33089);
or U45816 (N_45816,N_31715,N_32509);
nor U45817 (N_45817,N_33224,N_34947);
xnor U45818 (N_45818,N_35875,N_37254);
or U45819 (N_45819,N_31611,N_31997);
nand U45820 (N_45820,N_35689,N_33757);
and U45821 (N_45821,N_38017,N_33898);
nand U45822 (N_45822,N_34825,N_30862);
nor U45823 (N_45823,N_39708,N_34282);
xor U45824 (N_45824,N_30854,N_36791);
nand U45825 (N_45825,N_33760,N_36231);
or U45826 (N_45826,N_35006,N_34857);
xnor U45827 (N_45827,N_38085,N_32512);
or U45828 (N_45828,N_30810,N_36738);
or U45829 (N_45829,N_35714,N_33396);
or U45830 (N_45830,N_36063,N_30563);
xor U45831 (N_45831,N_35614,N_33777);
xor U45832 (N_45832,N_39007,N_37491);
xnor U45833 (N_45833,N_33668,N_34887);
nand U45834 (N_45834,N_30075,N_36259);
nand U45835 (N_45835,N_34467,N_39844);
and U45836 (N_45836,N_33082,N_32301);
or U45837 (N_45837,N_32882,N_37729);
and U45838 (N_45838,N_34730,N_39741);
nor U45839 (N_45839,N_30293,N_30141);
nand U45840 (N_45840,N_30284,N_34934);
nor U45841 (N_45841,N_39637,N_36312);
nand U45842 (N_45842,N_37527,N_35299);
nor U45843 (N_45843,N_38395,N_39111);
and U45844 (N_45844,N_38969,N_35350);
xor U45845 (N_45845,N_38279,N_37286);
or U45846 (N_45846,N_34505,N_39287);
or U45847 (N_45847,N_36250,N_37917);
or U45848 (N_45848,N_34090,N_30930);
nor U45849 (N_45849,N_36049,N_30174);
xor U45850 (N_45850,N_33467,N_33779);
nand U45851 (N_45851,N_34629,N_36525);
nor U45852 (N_45852,N_38268,N_36445);
or U45853 (N_45853,N_35143,N_32332);
xor U45854 (N_45854,N_37840,N_30614);
and U45855 (N_45855,N_39840,N_30904);
nor U45856 (N_45856,N_36020,N_37425);
nor U45857 (N_45857,N_33641,N_38869);
and U45858 (N_45858,N_33234,N_37715);
xor U45859 (N_45859,N_31065,N_31349);
nor U45860 (N_45860,N_32242,N_39924);
and U45861 (N_45861,N_36914,N_31638);
nor U45862 (N_45862,N_34832,N_33160);
and U45863 (N_45863,N_31872,N_36380);
or U45864 (N_45864,N_31817,N_38886);
and U45865 (N_45865,N_32949,N_35918);
or U45866 (N_45866,N_39797,N_34802);
xor U45867 (N_45867,N_36037,N_38401);
nand U45868 (N_45868,N_39632,N_30547);
and U45869 (N_45869,N_30389,N_38838);
nor U45870 (N_45870,N_30744,N_36174);
nor U45871 (N_45871,N_34522,N_39081);
or U45872 (N_45872,N_39448,N_37075);
nand U45873 (N_45873,N_32285,N_39376);
xor U45874 (N_45874,N_31566,N_39516);
nor U45875 (N_45875,N_39258,N_31472);
nor U45876 (N_45876,N_31521,N_31063);
or U45877 (N_45877,N_38068,N_37045);
xnor U45878 (N_45878,N_34941,N_36650);
nand U45879 (N_45879,N_39569,N_30604);
or U45880 (N_45880,N_34288,N_39442);
or U45881 (N_45881,N_30299,N_33256);
nor U45882 (N_45882,N_33455,N_31806);
or U45883 (N_45883,N_36851,N_31711);
xnor U45884 (N_45884,N_38317,N_33273);
nor U45885 (N_45885,N_33323,N_30152);
nor U45886 (N_45886,N_38330,N_36301);
xnor U45887 (N_45887,N_33112,N_34430);
xor U45888 (N_45888,N_35713,N_30759);
nor U45889 (N_45889,N_34125,N_31830);
xnor U45890 (N_45890,N_34065,N_39935);
nand U45891 (N_45891,N_33594,N_37424);
and U45892 (N_45892,N_31706,N_31646);
and U45893 (N_45893,N_34691,N_39618);
xnor U45894 (N_45894,N_37007,N_39682);
and U45895 (N_45895,N_33370,N_39212);
xnor U45896 (N_45896,N_32913,N_32328);
nor U45897 (N_45897,N_31660,N_37617);
nor U45898 (N_45898,N_33196,N_35555);
nor U45899 (N_45899,N_38801,N_33118);
or U45900 (N_45900,N_31095,N_38433);
nand U45901 (N_45901,N_38850,N_32122);
or U45902 (N_45902,N_31974,N_30165);
xnor U45903 (N_45903,N_34321,N_34427);
nand U45904 (N_45904,N_36274,N_35615);
xnor U45905 (N_45905,N_30462,N_33668);
nor U45906 (N_45906,N_34553,N_36824);
xor U45907 (N_45907,N_35660,N_36436);
nor U45908 (N_45908,N_32834,N_32370);
and U45909 (N_45909,N_30224,N_37654);
xor U45910 (N_45910,N_35890,N_32958);
xnor U45911 (N_45911,N_35344,N_33404);
and U45912 (N_45912,N_32281,N_37004);
or U45913 (N_45913,N_31632,N_33356);
and U45914 (N_45914,N_30720,N_32651);
nor U45915 (N_45915,N_36698,N_36738);
nand U45916 (N_45916,N_39997,N_30503);
xor U45917 (N_45917,N_39053,N_36839);
nand U45918 (N_45918,N_35550,N_34383);
nor U45919 (N_45919,N_33969,N_37346);
nand U45920 (N_45920,N_31387,N_30043);
xor U45921 (N_45921,N_30193,N_31950);
and U45922 (N_45922,N_37921,N_39074);
xnor U45923 (N_45923,N_36535,N_34558);
nand U45924 (N_45924,N_37220,N_32380);
xnor U45925 (N_45925,N_33106,N_34220);
nand U45926 (N_45926,N_35018,N_31515);
or U45927 (N_45927,N_39508,N_36700);
nand U45928 (N_45928,N_34609,N_33744);
nor U45929 (N_45929,N_30619,N_37979);
xnor U45930 (N_45930,N_36566,N_34365);
nor U45931 (N_45931,N_38557,N_36239);
xor U45932 (N_45932,N_32180,N_30140);
xor U45933 (N_45933,N_33418,N_35284);
nand U45934 (N_45934,N_33158,N_32057);
nor U45935 (N_45935,N_37105,N_37230);
nand U45936 (N_45936,N_34820,N_36145);
and U45937 (N_45937,N_36533,N_33411);
nor U45938 (N_45938,N_30836,N_31881);
or U45939 (N_45939,N_34469,N_38125);
xor U45940 (N_45940,N_36377,N_35659);
and U45941 (N_45941,N_31800,N_39881);
xor U45942 (N_45942,N_33210,N_33235);
nand U45943 (N_45943,N_38772,N_32465);
and U45944 (N_45944,N_36910,N_39443);
or U45945 (N_45945,N_36425,N_33563);
and U45946 (N_45946,N_33375,N_36135);
nand U45947 (N_45947,N_30983,N_33141);
or U45948 (N_45948,N_35970,N_39811);
or U45949 (N_45949,N_33488,N_34003);
nand U45950 (N_45950,N_35515,N_38546);
and U45951 (N_45951,N_34002,N_37274);
and U45952 (N_45952,N_32783,N_34046);
or U45953 (N_45953,N_38708,N_32715);
nand U45954 (N_45954,N_39121,N_37138);
nand U45955 (N_45955,N_36268,N_32593);
xor U45956 (N_45956,N_36045,N_37834);
nor U45957 (N_45957,N_39422,N_35058);
xor U45958 (N_45958,N_30095,N_34216);
nand U45959 (N_45959,N_32385,N_34291);
xnor U45960 (N_45960,N_36250,N_35805);
nor U45961 (N_45961,N_37073,N_34519);
xnor U45962 (N_45962,N_34532,N_30363);
nand U45963 (N_45963,N_36722,N_31430);
and U45964 (N_45964,N_39420,N_36881);
xor U45965 (N_45965,N_38717,N_32838);
nand U45966 (N_45966,N_32295,N_39540);
nor U45967 (N_45967,N_32903,N_31537);
nand U45968 (N_45968,N_33350,N_34315);
and U45969 (N_45969,N_33977,N_37256);
nand U45970 (N_45970,N_33806,N_37332);
nor U45971 (N_45971,N_32955,N_38575);
nor U45972 (N_45972,N_36311,N_36124);
nor U45973 (N_45973,N_37577,N_38147);
xor U45974 (N_45974,N_32582,N_31003);
and U45975 (N_45975,N_33527,N_39859);
or U45976 (N_45976,N_32992,N_36645);
nand U45977 (N_45977,N_30437,N_33603);
nor U45978 (N_45978,N_35613,N_30444);
nor U45979 (N_45979,N_34482,N_39341);
nand U45980 (N_45980,N_39028,N_30183);
nor U45981 (N_45981,N_38763,N_33636);
nand U45982 (N_45982,N_37013,N_38442);
xor U45983 (N_45983,N_33104,N_33056);
xor U45984 (N_45984,N_35827,N_38974);
nand U45985 (N_45985,N_31015,N_39928);
nand U45986 (N_45986,N_37190,N_38592);
or U45987 (N_45987,N_32498,N_31401);
or U45988 (N_45988,N_30381,N_36496);
xnor U45989 (N_45989,N_36076,N_30577);
nor U45990 (N_45990,N_32415,N_37668);
xnor U45991 (N_45991,N_36228,N_37890);
and U45992 (N_45992,N_38142,N_31174);
nand U45993 (N_45993,N_30418,N_38712);
nand U45994 (N_45994,N_35608,N_35098);
and U45995 (N_45995,N_35130,N_37976);
and U45996 (N_45996,N_32975,N_31874);
nor U45997 (N_45997,N_30478,N_35726);
nor U45998 (N_45998,N_38444,N_35213);
or U45999 (N_45999,N_39796,N_33878);
nor U46000 (N_46000,N_34053,N_36559);
nor U46001 (N_46001,N_32261,N_31264);
and U46002 (N_46002,N_36198,N_35601);
and U46003 (N_46003,N_35317,N_33038);
xor U46004 (N_46004,N_34917,N_31477);
xnor U46005 (N_46005,N_39017,N_36127);
nand U46006 (N_46006,N_38315,N_34410);
nor U46007 (N_46007,N_34804,N_32240);
nand U46008 (N_46008,N_35418,N_31426);
or U46009 (N_46009,N_34520,N_35181);
xnor U46010 (N_46010,N_32959,N_32687);
or U46011 (N_46011,N_32174,N_37807);
nand U46012 (N_46012,N_30653,N_34697);
xnor U46013 (N_46013,N_33665,N_33998);
nor U46014 (N_46014,N_39848,N_31936);
and U46015 (N_46015,N_38303,N_30826);
or U46016 (N_46016,N_35219,N_31215);
and U46017 (N_46017,N_36881,N_31313);
or U46018 (N_46018,N_31510,N_32254);
nor U46019 (N_46019,N_38327,N_34072);
or U46020 (N_46020,N_38385,N_37194);
or U46021 (N_46021,N_35323,N_33754);
xnor U46022 (N_46022,N_33007,N_31038);
nand U46023 (N_46023,N_38928,N_37227);
nor U46024 (N_46024,N_38246,N_37233);
nand U46025 (N_46025,N_36720,N_39479);
xnor U46026 (N_46026,N_38031,N_35992);
nand U46027 (N_46027,N_37613,N_30766);
and U46028 (N_46028,N_36860,N_38696);
or U46029 (N_46029,N_36618,N_34234);
nand U46030 (N_46030,N_35816,N_31341);
and U46031 (N_46031,N_36181,N_36349);
nor U46032 (N_46032,N_39084,N_37506);
nor U46033 (N_46033,N_32148,N_32489);
nand U46034 (N_46034,N_31839,N_38465);
or U46035 (N_46035,N_38424,N_37774);
xor U46036 (N_46036,N_39708,N_30610);
and U46037 (N_46037,N_33651,N_33376);
nand U46038 (N_46038,N_34919,N_34258);
nor U46039 (N_46039,N_32557,N_33587);
nand U46040 (N_46040,N_39589,N_33495);
or U46041 (N_46041,N_39484,N_32922);
xnor U46042 (N_46042,N_38586,N_34912);
and U46043 (N_46043,N_35177,N_38358);
xor U46044 (N_46044,N_39229,N_38362);
and U46045 (N_46045,N_34204,N_36602);
or U46046 (N_46046,N_39675,N_35716);
and U46047 (N_46047,N_31106,N_35405);
nor U46048 (N_46048,N_33688,N_35626);
xor U46049 (N_46049,N_30708,N_32746);
nor U46050 (N_46050,N_34895,N_30347);
and U46051 (N_46051,N_31550,N_30008);
nand U46052 (N_46052,N_39697,N_30766);
and U46053 (N_46053,N_34732,N_39846);
nor U46054 (N_46054,N_31311,N_34913);
xor U46055 (N_46055,N_35861,N_30596);
nor U46056 (N_46056,N_38919,N_31562);
nor U46057 (N_46057,N_36449,N_30995);
xnor U46058 (N_46058,N_31729,N_36929);
xnor U46059 (N_46059,N_32768,N_30749);
or U46060 (N_46060,N_35112,N_32655);
xnor U46061 (N_46061,N_30339,N_37504);
nor U46062 (N_46062,N_37384,N_34297);
nand U46063 (N_46063,N_37799,N_37168);
nor U46064 (N_46064,N_37119,N_39152);
or U46065 (N_46065,N_33519,N_31238);
nand U46066 (N_46066,N_36862,N_32786);
nand U46067 (N_46067,N_36043,N_39971);
and U46068 (N_46068,N_32542,N_36371);
xnor U46069 (N_46069,N_37091,N_38715);
nand U46070 (N_46070,N_37390,N_35797);
nor U46071 (N_46071,N_31500,N_38228);
nand U46072 (N_46072,N_31228,N_36311);
and U46073 (N_46073,N_34933,N_32976);
nor U46074 (N_46074,N_30513,N_37476);
and U46075 (N_46075,N_35381,N_33167);
and U46076 (N_46076,N_32346,N_35296);
and U46077 (N_46077,N_35557,N_38849);
or U46078 (N_46078,N_38170,N_33779);
or U46079 (N_46079,N_32108,N_30153);
nor U46080 (N_46080,N_33144,N_37794);
xnor U46081 (N_46081,N_34172,N_30968);
nor U46082 (N_46082,N_30322,N_38882);
xor U46083 (N_46083,N_38125,N_39651);
or U46084 (N_46084,N_30356,N_33892);
nand U46085 (N_46085,N_39321,N_34406);
nor U46086 (N_46086,N_35883,N_31380);
nor U46087 (N_46087,N_30112,N_35555);
or U46088 (N_46088,N_30565,N_36735);
nor U46089 (N_46089,N_34229,N_38914);
nand U46090 (N_46090,N_35891,N_39045);
nor U46091 (N_46091,N_37911,N_37723);
and U46092 (N_46092,N_35536,N_38234);
nand U46093 (N_46093,N_38128,N_32769);
and U46094 (N_46094,N_35714,N_35825);
nor U46095 (N_46095,N_36964,N_35687);
xor U46096 (N_46096,N_38688,N_38370);
xor U46097 (N_46097,N_36650,N_32627);
or U46098 (N_46098,N_32498,N_38242);
xnor U46099 (N_46099,N_36416,N_34473);
or U46100 (N_46100,N_37464,N_39602);
and U46101 (N_46101,N_32977,N_31688);
nand U46102 (N_46102,N_31513,N_37037);
nor U46103 (N_46103,N_31655,N_39609);
or U46104 (N_46104,N_38075,N_31591);
xnor U46105 (N_46105,N_34930,N_37770);
nand U46106 (N_46106,N_33140,N_36461);
or U46107 (N_46107,N_35631,N_31846);
and U46108 (N_46108,N_37808,N_37367);
nor U46109 (N_46109,N_37011,N_34193);
nor U46110 (N_46110,N_31032,N_35856);
nand U46111 (N_46111,N_32975,N_32745);
nor U46112 (N_46112,N_32620,N_31286);
or U46113 (N_46113,N_38563,N_39961);
nor U46114 (N_46114,N_35286,N_39770);
xor U46115 (N_46115,N_38744,N_34794);
and U46116 (N_46116,N_39888,N_32408);
nor U46117 (N_46117,N_30642,N_38379);
nor U46118 (N_46118,N_39513,N_37741);
nand U46119 (N_46119,N_34820,N_33380);
or U46120 (N_46120,N_37799,N_36957);
nor U46121 (N_46121,N_37294,N_30052);
nor U46122 (N_46122,N_39018,N_34351);
nor U46123 (N_46123,N_38648,N_32841);
or U46124 (N_46124,N_31171,N_34511);
nor U46125 (N_46125,N_36213,N_36175);
xor U46126 (N_46126,N_35862,N_31954);
nor U46127 (N_46127,N_35262,N_39976);
nand U46128 (N_46128,N_31360,N_35791);
xnor U46129 (N_46129,N_30145,N_30580);
and U46130 (N_46130,N_33688,N_36771);
and U46131 (N_46131,N_38089,N_31983);
xnor U46132 (N_46132,N_35471,N_39479);
nor U46133 (N_46133,N_30426,N_36084);
or U46134 (N_46134,N_39722,N_35967);
or U46135 (N_46135,N_35079,N_35045);
or U46136 (N_46136,N_34837,N_36380);
or U46137 (N_46137,N_38602,N_33299);
xnor U46138 (N_46138,N_37122,N_31931);
xnor U46139 (N_46139,N_33077,N_36235);
nor U46140 (N_46140,N_39913,N_35390);
nor U46141 (N_46141,N_33133,N_30402);
or U46142 (N_46142,N_31537,N_38495);
and U46143 (N_46143,N_32022,N_32632);
or U46144 (N_46144,N_31485,N_39168);
nand U46145 (N_46145,N_33097,N_38353);
and U46146 (N_46146,N_35097,N_33666);
xnor U46147 (N_46147,N_38293,N_30409);
and U46148 (N_46148,N_39438,N_33110);
and U46149 (N_46149,N_39697,N_37021);
or U46150 (N_46150,N_36699,N_33730);
xor U46151 (N_46151,N_36998,N_31178);
and U46152 (N_46152,N_38775,N_33173);
and U46153 (N_46153,N_30505,N_38850);
xnor U46154 (N_46154,N_38202,N_36501);
and U46155 (N_46155,N_39067,N_38418);
nand U46156 (N_46156,N_32672,N_31987);
nor U46157 (N_46157,N_34246,N_34822);
and U46158 (N_46158,N_33939,N_30108);
xor U46159 (N_46159,N_39165,N_39587);
xnor U46160 (N_46160,N_33051,N_31859);
nand U46161 (N_46161,N_36578,N_35196);
xnor U46162 (N_46162,N_39791,N_38150);
xnor U46163 (N_46163,N_34734,N_35905);
and U46164 (N_46164,N_30511,N_30137);
and U46165 (N_46165,N_31701,N_31158);
or U46166 (N_46166,N_32312,N_37035);
xnor U46167 (N_46167,N_37321,N_38401);
xor U46168 (N_46168,N_35791,N_35195);
or U46169 (N_46169,N_34936,N_30107);
or U46170 (N_46170,N_32101,N_31215);
nand U46171 (N_46171,N_35593,N_30614);
nor U46172 (N_46172,N_36415,N_31151);
and U46173 (N_46173,N_31823,N_31493);
or U46174 (N_46174,N_33523,N_32714);
and U46175 (N_46175,N_37052,N_32728);
nor U46176 (N_46176,N_30937,N_35023);
xnor U46177 (N_46177,N_31645,N_32716);
or U46178 (N_46178,N_37146,N_38377);
nor U46179 (N_46179,N_34000,N_33564);
and U46180 (N_46180,N_35060,N_39953);
xor U46181 (N_46181,N_34543,N_37229);
xnor U46182 (N_46182,N_30605,N_35199);
nand U46183 (N_46183,N_30736,N_39867);
xor U46184 (N_46184,N_30982,N_38411);
or U46185 (N_46185,N_34617,N_35412);
or U46186 (N_46186,N_35601,N_31740);
and U46187 (N_46187,N_33084,N_35586);
nor U46188 (N_46188,N_32849,N_31668);
or U46189 (N_46189,N_34711,N_34599);
nand U46190 (N_46190,N_37202,N_31988);
or U46191 (N_46191,N_38173,N_32249);
xnor U46192 (N_46192,N_37644,N_32543);
or U46193 (N_46193,N_30519,N_38774);
nand U46194 (N_46194,N_35745,N_30173);
xnor U46195 (N_46195,N_36254,N_32082);
and U46196 (N_46196,N_30136,N_30249);
nor U46197 (N_46197,N_39561,N_33535);
or U46198 (N_46198,N_38463,N_37792);
xor U46199 (N_46199,N_39629,N_38819);
or U46200 (N_46200,N_30505,N_38821);
nor U46201 (N_46201,N_37590,N_35472);
xor U46202 (N_46202,N_36839,N_35468);
xor U46203 (N_46203,N_35390,N_36529);
nor U46204 (N_46204,N_30535,N_36776);
or U46205 (N_46205,N_35241,N_33268);
nand U46206 (N_46206,N_33907,N_38366);
and U46207 (N_46207,N_32795,N_38696);
or U46208 (N_46208,N_30443,N_36073);
or U46209 (N_46209,N_30175,N_33503);
and U46210 (N_46210,N_38504,N_32085);
nand U46211 (N_46211,N_33510,N_39370);
and U46212 (N_46212,N_36583,N_34230);
xor U46213 (N_46213,N_39914,N_30972);
xnor U46214 (N_46214,N_37696,N_37689);
xor U46215 (N_46215,N_39271,N_38865);
nand U46216 (N_46216,N_30743,N_35747);
and U46217 (N_46217,N_30622,N_36020);
and U46218 (N_46218,N_36975,N_39030);
nor U46219 (N_46219,N_32208,N_30394);
xor U46220 (N_46220,N_30236,N_38123);
or U46221 (N_46221,N_38619,N_30221);
xor U46222 (N_46222,N_38527,N_36838);
and U46223 (N_46223,N_36821,N_32460);
and U46224 (N_46224,N_38679,N_34889);
and U46225 (N_46225,N_39823,N_38155);
and U46226 (N_46226,N_36325,N_34688);
or U46227 (N_46227,N_35524,N_37799);
nand U46228 (N_46228,N_39308,N_31003);
nor U46229 (N_46229,N_36435,N_30040);
nor U46230 (N_46230,N_34609,N_33989);
and U46231 (N_46231,N_37313,N_36290);
or U46232 (N_46232,N_32370,N_37732);
and U46233 (N_46233,N_32930,N_35082);
nor U46234 (N_46234,N_33379,N_35000);
nor U46235 (N_46235,N_38180,N_32193);
nand U46236 (N_46236,N_37111,N_30392);
nor U46237 (N_46237,N_36914,N_37505);
nand U46238 (N_46238,N_38022,N_38364);
nand U46239 (N_46239,N_38420,N_36965);
nor U46240 (N_46240,N_31810,N_34343);
or U46241 (N_46241,N_30924,N_34578);
xor U46242 (N_46242,N_34543,N_32802);
nor U46243 (N_46243,N_35478,N_31246);
or U46244 (N_46244,N_37702,N_32661);
xnor U46245 (N_46245,N_33383,N_31678);
nor U46246 (N_46246,N_36311,N_39409);
nor U46247 (N_46247,N_31448,N_33239);
xor U46248 (N_46248,N_38215,N_31295);
nand U46249 (N_46249,N_33173,N_35988);
nand U46250 (N_46250,N_34050,N_39413);
or U46251 (N_46251,N_37751,N_31181);
nand U46252 (N_46252,N_34541,N_39436);
or U46253 (N_46253,N_39305,N_37593);
and U46254 (N_46254,N_39008,N_39736);
or U46255 (N_46255,N_36377,N_34635);
and U46256 (N_46256,N_39203,N_33750);
or U46257 (N_46257,N_35680,N_35594);
nor U46258 (N_46258,N_34760,N_31263);
nor U46259 (N_46259,N_36948,N_31173);
nand U46260 (N_46260,N_31458,N_38417);
nand U46261 (N_46261,N_32119,N_38720);
nor U46262 (N_46262,N_33805,N_37739);
nand U46263 (N_46263,N_34464,N_32528);
and U46264 (N_46264,N_33238,N_36792);
nand U46265 (N_46265,N_30320,N_32365);
xor U46266 (N_46266,N_30449,N_32560);
xnor U46267 (N_46267,N_36748,N_33267);
nand U46268 (N_46268,N_34471,N_32905);
nand U46269 (N_46269,N_30494,N_39486);
nor U46270 (N_46270,N_30900,N_39967);
nor U46271 (N_46271,N_36349,N_31447);
nor U46272 (N_46272,N_30716,N_34837);
nor U46273 (N_46273,N_34917,N_33549);
nand U46274 (N_46274,N_34671,N_31747);
and U46275 (N_46275,N_33251,N_38061);
nor U46276 (N_46276,N_39548,N_33373);
and U46277 (N_46277,N_37388,N_39339);
and U46278 (N_46278,N_37324,N_39036);
and U46279 (N_46279,N_31853,N_37393);
and U46280 (N_46280,N_32420,N_38481);
or U46281 (N_46281,N_33104,N_34620);
and U46282 (N_46282,N_38005,N_33130);
xor U46283 (N_46283,N_32586,N_31789);
or U46284 (N_46284,N_34655,N_35563);
and U46285 (N_46285,N_30941,N_39491);
and U46286 (N_46286,N_30222,N_34130);
nor U46287 (N_46287,N_34236,N_32032);
nor U46288 (N_46288,N_39682,N_36810);
nor U46289 (N_46289,N_32524,N_35584);
nand U46290 (N_46290,N_34963,N_32525);
or U46291 (N_46291,N_36649,N_35360);
nor U46292 (N_46292,N_34805,N_32906);
and U46293 (N_46293,N_39920,N_36034);
or U46294 (N_46294,N_31286,N_37556);
nand U46295 (N_46295,N_32912,N_38385);
nand U46296 (N_46296,N_37196,N_35580);
and U46297 (N_46297,N_31669,N_38030);
and U46298 (N_46298,N_30065,N_31149);
nor U46299 (N_46299,N_31059,N_31709);
xnor U46300 (N_46300,N_38277,N_36866);
xnor U46301 (N_46301,N_33668,N_35869);
nor U46302 (N_46302,N_33060,N_35295);
or U46303 (N_46303,N_34061,N_33482);
or U46304 (N_46304,N_39227,N_35721);
and U46305 (N_46305,N_39100,N_32680);
nor U46306 (N_46306,N_32094,N_39418);
nor U46307 (N_46307,N_35075,N_34307);
or U46308 (N_46308,N_38029,N_39311);
and U46309 (N_46309,N_39647,N_34623);
or U46310 (N_46310,N_31808,N_32364);
xnor U46311 (N_46311,N_31039,N_35739);
or U46312 (N_46312,N_34144,N_34857);
nor U46313 (N_46313,N_31072,N_38317);
and U46314 (N_46314,N_31253,N_35650);
nor U46315 (N_46315,N_39379,N_39176);
nand U46316 (N_46316,N_37638,N_30251);
nor U46317 (N_46317,N_36091,N_36686);
or U46318 (N_46318,N_30601,N_33471);
xor U46319 (N_46319,N_37378,N_35794);
xor U46320 (N_46320,N_30925,N_39156);
xor U46321 (N_46321,N_39598,N_34214);
xor U46322 (N_46322,N_36742,N_33412);
xor U46323 (N_46323,N_30720,N_36047);
xor U46324 (N_46324,N_37349,N_38693);
nand U46325 (N_46325,N_39734,N_35061);
or U46326 (N_46326,N_38255,N_30370);
and U46327 (N_46327,N_34973,N_32864);
xor U46328 (N_46328,N_31740,N_31193);
nand U46329 (N_46329,N_35593,N_34055);
xor U46330 (N_46330,N_30236,N_39771);
xor U46331 (N_46331,N_32733,N_31866);
and U46332 (N_46332,N_31173,N_39122);
xnor U46333 (N_46333,N_33746,N_30490);
and U46334 (N_46334,N_30604,N_38272);
nand U46335 (N_46335,N_34370,N_38244);
nand U46336 (N_46336,N_37895,N_37583);
and U46337 (N_46337,N_38182,N_39483);
and U46338 (N_46338,N_34982,N_32991);
xor U46339 (N_46339,N_32875,N_39060);
and U46340 (N_46340,N_30390,N_37531);
and U46341 (N_46341,N_38565,N_34868);
or U46342 (N_46342,N_34699,N_38261);
or U46343 (N_46343,N_37513,N_35184);
nor U46344 (N_46344,N_39630,N_31016);
and U46345 (N_46345,N_33403,N_31639);
nor U46346 (N_46346,N_32020,N_30238);
or U46347 (N_46347,N_34899,N_37546);
nand U46348 (N_46348,N_30158,N_33224);
xor U46349 (N_46349,N_33413,N_34531);
and U46350 (N_46350,N_34691,N_32348);
nor U46351 (N_46351,N_36152,N_38627);
or U46352 (N_46352,N_37396,N_39106);
nor U46353 (N_46353,N_38182,N_31834);
nor U46354 (N_46354,N_33571,N_32675);
xor U46355 (N_46355,N_31680,N_32049);
or U46356 (N_46356,N_38383,N_35271);
nand U46357 (N_46357,N_34729,N_38817);
and U46358 (N_46358,N_36135,N_32762);
nor U46359 (N_46359,N_30994,N_37950);
nand U46360 (N_46360,N_36101,N_38221);
or U46361 (N_46361,N_31328,N_33384);
or U46362 (N_46362,N_31939,N_37260);
and U46363 (N_46363,N_37812,N_32579);
nand U46364 (N_46364,N_32304,N_33214);
nand U46365 (N_46365,N_39273,N_35435);
xnor U46366 (N_46366,N_33671,N_31928);
or U46367 (N_46367,N_36625,N_37578);
nor U46368 (N_46368,N_34137,N_39249);
and U46369 (N_46369,N_39989,N_38850);
nand U46370 (N_46370,N_30862,N_34753);
nand U46371 (N_46371,N_37976,N_32633);
nand U46372 (N_46372,N_30173,N_38764);
xnor U46373 (N_46373,N_35426,N_30230);
and U46374 (N_46374,N_30083,N_38729);
xor U46375 (N_46375,N_35767,N_31748);
or U46376 (N_46376,N_36623,N_35016);
nor U46377 (N_46377,N_30468,N_39971);
nand U46378 (N_46378,N_32256,N_31383);
or U46379 (N_46379,N_32551,N_30071);
xor U46380 (N_46380,N_38958,N_30510);
nor U46381 (N_46381,N_34325,N_38040);
nor U46382 (N_46382,N_33571,N_30985);
nand U46383 (N_46383,N_30440,N_33262);
xnor U46384 (N_46384,N_32265,N_35852);
or U46385 (N_46385,N_33424,N_35583);
or U46386 (N_46386,N_35086,N_35702);
nand U46387 (N_46387,N_31663,N_34265);
xnor U46388 (N_46388,N_35191,N_37941);
or U46389 (N_46389,N_33814,N_33022);
nand U46390 (N_46390,N_35502,N_31958);
nor U46391 (N_46391,N_31997,N_36628);
nor U46392 (N_46392,N_30981,N_31823);
nor U46393 (N_46393,N_33817,N_36499);
or U46394 (N_46394,N_32724,N_32545);
and U46395 (N_46395,N_32103,N_32835);
or U46396 (N_46396,N_35736,N_35413);
and U46397 (N_46397,N_30287,N_38607);
xnor U46398 (N_46398,N_33336,N_33558);
xnor U46399 (N_46399,N_38513,N_34107);
nor U46400 (N_46400,N_34111,N_38758);
nor U46401 (N_46401,N_30686,N_34932);
and U46402 (N_46402,N_30212,N_33630);
nor U46403 (N_46403,N_38131,N_35589);
nor U46404 (N_46404,N_38626,N_34998);
nor U46405 (N_46405,N_33669,N_30291);
or U46406 (N_46406,N_31748,N_31995);
xnor U46407 (N_46407,N_33539,N_31756);
nor U46408 (N_46408,N_36283,N_39773);
nand U46409 (N_46409,N_34304,N_35445);
or U46410 (N_46410,N_38184,N_36567);
nor U46411 (N_46411,N_35745,N_39006);
nand U46412 (N_46412,N_30782,N_33829);
and U46413 (N_46413,N_30781,N_34490);
or U46414 (N_46414,N_33775,N_32558);
nor U46415 (N_46415,N_39379,N_31722);
nor U46416 (N_46416,N_38363,N_39019);
or U46417 (N_46417,N_36477,N_38869);
nand U46418 (N_46418,N_39862,N_31657);
or U46419 (N_46419,N_39114,N_31355);
or U46420 (N_46420,N_37564,N_37828);
xor U46421 (N_46421,N_37210,N_34353);
and U46422 (N_46422,N_33024,N_32232);
or U46423 (N_46423,N_31493,N_32341);
and U46424 (N_46424,N_31850,N_33253);
nor U46425 (N_46425,N_31630,N_38263);
and U46426 (N_46426,N_37571,N_31819);
xor U46427 (N_46427,N_39160,N_37109);
or U46428 (N_46428,N_32117,N_30639);
nand U46429 (N_46429,N_39061,N_33217);
and U46430 (N_46430,N_37081,N_39489);
nor U46431 (N_46431,N_32616,N_31512);
nor U46432 (N_46432,N_37097,N_37426);
nor U46433 (N_46433,N_30112,N_34542);
and U46434 (N_46434,N_36731,N_35700);
and U46435 (N_46435,N_38516,N_33350);
nand U46436 (N_46436,N_36137,N_31186);
nand U46437 (N_46437,N_31152,N_37241);
nor U46438 (N_46438,N_30304,N_34934);
nand U46439 (N_46439,N_33690,N_39290);
nand U46440 (N_46440,N_36269,N_36673);
and U46441 (N_46441,N_35403,N_35529);
xor U46442 (N_46442,N_38981,N_37036);
xnor U46443 (N_46443,N_31034,N_38575);
nand U46444 (N_46444,N_33951,N_35978);
xnor U46445 (N_46445,N_34859,N_31987);
xor U46446 (N_46446,N_35937,N_32523);
or U46447 (N_46447,N_30139,N_33767);
xor U46448 (N_46448,N_37433,N_34623);
and U46449 (N_46449,N_36648,N_30613);
nand U46450 (N_46450,N_35092,N_37577);
nor U46451 (N_46451,N_33390,N_38892);
xnor U46452 (N_46452,N_37105,N_39807);
and U46453 (N_46453,N_39958,N_35153);
or U46454 (N_46454,N_33405,N_36933);
or U46455 (N_46455,N_39342,N_30946);
or U46456 (N_46456,N_31648,N_38457);
or U46457 (N_46457,N_36360,N_33325);
or U46458 (N_46458,N_35712,N_35351);
xnor U46459 (N_46459,N_31699,N_30694);
xnor U46460 (N_46460,N_31419,N_35152);
and U46461 (N_46461,N_34881,N_31060);
nand U46462 (N_46462,N_35532,N_32710);
or U46463 (N_46463,N_36981,N_35906);
nor U46464 (N_46464,N_31979,N_38520);
and U46465 (N_46465,N_33432,N_36413);
nor U46466 (N_46466,N_32914,N_37795);
or U46467 (N_46467,N_30084,N_37324);
and U46468 (N_46468,N_33078,N_36057);
and U46469 (N_46469,N_37240,N_39962);
nor U46470 (N_46470,N_32122,N_34255);
and U46471 (N_46471,N_32658,N_39222);
nor U46472 (N_46472,N_35521,N_31369);
nand U46473 (N_46473,N_39796,N_31573);
xor U46474 (N_46474,N_37847,N_36847);
and U46475 (N_46475,N_39975,N_34182);
nor U46476 (N_46476,N_30554,N_35603);
nor U46477 (N_46477,N_39668,N_32435);
or U46478 (N_46478,N_30292,N_33680);
nand U46479 (N_46479,N_32536,N_36008);
nor U46480 (N_46480,N_35255,N_31410);
and U46481 (N_46481,N_30894,N_39856);
nand U46482 (N_46482,N_30391,N_32530);
and U46483 (N_46483,N_31705,N_33213);
and U46484 (N_46484,N_31687,N_37491);
xor U46485 (N_46485,N_37719,N_35257);
or U46486 (N_46486,N_31770,N_30624);
nor U46487 (N_46487,N_37419,N_35119);
and U46488 (N_46488,N_38646,N_30368);
or U46489 (N_46489,N_34966,N_37275);
nor U46490 (N_46490,N_39896,N_31319);
or U46491 (N_46491,N_38643,N_38406);
nand U46492 (N_46492,N_31778,N_31037);
nor U46493 (N_46493,N_31314,N_39525);
xor U46494 (N_46494,N_30139,N_37951);
xnor U46495 (N_46495,N_31182,N_37746);
nand U46496 (N_46496,N_33703,N_31455);
or U46497 (N_46497,N_34586,N_34115);
xnor U46498 (N_46498,N_35098,N_36142);
or U46499 (N_46499,N_34457,N_36025);
nand U46500 (N_46500,N_30807,N_33052);
nor U46501 (N_46501,N_36232,N_33407);
xor U46502 (N_46502,N_32046,N_30175);
and U46503 (N_46503,N_31812,N_32298);
or U46504 (N_46504,N_38002,N_38233);
nand U46505 (N_46505,N_35419,N_34445);
nor U46506 (N_46506,N_39471,N_32501);
xor U46507 (N_46507,N_30548,N_33303);
or U46508 (N_46508,N_35994,N_34620);
nor U46509 (N_46509,N_30103,N_33605);
nand U46510 (N_46510,N_33617,N_35380);
xnor U46511 (N_46511,N_39604,N_35880);
nor U46512 (N_46512,N_30081,N_37688);
xor U46513 (N_46513,N_39322,N_37321);
and U46514 (N_46514,N_38239,N_30795);
xor U46515 (N_46515,N_34606,N_32075);
and U46516 (N_46516,N_32065,N_30279);
xor U46517 (N_46517,N_32779,N_35556);
and U46518 (N_46518,N_32820,N_32253);
nand U46519 (N_46519,N_38337,N_30843);
xnor U46520 (N_46520,N_38488,N_34590);
xnor U46521 (N_46521,N_38113,N_31433);
and U46522 (N_46522,N_37616,N_39639);
nand U46523 (N_46523,N_33065,N_36657);
or U46524 (N_46524,N_32933,N_31875);
and U46525 (N_46525,N_35784,N_37803);
nor U46526 (N_46526,N_39867,N_32417);
nand U46527 (N_46527,N_33601,N_39304);
nor U46528 (N_46528,N_34419,N_37335);
and U46529 (N_46529,N_37942,N_37346);
and U46530 (N_46530,N_35857,N_30370);
xor U46531 (N_46531,N_31412,N_34531);
nor U46532 (N_46532,N_35487,N_33917);
nor U46533 (N_46533,N_37610,N_37798);
or U46534 (N_46534,N_30442,N_32236);
nor U46535 (N_46535,N_33352,N_38924);
nor U46536 (N_46536,N_37662,N_34289);
xor U46537 (N_46537,N_36937,N_38410);
and U46538 (N_46538,N_36410,N_36793);
nor U46539 (N_46539,N_30506,N_32353);
and U46540 (N_46540,N_35153,N_30147);
and U46541 (N_46541,N_37377,N_36728);
and U46542 (N_46542,N_38781,N_36426);
xor U46543 (N_46543,N_34445,N_31642);
nor U46544 (N_46544,N_32449,N_33821);
xor U46545 (N_46545,N_30454,N_37727);
and U46546 (N_46546,N_31658,N_30736);
nor U46547 (N_46547,N_38901,N_35637);
or U46548 (N_46548,N_38417,N_37263);
nand U46549 (N_46549,N_37387,N_35889);
or U46550 (N_46550,N_33023,N_36490);
nor U46551 (N_46551,N_32090,N_32044);
xor U46552 (N_46552,N_31306,N_31340);
nor U46553 (N_46553,N_35262,N_39972);
or U46554 (N_46554,N_30762,N_34897);
xor U46555 (N_46555,N_38855,N_30903);
nand U46556 (N_46556,N_32041,N_32159);
and U46557 (N_46557,N_36081,N_36306);
xor U46558 (N_46558,N_38699,N_32549);
and U46559 (N_46559,N_34701,N_38162);
xor U46560 (N_46560,N_32215,N_34325);
nor U46561 (N_46561,N_33042,N_37402);
or U46562 (N_46562,N_32498,N_38399);
nor U46563 (N_46563,N_33423,N_38578);
or U46564 (N_46564,N_39522,N_34962);
nand U46565 (N_46565,N_32560,N_36322);
nor U46566 (N_46566,N_37890,N_35163);
nor U46567 (N_46567,N_30957,N_31099);
nand U46568 (N_46568,N_35243,N_36923);
nor U46569 (N_46569,N_30715,N_34084);
nor U46570 (N_46570,N_39758,N_32357);
nor U46571 (N_46571,N_36708,N_30249);
or U46572 (N_46572,N_36167,N_32365);
nor U46573 (N_46573,N_32003,N_32763);
nand U46574 (N_46574,N_38543,N_36220);
nand U46575 (N_46575,N_36318,N_38573);
and U46576 (N_46576,N_36704,N_30295);
and U46577 (N_46577,N_37534,N_37666);
xnor U46578 (N_46578,N_33636,N_38495);
or U46579 (N_46579,N_37599,N_36172);
or U46580 (N_46580,N_34566,N_38857);
and U46581 (N_46581,N_30845,N_34052);
xnor U46582 (N_46582,N_35632,N_31782);
nor U46583 (N_46583,N_39975,N_39436);
and U46584 (N_46584,N_37614,N_36177);
and U46585 (N_46585,N_30260,N_33870);
xor U46586 (N_46586,N_30675,N_39204);
nor U46587 (N_46587,N_30823,N_32236);
and U46588 (N_46588,N_32045,N_31163);
xnor U46589 (N_46589,N_36942,N_31143);
and U46590 (N_46590,N_34384,N_39966);
xor U46591 (N_46591,N_36355,N_30506);
and U46592 (N_46592,N_35919,N_36889);
and U46593 (N_46593,N_38138,N_38286);
xor U46594 (N_46594,N_37311,N_33080);
nor U46595 (N_46595,N_30513,N_36613);
nand U46596 (N_46596,N_32002,N_39245);
nand U46597 (N_46597,N_39982,N_34385);
and U46598 (N_46598,N_35660,N_36098);
nand U46599 (N_46599,N_31469,N_36867);
and U46600 (N_46600,N_33890,N_34629);
nand U46601 (N_46601,N_38071,N_33280);
and U46602 (N_46602,N_34127,N_31882);
nor U46603 (N_46603,N_34176,N_36769);
nand U46604 (N_46604,N_39518,N_34033);
and U46605 (N_46605,N_33845,N_39396);
nand U46606 (N_46606,N_30232,N_35690);
xnor U46607 (N_46607,N_36380,N_37557);
nor U46608 (N_46608,N_33749,N_36170);
nand U46609 (N_46609,N_30278,N_31736);
and U46610 (N_46610,N_31505,N_31785);
and U46611 (N_46611,N_37872,N_32483);
nand U46612 (N_46612,N_34060,N_30518);
nor U46613 (N_46613,N_36724,N_31586);
xnor U46614 (N_46614,N_37438,N_30298);
xor U46615 (N_46615,N_30431,N_34264);
nand U46616 (N_46616,N_33903,N_34934);
nor U46617 (N_46617,N_38429,N_35032);
and U46618 (N_46618,N_31369,N_37082);
nor U46619 (N_46619,N_38144,N_36198);
or U46620 (N_46620,N_37422,N_32397);
nand U46621 (N_46621,N_33858,N_36818);
xnor U46622 (N_46622,N_31153,N_32773);
or U46623 (N_46623,N_30047,N_30799);
nor U46624 (N_46624,N_34986,N_31627);
and U46625 (N_46625,N_36093,N_39039);
nand U46626 (N_46626,N_31394,N_37798);
or U46627 (N_46627,N_35413,N_34854);
xnor U46628 (N_46628,N_37790,N_35487);
nor U46629 (N_46629,N_35889,N_32739);
or U46630 (N_46630,N_30898,N_36618);
nor U46631 (N_46631,N_35547,N_32478);
xor U46632 (N_46632,N_34196,N_37386);
nand U46633 (N_46633,N_32593,N_32273);
xor U46634 (N_46634,N_37499,N_34133);
nand U46635 (N_46635,N_38758,N_30408);
and U46636 (N_46636,N_30752,N_30033);
and U46637 (N_46637,N_34117,N_38696);
or U46638 (N_46638,N_31285,N_38544);
xor U46639 (N_46639,N_37817,N_31458);
or U46640 (N_46640,N_35633,N_38843);
nor U46641 (N_46641,N_33915,N_35610);
or U46642 (N_46642,N_33976,N_32458);
or U46643 (N_46643,N_38502,N_34135);
xor U46644 (N_46644,N_38176,N_39868);
xnor U46645 (N_46645,N_33901,N_31628);
and U46646 (N_46646,N_31224,N_35195);
nor U46647 (N_46647,N_37720,N_35680);
or U46648 (N_46648,N_32612,N_39947);
or U46649 (N_46649,N_39059,N_33580);
nand U46650 (N_46650,N_39949,N_35387);
nor U46651 (N_46651,N_30423,N_38585);
nand U46652 (N_46652,N_30332,N_30321);
and U46653 (N_46653,N_39194,N_33671);
or U46654 (N_46654,N_32632,N_33181);
xnor U46655 (N_46655,N_35670,N_30963);
and U46656 (N_46656,N_35699,N_39669);
nand U46657 (N_46657,N_32050,N_36807);
and U46658 (N_46658,N_32156,N_32289);
and U46659 (N_46659,N_30415,N_31437);
nand U46660 (N_46660,N_33713,N_33310);
nand U46661 (N_46661,N_34668,N_31141);
or U46662 (N_46662,N_31676,N_35549);
nor U46663 (N_46663,N_37240,N_38751);
or U46664 (N_46664,N_35019,N_33169);
and U46665 (N_46665,N_33908,N_35305);
xnor U46666 (N_46666,N_33180,N_33616);
or U46667 (N_46667,N_32434,N_30358);
nand U46668 (N_46668,N_34690,N_39090);
and U46669 (N_46669,N_36517,N_35195);
and U46670 (N_46670,N_30294,N_38911);
nor U46671 (N_46671,N_37980,N_31948);
nor U46672 (N_46672,N_32346,N_38158);
or U46673 (N_46673,N_34888,N_32680);
or U46674 (N_46674,N_31789,N_35385);
or U46675 (N_46675,N_35965,N_38667);
nor U46676 (N_46676,N_34425,N_38127);
nand U46677 (N_46677,N_33730,N_35986);
nor U46678 (N_46678,N_30418,N_31695);
and U46679 (N_46679,N_37307,N_38739);
nor U46680 (N_46680,N_35632,N_39983);
and U46681 (N_46681,N_38596,N_37397);
or U46682 (N_46682,N_32096,N_39270);
xnor U46683 (N_46683,N_32482,N_30650);
xor U46684 (N_46684,N_33207,N_35650);
xnor U46685 (N_46685,N_37317,N_37387);
xnor U46686 (N_46686,N_33081,N_32307);
nand U46687 (N_46687,N_39384,N_36232);
xnor U46688 (N_46688,N_31267,N_37374);
and U46689 (N_46689,N_37049,N_38830);
xor U46690 (N_46690,N_30253,N_38956);
nand U46691 (N_46691,N_34924,N_35962);
xor U46692 (N_46692,N_31362,N_38590);
nor U46693 (N_46693,N_30823,N_36894);
xnor U46694 (N_46694,N_32168,N_39472);
nand U46695 (N_46695,N_36598,N_39731);
and U46696 (N_46696,N_39841,N_39679);
or U46697 (N_46697,N_39200,N_39227);
nor U46698 (N_46698,N_32109,N_32219);
nand U46699 (N_46699,N_31300,N_33114);
nand U46700 (N_46700,N_30277,N_30856);
nand U46701 (N_46701,N_30806,N_31962);
nor U46702 (N_46702,N_33618,N_32312);
xor U46703 (N_46703,N_35933,N_37829);
and U46704 (N_46704,N_35419,N_34354);
nand U46705 (N_46705,N_33559,N_31042);
or U46706 (N_46706,N_37812,N_39149);
or U46707 (N_46707,N_39410,N_30435);
nor U46708 (N_46708,N_34424,N_31443);
nand U46709 (N_46709,N_34221,N_37751);
xor U46710 (N_46710,N_30682,N_33483);
nor U46711 (N_46711,N_33410,N_30301);
nor U46712 (N_46712,N_39147,N_31349);
nor U46713 (N_46713,N_35919,N_35891);
nor U46714 (N_46714,N_35625,N_38259);
or U46715 (N_46715,N_38717,N_37955);
nor U46716 (N_46716,N_35873,N_38759);
nor U46717 (N_46717,N_38403,N_38516);
or U46718 (N_46718,N_36390,N_33024);
and U46719 (N_46719,N_31972,N_34053);
nand U46720 (N_46720,N_37407,N_33799);
or U46721 (N_46721,N_36865,N_30980);
or U46722 (N_46722,N_34786,N_39292);
nand U46723 (N_46723,N_36168,N_35660);
xnor U46724 (N_46724,N_37517,N_30649);
nand U46725 (N_46725,N_32477,N_38505);
xnor U46726 (N_46726,N_36792,N_35727);
or U46727 (N_46727,N_38353,N_30251);
nor U46728 (N_46728,N_38531,N_36664);
xnor U46729 (N_46729,N_38123,N_37514);
nor U46730 (N_46730,N_36517,N_37427);
nor U46731 (N_46731,N_35185,N_32863);
nand U46732 (N_46732,N_32894,N_37413);
nor U46733 (N_46733,N_37578,N_32276);
nand U46734 (N_46734,N_38077,N_35871);
or U46735 (N_46735,N_33130,N_31741);
nor U46736 (N_46736,N_31082,N_39832);
nor U46737 (N_46737,N_33359,N_38319);
and U46738 (N_46738,N_37424,N_36129);
nor U46739 (N_46739,N_32020,N_35738);
and U46740 (N_46740,N_30186,N_32226);
xnor U46741 (N_46741,N_38979,N_37473);
and U46742 (N_46742,N_34703,N_34896);
xnor U46743 (N_46743,N_33831,N_30759);
xor U46744 (N_46744,N_36848,N_37974);
or U46745 (N_46745,N_31041,N_36800);
nor U46746 (N_46746,N_35905,N_39275);
nand U46747 (N_46747,N_35675,N_37479);
nand U46748 (N_46748,N_39054,N_32176);
or U46749 (N_46749,N_38468,N_31610);
and U46750 (N_46750,N_37992,N_32792);
nand U46751 (N_46751,N_31232,N_32576);
or U46752 (N_46752,N_39957,N_37716);
or U46753 (N_46753,N_34633,N_34294);
nand U46754 (N_46754,N_33821,N_33076);
xor U46755 (N_46755,N_39576,N_30252);
nand U46756 (N_46756,N_32529,N_36151);
nor U46757 (N_46757,N_38863,N_33712);
nor U46758 (N_46758,N_39260,N_35315);
and U46759 (N_46759,N_36404,N_37177);
or U46760 (N_46760,N_32931,N_37597);
or U46761 (N_46761,N_38039,N_38431);
nand U46762 (N_46762,N_32471,N_35138);
and U46763 (N_46763,N_39542,N_30518);
and U46764 (N_46764,N_36815,N_32532);
xnor U46765 (N_46765,N_37772,N_34456);
or U46766 (N_46766,N_38978,N_33001);
nand U46767 (N_46767,N_33968,N_36198);
nor U46768 (N_46768,N_33039,N_37280);
or U46769 (N_46769,N_30858,N_35826);
nand U46770 (N_46770,N_34395,N_30962);
and U46771 (N_46771,N_33856,N_34895);
and U46772 (N_46772,N_31294,N_30143);
or U46773 (N_46773,N_36275,N_32348);
xor U46774 (N_46774,N_31568,N_32886);
xor U46775 (N_46775,N_34828,N_33549);
xnor U46776 (N_46776,N_35870,N_36358);
and U46777 (N_46777,N_39597,N_32423);
or U46778 (N_46778,N_38980,N_30162);
or U46779 (N_46779,N_35893,N_33553);
nand U46780 (N_46780,N_32321,N_38876);
nor U46781 (N_46781,N_37084,N_31399);
xnor U46782 (N_46782,N_33599,N_31632);
xnor U46783 (N_46783,N_39574,N_38854);
nor U46784 (N_46784,N_38618,N_38179);
nor U46785 (N_46785,N_35251,N_30636);
or U46786 (N_46786,N_32775,N_34503);
nand U46787 (N_46787,N_30157,N_32208);
nand U46788 (N_46788,N_33536,N_33939);
and U46789 (N_46789,N_35326,N_34231);
nor U46790 (N_46790,N_37394,N_30339);
or U46791 (N_46791,N_33543,N_36170);
nand U46792 (N_46792,N_30664,N_30892);
and U46793 (N_46793,N_37127,N_32107);
xor U46794 (N_46794,N_31204,N_36883);
xor U46795 (N_46795,N_36734,N_37266);
or U46796 (N_46796,N_31379,N_37223);
nor U46797 (N_46797,N_39885,N_38410);
nand U46798 (N_46798,N_34179,N_30532);
or U46799 (N_46799,N_32088,N_31453);
nor U46800 (N_46800,N_36020,N_36747);
or U46801 (N_46801,N_36539,N_33126);
nor U46802 (N_46802,N_38774,N_33245);
xnor U46803 (N_46803,N_34645,N_31139);
xor U46804 (N_46804,N_31791,N_39135);
nand U46805 (N_46805,N_38105,N_32904);
xnor U46806 (N_46806,N_32837,N_30978);
nor U46807 (N_46807,N_31455,N_39080);
nor U46808 (N_46808,N_36652,N_30718);
and U46809 (N_46809,N_34393,N_39348);
or U46810 (N_46810,N_31393,N_38093);
nand U46811 (N_46811,N_37922,N_32497);
nor U46812 (N_46812,N_38782,N_32174);
or U46813 (N_46813,N_36494,N_30841);
nor U46814 (N_46814,N_32809,N_32930);
or U46815 (N_46815,N_37879,N_36796);
xor U46816 (N_46816,N_38858,N_31890);
or U46817 (N_46817,N_32099,N_33244);
xor U46818 (N_46818,N_32410,N_39806);
xor U46819 (N_46819,N_38592,N_35834);
nand U46820 (N_46820,N_39318,N_30820);
and U46821 (N_46821,N_35847,N_39940);
nor U46822 (N_46822,N_30964,N_31497);
nor U46823 (N_46823,N_38239,N_38134);
xor U46824 (N_46824,N_36616,N_37808);
nand U46825 (N_46825,N_36669,N_31267);
or U46826 (N_46826,N_36314,N_34011);
nand U46827 (N_46827,N_31195,N_39171);
and U46828 (N_46828,N_37139,N_33875);
nor U46829 (N_46829,N_33467,N_37343);
or U46830 (N_46830,N_38960,N_34292);
or U46831 (N_46831,N_31395,N_33407);
or U46832 (N_46832,N_37875,N_38920);
nand U46833 (N_46833,N_38314,N_39244);
nand U46834 (N_46834,N_39352,N_39224);
or U46835 (N_46835,N_30124,N_33677);
and U46836 (N_46836,N_30979,N_36980);
or U46837 (N_46837,N_38076,N_33291);
xor U46838 (N_46838,N_31476,N_31041);
or U46839 (N_46839,N_36342,N_35923);
nand U46840 (N_46840,N_38468,N_38540);
xnor U46841 (N_46841,N_34999,N_32871);
nor U46842 (N_46842,N_38500,N_37486);
nor U46843 (N_46843,N_30859,N_37587);
nand U46844 (N_46844,N_33287,N_31689);
or U46845 (N_46845,N_33289,N_32488);
xnor U46846 (N_46846,N_39639,N_35255);
xor U46847 (N_46847,N_30024,N_32185);
xor U46848 (N_46848,N_32096,N_33364);
nor U46849 (N_46849,N_30636,N_31292);
xor U46850 (N_46850,N_30386,N_36724);
xnor U46851 (N_46851,N_36581,N_33808);
xnor U46852 (N_46852,N_32847,N_34299);
nor U46853 (N_46853,N_38310,N_31942);
and U46854 (N_46854,N_37754,N_31930);
nand U46855 (N_46855,N_37813,N_36442);
and U46856 (N_46856,N_38188,N_30306);
or U46857 (N_46857,N_34555,N_31627);
nand U46858 (N_46858,N_33896,N_39384);
or U46859 (N_46859,N_34140,N_30816);
xor U46860 (N_46860,N_32457,N_36282);
nand U46861 (N_46861,N_31072,N_37009);
nand U46862 (N_46862,N_32764,N_37357);
nand U46863 (N_46863,N_30819,N_35160);
nor U46864 (N_46864,N_38307,N_39499);
nand U46865 (N_46865,N_34832,N_34084);
xnor U46866 (N_46866,N_38891,N_31213);
or U46867 (N_46867,N_39739,N_38513);
nand U46868 (N_46868,N_36657,N_39715);
and U46869 (N_46869,N_31146,N_32134);
nand U46870 (N_46870,N_30285,N_30706);
nor U46871 (N_46871,N_33274,N_35081);
or U46872 (N_46872,N_35997,N_36226);
nor U46873 (N_46873,N_30776,N_37764);
and U46874 (N_46874,N_39864,N_39673);
and U46875 (N_46875,N_37457,N_39644);
nor U46876 (N_46876,N_39278,N_35550);
or U46877 (N_46877,N_37465,N_38089);
nor U46878 (N_46878,N_30562,N_32413);
nor U46879 (N_46879,N_30697,N_30239);
nand U46880 (N_46880,N_33832,N_37035);
and U46881 (N_46881,N_35500,N_32271);
xor U46882 (N_46882,N_39684,N_31789);
or U46883 (N_46883,N_35956,N_35656);
xnor U46884 (N_46884,N_38720,N_31601);
and U46885 (N_46885,N_33112,N_32164);
or U46886 (N_46886,N_34085,N_35440);
and U46887 (N_46887,N_33590,N_31259);
xnor U46888 (N_46888,N_35581,N_34034);
nand U46889 (N_46889,N_39944,N_36684);
and U46890 (N_46890,N_36166,N_37518);
nand U46891 (N_46891,N_33860,N_33811);
nor U46892 (N_46892,N_35280,N_33975);
and U46893 (N_46893,N_33531,N_36653);
nand U46894 (N_46894,N_34354,N_38195);
or U46895 (N_46895,N_32804,N_38702);
or U46896 (N_46896,N_34317,N_37513);
or U46897 (N_46897,N_36223,N_33781);
or U46898 (N_46898,N_30534,N_32198);
xnor U46899 (N_46899,N_34563,N_36957);
xor U46900 (N_46900,N_32090,N_35451);
or U46901 (N_46901,N_34074,N_31969);
and U46902 (N_46902,N_38853,N_36037);
nor U46903 (N_46903,N_32129,N_36207);
and U46904 (N_46904,N_35479,N_35364);
xnor U46905 (N_46905,N_38529,N_37030);
xor U46906 (N_46906,N_38860,N_35198);
nor U46907 (N_46907,N_30995,N_32324);
xor U46908 (N_46908,N_37070,N_30739);
xnor U46909 (N_46909,N_33281,N_34298);
and U46910 (N_46910,N_33778,N_32217);
or U46911 (N_46911,N_35686,N_31647);
and U46912 (N_46912,N_39435,N_35228);
or U46913 (N_46913,N_36003,N_37083);
xor U46914 (N_46914,N_37822,N_37743);
nand U46915 (N_46915,N_34228,N_37900);
nor U46916 (N_46916,N_34506,N_34549);
and U46917 (N_46917,N_32061,N_37991);
and U46918 (N_46918,N_30222,N_32198);
and U46919 (N_46919,N_31349,N_36660);
xor U46920 (N_46920,N_33227,N_32604);
nor U46921 (N_46921,N_33654,N_32356);
xnor U46922 (N_46922,N_39897,N_35978);
xor U46923 (N_46923,N_36639,N_30105);
nand U46924 (N_46924,N_38060,N_33807);
nand U46925 (N_46925,N_35049,N_33350);
and U46926 (N_46926,N_33080,N_37880);
nor U46927 (N_46927,N_38498,N_37998);
xor U46928 (N_46928,N_32264,N_32499);
nor U46929 (N_46929,N_32027,N_33476);
nand U46930 (N_46930,N_31425,N_33735);
nor U46931 (N_46931,N_39656,N_31797);
or U46932 (N_46932,N_30461,N_34525);
nor U46933 (N_46933,N_39926,N_37857);
and U46934 (N_46934,N_35783,N_37786);
and U46935 (N_46935,N_34174,N_33006);
nand U46936 (N_46936,N_30211,N_33799);
xor U46937 (N_46937,N_35172,N_37918);
nand U46938 (N_46938,N_34630,N_35496);
or U46939 (N_46939,N_31377,N_31584);
xnor U46940 (N_46940,N_31967,N_35161);
xor U46941 (N_46941,N_35754,N_31781);
xor U46942 (N_46942,N_34162,N_32397);
nor U46943 (N_46943,N_30176,N_35744);
nand U46944 (N_46944,N_37987,N_33978);
nor U46945 (N_46945,N_39358,N_31932);
and U46946 (N_46946,N_35880,N_38504);
or U46947 (N_46947,N_36297,N_35130);
xnor U46948 (N_46948,N_39689,N_30695);
or U46949 (N_46949,N_39492,N_32607);
xnor U46950 (N_46950,N_36308,N_36625);
nand U46951 (N_46951,N_32930,N_34315);
xor U46952 (N_46952,N_32559,N_35398);
nand U46953 (N_46953,N_37492,N_36993);
and U46954 (N_46954,N_34989,N_31363);
nor U46955 (N_46955,N_33208,N_33040);
nand U46956 (N_46956,N_31519,N_34244);
nand U46957 (N_46957,N_34813,N_38513);
xor U46958 (N_46958,N_30619,N_39932);
nand U46959 (N_46959,N_31706,N_37479);
nand U46960 (N_46960,N_33201,N_37576);
or U46961 (N_46961,N_31222,N_32001);
and U46962 (N_46962,N_31832,N_31653);
and U46963 (N_46963,N_37748,N_31799);
or U46964 (N_46964,N_39194,N_30212);
nor U46965 (N_46965,N_33105,N_37678);
nor U46966 (N_46966,N_38262,N_31379);
nand U46967 (N_46967,N_32107,N_37254);
xnor U46968 (N_46968,N_35518,N_38332);
xnor U46969 (N_46969,N_37117,N_34419);
or U46970 (N_46970,N_38445,N_32246);
nand U46971 (N_46971,N_33217,N_31430);
nand U46972 (N_46972,N_30260,N_31494);
nor U46973 (N_46973,N_33770,N_34532);
nor U46974 (N_46974,N_32743,N_38392);
nand U46975 (N_46975,N_38948,N_39571);
nor U46976 (N_46976,N_31760,N_35031);
nor U46977 (N_46977,N_39274,N_38795);
or U46978 (N_46978,N_35134,N_34278);
nand U46979 (N_46979,N_31240,N_37323);
xor U46980 (N_46980,N_30046,N_36355);
nand U46981 (N_46981,N_38704,N_30791);
nor U46982 (N_46982,N_38043,N_32794);
nor U46983 (N_46983,N_30478,N_37669);
or U46984 (N_46984,N_34651,N_39843);
nand U46985 (N_46985,N_30179,N_36566);
nor U46986 (N_46986,N_38329,N_38986);
xor U46987 (N_46987,N_36010,N_32333);
and U46988 (N_46988,N_37902,N_36598);
nor U46989 (N_46989,N_36674,N_36753);
or U46990 (N_46990,N_34436,N_34816);
and U46991 (N_46991,N_37789,N_32354);
and U46992 (N_46992,N_34091,N_33421);
nor U46993 (N_46993,N_32923,N_33059);
and U46994 (N_46994,N_31683,N_33328);
nand U46995 (N_46995,N_35439,N_31614);
or U46996 (N_46996,N_30991,N_32194);
and U46997 (N_46997,N_33147,N_37430);
nor U46998 (N_46998,N_30857,N_39456);
or U46999 (N_46999,N_37623,N_35183);
or U47000 (N_47000,N_38317,N_32948);
nor U47001 (N_47001,N_31184,N_35823);
and U47002 (N_47002,N_33669,N_31452);
nand U47003 (N_47003,N_38073,N_31787);
or U47004 (N_47004,N_36056,N_33682);
nand U47005 (N_47005,N_39542,N_30085);
nand U47006 (N_47006,N_33677,N_34625);
and U47007 (N_47007,N_35848,N_31070);
and U47008 (N_47008,N_36114,N_34810);
nand U47009 (N_47009,N_35531,N_31819);
nand U47010 (N_47010,N_32540,N_39125);
xor U47011 (N_47011,N_32529,N_37472);
nor U47012 (N_47012,N_34908,N_33438);
nor U47013 (N_47013,N_31171,N_37725);
and U47014 (N_47014,N_38582,N_34436);
xnor U47015 (N_47015,N_37726,N_36264);
nor U47016 (N_47016,N_39668,N_30069);
xnor U47017 (N_47017,N_33730,N_35727);
nor U47018 (N_47018,N_36064,N_37412);
nor U47019 (N_47019,N_38506,N_37333);
nor U47020 (N_47020,N_38705,N_33762);
xnor U47021 (N_47021,N_31012,N_30089);
xnor U47022 (N_47022,N_30408,N_38641);
nand U47023 (N_47023,N_32097,N_36644);
or U47024 (N_47024,N_31958,N_31980);
nand U47025 (N_47025,N_38753,N_37381);
nor U47026 (N_47026,N_31503,N_30459);
nand U47027 (N_47027,N_38381,N_38300);
or U47028 (N_47028,N_31824,N_39388);
or U47029 (N_47029,N_38172,N_33763);
nand U47030 (N_47030,N_36191,N_34269);
nor U47031 (N_47031,N_37998,N_30321);
or U47032 (N_47032,N_35946,N_32612);
xor U47033 (N_47033,N_38459,N_37730);
or U47034 (N_47034,N_38982,N_39928);
xnor U47035 (N_47035,N_36096,N_39372);
nor U47036 (N_47036,N_30799,N_33778);
and U47037 (N_47037,N_37006,N_36813);
or U47038 (N_47038,N_32679,N_36901);
xnor U47039 (N_47039,N_34673,N_38844);
or U47040 (N_47040,N_34297,N_38201);
and U47041 (N_47041,N_33807,N_30227);
nand U47042 (N_47042,N_37974,N_31673);
nand U47043 (N_47043,N_35362,N_33977);
nor U47044 (N_47044,N_38979,N_30474);
and U47045 (N_47045,N_30138,N_38109);
and U47046 (N_47046,N_33019,N_34842);
xor U47047 (N_47047,N_38109,N_39360);
nor U47048 (N_47048,N_33136,N_34817);
nand U47049 (N_47049,N_36451,N_39628);
xor U47050 (N_47050,N_38429,N_37156);
xnor U47051 (N_47051,N_33026,N_31435);
or U47052 (N_47052,N_35286,N_33444);
or U47053 (N_47053,N_35003,N_33002);
or U47054 (N_47054,N_33669,N_31736);
xor U47055 (N_47055,N_30284,N_31051);
nand U47056 (N_47056,N_32127,N_30506);
xnor U47057 (N_47057,N_31238,N_31824);
nand U47058 (N_47058,N_39978,N_34611);
xnor U47059 (N_47059,N_33036,N_33096);
and U47060 (N_47060,N_32233,N_38736);
nand U47061 (N_47061,N_37053,N_37231);
or U47062 (N_47062,N_31024,N_36922);
or U47063 (N_47063,N_33998,N_35752);
xnor U47064 (N_47064,N_33819,N_35089);
nand U47065 (N_47065,N_35202,N_31511);
nor U47066 (N_47066,N_37313,N_39942);
nand U47067 (N_47067,N_32370,N_33747);
xnor U47068 (N_47068,N_32662,N_37553);
nor U47069 (N_47069,N_32493,N_36783);
nor U47070 (N_47070,N_39781,N_39403);
and U47071 (N_47071,N_36173,N_31407);
nand U47072 (N_47072,N_38334,N_39270);
xnor U47073 (N_47073,N_33642,N_39207);
or U47074 (N_47074,N_31487,N_30605);
nor U47075 (N_47075,N_32819,N_36074);
or U47076 (N_47076,N_39964,N_39593);
or U47077 (N_47077,N_31256,N_38340);
nor U47078 (N_47078,N_31114,N_37742);
nor U47079 (N_47079,N_38358,N_33490);
or U47080 (N_47080,N_32666,N_33585);
nor U47081 (N_47081,N_35737,N_32430);
or U47082 (N_47082,N_37996,N_39349);
and U47083 (N_47083,N_39026,N_38507);
or U47084 (N_47084,N_38052,N_36674);
and U47085 (N_47085,N_30981,N_32247);
nor U47086 (N_47086,N_36999,N_35678);
and U47087 (N_47087,N_31135,N_38462);
nand U47088 (N_47088,N_33336,N_33636);
or U47089 (N_47089,N_38773,N_32791);
nor U47090 (N_47090,N_31755,N_35033);
xnor U47091 (N_47091,N_35618,N_36525);
xnor U47092 (N_47092,N_39033,N_36925);
nor U47093 (N_47093,N_34826,N_32597);
nor U47094 (N_47094,N_33456,N_34162);
nor U47095 (N_47095,N_31414,N_36394);
xnor U47096 (N_47096,N_34090,N_32088);
nor U47097 (N_47097,N_36641,N_34653);
nand U47098 (N_47098,N_39422,N_35798);
or U47099 (N_47099,N_36169,N_30657);
xnor U47100 (N_47100,N_32737,N_34125);
xnor U47101 (N_47101,N_32890,N_35421);
or U47102 (N_47102,N_31419,N_32804);
nand U47103 (N_47103,N_32099,N_36594);
nand U47104 (N_47104,N_30810,N_32645);
or U47105 (N_47105,N_31033,N_31481);
nand U47106 (N_47106,N_30011,N_31227);
nor U47107 (N_47107,N_34736,N_37776);
nand U47108 (N_47108,N_30424,N_33946);
xor U47109 (N_47109,N_31309,N_37802);
and U47110 (N_47110,N_34165,N_37007);
and U47111 (N_47111,N_38831,N_34775);
nand U47112 (N_47112,N_30654,N_35744);
nor U47113 (N_47113,N_32161,N_37592);
and U47114 (N_47114,N_37957,N_30768);
nand U47115 (N_47115,N_31477,N_35075);
and U47116 (N_47116,N_33801,N_33000);
nor U47117 (N_47117,N_31124,N_36193);
or U47118 (N_47118,N_32519,N_39494);
or U47119 (N_47119,N_37437,N_34493);
nand U47120 (N_47120,N_34247,N_32076);
nand U47121 (N_47121,N_33830,N_30345);
nand U47122 (N_47122,N_37363,N_35655);
or U47123 (N_47123,N_34670,N_37771);
or U47124 (N_47124,N_34011,N_36733);
or U47125 (N_47125,N_39180,N_38067);
nand U47126 (N_47126,N_34907,N_35088);
and U47127 (N_47127,N_30129,N_30533);
nor U47128 (N_47128,N_32721,N_35129);
nand U47129 (N_47129,N_32555,N_39579);
or U47130 (N_47130,N_36768,N_36714);
nor U47131 (N_47131,N_36774,N_31013);
xnor U47132 (N_47132,N_32034,N_39975);
nor U47133 (N_47133,N_31827,N_36880);
or U47134 (N_47134,N_35369,N_35100);
xor U47135 (N_47135,N_34493,N_37127);
xnor U47136 (N_47136,N_38704,N_35875);
xnor U47137 (N_47137,N_39756,N_38944);
or U47138 (N_47138,N_39120,N_30591);
nor U47139 (N_47139,N_33697,N_38528);
and U47140 (N_47140,N_36367,N_31888);
or U47141 (N_47141,N_31963,N_38319);
nand U47142 (N_47142,N_30097,N_31693);
and U47143 (N_47143,N_34423,N_33236);
and U47144 (N_47144,N_35583,N_37131);
nand U47145 (N_47145,N_34811,N_30707);
and U47146 (N_47146,N_31930,N_30878);
nand U47147 (N_47147,N_33791,N_31139);
and U47148 (N_47148,N_34601,N_30259);
nand U47149 (N_47149,N_35948,N_37308);
nand U47150 (N_47150,N_36399,N_33818);
xor U47151 (N_47151,N_32340,N_32566);
nand U47152 (N_47152,N_31629,N_34801);
or U47153 (N_47153,N_31171,N_37442);
nor U47154 (N_47154,N_38137,N_34307);
or U47155 (N_47155,N_35470,N_33778);
nor U47156 (N_47156,N_35092,N_37980);
nor U47157 (N_47157,N_34449,N_38064);
and U47158 (N_47158,N_37597,N_30569);
and U47159 (N_47159,N_37886,N_32530);
nand U47160 (N_47160,N_37367,N_37815);
nand U47161 (N_47161,N_32502,N_35869);
nand U47162 (N_47162,N_32916,N_30596);
nor U47163 (N_47163,N_32367,N_36859);
and U47164 (N_47164,N_30876,N_32760);
nor U47165 (N_47165,N_32796,N_39467);
nor U47166 (N_47166,N_37739,N_32822);
nor U47167 (N_47167,N_35809,N_35642);
nor U47168 (N_47168,N_31141,N_33482);
nor U47169 (N_47169,N_33798,N_35630);
nor U47170 (N_47170,N_35183,N_34113);
or U47171 (N_47171,N_37574,N_30673);
xor U47172 (N_47172,N_36143,N_31689);
xnor U47173 (N_47173,N_31786,N_38939);
or U47174 (N_47174,N_38127,N_33770);
nand U47175 (N_47175,N_32427,N_37697);
nor U47176 (N_47176,N_35477,N_39944);
or U47177 (N_47177,N_33128,N_34491);
nand U47178 (N_47178,N_37351,N_31495);
nand U47179 (N_47179,N_31197,N_31569);
xnor U47180 (N_47180,N_34380,N_38433);
and U47181 (N_47181,N_39328,N_35201);
nor U47182 (N_47182,N_39288,N_34963);
or U47183 (N_47183,N_34012,N_30372);
nor U47184 (N_47184,N_39849,N_30628);
nand U47185 (N_47185,N_35754,N_30865);
and U47186 (N_47186,N_32512,N_34728);
and U47187 (N_47187,N_31474,N_34081);
or U47188 (N_47188,N_33607,N_32046);
nand U47189 (N_47189,N_36609,N_39277);
nor U47190 (N_47190,N_35718,N_31018);
nand U47191 (N_47191,N_35399,N_33868);
nor U47192 (N_47192,N_37284,N_33254);
xnor U47193 (N_47193,N_33328,N_33349);
nor U47194 (N_47194,N_30122,N_30536);
or U47195 (N_47195,N_39076,N_35640);
or U47196 (N_47196,N_31069,N_30592);
or U47197 (N_47197,N_36042,N_37135);
nand U47198 (N_47198,N_37325,N_35419);
nand U47199 (N_47199,N_36752,N_34457);
xor U47200 (N_47200,N_34216,N_39889);
xnor U47201 (N_47201,N_30839,N_37746);
nor U47202 (N_47202,N_30294,N_30030);
or U47203 (N_47203,N_36894,N_36108);
nor U47204 (N_47204,N_32096,N_38945);
or U47205 (N_47205,N_33058,N_32389);
and U47206 (N_47206,N_37768,N_37847);
or U47207 (N_47207,N_37142,N_34141);
nand U47208 (N_47208,N_31439,N_39056);
or U47209 (N_47209,N_30812,N_39059);
xnor U47210 (N_47210,N_33238,N_38824);
or U47211 (N_47211,N_33233,N_34079);
nor U47212 (N_47212,N_32862,N_36452);
nor U47213 (N_47213,N_30555,N_38408);
or U47214 (N_47214,N_35714,N_32067);
and U47215 (N_47215,N_31792,N_35581);
and U47216 (N_47216,N_39527,N_38391);
nand U47217 (N_47217,N_33374,N_37006);
xor U47218 (N_47218,N_30425,N_35370);
nand U47219 (N_47219,N_36007,N_33197);
or U47220 (N_47220,N_30376,N_33464);
xor U47221 (N_47221,N_31575,N_32156);
nand U47222 (N_47222,N_33452,N_36974);
nand U47223 (N_47223,N_39414,N_32564);
nor U47224 (N_47224,N_36815,N_32920);
nor U47225 (N_47225,N_36835,N_30084);
nand U47226 (N_47226,N_33712,N_31205);
xnor U47227 (N_47227,N_36079,N_33047);
nand U47228 (N_47228,N_31690,N_34339);
nor U47229 (N_47229,N_31108,N_32928);
nor U47230 (N_47230,N_38876,N_37273);
or U47231 (N_47231,N_35722,N_33188);
nand U47232 (N_47232,N_34559,N_35407);
xor U47233 (N_47233,N_32181,N_34068);
and U47234 (N_47234,N_39764,N_36429);
xnor U47235 (N_47235,N_38011,N_36129);
nand U47236 (N_47236,N_31105,N_34008);
nand U47237 (N_47237,N_37172,N_36331);
or U47238 (N_47238,N_37745,N_38546);
nand U47239 (N_47239,N_34510,N_30588);
nor U47240 (N_47240,N_39958,N_36553);
or U47241 (N_47241,N_30567,N_35251);
xnor U47242 (N_47242,N_36401,N_39092);
or U47243 (N_47243,N_35640,N_30484);
nand U47244 (N_47244,N_39202,N_30991);
or U47245 (N_47245,N_38242,N_36912);
nor U47246 (N_47246,N_35131,N_32323);
and U47247 (N_47247,N_33229,N_31433);
nand U47248 (N_47248,N_33060,N_39773);
and U47249 (N_47249,N_36221,N_33477);
nand U47250 (N_47250,N_38952,N_35811);
xor U47251 (N_47251,N_32619,N_35164);
xnor U47252 (N_47252,N_34455,N_34258);
or U47253 (N_47253,N_34267,N_30429);
xor U47254 (N_47254,N_37401,N_36692);
xnor U47255 (N_47255,N_35785,N_32978);
and U47256 (N_47256,N_38407,N_30388);
xnor U47257 (N_47257,N_32258,N_32195);
nor U47258 (N_47258,N_38371,N_38036);
or U47259 (N_47259,N_36168,N_34147);
xnor U47260 (N_47260,N_31332,N_38436);
or U47261 (N_47261,N_30372,N_33712);
and U47262 (N_47262,N_35053,N_39611);
nand U47263 (N_47263,N_34587,N_31739);
nor U47264 (N_47264,N_37531,N_31806);
and U47265 (N_47265,N_36184,N_37689);
nand U47266 (N_47266,N_36432,N_34217);
xnor U47267 (N_47267,N_37039,N_35544);
nor U47268 (N_47268,N_31591,N_38218);
nand U47269 (N_47269,N_33735,N_30771);
xor U47270 (N_47270,N_37666,N_31148);
or U47271 (N_47271,N_31051,N_31676);
nand U47272 (N_47272,N_35088,N_37761);
and U47273 (N_47273,N_36922,N_37213);
nor U47274 (N_47274,N_30063,N_37792);
xnor U47275 (N_47275,N_33343,N_32856);
or U47276 (N_47276,N_30803,N_37865);
and U47277 (N_47277,N_31929,N_34629);
xor U47278 (N_47278,N_34142,N_33145);
xor U47279 (N_47279,N_35294,N_30748);
or U47280 (N_47280,N_33203,N_33840);
nand U47281 (N_47281,N_34463,N_32667);
or U47282 (N_47282,N_32184,N_35363);
or U47283 (N_47283,N_33186,N_31506);
nor U47284 (N_47284,N_33130,N_31206);
xor U47285 (N_47285,N_34547,N_34540);
or U47286 (N_47286,N_34334,N_37547);
xnor U47287 (N_47287,N_34449,N_30421);
and U47288 (N_47288,N_31943,N_38656);
and U47289 (N_47289,N_35691,N_37856);
and U47290 (N_47290,N_30823,N_37786);
nand U47291 (N_47291,N_33995,N_36213);
nor U47292 (N_47292,N_34737,N_38438);
nor U47293 (N_47293,N_34269,N_30583);
nand U47294 (N_47294,N_31071,N_32959);
and U47295 (N_47295,N_30225,N_36979);
xor U47296 (N_47296,N_31226,N_39830);
nand U47297 (N_47297,N_34433,N_39064);
and U47298 (N_47298,N_30394,N_36514);
nor U47299 (N_47299,N_32402,N_38116);
or U47300 (N_47300,N_34009,N_30448);
nand U47301 (N_47301,N_31893,N_34831);
nand U47302 (N_47302,N_37905,N_30187);
and U47303 (N_47303,N_33866,N_31537);
xor U47304 (N_47304,N_31965,N_37397);
nor U47305 (N_47305,N_31905,N_33373);
and U47306 (N_47306,N_37823,N_32980);
or U47307 (N_47307,N_38510,N_30244);
and U47308 (N_47308,N_33402,N_37754);
xor U47309 (N_47309,N_38078,N_35571);
or U47310 (N_47310,N_37530,N_37661);
xnor U47311 (N_47311,N_32484,N_30602);
or U47312 (N_47312,N_35124,N_35890);
or U47313 (N_47313,N_32901,N_34516);
and U47314 (N_47314,N_30158,N_31049);
xor U47315 (N_47315,N_35632,N_37569);
or U47316 (N_47316,N_34867,N_38187);
nand U47317 (N_47317,N_38432,N_33601);
nand U47318 (N_47318,N_33866,N_30268);
and U47319 (N_47319,N_36472,N_30044);
nor U47320 (N_47320,N_37579,N_31493);
nand U47321 (N_47321,N_39739,N_39230);
nor U47322 (N_47322,N_33819,N_32377);
xnor U47323 (N_47323,N_32651,N_32019);
nand U47324 (N_47324,N_35265,N_38001);
nor U47325 (N_47325,N_34085,N_32030);
xnor U47326 (N_47326,N_30160,N_31988);
nor U47327 (N_47327,N_37192,N_36182);
nand U47328 (N_47328,N_33194,N_39082);
xor U47329 (N_47329,N_36584,N_36614);
or U47330 (N_47330,N_38724,N_35025);
and U47331 (N_47331,N_36961,N_32001);
or U47332 (N_47332,N_37403,N_38363);
xor U47333 (N_47333,N_32162,N_31612);
xnor U47334 (N_47334,N_33028,N_33754);
nor U47335 (N_47335,N_31984,N_39434);
nand U47336 (N_47336,N_33105,N_36690);
or U47337 (N_47337,N_30996,N_34165);
and U47338 (N_47338,N_34318,N_38537);
xnor U47339 (N_47339,N_34527,N_30196);
and U47340 (N_47340,N_33352,N_33715);
nor U47341 (N_47341,N_36185,N_32162);
nand U47342 (N_47342,N_32698,N_30841);
nand U47343 (N_47343,N_35767,N_34180);
nand U47344 (N_47344,N_35752,N_38980);
or U47345 (N_47345,N_36662,N_33864);
and U47346 (N_47346,N_33479,N_33904);
xnor U47347 (N_47347,N_36053,N_32356);
nor U47348 (N_47348,N_31353,N_31578);
xor U47349 (N_47349,N_30123,N_34573);
or U47350 (N_47350,N_33729,N_34118);
xnor U47351 (N_47351,N_39822,N_33731);
xor U47352 (N_47352,N_31813,N_37116);
nand U47353 (N_47353,N_30437,N_31822);
nor U47354 (N_47354,N_31522,N_36932);
and U47355 (N_47355,N_30874,N_36318);
nand U47356 (N_47356,N_32552,N_31430);
nor U47357 (N_47357,N_30489,N_36868);
and U47358 (N_47358,N_33639,N_38188);
xor U47359 (N_47359,N_35166,N_35764);
xor U47360 (N_47360,N_33037,N_30105);
xnor U47361 (N_47361,N_30352,N_35821);
xor U47362 (N_47362,N_32526,N_36364);
or U47363 (N_47363,N_31559,N_36639);
nor U47364 (N_47364,N_39778,N_37613);
nor U47365 (N_47365,N_39643,N_31330);
xnor U47366 (N_47366,N_36121,N_34849);
or U47367 (N_47367,N_30818,N_30420);
nand U47368 (N_47368,N_33188,N_37403);
or U47369 (N_47369,N_39323,N_30512);
nor U47370 (N_47370,N_32496,N_32205);
and U47371 (N_47371,N_39218,N_38989);
nor U47372 (N_47372,N_39135,N_37785);
and U47373 (N_47373,N_33581,N_38221);
nor U47374 (N_47374,N_38917,N_39448);
nand U47375 (N_47375,N_33561,N_34115);
or U47376 (N_47376,N_30568,N_30406);
nand U47377 (N_47377,N_34794,N_32277);
or U47378 (N_47378,N_36646,N_35546);
or U47379 (N_47379,N_38133,N_33146);
nor U47380 (N_47380,N_39109,N_39410);
and U47381 (N_47381,N_30914,N_34490);
nor U47382 (N_47382,N_38334,N_30342);
or U47383 (N_47383,N_32666,N_31539);
and U47384 (N_47384,N_37744,N_32389);
nand U47385 (N_47385,N_38035,N_36321);
and U47386 (N_47386,N_33344,N_37776);
or U47387 (N_47387,N_38143,N_31495);
and U47388 (N_47388,N_39838,N_31615);
xnor U47389 (N_47389,N_30142,N_39928);
nand U47390 (N_47390,N_39817,N_37377);
nor U47391 (N_47391,N_32947,N_39633);
and U47392 (N_47392,N_31599,N_39570);
xnor U47393 (N_47393,N_32791,N_36719);
nand U47394 (N_47394,N_38644,N_39342);
nor U47395 (N_47395,N_31266,N_36610);
nand U47396 (N_47396,N_36020,N_37966);
nand U47397 (N_47397,N_34081,N_31701);
nand U47398 (N_47398,N_30588,N_39270);
nor U47399 (N_47399,N_32418,N_34177);
or U47400 (N_47400,N_33722,N_35790);
xor U47401 (N_47401,N_33425,N_38324);
xnor U47402 (N_47402,N_32525,N_30101);
nand U47403 (N_47403,N_36109,N_30089);
nor U47404 (N_47404,N_36752,N_30759);
and U47405 (N_47405,N_39139,N_35611);
xor U47406 (N_47406,N_34458,N_36775);
nand U47407 (N_47407,N_31410,N_30119);
xnor U47408 (N_47408,N_34187,N_39540);
xor U47409 (N_47409,N_31981,N_39064);
and U47410 (N_47410,N_30543,N_33907);
and U47411 (N_47411,N_38807,N_37913);
xor U47412 (N_47412,N_31415,N_36684);
xnor U47413 (N_47413,N_32857,N_34951);
xnor U47414 (N_47414,N_39381,N_39517);
or U47415 (N_47415,N_33316,N_37151);
and U47416 (N_47416,N_33456,N_31923);
or U47417 (N_47417,N_34638,N_37318);
and U47418 (N_47418,N_36475,N_35405);
nand U47419 (N_47419,N_31303,N_38813);
and U47420 (N_47420,N_32439,N_32941);
nand U47421 (N_47421,N_31218,N_33345);
or U47422 (N_47422,N_37827,N_34499);
and U47423 (N_47423,N_38302,N_39291);
nand U47424 (N_47424,N_36935,N_39025);
xnor U47425 (N_47425,N_39675,N_39580);
xnor U47426 (N_47426,N_37854,N_30822);
xor U47427 (N_47427,N_37789,N_36414);
xnor U47428 (N_47428,N_34011,N_32969);
and U47429 (N_47429,N_32027,N_31963);
or U47430 (N_47430,N_32366,N_37810);
nor U47431 (N_47431,N_32448,N_32220);
xor U47432 (N_47432,N_39570,N_35623);
xor U47433 (N_47433,N_32358,N_33943);
and U47434 (N_47434,N_37680,N_38715);
xnor U47435 (N_47435,N_38964,N_38717);
xnor U47436 (N_47436,N_35367,N_37346);
or U47437 (N_47437,N_31517,N_36327);
and U47438 (N_47438,N_36358,N_30811);
nor U47439 (N_47439,N_34816,N_30008);
or U47440 (N_47440,N_38022,N_32199);
xnor U47441 (N_47441,N_37429,N_33363);
or U47442 (N_47442,N_34483,N_35752);
or U47443 (N_47443,N_35753,N_37069);
and U47444 (N_47444,N_37476,N_37987);
and U47445 (N_47445,N_37191,N_39243);
nand U47446 (N_47446,N_35258,N_32602);
and U47447 (N_47447,N_32539,N_35412);
and U47448 (N_47448,N_34807,N_31079);
or U47449 (N_47449,N_36369,N_30307);
or U47450 (N_47450,N_30672,N_33459);
nor U47451 (N_47451,N_36739,N_30781);
or U47452 (N_47452,N_39307,N_38930);
or U47453 (N_47453,N_33174,N_38265);
nor U47454 (N_47454,N_38789,N_31088);
nand U47455 (N_47455,N_39064,N_35509);
nand U47456 (N_47456,N_35348,N_33806);
and U47457 (N_47457,N_38202,N_38265);
nand U47458 (N_47458,N_37031,N_34759);
nor U47459 (N_47459,N_32312,N_30611);
nor U47460 (N_47460,N_35329,N_36543);
nand U47461 (N_47461,N_37021,N_35490);
and U47462 (N_47462,N_32987,N_33347);
xor U47463 (N_47463,N_36893,N_37104);
or U47464 (N_47464,N_38378,N_33399);
or U47465 (N_47465,N_31234,N_31676);
and U47466 (N_47466,N_39583,N_39174);
xor U47467 (N_47467,N_37453,N_37452);
nand U47468 (N_47468,N_31406,N_38938);
nor U47469 (N_47469,N_33859,N_38973);
or U47470 (N_47470,N_32390,N_32336);
and U47471 (N_47471,N_36765,N_37043);
or U47472 (N_47472,N_30009,N_38669);
nor U47473 (N_47473,N_30629,N_35469);
xor U47474 (N_47474,N_35668,N_39674);
nand U47475 (N_47475,N_33478,N_39908);
nor U47476 (N_47476,N_36172,N_34070);
xnor U47477 (N_47477,N_33438,N_38215);
and U47478 (N_47478,N_36727,N_34656);
nand U47479 (N_47479,N_35144,N_30812);
and U47480 (N_47480,N_31662,N_31339);
xnor U47481 (N_47481,N_39234,N_39809);
xnor U47482 (N_47482,N_39065,N_37111);
nor U47483 (N_47483,N_31692,N_32702);
nand U47484 (N_47484,N_38740,N_35194);
and U47485 (N_47485,N_36550,N_34590);
nor U47486 (N_47486,N_32271,N_37157);
nor U47487 (N_47487,N_32487,N_36821);
or U47488 (N_47488,N_35581,N_30400);
or U47489 (N_47489,N_34433,N_30293);
nor U47490 (N_47490,N_33794,N_35588);
or U47491 (N_47491,N_37455,N_30889);
and U47492 (N_47492,N_31861,N_38074);
nand U47493 (N_47493,N_36982,N_36143);
nand U47494 (N_47494,N_33943,N_30386);
and U47495 (N_47495,N_30008,N_38848);
xor U47496 (N_47496,N_32872,N_39065);
xor U47497 (N_47497,N_36260,N_37860);
and U47498 (N_47498,N_35762,N_36932);
and U47499 (N_47499,N_34440,N_37822);
or U47500 (N_47500,N_35758,N_36037);
xnor U47501 (N_47501,N_39292,N_30324);
nor U47502 (N_47502,N_32111,N_35998);
and U47503 (N_47503,N_32785,N_37872);
nand U47504 (N_47504,N_35294,N_30636);
and U47505 (N_47505,N_32921,N_35321);
and U47506 (N_47506,N_39163,N_36384);
nand U47507 (N_47507,N_38279,N_38954);
xnor U47508 (N_47508,N_30581,N_33459);
or U47509 (N_47509,N_31345,N_32971);
nand U47510 (N_47510,N_32863,N_33959);
xnor U47511 (N_47511,N_35693,N_36160);
xnor U47512 (N_47512,N_30043,N_39539);
nor U47513 (N_47513,N_37215,N_37944);
and U47514 (N_47514,N_34098,N_32816);
or U47515 (N_47515,N_37161,N_37897);
nand U47516 (N_47516,N_39008,N_32557);
or U47517 (N_47517,N_36206,N_36948);
nand U47518 (N_47518,N_31754,N_39961);
and U47519 (N_47519,N_38985,N_34167);
and U47520 (N_47520,N_30818,N_31733);
xnor U47521 (N_47521,N_30802,N_37327);
nor U47522 (N_47522,N_35031,N_30992);
nand U47523 (N_47523,N_30740,N_34106);
and U47524 (N_47524,N_39122,N_37113);
nor U47525 (N_47525,N_39562,N_30558);
and U47526 (N_47526,N_36067,N_30093);
xor U47527 (N_47527,N_34239,N_37965);
nand U47528 (N_47528,N_32593,N_36421);
and U47529 (N_47529,N_35157,N_32391);
nand U47530 (N_47530,N_35372,N_38320);
nand U47531 (N_47531,N_39586,N_31389);
nand U47532 (N_47532,N_32688,N_38631);
xor U47533 (N_47533,N_35690,N_35471);
and U47534 (N_47534,N_35123,N_31105);
and U47535 (N_47535,N_38750,N_39920);
xnor U47536 (N_47536,N_33898,N_34762);
nor U47537 (N_47537,N_34785,N_37783);
or U47538 (N_47538,N_39555,N_33092);
xor U47539 (N_47539,N_31043,N_34976);
nor U47540 (N_47540,N_35937,N_35960);
and U47541 (N_47541,N_35361,N_33735);
nor U47542 (N_47542,N_36999,N_34658);
xor U47543 (N_47543,N_32578,N_32718);
nor U47544 (N_47544,N_35199,N_39338);
or U47545 (N_47545,N_35745,N_35648);
nand U47546 (N_47546,N_32438,N_34959);
xor U47547 (N_47547,N_39535,N_35328);
and U47548 (N_47548,N_33681,N_30045);
nor U47549 (N_47549,N_30024,N_38293);
or U47550 (N_47550,N_33393,N_39120);
xor U47551 (N_47551,N_38023,N_34675);
xor U47552 (N_47552,N_36578,N_39520);
or U47553 (N_47553,N_38212,N_30657);
xor U47554 (N_47554,N_35443,N_37135);
and U47555 (N_47555,N_35445,N_38827);
and U47556 (N_47556,N_34663,N_39020);
and U47557 (N_47557,N_39324,N_36257);
and U47558 (N_47558,N_30362,N_31624);
xnor U47559 (N_47559,N_35951,N_32723);
xor U47560 (N_47560,N_34189,N_38950);
nand U47561 (N_47561,N_30198,N_35693);
and U47562 (N_47562,N_36840,N_36428);
and U47563 (N_47563,N_30889,N_37977);
xnor U47564 (N_47564,N_31795,N_39852);
nor U47565 (N_47565,N_34054,N_37995);
or U47566 (N_47566,N_39164,N_31795);
nor U47567 (N_47567,N_38383,N_31445);
xnor U47568 (N_47568,N_33051,N_36944);
xnor U47569 (N_47569,N_32356,N_34371);
nand U47570 (N_47570,N_30464,N_32921);
and U47571 (N_47571,N_34585,N_34346);
or U47572 (N_47572,N_33228,N_31122);
nor U47573 (N_47573,N_36794,N_38974);
nor U47574 (N_47574,N_37152,N_36323);
and U47575 (N_47575,N_36431,N_33843);
nand U47576 (N_47576,N_36152,N_36467);
and U47577 (N_47577,N_33092,N_30117);
or U47578 (N_47578,N_36241,N_32635);
or U47579 (N_47579,N_38688,N_32917);
and U47580 (N_47580,N_37139,N_35185);
nand U47581 (N_47581,N_30746,N_39087);
nand U47582 (N_47582,N_39996,N_31091);
and U47583 (N_47583,N_35826,N_37269);
and U47584 (N_47584,N_32606,N_34529);
and U47585 (N_47585,N_37275,N_39364);
nand U47586 (N_47586,N_38161,N_37766);
or U47587 (N_47587,N_39223,N_31341);
nor U47588 (N_47588,N_36609,N_36014);
or U47589 (N_47589,N_33637,N_37909);
or U47590 (N_47590,N_34478,N_37166);
xnor U47591 (N_47591,N_36003,N_38124);
nor U47592 (N_47592,N_39396,N_39301);
nand U47593 (N_47593,N_35866,N_32221);
and U47594 (N_47594,N_33433,N_32492);
nand U47595 (N_47595,N_34171,N_35176);
nor U47596 (N_47596,N_38988,N_38899);
xnor U47597 (N_47597,N_33149,N_35423);
nor U47598 (N_47598,N_31458,N_32367);
and U47599 (N_47599,N_37101,N_32105);
nand U47600 (N_47600,N_34903,N_35867);
nand U47601 (N_47601,N_36428,N_32954);
xor U47602 (N_47602,N_39111,N_30550);
nor U47603 (N_47603,N_31741,N_36716);
nor U47604 (N_47604,N_35268,N_30228);
xnor U47605 (N_47605,N_31885,N_37392);
and U47606 (N_47606,N_38784,N_32038);
and U47607 (N_47607,N_30749,N_35852);
nand U47608 (N_47608,N_36456,N_36581);
nor U47609 (N_47609,N_37344,N_38600);
nor U47610 (N_47610,N_37606,N_35633);
and U47611 (N_47611,N_33568,N_37679);
xnor U47612 (N_47612,N_38058,N_36268);
and U47613 (N_47613,N_30561,N_34871);
nand U47614 (N_47614,N_34905,N_35196);
and U47615 (N_47615,N_35906,N_33187);
and U47616 (N_47616,N_30558,N_31022);
nand U47617 (N_47617,N_36021,N_31618);
nand U47618 (N_47618,N_32535,N_37321);
or U47619 (N_47619,N_32460,N_39644);
and U47620 (N_47620,N_36205,N_37842);
xor U47621 (N_47621,N_39938,N_37685);
and U47622 (N_47622,N_33234,N_35413);
nor U47623 (N_47623,N_39557,N_38132);
nand U47624 (N_47624,N_38693,N_33074);
nand U47625 (N_47625,N_31164,N_39685);
nor U47626 (N_47626,N_39293,N_34364);
nor U47627 (N_47627,N_32983,N_38572);
xor U47628 (N_47628,N_36289,N_32597);
xnor U47629 (N_47629,N_36513,N_38162);
and U47630 (N_47630,N_38978,N_37197);
and U47631 (N_47631,N_36034,N_34810);
or U47632 (N_47632,N_33873,N_30170);
or U47633 (N_47633,N_32880,N_30011);
and U47634 (N_47634,N_31279,N_33612);
nor U47635 (N_47635,N_35277,N_37362);
or U47636 (N_47636,N_37413,N_34086);
nor U47637 (N_47637,N_37792,N_36680);
or U47638 (N_47638,N_37331,N_32281);
and U47639 (N_47639,N_39717,N_36496);
xor U47640 (N_47640,N_30983,N_33020);
xor U47641 (N_47641,N_30975,N_31860);
nor U47642 (N_47642,N_34541,N_35692);
or U47643 (N_47643,N_39308,N_31509);
xor U47644 (N_47644,N_30756,N_39727);
nand U47645 (N_47645,N_32034,N_38949);
and U47646 (N_47646,N_31720,N_31424);
or U47647 (N_47647,N_37602,N_32657);
and U47648 (N_47648,N_33563,N_39301);
and U47649 (N_47649,N_37729,N_33308);
and U47650 (N_47650,N_38581,N_32118);
xnor U47651 (N_47651,N_31491,N_31695);
or U47652 (N_47652,N_38515,N_34280);
nand U47653 (N_47653,N_32516,N_37104);
or U47654 (N_47654,N_30778,N_31055);
nand U47655 (N_47655,N_34577,N_38969);
or U47656 (N_47656,N_34224,N_35091);
or U47657 (N_47657,N_36244,N_30987);
nand U47658 (N_47658,N_39307,N_30854);
xnor U47659 (N_47659,N_30884,N_32100);
or U47660 (N_47660,N_39087,N_39741);
nor U47661 (N_47661,N_30767,N_38021);
nand U47662 (N_47662,N_34117,N_39383);
nand U47663 (N_47663,N_30868,N_34142);
nor U47664 (N_47664,N_31396,N_34758);
nor U47665 (N_47665,N_35385,N_32545);
nand U47666 (N_47666,N_34385,N_36555);
nor U47667 (N_47667,N_35175,N_35635);
xnor U47668 (N_47668,N_37236,N_35313);
xnor U47669 (N_47669,N_38021,N_31269);
nor U47670 (N_47670,N_35928,N_35603);
nor U47671 (N_47671,N_38861,N_33396);
nor U47672 (N_47672,N_30515,N_38685);
nor U47673 (N_47673,N_31011,N_37916);
nor U47674 (N_47674,N_33207,N_33296);
nor U47675 (N_47675,N_32566,N_36824);
nand U47676 (N_47676,N_32582,N_30710);
xor U47677 (N_47677,N_39907,N_38337);
or U47678 (N_47678,N_32881,N_32849);
nand U47679 (N_47679,N_33131,N_30064);
nor U47680 (N_47680,N_32496,N_34057);
nor U47681 (N_47681,N_32740,N_35929);
nor U47682 (N_47682,N_36277,N_38254);
or U47683 (N_47683,N_35487,N_32400);
and U47684 (N_47684,N_30248,N_36825);
xnor U47685 (N_47685,N_33477,N_38715);
and U47686 (N_47686,N_34742,N_37014);
xnor U47687 (N_47687,N_31707,N_39834);
nor U47688 (N_47688,N_34841,N_32176);
or U47689 (N_47689,N_39140,N_37684);
xor U47690 (N_47690,N_36231,N_30837);
nand U47691 (N_47691,N_37216,N_39567);
nor U47692 (N_47692,N_36145,N_36459);
or U47693 (N_47693,N_31621,N_36194);
nor U47694 (N_47694,N_34605,N_32517);
nor U47695 (N_47695,N_38386,N_34496);
nor U47696 (N_47696,N_31223,N_33139);
nor U47697 (N_47697,N_33901,N_37187);
nor U47698 (N_47698,N_32805,N_31174);
or U47699 (N_47699,N_30339,N_36749);
nand U47700 (N_47700,N_35156,N_39307);
or U47701 (N_47701,N_39907,N_35622);
nor U47702 (N_47702,N_36138,N_34785);
and U47703 (N_47703,N_38725,N_33526);
xor U47704 (N_47704,N_39526,N_34518);
nor U47705 (N_47705,N_32557,N_30551);
nor U47706 (N_47706,N_39244,N_38368);
nand U47707 (N_47707,N_38157,N_35317);
or U47708 (N_47708,N_36030,N_33785);
xnor U47709 (N_47709,N_33003,N_36051);
nor U47710 (N_47710,N_38705,N_39341);
nor U47711 (N_47711,N_33721,N_39603);
and U47712 (N_47712,N_32780,N_36993);
xnor U47713 (N_47713,N_37225,N_36574);
nor U47714 (N_47714,N_32010,N_35539);
and U47715 (N_47715,N_32476,N_32614);
and U47716 (N_47716,N_39000,N_37926);
or U47717 (N_47717,N_39636,N_31474);
xnor U47718 (N_47718,N_39129,N_37349);
xnor U47719 (N_47719,N_38796,N_38225);
xor U47720 (N_47720,N_34825,N_31390);
nor U47721 (N_47721,N_34570,N_36034);
xor U47722 (N_47722,N_35556,N_38084);
nor U47723 (N_47723,N_35943,N_39502);
or U47724 (N_47724,N_32135,N_39664);
or U47725 (N_47725,N_32592,N_30171);
nor U47726 (N_47726,N_38131,N_33069);
or U47727 (N_47727,N_33501,N_30689);
and U47728 (N_47728,N_38235,N_37520);
nand U47729 (N_47729,N_31863,N_37382);
and U47730 (N_47730,N_35285,N_30679);
nor U47731 (N_47731,N_31813,N_38188);
nand U47732 (N_47732,N_30518,N_32927);
xnor U47733 (N_47733,N_31915,N_39610);
and U47734 (N_47734,N_34944,N_31981);
nor U47735 (N_47735,N_30742,N_33952);
nor U47736 (N_47736,N_37734,N_38876);
nor U47737 (N_47737,N_37909,N_38294);
and U47738 (N_47738,N_35640,N_38798);
nand U47739 (N_47739,N_31924,N_33719);
or U47740 (N_47740,N_30889,N_36294);
or U47741 (N_47741,N_34854,N_32571);
and U47742 (N_47742,N_30804,N_33262);
nor U47743 (N_47743,N_35288,N_35315);
and U47744 (N_47744,N_34794,N_37040);
and U47745 (N_47745,N_30399,N_32204);
or U47746 (N_47746,N_31907,N_36972);
nor U47747 (N_47747,N_32972,N_39827);
or U47748 (N_47748,N_37477,N_32860);
nor U47749 (N_47749,N_30013,N_38898);
nand U47750 (N_47750,N_35984,N_38398);
nor U47751 (N_47751,N_37757,N_37696);
and U47752 (N_47752,N_36939,N_32558);
and U47753 (N_47753,N_34236,N_31500);
xnor U47754 (N_47754,N_38591,N_30414);
nand U47755 (N_47755,N_36826,N_39613);
or U47756 (N_47756,N_39996,N_36849);
xor U47757 (N_47757,N_36366,N_33175);
or U47758 (N_47758,N_30090,N_35242);
nor U47759 (N_47759,N_34883,N_35754);
nand U47760 (N_47760,N_32456,N_37859);
nand U47761 (N_47761,N_34935,N_39257);
or U47762 (N_47762,N_33912,N_32830);
nand U47763 (N_47763,N_33959,N_36585);
xnor U47764 (N_47764,N_36535,N_37387);
xnor U47765 (N_47765,N_31240,N_32356);
or U47766 (N_47766,N_36184,N_39003);
and U47767 (N_47767,N_33133,N_32460);
or U47768 (N_47768,N_31949,N_38075);
xnor U47769 (N_47769,N_34862,N_32440);
nand U47770 (N_47770,N_34271,N_38197);
xnor U47771 (N_47771,N_37645,N_36347);
and U47772 (N_47772,N_33922,N_39387);
xnor U47773 (N_47773,N_35492,N_37581);
nand U47774 (N_47774,N_31085,N_31241);
and U47775 (N_47775,N_38637,N_39099);
and U47776 (N_47776,N_30744,N_39923);
xor U47777 (N_47777,N_32435,N_33829);
nor U47778 (N_47778,N_31068,N_35596);
nor U47779 (N_47779,N_39545,N_37752);
and U47780 (N_47780,N_31077,N_32814);
nand U47781 (N_47781,N_33861,N_36496);
xor U47782 (N_47782,N_38371,N_31851);
nand U47783 (N_47783,N_31755,N_31780);
and U47784 (N_47784,N_30307,N_35402);
nor U47785 (N_47785,N_37463,N_33253);
or U47786 (N_47786,N_34996,N_37252);
nand U47787 (N_47787,N_34552,N_30935);
or U47788 (N_47788,N_34887,N_39438);
nand U47789 (N_47789,N_30946,N_38480);
nor U47790 (N_47790,N_31696,N_30247);
nand U47791 (N_47791,N_38942,N_32914);
nor U47792 (N_47792,N_35524,N_35209);
xnor U47793 (N_47793,N_36198,N_31736);
or U47794 (N_47794,N_35659,N_33677);
nand U47795 (N_47795,N_35168,N_33570);
nor U47796 (N_47796,N_37031,N_39660);
and U47797 (N_47797,N_38133,N_33115);
xor U47798 (N_47798,N_32156,N_35724);
or U47799 (N_47799,N_31262,N_33928);
nand U47800 (N_47800,N_30305,N_39108);
nor U47801 (N_47801,N_37448,N_32054);
nand U47802 (N_47802,N_36303,N_36570);
nor U47803 (N_47803,N_33111,N_35487);
xor U47804 (N_47804,N_35666,N_35276);
and U47805 (N_47805,N_37032,N_33319);
or U47806 (N_47806,N_36123,N_33762);
and U47807 (N_47807,N_37901,N_39338);
xnor U47808 (N_47808,N_37682,N_33792);
nor U47809 (N_47809,N_38648,N_37153);
or U47810 (N_47810,N_35687,N_31845);
nand U47811 (N_47811,N_34383,N_32993);
nand U47812 (N_47812,N_36695,N_34469);
nand U47813 (N_47813,N_39091,N_37103);
nor U47814 (N_47814,N_33603,N_33728);
nand U47815 (N_47815,N_37048,N_37852);
and U47816 (N_47816,N_30850,N_36917);
nand U47817 (N_47817,N_37442,N_39795);
xnor U47818 (N_47818,N_37924,N_30891);
and U47819 (N_47819,N_39377,N_39922);
nand U47820 (N_47820,N_35642,N_30656);
or U47821 (N_47821,N_30142,N_36245);
and U47822 (N_47822,N_36740,N_31154);
xnor U47823 (N_47823,N_33919,N_30303);
nand U47824 (N_47824,N_34344,N_39818);
xor U47825 (N_47825,N_35277,N_30273);
xor U47826 (N_47826,N_35619,N_36287);
and U47827 (N_47827,N_35101,N_36165);
nand U47828 (N_47828,N_38185,N_39953);
and U47829 (N_47829,N_37655,N_30469);
or U47830 (N_47830,N_39755,N_39955);
and U47831 (N_47831,N_32870,N_32899);
or U47832 (N_47832,N_36470,N_35076);
nor U47833 (N_47833,N_31333,N_31797);
and U47834 (N_47834,N_35160,N_33306);
and U47835 (N_47835,N_35863,N_34428);
nand U47836 (N_47836,N_30195,N_36930);
or U47837 (N_47837,N_31358,N_36702);
nor U47838 (N_47838,N_38242,N_38565);
nor U47839 (N_47839,N_38630,N_31605);
or U47840 (N_47840,N_33777,N_38186);
nor U47841 (N_47841,N_35532,N_31090);
and U47842 (N_47842,N_39744,N_32151);
xor U47843 (N_47843,N_39402,N_31216);
nor U47844 (N_47844,N_32521,N_30028);
xor U47845 (N_47845,N_34909,N_37837);
and U47846 (N_47846,N_31116,N_34738);
nor U47847 (N_47847,N_38167,N_36537);
or U47848 (N_47848,N_32204,N_35021);
or U47849 (N_47849,N_30774,N_30565);
or U47850 (N_47850,N_37773,N_37779);
nand U47851 (N_47851,N_35148,N_33543);
xor U47852 (N_47852,N_33082,N_36997);
xor U47853 (N_47853,N_32686,N_35489);
or U47854 (N_47854,N_33668,N_38453);
nand U47855 (N_47855,N_38148,N_39762);
nor U47856 (N_47856,N_31943,N_35928);
or U47857 (N_47857,N_39395,N_36449);
or U47858 (N_47858,N_35732,N_33354);
nand U47859 (N_47859,N_30561,N_39287);
nor U47860 (N_47860,N_31608,N_39720);
xnor U47861 (N_47861,N_30285,N_34371);
and U47862 (N_47862,N_31007,N_31578);
and U47863 (N_47863,N_32472,N_33299);
or U47864 (N_47864,N_34954,N_39603);
nor U47865 (N_47865,N_34778,N_36456);
xnor U47866 (N_47866,N_30033,N_39029);
nor U47867 (N_47867,N_38244,N_33890);
or U47868 (N_47868,N_32286,N_35703);
or U47869 (N_47869,N_32987,N_36902);
xnor U47870 (N_47870,N_39298,N_33206);
and U47871 (N_47871,N_36426,N_32845);
nand U47872 (N_47872,N_34650,N_34661);
nor U47873 (N_47873,N_33223,N_39562);
nand U47874 (N_47874,N_31453,N_36825);
and U47875 (N_47875,N_37336,N_30922);
nand U47876 (N_47876,N_37094,N_31604);
xnor U47877 (N_47877,N_32331,N_39036);
nor U47878 (N_47878,N_38323,N_35017);
xor U47879 (N_47879,N_37058,N_30093);
nand U47880 (N_47880,N_32618,N_38124);
and U47881 (N_47881,N_35047,N_37826);
nand U47882 (N_47882,N_34059,N_36627);
and U47883 (N_47883,N_37203,N_33084);
nand U47884 (N_47884,N_34427,N_30793);
nor U47885 (N_47885,N_35786,N_38737);
or U47886 (N_47886,N_37690,N_36977);
nand U47887 (N_47887,N_31048,N_33846);
nor U47888 (N_47888,N_33465,N_34026);
nor U47889 (N_47889,N_38614,N_32324);
nor U47890 (N_47890,N_30363,N_33224);
nor U47891 (N_47891,N_38499,N_38231);
nor U47892 (N_47892,N_30218,N_32345);
xnor U47893 (N_47893,N_37110,N_37114);
xnor U47894 (N_47894,N_39977,N_34563);
xor U47895 (N_47895,N_32186,N_36683);
and U47896 (N_47896,N_32263,N_32624);
or U47897 (N_47897,N_38555,N_36750);
nor U47898 (N_47898,N_35266,N_35447);
or U47899 (N_47899,N_38664,N_37095);
or U47900 (N_47900,N_37629,N_39237);
nor U47901 (N_47901,N_39860,N_34182);
xor U47902 (N_47902,N_35626,N_37859);
and U47903 (N_47903,N_36363,N_31420);
nand U47904 (N_47904,N_39159,N_31014);
or U47905 (N_47905,N_31672,N_37246);
nand U47906 (N_47906,N_36814,N_34714);
nand U47907 (N_47907,N_39984,N_33728);
nand U47908 (N_47908,N_37269,N_31447);
and U47909 (N_47909,N_35838,N_30759);
nor U47910 (N_47910,N_35690,N_34721);
nor U47911 (N_47911,N_39223,N_39536);
xor U47912 (N_47912,N_36765,N_33954);
xor U47913 (N_47913,N_33623,N_30491);
nand U47914 (N_47914,N_33963,N_36445);
and U47915 (N_47915,N_30885,N_30736);
or U47916 (N_47916,N_31456,N_34881);
nand U47917 (N_47917,N_38759,N_34885);
or U47918 (N_47918,N_32809,N_37559);
or U47919 (N_47919,N_36564,N_30844);
and U47920 (N_47920,N_34444,N_37992);
and U47921 (N_47921,N_32036,N_30050);
xnor U47922 (N_47922,N_31748,N_39698);
nand U47923 (N_47923,N_36258,N_36110);
nand U47924 (N_47924,N_33759,N_39073);
and U47925 (N_47925,N_36270,N_32474);
xor U47926 (N_47926,N_38356,N_36561);
or U47927 (N_47927,N_34722,N_38541);
xor U47928 (N_47928,N_32870,N_31569);
nor U47929 (N_47929,N_31106,N_37192);
nand U47930 (N_47930,N_34153,N_36378);
or U47931 (N_47931,N_31120,N_33164);
or U47932 (N_47932,N_39814,N_37673);
nand U47933 (N_47933,N_30859,N_30862);
or U47934 (N_47934,N_39029,N_36706);
nor U47935 (N_47935,N_30732,N_36278);
nand U47936 (N_47936,N_37059,N_39671);
and U47937 (N_47937,N_35673,N_37945);
nand U47938 (N_47938,N_32834,N_39407);
or U47939 (N_47939,N_39433,N_32605);
nor U47940 (N_47940,N_37980,N_35168);
nand U47941 (N_47941,N_33868,N_39072);
xnor U47942 (N_47942,N_32023,N_36627);
xnor U47943 (N_47943,N_31805,N_38801);
or U47944 (N_47944,N_39562,N_39386);
or U47945 (N_47945,N_39376,N_33615);
and U47946 (N_47946,N_34632,N_33734);
nor U47947 (N_47947,N_30012,N_32947);
and U47948 (N_47948,N_33845,N_36729);
nor U47949 (N_47949,N_30834,N_33581);
nand U47950 (N_47950,N_32286,N_39239);
xnor U47951 (N_47951,N_32171,N_35565);
nand U47952 (N_47952,N_33517,N_30133);
nor U47953 (N_47953,N_31365,N_34380);
nor U47954 (N_47954,N_34427,N_34978);
xor U47955 (N_47955,N_35339,N_35924);
nand U47956 (N_47956,N_31145,N_39448);
or U47957 (N_47957,N_37134,N_31375);
nor U47958 (N_47958,N_38524,N_35489);
or U47959 (N_47959,N_36753,N_36771);
nor U47960 (N_47960,N_36161,N_32472);
xnor U47961 (N_47961,N_34113,N_31027);
and U47962 (N_47962,N_31132,N_38161);
xnor U47963 (N_47963,N_31454,N_34608);
or U47964 (N_47964,N_35107,N_37101);
nor U47965 (N_47965,N_32853,N_37428);
and U47966 (N_47966,N_36638,N_33633);
xnor U47967 (N_47967,N_31880,N_32284);
xor U47968 (N_47968,N_33467,N_37738);
or U47969 (N_47969,N_39588,N_33375);
and U47970 (N_47970,N_38084,N_33272);
nor U47971 (N_47971,N_34256,N_31990);
nand U47972 (N_47972,N_38771,N_36953);
or U47973 (N_47973,N_33599,N_35466);
or U47974 (N_47974,N_36758,N_36244);
nand U47975 (N_47975,N_33723,N_36596);
or U47976 (N_47976,N_37445,N_31089);
xor U47977 (N_47977,N_36646,N_38246);
xnor U47978 (N_47978,N_33552,N_36953);
nor U47979 (N_47979,N_35941,N_36067);
nor U47980 (N_47980,N_36584,N_33783);
nand U47981 (N_47981,N_39851,N_37038);
nor U47982 (N_47982,N_31348,N_31694);
xnor U47983 (N_47983,N_37146,N_39413);
nand U47984 (N_47984,N_37896,N_32091);
and U47985 (N_47985,N_39861,N_38868);
xnor U47986 (N_47986,N_33987,N_34034);
or U47987 (N_47987,N_31965,N_39672);
and U47988 (N_47988,N_34470,N_33442);
and U47989 (N_47989,N_39632,N_37365);
xnor U47990 (N_47990,N_35010,N_32568);
nor U47991 (N_47991,N_35887,N_33127);
nor U47992 (N_47992,N_39595,N_31759);
nand U47993 (N_47993,N_34531,N_30823);
nor U47994 (N_47994,N_33980,N_36641);
nand U47995 (N_47995,N_31783,N_39391);
or U47996 (N_47996,N_37259,N_32282);
or U47997 (N_47997,N_32493,N_32326);
and U47998 (N_47998,N_35411,N_30532);
or U47999 (N_47999,N_36420,N_37998);
nand U48000 (N_48000,N_31884,N_37772);
nand U48001 (N_48001,N_33526,N_33393);
xnor U48002 (N_48002,N_36430,N_36018);
or U48003 (N_48003,N_37589,N_32329);
and U48004 (N_48004,N_32882,N_32659);
and U48005 (N_48005,N_37461,N_30914);
xor U48006 (N_48006,N_38531,N_35905);
or U48007 (N_48007,N_30427,N_30766);
nand U48008 (N_48008,N_31987,N_38141);
and U48009 (N_48009,N_31096,N_33419);
nor U48010 (N_48010,N_36891,N_35512);
nand U48011 (N_48011,N_39865,N_32509);
xor U48012 (N_48012,N_39995,N_38971);
xor U48013 (N_48013,N_39970,N_39752);
and U48014 (N_48014,N_31157,N_35468);
nand U48015 (N_48015,N_39340,N_31557);
nor U48016 (N_48016,N_34864,N_38262);
or U48017 (N_48017,N_33938,N_30581);
xor U48018 (N_48018,N_37952,N_34177);
or U48019 (N_48019,N_32339,N_36745);
and U48020 (N_48020,N_33842,N_37134);
xnor U48021 (N_48021,N_38587,N_33562);
and U48022 (N_48022,N_31084,N_36217);
xor U48023 (N_48023,N_32714,N_31466);
nor U48024 (N_48024,N_35396,N_33752);
nor U48025 (N_48025,N_30469,N_35897);
nor U48026 (N_48026,N_32187,N_30540);
nand U48027 (N_48027,N_33520,N_30871);
nand U48028 (N_48028,N_39552,N_37491);
xnor U48029 (N_48029,N_39478,N_30175);
or U48030 (N_48030,N_32547,N_30108);
or U48031 (N_48031,N_38470,N_38919);
xnor U48032 (N_48032,N_35455,N_39793);
xnor U48033 (N_48033,N_33276,N_34159);
nand U48034 (N_48034,N_38809,N_35275);
xnor U48035 (N_48035,N_33865,N_36876);
and U48036 (N_48036,N_38073,N_30968);
xor U48037 (N_48037,N_36361,N_39584);
nand U48038 (N_48038,N_39722,N_31013);
xor U48039 (N_48039,N_38769,N_38917);
xnor U48040 (N_48040,N_35204,N_32202);
xor U48041 (N_48041,N_36107,N_39365);
nand U48042 (N_48042,N_37924,N_31222);
xnor U48043 (N_48043,N_39624,N_38326);
and U48044 (N_48044,N_31924,N_30071);
or U48045 (N_48045,N_32661,N_30714);
xor U48046 (N_48046,N_32641,N_36685);
nor U48047 (N_48047,N_32328,N_39226);
nor U48048 (N_48048,N_34038,N_33231);
or U48049 (N_48049,N_37738,N_33594);
and U48050 (N_48050,N_32007,N_33079);
or U48051 (N_48051,N_34342,N_39248);
nor U48052 (N_48052,N_31184,N_31649);
nand U48053 (N_48053,N_38787,N_38038);
or U48054 (N_48054,N_32835,N_34964);
nor U48055 (N_48055,N_33438,N_39264);
xnor U48056 (N_48056,N_32191,N_30244);
xor U48057 (N_48057,N_33223,N_30401);
nand U48058 (N_48058,N_39831,N_37783);
nand U48059 (N_48059,N_31191,N_31213);
and U48060 (N_48060,N_39192,N_34029);
or U48061 (N_48061,N_32098,N_34743);
nand U48062 (N_48062,N_39356,N_35705);
or U48063 (N_48063,N_37783,N_39649);
and U48064 (N_48064,N_33647,N_38933);
nand U48065 (N_48065,N_36352,N_38517);
or U48066 (N_48066,N_34958,N_35941);
and U48067 (N_48067,N_30406,N_38936);
and U48068 (N_48068,N_33885,N_31842);
or U48069 (N_48069,N_36746,N_32574);
xor U48070 (N_48070,N_32458,N_35637);
nand U48071 (N_48071,N_30727,N_30829);
or U48072 (N_48072,N_36779,N_33632);
nor U48073 (N_48073,N_32796,N_34297);
nand U48074 (N_48074,N_37188,N_39197);
nand U48075 (N_48075,N_37000,N_35144);
xnor U48076 (N_48076,N_38472,N_38167);
or U48077 (N_48077,N_31787,N_34981);
nor U48078 (N_48078,N_33269,N_35302);
nand U48079 (N_48079,N_32279,N_39370);
or U48080 (N_48080,N_31517,N_32533);
nand U48081 (N_48081,N_33798,N_39619);
xnor U48082 (N_48082,N_34332,N_34617);
xnor U48083 (N_48083,N_36041,N_33482);
nand U48084 (N_48084,N_33197,N_32957);
nand U48085 (N_48085,N_36434,N_30268);
xnor U48086 (N_48086,N_35565,N_39514);
xor U48087 (N_48087,N_35638,N_32344);
xor U48088 (N_48088,N_37089,N_37698);
xnor U48089 (N_48089,N_33037,N_31022);
xnor U48090 (N_48090,N_37432,N_36524);
or U48091 (N_48091,N_36856,N_34286);
xor U48092 (N_48092,N_36999,N_37673);
and U48093 (N_48093,N_38034,N_30422);
nor U48094 (N_48094,N_36905,N_35673);
xnor U48095 (N_48095,N_36199,N_35210);
and U48096 (N_48096,N_32689,N_37357);
or U48097 (N_48097,N_30524,N_37565);
nor U48098 (N_48098,N_38691,N_31555);
xnor U48099 (N_48099,N_31062,N_35040);
nand U48100 (N_48100,N_36215,N_33407);
nor U48101 (N_48101,N_35149,N_34177);
and U48102 (N_48102,N_33866,N_34240);
and U48103 (N_48103,N_33087,N_38253);
nor U48104 (N_48104,N_31875,N_33457);
nand U48105 (N_48105,N_32523,N_31875);
xor U48106 (N_48106,N_32233,N_38685);
or U48107 (N_48107,N_33797,N_36318);
and U48108 (N_48108,N_32308,N_32216);
and U48109 (N_48109,N_39237,N_36801);
or U48110 (N_48110,N_33284,N_32605);
and U48111 (N_48111,N_35539,N_36532);
nor U48112 (N_48112,N_30966,N_38158);
and U48113 (N_48113,N_30670,N_37310);
nor U48114 (N_48114,N_33659,N_30612);
xnor U48115 (N_48115,N_30984,N_33929);
and U48116 (N_48116,N_36157,N_37975);
nor U48117 (N_48117,N_31563,N_38244);
and U48118 (N_48118,N_38839,N_35553);
xor U48119 (N_48119,N_38589,N_31560);
and U48120 (N_48120,N_31818,N_33440);
xnor U48121 (N_48121,N_33184,N_31196);
and U48122 (N_48122,N_38294,N_34266);
nor U48123 (N_48123,N_37460,N_39482);
nor U48124 (N_48124,N_36285,N_39081);
nor U48125 (N_48125,N_38219,N_37895);
nand U48126 (N_48126,N_34168,N_36259);
nor U48127 (N_48127,N_38639,N_33944);
xnor U48128 (N_48128,N_33710,N_35759);
nand U48129 (N_48129,N_38529,N_31385);
and U48130 (N_48130,N_31950,N_31595);
nand U48131 (N_48131,N_38425,N_31422);
or U48132 (N_48132,N_31850,N_39992);
nand U48133 (N_48133,N_35835,N_33781);
or U48134 (N_48134,N_32145,N_38846);
xor U48135 (N_48135,N_39576,N_37416);
nor U48136 (N_48136,N_32424,N_35853);
and U48137 (N_48137,N_31625,N_32931);
and U48138 (N_48138,N_34442,N_37497);
xor U48139 (N_48139,N_31399,N_37374);
or U48140 (N_48140,N_39403,N_31915);
nor U48141 (N_48141,N_38017,N_31778);
xnor U48142 (N_48142,N_32579,N_36529);
and U48143 (N_48143,N_39811,N_38460);
nand U48144 (N_48144,N_35515,N_33033);
nor U48145 (N_48145,N_39345,N_37796);
nor U48146 (N_48146,N_36594,N_36481);
nor U48147 (N_48147,N_32600,N_38843);
nor U48148 (N_48148,N_30337,N_31298);
and U48149 (N_48149,N_35232,N_30330);
xor U48150 (N_48150,N_33128,N_38122);
or U48151 (N_48151,N_39784,N_39453);
nor U48152 (N_48152,N_36296,N_35240);
nor U48153 (N_48153,N_35871,N_38519);
or U48154 (N_48154,N_31041,N_38417);
xor U48155 (N_48155,N_37048,N_34107);
xnor U48156 (N_48156,N_34156,N_37394);
nand U48157 (N_48157,N_37057,N_38991);
nor U48158 (N_48158,N_33055,N_33888);
and U48159 (N_48159,N_36167,N_30578);
xnor U48160 (N_48160,N_31908,N_31821);
xor U48161 (N_48161,N_39009,N_36605);
nor U48162 (N_48162,N_39524,N_30464);
nor U48163 (N_48163,N_33691,N_35001);
nor U48164 (N_48164,N_37571,N_34383);
nand U48165 (N_48165,N_36258,N_39034);
or U48166 (N_48166,N_30005,N_34923);
nand U48167 (N_48167,N_34359,N_39367);
nand U48168 (N_48168,N_37506,N_38355);
nor U48169 (N_48169,N_38955,N_33405);
nand U48170 (N_48170,N_34944,N_39729);
or U48171 (N_48171,N_30737,N_37648);
and U48172 (N_48172,N_39927,N_34114);
nor U48173 (N_48173,N_36947,N_33897);
nor U48174 (N_48174,N_38584,N_32793);
and U48175 (N_48175,N_39046,N_34184);
and U48176 (N_48176,N_39474,N_34274);
or U48177 (N_48177,N_34461,N_39874);
nand U48178 (N_48178,N_32413,N_30822);
or U48179 (N_48179,N_38244,N_34210);
and U48180 (N_48180,N_35190,N_33782);
nand U48181 (N_48181,N_30212,N_34507);
and U48182 (N_48182,N_30319,N_34127);
or U48183 (N_48183,N_34744,N_37020);
nand U48184 (N_48184,N_36485,N_39587);
nor U48185 (N_48185,N_32299,N_37565);
and U48186 (N_48186,N_37275,N_34075);
nand U48187 (N_48187,N_36351,N_31462);
and U48188 (N_48188,N_30066,N_34914);
and U48189 (N_48189,N_34989,N_36464);
or U48190 (N_48190,N_39495,N_32422);
and U48191 (N_48191,N_39752,N_32217);
and U48192 (N_48192,N_38357,N_35039);
and U48193 (N_48193,N_33469,N_38562);
and U48194 (N_48194,N_38198,N_34377);
nor U48195 (N_48195,N_32050,N_37584);
xor U48196 (N_48196,N_39574,N_33521);
nand U48197 (N_48197,N_36650,N_38105);
or U48198 (N_48198,N_32346,N_30809);
nand U48199 (N_48199,N_39805,N_39744);
nor U48200 (N_48200,N_34035,N_33668);
or U48201 (N_48201,N_37541,N_35170);
and U48202 (N_48202,N_34229,N_39987);
and U48203 (N_48203,N_31579,N_34279);
nor U48204 (N_48204,N_38077,N_34793);
nor U48205 (N_48205,N_32271,N_33152);
or U48206 (N_48206,N_35438,N_38504);
xor U48207 (N_48207,N_34224,N_38923);
and U48208 (N_48208,N_35208,N_32499);
and U48209 (N_48209,N_33649,N_36178);
nand U48210 (N_48210,N_33611,N_30839);
or U48211 (N_48211,N_30397,N_30489);
or U48212 (N_48212,N_34953,N_36860);
nand U48213 (N_48213,N_32431,N_35687);
and U48214 (N_48214,N_37782,N_38110);
and U48215 (N_48215,N_37895,N_30335);
and U48216 (N_48216,N_36412,N_31499);
nand U48217 (N_48217,N_32795,N_39795);
xnor U48218 (N_48218,N_30220,N_30705);
and U48219 (N_48219,N_35801,N_35162);
xnor U48220 (N_48220,N_39717,N_36473);
or U48221 (N_48221,N_30287,N_34526);
or U48222 (N_48222,N_33829,N_38757);
or U48223 (N_48223,N_34659,N_37224);
xnor U48224 (N_48224,N_36969,N_34780);
and U48225 (N_48225,N_37611,N_32685);
and U48226 (N_48226,N_30510,N_36072);
nand U48227 (N_48227,N_35121,N_39980);
and U48228 (N_48228,N_35955,N_34379);
nor U48229 (N_48229,N_30787,N_35065);
xor U48230 (N_48230,N_39676,N_36160);
nor U48231 (N_48231,N_36153,N_37286);
xnor U48232 (N_48232,N_36016,N_33784);
xnor U48233 (N_48233,N_36095,N_35955);
nand U48234 (N_48234,N_35576,N_36763);
nor U48235 (N_48235,N_39665,N_30723);
nand U48236 (N_48236,N_31037,N_38191);
and U48237 (N_48237,N_34335,N_31299);
nor U48238 (N_48238,N_35735,N_38759);
xor U48239 (N_48239,N_33793,N_30320);
or U48240 (N_48240,N_37376,N_38225);
nand U48241 (N_48241,N_35417,N_37635);
nor U48242 (N_48242,N_39280,N_34969);
xnor U48243 (N_48243,N_33166,N_38047);
xnor U48244 (N_48244,N_34168,N_37125);
or U48245 (N_48245,N_34391,N_34207);
xor U48246 (N_48246,N_37323,N_37243);
and U48247 (N_48247,N_36992,N_38792);
nor U48248 (N_48248,N_35414,N_37677);
xor U48249 (N_48249,N_39460,N_38733);
nand U48250 (N_48250,N_31967,N_32949);
and U48251 (N_48251,N_38649,N_30232);
xor U48252 (N_48252,N_37301,N_30007);
nand U48253 (N_48253,N_36790,N_32120);
and U48254 (N_48254,N_34230,N_34068);
nand U48255 (N_48255,N_32229,N_30469);
and U48256 (N_48256,N_36307,N_31368);
and U48257 (N_48257,N_32488,N_33928);
nand U48258 (N_48258,N_33502,N_38320);
nor U48259 (N_48259,N_32299,N_32939);
or U48260 (N_48260,N_39957,N_33458);
or U48261 (N_48261,N_37539,N_38345);
nor U48262 (N_48262,N_32064,N_32865);
or U48263 (N_48263,N_37905,N_35716);
and U48264 (N_48264,N_31965,N_30740);
and U48265 (N_48265,N_38530,N_38449);
nand U48266 (N_48266,N_32762,N_32454);
nor U48267 (N_48267,N_31363,N_33682);
nor U48268 (N_48268,N_35979,N_38740);
xor U48269 (N_48269,N_35288,N_35938);
xor U48270 (N_48270,N_31797,N_35722);
xnor U48271 (N_48271,N_38938,N_33026);
nand U48272 (N_48272,N_38890,N_36915);
or U48273 (N_48273,N_38050,N_31883);
and U48274 (N_48274,N_36770,N_35959);
or U48275 (N_48275,N_39821,N_33674);
and U48276 (N_48276,N_36970,N_39491);
nand U48277 (N_48277,N_37742,N_32860);
or U48278 (N_48278,N_39170,N_35458);
or U48279 (N_48279,N_32001,N_30946);
nor U48280 (N_48280,N_37227,N_34713);
xor U48281 (N_48281,N_38550,N_38117);
and U48282 (N_48282,N_33129,N_37590);
and U48283 (N_48283,N_33856,N_39494);
or U48284 (N_48284,N_31937,N_33844);
xnor U48285 (N_48285,N_32297,N_35890);
or U48286 (N_48286,N_32646,N_32968);
or U48287 (N_48287,N_30785,N_37258);
and U48288 (N_48288,N_33184,N_39910);
and U48289 (N_48289,N_37327,N_34330);
xor U48290 (N_48290,N_34368,N_38462);
xor U48291 (N_48291,N_35072,N_34154);
nand U48292 (N_48292,N_35265,N_31479);
xnor U48293 (N_48293,N_34744,N_39722);
and U48294 (N_48294,N_39949,N_36378);
or U48295 (N_48295,N_39243,N_36898);
or U48296 (N_48296,N_36009,N_34732);
nor U48297 (N_48297,N_39453,N_39088);
nand U48298 (N_48298,N_33089,N_36399);
nor U48299 (N_48299,N_32004,N_30224);
nor U48300 (N_48300,N_33174,N_36630);
nor U48301 (N_48301,N_39269,N_30134);
nand U48302 (N_48302,N_39635,N_37255);
nand U48303 (N_48303,N_32379,N_39682);
or U48304 (N_48304,N_32095,N_34803);
and U48305 (N_48305,N_30901,N_39454);
and U48306 (N_48306,N_30538,N_39586);
nor U48307 (N_48307,N_31926,N_38947);
nor U48308 (N_48308,N_30066,N_32099);
nand U48309 (N_48309,N_36182,N_36021);
nor U48310 (N_48310,N_38978,N_31614);
or U48311 (N_48311,N_36726,N_35613);
nand U48312 (N_48312,N_39106,N_32733);
and U48313 (N_48313,N_37323,N_32626);
or U48314 (N_48314,N_30471,N_32898);
and U48315 (N_48315,N_38281,N_31207);
nand U48316 (N_48316,N_31124,N_31512);
xnor U48317 (N_48317,N_32767,N_36277);
nand U48318 (N_48318,N_38064,N_38313);
or U48319 (N_48319,N_35406,N_36902);
xor U48320 (N_48320,N_31442,N_34427);
or U48321 (N_48321,N_36531,N_31601);
xnor U48322 (N_48322,N_32430,N_34508);
nor U48323 (N_48323,N_32761,N_35563);
and U48324 (N_48324,N_30434,N_30757);
nand U48325 (N_48325,N_37444,N_33694);
nand U48326 (N_48326,N_39878,N_37904);
xor U48327 (N_48327,N_37870,N_34464);
nand U48328 (N_48328,N_34750,N_37984);
nand U48329 (N_48329,N_30246,N_37798);
or U48330 (N_48330,N_31105,N_33981);
nand U48331 (N_48331,N_39827,N_34345);
and U48332 (N_48332,N_32438,N_37338);
nand U48333 (N_48333,N_34410,N_37762);
xor U48334 (N_48334,N_35823,N_32699);
xnor U48335 (N_48335,N_34933,N_36436);
nand U48336 (N_48336,N_32783,N_36770);
and U48337 (N_48337,N_39284,N_30892);
xnor U48338 (N_48338,N_31104,N_34845);
or U48339 (N_48339,N_39073,N_33506);
nand U48340 (N_48340,N_34777,N_39862);
nand U48341 (N_48341,N_39953,N_38719);
and U48342 (N_48342,N_30349,N_30399);
xor U48343 (N_48343,N_33634,N_30183);
and U48344 (N_48344,N_38068,N_32330);
nand U48345 (N_48345,N_31967,N_32933);
nand U48346 (N_48346,N_31130,N_33578);
nor U48347 (N_48347,N_34558,N_34743);
or U48348 (N_48348,N_33289,N_30099);
nand U48349 (N_48349,N_36879,N_36480);
nor U48350 (N_48350,N_36784,N_37862);
xnor U48351 (N_48351,N_33202,N_31612);
or U48352 (N_48352,N_31805,N_32223);
nor U48353 (N_48353,N_36516,N_36213);
nor U48354 (N_48354,N_39156,N_34190);
and U48355 (N_48355,N_38083,N_32005);
nor U48356 (N_48356,N_31964,N_37761);
or U48357 (N_48357,N_32314,N_31189);
or U48358 (N_48358,N_35144,N_39582);
or U48359 (N_48359,N_33633,N_32108);
and U48360 (N_48360,N_39134,N_31521);
nor U48361 (N_48361,N_34698,N_37374);
xor U48362 (N_48362,N_35743,N_37330);
and U48363 (N_48363,N_33788,N_37061);
nor U48364 (N_48364,N_34479,N_38912);
nand U48365 (N_48365,N_33076,N_37461);
xor U48366 (N_48366,N_37418,N_32855);
xor U48367 (N_48367,N_36952,N_39782);
and U48368 (N_48368,N_38274,N_32430);
nor U48369 (N_48369,N_39436,N_30830);
nor U48370 (N_48370,N_30176,N_30714);
or U48371 (N_48371,N_39341,N_31480);
or U48372 (N_48372,N_35391,N_35098);
nor U48373 (N_48373,N_35240,N_38620);
nand U48374 (N_48374,N_34888,N_31281);
nor U48375 (N_48375,N_30577,N_33614);
and U48376 (N_48376,N_32639,N_30470);
and U48377 (N_48377,N_39531,N_35946);
and U48378 (N_48378,N_39131,N_37985);
nor U48379 (N_48379,N_39953,N_31977);
nand U48380 (N_48380,N_31518,N_34456);
or U48381 (N_48381,N_38687,N_32203);
or U48382 (N_48382,N_37092,N_34044);
xnor U48383 (N_48383,N_34855,N_35317);
and U48384 (N_48384,N_30731,N_37719);
and U48385 (N_48385,N_34051,N_34267);
nor U48386 (N_48386,N_34303,N_32147);
xor U48387 (N_48387,N_36017,N_39905);
nand U48388 (N_48388,N_39263,N_33505);
and U48389 (N_48389,N_35230,N_36261);
and U48390 (N_48390,N_35012,N_35975);
nand U48391 (N_48391,N_34712,N_34557);
nor U48392 (N_48392,N_33218,N_31190);
or U48393 (N_48393,N_32329,N_30151);
xor U48394 (N_48394,N_37090,N_38163);
xor U48395 (N_48395,N_33815,N_30521);
nand U48396 (N_48396,N_35237,N_38356);
and U48397 (N_48397,N_30188,N_36878);
or U48398 (N_48398,N_33425,N_39734);
nor U48399 (N_48399,N_38579,N_35337);
nor U48400 (N_48400,N_39342,N_32844);
nor U48401 (N_48401,N_38099,N_31444);
nor U48402 (N_48402,N_31332,N_32591);
or U48403 (N_48403,N_37024,N_33846);
xor U48404 (N_48404,N_32615,N_30730);
nor U48405 (N_48405,N_32525,N_36003);
and U48406 (N_48406,N_33638,N_33755);
and U48407 (N_48407,N_30381,N_36315);
or U48408 (N_48408,N_31537,N_37343);
or U48409 (N_48409,N_33347,N_39238);
nand U48410 (N_48410,N_39169,N_38645);
xnor U48411 (N_48411,N_30032,N_32264);
or U48412 (N_48412,N_37301,N_32724);
nor U48413 (N_48413,N_37955,N_31705);
nand U48414 (N_48414,N_32087,N_39402);
xor U48415 (N_48415,N_31002,N_38383);
nor U48416 (N_48416,N_31894,N_34932);
xnor U48417 (N_48417,N_37959,N_35508);
nand U48418 (N_48418,N_39039,N_31964);
or U48419 (N_48419,N_39032,N_36411);
nor U48420 (N_48420,N_39101,N_33466);
and U48421 (N_48421,N_37444,N_34646);
xnor U48422 (N_48422,N_39126,N_35343);
or U48423 (N_48423,N_30792,N_39021);
and U48424 (N_48424,N_39634,N_32823);
xor U48425 (N_48425,N_33818,N_36711);
or U48426 (N_48426,N_36730,N_38878);
and U48427 (N_48427,N_37155,N_36857);
xor U48428 (N_48428,N_30909,N_32965);
nor U48429 (N_48429,N_35009,N_39684);
or U48430 (N_48430,N_36040,N_31733);
and U48431 (N_48431,N_30182,N_33318);
nand U48432 (N_48432,N_31130,N_34051);
or U48433 (N_48433,N_34676,N_35748);
and U48434 (N_48434,N_36757,N_35255);
nand U48435 (N_48435,N_37974,N_33948);
nor U48436 (N_48436,N_35426,N_34238);
and U48437 (N_48437,N_37920,N_30185);
or U48438 (N_48438,N_39938,N_34577);
xor U48439 (N_48439,N_33969,N_30380);
nor U48440 (N_48440,N_32048,N_34808);
nor U48441 (N_48441,N_31123,N_39564);
nor U48442 (N_48442,N_33020,N_32570);
xnor U48443 (N_48443,N_31577,N_30482);
xor U48444 (N_48444,N_39210,N_32002);
nor U48445 (N_48445,N_39789,N_33884);
nand U48446 (N_48446,N_35978,N_31704);
nor U48447 (N_48447,N_31885,N_34154);
nand U48448 (N_48448,N_39717,N_30317);
or U48449 (N_48449,N_33709,N_38643);
and U48450 (N_48450,N_37737,N_38658);
and U48451 (N_48451,N_36504,N_31219);
nor U48452 (N_48452,N_35205,N_31719);
xor U48453 (N_48453,N_33625,N_32669);
or U48454 (N_48454,N_37916,N_30336);
xor U48455 (N_48455,N_35861,N_36865);
and U48456 (N_48456,N_34897,N_38941);
xor U48457 (N_48457,N_33906,N_30946);
nand U48458 (N_48458,N_37013,N_39080);
and U48459 (N_48459,N_38786,N_38491);
or U48460 (N_48460,N_33097,N_34741);
nand U48461 (N_48461,N_37218,N_30937);
nor U48462 (N_48462,N_30084,N_39100);
or U48463 (N_48463,N_39487,N_33440);
or U48464 (N_48464,N_34001,N_36070);
and U48465 (N_48465,N_36370,N_31048);
nand U48466 (N_48466,N_39195,N_36397);
nand U48467 (N_48467,N_30922,N_31596);
nor U48468 (N_48468,N_34634,N_34498);
and U48469 (N_48469,N_31495,N_38524);
or U48470 (N_48470,N_38400,N_35857);
nand U48471 (N_48471,N_33780,N_30998);
nor U48472 (N_48472,N_31640,N_38418);
nand U48473 (N_48473,N_38505,N_35281);
nor U48474 (N_48474,N_36211,N_39943);
nand U48475 (N_48475,N_35504,N_34335);
or U48476 (N_48476,N_33775,N_38945);
nor U48477 (N_48477,N_39107,N_37105);
and U48478 (N_48478,N_32188,N_37124);
nor U48479 (N_48479,N_34690,N_35692);
or U48480 (N_48480,N_38160,N_31659);
or U48481 (N_48481,N_38635,N_33040);
or U48482 (N_48482,N_37466,N_34352);
xor U48483 (N_48483,N_31200,N_38978);
and U48484 (N_48484,N_33890,N_30964);
or U48485 (N_48485,N_32359,N_33763);
and U48486 (N_48486,N_34270,N_38889);
and U48487 (N_48487,N_39393,N_33839);
xor U48488 (N_48488,N_32324,N_31814);
xor U48489 (N_48489,N_35241,N_36411);
nor U48490 (N_48490,N_39681,N_34482);
nand U48491 (N_48491,N_38531,N_39052);
nand U48492 (N_48492,N_37657,N_32183);
nand U48493 (N_48493,N_34497,N_32203);
nor U48494 (N_48494,N_32854,N_36524);
xnor U48495 (N_48495,N_36760,N_39660);
or U48496 (N_48496,N_31516,N_31915);
and U48497 (N_48497,N_34992,N_32499);
or U48498 (N_48498,N_32225,N_33355);
and U48499 (N_48499,N_35450,N_34540);
nor U48500 (N_48500,N_34424,N_32454);
and U48501 (N_48501,N_33086,N_33267);
or U48502 (N_48502,N_35833,N_35754);
nor U48503 (N_48503,N_33652,N_38691);
nand U48504 (N_48504,N_31364,N_33348);
xnor U48505 (N_48505,N_32032,N_33558);
nor U48506 (N_48506,N_34578,N_37072);
or U48507 (N_48507,N_34459,N_30707);
or U48508 (N_48508,N_38643,N_38706);
or U48509 (N_48509,N_30079,N_37574);
xor U48510 (N_48510,N_30162,N_32947);
nand U48511 (N_48511,N_38174,N_31881);
xnor U48512 (N_48512,N_39188,N_33686);
or U48513 (N_48513,N_33598,N_31176);
nand U48514 (N_48514,N_35998,N_39948);
xnor U48515 (N_48515,N_36703,N_31236);
and U48516 (N_48516,N_37492,N_33480);
nor U48517 (N_48517,N_35591,N_32329);
or U48518 (N_48518,N_31522,N_36453);
xor U48519 (N_48519,N_30623,N_37649);
xor U48520 (N_48520,N_33092,N_34717);
or U48521 (N_48521,N_35923,N_37818);
and U48522 (N_48522,N_39408,N_30224);
and U48523 (N_48523,N_38364,N_38904);
xnor U48524 (N_48524,N_36676,N_38868);
xnor U48525 (N_48525,N_32130,N_34535);
or U48526 (N_48526,N_30193,N_38347);
nor U48527 (N_48527,N_37915,N_30990);
and U48528 (N_48528,N_32459,N_32882);
nor U48529 (N_48529,N_36499,N_39282);
xor U48530 (N_48530,N_37606,N_33811);
nand U48531 (N_48531,N_35893,N_33097);
xor U48532 (N_48532,N_37956,N_39150);
nor U48533 (N_48533,N_39972,N_33021);
nand U48534 (N_48534,N_37636,N_36502);
and U48535 (N_48535,N_32270,N_30589);
or U48536 (N_48536,N_34324,N_38858);
and U48537 (N_48537,N_39660,N_33252);
nand U48538 (N_48538,N_34554,N_33867);
nand U48539 (N_48539,N_33838,N_37973);
xnor U48540 (N_48540,N_37146,N_37531);
and U48541 (N_48541,N_34675,N_37079);
nor U48542 (N_48542,N_38003,N_38948);
nor U48543 (N_48543,N_33717,N_38506);
nand U48544 (N_48544,N_35295,N_30483);
nand U48545 (N_48545,N_30873,N_38717);
xor U48546 (N_48546,N_35293,N_39109);
xor U48547 (N_48547,N_30030,N_38868);
or U48548 (N_48548,N_39683,N_34348);
nand U48549 (N_48549,N_31716,N_34185);
nor U48550 (N_48550,N_34129,N_36924);
nand U48551 (N_48551,N_34908,N_34330);
and U48552 (N_48552,N_37783,N_33106);
nor U48553 (N_48553,N_30520,N_39545);
nor U48554 (N_48554,N_31680,N_39052);
nand U48555 (N_48555,N_36616,N_39421);
and U48556 (N_48556,N_32736,N_36392);
nor U48557 (N_48557,N_34326,N_39276);
nor U48558 (N_48558,N_37719,N_33191);
or U48559 (N_48559,N_36827,N_31787);
xor U48560 (N_48560,N_33517,N_37950);
xor U48561 (N_48561,N_35678,N_30969);
xor U48562 (N_48562,N_35639,N_34009);
xnor U48563 (N_48563,N_31783,N_31053);
and U48564 (N_48564,N_39064,N_38447);
and U48565 (N_48565,N_30159,N_34682);
and U48566 (N_48566,N_39129,N_37369);
nand U48567 (N_48567,N_31563,N_38751);
nand U48568 (N_48568,N_38264,N_39083);
nand U48569 (N_48569,N_39635,N_31721);
or U48570 (N_48570,N_33651,N_39492);
nor U48571 (N_48571,N_39663,N_37172);
or U48572 (N_48572,N_31854,N_36313);
and U48573 (N_48573,N_39211,N_39314);
xnor U48574 (N_48574,N_39481,N_39947);
nand U48575 (N_48575,N_34249,N_39747);
nand U48576 (N_48576,N_34448,N_30451);
and U48577 (N_48577,N_32545,N_38649);
and U48578 (N_48578,N_35923,N_31993);
nor U48579 (N_48579,N_34663,N_38540);
nor U48580 (N_48580,N_38175,N_37600);
or U48581 (N_48581,N_39232,N_34923);
nor U48582 (N_48582,N_30451,N_32772);
nor U48583 (N_48583,N_35570,N_38408);
nand U48584 (N_48584,N_36247,N_35200);
nand U48585 (N_48585,N_32286,N_35319);
xnor U48586 (N_48586,N_33681,N_30756);
xor U48587 (N_48587,N_31049,N_34523);
or U48588 (N_48588,N_33213,N_38620);
xor U48589 (N_48589,N_38404,N_33062);
nor U48590 (N_48590,N_37976,N_33414);
and U48591 (N_48591,N_30708,N_38044);
and U48592 (N_48592,N_34991,N_39978);
nand U48593 (N_48593,N_33938,N_39065);
and U48594 (N_48594,N_38519,N_35881);
nand U48595 (N_48595,N_37832,N_32673);
xor U48596 (N_48596,N_35278,N_31488);
and U48597 (N_48597,N_32704,N_37457);
nand U48598 (N_48598,N_34460,N_31986);
xor U48599 (N_48599,N_32347,N_32338);
or U48600 (N_48600,N_36067,N_32444);
nand U48601 (N_48601,N_37872,N_39350);
nand U48602 (N_48602,N_36083,N_38790);
xnor U48603 (N_48603,N_30745,N_39826);
xnor U48604 (N_48604,N_39474,N_32211);
and U48605 (N_48605,N_37632,N_36035);
nor U48606 (N_48606,N_38231,N_34329);
and U48607 (N_48607,N_39015,N_37259);
and U48608 (N_48608,N_32748,N_38318);
or U48609 (N_48609,N_39991,N_36361);
and U48610 (N_48610,N_36550,N_34899);
nand U48611 (N_48611,N_35865,N_32468);
or U48612 (N_48612,N_37538,N_33791);
or U48613 (N_48613,N_30446,N_35696);
nor U48614 (N_48614,N_35095,N_37869);
nor U48615 (N_48615,N_35185,N_36455);
nor U48616 (N_48616,N_34183,N_31477);
and U48617 (N_48617,N_36514,N_31029);
or U48618 (N_48618,N_32502,N_36414);
or U48619 (N_48619,N_30475,N_39442);
nor U48620 (N_48620,N_33886,N_37116);
nand U48621 (N_48621,N_31202,N_31707);
nor U48622 (N_48622,N_33273,N_36879);
nor U48623 (N_48623,N_31745,N_33393);
nand U48624 (N_48624,N_37750,N_36977);
nand U48625 (N_48625,N_34194,N_35955);
or U48626 (N_48626,N_32146,N_31583);
or U48627 (N_48627,N_37116,N_33724);
nand U48628 (N_48628,N_30549,N_30969);
nand U48629 (N_48629,N_35293,N_37859);
or U48630 (N_48630,N_36882,N_35112);
or U48631 (N_48631,N_30147,N_33724);
xor U48632 (N_48632,N_39787,N_34717);
xor U48633 (N_48633,N_38119,N_34580);
nor U48634 (N_48634,N_36151,N_37168);
nor U48635 (N_48635,N_31555,N_34858);
nor U48636 (N_48636,N_34235,N_33782);
or U48637 (N_48637,N_39254,N_31284);
or U48638 (N_48638,N_36450,N_39023);
nor U48639 (N_48639,N_30521,N_34755);
or U48640 (N_48640,N_38391,N_36272);
xnor U48641 (N_48641,N_39621,N_37134);
and U48642 (N_48642,N_39969,N_33449);
xnor U48643 (N_48643,N_37537,N_31126);
nor U48644 (N_48644,N_38049,N_38562);
xnor U48645 (N_48645,N_35638,N_39278);
or U48646 (N_48646,N_33788,N_30485);
and U48647 (N_48647,N_35224,N_33482);
xnor U48648 (N_48648,N_32878,N_38793);
nor U48649 (N_48649,N_35030,N_36427);
nor U48650 (N_48650,N_32363,N_30971);
or U48651 (N_48651,N_33750,N_32996);
nor U48652 (N_48652,N_33990,N_32827);
and U48653 (N_48653,N_33652,N_31472);
nand U48654 (N_48654,N_30315,N_33318);
xor U48655 (N_48655,N_37832,N_33038);
or U48656 (N_48656,N_31457,N_33760);
xor U48657 (N_48657,N_35939,N_32387);
nand U48658 (N_48658,N_37846,N_35890);
or U48659 (N_48659,N_39231,N_39280);
nand U48660 (N_48660,N_32264,N_31478);
nor U48661 (N_48661,N_35051,N_39336);
nand U48662 (N_48662,N_30720,N_32134);
nand U48663 (N_48663,N_31581,N_38642);
nor U48664 (N_48664,N_39224,N_30273);
and U48665 (N_48665,N_31610,N_32270);
xor U48666 (N_48666,N_36214,N_37482);
or U48667 (N_48667,N_34594,N_32520);
nor U48668 (N_48668,N_34299,N_36156);
nor U48669 (N_48669,N_33831,N_38884);
and U48670 (N_48670,N_33102,N_37856);
or U48671 (N_48671,N_34874,N_39978);
nand U48672 (N_48672,N_37367,N_31855);
or U48673 (N_48673,N_36887,N_37355);
nand U48674 (N_48674,N_38056,N_34943);
xnor U48675 (N_48675,N_34719,N_38437);
nand U48676 (N_48676,N_33827,N_31850);
or U48677 (N_48677,N_33211,N_34897);
nor U48678 (N_48678,N_31603,N_32109);
and U48679 (N_48679,N_38651,N_35664);
nor U48680 (N_48680,N_34989,N_34769);
and U48681 (N_48681,N_30069,N_39782);
xnor U48682 (N_48682,N_33560,N_37024);
xnor U48683 (N_48683,N_39072,N_34075);
nand U48684 (N_48684,N_36373,N_31116);
nand U48685 (N_48685,N_31188,N_30430);
and U48686 (N_48686,N_39373,N_35675);
or U48687 (N_48687,N_38349,N_39409);
xor U48688 (N_48688,N_39942,N_38815);
xnor U48689 (N_48689,N_31507,N_39997);
nor U48690 (N_48690,N_38987,N_33417);
or U48691 (N_48691,N_30172,N_36322);
and U48692 (N_48692,N_36268,N_32293);
nand U48693 (N_48693,N_34788,N_30062);
and U48694 (N_48694,N_37570,N_32176);
and U48695 (N_48695,N_36740,N_33281);
xor U48696 (N_48696,N_39437,N_33246);
nand U48697 (N_48697,N_32612,N_37306);
nand U48698 (N_48698,N_32198,N_36597);
nand U48699 (N_48699,N_32094,N_30343);
and U48700 (N_48700,N_37353,N_33870);
nor U48701 (N_48701,N_31198,N_37804);
nor U48702 (N_48702,N_34839,N_36689);
xor U48703 (N_48703,N_33799,N_35482);
and U48704 (N_48704,N_36111,N_39351);
nor U48705 (N_48705,N_31585,N_39518);
xnor U48706 (N_48706,N_37726,N_36457);
or U48707 (N_48707,N_31382,N_38680);
and U48708 (N_48708,N_34509,N_35987);
nor U48709 (N_48709,N_31822,N_31741);
nand U48710 (N_48710,N_35030,N_38371);
or U48711 (N_48711,N_37878,N_31395);
or U48712 (N_48712,N_39947,N_37304);
nand U48713 (N_48713,N_37404,N_30785);
and U48714 (N_48714,N_37450,N_35918);
nand U48715 (N_48715,N_36272,N_31014);
nor U48716 (N_48716,N_30850,N_38347);
xor U48717 (N_48717,N_31690,N_37056);
nand U48718 (N_48718,N_33574,N_32555);
nor U48719 (N_48719,N_39386,N_36524);
nor U48720 (N_48720,N_37800,N_31048);
nand U48721 (N_48721,N_34811,N_35137);
and U48722 (N_48722,N_30849,N_34572);
xor U48723 (N_48723,N_35584,N_35613);
or U48724 (N_48724,N_38344,N_34364);
or U48725 (N_48725,N_30615,N_39571);
or U48726 (N_48726,N_39559,N_35548);
nand U48727 (N_48727,N_33478,N_31538);
and U48728 (N_48728,N_38107,N_38053);
nor U48729 (N_48729,N_39444,N_38212);
xnor U48730 (N_48730,N_38484,N_35606);
nand U48731 (N_48731,N_34840,N_30770);
xnor U48732 (N_48732,N_32247,N_34433);
nand U48733 (N_48733,N_32835,N_34024);
nor U48734 (N_48734,N_36920,N_37611);
nor U48735 (N_48735,N_35353,N_36938);
and U48736 (N_48736,N_36379,N_39863);
nand U48737 (N_48737,N_37265,N_33638);
or U48738 (N_48738,N_33524,N_38648);
nor U48739 (N_48739,N_35829,N_38758);
nor U48740 (N_48740,N_39423,N_30535);
and U48741 (N_48741,N_33968,N_39139);
nor U48742 (N_48742,N_32626,N_31349);
xnor U48743 (N_48743,N_36674,N_39386);
nand U48744 (N_48744,N_31549,N_34933);
xnor U48745 (N_48745,N_38089,N_33531);
and U48746 (N_48746,N_33546,N_34528);
nor U48747 (N_48747,N_35174,N_36382);
or U48748 (N_48748,N_32896,N_31903);
nand U48749 (N_48749,N_32306,N_38098);
nand U48750 (N_48750,N_37070,N_32400);
nand U48751 (N_48751,N_31619,N_37561);
nand U48752 (N_48752,N_35775,N_36649);
or U48753 (N_48753,N_33594,N_34157);
and U48754 (N_48754,N_39844,N_31739);
and U48755 (N_48755,N_38287,N_34589);
xor U48756 (N_48756,N_32293,N_34629);
nand U48757 (N_48757,N_35533,N_38557);
nor U48758 (N_48758,N_38457,N_32451);
or U48759 (N_48759,N_39226,N_31688);
nor U48760 (N_48760,N_32953,N_33855);
nor U48761 (N_48761,N_39326,N_38729);
and U48762 (N_48762,N_39299,N_30372);
and U48763 (N_48763,N_30201,N_30804);
nand U48764 (N_48764,N_38928,N_30137);
xor U48765 (N_48765,N_30034,N_37544);
and U48766 (N_48766,N_32878,N_30591);
or U48767 (N_48767,N_33631,N_30184);
nor U48768 (N_48768,N_34115,N_38055);
nor U48769 (N_48769,N_31933,N_34078);
or U48770 (N_48770,N_33197,N_35185);
xor U48771 (N_48771,N_33553,N_34006);
nor U48772 (N_48772,N_39845,N_32170);
and U48773 (N_48773,N_36645,N_35940);
xor U48774 (N_48774,N_36455,N_35551);
or U48775 (N_48775,N_39865,N_34707);
xor U48776 (N_48776,N_37138,N_34829);
nor U48777 (N_48777,N_30869,N_35772);
and U48778 (N_48778,N_37077,N_32539);
nor U48779 (N_48779,N_36013,N_36031);
nor U48780 (N_48780,N_31165,N_30124);
xnor U48781 (N_48781,N_36930,N_30827);
and U48782 (N_48782,N_35724,N_35932);
xnor U48783 (N_48783,N_39756,N_38094);
and U48784 (N_48784,N_37922,N_34829);
nor U48785 (N_48785,N_30092,N_39655);
or U48786 (N_48786,N_32300,N_38193);
nor U48787 (N_48787,N_36339,N_38842);
and U48788 (N_48788,N_30526,N_32317);
xor U48789 (N_48789,N_39350,N_37766);
or U48790 (N_48790,N_36993,N_37653);
xnor U48791 (N_48791,N_33932,N_37414);
xor U48792 (N_48792,N_35968,N_39187);
xor U48793 (N_48793,N_35506,N_32833);
nor U48794 (N_48794,N_32223,N_38844);
and U48795 (N_48795,N_35335,N_35689);
nor U48796 (N_48796,N_33914,N_32579);
nand U48797 (N_48797,N_38712,N_33698);
nand U48798 (N_48798,N_35735,N_32706);
xor U48799 (N_48799,N_38504,N_35881);
nor U48800 (N_48800,N_37286,N_34128);
or U48801 (N_48801,N_39299,N_39158);
nor U48802 (N_48802,N_33290,N_31911);
nand U48803 (N_48803,N_30060,N_32251);
nor U48804 (N_48804,N_35990,N_30348);
nand U48805 (N_48805,N_39542,N_35877);
xnor U48806 (N_48806,N_34903,N_32461);
or U48807 (N_48807,N_39995,N_36322);
or U48808 (N_48808,N_36554,N_30511);
or U48809 (N_48809,N_36011,N_37435);
and U48810 (N_48810,N_38383,N_33994);
nand U48811 (N_48811,N_38346,N_39601);
nand U48812 (N_48812,N_38041,N_32997);
xor U48813 (N_48813,N_35795,N_32247);
and U48814 (N_48814,N_34347,N_37045);
nor U48815 (N_48815,N_38700,N_37849);
and U48816 (N_48816,N_39027,N_33244);
nand U48817 (N_48817,N_34399,N_38559);
or U48818 (N_48818,N_39158,N_38797);
nand U48819 (N_48819,N_31159,N_36916);
or U48820 (N_48820,N_39974,N_38296);
and U48821 (N_48821,N_37834,N_31340);
nand U48822 (N_48822,N_33591,N_35997);
nor U48823 (N_48823,N_30160,N_36356);
xor U48824 (N_48824,N_39223,N_38677);
and U48825 (N_48825,N_34514,N_39874);
xnor U48826 (N_48826,N_37063,N_38193);
or U48827 (N_48827,N_35445,N_36370);
nand U48828 (N_48828,N_32928,N_37497);
xnor U48829 (N_48829,N_37025,N_36132);
nor U48830 (N_48830,N_35786,N_32467);
nor U48831 (N_48831,N_30403,N_39067);
xor U48832 (N_48832,N_35194,N_31271);
xor U48833 (N_48833,N_36682,N_34478);
xor U48834 (N_48834,N_37507,N_35222);
or U48835 (N_48835,N_38444,N_33170);
and U48836 (N_48836,N_31270,N_31847);
nor U48837 (N_48837,N_37482,N_30460);
xor U48838 (N_48838,N_36393,N_38506);
and U48839 (N_48839,N_31117,N_36137);
and U48840 (N_48840,N_36070,N_34916);
xor U48841 (N_48841,N_30314,N_39035);
xnor U48842 (N_48842,N_36834,N_36426);
or U48843 (N_48843,N_36967,N_35744);
nand U48844 (N_48844,N_30675,N_30491);
nor U48845 (N_48845,N_39868,N_32005);
xor U48846 (N_48846,N_31616,N_39525);
and U48847 (N_48847,N_37116,N_36532);
or U48848 (N_48848,N_37609,N_35709);
or U48849 (N_48849,N_31962,N_35742);
xnor U48850 (N_48850,N_33123,N_31258);
or U48851 (N_48851,N_31278,N_32857);
and U48852 (N_48852,N_32673,N_32416);
nand U48853 (N_48853,N_34339,N_38393);
nand U48854 (N_48854,N_34403,N_35712);
nor U48855 (N_48855,N_37763,N_30930);
or U48856 (N_48856,N_33867,N_39891);
nor U48857 (N_48857,N_32840,N_37205);
nand U48858 (N_48858,N_37717,N_36184);
or U48859 (N_48859,N_33480,N_34832);
or U48860 (N_48860,N_36792,N_39634);
nor U48861 (N_48861,N_39608,N_39416);
nor U48862 (N_48862,N_32225,N_35651);
nor U48863 (N_48863,N_36636,N_35854);
xnor U48864 (N_48864,N_38748,N_39625);
nor U48865 (N_48865,N_32622,N_30278);
and U48866 (N_48866,N_39403,N_38219);
or U48867 (N_48867,N_32169,N_33028);
or U48868 (N_48868,N_39758,N_35671);
xor U48869 (N_48869,N_36265,N_34261);
xor U48870 (N_48870,N_36035,N_36083);
xor U48871 (N_48871,N_34636,N_33486);
and U48872 (N_48872,N_32333,N_30205);
or U48873 (N_48873,N_35831,N_32804);
nand U48874 (N_48874,N_34886,N_36295);
nand U48875 (N_48875,N_34468,N_39034);
and U48876 (N_48876,N_34623,N_38069);
nand U48877 (N_48877,N_37947,N_39183);
xor U48878 (N_48878,N_37848,N_37911);
nand U48879 (N_48879,N_34757,N_38806);
nor U48880 (N_48880,N_37245,N_34613);
or U48881 (N_48881,N_34821,N_38455);
or U48882 (N_48882,N_36792,N_31215);
nand U48883 (N_48883,N_38451,N_30274);
nor U48884 (N_48884,N_32911,N_31011);
xnor U48885 (N_48885,N_33608,N_33680);
nand U48886 (N_48886,N_36456,N_31545);
nor U48887 (N_48887,N_34180,N_32098);
nand U48888 (N_48888,N_30063,N_33639);
xor U48889 (N_48889,N_32257,N_34949);
nor U48890 (N_48890,N_39076,N_39270);
nor U48891 (N_48891,N_39604,N_34351);
or U48892 (N_48892,N_32308,N_38368);
nor U48893 (N_48893,N_37008,N_37873);
nor U48894 (N_48894,N_33469,N_30669);
nand U48895 (N_48895,N_34107,N_34993);
or U48896 (N_48896,N_35530,N_39581);
and U48897 (N_48897,N_37445,N_33048);
nand U48898 (N_48898,N_37314,N_36645);
nand U48899 (N_48899,N_34568,N_34617);
nand U48900 (N_48900,N_31635,N_31004);
nand U48901 (N_48901,N_34347,N_33567);
or U48902 (N_48902,N_32209,N_31770);
nor U48903 (N_48903,N_36829,N_34948);
nor U48904 (N_48904,N_37326,N_34389);
or U48905 (N_48905,N_36382,N_37314);
or U48906 (N_48906,N_31229,N_33887);
or U48907 (N_48907,N_36089,N_34196);
xor U48908 (N_48908,N_33561,N_30014);
nand U48909 (N_48909,N_31356,N_35718);
and U48910 (N_48910,N_31054,N_30113);
nor U48911 (N_48911,N_39852,N_32670);
and U48912 (N_48912,N_32194,N_38922);
and U48913 (N_48913,N_33134,N_35937);
or U48914 (N_48914,N_36464,N_31968);
xnor U48915 (N_48915,N_30971,N_37636);
or U48916 (N_48916,N_35899,N_32003);
nand U48917 (N_48917,N_34976,N_39473);
or U48918 (N_48918,N_32549,N_37656);
xor U48919 (N_48919,N_30355,N_35381);
nand U48920 (N_48920,N_33953,N_30400);
xor U48921 (N_48921,N_35060,N_30239);
or U48922 (N_48922,N_36142,N_30839);
nor U48923 (N_48923,N_33822,N_37709);
nor U48924 (N_48924,N_31588,N_31843);
xor U48925 (N_48925,N_33671,N_34734);
nand U48926 (N_48926,N_39649,N_33673);
or U48927 (N_48927,N_30801,N_37501);
xnor U48928 (N_48928,N_34725,N_38599);
or U48929 (N_48929,N_37535,N_34447);
or U48930 (N_48930,N_38045,N_31475);
nor U48931 (N_48931,N_30336,N_30297);
nor U48932 (N_48932,N_35669,N_35895);
or U48933 (N_48933,N_36313,N_35876);
xnor U48934 (N_48934,N_38377,N_30953);
nor U48935 (N_48935,N_31123,N_39235);
and U48936 (N_48936,N_35840,N_36880);
xor U48937 (N_48937,N_39032,N_32008);
nand U48938 (N_48938,N_36126,N_38311);
nor U48939 (N_48939,N_34442,N_35736);
nand U48940 (N_48940,N_31919,N_33777);
nand U48941 (N_48941,N_33890,N_31400);
or U48942 (N_48942,N_37509,N_35474);
nand U48943 (N_48943,N_34923,N_37267);
nor U48944 (N_48944,N_38297,N_33734);
nand U48945 (N_48945,N_31529,N_30464);
nand U48946 (N_48946,N_37611,N_38436);
nand U48947 (N_48947,N_34269,N_35921);
or U48948 (N_48948,N_37656,N_36406);
or U48949 (N_48949,N_39051,N_33294);
nand U48950 (N_48950,N_36677,N_37733);
and U48951 (N_48951,N_32641,N_36005);
nor U48952 (N_48952,N_36398,N_39633);
xor U48953 (N_48953,N_33162,N_39110);
and U48954 (N_48954,N_34193,N_35552);
nand U48955 (N_48955,N_36258,N_36447);
xnor U48956 (N_48956,N_34133,N_36114);
or U48957 (N_48957,N_33667,N_33727);
and U48958 (N_48958,N_38006,N_30397);
nand U48959 (N_48959,N_39365,N_38458);
and U48960 (N_48960,N_36939,N_39571);
nor U48961 (N_48961,N_32313,N_38589);
or U48962 (N_48962,N_39325,N_35684);
xor U48963 (N_48963,N_38228,N_38628);
and U48964 (N_48964,N_31637,N_30300);
nor U48965 (N_48965,N_34144,N_33870);
xnor U48966 (N_48966,N_30280,N_36643);
and U48967 (N_48967,N_39972,N_32755);
xor U48968 (N_48968,N_38070,N_37051);
xor U48969 (N_48969,N_33539,N_30501);
and U48970 (N_48970,N_38146,N_37839);
xor U48971 (N_48971,N_31536,N_32679);
nor U48972 (N_48972,N_36532,N_34004);
or U48973 (N_48973,N_35527,N_31857);
xnor U48974 (N_48974,N_35586,N_36678);
or U48975 (N_48975,N_36834,N_35228);
and U48976 (N_48976,N_38705,N_35830);
and U48977 (N_48977,N_39726,N_38593);
and U48978 (N_48978,N_35241,N_37792);
or U48979 (N_48979,N_34659,N_37205);
or U48980 (N_48980,N_30388,N_32211);
or U48981 (N_48981,N_39203,N_34468);
or U48982 (N_48982,N_38166,N_32016);
and U48983 (N_48983,N_31030,N_36104);
nand U48984 (N_48984,N_38299,N_35656);
nand U48985 (N_48985,N_39309,N_33331);
and U48986 (N_48986,N_37016,N_38721);
nand U48987 (N_48987,N_33075,N_30189);
xor U48988 (N_48988,N_33909,N_36643);
xor U48989 (N_48989,N_32900,N_37070);
and U48990 (N_48990,N_35484,N_36682);
xnor U48991 (N_48991,N_35264,N_34714);
or U48992 (N_48992,N_38952,N_32192);
nand U48993 (N_48993,N_36078,N_31688);
and U48994 (N_48994,N_34499,N_33540);
xnor U48995 (N_48995,N_33120,N_35045);
xnor U48996 (N_48996,N_30541,N_38612);
and U48997 (N_48997,N_33917,N_30142);
and U48998 (N_48998,N_33431,N_34022);
nor U48999 (N_48999,N_33212,N_34460);
xor U49000 (N_49000,N_36062,N_37530);
nor U49001 (N_49001,N_35559,N_36797);
nor U49002 (N_49002,N_35004,N_35881);
nand U49003 (N_49003,N_39530,N_37324);
and U49004 (N_49004,N_32325,N_30324);
xor U49005 (N_49005,N_37377,N_31750);
xor U49006 (N_49006,N_37798,N_32949);
or U49007 (N_49007,N_31590,N_34586);
xor U49008 (N_49008,N_39213,N_39884);
nor U49009 (N_49009,N_37287,N_35232);
nand U49010 (N_49010,N_39027,N_33836);
xnor U49011 (N_49011,N_38063,N_30182);
or U49012 (N_49012,N_31898,N_32185);
or U49013 (N_49013,N_35770,N_37247);
or U49014 (N_49014,N_35009,N_31905);
and U49015 (N_49015,N_36218,N_31496);
or U49016 (N_49016,N_36976,N_32349);
or U49017 (N_49017,N_33471,N_31860);
nand U49018 (N_49018,N_32421,N_35652);
or U49019 (N_49019,N_34413,N_39933);
or U49020 (N_49020,N_38399,N_35650);
and U49021 (N_49021,N_39522,N_36753);
nor U49022 (N_49022,N_34270,N_37791);
nand U49023 (N_49023,N_36710,N_38950);
xnor U49024 (N_49024,N_38559,N_38225);
nand U49025 (N_49025,N_36818,N_31649);
xnor U49026 (N_49026,N_32303,N_32197);
and U49027 (N_49027,N_37514,N_33841);
xnor U49028 (N_49028,N_31824,N_39822);
nor U49029 (N_49029,N_38706,N_33118);
xnor U49030 (N_49030,N_36819,N_31441);
or U49031 (N_49031,N_36040,N_39081);
or U49032 (N_49032,N_34103,N_34708);
and U49033 (N_49033,N_32795,N_35539);
and U49034 (N_49034,N_30888,N_39621);
or U49035 (N_49035,N_31951,N_36812);
nand U49036 (N_49036,N_35695,N_35583);
xor U49037 (N_49037,N_34691,N_30226);
and U49038 (N_49038,N_39625,N_31786);
or U49039 (N_49039,N_38220,N_35718);
nand U49040 (N_49040,N_32834,N_33115);
nor U49041 (N_49041,N_32516,N_32510);
xnor U49042 (N_49042,N_35218,N_38198);
or U49043 (N_49043,N_30922,N_36981);
nand U49044 (N_49044,N_37998,N_39080);
nand U49045 (N_49045,N_33882,N_36327);
nand U49046 (N_49046,N_32346,N_35901);
and U49047 (N_49047,N_39166,N_33965);
nand U49048 (N_49048,N_32243,N_39837);
or U49049 (N_49049,N_37773,N_35947);
nand U49050 (N_49050,N_32415,N_35194);
nor U49051 (N_49051,N_32198,N_33604);
xnor U49052 (N_49052,N_30915,N_38302);
xor U49053 (N_49053,N_35388,N_31023);
or U49054 (N_49054,N_37057,N_30190);
nand U49055 (N_49055,N_39232,N_33005);
nor U49056 (N_49056,N_34521,N_32792);
or U49057 (N_49057,N_34909,N_39315);
nand U49058 (N_49058,N_37151,N_36549);
or U49059 (N_49059,N_32583,N_36341);
nand U49060 (N_49060,N_37273,N_34285);
xnor U49061 (N_49061,N_39704,N_39777);
nor U49062 (N_49062,N_36467,N_30365);
xnor U49063 (N_49063,N_31444,N_35192);
and U49064 (N_49064,N_38391,N_34375);
or U49065 (N_49065,N_31583,N_36080);
nor U49066 (N_49066,N_33375,N_39106);
xnor U49067 (N_49067,N_39898,N_36760);
nor U49068 (N_49068,N_32695,N_38506);
nand U49069 (N_49069,N_35820,N_36737);
nor U49070 (N_49070,N_32535,N_35345);
and U49071 (N_49071,N_36445,N_38359);
xnor U49072 (N_49072,N_37701,N_37047);
nor U49073 (N_49073,N_35300,N_36443);
nor U49074 (N_49074,N_36906,N_39000);
or U49075 (N_49075,N_33226,N_34388);
or U49076 (N_49076,N_31634,N_34260);
nand U49077 (N_49077,N_33361,N_38251);
and U49078 (N_49078,N_32360,N_31199);
nor U49079 (N_49079,N_35469,N_38836);
and U49080 (N_49080,N_39640,N_36539);
and U49081 (N_49081,N_39485,N_38155);
xor U49082 (N_49082,N_37779,N_39168);
nand U49083 (N_49083,N_37668,N_30032);
nand U49084 (N_49084,N_38341,N_38282);
nor U49085 (N_49085,N_35493,N_36580);
xnor U49086 (N_49086,N_37051,N_37588);
and U49087 (N_49087,N_32908,N_38843);
nor U49088 (N_49088,N_30169,N_30617);
nand U49089 (N_49089,N_38717,N_30586);
or U49090 (N_49090,N_35107,N_36492);
nor U49091 (N_49091,N_39556,N_32693);
xnor U49092 (N_49092,N_39476,N_32956);
and U49093 (N_49093,N_34949,N_39192);
nand U49094 (N_49094,N_34845,N_36912);
or U49095 (N_49095,N_32076,N_30745);
nand U49096 (N_49096,N_39459,N_38383);
and U49097 (N_49097,N_37741,N_30945);
nand U49098 (N_49098,N_31767,N_33402);
and U49099 (N_49099,N_33707,N_38579);
xor U49100 (N_49100,N_39489,N_33177);
nand U49101 (N_49101,N_31662,N_34697);
and U49102 (N_49102,N_32971,N_39866);
nor U49103 (N_49103,N_34248,N_37232);
nor U49104 (N_49104,N_36511,N_31339);
nor U49105 (N_49105,N_30088,N_38413);
and U49106 (N_49106,N_37756,N_33996);
nor U49107 (N_49107,N_39822,N_35004);
xor U49108 (N_49108,N_31822,N_31381);
nand U49109 (N_49109,N_34721,N_38297);
nand U49110 (N_49110,N_33714,N_32430);
and U49111 (N_49111,N_38960,N_32750);
nand U49112 (N_49112,N_31364,N_39513);
xor U49113 (N_49113,N_37372,N_34192);
nor U49114 (N_49114,N_32189,N_38456);
nor U49115 (N_49115,N_38669,N_34582);
nand U49116 (N_49116,N_32959,N_35070);
xor U49117 (N_49117,N_34230,N_34325);
and U49118 (N_49118,N_36014,N_30928);
or U49119 (N_49119,N_33435,N_37301);
nor U49120 (N_49120,N_33613,N_31533);
nand U49121 (N_49121,N_35130,N_39882);
xnor U49122 (N_49122,N_37082,N_38653);
or U49123 (N_49123,N_33398,N_38603);
xor U49124 (N_49124,N_32155,N_30168);
or U49125 (N_49125,N_39914,N_34385);
and U49126 (N_49126,N_34301,N_33017);
and U49127 (N_49127,N_30271,N_35492);
nor U49128 (N_49128,N_38743,N_38711);
nand U49129 (N_49129,N_39376,N_37028);
or U49130 (N_49130,N_36199,N_34169);
and U49131 (N_49131,N_37289,N_33147);
and U49132 (N_49132,N_37635,N_37538);
xnor U49133 (N_49133,N_34644,N_37700);
or U49134 (N_49134,N_32254,N_31920);
xor U49135 (N_49135,N_38420,N_33077);
nand U49136 (N_49136,N_34902,N_39445);
xor U49137 (N_49137,N_31897,N_34644);
nand U49138 (N_49138,N_30696,N_37350);
nor U49139 (N_49139,N_39180,N_36156);
or U49140 (N_49140,N_37265,N_30117);
nor U49141 (N_49141,N_32496,N_38234);
nand U49142 (N_49142,N_35338,N_30096);
xor U49143 (N_49143,N_38177,N_36633);
xnor U49144 (N_49144,N_32703,N_36461);
and U49145 (N_49145,N_39253,N_31841);
nor U49146 (N_49146,N_38836,N_31089);
nor U49147 (N_49147,N_31724,N_35406);
nor U49148 (N_49148,N_30803,N_30255);
xor U49149 (N_49149,N_37247,N_39165);
xnor U49150 (N_49150,N_30706,N_37465);
nand U49151 (N_49151,N_38325,N_36296);
nand U49152 (N_49152,N_38575,N_37005);
nand U49153 (N_49153,N_34283,N_36885);
xor U49154 (N_49154,N_36508,N_30013);
nor U49155 (N_49155,N_31043,N_38782);
nand U49156 (N_49156,N_36562,N_39895);
or U49157 (N_49157,N_36615,N_31989);
and U49158 (N_49158,N_37863,N_39697);
nand U49159 (N_49159,N_31339,N_38847);
nand U49160 (N_49160,N_32960,N_30409);
nor U49161 (N_49161,N_38955,N_38180);
or U49162 (N_49162,N_34112,N_34289);
nand U49163 (N_49163,N_39357,N_31702);
nand U49164 (N_49164,N_38424,N_35644);
nand U49165 (N_49165,N_39112,N_34413);
xnor U49166 (N_49166,N_33955,N_36359);
or U49167 (N_49167,N_31659,N_33560);
nor U49168 (N_49168,N_39732,N_39138);
and U49169 (N_49169,N_35901,N_36033);
and U49170 (N_49170,N_32429,N_36986);
xnor U49171 (N_49171,N_32243,N_34282);
nand U49172 (N_49172,N_38416,N_32698);
nand U49173 (N_49173,N_37646,N_38028);
nor U49174 (N_49174,N_35583,N_33291);
or U49175 (N_49175,N_30213,N_36163);
and U49176 (N_49176,N_33172,N_38782);
or U49177 (N_49177,N_35354,N_32669);
or U49178 (N_49178,N_31658,N_31228);
and U49179 (N_49179,N_31754,N_30465);
or U49180 (N_49180,N_32915,N_33557);
or U49181 (N_49181,N_36200,N_39363);
nor U49182 (N_49182,N_30858,N_39579);
nand U49183 (N_49183,N_37352,N_39621);
and U49184 (N_49184,N_34154,N_34625);
xor U49185 (N_49185,N_30891,N_36419);
xor U49186 (N_49186,N_32901,N_31860);
or U49187 (N_49187,N_33844,N_33422);
and U49188 (N_49188,N_35951,N_34273);
xor U49189 (N_49189,N_37243,N_31727);
nand U49190 (N_49190,N_30951,N_33331);
xnor U49191 (N_49191,N_38710,N_30975);
and U49192 (N_49192,N_37092,N_30439);
nor U49193 (N_49193,N_36952,N_38487);
xnor U49194 (N_49194,N_30757,N_35523);
and U49195 (N_49195,N_35772,N_37424);
nand U49196 (N_49196,N_39344,N_35102);
xor U49197 (N_49197,N_35387,N_38629);
nor U49198 (N_49198,N_34648,N_38359);
and U49199 (N_49199,N_34341,N_34198);
and U49200 (N_49200,N_37139,N_34849);
nor U49201 (N_49201,N_30795,N_34081);
nand U49202 (N_49202,N_35805,N_34794);
xnor U49203 (N_49203,N_30881,N_34819);
nor U49204 (N_49204,N_32805,N_33072);
xnor U49205 (N_49205,N_30276,N_32752);
nand U49206 (N_49206,N_34447,N_30386);
nor U49207 (N_49207,N_32523,N_31512);
nand U49208 (N_49208,N_30956,N_39422);
nor U49209 (N_49209,N_32236,N_38000);
nor U49210 (N_49210,N_38059,N_33027);
nor U49211 (N_49211,N_30134,N_34006);
or U49212 (N_49212,N_30616,N_36873);
xor U49213 (N_49213,N_30446,N_34022);
nand U49214 (N_49214,N_36417,N_32478);
xor U49215 (N_49215,N_33767,N_37102);
xnor U49216 (N_49216,N_33274,N_33680);
nand U49217 (N_49217,N_39958,N_31972);
nand U49218 (N_49218,N_33033,N_39635);
and U49219 (N_49219,N_37057,N_33887);
nor U49220 (N_49220,N_30841,N_34550);
and U49221 (N_49221,N_36278,N_32207);
nor U49222 (N_49222,N_35126,N_30765);
nor U49223 (N_49223,N_38414,N_38614);
and U49224 (N_49224,N_34176,N_38384);
xor U49225 (N_49225,N_33242,N_38958);
nand U49226 (N_49226,N_31404,N_39474);
nand U49227 (N_49227,N_34478,N_38866);
nor U49228 (N_49228,N_39475,N_33482);
nor U49229 (N_49229,N_39004,N_38357);
xor U49230 (N_49230,N_30923,N_39451);
nand U49231 (N_49231,N_34783,N_37102);
xnor U49232 (N_49232,N_33370,N_37571);
and U49233 (N_49233,N_31497,N_34288);
xor U49234 (N_49234,N_35340,N_33075);
and U49235 (N_49235,N_31219,N_32452);
or U49236 (N_49236,N_35359,N_36044);
xor U49237 (N_49237,N_32541,N_39247);
nor U49238 (N_49238,N_37926,N_37888);
and U49239 (N_49239,N_39174,N_37419);
or U49240 (N_49240,N_38452,N_38752);
or U49241 (N_49241,N_34569,N_36782);
or U49242 (N_49242,N_30554,N_31589);
or U49243 (N_49243,N_34543,N_39038);
or U49244 (N_49244,N_33154,N_33555);
or U49245 (N_49245,N_39190,N_39397);
nor U49246 (N_49246,N_30780,N_37603);
or U49247 (N_49247,N_32156,N_34675);
xnor U49248 (N_49248,N_30058,N_36413);
xor U49249 (N_49249,N_31329,N_38542);
or U49250 (N_49250,N_35405,N_32380);
and U49251 (N_49251,N_34343,N_38336);
nand U49252 (N_49252,N_35593,N_38669);
xnor U49253 (N_49253,N_33057,N_34744);
and U49254 (N_49254,N_31554,N_38242);
and U49255 (N_49255,N_30334,N_37988);
xnor U49256 (N_49256,N_36561,N_33981);
nand U49257 (N_49257,N_34304,N_39476);
and U49258 (N_49258,N_32483,N_34358);
nor U49259 (N_49259,N_31802,N_39259);
nor U49260 (N_49260,N_38012,N_36554);
and U49261 (N_49261,N_37412,N_35593);
nand U49262 (N_49262,N_33424,N_34249);
and U49263 (N_49263,N_37360,N_32686);
nor U49264 (N_49264,N_36208,N_30723);
and U49265 (N_49265,N_32324,N_31992);
nor U49266 (N_49266,N_39245,N_32027);
nand U49267 (N_49267,N_31798,N_35715);
nor U49268 (N_49268,N_35958,N_32430);
or U49269 (N_49269,N_39126,N_33866);
nor U49270 (N_49270,N_31101,N_36075);
nand U49271 (N_49271,N_34653,N_32656);
nor U49272 (N_49272,N_35994,N_30667);
and U49273 (N_49273,N_37745,N_37516);
nand U49274 (N_49274,N_37793,N_32987);
nor U49275 (N_49275,N_31524,N_33557);
nand U49276 (N_49276,N_34038,N_39733);
nor U49277 (N_49277,N_30287,N_30278);
nand U49278 (N_49278,N_34607,N_37511);
nand U49279 (N_49279,N_30906,N_39187);
and U49280 (N_49280,N_31926,N_32947);
nor U49281 (N_49281,N_32842,N_39553);
xnor U49282 (N_49282,N_38833,N_34399);
nand U49283 (N_49283,N_31441,N_37483);
or U49284 (N_49284,N_35714,N_33846);
nand U49285 (N_49285,N_36521,N_32132);
nand U49286 (N_49286,N_31490,N_35499);
and U49287 (N_49287,N_34957,N_38903);
nand U49288 (N_49288,N_38089,N_35541);
nand U49289 (N_49289,N_35962,N_38254);
and U49290 (N_49290,N_34078,N_37824);
nand U49291 (N_49291,N_32873,N_30308);
nand U49292 (N_49292,N_35891,N_38572);
nor U49293 (N_49293,N_38587,N_35784);
nand U49294 (N_49294,N_38153,N_35366);
and U49295 (N_49295,N_32395,N_33318);
and U49296 (N_49296,N_32161,N_39898);
xor U49297 (N_49297,N_32504,N_33997);
nand U49298 (N_49298,N_37230,N_39692);
or U49299 (N_49299,N_34961,N_30026);
nor U49300 (N_49300,N_37418,N_32585);
xnor U49301 (N_49301,N_34557,N_32159);
nand U49302 (N_49302,N_30822,N_39809);
nand U49303 (N_49303,N_37930,N_32719);
nand U49304 (N_49304,N_34111,N_31858);
or U49305 (N_49305,N_34544,N_33729);
nor U49306 (N_49306,N_36261,N_32453);
nand U49307 (N_49307,N_38309,N_34052);
nor U49308 (N_49308,N_36187,N_38822);
and U49309 (N_49309,N_32807,N_30090);
and U49310 (N_49310,N_31505,N_30755);
or U49311 (N_49311,N_30646,N_39157);
nand U49312 (N_49312,N_31726,N_37861);
or U49313 (N_49313,N_30654,N_31702);
nor U49314 (N_49314,N_32605,N_38064);
and U49315 (N_49315,N_30711,N_33070);
nor U49316 (N_49316,N_35025,N_39519);
and U49317 (N_49317,N_36890,N_37422);
xnor U49318 (N_49318,N_33502,N_37174);
nor U49319 (N_49319,N_39533,N_37987);
nor U49320 (N_49320,N_34115,N_34575);
xnor U49321 (N_49321,N_38106,N_37383);
or U49322 (N_49322,N_35811,N_31331);
and U49323 (N_49323,N_39451,N_32732);
or U49324 (N_49324,N_34071,N_34698);
or U49325 (N_49325,N_33679,N_38681);
nand U49326 (N_49326,N_39671,N_39869);
nor U49327 (N_49327,N_37298,N_37058);
and U49328 (N_49328,N_36593,N_38802);
xnor U49329 (N_49329,N_35187,N_36928);
xnor U49330 (N_49330,N_30540,N_31623);
nand U49331 (N_49331,N_31978,N_33358);
nor U49332 (N_49332,N_32013,N_34432);
nor U49333 (N_49333,N_38595,N_39379);
nand U49334 (N_49334,N_31303,N_38674);
xnor U49335 (N_49335,N_38126,N_31725);
or U49336 (N_49336,N_32527,N_34112);
nand U49337 (N_49337,N_35259,N_31648);
nand U49338 (N_49338,N_35410,N_31599);
xor U49339 (N_49339,N_39101,N_36770);
or U49340 (N_49340,N_30598,N_33530);
and U49341 (N_49341,N_39991,N_37244);
and U49342 (N_49342,N_35044,N_38342);
xor U49343 (N_49343,N_38911,N_38279);
nand U49344 (N_49344,N_34353,N_34650);
nor U49345 (N_49345,N_34931,N_38748);
nor U49346 (N_49346,N_39247,N_36034);
nor U49347 (N_49347,N_39886,N_37754);
nand U49348 (N_49348,N_33253,N_34693);
nand U49349 (N_49349,N_37452,N_34278);
or U49350 (N_49350,N_30868,N_32308);
and U49351 (N_49351,N_32273,N_35824);
nor U49352 (N_49352,N_37277,N_35600);
nor U49353 (N_49353,N_36754,N_32146);
nand U49354 (N_49354,N_32694,N_37068);
nor U49355 (N_49355,N_32310,N_36010);
or U49356 (N_49356,N_38674,N_30616);
and U49357 (N_49357,N_35739,N_32611);
or U49358 (N_49358,N_32946,N_32560);
nand U49359 (N_49359,N_36514,N_34543);
nor U49360 (N_49360,N_33158,N_31564);
xnor U49361 (N_49361,N_39804,N_37672);
or U49362 (N_49362,N_35485,N_33613);
and U49363 (N_49363,N_38137,N_34463);
nand U49364 (N_49364,N_39395,N_38523);
and U49365 (N_49365,N_32337,N_38722);
and U49366 (N_49366,N_33635,N_37110);
xor U49367 (N_49367,N_39090,N_30557);
nor U49368 (N_49368,N_38566,N_36544);
and U49369 (N_49369,N_38562,N_34376);
and U49370 (N_49370,N_34036,N_32865);
nand U49371 (N_49371,N_33055,N_30596);
xor U49372 (N_49372,N_35305,N_33509);
nand U49373 (N_49373,N_33160,N_34728);
nand U49374 (N_49374,N_34363,N_30181);
nand U49375 (N_49375,N_32195,N_36023);
nor U49376 (N_49376,N_37184,N_39764);
nand U49377 (N_49377,N_33601,N_31212);
and U49378 (N_49378,N_38711,N_32425);
nand U49379 (N_49379,N_30248,N_39337);
xnor U49380 (N_49380,N_35219,N_36912);
or U49381 (N_49381,N_35304,N_38710);
xor U49382 (N_49382,N_32957,N_39948);
or U49383 (N_49383,N_30425,N_39134);
xor U49384 (N_49384,N_35767,N_34920);
nand U49385 (N_49385,N_34481,N_39743);
nor U49386 (N_49386,N_38155,N_36377);
xnor U49387 (N_49387,N_31952,N_32370);
nand U49388 (N_49388,N_33458,N_34968);
xor U49389 (N_49389,N_37971,N_35987);
nand U49390 (N_49390,N_38827,N_38439);
nor U49391 (N_49391,N_30662,N_38349);
and U49392 (N_49392,N_35091,N_38159);
and U49393 (N_49393,N_32653,N_39195);
or U49394 (N_49394,N_34431,N_32427);
nand U49395 (N_49395,N_32348,N_30674);
nand U49396 (N_49396,N_31857,N_32939);
or U49397 (N_49397,N_39782,N_31518);
nand U49398 (N_49398,N_31303,N_37897);
nand U49399 (N_49399,N_31639,N_39411);
and U49400 (N_49400,N_39762,N_37128);
nor U49401 (N_49401,N_30419,N_35437);
xnor U49402 (N_49402,N_32660,N_31523);
or U49403 (N_49403,N_31995,N_30904);
nand U49404 (N_49404,N_38230,N_39647);
or U49405 (N_49405,N_31385,N_39177);
and U49406 (N_49406,N_39190,N_36110);
or U49407 (N_49407,N_38730,N_32258);
and U49408 (N_49408,N_38849,N_39552);
xor U49409 (N_49409,N_30366,N_37613);
nand U49410 (N_49410,N_34234,N_36272);
or U49411 (N_49411,N_32378,N_32990);
nand U49412 (N_49412,N_31047,N_37555);
nor U49413 (N_49413,N_39607,N_31501);
xnor U49414 (N_49414,N_30799,N_34806);
nor U49415 (N_49415,N_34815,N_33270);
and U49416 (N_49416,N_35901,N_39559);
nand U49417 (N_49417,N_34765,N_36225);
nand U49418 (N_49418,N_31556,N_31470);
xor U49419 (N_49419,N_32884,N_39248);
nor U49420 (N_49420,N_33854,N_35437);
or U49421 (N_49421,N_38446,N_39584);
nand U49422 (N_49422,N_37042,N_39613);
nand U49423 (N_49423,N_33011,N_32590);
and U49424 (N_49424,N_33567,N_39411);
and U49425 (N_49425,N_30890,N_39544);
nor U49426 (N_49426,N_39763,N_39627);
xnor U49427 (N_49427,N_39118,N_36621);
nor U49428 (N_49428,N_37294,N_32234);
nor U49429 (N_49429,N_30122,N_38346);
and U49430 (N_49430,N_39441,N_37409);
xnor U49431 (N_49431,N_32749,N_37669);
nor U49432 (N_49432,N_38186,N_34199);
or U49433 (N_49433,N_31999,N_38954);
nor U49434 (N_49434,N_35468,N_31817);
or U49435 (N_49435,N_31247,N_34996);
nor U49436 (N_49436,N_34781,N_30055);
and U49437 (N_49437,N_38674,N_30456);
and U49438 (N_49438,N_35952,N_37560);
nand U49439 (N_49439,N_38053,N_38488);
nor U49440 (N_49440,N_36317,N_31601);
xnor U49441 (N_49441,N_35737,N_33048);
nor U49442 (N_49442,N_33911,N_37109);
or U49443 (N_49443,N_33414,N_31790);
and U49444 (N_49444,N_31657,N_32980);
nor U49445 (N_49445,N_31394,N_36894);
xor U49446 (N_49446,N_36530,N_37232);
and U49447 (N_49447,N_30353,N_38173);
and U49448 (N_49448,N_36778,N_31292);
xnor U49449 (N_49449,N_31195,N_38718);
nor U49450 (N_49450,N_39789,N_39757);
xor U49451 (N_49451,N_30976,N_31229);
nor U49452 (N_49452,N_34773,N_39563);
nand U49453 (N_49453,N_33547,N_36306);
and U49454 (N_49454,N_39842,N_34357);
or U49455 (N_49455,N_36331,N_36698);
or U49456 (N_49456,N_38111,N_30361);
nor U49457 (N_49457,N_38760,N_37557);
nor U49458 (N_49458,N_35269,N_33931);
or U49459 (N_49459,N_39974,N_34916);
xnor U49460 (N_49460,N_30989,N_38879);
or U49461 (N_49461,N_39903,N_32893);
and U49462 (N_49462,N_36486,N_39098);
and U49463 (N_49463,N_33103,N_36110);
nand U49464 (N_49464,N_38722,N_32126);
nor U49465 (N_49465,N_33700,N_35752);
nor U49466 (N_49466,N_39684,N_31530);
nor U49467 (N_49467,N_39291,N_31047);
nand U49468 (N_49468,N_37106,N_36481);
and U49469 (N_49469,N_37265,N_39676);
and U49470 (N_49470,N_32685,N_34448);
nand U49471 (N_49471,N_32139,N_33930);
nor U49472 (N_49472,N_31093,N_37466);
xnor U49473 (N_49473,N_37870,N_39547);
nand U49474 (N_49474,N_35255,N_37346);
or U49475 (N_49475,N_34491,N_34913);
or U49476 (N_49476,N_39274,N_30940);
and U49477 (N_49477,N_32838,N_38417);
and U49478 (N_49478,N_37166,N_34772);
or U49479 (N_49479,N_30861,N_31241);
and U49480 (N_49480,N_30288,N_30903);
nor U49481 (N_49481,N_36273,N_35415);
nand U49482 (N_49482,N_37664,N_37829);
and U49483 (N_49483,N_32034,N_31917);
nor U49484 (N_49484,N_34745,N_32195);
nand U49485 (N_49485,N_30712,N_33371);
or U49486 (N_49486,N_32850,N_38838);
nor U49487 (N_49487,N_36385,N_32324);
nand U49488 (N_49488,N_39500,N_35831);
or U49489 (N_49489,N_35782,N_30794);
nand U49490 (N_49490,N_33475,N_33358);
xnor U49491 (N_49491,N_39942,N_33067);
nor U49492 (N_49492,N_38103,N_34427);
xor U49493 (N_49493,N_34149,N_33877);
nand U49494 (N_49494,N_39004,N_36917);
or U49495 (N_49495,N_38873,N_32399);
and U49496 (N_49496,N_34470,N_33727);
nor U49497 (N_49497,N_33832,N_35793);
or U49498 (N_49498,N_37083,N_36280);
or U49499 (N_49499,N_33259,N_30894);
nor U49500 (N_49500,N_34908,N_32470);
nand U49501 (N_49501,N_32545,N_37537);
nor U49502 (N_49502,N_30734,N_38509);
nor U49503 (N_49503,N_34264,N_31655);
and U49504 (N_49504,N_33779,N_36828);
or U49505 (N_49505,N_36010,N_39723);
xor U49506 (N_49506,N_36276,N_32319);
and U49507 (N_49507,N_37192,N_37002);
or U49508 (N_49508,N_37867,N_39238);
or U49509 (N_49509,N_36256,N_31641);
or U49510 (N_49510,N_34463,N_34551);
and U49511 (N_49511,N_32885,N_30195);
xor U49512 (N_49512,N_32799,N_34353);
or U49513 (N_49513,N_37187,N_39598);
nor U49514 (N_49514,N_39788,N_33006);
nand U49515 (N_49515,N_32787,N_32364);
and U49516 (N_49516,N_32196,N_35998);
or U49517 (N_49517,N_32149,N_30244);
nor U49518 (N_49518,N_35905,N_31990);
xor U49519 (N_49519,N_34529,N_39437);
nand U49520 (N_49520,N_37173,N_31780);
or U49521 (N_49521,N_30812,N_34391);
xor U49522 (N_49522,N_39585,N_31045);
or U49523 (N_49523,N_33449,N_38851);
nand U49524 (N_49524,N_35453,N_34166);
xnor U49525 (N_49525,N_35142,N_30828);
xor U49526 (N_49526,N_31855,N_38120);
or U49527 (N_49527,N_33669,N_32441);
or U49528 (N_49528,N_33721,N_35885);
nor U49529 (N_49529,N_37859,N_34068);
nand U49530 (N_49530,N_30437,N_35245);
xor U49531 (N_49531,N_35293,N_38270);
nand U49532 (N_49532,N_39810,N_35023);
nand U49533 (N_49533,N_38994,N_39091);
and U49534 (N_49534,N_38001,N_39758);
xnor U49535 (N_49535,N_39073,N_31424);
nor U49536 (N_49536,N_33515,N_32258);
xor U49537 (N_49537,N_35830,N_32315);
xor U49538 (N_49538,N_39281,N_32548);
nand U49539 (N_49539,N_32085,N_34653);
nand U49540 (N_49540,N_39850,N_31489);
and U49541 (N_49541,N_36498,N_32119);
nand U49542 (N_49542,N_32980,N_37191);
and U49543 (N_49543,N_34083,N_39932);
or U49544 (N_49544,N_33227,N_38097);
nand U49545 (N_49545,N_39314,N_39371);
nand U49546 (N_49546,N_31638,N_31342);
nor U49547 (N_49547,N_38006,N_38064);
and U49548 (N_49548,N_36922,N_34651);
nor U49549 (N_49549,N_35876,N_30652);
nor U49550 (N_49550,N_39300,N_36187);
and U49551 (N_49551,N_31781,N_34432);
xnor U49552 (N_49552,N_36263,N_37741);
or U49553 (N_49553,N_32302,N_37529);
xor U49554 (N_49554,N_30477,N_30969);
nand U49555 (N_49555,N_39814,N_30955);
and U49556 (N_49556,N_30930,N_39506);
xnor U49557 (N_49557,N_36827,N_34407);
nand U49558 (N_49558,N_39938,N_36184);
xor U49559 (N_49559,N_34143,N_35025);
xnor U49560 (N_49560,N_36543,N_35566);
nor U49561 (N_49561,N_34710,N_32718);
nor U49562 (N_49562,N_35365,N_31312);
nand U49563 (N_49563,N_34382,N_32415);
and U49564 (N_49564,N_38512,N_36514);
and U49565 (N_49565,N_34118,N_37236);
nor U49566 (N_49566,N_38027,N_39029);
nor U49567 (N_49567,N_34647,N_38687);
or U49568 (N_49568,N_30383,N_30984);
nor U49569 (N_49569,N_34656,N_34197);
xor U49570 (N_49570,N_31565,N_31257);
and U49571 (N_49571,N_36590,N_34543);
nand U49572 (N_49572,N_31021,N_30391);
nor U49573 (N_49573,N_37312,N_31548);
and U49574 (N_49574,N_38756,N_35256);
xnor U49575 (N_49575,N_30055,N_35284);
xor U49576 (N_49576,N_31821,N_39990);
nand U49577 (N_49577,N_36372,N_34498);
nand U49578 (N_49578,N_30713,N_37707);
xnor U49579 (N_49579,N_36771,N_30511);
nor U49580 (N_49580,N_34266,N_37708);
and U49581 (N_49581,N_39510,N_36260);
and U49582 (N_49582,N_36829,N_32530);
nor U49583 (N_49583,N_36903,N_38656);
or U49584 (N_49584,N_38006,N_31329);
or U49585 (N_49585,N_30849,N_37778);
nor U49586 (N_49586,N_37462,N_31149);
nor U49587 (N_49587,N_31313,N_31807);
nand U49588 (N_49588,N_39604,N_35549);
nand U49589 (N_49589,N_35285,N_35555);
or U49590 (N_49590,N_37183,N_34676);
xor U49591 (N_49591,N_39343,N_33208);
or U49592 (N_49592,N_36115,N_31252);
and U49593 (N_49593,N_34550,N_38597);
nand U49594 (N_49594,N_32320,N_31431);
nand U49595 (N_49595,N_36426,N_31573);
nor U49596 (N_49596,N_37780,N_39340);
and U49597 (N_49597,N_33366,N_30057);
or U49598 (N_49598,N_31048,N_39198);
or U49599 (N_49599,N_31854,N_34503);
xor U49600 (N_49600,N_33321,N_39367);
or U49601 (N_49601,N_32323,N_36848);
nand U49602 (N_49602,N_35816,N_36799);
or U49603 (N_49603,N_37203,N_36529);
or U49604 (N_49604,N_34766,N_34681);
nor U49605 (N_49605,N_37162,N_31455);
or U49606 (N_49606,N_33832,N_32028);
nor U49607 (N_49607,N_39759,N_37537);
xor U49608 (N_49608,N_39542,N_32200);
nor U49609 (N_49609,N_33292,N_37702);
xnor U49610 (N_49610,N_35805,N_38155);
xnor U49611 (N_49611,N_39916,N_34261);
nand U49612 (N_49612,N_33144,N_34071);
xor U49613 (N_49613,N_32290,N_30779);
nor U49614 (N_49614,N_35441,N_36064);
nand U49615 (N_49615,N_32349,N_32088);
or U49616 (N_49616,N_33939,N_35026);
xnor U49617 (N_49617,N_38829,N_32662);
xnor U49618 (N_49618,N_35648,N_35530);
nor U49619 (N_49619,N_38296,N_36554);
or U49620 (N_49620,N_34943,N_37211);
xnor U49621 (N_49621,N_35919,N_36176);
and U49622 (N_49622,N_30268,N_36997);
and U49623 (N_49623,N_39571,N_33196);
and U49624 (N_49624,N_39285,N_31471);
nand U49625 (N_49625,N_33457,N_33445);
xor U49626 (N_49626,N_37313,N_36947);
nor U49627 (N_49627,N_31025,N_35966);
or U49628 (N_49628,N_35347,N_37874);
nand U49629 (N_49629,N_35890,N_31585);
or U49630 (N_49630,N_32780,N_36976);
nor U49631 (N_49631,N_31590,N_30157);
and U49632 (N_49632,N_38112,N_38067);
nand U49633 (N_49633,N_32352,N_33724);
xor U49634 (N_49634,N_32513,N_35517);
or U49635 (N_49635,N_30151,N_33576);
nand U49636 (N_49636,N_33030,N_39878);
xnor U49637 (N_49637,N_37109,N_35451);
nor U49638 (N_49638,N_39508,N_35312);
nor U49639 (N_49639,N_38661,N_33505);
or U49640 (N_49640,N_30493,N_33234);
and U49641 (N_49641,N_33825,N_34534);
nor U49642 (N_49642,N_30842,N_39316);
nor U49643 (N_49643,N_30017,N_32965);
nand U49644 (N_49644,N_31823,N_35453);
and U49645 (N_49645,N_31534,N_39517);
xor U49646 (N_49646,N_38569,N_37440);
nand U49647 (N_49647,N_31240,N_33263);
nand U49648 (N_49648,N_35493,N_39553);
and U49649 (N_49649,N_36484,N_38112);
nor U49650 (N_49650,N_38177,N_36323);
nand U49651 (N_49651,N_31500,N_30070);
nand U49652 (N_49652,N_33821,N_36879);
and U49653 (N_49653,N_34790,N_32152);
nand U49654 (N_49654,N_31979,N_32614);
nand U49655 (N_49655,N_33636,N_34280);
and U49656 (N_49656,N_33373,N_34562);
nand U49657 (N_49657,N_35322,N_31710);
xnor U49658 (N_49658,N_33633,N_37009);
and U49659 (N_49659,N_33958,N_32484);
xnor U49660 (N_49660,N_37695,N_35977);
xor U49661 (N_49661,N_39036,N_36114);
nand U49662 (N_49662,N_30719,N_36913);
or U49663 (N_49663,N_37146,N_31618);
or U49664 (N_49664,N_34792,N_30097);
or U49665 (N_49665,N_31103,N_37248);
xnor U49666 (N_49666,N_32558,N_33501);
nand U49667 (N_49667,N_36923,N_38725);
nand U49668 (N_49668,N_32188,N_36348);
nor U49669 (N_49669,N_39324,N_36966);
or U49670 (N_49670,N_34731,N_36576);
nand U49671 (N_49671,N_39684,N_38073);
and U49672 (N_49672,N_37872,N_35256);
nor U49673 (N_49673,N_36388,N_33130);
nor U49674 (N_49674,N_36171,N_39682);
nor U49675 (N_49675,N_38030,N_32940);
xnor U49676 (N_49676,N_35877,N_36801);
nand U49677 (N_49677,N_36972,N_36444);
or U49678 (N_49678,N_36797,N_33135);
or U49679 (N_49679,N_33555,N_31574);
nor U49680 (N_49680,N_33717,N_34675);
and U49681 (N_49681,N_39690,N_34008);
or U49682 (N_49682,N_32023,N_39550);
xnor U49683 (N_49683,N_37125,N_37135);
nand U49684 (N_49684,N_30730,N_33828);
nand U49685 (N_49685,N_36942,N_32115);
nor U49686 (N_49686,N_30146,N_39845);
nor U49687 (N_49687,N_30370,N_31453);
nand U49688 (N_49688,N_35170,N_33533);
nand U49689 (N_49689,N_35501,N_39763);
nor U49690 (N_49690,N_35014,N_35016);
xor U49691 (N_49691,N_33014,N_36954);
and U49692 (N_49692,N_38480,N_30379);
and U49693 (N_49693,N_30719,N_36839);
nand U49694 (N_49694,N_30284,N_34942);
xor U49695 (N_49695,N_35671,N_33852);
xnor U49696 (N_49696,N_35062,N_39241);
or U49697 (N_49697,N_30695,N_38335);
nand U49698 (N_49698,N_35591,N_36261);
nand U49699 (N_49699,N_31718,N_32876);
xor U49700 (N_49700,N_36107,N_37721);
xor U49701 (N_49701,N_30140,N_30978);
or U49702 (N_49702,N_38933,N_32673);
xnor U49703 (N_49703,N_32164,N_38607);
nand U49704 (N_49704,N_32892,N_31275);
nand U49705 (N_49705,N_39113,N_36639);
nor U49706 (N_49706,N_30782,N_31405);
nor U49707 (N_49707,N_39339,N_35457);
xnor U49708 (N_49708,N_38132,N_30982);
xnor U49709 (N_49709,N_36250,N_33372);
nor U49710 (N_49710,N_38248,N_30204);
or U49711 (N_49711,N_32356,N_33482);
xor U49712 (N_49712,N_34662,N_30123);
nor U49713 (N_49713,N_35307,N_39109);
or U49714 (N_49714,N_38627,N_32837);
nand U49715 (N_49715,N_38415,N_31732);
or U49716 (N_49716,N_32151,N_36528);
and U49717 (N_49717,N_32659,N_38263);
or U49718 (N_49718,N_35257,N_33139);
and U49719 (N_49719,N_36168,N_36161);
or U49720 (N_49720,N_35200,N_30501);
or U49721 (N_49721,N_34786,N_32422);
and U49722 (N_49722,N_31282,N_35188);
or U49723 (N_49723,N_32720,N_39488);
xor U49724 (N_49724,N_31435,N_33324);
xor U49725 (N_49725,N_35917,N_36901);
or U49726 (N_49726,N_37127,N_39038);
and U49727 (N_49727,N_35391,N_35223);
nor U49728 (N_49728,N_39651,N_34774);
nand U49729 (N_49729,N_31560,N_30142);
nor U49730 (N_49730,N_30721,N_32952);
and U49731 (N_49731,N_31546,N_32322);
nor U49732 (N_49732,N_34523,N_32741);
or U49733 (N_49733,N_33880,N_32919);
and U49734 (N_49734,N_34372,N_30293);
nor U49735 (N_49735,N_30094,N_30229);
and U49736 (N_49736,N_39448,N_37982);
nor U49737 (N_49737,N_32687,N_34379);
and U49738 (N_49738,N_31267,N_37241);
xor U49739 (N_49739,N_39987,N_32025);
and U49740 (N_49740,N_30831,N_39623);
nor U49741 (N_49741,N_37927,N_32390);
xnor U49742 (N_49742,N_31720,N_32677);
and U49743 (N_49743,N_39709,N_31722);
nand U49744 (N_49744,N_34429,N_34475);
or U49745 (N_49745,N_39743,N_38243);
nor U49746 (N_49746,N_30772,N_32356);
xnor U49747 (N_49747,N_34656,N_36978);
xor U49748 (N_49748,N_35184,N_38989);
nand U49749 (N_49749,N_33821,N_30380);
nand U49750 (N_49750,N_33407,N_35464);
or U49751 (N_49751,N_33426,N_35494);
and U49752 (N_49752,N_31032,N_38964);
xor U49753 (N_49753,N_36318,N_30122);
and U49754 (N_49754,N_34987,N_31383);
and U49755 (N_49755,N_33509,N_34059);
or U49756 (N_49756,N_34389,N_32864);
xor U49757 (N_49757,N_36313,N_39715);
nand U49758 (N_49758,N_35160,N_37755);
or U49759 (N_49759,N_33248,N_35855);
and U49760 (N_49760,N_33701,N_34776);
xor U49761 (N_49761,N_34206,N_38159);
and U49762 (N_49762,N_30815,N_33012);
and U49763 (N_49763,N_31943,N_35191);
or U49764 (N_49764,N_38742,N_39222);
or U49765 (N_49765,N_36401,N_37158);
nand U49766 (N_49766,N_33591,N_33729);
nor U49767 (N_49767,N_35005,N_32488);
and U49768 (N_49768,N_31859,N_39831);
xnor U49769 (N_49769,N_35924,N_38402);
nand U49770 (N_49770,N_30581,N_33253);
nand U49771 (N_49771,N_37697,N_32592);
and U49772 (N_49772,N_32559,N_38637);
nor U49773 (N_49773,N_35092,N_37630);
and U49774 (N_49774,N_30123,N_37984);
nor U49775 (N_49775,N_36458,N_38297);
and U49776 (N_49776,N_30920,N_32557);
and U49777 (N_49777,N_31955,N_35136);
nor U49778 (N_49778,N_37657,N_38280);
nor U49779 (N_49779,N_34633,N_34745);
or U49780 (N_49780,N_36559,N_30195);
xnor U49781 (N_49781,N_30391,N_37741);
or U49782 (N_49782,N_39752,N_38787);
and U49783 (N_49783,N_32530,N_38171);
and U49784 (N_49784,N_33914,N_37549);
xor U49785 (N_49785,N_36195,N_36454);
xnor U49786 (N_49786,N_34015,N_34046);
or U49787 (N_49787,N_39230,N_34680);
nand U49788 (N_49788,N_35593,N_39663);
and U49789 (N_49789,N_33545,N_39827);
or U49790 (N_49790,N_38052,N_35132);
and U49791 (N_49791,N_38290,N_30421);
xnor U49792 (N_49792,N_35020,N_33336);
xor U49793 (N_49793,N_34180,N_33044);
nor U49794 (N_49794,N_33366,N_38703);
nand U49795 (N_49795,N_31599,N_34868);
xnor U49796 (N_49796,N_36891,N_33881);
nand U49797 (N_49797,N_34675,N_39244);
and U49798 (N_49798,N_31241,N_38941);
or U49799 (N_49799,N_34481,N_31540);
nand U49800 (N_49800,N_31827,N_32269);
xnor U49801 (N_49801,N_35116,N_32148);
and U49802 (N_49802,N_31993,N_31999);
and U49803 (N_49803,N_36133,N_31495);
nor U49804 (N_49804,N_38443,N_30674);
and U49805 (N_49805,N_34274,N_31822);
xor U49806 (N_49806,N_36379,N_36487);
xor U49807 (N_49807,N_36631,N_34021);
nor U49808 (N_49808,N_37151,N_34172);
and U49809 (N_49809,N_36003,N_33404);
nand U49810 (N_49810,N_31163,N_33439);
xnor U49811 (N_49811,N_30941,N_33779);
and U49812 (N_49812,N_38604,N_34135);
nor U49813 (N_49813,N_33096,N_32568);
or U49814 (N_49814,N_38156,N_39173);
nor U49815 (N_49815,N_32250,N_39306);
or U49816 (N_49816,N_32893,N_30216);
and U49817 (N_49817,N_39021,N_33582);
nand U49818 (N_49818,N_31227,N_37624);
nor U49819 (N_49819,N_39224,N_32293);
xor U49820 (N_49820,N_39218,N_37399);
and U49821 (N_49821,N_34248,N_39392);
and U49822 (N_49822,N_34572,N_34005);
nand U49823 (N_49823,N_36125,N_32820);
nand U49824 (N_49824,N_38896,N_36351);
xor U49825 (N_49825,N_37077,N_36644);
xnor U49826 (N_49826,N_39521,N_33247);
xor U49827 (N_49827,N_35903,N_36340);
xnor U49828 (N_49828,N_38594,N_37848);
and U49829 (N_49829,N_33577,N_36351);
xnor U49830 (N_49830,N_34461,N_39872);
xnor U49831 (N_49831,N_36273,N_37362);
and U49832 (N_49832,N_34019,N_32262);
nand U49833 (N_49833,N_39833,N_37325);
nand U49834 (N_49834,N_38952,N_37922);
and U49835 (N_49835,N_34109,N_34789);
nor U49836 (N_49836,N_32971,N_30237);
xnor U49837 (N_49837,N_37901,N_38837);
or U49838 (N_49838,N_33382,N_34273);
or U49839 (N_49839,N_33784,N_36768);
and U49840 (N_49840,N_30766,N_31110);
or U49841 (N_49841,N_32731,N_37427);
nor U49842 (N_49842,N_33016,N_33307);
nand U49843 (N_49843,N_35404,N_34434);
xor U49844 (N_49844,N_32151,N_33025);
xnor U49845 (N_49845,N_31521,N_39954);
xnor U49846 (N_49846,N_37777,N_37480);
nor U49847 (N_49847,N_37596,N_38996);
and U49848 (N_49848,N_36048,N_37478);
or U49849 (N_49849,N_31771,N_30267);
or U49850 (N_49850,N_32805,N_38317);
and U49851 (N_49851,N_33545,N_34580);
or U49852 (N_49852,N_34973,N_35573);
xnor U49853 (N_49853,N_32648,N_37891);
nor U49854 (N_49854,N_39772,N_38560);
xnor U49855 (N_49855,N_34576,N_38600);
and U49856 (N_49856,N_39215,N_34821);
and U49857 (N_49857,N_34334,N_36031);
xnor U49858 (N_49858,N_37091,N_32936);
nand U49859 (N_49859,N_38254,N_36335);
xor U49860 (N_49860,N_30321,N_39691);
xor U49861 (N_49861,N_31771,N_34542);
nor U49862 (N_49862,N_34643,N_38967);
and U49863 (N_49863,N_34632,N_30600);
nor U49864 (N_49864,N_34538,N_31835);
xor U49865 (N_49865,N_32967,N_38354);
nand U49866 (N_49866,N_38384,N_38171);
nand U49867 (N_49867,N_30931,N_31070);
or U49868 (N_49868,N_30445,N_33524);
xor U49869 (N_49869,N_35240,N_35126);
and U49870 (N_49870,N_31948,N_32526);
xor U49871 (N_49871,N_39634,N_39224);
and U49872 (N_49872,N_38336,N_34180);
nor U49873 (N_49873,N_30207,N_32262);
nand U49874 (N_49874,N_30944,N_33971);
nand U49875 (N_49875,N_38245,N_34206);
nand U49876 (N_49876,N_32587,N_35536);
nor U49877 (N_49877,N_30372,N_38456);
nor U49878 (N_49878,N_39596,N_33839);
nor U49879 (N_49879,N_36150,N_33008);
or U49880 (N_49880,N_39627,N_36340);
or U49881 (N_49881,N_30324,N_35744);
or U49882 (N_49882,N_32356,N_32272);
or U49883 (N_49883,N_34044,N_39327);
or U49884 (N_49884,N_36195,N_37508);
or U49885 (N_49885,N_35737,N_30471);
and U49886 (N_49886,N_35401,N_34176);
and U49887 (N_49887,N_34172,N_35940);
nand U49888 (N_49888,N_30862,N_36910);
nand U49889 (N_49889,N_34032,N_35236);
and U49890 (N_49890,N_39813,N_32873);
nor U49891 (N_49891,N_38949,N_38776);
xor U49892 (N_49892,N_30155,N_36222);
or U49893 (N_49893,N_37215,N_34080);
or U49894 (N_49894,N_33300,N_38861);
or U49895 (N_49895,N_34118,N_33480);
nand U49896 (N_49896,N_39538,N_30923);
or U49897 (N_49897,N_32784,N_34506);
xnor U49898 (N_49898,N_39645,N_31084);
nand U49899 (N_49899,N_31577,N_38536);
xor U49900 (N_49900,N_34480,N_31923);
nor U49901 (N_49901,N_30007,N_34499);
nor U49902 (N_49902,N_34010,N_31892);
or U49903 (N_49903,N_34991,N_32617);
xnor U49904 (N_49904,N_37813,N_33745);
or U49905 (N_49905,N_34372,N_39262);
or U49906 (N_49906,N_33765,N_33708);
and U49907 (N_49907,N_36397,N_37809);
or U49908 (N_49908,N_31332,N_30187);
xnor U49909 (N_49909,N_39465,N_38496);
nand U49910 (N_49910,N_34252,N_32939);
xor U49911 (N_49911,N_33924,N_31604);
nand U49912 (N_49912,N_30784,N_30936);
and U49913 (N_49913,N_31297,N_38150);
xnor U49914 (N_49914,N_32392,N_32277);
nand U49915 (N_49915,N_37651,N_37789);
or U49916 (N_49916,N_31217,N_38130);
and U49917 (N_49917,N_33527,N_38322);
nor U49918 (N_49918,N_33329,N_30207);
and U49919 (N_49919,N_37484,N_32868);
nor U49920 (N_49920,N_38449,N_30646);
or U49921 (N_49921,N_32268,N_38453);
xnor U49922 (N_49922,N_38963,N_33274);
and U49923 (N_49923,N_33141,N_32194);
or U49924 (N_49924,N_39306,N_39245);
and U49925 (N_49925,N_34165,N_35753);
nand U49926 (N_49926,N_37626,N_31351);
or U49927 (N_49927,N_30256,N_31676);
or U49928 (N_49928,N_37347,N_39896);
nand U49929 (N_49929,N_36747,N_30002);
and U49930 (N_49930,N_35586,N_35133);
xnor U49931 (N_49931,N_30873,N_31612);
nand U49932 (N_49932,N_33547,N_33340);
and U49933 (N_49933,N_36570,N_37435);
nand U49934 (N_49934,N_34869,N_30553);
and U49935 (N_49935,N_34786,N_39382);
and U49936 (N_49936,N_35806,N_30824);
nand U49937 (N_49937,N_37274,N_31377);
nand U49938 (N_49938,N_38393,N_36674);
xnor U49939 (N_49939,N_36290,N_30324);
nor U49940 (N_49940,N_39788,N_38745);
or U49941 (N_49941,N_35219,N_33522);
nor U49942 (N_49942,N_30400,N_33303);
xnor U49943 (N_49943,N_35109,N_39355);
or U49944 (N_49944,N_31299,N_39177);
nand U49945 (N_49945,N_39737,N_37823);
nand U49946 (N_49946,N_34908,N_31223);
and U49947 (N_49947,N_39444,N_34855);
nand U49948 (N_49948,N_35305,N_34027);
xor U49949 (N_49949,N_32221,N_39931);
nor U49950 (N_49950,N_34466,N_30586);
nand U49951 (N_49951,N_37590,N_34517);
and U49952 (N_49952,N_35078,N_35617);
and U49953 (N_49953,N_32317,N_36644);
and U49954 (N_49954,N_38618,N_36457);
nand U49955 (N_49955,N_37331,N_38633);
nand U49956 (N_49956,N_32471,N_33961);
or U49957 (N_49957,N_39942,N_39751);
nand U49958 (N_49958,N_35994,N_37902);
and U49959 (N_49959,N_34269,N_33563);
xor U49960 (N_49960,N_37257,N_35731);
and U49961 (N_49961,N_34978,N_31961);
and U49962 (N_49962,N_32085,N_38412);
xnor U49963 (N_49963,N_38214,N_34494);
xnor U49964 (N_49964,N_34967,N_35308);
and U49965 (N_49965,N_38597,N_31752);
and U49966 (N_49966,N_34790,N_30183);
xnor U49967 (N_49967,N_38757,N_39347);
nand U49968 (N_49968,N_33466,N_36132);
xor U49969 (N_49969,N_32009,N_32163);
and U49970 (N_49970,N_30369,N_38903);
nor U49971 (N_49971,N_31662,N_38426);
or U49972 (N_49972,N_31257,N_39450);
xnor U49973 (N_49973,N_36097,N_36760);
or U49974 (N_49974,N_31467,N_33683);
nand U49975 (N_49975,N_38755,N_35936);
and U49976 (N_49976,N_36675,N_33255);
xnor U49977 (N_49977,N_39944,N_35718);
and U49978 (N_49978,N_38311,N_38363);
nand U49979 (N_49979,N_33007,N_32649);
nand U49980 (N_49980,N_34768,N_30394);
nand U49981 (N_49981,N_36989,N_37008);
xnor U49982 (N_49982,N_30265,N_34004);
or U49983 (N_49983,N_30745,N_35086);
nor U49984 (N_49984,N_39053,N_36530);
nand U49985 (N_49985,N_31194,N_37362);
nand U49986 (N_49986,N_31269,N_39920);
xnor U49987 (N_49987,N_34159,N_35762);
xor U49988 (N_49988,N_35329,N_33877);
or U49989 (N_49989,N_34812,N_34121);
nand U49990 (N_49990,N_32585,N_30087);
xor U49991 (N_49991,N_38256,N_32335);
nor U49992 (N_49992,N_35494,N_36496);
xnor U49993 (N_49993,N_30064,N_38582);
nor U49994 (N_49994,N_34359,N_35632);
nor U49995 (N_49995,N_36992,N_35459);
and U49996 (N_49996,N_34410,N_35119);
and U49997 (N_49997,N_32288,N_35394);
or U49998 (N_49998,N_39818,N_36727);
and U49999 (N_49999,N_30635,N_31749);
xnor UO_0 (O_0,N_45628,N_45506);
and UO_1 (O_1,N_45781,N_44712);
and UO_2 (O_2,N_48664,N_45923);
and UO_3 (O_3,N_45022,N_42031);
nand UO_4 (O_4,N_48871,N_46804);
and UO_5 (O_5,N_47203,N_40168);
nor UO_6 (O_6,N_49381,N_42152);
xor UO_7 (O_7,N_48600,N_40493);
nor UO_8 (O_8,N_42801,N_49211);
xnor UO_9 (O_9,N_48288,N_44625);
and UO_10 (O_10,N_40021,N_45046);
nor UO_11 (O_11,N_44582,N_41647);
xor UO_12 (O_12,N_43890,N_42915);
or UO_13 (O_13,N_46287,N_41469);
nand UO_14 (O_14,N_49926,N_49475);
or UO_15 (O_15,N_49580,N_40056);
xor UO_16 (O_16,N_44982,N_40861);
nor UO_17 (O_17,N_45836,N_40625);
nor UO_18 (O_18,N_45513,N_40496);
nand UO_19 (O_19,N_43907,N_41687);
or UO_20 (O_20,N_46256,N_45716);
or UO_21 (O_21,N_43814,N_42631);
and UO_22 (O_22,N_43322,N_44150);
or UO_23 (O_23,N_44770,N_47905);
nor UO_24 (O_24,N_49500,N_43952);
and UO_25 (O_25,N_41220,N_46971);
and UO_26 (O_26,N_41553,N_42448);
or UO_27 (O_27,N_46389,N_47875);
xor UO_28 (O_28,N_48864,N_47748);
or UO_29 (O_29,N_43235,N_41391);
nor UO_30 (O_30,N_40362,N_49966);
or UO_31 (O_31,N_47708,N_45977);
xnor UO_32 (O_32,N_43465,N_42617);
or UO_33 (O_33,N_46867,N_49621);
nor UO_34 (O_34,N_40212,N_44321);
xor UO_35 (O_35,N_42501,N_47328);
nand UO_36 (O_36,N_40446,N_49662);
nand UO_37 (O_37,N_48742,N_48477);
and UO_38 (O_38,N_45003,N_48370);
nand UO_39 (O_39,N_48439,N_42870);
and UO_40 (O_40,N_48497,N_42889);
and UO_41 (O_41,N_45015,N_45712);
or UO_42 (O_42,N_45432,N_40980);
nand UO_43 (O_43,N_45135,N_48475);
nor UO_44 (O_44,N_43534,N_49736);
nor UO_45 (O_45,N_42083,N_48251);
or UO_46 (O_46,N_47744,N_46460);
nor UO_47 (O_47,N_40876,N_48471);
xor UO_48 (O_48,N_41385,N_49937);
nor UO_49 (O_49,N_40550,N_45839);
xor UO_50 (O_50,N_42541,N_41656);
xnor UO_51 (O_51,N_43216,N_45793);
nand UO_52 (O_52,N_42565,N_40488);
xnor UO_53 (O_53,N_44659,N_48143);
or UO_54 (O_54,N_43318,N_40816);
nor UO_55 (O_55,N_47428,N_45855);
or UO_56 (O_56,N_41923,N_48934);
nor UO_57 (O_57,N_47721,N_44389);
or UO_58 (O_58,N_48713,N_45649);
nor UO_59 (O_59,N_44640,N_43272);
nor UO_60 (O_60,N_48955,N_46757);
nor UO_61 (O_61,N_42757,N_47626);
xnor UO_62 (O_62,N_46887,N_43419);
nand UO_63 (O_63,N_41456,N_41154);
nand UO_64 (O_64,N_40755,N_40400);
nor UO_65 (O_65,N_41188,N_46444);
and UO_66 (O_66,N_49668,N_45311);
and UO_67 (O_67,N_44945,N_40581);
nor UO_68 (O_68,N_49839,N_44858);
and UO_69 (O_69,N_46664,N_48583);
or UO_70 (O_70,N_41077,N_45884);
and UO_71 (O_71,N_46266,N_47851);
and UO_72 (O_72,N_43374,N_49469);
xor UO_73 (O_73,N_41216,N_46479);
nor UO_74 (O_74,N_43683,N_43881);
and UO_75 (O_75,N_40354,N_47491);
or UO_76 (O_76,N_40392,N_42937);
and UO_77 (O_77,N_40316,N_46409);
nor UO_78 (O_78,N_42894,N_45479);
nor UO_79 (O_79,N_49782,N_49635);
or UO_80 (O_80,N_42092,N_47877);
xor UO_81 (O_81,N_41831,N_43191);
nand UO_82 (O_82,N_45965,N_45430);
and UO_83 (O_83,N_44957,N_48855);
and UO_84 (O_84,N_41938,N_40420);
and UO_85 (O_85,N_49436,N_41406);
xnor UO_86 (O_86,N_44428,N_49395);
and UO_87 (O_87,N_48595,N_42508);
xnor UO_88 (O_88,N_42093,N_42466);
and UO_89 (O_89,N_46611,N_46120);
nor UO_90 (O_90,N_40835,N_40210);
nor UO_91 (O_91,N_44748,N_49717);
or UO_92 (O_92,N_49905,N_40030);
xnor UO_93 (O_93,N_40782,N_43623);
or UO_94 (O_94,N_45767,N_42648);
and UO_95 (O_95,N_40925,N_45984);
nor UO_96 (O_96,N_47754,N_44280);
and UO_97 (O_97,N_49341,N_48052);
and UO_98 (O_98,N_46206,N_42884);
and UO_99 (O_99,N_46468,N_40343);
xnor UO_100 (O_100,N_40186,N_49578);
nand UO_101 (O_101,N_43455,N_47294);
and UO_102 (O_102,N_44112,N_41820);
xnor UO_103 (O_103,N_42759,N_42951);
xor UO_104 (O_104,N_43369,N_46902);
nand UO_105 (O_105,N_46638,N_49311);
and UO_106 (O_106,N_42040,N_43726);
and UO_107 (O_107,N_46602,N_44794);
nor UO_108 (O_108,N_42552,N_47479);
nor UO_109 (O_109,N_44898,N_48619);
or UO_110 (O_110,N_40218,N_44981);
and UO_111 (O_111,N_49128,N_42649);
and UO_112 (O_112,N_45285,N_49622);
xor UO_113 (O_113,N_49454,N_40465);
xor UO_114 (O_114,N_42816,N_47122);
and UO_115 (O_115,N_41185,N_48392);
and UO_116 (O_116,N_43287,N_40929);
or UO_117 (O_117,N_49760,N_47917);
nor UO_118 (O_118,N_45252,N_40649);
xnor UO_119 (O_119,N_42133,N_46192);
xnor UO_120 (O_120,N_41743,N_46617);
or UO_121 (O_121,N_40371,N_43067);
xnor UO_122 (O_122,N_45010,N_41764);
or UO_123 (O_123,N_49490,N_44587);
and UO_124 (O_124,N_44535,N_44578);
xor UO_125 (O_125,N_49989,N_45248);
xor UO_126 (O_126,N_43462,N_46306);
nand UO_127 (O_127,N_49809,N_45589);
nor UO_128 (O_128,N_41410,N_47272);
nand UO_129 (O_129,N_48333,N_40197);
and UO_130 (O_130,N_41095,N_40386);
and UO_131 (O_131,N_49555,N_48078);
and UO_132 (O_132,N_40374,N_41380);
and UO_133 (O_133,N_44278,N_46429);
nor UO_134 (O_134,N_40334,N_47677);
nand UO_135 (O_135,N_47679,N_42997);
xnor UO_136 (O_136,N_47610,N_47115);
xor UO_137 (O_137,N_45104,N_48823);
or UO_138 (O_138,N_46368,N_42583);
nand UO_139 (O_139,N_45811,N_47181);
xor UO_140 (O_140,N_48993,N_44384);
or UO_141 (O_141,N_42630,N_48950);
nor UO_142 (O_142,N_44990,N_41986);
nand UO_143 (O_143,N_48838,N_40448);
nor UO_144 (O_144,N_44061,N_46693);
xor UO_145 (O_145,N_42783,N_49978);
nand UO_146 (O_146,N_41419,N_47755);
or UO_147 (O_147,N_45857,N_48045);
nand UO_148 (O_148,N_42166,N_40079);
and UO_149 (O_149,N_44148,N_40127);
xnor UO_150 (O_150,N_46519,N_44049);
xnor UO_151 (O_151,N_47629,N_47436);
xnor UO_152 (O_152,N_40416,N_41326);
and UO_153 (O_153,N_41783,N_43756);
or UO_154 (O_154,N_49990,N_48830);
and UO_155 (O_155,N_46772,N_47298);
and UO_156 (O_156,N_41407,N_43069);
or UO_157 (O_157,N_47553,N_48640);
xor UO_158 (O_158,N_49568,N_40007);
xor UO_159 (O_159,N_44452,N_40434);
xor UO_160 (O_160,N_45256,N_49970);
xnor UO_161 (O_161,N_42538,N_46874);
nor UO_162 (O_162,N_45308,N_42850);
or UO_163 (O_163,N_44129,N_46196);
or UO_164 (O_164,N_44759,N_46024);
xnor UO_165 (O_165,N_45455,N_40287);
xnor UO_166 (O_166,N_41784,N_49107);
nand UO_167 (O_167,N_43492,N_43178);
and UO_168 (O_168,N_47526,N_46722);
xnor UO_169 (O_169,N_48484,N_49841);
xnor UO_170 (O_170,N_47440,N_49589);
nand UO_171 (O_171,N_43509,N_46639);
nand UO_172 (O_172,N_47676,N_46286);
or UO_173 (O_173,N_46093,N_40779);
xor UO_174 (O_174,N_45909,N_42690);
nand UO_175 (O_175,N_40621,N_44971);
nor UO_176 (O_176,N_42163,N_49875);
or UO_177 (O_177,N_46130,N_47042);
nand UO_178 (O_178,N_43280,N_44414);
nor UO_179 (O_179,N_40813,N_44015);
nor UO_180 (O_180,N_46158,N_43147);
xnor UO_181 (O_181,N_44160,N_47004);
xor UO_182 (O_182,N_46386,N_40901);
nand UO_183 (O_183,N_43669,N_46812);
nand UO_184 (O_184,N_49288,N_43131);
nand UO_185 (O_185,N_40028,N_48554);
nand UO_186 (O_186,N_41473,N_46305);
and UO_187 (O_187,N_43561,N_47194);
nand UO_188 (O_188,N_49797,N_43415);
or UO_189 (O_189,N_48271,N_48083);
or UO_190 (O_190,N_40988,N_41853);
nand UO_191 (O_191,N_46347,N_41817);
xnor UO_192 (O_192,N_44098,N_48712);
or UO_193 (O_193,N_48418,N_47078);
or UO_194 (O_194,N_44687,N_42881);
or UO_195 (O_195,N_45822,N_46498);
and UO_196 (O_196,N_44008,N_46543);
xnor UO_197 (O_197,N_44092,N_47333);
and UO_198 (O_198,N_49856,N_40768);
and UO_199 (O_199,N_47840,N_42475);
xor UO_200 (O_200,N_43803,N_42480);
and UO_201 (O_201,N_44437,N_43478);
nor UO_202 (O_202,N_44466,N_45730);
nand UO_203 (O_203,N_42286,N_49237);
xor UO_204 (O_204,N_46587,N_49804);
xnor UO_205 (O_205,N_45496,N_47397);
nand UO_206 (O_206,N_43159,N_44871);
nor UO_207 (O_207,N_47992,N_47098);
or UO_208 (O_208,N_44525,N_48531);
xnor UO_209 (O_209,N_44863,N_40575);
nor UO_210 (O_210,N_41600,N_44139);
or UO_211 (O_211,N_41157,N_41305);
nor UO_212 (O_212,N_46048,N_40244);
nand UO_213 (O_213,N_46210,N_43372);
xnor UO_214 (O_214,N_46145,N_40892);
nor UO_215 (O_215,N_40987,N_40899);
or UO_216 (O_216,N_40827,N_44506);
or UO_217 (O_217,N_41014,N_48468);
xnor UO_218 (O_218,N_45366,N_44809);
nand UO_219 (O_219,N_41362,N_48327);
or UO_220 (O_220,N_47522,N_44311);
nand UO_221 (O_221,N_43793,N_40013);
or UO_222 (O_222,N_43924,N_46432);
xnor UO_223 (O_223,N_42684,N_46885);
nand UO_224 (O_224,N_48691,N_44545);
or UO_225 (O_225,N_49719,N_44084);
or UO_226 (O_226,N_45111,N_43826);
nand UO_227 (O_227,N_44928,N_47608);
nor UO_228 (O_228,N_44433,N_41508);
nand UO_229 (O_229,N_40658,N_42703);
xor UO_230 (O_230,N_40541,N_47923);
and UO_231 (O_231,N_43698,N_40499);
or UO_232 (O_232,N_42640,N_48079);
nand UO_233 (O_233,N_43718,N_41863);
nand UO_234 (O_234,N_49504,N_41822);
xor UO_235 (O_235,N_48215,N_40754);
nand UO_236 (O_236,N_48164,N_46978);
nand UO_237 (O_237,N_44108,N_42071);
xor UO_238 (O_238,N_44217,N_49376);
xnor UO_239 (O_239,N_49427,N_44403);
xnor UO_240 (O_240,N_49921,N_45808);
nor UO_241 (O_241,N_44592,N_46556);
and UO_242 (O_242,N_46068,N_48951);
xnor UO_243 (O_243,N_44810,N_44169);
and UO_244 (O_244,N_40549,N_45665);
or UO_245 (O_245,N_41937,N_45530);
nand UO_246 (O_246,N_48416,N_49125);
nand UO_247 (O_247,N_42377,N_45096);
or UO_248 (O_248,N_49429,N_47276);
nand UO_249 (O_249,N_45355,N_44542);
nor UO_250 (O_250,N_41983,N_49209);
nor UO_251 (O_251,N_47046,N_44869);
and UO_252 (O_252,N_47577,N_46066);
xor UO_253 (O_253,N_43784,N_45615);
nand UO_254 (O_254,N_48239,N_43036);
nor UO_255 (O_255,N_41205,N_44132);
or UO_256 (O_256,N_45208,N_46296);
nor UO_257 (O_257,N_46064,N_41344);
xor UO_258 (O_258,N_47396,N_44505);
or UO_259 (O_259,N_46582,N_44448);
xor UO_260 (O_260,N_47492,N_41311);
and UO_261 (O_261,N_47344,N_43151);
and UO_262 (O_262,N_41346,N_41012);
and UO_263 (O_263,N_44864,N_49379);
xor UO_264 (O_264,N_41262,N_42109);
and UO_265 (O_265,N_47467,N_48962);
xnor UO_266 (O_266,N_46688,N_45017);
xnor UO_267 (O_267,N_41067,N_49026);
or UO_268 (O_268,N_47883,N_40093);
nor UO_269 (O_269,N_41858,N_44091);
nor UO_270 (O_270,N_45931,N_49561);
nand UO_271 (O_271,N_45429,N_41897);
nor UO_272 (O_272,N_41792,N_40332);
nand UO_273 (O_273,N_45287,N_47488);
and UO_274 (O_274,N_47569,N_47798);
xnor UO_275 (O_275,N_48602,N_42808);
xnor UO_276 (O_276,N_44744,N_41234);
and UO_277 (O_277,N_47480,N_43730);
xnor UO_278 (O_278,N_44096,N_43734);
nand UO_279 (O_279,N_49949,N_48882);
nand UO_280 (O_280,N_42341,N_47293);
xor UO_281 (O_281,N_40729,N_40762);
xnor UO_282 (O_282,N_48103,N_46061);
or UO_283 (O_283,N_48588,N_47030);
or UO_284 (O_284,N_46336,N_40613);
xnor UO_285 (O_285,N_47937,N_46790);
xnor UO_286 (O_286,N_49864,N_44265);
nand UO_287 (O_287,N_40132,N_46233);
xor UO_288 (O_288,N_46739,N_42202);
nand UO_289 (O_289,N_40545,N_44698);
xor UO_290 (O_290,N_42683,N_42800);
nand UO_291 (O_291,N_49629,N_45200);
and UO_292 (O_292,N_47505,N_40863);
or UO_293 (O_293,N_43312,N_41423);
nor UO_294 (O_294,N_44165,N_40269);
nor UO_295 (O_295,N_42278,N_41935);
or UO_296 (O_296,N_49424,N_42151);
nand UO_297 (O_297,N_45748,N_49838);
nor UO_298 (O_298,N_45858,N_46465);
and UO_299 (O_299,N_43172,N_46888);
or UO_300 (O_300,N_46480,N_48750);
or UO_301 (O_301,N_46509,N_44290);
or UO_302 (O_302,N_47906,N_47006);
nand UO_303 (O_303,N_40483,N_44675);
xor UO_304 (O_304,N_43763,N_43457);
and UO_305 (O_305,N_43023,N_48262);
nand UO_306 (O_306,N_44873,N_49616);
and UO_307 (O_307,N_45026,N_44881);
nand UO_308 (O_308,N_46754,N_41644);
xor UO_309 (O_309,N_40089,N_43508);
or UO_310 (O_310,N_45130,N_44848);
and UO_311 (O_311,N_46928,N_41733);
nand UO_312 (O_312,N_42191,N_49811);
nor UO_313 (O_313,N_47297,N_49503);
nor UO_314 (O_314,N_44522,N_44313);
or UO_315 (O_315,N_43746,N_46092);
nand UO_316 (O_316,N_44146,N_42476);
and UO_317 (O_317,N_48532,N_41487);
or UO_318 (O_318,N_42198,N_41231);
or UO_319 (O_319,N_49312,N_44082);
xor UO_320 (O_320,N_42619,N_48144);
nand UO_321 (O_321,N_41823,N_42966);
nand UO_322 (O_322,N_45899,N_40644);
nand UO_323 (O_323,N_48862,N_46099);
xor UO_324 (O_324,N_41363,N_47562);
nor UO_325 (O_325,N_47730,N_40681);
nor UO_326 (O_326,N_49860,N_47172);
nor UO_327 (O_327,N_41283,N_47392);
nor UO_328 (O_328,N_44793,N_48833);
and UO_329 (O_329,N_47874,N_43264);
nand UO_330 (O_330,N_43776,N_46027);
nand UO_331 (O_331,N_44067,N_42730);
nor UO_332 (O_332,N_40588,N_49681);
or UO_333 (O_333,N_40839,N_47360);
nor UO_334 (O_334,N_45450,N_49508);
or UO_335 (O_335,N_47274,N_42946);
or UO_336 (O_336,N_43005,N_47349);
or UO_337 (O_337,N_43240,N_48959);
and UO_338 (O_338,N_47558,N_43072);
nand UO_339 (O_339,N_41123,N_40232);
and UO_340 (O_340,N_42605,N_40195);
and UO_341 (O_341,N_44654,N_45750);
nor UO_342 (O_342,N_49098,N_41511);
xor UO_343 (O_343,N_49847,N_41444);
nand UO_344 (O_344,N_45655,N_43161);
or UO_345 (O_345,N_47997,N_46669);
nor UO_346 (O_346,N_46244,N_41752);
and UO_347 (O_347,N_47289,N_47720);
or UO_348 (O_348,N_43435,N_41393);
or UO_349 (O_349,N_49346,N_46065);
and UO_350 (O_350,N_48305,N_40450);
nand UO_351 (O_351,N_46416,N_45663);
and UO_352 (O_352,N_49979,N_40801);
xnor UO_353 (O_353,N_48992,N_48301);
nor UO_354 (O_354,N_44738,N_44603);
or UO_355 (O_355,N_41513,N_45986);
nor UO_356 (O_356,N_41786,N_44016);
nor UO_357 (O_357,N_41850,N_49333);
nor UO_358 (O_358,N_46270,N_45196);
nand UO_359 (O_359,N_47408,N_47785);
or UO_360 (O_360,N_48979,N_45277);
nor UO_361 (O_361,N_42204,N_44152);
xnor UO_362 (O_362,N_45861,N_40272);
nand UO_363 (O_363,N_47654,N_48201);
xor UO_364 (O_364,N_41144,N_46457);
nand UO_365 (O_365,N_46743,N_44376);
xor UO_366 (O_366,N_43150,N_41379);
or UO_367 (O_367,N_49851,N_49798);
or UO_368 (O_368,N_49673,N_47576);
or UO_369 (O_369,N_49925,N_44649);
and UO_370 (O_370,N_45772,N_45136);
xnor UO_371 (O_371,N_47804,N_47597);
xor UO_372 (O_372,N_49417,N_46863);
nor UO_373 (O_373,N_46545,N_49924);
and UO_374 (O_374,N_47326,N_44259);
xor UO_375 (O_375,N_44474,N_42797);
xnor UO_376 (O_376,N_47793,N_42055);
nand UO_377 (O_377,N_46697,N_40080);
or UO_378 (O_378,N_47153,N_46692);
and UO_379 (O_379,N_47083,N_46417);
nor UO_380 (O_380,N_43311,N_42081);
xnor UO_381 (O_381,N_44285,N_42811);
nor UO_382 (O_382,N_49126,N_41491);
nor UO_383 (O_383,N_40590,N_46317);
nor UO_384 (O_384,N_48798,N_40856);
nor UO_385 (O_385,N_49339,N_40534);
nand UO_386 (O_386,N_47617,N_48429);
nand UO_387 (O_387,N_43886,N_43001);
xor UO_388 (O_388,N_42749,N_42639);
and UO_389 (O_389,N_41055,N_46658);
nor UO_390 (O_390,N_45850,N_46226);
or UO_391 (O_391,N_46109,N_40918);
xor UO_392 (O_392,N_42642,N_45033);
xor UO_393 (O_393,N_46010,N_47635);
nor UO_394 (O_394,N_49695,N_47896);
or UO_395 (O_395,N_45073,N_49940);
nor UO_396 (O_396,N_43047,N_42100);
or UO_397 (O_397,N_41825,N_49920);
nand UO_398 (O_398,N_47501,N_42036);
xnor UO_399 (O_399,N_41399,N_44880);
and UO_400 (O_400,N_43286,N_40971);
xnor UO_401 (O_401,N_41452,N_42943);
xor UO_402 (O_402,N_49972,N_47530);
nor UO_403 (O_403,N_46079,N_47380);
nor UO_404 (O_404,N_45658,N_44622);
nor UO_405 (O_405,N_41663,N_49711);
and UO_406 (O_406,N_46393,N_48469);
xnor UO_407 (O_407,N_41778,N_49184);
xor UO_408 (O_408,N_45693,N_46659);
nand UO_409 (O_409,N_45675,N_45148);
and UO_410 (O_410,N_41099,N_41299);
nand UO_411 (O_411,N_41713,N_49388);
xor UO_412 (O_412,N_45947,N_45946);
nor UO_413 (O_413,N_43461,N_41125);
or UO_414 (O_414,N_46440,N_47671);
xor UO_415 (O_415,N_40740,N_48749);
and UO_416 (O_416,N_47656,N_45768);
or UO_417 (O_417,N_49603,N_47070);
or UO_418 (O_418,N_46958,N_42868);
nand UO_419 (O_419,N_41912,N_40006);
nor UO_420 (O_420,N_46359,N_48267);
xor UO_421 (O_421,N_43368,N_40043);
and UO_422 (O_422,N_42579,N_46940);
nor UO_423 (O_423,N_43733,N_40363);
nand UO_424 (O_424,N_41948,N_41576);
nand UO_425 (O_425,N_48641,N_44019);
xnor UO_426 (O_426,N_40598,N_41498);
or UO_427 (O_427,N_42836,N_48275);
xnor UO_428 (O_428,N_47513,N_46459);
nand UO_429 (O_429,N_40470,N_40910);
xnor UO_430 (O_430,N_48024,N_46579);
nand UO_431 (O_431,N_40207,N_47000);
nand UO_432 (O_432,N_49428,N_45000);
nand UO_433 (O_433,N_45162,N_42398);
nor UO_434 (O_434,N_48104,N_46161);
nand UO_435 (O_435,N_40340,N_49242);
nor UO_436 (O_436,N_48897,N_40278);
nor UO_437 (O_437,N_41943,N_48286);
nor UO_438 (O_438,N_46211,N_47702);
xnor UO_439 (O_439,N_48702,N_44127);
and UO_440 (O_440,N_43453,N_41076);
nand UO_441 (O_441,N_44661,N_47077);
or UO_442 (O_442,N_48382,N_46728);
xor UO_443 (O_443,N_43610,N_48661);
and UO_444 (O_444,N_44270,N_43602);
or UO_445 (O_445,N_40140,N_47481);
xnor UO_446 (O_446,N_40557,N_45805);
or UO_447 (O_447,N_45543,N_44012);
and UO_448 (O_448,N_44037,N_40643);
nor UO_449 (O_449,N_47761,N_48085);
xor UO_450 (O_450,N_45701,N_44696);
xor UO_451 (O_451,N_40002,N_49173);
or UO_452 (O_452,N_47709,N_44151);
nand UO_453 (O_453,N_47788,N_45217);
or UO_454 (O_454,N_45131,N_41910);
nor UO_455 (O_455,N_44876,N_45336);
and UO_456 (O_456,N_40855,N_49667);
nand UO_457 (O_457,N_42962,N_44763);
nor UO_458 (O_458,N_40066,N_49626);
nand UO_459 (O_459,N_45207,N_48081);
nand UO_460 (O_460,N_40605,N_40133);
nor UO_461 (O_461,N_44318,N_40769);
and UO_462 (O_462,N_48246,N_46000);
nand UO_463 (O_463,N_45960,N_45956);
nor UO_464 (O_464,N_46029,N_46522);
nor UO_465 (O_465,N_45254,N_47706);
nor UO_466 (O_466,N_46581,N_46787);
and UO_467 (O_467,N_45614,N_41832);
and UO_468 (O_468,N_42600,N_43749);
xor UO_469 (O_469,N_42548,N_42130);
xnor UO_470 (O_470,N_42450,N_46549);
or UO_471 (O_471,N_40919,N_46926);
and UO_472 (O_472,N_49577,N_43234);
and UO_473 (O_473,N_45827,N_46148);
or UO_474 (O_474,N_45508,N_41502);
nand UO_475 (O_475,N_44296,N_42387);
xnor UO_476 (O_476,N_41848,N_42587);
nand UO_477 (O_477,N_49282,N_42078);
xor UO_478 (O_478,N_42473,N_41213);
nor UO_479 (O_479,N_47192,N_46920);
or UO_480 (O_480,N_40923,N_43402);
nor UO_481 (O_481,N_42142,N_43083);
nor UO_482 (O_482,N_41602,N_48582);
or UO_483 (O_483,N_42149,N_45690);
or UO_484 (O_484,N_41988,N_40686);
nand UO_485 (O_485,N_45145,N_47154);
nor UO_486 (O_486,N_48840,N_40521);
nor UO_487 (O_487,N_47589,N_46195);
xor UO_488 (O_488,N_43898,N_43688);
nand UO_489 (O_489,N_42070,N_49732);
nor UO_490 (O_490,N_48389,N_46532);
nor UO_491 (O_491,N_46486,N_48774);
xnor UO_492 (O_492,N_41302,N_41535);
xnor UO_493 (O_493,N_46102,N_45498);
and UO_494 (O_494,N_40129,N_49048);
nand UO_495 (O_495,N_49448,N_49235);
nor UO_496 (O_496,N_45422,N_44657);
xnor UO_497 (O_497,N_46770,N_49111);
or UO_498 (O_498,N_47002,N_42610);
nor UO_499 (O_499,N_49714,N_43471);
or UO_500 (O_500,N_41306,N_42712);
nand UO_501 (O_501,N_47956,N_48023);
xnor UO_502 (O_502,N_46308,N_48254);
nand UO_503 (O_503,N_49687,N_43021);
nand UO_504 (O_504,N_46964,N_43401);
or UO_505 (O_505,N_40949,N_45698);
xor UO_506 (O_506,N_48891,N_40103);
and UO_507 (O_507,N_41135,N_49205);
or UO_508 (O_508,N_45672,N_49226);
xor UO_509 (O_509,N_40837,N_45290);
xor UO_510 (O_510,N_41160,N_41737);
nand UO_511 (O_511,N_48378,N_43042);
nor UO_512 (O_512,N_46261,N_44606);
and UO_513 (O_513,N_40073,N_45079);
nor UO_514 (O_514,N_41013,N_46974);
nand UO_515 (O_515,N_42644,N_49815);
nand UO_516 (O_516,N_44394,N_43873);
xor UO_517 (O_517,N_49538,N_45623);
and UO_518 (O_518,N_49823,N_42832);
or UO_519 (O_519,N_48690,N_43175);
or UO_520 (O_520,N_40208,N_45798);
and UO_521 (O_521,N_46820,N_46028);
and UO_522 (O_522,N_42073,N_48295);
nor UO_523 (O_523,N_48888,N_42023);
nand UO_524 (O_524,N_49514,N_44253);
nand UO_525 (O_525,N_40883,N_41307);
and UO_526 (O_526,N_44523,N_41340);
nor UO_527 (O_527,N_41691,N_42063);
or UO_528 (O_528,N_49192,N_40459);
nand UO_529 (O_529,N_49214,N_41484);
nor UO_530 (O_530,N_46025,N_40457);
or UO_531 (O_531,N_45892,N_49170);
nand UO_532 (O_532,N_46205,N_49742);
nand UO_533 (O_533,N_43527,N_44663);
nand UO_534 (O_534,N_41319,N_42465);
or UO_535 (O_535,N_41547,N_46273);
xor UO_536 (O_536,N_43041,N_48542);
or UO_537 (O_537,N_42233,N_41247);
nor UO_538 (O_538,N_49982,N_42782);
xor UO_539 (O_539,N_42028,N_44776);
nand UO_540 (O_540,N_40906,N_41207);
nor UO_541 (O_541,N_41128,N_46574);
and UO_542 (O_542,N_44136,N_49273);
or UO_543 (O_543,N_48000,N_40756);
xor UO_544 (O_544,N_41303,N_40728);
nand UO_545 (O_545,N_40027,N_41392);
xnor UO_546 (O_546,N_44121,N_43104);
nor UO_547 (O_547,N_42510,N_42741);
and UO_548 (O_548,N_47945,N_48125);
xnor UO_549 (O_549,N_46765,N_49343);
nand UO_550 (O_550,N_47039,N_43289);
nand UO_551 (O_551,N_49482,N_47095);
nand UO_552 (O_552,N_42150,N_48571);
and UO_553 (O_553,N_43671,N_46184);
or UO_554 (O_554,N_49656,N_41945);
nor UO_555 (O_555,N_49426,N_41738);
or UO_556 (O_556,N_42732,N_41523);
nand UO_557 (O_557,N_46809,N_46246);
nand UO_558 (O_558,N_48629,N_47867);
or UO_559 (O_559,N_42696,N_49552);
nand UO_560 (O_560,N_41023,N_44652);
or UO_561 (O_561,N_42311,N_47285);
nor UO_562 (O_562,N_42553,N_46796);
and UO_563 (O_563,N_48425,N_40561);
xor UO_564 (O_564,N_43624,N_42240);
or UO_565 (O_565,N_43837,N_40412);
and UO_566 (O_566,N_46232,N_45279);
or UO_567 (O_567,N_44517,N_42418);
nor UO_568 (O_568,N_48634,N_48617);
or UO_569 (O_569,N_45350,N_49605);
or UO_570 (O_570,N_47430,N_48501);
or UO_571 (O_571,N_40710,N_47722);
and UO_572 (O_572,N_41565,N_40310);
nand UO_573 (O_573,N_48687,N_44182);
xor UO_574 (O_574,N_49624,N_46123);
or UO_575 (O_575,N_47193,N_44177);
and UO_576 (O_576,N_41121,N_46725);
nand UO_577 (O_577,N_48193,N_41486);
and UO_578 (O_578,N_44058,N_44579);
and UO_579 (O_579,N_40169,N_49915);
nand UO_580 (O_580,N_44817,N_41463);
xor UO_581 (O_581,N_40514,N_48220);
nor UO_582 (O_582,N_47704,N_43953);
xnor UO_583 (O_583,N_45987,N_48827);
xor UO_584 (O_584,N_45597,N_40823);
nor UO_585 (O_585,N_46370,N_49109);
nor UO_586 (O_586,N_43473,N_40693);
nor UO_587 (O_587,N_45188,N_47852);
or UO_588 (O_588,N_49554,N_49861);
or UO_589 (O_589,N_47832,N_48480);
and UO_590 (O_590,N_44107,N_47541);
nor UO_591 (O_591,N_41949,N_41699);
or UO_592 (O_592,N_41971,N_45546);
nand UO_593 (O_593,N_44555,N_42216);
or UO_594 (O_594,N_48062,N_41053);
nand UO_595 (O_595,N_48806,N_46986);
and UO_596 (O_596,N_49544,N_46191);
xor UO_597 (O_597,N_48026,N_48005);
and UO_598 (O_598,N_47355,N_43841);
nand UO_599 (O_599,N_42705,N_49378);
nor UO_600 (O_600,N_43363,N_46657);
xnor UO_601 (O_601,N_40206,N_47155);
nand UO_602 (O_602,N_42655,N_42351);
nor UO_603 (O_603,N_40337,N_43004);
nor UO_604 (O_604,N_40739,N_43025);
and UO_605 (O_605,N_48910,N_42447);
nand UO_606 (O_606,N_42950,N_45968);
xnor UO_607 (O_607,N_46767,N_45620);
or UO_608 (O_608,N_45967,N_43708);
nand UO_609 (O_609,N_47710,N_46778);
nand UO_610 (O_610,N_46450,N_42357);
or UO_611 (O_611,N_48947,N_46763);
xor UO_612 (O_612,N_44494,N_46451);
xnor UO_613 (O_613,N_46311,N_44340);
or UO_614 (O_614,N_48908,N_45125);
or UO_615 (O_615,N_42439,N_41066);
or UO_616 (O_616,N_41233,N_47803);
nand UO_617 (O_617,N_46405,N_40518);
nand UO_618 (O_618,N_49611,N_49308);
nor UO_619 (O_619,N_48006,N_49392);
xor UO_620 (O_620,N_49618,N_43171);
nor UO_621 (O_621,N_41725,N_46255);
or UO_622 (O_622,N_44803,N_40718);
and UO_623 (O_623,N_44935,N_48820);
or UO_624 (O_624,N_45762,N_41997);
nand UO_625 (O_625,N_47108,N_49976);
and UO_626 (O_626,N_43361,N_40098);
nor UO_627 (O_627,N_49094,N_47449);
xnor UO_628 (O_628,N_43120,N_45774);
or UO_629 (O_629,N_48444,N_47843);
and UO_630 (O_630,N_47510,N_43008);
nand UO_631 (O_631,N_46400,N_42974);
nand UO_632 (O_632,N_40974,N_48847);
nand UO_633 (O_633,N_40713,N_45696);
nor UO_634 (O_634,N_47146,N_40821);
nor UO_635 (O_635,N_46798,N_47498);
xnor UO_636 (O_636,N_42795,N_40311);
and UO_637 (O_637,N_44059,N_45587);
and UO_638 (O_638,N_44183,N_43028);
and UO_639 (O_639,N_45788,N_48939);
nor UO_640 (O_640,N_44899,N_48351);
and UO_641 (O_641,N_42293,N_46052);
xor UO_642 (O_642,N_44462,N_48021);
nor UO_643 (O_643,N_47955,N_48145);
xor UO_644 (O_644,N_49524,N_49942);
or UO_645 (O_645,N_42321,N_46839);
or UO_646 (O_646,N_41400,N_44521);
nand UO_647 (O_647,N_48553,N_41228);
or UO_648 (O_648,N_47354,N_43487);
or UO_649 (O_649,N_41619,N_45474);
nor UO_650 (O_650,N_43332,N_40165);
nand UO_651 (O_651,N_46467,N_40673);
nand UO_652 (O_652,N_45330,N_46988);
nand UO_653 (O_653,N_45705,N_44838);
or UO_654 (O_654,N_45988,N_40626);
xnor UO_655 (O_655,N_46004,N_45085);
nor UO_656 (O_656,N_43867,N_43851);
or UO_657 (O_657,N_42701,N_48438);
nor UO_658 (O_658,N_40912,N_42921);
nand UO_659 (O_659,N_40528,N_48487);
nand UO_660 (O_660,N_47539,N_48597);
xnor UO_661 (O_661,N_46720,N_49836);
or UO_662 (O_662,N_43111,N_48424);
nand UO_663 (O_663,N_43944,N_49833);
xnor UO_664 (O_664,N_41990,N_44194);
or UO_665 (O_665,N_47952,N_41610);
nand UO_666 (O_666,N_47944,N_47422);
nor UO_667 (O_667,N_47425,N_49528);
nor UO_668 (O_668,N_46632,N_41604);
or UO_669 (O_669,N_47024,N_40182);
xor UO_670 (O_670,N_46458,N_43910);
and UO_671 (O_671,N_41641,N_44581);
nand UO_672 (O_672,N_45770,N_41730);
nand UO_673 (O_673,N_42122,N_49479);
or UO_674 (O_674,N_49198,N_49916);
or UO_675 (O_675,N_47978,N_43866);
nor UO_676 (O_676,N_44563,N_47693);
nand UO_677 (O_677,N_48043,N_42678);
or UO_678 (O_678,N_40783,N_42312);
and UO_679 (O_679,N_45274,N_42392);
nand UO_680 (O_680,N_48814,N_45189);
and UO_681 (O_681,N_43931,N_46568);
or UO_682 (O_682,N_44784,N_48008);
nor UO_683 (O_683,N_47322,N_46116);
or UO_684 (O_684,N_40335,N_41507);
and UO_685 (O_685,N_43503,N_42964);
or UO_686 (O_686,N_41914,N_45864);
xor UO_687 (O_687,N_40858,N_45486);
or UO_688 (O_688,N_47841,N_41413);
nor UO_689 (O_689,N_46643,N_46034);
xor UO_690 (O_690,N_47582,N_48207);
xor UO_691 (O_691,N_45371,N_49829);
nor UO_692 (O_692,N_44878,N_44043);
nor UO_693 (O_693,N_45160,N_47143);
nand UO_694 (O_694,N_44293,N_43142);
nand UO_695 (O_695,N_43817,N_42470);
nand UO_696 (O_696,N_42702,N_49160);
nand UO_697 (O_697,N_45659,N_40772);
nor UO_698 (O_698,N_47604,N_40106);
or UO_699 (O_699,N_49330,N_45807);
and UO_700 (O_700,N_46495,N_41929);
and UO_701 (O_701,N_40185,N_46751);
or UO_702 (O_702,N_49871,N_45542);
nor UO_703 (O_703,N_47971,N_49646);
nor UO_704 (O_704,N_48753,N_41100);
nand UO_705 (O_705,N_47054,N_43375);
nand UO_706 (O_706,N_46338,N_41904);
and UO_707 (O_707,N_42751,N_40432);
nor UO_708 (O_708,N_49459,N_41292);
nor UO_709 (O_709,N_40831,N_48666);
xnor UO_710 (O_710,N_42986,N_43052);
nand UO_711 (O_711,N_42560,N_41252);
nand UO_712 (O_712,N_40844,N_41316);
nor UO_713 (O_713,N_41688,N_46049);
nor UO_714 (O_714,N_49933,N_49502);
nor UO_715 (O_715,N_41017,N_43968);
or UO_716 (O_716,N_45873,N_41147);
xor UO_717 (O_717,N_42830,N_44287);
nand UO_718 (O_718,N_48802,N_48307);
nor UO_719 (O_719,N_48338,N_46199);
and UO_720 (O_720,N_43815,N_47187);
and UO_721 (O_721,N_49169,N_49532);
nor UO_722 (O_722,N_41040,N_47237);
nor UO_723 (O_723,N_40829,N_44347);
xnor UO_724 (O_724,N_46551,N_49958);
or UO_725 (O_725,N_46180,N_40825);
or UO_726 (O_726,N_46590,N_44736);
or UO_727 (O_727,N_46288,N_40131);
xnor UO_728 (O_728,N_47596,N_44877);
nand UO_729 (O_729,N_47605,N_49020);
xor UO_730 (O_730,N_42505,N_41985);
and UO_731 (O_731,N_47468,N_48917);
nor UO_732 (O_732,N_49334,N_40085);
and UO_733 (O_733,N_40476,N_48391);
xnor UO_734 (O_734,N_47999,N_49283);
and UO_735 (O_735,N_48340,N_42156);
or UO_736 (O_736,N_42818,N_46411);
nor UO_737 (O_737,N_45591,N_47036);
and UO_738 (O_738,N_43994,N_48188);
or UO_739 (O_739,N_40840,N_41864);
and UO_740 (O_740,N_42434,N_40149);
and UO_741 (O_741,N_41981,N_46494);
or UO_742 (O_742,N_47097,N_45934);
or UO_743 (O_743,N_47764,N_44074);
nor UO_744 (O_744,N_43999,N_40607);
nor UO_745 (O_745,N_40437,N_41617);
nor UO_746 (O_746,N_43828,N_46755);
xnor UO_747 (O_747,N_48813,N_44002);
and UO_748 (O_748,N_47767,N_42596);
xnor UO_749 (O_749,N_45216,N_46661);
and UO_750 (O_750,N_46481,N_43647);
nand UO_751 (O_751,N_45457,N_44629);
nor UO_752 (O_752,N_46965,N_47371);
and UO_753 (O_753,N_41762,N_47601);
or UO_754 (O_754,N_42512,N_45197);
and UO_755 (O_755,N_46908,N_49523);
nor UO_756 (O_756,N_43221,N_43790);
nand UO_757 (O_757,N_44934,N_45375);
xnor UO_758 (O_758,N_48073,N_47540);
or UO_759 (O_759,N_41171,N_42589);
nand UO_760 (O_760,N_40221,N_44178);
nand UO_761 (O_761,N_42119,N_40860);
nand UO_762 (O_762,N_49906,N_43921);
xor UO_763 (O_763,N_41952,N_42030);
xnor UO_764 (O_764,N_46072,N_43644);
nor UO_765 (O_765,N_47021,N_42226);
nand UO_766 (O_766,N_45813,N_42592);
or UO_767 (O_767,N_41458,N_40647);
and UO_768 (O_768,N_44367,N_41238);
nand UO_769 (O_769,N_49010,N_40556);
nand UO_770 (O_770,N_43124,N_46649);
nor UO_771 (O_771,N_47670,N_43592);
nor UO_772 (O_772,N_47489,N_45837);
nor UO_773 (O_773,N_47810,N_41712);
xor UO_774 (O_774,N_40211,N_42554);
xor UO_775 (O_775,N_40895,N_47472);
nor UO_776 (O_776,N_44569,N_45684);
nor UO_777 (O_777,N_42675,N_46019);
nand UO_778 (O_778,N_49941,N_46823);
or UO_779 (O_779,N_42207,N_43279);
or UO_780 (O_780,N_45440,N_47001);
nor UO_781 (O_781,N_41210,N_46516);
xor UO_782 (O_782,N_45896,N_44328);
nand UO_783 (O_783,N_48615,N_46089);
nand UO_784 (O_784,N_48231,N_40992);
xnor UO_785 (O_785,N_44669,N_47584);
nor UO_786 (O_786,N_42429,N_45702);
nand UO_787 (O_787,N_44823,N_48137);
xnor UO_788 (O_788,N_47789,N_45019);
and UO_789 (O_789,N_49375,N_46845);
nor UO_790 (O_790,N_49249,N_47110);
nand UO_791 (O_791,N_43879,N_49563);
nor UO_792 (O_792,N_43182,N_45212);
or UO_793 (O_793,N_44573,N_46997);
nor UO_794 (O_794,N_46848,N_43622);
or UO_795 (O_795,N_43946,N_48705);
nor UO_796 (O_796,N_41248,N_43554);
xnor UO_797 (O_797,N_42274,N_47628);
or UO_798 (O_798,N_43981,N_45936);
and UO_799 (O_799,N_45134,N_41556);
or UO_800 (O_800,N_47282,N_44275);
nand UO_801 (O_801,N_41324,N_47549);
nand UO_802 (O_802,N_40341,N_40256);
nand UO_803 (O_803,N_45183,N_45261);
xnor UO_804 (O_804,N_46009,N_43245);
nand UO_805 (O_805,N_46357,N_41531);
or UO_806 (O_806,N_45914,N_41675);
xnor UO_807 (O_807,N_40262,N_48909);
nor UO_808 (O_808,N_46857,N_42817);
nand UO_809 (O_809,N_47643,N_48772);
nand UO_810 (O_810,N_47771,N_40397);
nor UO_811 (O_811,N_43237,N_45139);
nor UO_812 (O_812,N_47845,N_43571);
and UO_813 (O_813,N_49152,N_40938);
nand UO_814 (O_814,N_40411,N_48442);
nor UO_815 (O_815,N_49301,N_48561);
nor UO_816 (O_816,N_46078,N_45066);
nor UO_817 (O_817,N_41048,N_40032);
nand UO_818 (O_818,N_41944,N_40041);
xnor UO_819 (O_819,N_48815,N_41785);
and UO_820 (O_820,N_48521,N_48983);
nor UO_821 (O_821,N_44171,N_43317);
nand UO_822 (O_822,N_42428,N_44289);
nand UO_823 (O_823,N_42499,N_42065);
nand UO_824 (O_824,N_46283,N_45608);
nand UO_825 (O_825,N_42542,N_44094);
nor UO_826 (O_826,N_44734,N_43039);
nor UO_827 (O_827,N_42059,N_48948);
or UO_828 (O_828,N_46492,N_46605);
nor UO_829 (O_829,N_48014,N_43811);
and UO_830 (O_830,N_46913,N_41211);
or UO_831 (O_831,N_41163,N_43576);
or UO_832 (O_832,N_44338,N_48892);
and UO_833 (O_833,N_41010,N_42302);
nand UO_834 (O_834,N_49314,N_49243);
nand UO_835 (O_835,N_46901,N_40595);
or UO_836 (O_836,N_47975,N_42849);
xnor UO_837 (O_837,N_41057,N_47287);
or UO_838 (O_838,N_45283,N_49442);
xnor UO_839 (O_839,N_41494,N_43857);
nand UO_840 (O_840,N_42845,N_46514);
and UO_841 (O_841,N_44111,N_45879);
or UO_842 (O_842,N_40019,N_44958);
and UO_843 (O_843,N_43648,N_45044);
and UO_844 (O_844,N_41866,N_44682);
xor UO_845 (O_845,N_42815,N_44758);
xor UO_846 (O_846,N_48413,N_40254);
nor UO_847 (O_847,N_48662,N_43497);
nand UO_848 (O_848,N_44679,N_47268);
nand UO_849 (O_849,N_44301,N_46929);
or UO_850 (O_850,N_42669,N_48124);
xor UO_851 (O_851,N_47518,N_41232);
xnor UO_852 (O_852,N_40678,N_46182);
nor UO_853 (O_853,N_44159,N_43626);
and UO_854 (O_854,N_47929,N_48055);
nand UO_855 (O_855,N_44256,N_46817);
nor UO_856 (O_856,N_45435,N_41460);
xnor UO_857 (O_857,N_41963,N_46882);
and UO_858 (O_858,N_49790,N_42707);
nor UO_859 (O_859,N_49670,N_45939);
and UO_860 (O_860,N_46380,N_42556);
xnor UO_861 (O_861,N_44288,N_49513);
nor UO_862 (O_862,N_40158,N_42049);
or UO_863 (O_863,N_45531,N_47685);
nand UO_864 (O_864,N_41824,N_49167);
nor UO_865 (O_865,N_46474,N_46404);
or UO_866 (O_866,N_45412,N_48680);
nand UO_867 (O_867,N_48980,N_40543);
and UO_868 (O_868,N_46264,N_47692);
nor UO_869 (O_869,N_45106,N_47056);
nand UO_870 (O_870,N_41428,N_47622);
xnor UO_871 (O_871,N_42555,N_41177);
nand UO_872 (O_872,N_49907,N_40736);
nand UO_873 (O_873,N_46391,N_47139);
and UO_874 (O_874,N_41165,N_48796);
nand UO_875 (O_875,N_47448,N_43560);
xor UO_876 (O_876,N_47114,N_43839);
nor UO_877 (O_877,N_45242,N_46512);
or UO_878 (O_878,N_49363,N_46260);
or UO_879 (O_879,N_40777,N_46699);
nor UO_880 (O_880,N_41168,N_42183);
nor UO_881 (O_881,N_44833,N_43581);
xor UO_882 (O_882,N_41807,N_44163);
xor UO_883 (O_883,N_41244,N_40805);
nand UO_884 (O_884,N_41272,N_48448);
nand UO_885 (O_885,N_48135,N_40264);
xor UO_886 (O_886,N_46342,N_49059);
or UO_887 (O_887,N_48508,N_45158);
nand UO_888 (O_888,N_48181,N_49164);
or UO_889 (O_889,N_43380,N_40653);
and UO_890 (O_890,N_42105,N_41493);
nand UO_891 (O_891,N_47863,N_42612);
xor UO_892 (O_892,N_47969,N_48789);
or UO_893 (O_893,N_43699,N_43187);
nand UO_894 (O_894,N_45438,N_48626);
nor UO_895 (O_895,N_47946,N_45081);
or UO_896 (O_896,N_46559,N_43156);
or UO_897 (O_897,N_47124,N_45806);
nand UO_898 (O_898,N_47953,N_46853);
and UO_899 (O_899,N_46810,N_48383);
or UO_900 (O_900,N_43014,N_42693);
nand UO_901 (O_901,N_43964,N_40968);
xnor UO_902 (O_902,N_49943,N_47745);
or UO_903 (O_903,N_48819,N_47550);
xor UO_904 (O_904,N_46209,N_44609);
nand UO_905 (O_905,N_48064,N_44047);
and UO_906 (O_906,N_49305,N_49666);
nor UO_907 (O_907,N_47446,N_40716);
and UO_908 (O_908,N_40554,N_48237);
or UO_909 (O_909,N_42015,N_48544);
and UO_910 (O_910,N_44550,N_40478);
xor UO_911 (O_911,N_43288,N_41563);
nand UO_912 (O_912,N_45695,N_44722);
nor UO_913 (O_913,N_42791,N_41830);
and UO_914 (O_914,N_45624,N_48911);
and UO_915 (O_915,N_42464,N_42248);
and UO_916 (O_916,N_48527,N_46142);
or UO_917 (O_917,N_49187,N_46291);
or UO_918 (O_918,N_41058,N_43407);
and UO_919 (O_919,N_44919,N_40836);
and UO_920 (O_920,N_45692,N_45601);
nand UO_921 (O_921,N_41039,N_43646);
and UO_922 (O_922,N_45582,N_41481);
nand UO_923 (O_923,N_40290,N_45726);
or UO_924 (O_924,N_40231,N_40724);
or UO_925 (O_925,N_43054,N_44297);
or UO_926 (O_926,N_42896,N_49977);
nor UO_927 (O_927,N_47820,N_44319);
and UO_928 (O_928,N_48270,N_47466);
xor UO_929 (O_929,N_40241,N_40843);
xnor UO_930 (O_930,N_43740,N_45177);
or UO_931 (O_931,N_40147,N_40464);
nand UO_932 (O_932,N_45054,N_43316);
and UO_933 (O_933,N_44499,N_45867);
xor UO_934 (O_934,N_40492,N_42873);
or UO_935 (O_935,N_47026,N_45547);
and UO_936 (O_936,N_46730,N_47250);
xor UO_937 (O_937,N_40361,N_41151);
nand UO_938 (O_938,N_43838,N_41964);
xnor UO_939 (O_939,N_46150,N_44549);
or UO_940 (O_940,N_44608,N_42528);
xnor UO_941 (O_941,N_42588,N_42303);
nand UO_942 (O_942,N_41596,N_47739);
nand UO_943 (O_943,N_48585,N_44457);
nand UO_944 (O_944,N_44488,N_42039);
nand UO_945 (O_945,N_46144,N_48765);
xor UO_946 (O_946,N_41142,N_41632);
and UO_947 (O_947,N_49430,N_48194);
nand UO_948 (O_948,N_41320,N_46834);
nor UO_949 (O_949,N_44825,N_44017);
xnor UO_950 (O_950,N_45859,N_48841);
xor UO_951 (O_951,N_41284,N_46083);
or UO_952 (O_952,N_44354,N_42967);
and UO_953 (O_953,N_45970,N_43445);
xnor UO_954 (O_954,N_42955,N_41710);
xnor UO_955 (O_955,N_42762,N_49190);
nor UO_956 (O_956,N_44087,N_41298);
or UO_957 (O_957,N_45032,N_48373);
nor UO_958 (O_958,N_48618,N_40497);
xnor UO_959 (O_959,N_48660,N_41331);
nand UO_960 (O_960,N_40145,N_45152);
or UO_961 (O_961,N_49206,N_48563);
and UO_962 (O_962,N_41921,N_47493);
and UO_963 (O_963,N_42047,N_44269);
or UO_964 (O_964,N_46515,N_47032);
nor UO_965 (O_965,N_44619,N_41367);
nand UO_966 (O_966,N_48879,N_42228);
or UO_967 (O_967,N_42694,N_45504);
xnor UO_968 (O_968,N_44441,N_41261);
and UO_969 (O_969,N_45824,N_45039);
nand UO_970 (O_970,N_48859,N_42462);
nor UO_971 (O_971,N_41333,N_49180);
nand UO_972 (O_972,N_46324,N_44678);
xnor UO_973 (O_973,N_40494,N_45021);
nor UO_974 (O_974,N_40928,N_44262);
nand UO_975 (O_975,N_43122,N_41145);
nand UO_976 (O_976,N_40029,N_41343);
nor UO_977 (O_977,N_46310,N_43333);
xor UO_978 (O_978,N_45856,N_49689);
xnor UO_979 (O_979,N_42295,N_47825);
nand UO_980 (O_980,N_42352,N_46620);
nor UO_981 (O_981,N_40121,N_46912);
or UO_982 (O_982,N_45272,N_45998);
xor UO_983 (O_983,N_47052,N_41411);
nor UO_984 (O_984,N_46969,N_49515);
nand UO_985 (O_985,N_49511,N_49197);
nand UO_986 (O_986,N_42443,N_42225);
nor UO_987 (O_987,N_46200,N_47947);
and UO_988 (O_988,N_41650,N_40570);
or UO_989 (O_989,N_41424,N_42613);
or UO_990 (O_990,N_44942,N_49885);
xnor UO_991 (O_991,N_42810,N_45609);
nand UO_992 (O_992,N_47811,N_49510);
nor UO_993 (O_993,N_47528,N_44463);
xnor UO_994 (O_994,N_42679,N_49904);
or UO_995 (O_995,N_40503,N_41153);
nand UO_996 (O_996,N_41334,N_43270);
nand UO_997 (O_997,N_48408,N_46682);
xnor UO_998 (O_998,N_44041,N_43421);
and UO_999 (O_999,N_47431,N_43666);
nand UO_1000 (O_1000,N_47461,N_43805);
nor UO_1001 (O_1001,N_49340,N_44460);
or UO_1002 (O_1002,N_41445,N_49509);
or UO_1003 (O_1003,N_47889,N_46769);
nand UO_1004 (O_1004,N_42268,N_42609);
nor UO_1005 (O_1005,N_44254,N_46502);
nor UO_1006 (O_1006,N_45510,N_41614);
or UO_1007 (O_1007,N_40377,N_43495);
and UO_1008 (O_1008,N_42223,N_48787);
or UO_1009 (O_1009,N_48533,N_43416);
and UO_1010 (O_1010,N_47583,N_48367);
or UO_1011 (O_1011,N_49846,N_46133);
and UO_1012 (O_1012,N_43432,N_46146);
xor UO_1013 (O_1013,N_48344,N_46301);
or UO_1014 (O_1014,N_44064,N_42852);
and UO_1015 (O_1015,N_46794,N_44807);
nand UO_1016 (O_1016,N_47105,N_48938);
nor UO_1017 (O_1017,N_41161,N_42835);
or UO_1018 (O_1018,N_46711,N_46565);
or UO_1019 (O_1019,N_45462,N_42237);
or UO_1020 (O_1020,N_41377,N_47762);
nand UO_1021 (O_1021,N_43545,N_43573);
nand UO_1022 (O_1022,N_46702,N_44813);
and UO_1023 (O_1023,N_43321,N_42365);
nand UO_1024 (O_1024,N_46082,N_40405);
nor UO_1025 (O_1025,N_49046,N_47980);
and UO_1026 (O_1026,N_46156,N_49063);
nand UO_1027 (O_1027,N_46031,N_46861);
xor UO_1028 (O_1028,N_43026,N_47086);
and UO_1029 (O_1029,N_49389,N_43701);
xnor UO_1030 (O_1030,N_44642,N_45654);
or UO_1031 (O_1031,N_46285,N_46819);
nand UO_1032 (O_1032,N_49993,N_49543);
nand UO_1033 (O_1033,N_47578,N_46795);
or UO_1034 (O_1034,N_48289,N_47031);
nand UO_1035 (O_1035,N_41347,N_47211);
xnor UO_1036 (O_1036,N_41093,N_44874);
nand UO_1037 (O_1037,N_48076,N_44762);
xnor UO_1038 (O_1038,N_41906,N_46299);
xor UO_1039 (O_1039,N_49232,N_45167);
nor UO_1040 (O_1040,N_40054,N_49451);
nor UO_1041 (O_1041,N_49406,N_42306);
or UO_1042 (O_1042,N_43294,N_48121);
nand UO_1043 (O_1043,N_40788,N_45418);
or UO_1044 (O_1044,N_40279,N_45802);
or UO_1045 (O_1045,N_43426,N_46676);
nor UO_1046 (O_1046,N_49422,N_42779);
nor UO_1047 (O_1047,N_42046,N_49795);
or UO_1048 (O_1048,N_40789,N_47680);
or UO_1049 (O_1049,N_45577,N_41170);
or UO_1050 (O_1050,N_44860,N_48038);
or UO_1051 (O_1051,N_44315,N_49471);
nor UO_1052 (O_1052,N_48930,N_48435);
nor UO_1053 (O_1053,N_44447,N_44027);
nor UO_1054 (O_1054,N_41050,N_48130);
xor UO_1055 (O_1055,N_45666,N_43510);
or UO_1056 (O_1056,N_41810,N_43422);
or UO_1057 (O_1057,N_49615,N_46962);
or UO_1058 (O_1058,N_44118,N_49702);
nor UO_1059 (O_1059,N_41538,N_41357);
and UO_1060 (O_1060,N_41222,N_42718);
nor UO_1061 (O_1061,N_44103,N_47251);
nand UO_1062 (O_1062,N_41651,N_40014);
nor UO_1063 (O_1063,N_46942,N_40958);
xnor UO_1064 (O_1064,N_48966,N_48828);
or UO_1065 (O_1065,N_49357,N_49228);
or UO_1066 (O_1066,N_49225,N_41871);
nor UO_1067 (O_1067,N_44119,N_43723);
nor UO_1068 (O_1068,N_48972,N_49291);
and UO_1069 (O_1069,N_43865,N_40441);
xnor UO_1070 (O_1070,N_42859,N_42468);
or UO_1071 (O_1071,N_40506,N_46589);
nand UO_1072 (O_1072,N_45982,N_41860);
xor UO_1073 (O_1073,N_45901,N_42517);
nand UO_1074 (O_1074,N_44539,N_46352);
nand UO_1075 (O_1075,N_48569,N_44792);
and UO_1076 (O_1076,N_44388,N_46497);
or UO_1077 (O_1077,N_42205,N_42048);
nand UO_1078 (O_1078,N_46488,N_40418);
nand UO_1079 (O_1079,N_49880,N_47337);
or UO_1080 (O_1080,N_41101,N_44100);
or UO_1081 (O_1081,N_48821,N_48603);
and UO_1082 (O_1082,N_42355,N_42918);
nor UO_1083 (O_1083,N_45434,N_40596);
nor UO_1084 (O_1084,N_40606,N_45571);
or UO_1085 (O_1085,N_46915,N_48282);
xor UO_1086 (O_1086,N_48816,N_46781);
and UO_1087 (O_1087,N_46193,N_42668);
nand UO_1088 (O_1088,N_44113,N_46464);
nand UO_1089 (O_1089,N_43203,N_44248);
and UO_1090 (O_1090,N_49720,N_48697);
nor UO_1091 (O_1091,N_46761,N_44806);
and UO_1092 (O_1092,N_44497,N_47118);
nor UO_1093 (O_1093,N_41957,N_48041);
and UO_1094 (O_1094,N_41580,N_43357);
and UO_1095 (O_1095,N_48737,N_48184);
or UO_1096 (O_1096,N_48803,N_46208);
or UO_1097 (O_1097,N_41181,N_47395);
or UO_1098 (O_1098,N_43988,N_49546);
nand UO_1099 (O_1099,N_45227,N_45205);
nand UO_1100 (O_1100,N_49011,N_40787);
xnor UO_1101 (O_1101,N_49685,N_46626);
or UO_1102 (O_1102,N_46496,N_41141);
and UO_1103 (O_1103,N_41328,N_48534);
xnor UO_1104 (O_1104,N_49185,N_48138);
and UO_1105 (O_1105,N_45868,N_48257);
xnor UO_1106 (O_1106,N_43466,N_43572);
nand UO_1107 (O_1107,N_46074,N_40880);
or UO_1108 (O_1108,N_48368,N_42953);
nand UO_1109 (O_1109,N_49984,N_40404);
nand UO_1110 (O_1110,N_46563,N_43597);
nor UO_1111 (O_1111,N_45024,N_47965);
nor UO_1112 (O_1112,N_48492,N_46837);
and UO_1113 (O_1113,N_48199,N_42399);
xor UO_1114 (O_1114,N_44018,N_44747);
and UO_1115 (O_1115,N_41795,N_47503);
nand UO_1116 (O_1116,N_45776,N_48912);
nor UO_1117 (O_1117,N_49044,N_49800);
and UO_1118 (O_1118,N_44634,N_44520);
or UO_1119 (O_1119,N_48230,N_48846);
nor UO_1120 (O_1120,N_48799,N_49455);
nor UO_1121 (O_1121,N_40802,N_49522);
nand UO_1122 (O_1122,N_42627,N_48003);
and UO_1123 (O_1123,N_41004,N_45607);
nand UO_1124 (O_1124,N_47546,N_43086);
and UO_1125 (O_1125,N_44756,N_42400);
and UO_1126 (O_1126,N_40243,N_41758);
xnor UO_1127 (O_1127,N_41126,N_47304);
and UO_1128 (O_1128,N_40646,N_45651);
nor UO_1129 (O_1129,N_48822,N_49730);
or UO_1130 (O_1130,N_42880,N_45954);
xor UO_1131 (O_1131,N_49457,N_48875);
xor UO_1132 (O_1132,N_46598,N_46241);
nor UO_1133 (O_1133,N_42963,N_45373);
nor UO_1134 (O_1134,N_48356,N_41961);
or UO_1135 (O_1135,N_40579,N_41260);
xnor UO_1136 (O_1136,N_40376,N_43377);
or UO_1137 (O_1137,N_44451,N_43892);
nand UO_1138 (O_1138,N_48851,N_48667);
nor UO_1139 (O_1139,N_41558,N_49402);
and UO_1140 (O_1140,N_43049,N_47352);
and UO_1141 (O_1141,N_42419,N_44051);
nor UO_1142 (O_1142,N_47694,N_45952);
nor UO_1143 (O_1143,N_41243,N_41267);
nor UO_1144 (O_1144,N_45525,N_48365);
nor UO_1145 (O_1145,N_41927,N_40303);
xor UO_1146 (O_1146,N_45057,N_48986);
xor UO_1147 (O_1147,N_49721,N_40820);
nand UO_1148 (O_1148,N_44996,N_41621);
and UO_1149 (O_1149,N_44021,N_45595);
or UO_1150 (O_1150,N_48190,N_46873);
and UO_1151 (O_1151,N_49257,N_46791);
xor UO_1152 (O_1152,N_49850,N_48401);
or UO_1153 (O_1153,N_46374,N_44730);
or UO_1154 (O_1154,N_40137,N_40941);
xnor UO_1155 (O_1155,N_49892,N_42664);
nand UO_1156 (O_1156,N_42754,N_42670);
xor UO_1157 (O_1157,N_47729,N_46972);
xor UO_1158 (O_1158,N_49274,N_41018);
nand UO_1159 (O_1159,N_47662,N_42118);
xor UO_1160 (O_1160,N_42531,N_46167);
xor UO_1161 (O_1161,N_46106,N_47234);
xnor UO_1162 (O_1162,N_40306,N_42271);
or UO_1163 (O_1163,N_42123,N_47827);
nand UO_1164 (O_1164,N_46591,N_41900);
and UO_1165 (O_1165,N_45619,N_45828);
or UO_1166 (O_1166,N_42252,N_44729);
or UO_1167 (O_1167,N_48169,N_41459);
xnor UO_1168 (O_1168,N_44258,N_49703);
xnor UO_1169 (O_1169,N_40676,N_47900);
and UO_1170 (O_1170,N_41280,N_40435);
nand UO_1171 (O_1171,N_41182,N_44954);
xnor UO_1172 (O_1172,N_43273,N_44052);
and UO_1173 (O_1173,N_43404,N_47494);
nor UO_1174 (O_1174,N_45581,N_49367);
xnor UO_1175 (O_1175,N_40261,N_43526);
nor UO_1176 (O_1176,N_48094,N_44044);
or UO_1177 (O_1177,N_42145,N_43860);
or UO_1178 (O_1178,N_46724,N_48472);
nand UO_1179 (O_1179,N_46235,N_48372);
xnor UO_1180 (O_1180,N_41110,N_46331);
nand UO_1181 (O_1181,N_40101,N_45515);
and UO_1182 (O_1182,N_47129,N_42244);
or UO_1183 (O_1183,N_48885,N_40569);
or UO_1184 (O_1184,N_44929,N_41700);
nor UO_1185 (O_1185,N_40017,N_42339);
nand UO_1186 (O_1186,N_47123,N_44691);
and UO_1187 (O_1187,N_43209,N_40318);
xor UO_1188 (O_1188,N_43737,N_48366);
xor UO_1189 (O_1189,N_42722,N_42546);
nand UO_1190 (O_1190,N_49078,N_43507);
and UO_1191 (O_1191,N_47652,N_42219);
xor UO_1192 (O_1192,N_40146,N_47261);
nor UO_1193 (O_1193,N_49137,N_44473);
or UO_1194 (O_1194,N_40991,N_48285);
nor UO_1195 (O_1195,N_43087,N_44959);
xor UO_1196 (O_1196,N_48221,N_48608);
nor UO_1197 (O_1197,N_43185,N_44271);
nor UO_1198 (O_1198,N_43257,N_44733);
xor UO_1199 (O_1199,N_48160,N_43941);
xor UO_1200 (O_1200,N_46040,N_46967);
nand UO_1201 (O_1201,N_49796,N_45387);
or UO_1202 (O_1202,N_45410,N_42102);
nand UO_1203 (O_1203,N_45778,N_43463);
xor UO_1204 (O_1204,N_43206,N_45391);
nor UO_1205 (O_1205,N_49394,N_45075);
and UO_1206 (O_1206,N_48153,N_49366);
xor UO_1207 (O_1207,N_45402,N_42822);
nor UO_1208 (O_1208,N_48520,N_41317);
nand UO_1209 (O_1209,N_42927,N_40993);
xor UO_1210 (O_1210,N_42521,N_47573);
and UO_1211 (O_1211,N_47859,N_45176);
or UO_1212 (O_1212,N_48621,N_42895);
nand UO_1213 (O_1213,N_41546,N_48291);
or UO_1214 (O_1214,N_48397,N_40064);
nor UO_1215 (O_1215,N_47273,N_49066);
and UO_1216 (O_1216,N_45989,N_43556);
and UO_1217 (O_1217,N_47886,N_49093);
xnor UO_1218 (O_1218,N_41721,N_43514);
or UO_1219 (O_1219,N_45109,N_40422);
or UO_1220 (O_1220,N_43830,N_45122);
or UO_1221 (O_1221,N_44716,N_45413);
nor UO_1222 (O_1222,N_41148,N_43146);
nand UO_1223 (O_1223,N_49696,N_45603);
nand UO_1224 (O_1224,N_42243,N_43891);
nor UO_1225 (O_1225,N_45063,N_49909);
nand UO_1226 (O_1226,N_44529,N_41175);
nand UO_1227 (O_1227,N_40036,N_47168);
nor UO_1228 (O_1228,N_47757,N_45078);
or UO_1229 (O_1229,N_40870,N_42929);
and UO_1230 (O_1230,N_43157,N_49655);
xnor UO_1231 (O_1231,N_43406,N_41060);
or UO_1232 (O_1232,N_48332,N_41008);
or UO_1233 (O_1233,N_40205,N_43019);
or UO_1234 (O_1234,N_48623,N_48502);
nor UO_1235 (O_1235,N_40620,N_44295);
nand UO_1236 (O_1236,N_42977,N_40853);
nand UO_1237 (O_1237,N_46007,N_47807);
nand UO_1238 (O_1238,N_48878,N_43411);
xor UO_1239 (O_1239,N_43846,N_44427);
and UO_1240 (O_1240,N_48818,N_46041);
nand UO_1241 (O_1241,N_46412,N_48210);
or UO_1242 (O_1242,N_47260,N_49092);
nand UO_1243 (O_1243,N_49156,N_41802);
or UO_1244 (O_1244,N_43085,N_49583);
or UO_1245 (O_1245,N_46732,N_47350);
xor UO_1246 (O_1246,N_44472,N_44464);
nand UO_1247 (O_1247,N_45008,N_41288);
and UO_1248 (O_1248,N_43105,N_48536);
and UO_1249 (O_1249,N_47100,N_48785);
and UO_1250 (O_1250,N_48782,N_46910);
and UO_1251 (O_1251,N_45826,N_49781);
or UO_1252 (O_1252,N_48771,N_47053);
nor UO_1253 (O_1253,N_43334,N_45400);
and UO_1254 (O_1254,N_45612,N_41191);
nor UO_1255 (O_1255,N_45289,N_42804);
nand UO_1256 (O_1256,N_47270,N_40511);
and UO_1257 (O_1257,N_47831,N_44137);
and UO_1258 (O_1258,N_49994,N_47400);
nand UO_1259 (O_1259,N_48312,N_49709);
or UO_1260 (O_1260,N_41796,N_41826);
nor UO_1261 (O_1261,N_42446,N_47735);
or UO_1262 (O_1262,N_49210,N_44852);
xor UO_1263 (O_1263,N_40118,N_45880);
and UO_1264 (O_1264,N_42635,N_42686);
nand UO_1265 (O_1265,N_41593,N_41054);
nor UO_1266 (O_1266,N_45324,N_40586);
nand UO_1267 (O_1267,N_47587,N_43736);
or UO_1268 (O_1268,N_42500,N_49127);
nor UO_1269 (O_1269,N_45238,N_45629);
xor UO_1270 (O_1270,N_41630,N_42594);
and UO_1271 (O_1271,N_41042,N_48514);
nor UO_1272 (O_1272,N_41082,N_41372);
and UO_1273 (O_1273,N_40217,N_48676);
or UO_1274 (O_1274,N_45707,N_42485);
nand UO_1275 (O_1275,N_47249,N_49954);
and UO_1276 (O_1276,N_44072,N_45519);
nand UO_1277 (O_1277,N_40933,N_44205);
xor UO_1278 (O_1278,N_44847,N_43779);
and UO_1279 (O_1279,N_41599,N_40237);
xnor UO_1280 (O_1280,N_47703,N_44356);
or UO_1281 (O_1281,N_44411,N_48495);
and UO_1282 (O_1282,N_41117,N_46453);
or UO_1283 (O_1283,N_44470,N_40480);
and UO_1284 (O_1284,N_43785,N_40632);
nor UO_1285 (O_1285,N_47419,N_43285);
nor UO_1286 (O_1286,N_45842,N_43119);
nor UO_1287 (O_1287,N_47170,N_49918);
xnor UO_1288 (O_1288,N_46975,N_45220);
xnor UO_1289 (O_1289,N_42087,N_45295);
nor UO_1290 (O_1290,N_42294,N_43993);
or UO_1291 (O_1291,N_49360,N_42124);
nor UO_1292 (O_1292,N_46526,N_41777);
nand UO_1293 (O_1293,N_44889,N_47085);
xnor UO_1294 (O_1294,N_42035,N_45447);
nand UO_1295 (O_1295,N_41477,N_49446);
nor UO_1296 (O_1296,N_42265,N_49686);
nand UO_1297 (O_1297,N_49296,N_46013);
xor UO_1298 (O_1298,N_45354,N_45288);
or UO_1299 (O_1299,N_42350,N_45265);
and UO_1300 (O_1300,N_48794,N_46298);
nor UO_1301 (O_1301,N_46105,N_45804);
nor UO_1302 (O_1302,N_47802,N_45154);
and UO_1303 (O_1303,N_44562,N_49956);
nand UO_1304 (O_1304,N_40001,N_41659);
xnor UO_1305 (O_1305,N_43158,N_49443);
or UO_1306 (O_1306,N_40797,N_43799);
xnor UO_1307 (O_1307,N_43914,N_49401);
nand UO_1308 (O_1308,N_49516,N_42618);
nand UO_1309 (O_1309,N_47196,N_44294);
nor UO_1310 (O_1310,N_48142,N_46418);
nor UO_1311 (O_1311,N_43403,N_43658);
xnor UO_1312 (O_1312,N_40758,N_44324);
or UO_1313 (O_1313,N_40451,N_40666);
or UO_1314 (O_1314,N_42287,N_45870);
xor UO_1315 (O_1315,N_41447,N_42262);
or UO_1316 (O_1316,N_46442,N_46425);
or UO_1317 (O_1317,N_48775,N_49238);
or UO_1318 (O_1318,N_44554,N_48430);
nor UO_1319 (O_1319,N_46576,N_49591);
nand UO_1320 (O_1320,N_40473,N_43251);
nor UO_1321 (O_1321,N_45669,N_44602);
or UO_1322 (O_1322,N_43293,N_47214);
nor UO_1323 (O_1323,N_44162,N_44842);
xnor UO_1324 (O_1324,N_47087,N_46875);
xor UO_1325 (O_1325,N_47246,N_46673);
nor UO_1326 (O_1326,N_46435,N_43476);
xor UO_1327 (O_1327,N_41255,N_41585);
and UO_1328 (O_1328,N_48769,N_40180);
xor UO_1329 (O_1329,N_41278,N_47663);
or UO_1330 (O_1330,N_45439,N_48973);
and UO_1331 (O_1331,N_49279,N_40099);
nor UO_1332 (O_1332,N_46766,N_49967);
nor UO_1333 (O_1333,N_45819,N_45598);
nor UO_1334 (O_1334,N_47659,N_43439);
nand UO_1335 (O_1335,N_40559,N_46640);
and UO_1336 (O_1336,N_46367,N_40572);
nand UO_1337 (O_1337,N_49560,N_45745);
and UO_1338 (O_1338,N_41960,N_46630);
nor UO_1339 (O_1339,N_41901,N_42591);
or UO_1340 (O_1340,N_47842,N_49318);
nand UO_1341 (O_1341,N_44116,N_43744);
and UO_1342 (O_1342,N_42725,N_40796);
or UO_1343 (O_1343,N_44022,N_41341);
and UO_1344 (O_1344,N_47599,N_46993);
and UO_1345 (O_1345,N_45815,N_40203);
and UO_1346 (O_1346,N_44033,N_44930);
nor UO_1347 (O_1347,N_45681,N_42332);
nand UO_1348 (O_1348,N_40851,N_40498);
nand UO_1349 (O_1349,N_43696,N_47856);
nand UO_1350 (O_1350,N_46186,N_49600);
or UO_1351 (O_1351,N_45113,N_47858);
or UO_1352 (O_1352,N_42537,N_47415);
nor UO_1353 (O_1353,N_42736,N_47175);
xor UO_1354 (O_1354,N_47064,N_44568);
or UO_1355 (O_1355,N_49822,N_44788);
xor UO_1356 (O_1356,N_46647,N_47404);
nor UO_1357 (O_1357,N_49759,N_44941);
nor UO_1358 (O_1358,N_46454,N_40648);
nand UO_1359 (O_1359,N_44413,N_40916);
nor UO_1360 (O_1360,N_45572,N_44888);
or UO_1361 (O_1361,N_41799,N_45477);
xor UO_1362 (O_1362,N_48283,N_42577);
nor UO_1363 (O_1363,N_45906,N_42923);
xnor UO_1364 (O_1364,N_46187,N_48460);
nand UO_1365 (O_1365,N_43164,N_48952);
nand UO_1366 (O_1366,N_44211,N_43930);
and UO_1367 (O_1367,N_45799,N_46529);
or UO_1368 (O_1368,N_43376,N_41633);
and UO_1369 (O_1369,N_46243,N_42099);
nor UO_1370 (O_1370,N_44897,N_46953);
nor UO_1371 (O_1371,N_46762,N_43585);
xor UO_1372 (O_1372,N_47368,N_46043);
or UO_1373 (O_1373,N_41337,N_46204);
and UO_1374 (O_1374,N_42843,N_46039);
or UO_1375 (O_1375,N_48080,N_43452);
and UO_1376 (O_1376,N_43296,N_45613);
and UO_1377 (O_1377,N_46650,N_43939);
or UO_1378 (O_1378,N_45792,N_46295);
xnor UO_1379 (O_1379,N_48715,N_45029);
nand UO_1380 (O_1380,N_41408,N_46415);
and UO_1381 (O_1381,N_48427,N_40150);
nor UO_1382 (O_1382,N_48150,N_45211);
or UO_1383 (O_1383,N_43308,N_45458);
nor UO_1384 (O_1384,N_47200,N_41545);
nand UO_1385 (O_1385,N_40688,N_44189);
nor UO_1386 (O_1386,N_49579,N_49269);
or UO_1387 (O_1387,N_46548,N_43388);
and UO_1388 (O_1388,N_41415,N_47976);
xnor UO_1389 (O_1389,N_49328,N_48151);
and UO_1390 (O_1390,N_46721,N_42184);
nor UO_1391 (O_1391,N_48186,N_47950);
or UO_1392 (O_1392,N_43665,N_47015);
and UO_1393 (O_1393,N_43725,N_49520);
nand UO_1394 (O_1394,N_47117,N_44660);
and UO_1395 (O_1395,N_41162,N_42478);
nor UO_1396 (O_1396,N_45888,N_47515);
and UO_1397 (O_1397,N_40752,N_44279);
nand UO_1398 (O_1398,N_45723,N_49342);
and UO_1399 (O_1399,N_43496,N_43552);
or UO_1400 (O_1400,N_48762,N_41645);
nand UO_1401 (O_1401,N_45363,N_44831);
nand UO_1402 (O_1402,N_46990,N_45454);
nand UO_1403 (O_1403,N_40548,N_46961);
and UO_1404 (O_1404,N_43190,N_49467);
or UO_1405 (O_1405,N_48935,N_44800);
nor UO_1406 (O_1406,N_48462,N_49004);
xnor UO_1407 (O_1407,N_42770,N_41898);
or UO_1408 (O_1408,N_43153,N_41834);
nor UO_1409 (O_1409,N_49529,N_42563);
and UO_1410 (O_1410,N_44624,N_41709);
nand UO_1411 (O_1411,N_40955,N_46740);
xnor UO_1412 (O_1412,N_46992,N_43342);
nand UO_1413 (O_1413,N_49142,N_43225);
or UO_1414 (O_1414,N_41061,N_47967);
nor UO_1415 (O_1415,N_47611,N_46333);
nand UO_1416 (O_1416,N_49348,N_41421);
or UO_1417 (O_1417,N_46843,N_43232);
xor UO_1418 (O_1418,N_48504,N_44623);
nor UO_1419 (O_1419,N_48359,N_44442);
or UO_1420 (O_1420,N_40824,N_47661);
or UO_1421 (O_1421,N_45810,N_43082);
or UO_1422 (O_1422,N_46566,N_43532);
nor UO_1423 (O_1423,N_44591,N_41670);
nand UO_1424 (O_1424,N_48314,N_41258);
or UO_1425 (O_1425,N_48699,N_41766);
or UO_1426 (O_1426,N_44102,N_43722);
and UO_1427 (O_1427,N_43777,N_46188);
nand UO_1428 (O_1428,N_42695,N_41793);
nand UO_1429 (O_1429,N_49986,N_48159);
xnor UO_1430 (O_1430,N_46077,N_45098);
and UO_1431 (O_1431,N_44068,N_40487);
nand UO_1432 (O_1432,N_44524,N_40902);
nand UO_1433 (O_1433,N_47766,N_46202);
nor UO_1434 (O_1434,N_46957,N_42239);
xnor UO_1435 (O_1435,N_40770,N_46343);
nand UO_1436 (O_1436,N_40563,N_40618);
nand UO_1437 (O_1437,N_41208,N_41083);
nand UO_1438 (O_1438,N_48831,N_41865);
nor UO_1439 (O_1439,N_40449,N_47286);
and UO_1440 (O_1440,N_40738,N_48030);
nor UO_1441 (O_1441,N_48873,N_43906);
and UO_1442 (O_1442,N_49439,N_46215);
and UO_1443 (O_1443,N_41578,N_44154);
or UO_1444 (O_1444,N_42173,N_42771);
nor UO_1445 (O_1445,N_47382,N_42979);
or UO_1446 (O_1446,N_41131,N_40198);
xnor UO_1447 (O_1447,N_49466,N_40504);
nor UO_1448 (O_1448,N_40462,N_42982);
or UO_1449 (O_1449,N_43467,N_48652);
or UO_1450 (O_1450,N_42376,N_42421);
and UO_1451 (O_1451,N_40994,N_49476);
nand UO_1452 (O_1452,N_45847,N_45490);
and UO_1453 (O_1453,N_45637,N_44385);
nor UO_1454 (O_1454,N_42057,N_44228);
nor UO_1455 (O_1455,N_48213,N_41088);
nand UO_1456 (O_1456,N_45554,N_42677);
or UO_1457 (O_1457,N_41892,N_49068);
or UO_1458 (O_1458,N_47240,N_46363);
nand UO_1459 (O_1459,N_42971,N_44845);
nor UO_1460 (O_1460,N_40553,N_46131);
nor UO_1461 (O_1461,N_43728,N_45809);
and UO_1462 (O_1462,N_48631,N_41649);
xor UO_1463 (O_1463,N_49362,N_41025);
nand UO_1464 (O_1464,N_45203,N_49140);
or UO_1465 (O_1465,N_44056,N_45370);
nand UO_1466 (O_1466,N_49344,N_43650);
and UO_1467 (O_1467,N_46500,N_42002);
and UO_1468 (O_1468,N_44586,N_46212);
or UO_1469 (O_1469,N_41682,N_45599);
nor UO_1470 (O_1470,N_49019,N_40213);
xor UO_1471 (O_1471,N_47690,N_48118);
or UO_1472 (O_1472,N_42700,N_49022);
nand UO_1473 (O_1473,N_48403,N_44156);
nor UO_1474 (O_1474,N_45213,N_48012);
nand UO_1475 (O_1475,N_43635,N_49133);
and UO_1476 (O_1476,N_49679,N_44717);
xor UO_1477 (O_1477,N_46807,N_49945);
and UO_1478 (O_1478,N_49704,N_44779);
nand UO_1479 (O_1479,N_49682,N_45463);
xnor UO_1480 (O_1480,N_44443,N_43079);
and UO_1481 (O_1481,N_48638,N_44818);
or UO_1482 (O_1482,N_44143,N_43013);
xor UO_1483 (O_1483,N_45580,N_47908);
and UO_1484 (O_1484,N_44732,N_41965);
xnor UO_1485 (O_1485,N_40509,N_40977);
xor UO_1486 (O_1486,N_40225,N_49369);
and UO_1487 (O_1487,N_44204,N_45084);
and UO_1488 (O_1488,N_42659,N_40284);
nand UO_1489 (O_1489,N_46428,N_47559);
xnor UO_1490 (O_1490,N_40088,N_44028);
nand UO_1491 (O_1491,N_46518,N_40025);
or UO_1492 (O_1492,N_41285,N_49859);
and UO_1493 (O_1493,N_48428,N_48896);
xnor UO_1494 (O_1494,N_44688,N_49997);
xnor UO_1495 (O_1495,N_42723,N_47733);
nand UO_1496 (O_1496,N_46321,N_45604);
xor UO_1497 (O_1497,N_46637,N_47712);
and UO_1498 (O_1498,N_48249,N_47907);
nand UO_1499 (O_1499,N_48748,N_47324);
nand UO_1500 (O_1500,N_48899,N_45821);
xnor UO_1501 (O_1501,N_45303,N_45253);
nand UO_1502 (O_1502,N_47280,N_40201);
nor UO_1503 (O_1503,N_40874,N_45481);
nor UO_1504 (O_1504,N_48906,N_42385);
or UO_1505 (O_1505,N_42854,N_48777);
nand UO_1506 (O_1506,N_49733,N_46642);
nand UO_1507 (O_1507,N_49865,N_42452);
xor UO_1508 (O_1508,N_47336,N_40087);
or UO_1509 (O_1509,N_46323,N_46353);
or UO_1510 (O_1510,N_49749,N_46542);
or UO_1511 (O_1511,N_45299,N_43872);
nand UO_1512 (O_1512,N_41899,N_43996);
and UO_1513 (O_1513,N_41917,N_42169);
or UO_1514 (O_1514,N_42186,N_43358);
xor UO_1515 (O_1515,N_45362,N_48458);
nor UO_1516 (O_1516,N_44088,N_44701);
nor UO_1517 (O_1517,N_47855,N_45832);
nand UO_1518 (O_1518,N_46930,N_48148);
and UO_1519 (O_1519,N_42930,N_41251);
nor UO_1520 (O_1520,N_43616,N_40555);
nor UO_1521 (O_1521,N_47376,N_43278);
xnor UO_1522 (O_1522,N_44920,N_46140);
and UO_1523 (O_1523,N_49480,N_45268);
and UO_1524 (O_1524,N_40745,N_46371);
or UO_1525 (O_1525,N_48708,N_47367);
nor UO_1526 (O_1526,N_48581,N_48422);
xnor UO_1527 (O_1527,N_43922,N_46689);
xnor UO_1528 (O_1528,N_40388,N_45963);
nand UO_1529 (O_1529,N_44993,N_41577);
nor UO_1530 (O_1530,N_47655,N_43290);
nor UO_1531 (O_1531,N_47713,N_45575);
nand UO_1532 (O_1532,N_44063,N_44174);
and UO_1533 (O_1533,N_42251,N_40077);
nor UO_1534 (O_1534,N_43428,N_40760);
or UO_1535 (O_1535,N_49036,N_42431);
nor UO_1536 (O_1536,N_46012,N_47378);
and UO_1537 (O_1537,N_42960,N_44225);
or UO_1538 (O_1538,N_45862,N_45893);
and UO_1539 (O_1539,N_40807,N_47255);
nand UO_1540 (O_1540,N_40706,N_48682);
nand UO_1541 (O_1541,N_49649,N_48202);
or UO_1542 (O_1542,N_47176,N_45548);
xnor UO_1543 (O_1543,N_48470,N_46087);
nand UO_1544 (O_1544,N_42704,N_47830);
and UO_1545 (O_1545,N_49863,N_49973);
or UO_1546 (O_1546,N_48594,N_41195);
and UO_1547 (O_1547,N_44862,N_46789);
nand UO_1548 (O_1548,N_49265,N_46263);
nor UO_1549 (O_1549,N_45497,N_44106);
xnor UO_1550 (O_1550,N_40040,N_46303);
and UO_1551 (O_1551,N_48522,N_43135);
nand UO_1552 (O_1552,N_48109,N_40990);
nor UO_1553 (O_1553,N_44965,N_47669);
and UO_1554 (O_1554,N_48212,N_45045);
and UO_1555 (O_1555,N_44767,N_40624);
nor UO_1556 (O_1556,N_40015,N_41611);
or UO_1557 (O_1557,N_41090,N_46085);
xor UO_1558 (O_1558,N_44546,N_47416);
nor UO_1559 (O_1559,N_40104,N_40965);
nor UO_1560 (O_1560,N_48645,N_48406);
nand UO_1561 (O_1561,N_49060,N_49486);
nand UO_1562 (O_1562,N_43908,N_43351);
nor UO_1563 (O_1563,N_44768,N_40757);
and UO_1564 (O_1564,N_49115,N_45834);
or UO_1565 (O_1565,N_41975,N_45444);
xnor UO_1566 (O_1566,N_45911,N_48746);
or UO_1567 (O_1567,N_48596,N_46717);
nand UO_1568 (O_1568,N_43707,N_45704);
nor UO_1569 (O_1569,N_45335,N_48317);
and UO_1570 (O_1570,N_49900,N_43107);
or UO_1571 (O_1571,N_47580,N_43747);
nor UO_1572 (O_1572,N_42249,N_44487);
nand UO_1573 (O_1573,N_47456,N_43692);
nor UO_1574 (O_1574,N_47959,N_42425);
and UO_1575 (O_1575,N_48387,N_41313);
nand UO_1576 (O_1576,N_47674,N_44128);
nand UO_1577 (O_1577,N_42507,N_40744);
and UO_1578 (O_1578,N_45957,N_47966);
nor UO_1579 (O_1579,N_45505,N_46738);
and UO_1580 (O_1580,N_47447,N_40360);
nand UO_1581 (O_1581,N_49938,N_40866);
and UO_1582 (O_1582,N_49534,N_49083);
and UO_1583 (O_1583,N_40578,N_48385);
nand UO_1584 (O_1584,N_40966,N_47615);
or UO_1585 (O_1585,N_44444,N_43115);
nand UO_1586 (O_1586,N_48555,N_42422);
or UO_1587 (O_1587,N_40691,N_45302);
nand UO_1588 (O_1588,N_41376,N_48506);
and UO_1589 (O_1589,N_48858,N_43529);
nand UO_1590 (O_1590,N_48091,N_46067);
or UO_1591 (O_1591,N_42308,N_43703);
and UO_1592 (O_1592,N_40608,N_40194);
or UO_1593 (O_1593,N_46694,N_40291);
xor UO_1594 (O_1594,N_41206,N_49110);
and UO_1595 (O_1595,N_45489,N_46835);
or UO_1596 (O_1596,N_47979,N_46318);
nor UO_1597 (O_1597,N_45761,N_42343);
xnor UO_1598 (O_1598,N_42384,N_49910);
nor UO_1599 (O_1599,N_48066,N_49824);
xnor UO_1600 (O_1600,N_41660,N_49413);
or UO_1601 (O_1601,N_45526,N_46332);
and UO_1602 (O_1602,N_44992,N_44931);
or UO_1603 (O_1603,N_49248,N_40157);
and UO_1604 (O_1604,N_40519,N_44667);
nand UO_1605 (O_1605,N_48260,N_45328);
nor UO_1606 (O_1606,N_44393,N_42121);
and UO_1607 (O_1607,N_48059,N_46775);
and UO_1608 (O_1608,N_48788,N_45077);
or UO_1609 (O_1609,N_45922,N_42012);
and UO_1610 (O_1610,N_43518,N_46830);
nor UO_1611 (O_1611,N_47379,N_43804);
nor UO_1612 (O_1612,N_46939,N_48734);
xnor UO_1613 (O_1613,N_44266,N_43651);
or UO_1614 (O_1614,N_43818,N_41591);
and UO_1615 (O_1615,N_49207,N_47188);
xor UO_1616 (O_1616,N_49390,N_43155);
or UO_1617 (O_1617,N_47135,N_40452);
xnor UO_1618 (O_1618,N_48240,N_47768);
and UO_1619 (O_1619,N_43760,N_46407);
xor UO_1620 (O_1620,N_45121,N_42214);
and UO_1621 (O_1621,N_41027,N_43345);
and UO_1622 (O_1622,N_40142,N_49143);
nand UO_1623 (O_1623,N_46525,N_42882);
xor UO_1624 (O_1624,N_49267,N_47911);
and UO_1625 (O_1625,N_45625,N_42838);
nor UO_1626 (O_1626,N_42753,N_48900);
nor UO_1627 (O_1627,N_40909,N_47266);
xor UO_1628 (O_1628,N_42427,N_47029);
and UO_1629 (O_1629,N_48293,N_43854);
nor UO_1630 (O_1630,N_47402,N_48960);
xor UO_1631 (O_1631,N_41550,N_44883);
and UO_1632 (O_1632,N_46715,N_48132);
nand UO_1633 (O_1633,N_40074,N_43762);
nand UO_1634 (O_1634,N_46373,N_47780);
xor UO_1635 (O_1635,N_46712,N_44953);
nand UO_1636 (O_1636,N_46841,N_46687);
nand UO_1637 (O_1637,N_42272,N_40546);
and UO_1638 (O_1638,N_41978,N_45876);
xor UO_1639 (O_1639,N_40274,N_45117);
or UO_1640 (O_1640,N_44861,N_46897);
and UO_1641 (O_1641,N_43566,N_48017);
or UO_1642 (O_1642,N_48234,N_44694);
or UO_1643 (O_1643,N_46714,N_46149);
nor UO_1644 (O_1644,N_48795,N_42839);
and UO_1645 (O_1645,N_44938,N_41532);
xnor UO_1646 (O_1646,N_47169,N_49778);
and UO_1647 (O_1647,N_43230,N_44968);
xor UO_1648 (O_1648,N_49772,N_49914);
xor UO_1649 (O_1649,N_40505,N_46616);
nand UO_1650 (O_1650,N_42863,N_45071);
nand UO_1651 (O_1651,N_45769,N_49032);
nor UO_1652 (O_1652,N_41772,N_44872);
and UO_1653 (O_1653,N_41359,N_46899);
or UO_1654 (O_1654,N_49746,N_40617);
and UO_1655 (O_1655,N_46088,N_46998);
or UO_1656 (O_1656,N_47882,N_46268);
nand UO_1657 (O_1657,N_45780,N_47977);
and UO_1658 (O_1658,N_43834,N_46718);
and UO_1659 (O_1659,N_47302,N_49912);
and UO_1660 (O_1660,N_42382,N_41695);
xnor UO_1661 (O_1661,N_45141,N_43689);
and UO_1662 (O_1662,N_48872,N_47731);
nand UO_1663 (O_1663,N_42994,N_46037);
nor UO_1664 (O_1664,N_48053,N_48180);
xor UO_1665 (O_1665,N_46865,N_44144);
xnor UO_1666 (O_1666,N_46387,N_40436);
and UO_1667 (O_1667,N_45437,N_40062);
nand UO_1668 (O_1668,N_43241,N_46104);
nor UO_1669 (O_1669,N_43010,N_42378);
nand UO_1670 (O_1670,N_47897,N_46886);
or UO_1671 (O_1671,N_47728,N_48633);
and UO_1672 (O_1672,N_40238,N_48035);
xnor UO_1673 (O_1673,N_43609,N_43742);
nor UO_1674 (O_1674,N_41465,N_48889);
xor UO_1675 (O_1675,N_45461,N_44913);
and UO_1676 (O_1676,N_49136,N_48865);
nor UO_1677 (O_1677,N_42585,N_40631);
or UO_1678 (O_1678,N_44155,N_49435);
nand UO_1679 (O_1679,N_42944,N_49189);
and UO_1680 (O_1680,N_46524,N_42862);
nand UO_1681 (O_1681,N_46399,N_46960);
nand UO_1682 (O_1682,N_48719,N_41575);
or UO_1683 (O_1683,N_48447,N_42129);
xnor UO_1684 (O_1684,N_42728,N_42380);
nand UO_1685 (O_1685,N_49565,N_47050);
and UO_1686 (O_1686,N_43593,N_43385);
xnor UO_1687 (O_1687,N_41536,N_42535);
or UO_1688 (O_1688,N_47613,N_44508);
nand UO_1689 (O_1689,N_40799,N_44314);
and UO_1690 (O_1690,N_48854,N_41374);
or UO_1691 (O_1691,N_43017,N_41761);
or UO_1692 (O_1692,N_40900,N_48431);
xor UO_1693 (O_1693,N_47473,N_41158);
or UO_1694 (O_1694,N_44865,N_40707);
or UO_1695 (O_1695,N_46553,N_43980);
and UO_1696 (O_1696,N_48489,N_48056);
xnor UO_1697 (O_1697,N_43883,N_47727);
nor UO_1698 (O_1698,N_45757,N_45352);
or UO_1699 (O_1699,N_40155,N_47983);
or UO_1700 (O_1700,N_48604,N_48564);
or UO_1701 (O_1701,N_48276,N_46022);
nand UO_1702 (O_1702,N_44887,N_47254);
and UO_1703 (O_1703,N_43179,N_45997);
xor UO_1704 (O_1704,N_49497,N_48836);
xor UO_1705 (O_1705,N_43752,N_40976);
and UO_1706 (O_1706,N_47717,N_49968);
xnor UO_1707 (O_1707,N_49498,N_45118);
nor UO_1708 (O_1708,N_45785,N_45257);
nor UO_1709 (O_1709,N_41993,N_40406);
nor UO_1710 (O_1710,N_45102,N_46001);
or UO_1711 (O_1711,N_40513,N_43174);
xor UO_1712 (O_1712,N_40566,N_48371);
and UO_1713 (O_1713,N_43608,N_41844);
nor UO_1714 (O_1714,N_48915,N_41200);
and UO_1715 (O_1715,N_49444,N_46493);
xor UO_1716 (O_1716,N_42259,N_44867);
or UO_1717 (O_1717,N_48217,N_48644);
or UO_1718 (O_1718,N_43031,N_44449);
nor UO_1719 (O_1719,N_43033,N_47236);
xnor UO_1720 (O_1720,N_45451,N_41598);
nand UO_1721 (O_1721,N_41922,N_46091);
or UO_1722 (O_1722,N_46991,N_41063);
or UO_1723 (O_1723,N_43977,N_42871);
nand UO_1724 (O_1724,N_41704,N_47864);
or UO_1725 (O_1725,N_41035,N_45560);
and UO_1726 (O_1726,N_40508,N_43450);
xnor UO_1727 (O_1727,N_49722,N_48829);
or UO_1728 (O_1728,N_45060,N_45677);
and UO_1729 (O_1729,N_48485,N_46101);
nor UO_1730 (O_1730,N_45415,N_47119);
nand UO_1731 (O_1731,N_49852,N_47157);
xnor UO_1732 (O_1732,N_44773,N_42456);
and UO_1733 (O_1733,N_40141,N_45340);
and UO_1734 (O_1734,N_40589,N_48022);
nor UO_1735 (O_1735,N_44596,N_43046);
and UO_1736 (O_1736,N_41942,N_48071);
xor UO_1737 (O_1737,N_40065,N_45877);
xnor UO_1738 (O_1738,N_48946,N_46641);
and UO_1739 (O_1739,N_46831,N_43177);
and UO_1740 (O_1740,N_47410,N_41939);
nor UO_1741 (O_1741,N_40656,N_48997);
or UO_1742 (O_1742,N_48866,N_47088);
or UO_1743 (O_1743,N_43292,N_47391);
xor UO_1744 (O_1744,N_43359,N_45180);
xnor UO_1745 (O_1745,N_43056,N_40512);
nor UO_1746 (O_1746,N_44832,N_46377);
nand UO_1747 (O_1747,N_49965,N_47833);
nor UO_1748 (O_1748,N_48027,N_45897);
xnor UO_1749 (O_1749,N_46674,N_46513);
or UO_1750 (O_1750,N_46904,N_45553);
or UO_1751 (O_1751,N_41085,N_40461);
and UO_1752 (O_1752,N_48861,N_48685);
or UO_1753 (O_1753,N_44471,N_48171);
nand UO_1754 (O_1754,N_43896,N_44766);
or UO_1755 (O_1755,N_44436,N_49370);
nor UO_1756 (O_1756,N_42004,N_41877);
nor UO_1757 (O_1757,N_40944,N_45933);
or UO_1758 (O_1758,N_47645,N_40012);
xor UO_1759 (O_1759,N_44377,N_44791);
or UO_1760 (O_1760,N_45333,N_45605);
nand UO_1761 (O_1761,N_46856,N_49988);
or UO_1762 (O_1762,N_42990,N_49660);
or UO_1763 (O_1763,N_47565,N_49374);
nor UO_1764 (O_1764,N_40803,N_40245);
and UO_1765 (O_1765,N_47594,N_42458);
nand UO_1766 (O_1766,N_46706,N_46635);
xor UO_1767 (O_1767,N_44045,N_41266);
nand UO_1768 (O_1768,N_46925,N_40067);
xnor UO_1769 (O_1769,N_49598,N_46523);
and UO_1770 (O_1770,N_44386,N_42112);
xor UO_1771 (O_1771,N_41270,N_47560);
or UO_1772 (O_1772,N_41742,N_42187);
xor UO_1773 (O_1773,N_49163,N_46764);
xor UO_1774 (O_1774,N_48923,N_45339);
or UO_1775 (O_1775,N_48850,N_45403);
xor UO_1776 (O_1776,N_49359,N_44950);
or UO_1777 (O_1777,N_49321,N_44927);
xnor UO_1778 (O_1778,N_41729,N_48612);
nor UO_1779 (O_1779,N_41746,N_49313);
and UO_1780 (O_1780,N_40365,N_47066);
and UO_1781 (O_1781,N_41476,N_41562);
nor UO_1782 (O_1782,N_42735,N_42665);
nand UO_1783 (O_1783,N_40053,N_43840);
xor UO_1784 (O_1784,N_40321,N_45752);
xor UO_1785 (O_1785,N_48096,N_41674);
and UO_1786 (O_1786,N_47912,N_47082);
and UO_1787 (O_1787,N_45635,N_49923);
and UO_1788 (O_1788,N_40792,N_40364);
or UO_1789 (O_1789,N_46073,N_45961);
nand UO_1790 (O_1790,N_47838,N_45534);
and UO_1791 (O_1791,N_46096,N_46227);
and UO_1792 (O_1792,N_41435,N_49643);
and UO_1793 (O_1793,N_48625,N_47284);
xor UO_1794 (O_1794,N_45317,N_40571);
xnor UO_1795 (O_1795,N_43275,N_43094);
nand UO_1796 (O_1796,N_46325,N_43091);
or UO_1797 (O_1797,N_40193,N_41224);
xor UO_1798 (O_1798,N_44024,N_48756);
or UO_1799 (O_1799,N_45023,N_45394);
or UO_1800 (O_1800,N_46327,N_40174);
nand UO_1801 (O_1801,N_46139,N_46477);
nor UO_1802 (O_1802,N_43173,N_43682);
or UO_1803 (O_1803,N_42925,N_40943);
xor UO_1804 (O_1804,N_45985,N_49031);
nand UO_1805 (O_1805,N_43548,N_40599);
and UO_1806 (O_1806,N_48325,N_48256);
nor UO_1807 (O_1807,N_43400,N_48974);
and UO_1808 (O_1808,N_47935,N_48410);
nor UO_1809 (O_1809,N_46741,N_41745);
and UO_1810 (O_1810,N_49204,N_42494);
and UO_1811 (O_1811,N_43844,N_49974);
xnor UO_1812 (O_1812,N_47586,N_42299);
and UO_1813 (O_1813,N_44884,N_49400);
nor UO_1814 (O_1814,N_48877,N_42614);
nor UO_1815 (O_1815,N_48070,N_47821);
or UO_1816 (O_1816,N_41038,N_47177);
nand UO_1817 (O_1817,N_41979,N_43349);
or UO_1818 (O_1818,N_47027,N_41021);
nor UO_1819 (O_1819,N_46369,N_47743);
nand UO_1820 (O_1820,N_42388,N_45187);
xor UO_1821 (O_1821,N_42054,N_49971);
or UO_1822 (O_1822,N_43511,N_48302);
nor UO_1823 (O_1823,N_49951,N_42805);
xnor UO_1824 (O_1824,N_48711,N_42296);
and UO_1825 (O_1825,N_44459,N_46097);
or UO_1826 (O_1826,N_45765,N_42920);
nor UO_1827 (O_1827,N_41759,N_49625);
and UO_1828 (O_1828,N_43138,N_42806);
or UO_1829 (O_1829,N_47245,N_48575);
xnor UO_1830 (O_1830,N_44790,N_47308);
or UO_1831 (O_1831,N_49387,N_42496);
and UO_1832 (O_1832,N_46633,N_47746);
or UO_1833 (O_1833,N_43226,N_44697);
xnor UO_1834 (O_1834,N_44235,N_40793);
nor UO_1835 (O_1835,N_40111,N_48954);
and UO_1836 (O_1836,N_45823,N_43224);
or UO_1837 (O_1837,N_48139,N_48573);
nand UO_1838 (O_1838,N_40674,N_47719);
or UO_1839 (O_1839,N_44402,N_48206);
or UO_1840 (O_1840,N_42394,N_49091);
and UO_1841 (O_1841,N_42626,N_42856);
nand UO_1842 (O_1842,N_49569,N_49713);
nor UO_1843 (O_1843,N_48976,N_45114);
and UO_1844 (O_1844,N_45913,N_45584);
or UO_1845 (O_1845,N_47753,N_49295);
nand UO_1846 (O_1846,N_48197,N_47403);
xor UO_1847 (O_1847,N_48229,N_47405);
or UO_1848 (O_1848,N_49410,N_46129);
nor UO_1849 (O_1849,N_40695,N_42329);
or UO_1850 (O_1850,N_41658,N_48523);
nor UO_1851 (O_1851,N_43515,N_49352);
or UO_1852 (O_1852,N_49594,N_46955);
or UO_1853 (O_1853,N_45460,N_48316);
and UO_1854 (O_1854,N_41774,N_47529);
nand UO_1855 (O_1855,N_43659,N_46756);
nor UO_1856 (O_1856,N_49405,N_41429);
or UO_1857 (O_1857,N_44277,N_44003);
nor UO_1858 (O_1858,N_49983,N_43197);
or UO_1859 (O_1859,N_41925,N_47149);
nand UO_1860 (O_1860,N_41947,N_42890);
xnor UO_1861 (O_1861,N_47490,N_43268);
nor UO_1862 (O_1862,N_42127,N_46700);
nand UO_1863 (O_1863,N_43926,N_45544);
nor UO_1864 (O_1864,N_44426,N_46328);
nand UO_1865 (O_1865,N_47487,N_42304);
xnor UO_1866 (O_1866,N_43850,N_48937);
xnor UO_1867 (O_1867,N_41433,N_40852);
xnor UO_1868 (O_1868,N_41179,N_44490);
nor UO_1869 (O_1869,N_46606,N_40300);
nand UO_1870 (O_1870,N_41816,N_40525);
or UO_1871 (O_1871,N_48894,N_40891);
and UO_1872 (O_1872,N_43574,N_46944);
or UO_1873 (O_1873,N_43075,N_46981);
nand UO_1874 (O_1874,N_41852,N_49957);
xnor UO_1875 (O_1875,N_41588,N_49432);
or UO_1876 (O_1876,N_40160,N_46030);
or UO_1877 (O_1877,N_49980,N_49872);
or UO_1878 (O_1878,N_48637,N_42134);
nand UO_1879 (O_1879,N_41183,N_43915);
or UO_1880 (O_1880,N_43048,N_46033);
nand UO_1881 (O_1881,N_49672,N_45321);
and UO_1882 (O_1882,N_42650,N_44272);
nor UO_1883 (O_1883,N_45478,N_43096);
or UO_1884 (O_1884,N_44924,N_41464);
xnor UO_1885 (O_1885,N_44940,N_47921);
nand UO_1886 (O_1886,N_42907,N_40597);
and UO_1887 (O_1887,N_43195,N_49105);
or UO_1888 (O_1888,N_49718,N_40766);
and UO_1889 (O_1889,N_44418,N_44988);
xor UO_1890 (O_1890,N_47536,N_46143);
or UO_1891 (O_1891,N_47179,N_47025);
and UO_1892 (O_1892,N_46294,N_45182);
nor UO_1893 (O_1893,N_46868,N_48628);
nor UO_1894 (O_1894,N_47229,N_43210);
nor UO_1895 (O_1895,N_41074,N_42033);
or UO_1896 (O_1896,N_47058,N_40791);
xor UO_1897 (O_1897,N_46320,N_41741);
nor UO_1898 (O_1898,N_45240,N_47805);
and UO_1899 (O_1899,N_43000,N_49123);
xor UO_1900 (O_1900,N_45527,N_49612);
or UO_1901 (O_1901,N_48376,N_40317);
nand UO_1902 (O_1902,N_47090,N_47800);
xnor UO_1903 (O_1903,N_47839,N_44666);
xnor UO_1904 (O_1904,N_47092,N_49628);
xnor UO_1905 (O_1905,N_48292,N_49013);
nor UO_1906 (O_1906,N_40664,N_44373);
or UO_1907 (O_1907,N_44062,N_44038);
and UO_1908 (O_1908,N_42250,N_42264);
nand UO_1909 (O_1909,N_44952,N_43663);
or UO_1910 (O_1910,N_40281,N_45993);
nor UO_1911 (O_1911,N_46665,N_49981);
xor UO_1912 (O_1912,N_47511,N_45294);
or UO_1913 (O_1913,N_43489,N_47080);
or UO_1914 (O_1914,N_46671,N_42199);
or UO_1915 (O_1915,N_47653,N_49445);
or UO_1916 (O_1916,N_41974,N_40733);
xnor UO_1917 (O_1917,N_48157,N_42502);
nor UO_1918 (O_1918,N_40905,N_45621);
nor UO_1919 (O_1919,N_49913,N_49636);
nor UO_1920 (O_1920,N_48250,N_47414);
or UO_1921 (O_1921,N_40771,N_44255);
nand UO_1922 (O_1922,N_47353,N_46322);
nand UO_1923 (O_1923,N_43071,N_45016);
nand UO_1924 (O_1924,N_40447,N_47385);
or UO_1925 (O_1925,N_46752,N_46050);
nor UO_1926 (O_1926,N_49869,N_42348);
nor UO_1927 (O_1927,N_42652,N_46893);
nor UO_1928 (O_1928,N_41499,N_48354);
nand UO_1929 (O_1929,N_45058,N_44425);
or UO_1930 (O_1930,N_45127,N_44984);
or UO_1931 (O_1931,N_45647,N_41137);
and UO_1932 (O_1932,N_47949,N_44689);
and UO_1933 (O_1933,N_41749,N_44320);
nor UO_1934 (O_1934,N_45035,N_42224);
nor UO_1935 (O_1935,N_47166,N_45322);
xnor UO_1936 (O_1936,N_46890,N_49212);
or UO_1937 (O_1937,N_41924,N_45747);
and UO_1938 (O_1938,N_43583,N_47338);
nand UO_1939 (O_1939,N_49697,N_46829);
or UO_1940 (O_1940,N_41345,N_49141);
nor UO_1941 (O_1941,N_49601,N_48390);
xnor UO_1942 (O_1942,N_47065,N_46046);
and UO_1943 (O_1943,N_48309,N_43687);
xor UO_1944 (O_1944,N_45009,N_48377);
nor UO_1945 (O_1945,N_42789,N_49391);
nor UO_1946 (O_1946,N_48219,N_42171);
and UO_1947 (O_1947,N_43771,N_47167);
or UO_1948 (O_1948,N_47542,N_47623);
and UO_1949 (O_1949,N_43677,N_42104);
nand UO_1950 (O_1950,N_46279,N_46573);
nor UO_1951 (O_1951,N_44727,N_42147);
nor UO_1952 (O_1952,N_48499,N_45329);
xor UO_1953 (O_1953,N_42761,N_42790);
nor UO_1954 (O_1954,N_46217,N_47267);
nand UO_1955 (O_1955,N_48505,N_42996);
nand UO_1956 (O_1956,N_47173,N_43144);
or UO_1957 (O_1957,N_49545,N_49810);
nor UO_1958 (O_1958,N_40251,N_46833);
nand UO_1959 (O_1959,N_44617,N_42368);
and UO_1960 (O_1960,N_48252,N_44975);
or UO_1961 (O_1961,N_47040,N_48981);
and UO_1962 (O_1962,N_42132,N_44853);
xnor UO_1963 (O_1963,N_42433,N_43695);
nand UO_1964 (O_1964,N_47386,N_44822);
xnor UO_1965 (O_1965,N_40176,N_49826);
xor UO_1966 (O_1966,N_49588,N_46427);
or UO_1967 (O_1967,N_41152,N_42687);
xor UO_1968 (O_1968,N_44395,N_43339);
and UO_1969 (O_1969,N_48538,N_49710);
nand UO_1970 (O_1970,N_49608,N_46517);
and UO_1971 (O_1971,N_41047,N_47047);
nor UO_1972 (O_1972,N_44124,N_44757);
and UO_1973 (O_1973,N_47342,N_43667);
or UO_1974 (O_1974,N_49813,N_43486);
and UO_1975 (O_1975,N_41485,N_44379);
and UO_1976 (O_1976,N_44949,N_46395);
nand UO_1977 (O_1977,N_48119,N_40120);
and UO_1978 (O_1978,N_44856,N_44298);
xnor UO_1979 (O_1979,N_49447,N_44140);
or UO_1980 (O_1980,N_44778,N_45169);
xor UO_1981 (O_1981,N_45653,N_40280);
nor UO_1982 (O_1982,N_45226,N_46996);
xor UO_1983 (O_1983,N_48738,N_40961);
nor UO_1984 (O_1984,N_49665,N_49055);
nand UO_1985 (O_1985,N_48677,N_44439);
and UO_1986 (O_1986,N_48919,N_49779);
nor UO_1987 (O_1987,N_40170,N_42085);
xnor UO_1988 (O_1988,N_40403,N_48029);
and UO_1989 (O_1989,N_47271,N_42136);
and UO_1990 (O_1990,N_46470,N_48651);
or UO_1991 (O_1991,N_40638,N_41045);
xor UO_1992 (O_1992,N_48593,N_48009);
nor UO_1993 (O_1993,N_44909,N_47325);
and UO_1994 (O_1994,N_45425,N_46881);
nor UO_1995 (O_1995,N_42125,N_40871);
nor UO_1996 (O_1996,N_46539,N_49631);
nand UO_1997 (O_1997,N_46384,N_44327);
nand UO_1998 (O_1998,N_42991,N_43438);
xnor UO_1999 (O_1999,N_40396,N_42869);
and UO_2000 (O_2000,N_43949,N_45562);
xor UO_2001 (O_2001,N_40650,N_45292);
and UO_2002 (O_2002,N_42931,N_41348);
xor UO_2003 (O_2003,N_45521,N_49897);
or UO_2004 (O_2004,N_49000,N_47013);
nand UO_2005 (O_2005,N_42796,N_49324);
or UO_2006 (O_2006,N_47195,N_49521);
and UO_2007 (O_2007,N_49819,N_49674);
and UO_2008 (O_2008,N_49590,N_40727);
nand UO_2009 (O_2009,N_41286,N_49888);
nand UO_2010 (O_2010,N_41954,N_44751);
and UO_2011 (O_2011,N_43324,N_48586);
or UO_2012 (O_2012,N_46340,N_46836);
nor UO_2013 (O_2013,N_43393,N_45170);
nor UO_2014 (O_2014,N_43200,N_44199);
xor UO_2015 (O_2015,N_45812,N_48659);
xor UO_2016 (O_2016,N_43460,N_42178);
nand UO_2017 (O_2017,N_47741,N_49088);
nor UO_2018 (O_2018,N_44662,N_42086);
nor UO_2019 (O_2019,N_41827,N_49581);
nand UO_2020 (O_2020,N_41308,N_48384);
xnor UO_2021 (O_2021,N_42300,N_49245);
nand UO_2022 (O_2022,N_45384,N_48244);
nand UO_2023 (O_2023,N_47496,N_48346);
nor UO_2024 (O_2024,N_49541,N_44643);
nor UO_2025 (O_2025,N_47144,N_44570);
nor UO_2026 (O_2026,N_46134,N_44161);
xor UO_2027 (O_2027,N_49494,N_48920);
nor UO_2028 (O_2028,N_46154,N_44637);
and UO_2029 (O_2029,N_43808,N_44557);
nor UO_2030 (O_2030,N_41265,N_44434);
xnor UO_2031 (O_2031,N_47987,N_48395);
nand UO_2032 (O_2032,N_49927,N_47248);
nand UO_2033 (O_2033,N_41902,N_49783);
xor UO_2034 (O_2034,N_46943,N_43379);
nand UO_2035 (O_2035,N_41775,N_40190);
nor UO_2036 (O_2036,N_48958,N_46678);
or UO_2037 (O_2037,N_43327,N_49347);
xnor UO_2038 (O_2038,N_48113,N_43878);
and UO_2039 (O_2039,N_45298,N_45920);
nand UO_2040 (O_2040,N_49028,N_46051);
and UO_2041 (O_2041,N_43987,N_49331);
xnor UO_2042 (O_2042,N_46636,N_43751);
or UO_2043 (O_2043,N_43965,N_40350);
or UO_2044 (O_2044,N_49519,N_42114);
nor UO_2045 (O_2045,N_44656,N_49303);
nand UO_2046 (O_2046,N_41714,N_45727);
nor UO_2047 (O_2047,N_41196,N_40107);
or UO_2048 (O_2048,N_40726,N_47365);
nand UO_2049 (O_2049,N_45725,N_40998);
xnor UO_2050 (O_2050,N_47227,N_49999);
nor UO_2051 (O_2051,N_48350,N_48616);
and UO_2052 (O_2052,N_40875,N_41172);
and UO_2053 (O_2053,N_45229,N_40458);
and UO_2054 (O_2054,N_43383,N_42860);
xnor UO_2055 (O_2055,N_46625,N_45356);
or UO_2056 (O_2056,N_48674,N_44613);
nand UO_2057 (O_2057,N_41895,N_48513);
and UO_2058 (O_2058,N_45210,N_46949);
nor UO_2059 (O_2059,N_44196,N_42331);
nor UO_2060 (O_2060,N_46878,N_45309);
xor UO_2061 (O_2061,N_46152,N_47321);
xor UO_2062 (O_2062,N_43917,N_47256);
or UO_2063 (O_2063,N_41052,N_49535);
nor UO_2064 (O_2064,N_47262,N_42172);
and UO_2065 (O_2065,N_40651,N_48208);
and UO_2066 (O_2066,N_48730,N_47497);
and UO_2067 (O_2067,N_42058,N_47257);
or UO_2068 (O_2068,N_48921,N_45549);
xor UO_2069 (O_2069,N_43118,N_48037);
nand UO_2070 (O_2070,N_47572,N_48284);
and UO_2071 (O_2071,N_40398,N_46284);
xor UO_2072 (O_2072,N_44951,N_40299);
and UO_2073 (O_2073,N_46018,N_49255);
and UO_2074 (O_2074,N_49671,N_49715);
nand UO_2075 (O_2075,N_44572,N_43724);
or UO_2076 (O_2076,N_46396,N_45353);
or UO_2077 (O_2077,N_42336,N_46036);
nor UO_2078 (O_2078,N_42784,N_44336);
and UO_2079 (O_2079,N_45865,N_46011);
nand UO_2080 (O_2080,N_42042,N_43678);
nor UO_2081 (O_2081,N_43768,N_43835);
xor UO_2082 (O_2082,N_40484,N_45740);
nor UO_2083 (O_2083,N_46758,N_49644);
and UO_2084 (O_2084,N_48086,N_49792);
nand UO_2085 (O_2085,N_46607,N_48402);
or UO_2086 (O_2086,N_47718,N_47451);
xnor UO_2087 (O_2087,N_45835,N_49707);
nand UO_2088 (O_2088,N_40368,N_42616);
or UO_2089 (O_2089,N_42003,N_42242);
xor UO_2090 (O_2090,N_49777,N_49828);
or UO_2091 (O_2091,N_47126,N_45512);
nor UO_2092 (O_2092,N_48112,N_40888);
and UO_2093 (O_2093,N_47777,N_40091);
xnor UO_2094 (O_2094,N_44560,N_46491);
xor UO_2095 (O_2095,N_47990,N_40685);
xor UO_2096 (O_2096,N_44210,N_47606);
nor UO_2097 (O_2097,N_47390,N_48987);
or UO_2098 (O_2098,N_44478,N_42025);
nor UO_2099 (O_2099,N_40222,N_48670);
nor UO_2100 (O_2100,N_41322,N_48845);
nor UO_2101 (O_2101,N_40804,N_40830);
nor UO_2102 (O_2102,N_41867,N_49222);
nand UO_2103 (O_2103,N_44420,N_40163);
and UO_2104 (O_2104,N_40084,N_49526);
nand UO_2105 (O_2105,N_48647,N_43643);
xnor UO_2106 (O_2106,N_47551,N_44109);
and UO_2107 (O_2107,N_43925,N_47444);
or UO_2108 (O_2108,N_42103,N_47500);
nor UO_2109 (O_2109,N_40453,N_43101);
xor UO_2110 (O_2110,N_41446,N_42442);
nor UO_2111 (O_2111,N_45266,N_49774);
nand UO_2112 (O_2112,N_40239,N_43824);
nand UO_2113 (O_2113,N_46485,N_41219);
or UO_2114 (O_2114,N_40068,N_47190);
nor UO_2115 (O_2115,N_44372,N_40747);
nor UO_2116 (O_2116,N_45715,N_45331);
and UO_2117 (O_2117,N_42463,N_41991);
nor UO_2118 (O_2118,N_47433,N_42846);
or UO_2119 (O_2119,N_49738,N_43764);
or UO_2120 (O_2120,N_46956,N_42328);
nand UO_2121 (O_2121,N_44093,N_44387);
and UO_2122 (O_2122,N_46880,N_49382);
nor UO_2123 (O_2123,N_42432,N_46354);
xor UO_2124 (O_2124,N_46554,N_44286);
or UO_2125 (O_2125,N_45689,N_41883);
xor UO_2126 (O_2126,N_46705,N_43168);
nor UO_2127 (O_2127,N_43276,N_43633);
and UO_2128 (O_2128,N_44283,N_44946);
xor UO_2129 (O_2129,N_43424,N_45396);
or UO_2130 (O_2130,N_40156,N_49158);
and UO_2131 (O_2131,N_45427,N_45282);
nand UO_2132 (O_2132,N_43213,N_41217);
and UO_2133 (O_2133,N_49992,N_40978);
nor UO_2134 (O_2134,N_42270,N_48860);
nand UO_2135 (O_2135,N_49112,N_43059);
xor UO_2136 (O_2136,N_47151,N_44799);
nor UO_2137 (O_2137,N_48097,N_49084);
and UO_2138 (O_2138,N_43547,N_40123);
or UO_2139 (O_2139,N_41386,N_43672);
nand UO_2140 (O_2140,N_48766,N_47226);
or UO_2141 (O_2141,N_47787,N_40741);
nor UO_2142 (O_2142,N_43997,N_47668);
xor UO_2143 (O_2143,N_42906,N_48767);
xnor UO_2144 (O_2144,N_42933,N_47197);
nand UO_2145 (O_2145,N_49017,N_40472);
xor UO_2146 (O_2146,N_49179,N_44467);
nor UO_2147 (O_2147,N_49728,N_45760);
and UO_2148 (O_2148,N_41970,N_48587);
or UO_2149 (O_2149,N_47007,N_44857);
nand UO_2150 (O_2150,N_48108,N_45645);
nand UO_2151 (O_2151,N_44198,N_40081);
nor UO_2152 (O_2152,N_44219,N_40289);
and UO_2153 (O_2153,N_49322,N_41492);
nor UO_2154 (O_2154,N_41332,N_43239);
nand UO_2155 (O_2155,N_46160,N_48579);
xor UO_2156 (O_2156,N_44745,N_45107);
xnor UO_2157 (O_2157,N_46267,N_45791);
or UO_2158 (O_2158,N_44685,N_40868);
nand UO_2159 (O_2159,N_43684,N_40817);
nand UO_2160 (O_2160,N_40663,N_42326);
nor UO_2161 (O_2161,N_44453,N_41767);
nand UO_2162 (O_2162,N_46544,N_46490);
xor UO_2163 (O_2163,N_41525,N_45905);
xnor UO_2164 (O_2164,N_44495,N_49767);
or UO_2165 (O_2165,N_42305,N_48228);
and UO_2166 (O_2166,N_41718,N_43810);
and UO_2167 (O_2167,N_49597,N_44500);
nor UO_2168 (O_2168,N_46484,N_41478);
xor UO_2169 (O_2169,N_49996,N_43328);
xor UO_2170 (O_2170,N_46375,N_47278);
nand UO_2171 (O_2171,N_43504,N_48419);
and UO_2172 (O_2172,N_47238,N_46924);
or UO_2173 (O_2173,N_47826,N_46172);
or UO_2174 (O_2174,N_41230,N_45563);
nand UO_2175 (O_2175,N_42989,N_43472);
or UO_2176 (O_2176,N_40882,N_49987);
or UO_2177 (O_2177,N_46784,N_49297);
and UO_2178 (O_2178,N_40567,N_41026);
nand UO_2179 (O_2179,N_46569,N_45043);
xnor UO_2180 (O_2180,N_40655,N_40369);
nor UO_2181 (O_2181,N_47561,N_41483);
nor UO_2182 (O_2182,N_47758,N_46258);
nor UO_2183 (O_2183,N_40609,N_45377);
or UO_2184 (O_2184,N_45585,N_45133);
or UO_2185 (O_2185,N_46852,N_41355);
and UO_2186 (O_2186,N_42032,N_47544);
or UO_2187 (O_2187,N_44032,N_45381);
nor UO_2188 (O_2188,N_43961,N_43050);
and UO_2189 (O_2189,N_46547,N_41701);
nor UO_2190 (O_2190,N_47904,N_45640);
xnor UO_2191 (O_2191,N_43657,N_49087);
nor UO_2192 (O_2192,N_41805,N_47634);
xor UO_2193 (O_2193,N_44820,N_44195);
and UO_2194 (O_2194,N_48811,N_49606);
and UO_2195 (O_2195,N_46660,N_46218);
xnor UO_2196 (O_2196,N_42279,N_44835);
nor UO_2197 (O_2197,N_43544,N_42533);
nor UO_2198 (O_2198,N_42051,N_46555);
nand UO_2199 (O_2199,N_41870,N_41567);
and UO_2200 (O_2200,N_42477,N_46963);
nor UO_2201 (O_2201,N_46274,N_41789);
or UO_2202 (O_2202,N_43923,N_41623);
and UO_2203 (O_2203,N_42115,N_42647);
and UO_2204 (O_2204,N_41253,N_41811);
nor UO_2205 (O_2205,N_45763,N_41282);
nor UO_2206 (O_2206,N_47017,N_46062);
nand UO_2207 (O_2207,N_44752,N_43522);
and UO_2208 (O_2208,N_47140,N_45193);
nor UO_2209 (O_2209,N_46825,N_44576);
xor UO_2210 (O_2210,N_44005,N_41574);
nand UO_2211 (O_2211,N_44456,N_46677);
or UO_2212 (O_2212,N_41402,N_45919);
and UO_2213 (O_2213,N_49936,N_41364);
xor UO_2214 (O_2214,N_41197,N_40781);
nand UO_2215 (O_2215,N_48654,N_40202);
nor UO_2216 (O_2216,N_41643,N_40342);
nand UO_2217 (O_2217,N_47644,N_45201);
or UO_2218 (O_2218,N_49932,N_43717);
or UO_2219 (O_2219,N_41390,N_48347);
nor UO_2220 (O_2220,N_44477,N_40564);
or UO_2221 (O_2221,N_44382,N_44123);
and UO_2222 (O_2222,N_40050,N_49595);
nor UO_2223 (O_2223,N_42165,N_41081);
xor UO_2224 (O_2224,N_45007,N_42285);
and UO_2225 (O_2225,N_44715,N_42803);
nand UO_2226 (O_2226,N_44209,N_48409);
or UO_2227 (O_2227,N_49855,N_44612);
xor UO_2228 (O_2228,N_47038,N_42586);
xnor UO_2229 (O_2229,N_45817,N_41470);
and UO_2230 (O_2230,N_48743,N_45955);
or UO_2231 (O_2231,N_44215,N_41115);
or UO_2232 (O_2232,N_46023,N_41453);
nand UO_2233 (O_2233,N_40679,N_44300);
or UO_2234 (O_2234,N_49922,N_42834);
xor UO_2235 (O_2235,N_49868,N_41003);
and UO_2236 (O_2236,N_47137,N_40742);
or UO_2237 (O_2237,N_44208,N_47089);
nor UO_2238 (O_2238,N_45442,N_41321);
xnor UO_2239 (O_2239,N_41318,N_48780);
nand UO_2240 (O_2240,N_47156,N_45797);
nor UO_2241 (O_2241,N_47463,N_47581);
xor UO_2242 (O_2242,N_45456,N_43060);
nand UO_2243 (O_2243,N_44690,N_42691);
nor UO_2244 (O_2244,N_41966,N_42595);
nand UO_2245 (O_2245,N_41073,N_41524);
nand UO_2246 (O_2246,N_49886,N_44252);
and UO_2247 (O_2247,N_41065,N_46871);
nor UO_2248 (O_2248,N_49693,N_42158);
or UO_2249 (O_2249,N_40491,N_46489);
nor UO_2250 (O_2250,N_45385,N_46433);
nand UO_2251 (O_2251,N_47186,N_41143);
or UO_2252 (O_2252,N_44814,N_45186);
nand UO_2253 (O_2253,N_47861,N_48693);
nor UO_2254 (O_2254,N_44670,N_47647);
or UO_2255 (O_2255,N_49784,N_41638);
nor UO_2256 (O_2256,N_43412,N_43531);
nand UO_2257 (O_2257,N_46275,N_45962);
nand UO_2258 (O_2258,N_43355,N_42598);
nor UO_2259 (O_2259,N_46876,N_42975);
nand UO_2260 (O_2260,N_46652,N_49012);
or UO_2261 (O_2261,N_42629,N_46976);
and UO_2262 (O_2262,N_49645,N_44325);
or UO_2263 (O_2263,N_40529,N_44849);
and UO_2264 (O_2264,N_40399,N_45751);
nand UO_2265 (O_2265,N_46849,N_47765);
nor UO_2266 (O_2266,N_41297,N_41198);
xor UO_2267 (O_2267,N_48218,N_45616);
and UO_2268 (O_2268,N_47776,N_45790);
xor UO_2269 (O_2269,N_47683,N_47022);
xor UO_2270 (O_2270,N_42141,N_45803);
or UO_2271 (O_2271,N_46683,N_47981);
nand UO_2272 (O_2272,N_43711,N_45004);
and UO_2273 (O_2273,N_44332,N_40774);
and UO_2274 (O_2274,N_45480,N_48031);
or UO_2275 (O_2275,N_46895,N_41646);
nand UO_2276 (O_2276,N_47418,N_45925);
nand UO_2277 (O_2277,N_49114,N_43356);
xor UO_2278 (O_2278,N_41605,N_44639);
nor UO_2279 (O_2279,N_47148,N_49384);
and UO_2280 (O_2280,N_45894,N_43588);
nand UO_2281 (O_2281,N_41950,N_42486);
xor UO_2282 (O_2282,N_41382,N_49903);
xor UO_2283 (O_2283,N_43516,N_47862);
nor UO_2284 (O_2284,N_49102,N_41681);
nor UO_2285 (O_2285,N_41310,N_48931);
and UO_2286 (O_2286,N_46612,N_44339);
and UO_2287 (O_2287,N_49740,N_47434);
xnor UO_2288 (O_2288,N_40611,N_46194);
nand UO_2289 (O_2289,N_48709,N_40775);
nand UO_2290 (O_2290,N_48233,N_40183);
or UO_2291 (O_2291,N_46937,N_47523);
and UO_2292 (O_2292,N_40250,N_48558);
xnor UO_2293 (O_2293,N_45978,N_48849);
xor UO_2294 (O_2294,N_49575,N_41903);
and UO_2295 (O_2295,N_47773,N_41672);
and UO_2296 (O_2296,N_43384,N_49208);
nor UO_2297 (O_2297,N_44551,N_46117);
and UO_2298 (O_2298,N_40633,N_40258);
or UO_2299 (O_2299,N_43782,N_46903);
and UO_2300 (O_2300,N_44749,N_46970);
nand UO_2301 (O_2301,N_41389,N_40355);
nor UO_2302 (O_2302,N_40357,N_40527);
nor UO_2303 (O_2303,N_40750,N_47749);
xnor UO_2304 (O_2304,N_40349,N_49757);
or UO_2305 (O_2305,N_44750,N_42254);
and UO_2306 (O_2306,N_42887,N_45091);
nor UO_2307 (O_2307,N_41329,N_49962);
nor UO_2308 (O_2308,N_47477,N_47848);
or UO_2309 (O_2309,N_41999,N_45151);
nand UO_2310 (O_2310,N_41420,N_44206);
nor UO_2311 (O_2311,N_47516,N_49251);
nor UO_2312 (O_2312,N_42928,N_48778);
xnor UO_2313 (O_2313,N_42540,N_40009);
nor UO_2314 (O_2314,N_44030,N_43766);
nor UO_2315 (O_2315,N_45555,N_49286);
xor UO_2316 (O_2316,N_47295,N_45344);
nor UO_2317 (O_2317,N_40911,N_45245);
xor UO_2318 (O_2318,N_43077,N_44709);
and UO_2319 (O_2319,N_41847,N_46108);
nand UO_2320 (O_2320,N_43897,N_48905);
nor UO_2321 (O_2321,N_42391,N_42646);
xnor UO_2322 (O_2322,N_41114,N_49794);
xnor UO_2323 (O_2323,N_41212,N_42193);
or UO_2324 (O_2324,N_42812,N_46860);
and UO_2325 (O_2325,N_46870,N_47876);
or UO_2326 (O_2326,N_42200,N_49948);
nand UO_2327 (O_2327,N_45709,N_48238);
nor UO_2328 (O_2328,N_46253,N_42988);
nor UO_2329 (O_2329,N_49364,N_44721);
nand UO_2330 (O_2330,N_47616,N_43262);
nor UO_2331 (O_2331,N_46456,N_41653);
xor UO_2332 (O_2332,N_41551,N_46780);
nor UO_2333 (O_2333,N_45794,N_42283);
and UO_2334 (O_2334,N_47109,N_42016);
or UO_2335 (O_2335,N_40271,N_48843);
xor UO_2336 (O_2336,N_48474,N_49263);
xnor UO_2337 (O_2337,N_43032,N_42680);
xnor UO_2338 (O_2338,N_43214,N_48016);
or UO_2339 (O_2339,N_48433,N_49753);
xnor UO_2340 (O_2340,N_40097,N_41679);
and UO_2341 (O_2341,N_48591,N_46663);
nor UO_2342 (O_2342,N_43100,N_44454);
xor UO_2343 (O_2343,N_47957,N_49743);
or UO_2344 (O_2344,N_41338,N_48077);
nand UO_2345 (O_2345,N_40940,N_44821);
and UO_2346 (O_2346,N_40022,N_47356);
or UO_2347 (O_2347,N_47872,N_46776);
and UO_2348 (O_2348,N_41771,N_46584);
nand UO_2349 (O_2349,N_49221,N_45667);
nand UO_2350 (O_2350,N_49227,N_45736);
nor UO_2351 (O_2351,N_47160,N_45116);
and UO_2352 (O_2352,N_46316,N_46302);
nor UO_2353 (O_2353,N_43009,N_44548);
or UO_2354 (O_2354,N_49415,N_46537);
and UO_2355 (O_2355,N_42566,N_44518);
and UO_2356 (O_2356,N_46179,N_44519);
nor UO_2357 (O_2357,N_45680,N_41933);
and UO_2358 (O_2358,N_43714,N_45053);
or UO_2359 (O_2359,N_43162,N_45685);
nand UO_2360 (O_2360,N_42593,N_45359);
nand UO_2361 (O_2361,N_44362,N_43070);
xnor UO_2362 (O_2362,N_47502,N_42426);
xnor UO_2363 (O_2363,N_47218,N_49512);
and UO_2364 (O_2364,N_44599,N_43305);
or UO_2365 (O_2365,N_49734,N_47283);
nor UO_2366 (O_2366,N_40353,N_45535);
nor UO_2367 (O_2367,N_43002,N_47991);
or UO_2368 (O_2368,N_47928,N_43260);
nand UO_2369 (O_2369,N_48120,N_46801);
xnor UO_2370 (O_2370,N_45028,N_42932);
xnor UO_2371 (O_2371,N_45706,N_44537);
and UO_2372 (O_2372,N_41239,N_42766);
and UO_2373 (O_2373,N_45524,N_40428);
xnor UO_2374 (O_2374,N_46330,N_46174);
nor UO_2375 (O_2375,N_43632,N_44607);
and UO_2376 (O_2376,N_47162,N_42241);
nand UO_2377 (O_2377,N_45048,N_46366);
or UO_2378 (O_2378,N_47347,N_43577);
nand UO_2379 (O_2379,N_45679,N_47640);
or UO_2380 (O_2380,N_44846,N_46686);
nand UO_2381 (O_2381,N_49862,N_44302);
and UO_2382 (O_2382,N_48967,N_48810);
nor UO_2383 (O_2383,N_48926,N_44890);
and UO_2384 (O_2384,N_43474,N_48655);
nor UO_2385 (O_2385,N_46646,N_46070);
or UO_2386 (O_2386,N_45711,N_41854);
or UO_2387 (O_2387,N_48636,N_43485);
xor UO_2388 (O_2388,N_41315,N_49599);
nand UO_2389 (O_2389,N_49033,N_46851);
nor UO_2390 (O_2390,N_42785,N_42840);
or UO_2391 (O_2391,N_47116,N_43454);
nand UO_2392 (O_2392,N_42231,N_47319);
nand UO_2393 (O_2393,N_44484,N_40751);
nor UO_2394 (O_2394,N_45445,N_43759);
or UO_2395 (O_2395,N_41257,N_48898);
nor UO_2396 (O_2396,N_44808,N_46985);
or UO_2397 (O_2397,N_45948,N_47432);
xor UO_2398 (O_2398,N_44317,N_42050);
nor UO_2399 (O_2399,N_42908,N_45664);
nor UO_2400 (O_2400,N_41542,N_49818);
or UO_2401 (O_2401,N_47711,N_46599);
or UO_2402 (O_2402,N_43121,N_46938);
and UO_2403 (O_2403,N_49239,N_42603);
nand UO_2404 (O_2404,N_48607,N_48336);
nand UO_2405 (O_2405,N_42309,N_46588);
nand UO_2406 (O_2406,N_42056,N_44829);
and UO_2407 (O_2407,N_40960,N_43181);
nand UO_2408 (O_2408,N_48357,N_45728);
or UO_2409 (O_2409,N_47215,N_41750);
xor UO_2410 (O_2410,N_48733,N_49150);
and UO_2411 (O_2411,N_41818,N_40832);
or UO_2412 (O_2412,N_49462,N_43192);
or UO_2413 (O_2413,N_46681,N_42706);
or UO_2414 (O_2414,N_49177,N_43710);
or UO_2415 (O_2415,N_43656,N_45674);
xor UO_2416 (O_2416,N_46952,N_40083);
nor UO_2417 (O_2417,N_42181,N_42027);
and UO_2418 (O_2418,N_47527,N_44985);
xor UO_2419 (O_2419,N_42410,N_44352);
nand UO_2420 (O_2420,N_48020,N_41555);
xnor UO_2421 (O_2421,N_42320,N_42479);
or UO_2422 (O_2422,N_43936,N_47779);
or UO_2423 (O_2423,N_45829,N_45964);
nand UO_2424 (O_2424,N_44164,N_49049);
or UO_2425 (O_2425,N_48874,N_48463);
and UO_2426 (O_2426,N_49183,N_42601);
and UO_2427 (O_2427,N_42743,N_45898);
or UO_2428 (O_2428,N_46883,N_45464);
nor UO_2429 (O_2429,N_44223,N_45198);
or UO_2430 (O_2430,N_41719,N_44400);
nor UO_2431 (O_2431,N_47346,N_43957);
or UO_2432 (O_2432,N_45969,N_41398);
nor UO_2433 (O_2433,N_40930,N_43887);
or UO_2434 (O_2434,N_45682,N_48566);
nand UO_2435 (O_2435,N_45013,N_49518);
nor UO_2436 (O_2436,N_49985,N_46528);
or UO_2437 (O_2437,N_42221,N_41075);
nand UO_2438 (O_2438,N_41497,N_46627);
and UO_2439 (O_2439,N_42980,N_48943);
nor UO_2440 (O_2440,N_45345,N_47306);
and UO_2441 (O_2441,N_43856,N_41849);
xnor UO_2442 (O_2442,N_49723,N_43246);
nor UO_2443 (O_2443,N_46916,N_42291);
nand UO_2444 (O_2444,N_48932,N_48122);
or UO_2445 (O_2445,N_42201,N_41436);
xor UO_2446 (O_2446,N_46731,N_41856);
and UO_2447 (O_2447,N_48526,N_46183);
or UO_2448 (O_2448,N_42190,N_46355);
nand UO_2449 (O_2449,N_46608,N_41973);
or UO_2450 (O_2450,N_47925,N_48364);
nand UO_2451 (O_2451,N_41330,N_48903);
or UO_2452 (O_2452,N_42833,N_42607);
or UO_2453 (O_2453,N_49220,N_49001);
or UO_2454 (O_2454,N_42445,N_41637);
nor UO_2455 (O_2455,N_42978,N_45161);
nand UO_2456 (O_2456,N_40502,N_46312);
nor UO_2457 (O_2457,N_42356,N_47931);
nor UO_2458 (O_2458,N_47460,N_47700);
or UO_2459 (O_2459,N_45475,N_48129);
or UO_2460 (O_2460,N_45973,N_47564);
and UO_2461 (O_2461,N_45380,N_43423);
xnor UO_2462 (O_2462,N_49487,N_47427);
or UO_2463 (O_2463,N_42232,N_46623);
or UO_2464 (O_2464,N_41896,N_43568);
or UO_2465 (O_2465,N_42911,N_40600);
nor UO_2466 (O_2466,N_41079,N_49708);
nor UO_2467 (O_2467,N_45086,N_47291);
or UO_2468 (O_2468,N_40637,N_49223);
nor UO_2469 (O_2469,N_49290,N_43831);
or UO_2470 (O_2470,N_44960,N_45644);
or UO_2471 (O_2471,N_45773,N_47010);
nand UO_2472 (O_2472,N_47387,N_41583);
xnor UO_2473 (O_2473,N_49506,N_49566);
nor UO_2474 (O_2474,N_49356,N_42651);
and UO_2475 (O_2475,N_45502,N_43261);
or UO_2476 (O_2476,N_46918,N_48272);
and UO_2477 (O_2477,N_42288,N_41371);
nand UO_2478 (O_2478,N_48961,N_42453);
nor UO_2479 (O_2479,N_47817,N_42180);
and UO_2480 (O_2480,N_48437,N_47650);
nand UO_2481 (O_2481,N_44046,N_40517);
xor UO_2482 (O_2482,N_42009,N_43513);
xor UO_2483 (O_2483,N_45347,N_49216);
nor UO_2484 (O_2484,N_44221,N_44614);
nor UO_2485 (O_2485,N_41698,N_45470);
nor UO_2486 (O_2486,N_44785,N_40690);
and UO_2487 (O_2487,N_40584,N_47624);
nand UO_2488 (O_2488,N_44653,N_40333);
nor UO_2489 (O_2489,N_45820,N_44693);
and UO_2490 (O_2490,N_42182,N_41059);
and UO_2491 (O_2491,N_44406,N_40964);
xnor UO_2492 (O_2492,N_43863,N_46224);
xnor UO_2493 (O_2493,N_48606,N_40628);
nor UO_2494 (O_2494,N_40391,N_46125);
xnor UO_2495 (O_2495,N_44095,N_45714);
or UO_2496 (O_2496,N_43565,N_49653);
nor UO_2497 (O_2497,N_43829,N_43201);
nand UO_2498 (O_2498,N_46600,N_43018);
xnor UO_2499 (O_2499,N_49630,N_43557);
and UO_2500 (O_2500,N_49775,N_48893);
nand UO_2501 (O_2501,N_43884,N_43761);
xnor UO_2502 (O_2502,N_41353,N_49570);
nand UO_2503 (O_2503,N_48176,N_41291);
nand UO_2504 (O_2504,N_42203,N_49816);
or UO_2505 (O_2505,N_47903,N_44440);
nor UO_2506 (O_2506,N_49659,N_47464);
nand UO_2507 (O_2507,N_42941,N_42420);
xnor UO_2508 (O_2508,N_40224,N_43430);
and UO_2509 (O_2509,N_40623,N_40108);
or UO_2510 (O_2510,N_48996,N_42072);
xor UO_2511 (O_2511,N_40117,N_43390);
nand UO_2512 (O_2512,N_46419,N_45618);
nand UO_2513 (O_2513,N_48671,N_44538);
nand UO_2514 (O_2514,N_42213,N_42606);
and UO_2515 (O_2515,N_40322,N_41138);
or UO_2516 (O_2516,N_48540,N_40986);
xor UO_2517 (O_2517,N_48924,N_48396);
and UO_2518 (O_2518,N_48339,N_40699);
xnor UO_2519 (O_2519,N_40063,N_43681);
and UO_2520 (O_2520,N_44333,N_42570);
nand UO_2521 (O_2521,N_43543,N_40808);
nand UO_2522 (O_2522,N_44261,N_49558);
xnor UO_2523 (O_2523,N_40192,N_42851);
nor UO_2524 (O_2524,N_44966,N_41189);
or UO_2525 (O_2525,N_43780,N_45424);
nor UO_2526 (O_2526,N_44308,N_41451);
nand UO_2527 (O_2527,N_40308,N_43029);
xor UO_2528 (O_2528,N_41087,N_47736);
nand UO_2529 (O_2529,N_40060,N_45627);
xnor UO_2530 (O_2530,N_49072,N_45473);
xnor UO_2531 (O_2531,N_41748,N_43832);
xor UO_2532 (O_2532,N_47943,N_44680);
xnor UO_2533 (O_2533,N_49253,N_45731);
nor UO_2534 (O_2534,N_41300,N_40957);
nor UO_2535 (O_2535,N_47426,N_42814);
xnor UO_2536 (O_2536,N_43750,N_40806);
xor UO_2537 (O_2537,N_40732,N_40427);
nor UO_2538 (O_2538,N_45816,N_46282);
and UO_2539 (O_2539,N_48049,N_47235);
nand UO_2540 (O_2540,N_47822,N_40952);
and UO_2541 (O_2541,N_46662,N_44050);
nor UO_2542 (O_2542,N_48590,N_45174);
xnor UO_2543 (O_2543,N_44893,N_42461);
or UO_2544 (O_2544,N_43166,N_49786);
and UO_2545 (O_2545,N_40347,N_42481);
nand UO_2546 (O_2546,N_45449,N_42371);
nand UO_2547 (O_2547,N_49991,N_43712);
xor UO_2548 (O_2548,N_43263,N_43951);
nor UO_2549 (O_2549,N_47538,N_40270);
or UO_2550 (O_2550,N_42383,N_49315);
and UO_2551 (O_2551,N_49270,N_49449);
or UO_2552 (O_2552,N_49039,N_49194);
or UO_2553 (O_2553,N_44995,N_43990);
nor UO_2554 (O_2554,N_49383,N_43291);
xor UO_2555 (O_2555,N_46695,N_45327);
nor UO_2556 (O_2556,N_48449,N_49176);
or UO_2557 (O_2557,N_46651,N_47074);
and UO_2558 (O_2558,N_41840,N_49831);
and UO_2559 (O_2559,N_48725,N_47598);
nand UO_2560 (O_2560,N_45191,N_45860);
and UO_2561 (O_2561,N_47183,N_48054);
nand UO_2562 (O_2562,N_45110,N_42948);
and UO_2563 (O_2563,N_40328,N_49890);
or UO_2564 (O_2564,N_47132,N_49070);
and UO_2565 (O_2565,N_49178,N_40530);
nand UO_2566 (O_2566,N_45610,N_47121);
xnor UO_2567 (O_2567,N_45306,N_42126);
xor UO_2568 (O_2568,N_43791,N_43204);
or UO_2569 (O_2569,N_47970,N_40277);
nor UO_2570 (O_2570,N_44633,N_46813);
and UO_2571 (O_2571,N_45737,N_44086);
nor UO_2572 (O_2572,N_43347,N_46408);
or UO_2573 (O_2573,N_49812,N_48732);
or UO_2574 (O_2574,N_40936,N_44401);
or UO_2575 (O_2575,N_49419,N_41564);
xnor UO_2576 (O_2576,N_43266,N_43852);
nor UO_2577 (O_2577,N_49489,N_47441);
xnor UO_2578 (O_2578,N_45719,N_46038);
xnor UO_2579 (O_2579,N_44145,N_45230);
or UO_2580 (O_2580,N_48450,N_44007);
nand UO_2581 (O_2581,N_45244,N_44834);
xnor UO_2582 (O_2582,N_49131,N_49037);
and UO_2583 (O_2583,N_41107,N_43520);
nor UO_2584 (O_2584,N_46111,N_42227);
or UO_2585 (O_2585,N_42327,N_40857);
and UO_2586 (O_2586,N_47639,N_43933);
nor UO_2587 (O_2587,N_45143,N_42913);
and UO_2588 (O_2588,N_48776,N_41091);
nand UO_2589 (O_2589,N_41397,N_43709);
and UO_2590 (O_2590,N_40312,N_47133);
nand UO_2591 (O_2591,N_41360,N_45697);
nor UO_2592 (O_2592,N_44485,N_41753);
nor UO_2593 (O_2593,N_40495,N_46703);
or UO_2594 (O_2594,N_49199,N_44114);
nand UO_2595 (O_2595,N_41509,N_41518);
or UO_2596 (O_2596,N_40896,N_42959);
xnor UO_2597 (O_2597,N_45636,N_42396);
nand UO_2598 (O_2598,N_43935,N_49181);
xor UO_2599 (O_2599,N_41724,N_43603);
nor UO_2600 (O_2600,N_48034,N_49964);
nand UO_2601 (O_2601,N_44374,N_45994);
xnor UO_2602 (O_2602,N_40094,N_42632);
or UO_2603 (O_2603,N_49785,N_44299);
xnor UO_2604 (O_2604,N_48736,N_48421);
and UO_2605 (O_2605,N_46289,N_48481);
nand UO_2606 (O_2606,N_49758,N_45250);
nand UO_2607 (O_2607,N_43405,N_44514);
nor UO_2608 (O_2608,N_41002,N_49349);
and UO_2609 (O_2609,N_41837,N_42052);
or UO_2610 (O_2610,N_44955,N_49633);
and UO_2611 (O_2611,N_43903,N_43099);
nand UO_2612 (O_2612,N_47996,N_47786);
or UO_2613 (O_2613,N_47228,N_43584);
xnor UO_2614 (O_2614,N_46854,N_42282);
xnor UO_2615 (O_2615,N_42266,N_43876);
xor UO_2616 (O_2616,N_45999,N_45926);
and UO_2617 (O_2617,N_44493,N_43536);
or UO_2618 (O_2618,N_44120,N_46392);
and UO_2619 (O_2619,N_48098,N_49403);
nand UO_2620 (O_2620,N_47223,N_47508);
nor UO_2621 (O_2621,N_44065,N_42709);
nand UO_2622 (O_2622,N_42663,N_46987);
nand UO_2623 (O_2623,N_46535,N_45469);
xor UO_2624 (O_2624,N_41279,N_42397);
and UO_2625 (O_2625,N_46747,N_47824);
xor UO_2626 (O_2626,N_43674,N_44969);
xor UO_2627 (O_2627,N_47619,N_40660);
and UO_2628 (O_2628,N_40489,N_48509);
nand UO_2629 (O_2629,N_45297,N_47850);
nand UO_2630 (O_2630,N_41932,N_46567);
nor UO_2631 (O_2631,N_44422,N_41225);
xnor UO_2632 (O_2632,N_47343,N_41223);
nand UO_2633 (O_2633,N_44131,N_47023);
nor UO_2634 (O_2634,N_47296,N_43578);
xor UO_2635 (O_2635,N_40538,N_48101);
nand UO_2636 (O_2636,N_48942,N_40723);
or UO_2637 (O_2637,N_49300,N_48809);
nand UO_2638 (O_2638,N_40669,N_42454);
and UO_2639 (O_2639,N_47701,N_46219);
or UO_2640 (O_2640,N_44168,N_48440);
or UO_2641 (O_2641,N_43446,N_44075);
and UO_2642 (O_2642,N_45468,N_44906);
and UO_2643 (O_2643,N_47873,N_42013);
nand UO_2644 (O_2644,N_49287,N_45369);
and UO_2645 (O_2645,N_49934,N_41639);
and UO_2646 (O_2646,N_49596,N_49256);
and UO_2647 (O_2647,N_47556,N_43877);
nand UO_2648 (O_2648,N_49843,N_43533);
xnor UO_2649 (O_2649,N_41782,N_41369);
nand UO_2650 (O_2650,N_44483,N_44772);
nand UO_2651 (O_2651,N_44564,N_45771);
nor UO_2652 (O_2652,N_49817,N_44944);
xor UO_2653 (O_2653,N_45518,N_40814);
nor UO_2654 (O_2654,N_47895,N_42404);
nor UO_2655 (O_2655,N_43506,N_45472);
nand UO_2656 (O_2656,N_44057,N_40144);
nor UO_2657 (O_2657,N_40730,N_41037);
nand UO_2658 (O_2658,N_40151,N_47920);
or UO_2659 (O_2659,N_43706,N_43691);
nor UO_2660 (O_2660,N_46603,N_48274);
xnor UO_2661 (O_2661,N_45495,N_44632);
xnor UO_2662 (O_2662,N_49345,N_41951);
and UO_2663 (O_2663,N_43448,N_48562);
xor UO_2664 (O_2664,N_45800,N_40177);
nand UO_2665 (O_2665,N_44577,N_41439);
xor UO_2666 (O_2666,N_49371,N_44781);
xor UO_2667 (O_2667,N_40516,N_48255);
nor UO_2668 (O_2668,N_45108,N_48236);
and UO_2669 (O_2669,N_41594,N_45633);
or UO_2670 (O_2670,N_49075,N_44509);
and UO_2671 (O_2671,N_43007,N_42550);
xor UO_2672 (O_2672,N_45249,N_43256);
xnor UO_2673 (O_2673,N_49854,N_47637);
and UO_2674 (O_2674,N_40100,N_48791);
xor UO_2675 (O_2675,N_44836,N_44212);
nand UO_2676 (O_2676,N_45218,N_43794);
and UO_2677 (O_2677,N_49898,N_42874);
nor UO_2678 (O_2678,N_41133,N_42938);
xnor UO_2679 (O_2679,N_45721,N_45594);
nor UO_2680 (O_2680,N_49234,N_47332);
and UO_2681 (O_2681,N_49202,N_44391);
and UO_2682 (O_2682,N_45124,N_46362);
xnor UO_2683 (O_2683,N_48050,N_48355);
xnor UO_2684 (O_2684,N_49641,N_46406);
or UO_2685 (O_2685,N_49431,N_40044);
and UO_2686 (O_2686,N_41828,N_45796);
nand UO_2687 (O_2687,N_49461,N_48140);
xnor UO_2688 (O_2688,N_47495,N_49203);
or UO_2689 (O_2689,N_41335,N_44917);
nand UO_2690 (O_2690,N_41214,N_45069);
nand UO_2691 (O_2691,N_49230,N_40734);
nand UO_2692 (O_2692,N_43971,N_48764);
xnor UO_2693 (O_2693,N_46822,N_48162);
nand UO_2694 (O_2694,N_41640,N_43233);
xnor UO_2695 (O_2695,N_41510,N_44166);
nand UO_2696 (O_2696,N_43183,N_45097);
nor UO_2697 (O_2697,N_44668,N_41813);
xor UO_2698 (O_2698,N_40641,N_48211);
nor UO_2699 (O_2699,N_43934,N_43611);
nand UO_2700 (O_2700,N_43613,N_43579);
xor UO_2701 (O_2701,N_46445,N_48543);
nor UO_2702 (O_2702,N_43991,N_49533);
and UO_2703 (O_2703,N_48473,N_45930);
nor UO_2704 (O_2704,N_43732,N_45491);
or UO_2705 (O_2705,N_44138,N_41661);
and UO_2706 (O_2706,N_44229,N_40841);
xnor UO_2707 (O_2707,N_43600,N_49104);
nor UO_2708 (O_2708,N_42044,N_49231);
and UO_2709 (O_2709,N_49138,N_48611);
or UO_2710 (O_2710,N_46225,N_42865);
or UO_2711 (O_2711,N_45374,N_42437);
xnor UO_2712 (O_2712,N_45945,N_43470);
nand UO_2713 (O_2713,N_40748,N_46055);
nor UO_2714 (O_2714,N_49478,N_40339);
and UO_2715 (O_2715,N_46696,N_42353);
and UO_2716 (O_2716,N_41122,N_47618);
xnor UO_2717 (O_2717,N_49751,N_45691);
nand UO_2718 (O_2718,N_40345,N_41955);
xnor UO_2719 (O_2719,N_42229,N_40671);
and UO_2720 (O_2720,N_41794,N_45348);
xnor UO_2721 (O_2721,N_49373,N_43738);
nand UO_2722 (O_2722,N_41227,N_48133);
xor UO_2723 (O_2723,N_42000,N_45001);
nand UO_2724 (O_2724,N_43012,N_43058);
nand UO_2725 (O_2725,N_46103,N_44036);
nor UO_2726 (O_2726,N_40325,N_41731);
nor UO_2727 (O_2727,N_45622,N_40477);
nor UO_2728 (O_2728,N_48622,N_45318);
or UO_2729 (O_2729,N_43081,N_43016);
nor UO_2730 (O_2730,N_41930,N_47442);
xor UO_2731 (O_2731,N_41488,N_47063);
xnor UO_2732 (O_2732,N_41441,N_41005);
xor UO_2733 (O_2733,N_41105,N_48643);
nor UO_2734 (O_2734,N_45052,N_42984);
nor UO_2735 (O_2735,N_46165,N_49610);
and UO_2736 (O_2736,N_43676,N_47866);
or UO_2737 (O_2737,N_44719,N_42091);
nor UO_2738 (O_2738,N_48883,N_40023);
nand UO_2739 (O_2739,N_43011,N_48863);
xor UO_2740 (O_2740,N_47916,N_46141);
and UO_2741 (O_2741,N_43304,N_42155);
or UO_2742 (O_2742,N_44184,N_42011);
xnor UO_2743 (O_2743,N_43313,N_43820);
or UO_2744 (O_2744,N_44665,N_42143);
and UO_2745 (O_2745,N_49008,N_42794);
xor UO_2746 (O_2746,N_45710,N_42799);
and UO_2747 (O_2747,N_42263,N_44650);
and UO_2748 (O_2748,N_48069,N_42330);
and UO_2749 (O_2749,N_49409,N_42901);
xor UO_2750 (O_2750,N_49950,N_48826);
nor UO_2751 (O_2751,N_46941,N_45383);
and UO_2752 (O_2752,N_49531,N_41723);
and UO_2753 (O_2753,N_44010,N_48100);
nor UO_2754 (O_2754,N_44482,N_45908);
or UO_2755 (O_2755,N_46426,N_47932);
nand UO_2756 (O_2756,N_44249,N_47750);
xnor UO_2757 (O_2757,N_40601,N_42120);
nor UO_2758 (O_2758,N_49135,N_43505);
xnor UO_2759 (O_2759,N_42162,N_48280);
or UO_2760 (O_2760,N_43309,N_44903);
xnor UO_2761 (O_2761,N_48758,N_44083);
nand UO_2762 (O_2762,N_40552,N_47483);
xnor UO_2763 (O_2763,N_42095,N_45944);
and UO_2764 (O_2764,N_43125,N_45520);
nor UO_2765 (O_2765,N_40090,N_49998);
nor UO_2766 (O_2766,N_42487,N_47614);
nor UO_2767 (O_2767,N_47161,N_48381);
nor UO_2768 (O_2768,N_49574,N_43940);
or UO_2769 (O_2769,N_48445,N_44237);
and UO_2770 (O_2770,N_40731,N_42024);
or UO_2771 (O_2771,N_49453,N_48192);
nor UO_2772 (O_2772,N_47455,N_44421);
nor UO_2773 (O_2773,N_42699,N_42034);
xor UO_2774 (O_2774,N_45830,N_44513);
nor UO_2775 (O_2775,N_42197,N_43199);
nor UO_2776 (O_2776,N_46326,N_40917);
and UO_2777 (O_2777,N_47323,N_42756);
or UO_2778 (O_2778,N_40301,N_41136);
or UO_2779 (O_2779,N_41503,N_41815);
xnor UO_2780 (O_2780,N_47537,N_48491);
and UO_2781 (O_2781,N_46610,N_43625);
nor UO_2782 (O_2782,N_42714,N_44567);
xor UO_2783 (O_2783,N_43165,N_46538);
nor UO_2784 (O_2784,N_42692,N_48165);
nand UO_2785 (O_2785,N_41468,N_49678);
nand UO_2786 (O_2786,N_41953,N_45251);
and UO_2787 (O_2787,N_40547,N_48729);
nand UO_2788 (O_2788,N_41401,N_49118);
and UO_2789 (O_2789,N_42551,N_48834);
nand UO_2790 (O_2790,N_40684,N_48323);
nand UO_2791 (O_2791,N_49307,N_46733);
nand UO_2792 (O_2792,N_41801,N_49106);
xor UO_2793 (O_2793,N_49281,N_40602);
or UO_2794 (O_2794,N_45943,N_41915);
nor UO_2795 (O_2795,N_47919,N_49939);
nor UO_2796 (O_2796,N_42961,N_41851);
xor UO_2797 (O_2797,N_46222,N_48296);
nor UO_2798 (O_2798,N_41888,N_45202);
or UO_2799 (O_2799,N_42490,N_42515);
or UO_2800 (O_2800,N_45921,N_45137);
or UO_2801 (O_2801,N_46346,N_44190);
nor UO_2802 (O_2802,N_40026,N_44099);
nand UO_2803 (O_2803,N_47585,N_40092);
nor UO_2804 (O_2804,N_41350,N_44646);
nand UO_2805 (O_2805,N_49499,N_46293);
and UO_2806 (O_2806,N_45849,N_45262);
nand UO_2807 (O_2807,N_42195,N_49252);
or UO_2808 (O_2808,N_48047,N_48042);
xnor UO_2809 (O_2809,N_40657,N_40634);
and UO_2810 (O_2810,N_49911,N_44541);
or UO_2811 (O_2811,N_45419,N_44932);
nand UO_2812 (O_2812,N_41561,N_40167);
and UO_2813 (O_2813,N_46098,N_46846);
nand UO_2814 (O_2814,N_46262,N_44686);
or UO_2815 (O_2815,N_45338,N_44943);
nor UO_2816 (O_2816,N_40082,N_46531);
nand UO_2817 (O_2817,N_44307,N_46768);
nor UO_2818 (O_2818,N_46335,N_48510);
or UO_2819 (O_2819,N_42853,N_49292);
nand UO_2820 (O_2820,N_47760,N_44346);
xnor UO_2821 (O_2821,N_41430,N_46858);
xor UO_2822 (O_2822,N_43998,N_47084);
and UO_2823 (O_2823,N_40370,N_47044);
nand UO_2824 (O_2824,N_44671,N_43772);
and UO_2825 (O_2825,N_44089,N_46777);
nor UO_2826 (O_2826,N_49623,N_46821);
xnor UO_2827 (O_2827,N_43735,N_42497);
and UO_2828 (O_2828,N_43982,N_45221);
nand UO_2829 (O_2829,N_49397,N_46840);
and UO_2830 (O_2830,N_43367,N_42206);
and UO_2831 (O_2831,N_43660,N_48166);
and UO_2832 (O_2832,N_41032,N_49468);
xnor UO_2833 (O_2833,N_49584,N_43408);
xnor UO_2834 (O_2834,N_41634,N_47320);
nor UO_2835 (O_2835,N_44239,N_43668);
or UO_2836 (O_2836,N_48490,N_41755);
xnor UO_2837 (O_2837,N_47034,N_47570);
and UO_2838 (O_2838,N_40011,N_42545);
xor UO_2839 (O_2839,N_45641,N_49200);
nor UO_2840 (O_2840,N_40849,N_41622);
xor UO_2841 (O_2841,N_47936,N_45545);
and UO_2842 (O_2842,N_44900,N_48995);
xnor UO_2843 (O_2843,N_44764,N_44175);
nor UO_2844 (O_2844,N_47204,N_44323);
or UO_2845 (O_2845,N_42547,N_43037);
or UO_2846 (O_2846,N_46271,N_43995);
or UO_2847 (O_2847,N_44534,N_41773);
and UO_2848 (O_2848,N_46203,N_41781);
xor UO_2849 (O_2849,N_48436,N_45407);
and UO_2850 (O_2850,N_48106,N_49745);
nand UO_2851 (O_2851,N_48792,N_40945);
nor UO_2852 (O_2852,N_43652,N_48182);
xor UO_2853 (O_2853,N_47783,N_48550);
xnor UO_2854 (O_2854,N_42968,N_42088);
nand UO_2855 (O_2855,N_42067,N_48605);
and UO_2856 (O_2856,N_47243,N_42375);
and UO_2857 (O_2857,N_43228,N_43219);
nor UO_2858 (O_2858,N_40926,N_40382);
nor UO_2859 (O_2859,N_45126,N_42379);
nor UO_2860 (O_2860,N_43417,N_46900);
xor UO_2861 (O_2861,N_46719,N_49586);
and UO_2862 (O_2862,N_47686,N_45263);
nor UO_2863 (O_2863,N_41570,N_48723);
xor UO_2864 (O_2864,N_42362,N_40046);
nand UO_2865 (O_2865,N_45070,N_46080);
nand UO_2866 (O_2866,N_48065,N_45149);
or UO_2867 (O_2867,N_42742,N_46619);
nor UO_2868 (O_2868,N_41797,N_47998);
nor UO_2869 (O_2869,N_47423,N_41414);
nand UO_2870 (O_2870,N_41443,N_47198);
and UO_2871 (O_2871,N_40356,N_48639);
nand UO_2872 (O_2872,N_48310,N_49280);
nor UO_2873 (O_2873,N_45365,N_41296);
and UO_2874 (O_2874,N_43102,N_45844);
xor UO_2875 (O_2875,N_46112,N_43469);
nand UO_2876 (O_2876,N_44540,N_43702);
or UO_2877 (O_2877,N_42361,N_46583);
and UO_2878 (O_2878,N_48517,N_47836);
nand UO_2879 (O_2879,N_48264,N_41500);
xor UO_2880 (O_2880,N_48278,N_42359);
and UO_2881 (O_2881,N_44371,N_48572);
and UO_2882 (O_2882,N_46614,N_46382);
nand UO_2883 (O_2883,N_43451,N_45051);
and UO_2884 (O_2884,N_41031,N_40979);
nor UO_2885 (O_2885,N_45483,N_48263);
and UO_2886 (O_2886,N_40159,N_48114);
nand UO_2887 (O_2887,N_48007,N_45364);
xnor UO_2888 (O_2888,N_43130,N_42954);
and UO_2889 (O_2889,N_47330,N_48904);
nor UO_2890 (O_2890,N_43088,N_40110);
nand UO_2891 (O_2891,N_47307,N_42144);
nor UO_2892 (O_2892,N_41936,N_46472);
and UO_2893 (O_2893,N_45199,N_47005);
or UO_2894 (O_2894,N_46645,N_43806);
and UO_2895 (O_2895,N_41504,N_46644);
and UO_2896 (O_2896,N_44197,N_49877);
xnor UO_2897 (O_2897,N_46017,N_46805);
or UO_2898 (O_2898,N_45783,N_41201);
nor UO_2899 (O_2899,N_42273,N_48703);
nand UO_2900 (O_2900,N_42520,N_42469);
or UO_2901 (O_2901,N_44910,N_45215);
nand UO_2902 (O_2902,N_40565,N_45059);
or UO_2903 (O_2903,N_47178,N_45742);
or UO_2904 (O_2904,N_48216,N_45062);
or UO_2905 (O_2905,N_42622,N_42544);
nor UO_2906 (O_2906,N_48844,N_43589);
and UO_2907 (O_2907,N_47714,N_46414);
nor UO_2908 (O_2908,N_48253,N_41396);
xor UO_2909 (O_2909,N_45779,N_42866);
and UO_2910 (O_2910,N_46609,N_43954);
and UO_2911 (O_2911,N_46229,N_40735);
nand UO_2912 (O_2912,N_48518,N_43456);
xor UO_2913 (O_2913,N_48001,N_42390);
or UO_2914 (O_2914,N_41572,N_42194);
nand UO_2915 (O_2915,N_44695,N_47665);
nor UO_2916 (O_2916,N_43482,N_46436);
nand UO_2917 (O_2917,N_47003,N_41635);
or UO_2918 (O_2918,N_44630,N_47726);
nor UO_2919 (O_2919,N_41543,N_44125);
xnor UO_2920 (O_2920,N_41920,N_49808);
or UO_2921 (O_2921,N_44446,N_40384);
nor UO_2922 (O_2922,N_47770,N_40761);
and UO_2923 (O_2923,N_40629,N_49271);
xor UO_2924 (O_2924,N_46119,N_45378);
nor UO_2925 (O_2925,N_41879,N_48589);
or UO_2926 (O_2926,N_45246,N_49484);
and UO_2927 (O_2927,N_47011,N_41388);
or UO_2928 (O_2928,N_48837,N_41855);
or UO_2929 (O_2929,N_48335,N_49086);
xor UO_2930 (O_2930,N_45718,N_42064);
xnor UO_2931 (O_2931,N_44916,N_48226);
xnor UO_2932 (O_2932,N_43827,N_42082);
and UO_2933 (O_2933,N_41763,N_44381);
nand UO_2934 (O_2934,N_44904,N_48152);
and UO_2935 (O_2935,N_49975,N_40551);
and UO_2936 (O_2936,N_48857,N_47751);
or UO_2937 (O_2937,N_40931,N_42435);
or UO_2938 (O_2938,N_45431,N_45337);
xnor UO_2939 (O_2939,N_44638,N_40273);
nor UO_2940 (O_2940,N_43719,N_47388);
nor UO_2941 (O_2941,N_43662,N_48279);
and UO_2942 (O_2942,N_40430,N_42061);
or UO_2943 (O_2943,N_40778,N_47881);
or UO_2944 (O_2944,N_44627,N_46075);
xor UO_2945 (O_2945,N_47035,N_46238);
and UO_2946 (O_2946,N_47973,N_46891);
xor UO_2947 (O_2947,N_46058,N_44651);
or UO_2948 (O_2948,N_45883,N_41686);
and UO_2949 (O_2949,N_46931,N_48358);
nand UO_2950 (O_2950,N_44244,N_41112);
nor UO_2951 (O_2951,N_43535,N_48751);
and UO_2952 (O_2952,N_43861,N_45889);
and UO_2953 (O_2953,N_48205,N_45972);
or UO_2954 (O_2954,N_40913,N_42875);
nand UO_2955 (O_2955,N_45239,N_45632);
or UO_2956 (O_2956,N_41998,N_48929);
xnor UO_2957 (O_2957,N_42549,N_48167);
xnor UO_2958 (O_2958,N_45315,N_45453);
and UO_2959 (O_2959,N_48656,N_40953);
xnor UO_2960 (O_2960,N_41559,N_43664);
nand UO_2961 (O_2961,N_46339,N_40407);
or UO_2962 (O_2962,N_47853,N_42672);
or UO_2963 (O_2963,N_49607,N_45552);
and UO_2964 (O_2964,N_48241,N_45734);
nand UO_2965 (O_2965,N_49034,N_47420);
or UO_2966 (O_2966,N_44989,N_46081);
or UO_2967 (O_2967,N_40786,N_43955);
nor UO_2968 (O_2968,N_49492,N_44802);
xnor UO_2969 (O_2969,N_43108,N_40773);
or UO_2970 (O_2970,N_44705,N_43447);
xnor UO_2971 (O_2971,N_42872,N_42777);
nand UO_2972 (O_2972,N_45838,N_47555);
nor UO_2973 (O_2973,N_43549,N_42752);
or UO_2974 (O_2974,N_48092,N_41620);
xor UO_2975 (O_2975,N_47299,N_47484);
xnor UO_2976 (O_2976,N_40951,N_41740);
and UO_2977 (O_2977,N_44839,N_43880);
xnor UO_2978 (O_2978,N_41685,N_48969);
and UO_2979 (O_2979,N_47112,N_43398);
nand UO_2980 (O_2980,N_44179,N_49485);
xor UO_2981 (O_2981,N_44844,N_41395);
and UO_2982 (O_2982,N_44233,N_40946);
nand UO_2983 (O_2983,N_40415,N_48706);
and UO_2984 (O_2984,N_40627,N_47837);
xnor UO_2985 (O_2985,N_42363,N_42413);
nand UO_2986 (O_2986,N_45958,N_46110);
and UO_2987 (O_2987,N_44737,N_40507);
and UO_2988 (O_2988,N_41571,N_49027);
and UO_2989 (O_2989,N_49557,N_44594);
nand UO_2990 (O_2990,N_43819,N_41242);
xor UO_2991 (O_2991,N_43601,N_41530);
or UO_2992 (O_2992,N_47093,N_40115);
and UO_2993 (O_2993,N_41664,N_42298);
nor UO_2994 (O_2994,N_45236,N_49166);
xnor UO_2995 (O_2995,N_49258,N_48223);
nor UO_2996 (O_2996,N_41568,N_49045);
or UO_2997 (O_2997,N_40704,N_43227);
xnor UO_2998 (O_2998,N_40922,N_49658);
xor UO_2999 (O_2999,N_40668,N_45871);
nor UO_3000 (O_3000,N_44532,N_48696);
nor UO_3001 (O_3001,N_49866,N_45360);
and UO_3002 (O_3002,N_43282,N_41821);
xnor UO_3003 (O_3003,N_45782,N_47470);
nor UO_3004 (O_3004,N_40914,N_41466);
or UO_3005 (O_3005,N_40417,N_45724);
nor UO_3006 (O_3006,N_47094,N_44203);
or UO_3007 (O_3007,N_42493,N_45720);
nand UO_3008 (O_3008,N_41887,N_41235);
nand UO_3009 (O_3009,N_40722,N_45743);
xor UO_3010 (O_3010,N_46122,N_40148);
nor UO_3011 (O_3011,N_47253,N_48945);
xor UO_3012 (O_3012,N_44620,N_44998);
nor UO_3013 (O_3013,N_42345,N_48179);
nand UO_3014 (O_3014,N_46443,N_43062);
or UO_3015 (O_3015,N_42689,N_44130);
or UO_3016 (O_3016,N_47438,N_49134);
nand UO_3017 (O_3017,N_45343,N_49677);
nand UO_3018 (O_3018,N_41514,N_44796);
xnor UO_3019 (O_3019,N_48807,N_44181);
xnor UO_3020 (O_3020,N_44104,N_49820);
or UO_3021 (O_3021,N_41684,N_42374);
xor UO_3022 (O_3022,N_43244,N_47868);
or UO_3023 (O_3023,N_41928,N_44786);
and UO_3024 (O_3024,N_41708,N_47796);
or UO_3025 (O_3025,N_45304,N_49005);
and UO_3026 (O_3026,N_41517,N_43110);
or UO_3027 (O_3027,N_49473,N_42037);
nor UO_3028 (O_3028,N_48800,N_45264);
xor UO_3029 (O_3029,N_48881,N_48856);
nor UO_3030 (O_3030,N_45034,N_44180);
and UO_3031 (O_3031,N_46782,N_47230);
nor UO_3032 (O_3032,N_44795,N_45949);
or UO_3033 (O_3033,N_42888,N_45996);
or UO_3034 (O_3034,N_41890,N_48432);
xor UO_3035 (O_3035,N_48156,N_48414);
or UO_3036 (O_3036,N_43519,N_45559);
nor UO_3037 (O_3037,N_44070,N_40636);
xor UO_3038 (O_3038,N_44334,N_41336);
nand UO_3039 (O_3039,N_44672,N_48441);
nor UO_3040 (O_3040,N_40260,N_49525);
or UO_3041 (O_3041,N_49042,N_40524);
or UO_3042 (O_3042,N_49254,N_49191);
and UO_3043 (O_3043,N_42825,N_41019);
and UO_3044 (O_3044,N_43346,N_43114);
xnor UO_3045 (O_3045,N_44360,N_48683);
nand UO_3046 (O_3046,N_46473,N_47358);
and UO_3047 (O_3047,N_49071,N_44684);
xor UO_3048 (O_3048,N_49744,N_41139);
and UO_3049 (O_3049,N_45758,N_46983);
or UO_3050 (O_3050,N_47756,N_47201);
nor UO_3051 (O_3051,N_43143,N_44364);
nor UO_3052 (O_3052,N_46356,N_40838);
xnor UO_3053 (O_3053,N_43754,N_40401);
nor UO_3054 (O_3054,N_47547,N_45854);
and UO_3055 (O_3055,N_41627,N_40327);
nor UO_3056 (O_3056,N_44911,N_44628);
nand UO_3057 (O_3057,N_48482,N_49404);
xor UO_3058 (O_3058,N_43154,N_44914);
or UO_3059 (O_3059,N_42900,N_46162);
nand UO_3060 (O_3060,N_46265,N_46578);
xor UO_3061 (O_3061,N_46449,N_41489);
and UO_3062 (O_3062,N_48808,N_47664);
nor UO_3063 (O_3063,N_46277,N_45140);
nor UO_3064 (O_3064,N_42280,N_41618);
xor UO_3065 (O_3065,N_48657,N_47147);
nand UO_3066 (O_3066,N_44677,N_48232);
xor UO_3067 (O_3067,N_41069,N_46575);
and UO_3068 (O_3068,N_48964,N_43387);
or UO_3069 (O_3069,N_46452,N_43680);
nor UO_3070 (O_3070,N_44416,N_46604);
xnor UO_3071 (O_3071,N_48040,N_43586);
nand UO_3072 (O_3072,N_45708,N_43700);
nor UO_3073 (O_3073,N_40812,N_47020);
and UO_3074 (O_3074,N_46269,N_49669);
nand UO_3075 (O_3075,N_46907,N_40604);
nor UO_3076 (O_3076,N_49354,N_44711);
xor UO_3077 (O_3077,N_43638,N_45648);
and UO_3078 (O_3078,N_45686,N_41450);
and UO_3079 (O_3079,N_40746,N_41293);
nand UO_3080 (O_3080,N_42731,N_40582);
or UO_3081 (O_3081,N_43900,N_44073);
or UO_3082 (O_3082,N_43901,N_40907);
or UO_3083 (O_3083,N_47300,N_45185);
and UO_3084 (O_3084,N_49873,N_47060);
xor UO_3085 (O_3085,N_49411,N_48258);
nand UO_3086 (O_3086,N_42893,N_41941);
and UO_3087 (O_3087,N_41056,N_44531);
or UO_3088 (O_3088,N_41919,N_41806);
and UO_3089 (O_3089,N_44380,N_43758);
nand UO_3090 (O_3090,N_49052,N_49747);
xor UO_3091 (O_3091,N_48825,N_44264);
xor UO_3092 (O_3092,N_44891,N_41521);
nand UO_3093 (O_3093,N_45673,N_43093);
xor UO_3094 (O_3094,N_41132,N_40737);
nor UO_3095 (O_3095,N_40307,N_43366);
nand UO_3096 (O_3096,N_44704,N_43027);
or UO_3097 (O_3097,N_41404,N_42503);
and UO_3098 (O_3098,N_49803,N_44013);
nand UO_3099 (O_3099,N_48324,N_47782);
or UO_3100 (O_3100,N_49664,N_43208);
xor UO_3101 (O_3101,N_42636,N_45509);
nor UO_3102 (O_3102,N_45014,N_44383);
nand UO_3103 (O_3103,N_42564,N_47191);
nor UO_3104 (O_3104,N_43323,N_49537);
nor UO_3105 (O_3105,N_42176,N_43590);
or UO_3106 (O_3106,N_43767,N_42212);
xor UO_3107 (O_3107,N_43992,N_42715);
and UO_3108 (O_3108,N_46760,N_40886);
nor UO_3109 (O_3109,N_45735,N_47924);
and UO_3110 (O_3110,N_41072,N_48868);
and UO_3111 (O_3111,N_46044,N_49652);
nor UO_3112 (O_3112,N_48273,N_40937);
and UO_3113 (O_3113,N_42349,N_40859);
nand UO_3114 (O_3114,N_41668,N_48884);
nor UO_3115 (O_3115,N_40351,N_46060);
nor UO_3116 (O_3116,N_49675,N_41592);
nor UO_3117 (O_3117,N_45219,N_49053);
and UO_3118 (O_3118,N_40293,N_44263);
or UO_3119 (O_3119,N_45863,N_46771);
and UO_3120 (O_3120,N_43184,N_44408);
nor UO_3121 (O_3121,N_42844,N_46221);
or UO_3122 (O_3122,N_49460,N_44547);
xnor UO_3123 (O_3123,N_41049,N_43919);
nor UO_3124 (O_3124,N_40031,N_49365);
or UO_3125 (O_3125,N_46506,N_43253);
or UO_3126 (O_3126,N_43249,N_48147);
nand UO_3127 (O_3127,N_43661,N_41361);
xor UO_3128 (O_3128,N_43715,N_44879);
nand UO_3129 (O_3129,N_42236,N_47247);
xor UO_3130 (O_3130,N_47885,N_46914);
or UO_3131 (O_3131,N_48493,N_41552);
or UO_3132 (O_3132,N_41015,N_46704);
nand UO_3133 (O_3133,N_41636,N_44331);
xnor UO_3134 (O_3134,N_46446,N_42916);
and UO_3135 (O_3135,N_49787,N_43481);
nand UO_3136 (O_3136,N_47125,N_46994);
or UO_3137 (O_3137,N_49830,N_44979);
or UO_3138 (O_3138,N_42131,N_48546);
and UO_3139 (O_3139,N_46483,N_48658);
xor UO_3140 (O_3140,N_41526,N_43193);
and UO_3141 (O_3141,N_46510,N_40216);
and UO_3142 (O_3142,N_40020,N_43979);
nand UO_3143 (O_3143,N_43169,N_46558);
and UO_3144 (O_3144,N_43298,N_42958);
nand UO_3145 (O_3145,N_41405,N_44530);
and UO_3146 (O_3146,N_43621,N_47071);
nor UO_3147 (O_3147,N_40143,N_44987);
and UO_3148 (O_3148,N_41597,N_47566);
xnor UO_3149 (O_3149,N_44048,N_47288);
nand UO_3150 (O_3150,N_47208,N_40052);
and UO_3151 (O_3151,N_48761,N_46877);
and UO_3152 (O_3152,N_49556,N_48576);
and UO_3153 (O_3153,N_48337,N_48177);
nor UO_3154 (O_3154,N_43409,N_49081);
xor UO_3155 (O_3155,N_45061,N_41655);
nand UO_3156 (O_3156,N_41442,N_44469);
nor UO_3157 (O_3157,N_46802,N_40171);
nor UO_3158 (O_3158,N_44430,N_42111);
or UO_3159 (O_3159,N_42855,N_45746);
or UO_3160 (O_3160,N_48707,N_49229);
and UO_3161 (O_3161,N_40359,N_48457);
nor UO_3162 (O_3162,N_46137,N_41467);
nand UO_3163 (O_3163,N_48203,N_40522);
nand UO_3164 (O_3164,N_45258,N_41689);
nor UO_3165 (O_3165,N_41705,N_47317);
xor UO_3166 (O_3166,N_40234,N_48852);
xor UO_3167 (O_3167,N_48455,N_43145);
or UO_3168 (O_3168,N_43649,N_40282);
xnor UO_3169 (O_3169,N_44787,N_40672);
or UO_3170 (O_3170,N_41581,N_41412);
nor UO_3171 (O_3171,N_41728,N_49155);
nand UO_3172 (O_3172,N_43217,N_47244);
nand UO_3173 (O_3173,N_44896,N_45566);
nor UO_3174 (O_3174,N_43525,N_43670);
or UO_3175 (O_3175,N_45699,N_40719);
nor UO_3176 (O_3176,N_43874,N_41226);
xor UO_3177 (O_3177,N_45314,N_40204);
or UO_3178 (O_3178,N_45875,N_45293);
and UO_3179 (O_3179,N_42698,N_43061);
or UO_3180 (O_3180,N_44947,N_40166);
nor UO_3181 (O_3181,N_48519,N_47263);
nor UO_3182 (O_3182,N_41862,N_44055);
or UO_3183 (O_3183,N_45184,N_45528);
or UO_3184 (O_3184,N_46541,N_47595);
nand UO_3185 (O_3185,N_44556,N_46618);
or UO_3186 (O_3186,N_44455,N_45557);
nand UO_3187 (O_3187,N_40008,N_47224);
nand UO_3188 (O_3188,N_41106,N_46932);
nor UO_3189 (O_3189,N_40764,N_41471);
nand UO_3190 (O_3190,N_49893,N_48541);
nor UO_3191 (O_3191,N_44580,N_44133);
nand UO_3192 (O_3192,N_42625,N_45132);
and UO_3193 (O_3193,N_44885,N_46680);
xnor UO_3194 (O_3194,N_47016,N_44126);
nor UO_3195 (O_3195,N_42041,N_41669);
xor UO_3196 (O_3196,N_40024,N_47954);
or UO_3197 (O_3197,N_40268,N_45981);
and UO_3198 (O_3198,N_47678,N_41496);
xor UO_3199 (O_3199,N_41089,N_44997);
xnor UO_3200 (O_3200,N_46621,N_42599);
nand UO_3201 (O_3201,N_43538,N_46806);
and UO_3202 (O_3202,N_48294,N_47062);
xor UO_3203 (O_3203,N_45775,N_42972);
xor UO_3204 (O_3204,N_46248,N_45159);
or UO_3205 (O_3205,N_48299,N_48342);
or UO_3206 (O_3206,N_47860,N_44282);
and UO_3207 (O_3207,N_42654,N_41654);
or UO_3208 (O_3208,N_43236,N_41808);
xnor UO_3209 (O_3209,N_42905,N_45401);
nor UO_3210 (O_3210,N_48304,N_47891);
or UO_3211 (O_3211,N_44544,N_41356);
nand UO_3212 (O_3212,N_48268,N_42615);
nand UO_3213 (O_3213,N_44725,N_47649);
and UO_3214 (O_3214,N_44742,N_44480);
or UO_3215 (O_3215,N_45234,N_45276);
xor UO_3216 (O_3216,N_44191,N_40544);
or UO_3217 (O_3217,N_45974,N_41857);
xor UO_3218 (O_3218,N_42167,N_43757);
nor UO_3219 (O_3219,N_42769,N_48936);
and UO_3220 (O_3220,N_42877,N_49620);
or UO_3221 (O_3221,N_49776,N_44753);
xnor UO_3222 (O_3222,N_41984,N_47182);
xor UO_3223 (O_3223,N_42358,N_48369);
xnor UO_3224 (O_3224,N_47725,N_46748);
or UO_3225 (O_3225,N_42460,N_41124);
nor UO_3226 (O_3226,N_45296,N_45471);
or UO_3227 (O_3227,N_45983,N_42819);
nand UO_3228 (O_3228,N_44491,N_48567);
nand UO_3229 (O_3229,N_44260,N_40402);
nor UO_3230 (O_3230,N_49881,N_43418);
or UO_3231 (O_3231,N_46276,N_43140);
nor UO_3232 (O_3232,N_41184,N_42467);
nand UO_3233 (O_3233,N_42660,N_46471);
xor UO_3234 (O_3234,N_45533,N_45307);
and UO_3235 (O_3235,N_46744,N_40122);
nand UO_3236 (O_3236,N_48149,N_46234);
and UO_3237 (O_3237,N_41667,N_43464);
and UO_3238 (O_3238,N_47705,N_46729);
nand UO_3239 (O_3239,N_45049,N_40981);
and UO_3240 (O_3240,N_43888,N_40326);
nor UO_3241 (O_3241,N_49260,N_40593);
nand UO_3242 (O_3242,N_42682,N_40055);
xnor UO_3243 (O_3243,N_47277,N_48971);
nor UO_3244 (O_3244,N_40630,N_43916);
nand UO_3245 (O_3245,N_44479,N_43303);
or UO_3246 (O_3246,N_43163,N_47563);
xor UO_3247 (O_3247,N_49902,N_49699);
and UO_3248 (O_3248,N_43786,N_41064);
nand UO_3249 (O_3249,N_46499,N_42674);
nor UO_3250 (O_3250,N_45916,N_41607);
or UO_3251 (O_3251,N_48102,N_42504);
xnor UO_3252 (O_3252,N_40842,N_44595);
nor UO_3253 (O_3253,N_46511,N_46947);
xor UO_3254 (O_3254,N_49054,N_48918);
xor UO_3255 (O_3255,N_46934,N_45395);
xnor UO_3256 (O_3256,N_41874,N_44200);
nor UO_3257 (O_3257,N_47075,N_41996);
or UO_3258 (O_3258,N_43132,N_43551);
nand UO_3259 (O_3259,N_49433,N_42096);
nor UO_3260 (O_3260,N_42802,N_47716);
or UO_3261 (O_3261,N_41765,N_49246);
and UO_3262 (O_3262,N_47520,N_42373);
nand UO_3263 (O_3263,N_48773,N_43112);
nand UO_3264 (O_3264,N_41339,N_49077);
xnor UO_3265 (O_3265,N_43822,N_40113);
or UO_3266 (O_3266,N_49731,N_44925);
nand UO_3267 (O_3267,N_49737,N_44967);
or UO_3268 (O_3268,N_44330,N_43739);
nor UO_3269 (O_3269,N_43909,N_48989);
or UO_3270 (O_3270,N_43283,N_45115);
or UO_3271 (O_3271,N_43904,N_47103);
nand UO_3272 (O_3272,N_49464,N_42005);
or UO_3273 (O_3273,N_49165,N_49145);
and UO_3274 (O_3274,N_47989,N_43068);
nand UO_3275 (O_3275,N_42372,N_46201);
nor UO_3276 (O_3276,N_43080,N_46056);
nand UO_3277 (O_3277,N_41457,N_42558);
nand UO_3278 (O_3278,N_48398,N_46735);
and UO_3279 (O_3279,N_43250,N_43229);
and UO_3280 (O_3280,N_46114,N_45281);
nand UO_3281 (O_3281,N_47312,N_40680);
nand UO_3282 (O_3282,N_44170,N_44135);
xor UO_3283 (O_3283,N_47902,N_43189);
nor UO_3284 (O_3284,N_44417,N_43044);
nor UO_3285 (O_3285,N_44769,N_40725);
nand UO_3286 (O_3286,N_45399,N_49741);
and UO_3287 (O_3287,N_49236,N_46580);
or UO_3288 (O_3288,N_46753,N_43612);
and UO_3289 (O_3289,N_42370,N_43541);
nor UO_3290 (O_3290,N_40042,N_44561);
and UO_3291 (O_3291,N_48412,N_45687);
and UO_3292 (O_3292,N_45150,N_41264);
nor UO_3293 (O_3293,N_46980,N_41236);
and UO_3294 (O_3294,N_48087,N_49067);
xnor UO_3295 (O_3295,N_49768,N_45214);
xnor UO_3296 (O_3296,N_47412,N_40421);
nand UO_3297 (O_3297,N_41199,N_44291);
and UO_3298 (O_3298,N_40051,N_43055);
and UO_3299 (O_3299,N_43242,N_46063);
and UO_3300 (O_3300,N_48988,N_42222);
and UO_3301 (O_3301,N_40712,N_41479);
or UO_3302 (O_3302,N_40154,N_43299);
nand UO_3303 (O_3303,N_45172,N_47636);
xnor UO_3304 (O_3304,N_40865,N_46169);
nand UO_3305 (O_3305,N_41882,N_48204);
and UO_3306 (O_3306,N_40175,N_49201);
or UO_3307 (O_3307,N_49748,N_42414);
xnor UO_3308 (O_3308,N_43222,N_49276);
or UO_3309 (O_3309,N_46869,N_46710);
xor UO_3310 (O_3310,N_44859,N_45397);
and UO_3311 (O_3311,N_42848,N_41780);
xnor UO_3312 (O_3312,N_40366,N_47915);
xnor UO_3313 (O_3313,N_41426,N_47507);
and UO_3314 (O_3314,N_42793,N_44322);
or UO_3315 (O_3315,N_44142,N_43755);
nand UO_3316 (O_3316,N_42523,N_47898);
or UO_3317 (O_3317,N_48916,N_46797);
nor UO_3318 (O_3318,N_40057,N_42230);
nor UO_3319 (O_3319,N_45903,N_41690);
nor UO_3320 (O_3320,N_42628,N_41294);
nand UO_3321 (O_3321,N_42965,N_43477);
or UO_3322 (O_3322,N_44397,N_44431);
or UO_3323 (O_3323,N_45872,N_43567);
nor UO_3324 (O_3324,N_42773,N_41881);
nor UO_3325 (O_3325,N_49793,N_45787);
nand UO_3326 (O_3326,N_49540,N_41836);
xnor UO_3327 (O_3327,N_40969,N_43074);
xnor UO_3328 (O_3328,N_40112,N_40659);
and UO_3329 (O_3329,N_48698,N_44405);
or UO_3330 (O_3330,N_47941,N_48547);
nor UO_3331 (O_3331,N_47673,N_47675);
nand UO_3332 (O_3332,N_46297,N_49474);
nand UO_3333 (O_3333,N_49632,N_46653);
nand UO_3334 (O_3334,N_43160,N_45120);
or UO_3335 (O_3335,N_42623,N_43765);
xnor UO_3336 (O_3336,N_43929,N_46379);
nand UO_3337 (O_3337,N_42340,N_48578);
xnor UO_3338 (O_3338,N_48953,N_43399);
and UO_3339 (O_3339,N_42405,N_49676);
and UO_3340 (O_3340,N_41097,N_47939);
nand UO_3341 (O_3341,N_42323,N_49372);
or UO_3342 (O_3342,N_46521,N_40409);
xor UO_3343 (O_3343,N_42277,N_47543);
nand UO_3344 (O_3344,N_41119,N_47823);
nand UO_3345 (O_3345,N_44528,N_41034);
xnor UO_3346 (O_3346,N_47579,N_48089);
nor UO_3347 (O_3347,N_48123,N_46562);
or UO_3348 (O_3348,N_49770,N_45171);
nor UO_3349 (O_3349,N_42969,N_42290);
nand UO_3350 (O_3350,N_44345,N_48999);
nand UO_3351 (O_3351,N_49168,N_47279);
or UO_3352 (O_3352,N_44566,N_48797);
nor UO_3353 (O_3353,N_49690,N_48420);
or UO_3354 (O_3354,N_47737,N_47363);
nand UO_3355 (O_3355,N_47790,N_49408);
nand UO_3356 (O_3356,N_44706,N_45738);
and UO_3357 (O_3357,N_44399,N_49799);
or UO_3358 (O_3358,N_43336,N_47994);
and UO_3359 (O_3359,N_42438,N_43885);
or UO_3360 (O_3360,N_42455,N_45005);
xor UO_3361 (O_3361,N_44031,N_42281);
nor UO_3362 (O_3362,N_42159,N_42780);
nor UO_3363 (O_3363,N_44575,N_45979);
nand UO_3364 (O_3364,N_43340,N_41368);
and UO_3365 (O_3365,N_40709,N_47429);
or UO_3366 (O_3366,N_43205,N_41263);
or UO_3367 (O_3367,N_43215,N_41180);
nand UO_3368 (O_3368,N_48352,N_44837);
nand UO_3369 (O_3369,N_43679,N_42524);
xor UO_3370 (O_3370,N_40295,N_43787);
and UO_3371 (O_3371,N_49849,N_48465);
nand UO_3372 (O_3372,N_40249,N_45406);
nand UO_3373 (O_3373,N_42879,N_45087);
or UO_3374 (O_3374,N_41734,N_48105);
or UO_3375 (O_3375,N_45325,N_42747);
xor UO_3376 (O_3376,N_40292,N_42471);
nand UO_3377 (O_3377,N_43848,N_41776);
nor UO_3378 (O_3378,N_43129,N_41416);
nor UO_3379 (O_3379,N_45243,N_49043);
and UO_3380 (O_3380,N_40535,N_41992);
nor UO_3381 (O_3381,N_44912,N_46136);
nand UO_3382 (O_3382,N_43391,N_40161);
and UO_3383 (O_3383,N_43494,N_46069);
or UO_3384 (O_3384,N_47791,N_48853);
nor UO_3385 (O_3385,N_47315,N_47478);
or UO_3386 (O_3386,N_41022,N_44246);
nor UO_3387 (O_3387,N_47184,N_40717);
nor UO_3388 (O_3388,N_44735,N_48315);
xnor UO_3389 (O_3389,N_45602,N_43642);
or UO_3390 (O_3390,N_48362,N_44720);
or UO_3391 (O_3391,N_48175,N_42638);
or UO_3392 (O_3392,N_41314,N_45074);
nor UO_3393 (O_3393,N_43871,N_47887);
and UO_3394 (O_3394,N_46982,N_41432);
xnor UO_3395 (O_3395,N_43034,N_42366);
nor UO_3396 (O_3396,N_42745,N_40319);
or UO_3397 (O_3397,N_44543,N_40694);
nand UO_3398 (O_3398,N_48570,N_44025);
or UO_3399 (O_3399,N_40996,N_46413);
xor UO_3400 (O_3400,N_49336,N_49959);
nand UO_3401 (O_3401,N_46927,N_41425);
xnor UO_3402 (O_3402,N_42498,N_46178);
and UO_3403 (O_3403,N_40444,N_46439);
xnor UO_3404 (O_3404,N_43802,N_46800);
and UO_3405 (O_3405,N_47398,N_44034);
or UO_3406 (O_3406,N_42821,N_45379);
and UO_3407 (O_3407,N_44185,N_48867);
nand UO_3408 (O_3408,N_43350,N_49175);
xor UO_3409 (O_3409,N_48168,N_41190);
nor UO_3410 (O_3410,N_40904,N_45570);
nor UO_3411 (O_3411,N_46945,N_41096);
and UO_3412 (O_3412,N_41204,N_44728);
and UO_3413 (O_3413,N_40242,N_46959);
nand UO_3414 (O_3414,N_47265,N_47806);
nand UO_3415 (O_3415,N_41676,N_44335);
and UO_3416 (O_3416,N_46315,N_48248);
or UO_3417 (O_3417,N_45112,N_46230);
nand UO_3418 (O_3418,N_49325,N_47012);
and UO_3419 (O_3419,N_43211,N_45090);
and UO_3420 (O_3420,N_45529,N_48466);
nor UO_3421 (O_3421,N_43499,N_44398);
nor UO_3422 (O_3422,N_41579,N_46239);
nand UO_3423 (O_3423,N_43558,N_48464);
or UO_3424 (O_3424,N_45092,N_41178);
or UO_3425 (O_3425,N_48297,N_40367);
and UO_3426 (O_3426,N_49694,N_45940);
and UO_3427 (O_3427,N_49683,N_48074);
or UO_3428 (O_3428,N_46896,N_43587);
and UO_3429 (O_3429,N_40587,N_48692);
nor UO_3430 (O_3430,N_47068,N_46727);
nand UO_3431 (O_3431,N_44326,N_43894);
and UO_3432 (O_3432,N_44923,N_46552);
nand UO_3433 (O_3433,N_43630,N_48535);
and UO_3434 (O_3434,N_49440,N_44700);
and UO_3435 (O_3435,N_44486,N_48407);
or UO_3436 (O_3436,N_45517,N_40884);
nor UO_3437 (O_3437,N_47327,N_48195);
or UO_3438 (O_3438,N_45291,N_46231);
nor UO_3439 (O_3439,N_44870,N_43097);
and UO_3440 (O_3440,N_43459,N_45561);
xnor UO_3441 (O_3441,N_47145,N_40982);
nor UO_3442 (O_3442,N_42367,N_45072);
nand UO_3443 (O_3443,N_43654,N_47130);
xor UO_3444 (O_3444,N_43809,N_47603);
or UO_3445 (O_3445,N_46667,N_48998);
nand UO_3446 (O_3446,N_48524,N_45924);
and UO_3447 (O_3447,N_48779,N_45155);
nor UO_3448 (O_3448,N_42561,N_48824);
nor UO_3449 (O_3449,N_41325,N_44775);
nor UO_3450 (O_3450,N_40037,N_48088);
nand UO_3451 (O_3451,N_42043,N_40915);
and UO_3452 (O_3452,N_44363,N_47797);
nand UO_3453 (O_3453,N_43972,N_47554);
nand UO_3454 (O_3454,N_41084,N_40967);
and UO_3455 (O_3455,N_42662,N_48196);
and UO_3456 (O_3456,N_46469,N_49035);
xor UO_3457 (O_3457,N_49117,N_41736);
nand UO_3458 (O_3458,N_41587,N_49038);
nand UO_3459 (O_3459,N_42068,N_44604);
nand UO_3460 (O_3460,N_47995,N_42492);
nand UO_3461 (O_3461,N_44827,N_48895);
nand UO_3462 (O_3462,N_41803,N_43354);
nand UO_3463 (O_3463,N_49549,N_45852);
nand UO_3464 (O_3464,N_44901,N_46966);
nand UO_3465 (O_3465,N_47142,N_40927);
nand UO_3466 (O_3466,N_48128,N_45990);
nor UO_3467 (O_3467,N_45975,N_40810);
or UO_3468 (O_3468,N_45749,N_42713);
nor UO_3469 (O_3469,N_46344,N_42621);
nand UO_3470 (O_3470,N_46629,N_43123);
nor UO_3471 (O_3471,N_48551,N_42472);
or UO_3472 (O_3472,N_42842,N_40442);
or UO_3473 (O_3473,N_41146,N_40635);
or UO_3474 (O_3474,N_40667,N_40848);
nor UO_3475 (O_3475,N_43353,N_44644);
xnor UO_3476 (O_3476,N_49604,N_48963);
and UO_3477 (O_3477,N_44081,N_48529);
xnor UO_3478 (O_3478,N_42543,N_47377);
or UO_3479 (O_3479,N_49076,N_48801);
nand UO_3480 (O_3480,N_48222,N_48735);
and UO_3481 (O_3481,N_44655,N_40698);
xor UO_3482 (O_3482,N_49477,N_49323);
nor UO_3483 (O_3483,N_43137,N_43956);
nor UO_3484 (O_3484,N_45656,N_42837);
and UO_3485 (O_3485,N_43443,N_47019);
xnor UO_3486 (O_3486,N_43449,N_47303);
nor UO_3487 (O_3487,N_48584,N_48516);
nor UO_3488 (O_3488,N_48839,N_47666);
xnor UO_3489 (O_3489,N_47738,N_41913);
xor UO_3490 (O_3490,N_48329,N_42175);
and UO_3491 (O_3491,N_45900,N_47633);
or UO_3492 (O_3492,N_49047,N_48790);
nand UO_3493 (O_3493,N_46177,N_40765);
or UO_3494 (O_3494,N_48755,N_46376);
nand UO_3495 (O_3495,N_47884,N_45408);
nand UO_3496 (O_3496,N_42526,N_47018);
nand UO_3497 (O_3497,N_43741,N_40490);
or UO_3498 (O_3498,N_49769,N_44584);
nor UO_3499 (O_3499,N_42858,N_49754);
xor UO_3500 (O_3500,N_45845,N_41274);
or UO_3501 (O_3501,N_48353,N_45095);
nor UO_3502 (O_3502,N_44220,N_42935);
xnor UO_3503 (O_3503,N_46707,N_49756);
xnor UO_3504 (O_3504,N_42597,N_48060);
xor UO_3505 (O_3505,N_48443,N_43051);
or UO_3506 (O_3506,N_42685,N_40893);
xor UO_3507 (O_3507,N_44366,N_49310);
or UO_3508 (O_3508,N_40743,N_47914);
and UO_3509 (O_3509,N_42137,N_42316);
nand UO_3510 (O_3510,N_43207,N_40539);
and UO_3511 (O_3511,N_43434,N_47784);
nand UO_3512 (O_3512,N_45878,N_47571);
nand UO_3513 (O_3513,N_41744,N_46815);
nand UO_3514 (O_3514,N_45103,N_40784);
or UO_3515 (O_3515,N_49773,N_41102);
and UO_3516 (O_3516,N_46948,N_48539);
or UO_3517 (O_3517,N_49780,N_44029);
and UO_3518 (O_3518,N_44621,N_46501);
nor UO_3519 (O_3519,N_46173,N_43133);
and UO_3520 (O_3520,N_45082,N_40200);
nand UO_3521 (O_3521,N_44830,N_43836);
or UO_3522 (O_3522,N_47138,N_43855);
or UO_3523 (O_3523,N_42673,N_46107);
nor UO_3524 (O_3524,N_41843,N_47458);
xor UO_3525 (O_3525,N_47632,N_40423);
nand UO_3526 (O_3526,N_46059,N_48269);
nand UO_3527 (O_3527,N_41516,N_49129);
xnor UO_3528 (O_3528,N_49960,N_40034);
and UO_3529 (O_3529,N_46189,N_49217);
nand UO_3530 (O_3530,N_44828,N_49097);
nor UO_3531 (O_3531,N_42750,N_41078);
nand UO_3532 (O_3532,N_41000,N_41240);
and UO_3533 (O_3533,N_44674,N_46788);
or UO_3534 (O_3534,N_42066,N_49789);
nor UO_3535 (O_3535,N_47374,N_45270);
xnor UO_3536 (O_3536,N_47453,N_45668);
xor UO_3537 (O_3537,N_44797,N_47445);
xor UO_3538 (O_3538,N_43969,N_44926);
nor UO_3539 (O_3539,N_48559,N_42369);
xnor UO_3540 (O_3540,N_41281,N_46166);
nand UO_3541 (O_3541,N_47158,N_48247);
or UO_3542 (O_3542,N_49380,N_49657);
nand UO_3543 (O_3543,N_46361,N_44994);
xnor UO_3544 (O_3544,N_42170,N_48646);
or UO_3545 (O_3545,N_44681,N_45739);
or UO_3546 (O_3546,N_48672,N_47450);
and UO_3547 (O_3547,N_43958,N_48754);
or UO_3548 (O_3548,N_48528,N_49470);
or UO_3549 (O_3549,N_48673,N_40283);
and UO_3550 (O_3550,N_48107,N_40603);
or UO_3551 (O_3551,N_41462,N_43774);
or UO_3552 (O_3552,N_49025,N_47672);
or UO_3553 (O_3553,N_45661,N_45271);
and UO_3554 (O_3554,N_43128,N_48452);
nor UO_3555 (O_3555,N_47968,N_42719);
xor UO_3556 (O_3556,N_44060,N_46951);
and UO_3557 (O_3557,N_41522,N_46430);
or UO_3558 (O_3558,N_41529,N_43713);
nor UO_3559 (O_3559,N_45536,N_46100);
nor UO_3560 (O_3560,N_44214,N_48601);
nand UO_3561 (O_3561,N_45777,N_48548);
xor UO_3562 (O_3562,N_45138,N_46365);
and UO_3563 (O_3563,N_43064,N_48063);
nand UO_3564 (O_3564,N_40759,N_41229);
and UO_3565 (O_3565,N_43864,N_40573);
or UO_3566 (O_3566,N_45959,N_40471);
nand UO_3567 (O_3567,N_47642,N_45485);
nand UO_3568 (O_3568,N_42826,N_43127);
nand UO_3569 (O_3569,N_41495,N_45590);
or UO_3570 (O_3570,N_42010,N_43753);
nand UO_3571 (O_3571,N_43945,N_48068);
nor UO_3572 (O_3572,N_48665,N_42060);
or UO_3573 (O_3573,N_47724,N_42902);
nor UO_3574 (O_3574,N_46420,N_46536);
nor UO_3575 (O_3575,N_45639,N_41868);
or UO_3576 (O_3576,N_47857,N_43441);
nand UO_3577 (O_3577,N_43595,N_48720);
and UO_3578 (O_3578,N_40018,N_44348);
or UO_3579 (O_3579,N_41891,N_42260);
or UO_3580 (O_3580,N_43139,N_40164);
nand UO_3581 (O_3581,N_42661,N_49501);
or UO_3582 (O_3582,N_46838,N_48870);
xor UO_3583 (O_3583,N_41677,N_46351);
nor UO_3584 (O_3584,N_42324,N_42337);
nor UO_3585 (O_3585,N_41609,N_42045);
xnor UO_3586 (O_3586,N_45349,N_47964);
nand UO_3587 (O_3587,N_43491,N_42310);
nor UO_3588 (O_3588,N_44964,N_44117);
nor UO_3589 (O_3589,N_45789,N_43875);
xnor UO_3590 (O_3590,N_40763,N_45630);
or UO_3591 (O_3591,N_47715,N_43720);
nor UO_3592 (O_3592,N_49895,N_42246);
and UO_3593 (O_3593,N_49079,N_43605);
and UO_3594 (O_3594,N_45676,N_43065);
xnor UO_3595 (O_3595,N_48832,N_41187);
or UO_3596 (O_3596,N_46422,N_47233);
nand UO_3597 (O_3597,N_41193,N_44358);
xnor UO_3598 (O_3598,N_45882,N_42116);
nor UO_3599 (O_3599,N_48400,N_46505);
nor UO_3600 (O_3600,N_46984,N_46337);
xor UO_3601 (O_3601,N_45446,N_41908);
or UO_3602 (O_3602,N_42021,N_47384);
or UO_3603 (O_3603,N_44468,N_41256);
and UO_3604 (O_3604,N_47854,N_42179);
or UO_3605 (O_3605,N_42910,N_40542);
nand UO_3606 (O_3606,N_44465,N_48580);
and UO_3607 (O_3607,N_49919,N_48328);
xnor UO_3608 (O_3608,N_44378,N_49827);
or UO_3609 (O_3609,N_40378,N_48496);
nand UO_3610 (O_3610,N_46634,N_45392);
or UO_3611 (O_3611,N_42440,N_49219);
or UO_3612 (O_3612,N_46745,N_45166);
xnor UO_3613 (O_3613,N_46691,N_49399);
and UO_3614 (O_3614,N_47127,N_46076);
and UO_3615 (O_3615,N_42657,N_42423);
nor UO_3616 (O_3616,N_49149,N_43006);
and UO_3617 (O_3617,N_44077,N_43148);
nand UO_3618 (O_3618,N_45088,N_47940);
or UO_3619 (O_3619,N_46596,N_43704);
nor UO_3620 (O_3620,N_42511,N_48158);
xor UO_3621 (O_3621,N_42495,N_40408);
xnor UO_3622 (O_3622,N_40219,N_46281);
nor UO_3623 (O_3623,N_49700,N_47069);
xnor UO_3624 (O_3624,N_42403,N_40467);
xnor UO_3625 (O_3625,N_43769,N_41706);
or UO_3626 (O_3626,N_43962,N_49654);
and UO_3627 (O_3627,N_41582,N_41437);
and UO_3628 (O_3628,N_43330,N_44292);
or UO_3629 (O_3629,N_40039,N_45753);
nand UO_3630 (O_3630,N_48549,N_48028);
nand UO_3631 (O_3631,N_43524,N_43800);
xnor UO_3632 (O_3632,N_42106,N_43783);
or UO_3633 (O_3633,N_41629,N_48704);
or UO_3634 (O_3634,N_42424,N_47361);
xnor UO_3635 (O_3635,N_44553,N_48515);
nand UO_3636 (O_3636,N_40220,N_47592);
nand UO_3637 (O_3637,N_44936,N_41024);
and UO_3638 (O_3638,N_41770,N_49472);
and UO_3639 (O_3639,N_46933,N_48727);
nand UO_3640 (O_3640,N_49277,N_45938);
xnor UO_3641 (O_3641,N_44268,N_44053);
nor UO_3642 (O_3642,N_43627,N_43396);
or UO_3643 (O_3643,N_43343,N_42177);
nand UO_3644 (O_3644,N_46341,N_41455);
nor UO_3645 (O_3645,N_43325,N_45670);
or UO_3646 (O_3646,N_48627,N_49153);
nand UO_3647 (O_3647,N_48770,N_47457);
and UO_3648 (O_3648,N_41842,N_45237);
or UO_3649 (O_3649,N_40414,N_43918);
nor UO_3650 (O_3650,N_43116,N_44231);
xor UO_3651 (O_3651,N_48067,N_45541);
nor UO_3652 (O_3652,N_41174,N_40259);
and UO_3653 (O_3653,N_40336,N_49587);
nand UO_3654 (O_3654,N_43043,N_48322);
xnor UO_3655 (O_3655,N_49548,N_47206);
nor UO_3656 (O_3656,N_44461,N_49162);
or UO_3657 (O_3657,N_43555,N_41527);
xnor UO_3658 (O_3658,N_46045,N_45417);
nand UO_3659 (O_3659,N_44390,N_40265);
or UO_3660 (O_3660,N_42441,N_44274);
xor UO_3661 (O_3661,N_43502,N_49867);
nand UO_3662 (O_3662,N_40372,N_48642);
or UO_3663 (O_3663,N_45717,N_45305);
and UO_3664 (O_3664,N_43364,N_42917);
xor UO_3665 (O_3665,N_41129,N_48650);
or UO_3666 (O_3666,N_46816,N_43859);
nand UO_3667 (O_3667,N_47828,N_47375);
nor UO_3668 (O_3668,N_41885,N_41812);
nand UO_3669 (O_3669,N_45831,N_41474);
or UO_3670 (O_3670,N_42559,N_40702);
and UO_3671 (O_3671,N_42075,N_41104);
nand UO_3672 (O_3672,N_43975,N_46803);
xnor UO_3673 (O_3673,N_40419,N_41980);
xor UO_3674 (O_3674,N_47871,N_45041);
and UO_3675 (O_3675,N_48478,N_42737);
xor UO_3676 (O_3676,N_43458,N_41628);
or UO_3677 (O_3677,N_48975,N_47213);
and UO_3678 (O_3678,N_45310,N_49188);
or UO_3679 (O_3679,N_41352,N_42245);
nor UO_3680 (O_3680,N_43089,N_45055);
or UO_3681 (O_3681,N_41926,N_49285);
or UO_3682 (O_3682,N_47814,N_46424);
or UO_3683 (O_3683,N_47072,N_40425);
or UO_3684 (O_3684,N_41884,N_46272);
nor UO_3685 (O_3685,N_44344,N_46520);
and UO_3686 (O_3686,N_49006,N_47808);
nand UO_3687 (O_3687,N_49130,N_48686);
xor UO_3688 (O_3688,N_42658,N_41869);
nor UO_3689 (O_3689,N_45586,N_41539);
and UO_3690 (O_3690,N_48375,N_49425);
or UO_3691 (O_3691,N_41071,N_49634);
or UO_3692 (O_3692,N_49692,N_47532);
and UO_3693 (O_3693,N_42716,N_41995);
and UO_3694 (O_3694,N_41711,N_44186);
and UO_3695 (O_3695,N_40438,N_47340);
and UO_3696 (O_3696,N_46898,N_47972);
xor UO_3697 (O_3697,N_43653,N_46213);
nand UO_3698 (O_3698,N_43223,N_47486);
or UO_3699 (O_3699,N_44741,N_42763);
or UO_3700 (O_3700,N_49218,N_47048);
nor UO_3701 (O_3701,N_41603,N_46364);
or UO_3702 (O_3702,N_46482,N_44429);
and UO_3703 (O_3703,N_49124,N_47557);
xor UO_3704 (O_3704,N_42904,N_47120);
and UO_3705 (O_3705,N_47696,N_44918);
nor UO_3706 (O_3706,N_40705,N_43537);
xnor UO_3707 (O_3707,N_45841,N_46654);
or UO_3708 (O_3708,N_47242,N_47732);
nand UO_3709 (O_3709,N_45128,N_40196);
nor UO_3710 (O_3710,N_49844,N_40989);
nor UO_3711 (O_3711,N_43392,N_47212);
nor UO_3712 (O_3712,N_46850,N_44303);
and UO_3713 (O_3713,N_49193,N_46054);
nor UO_3714 (O_3714,N_44236,N_49023);
xor UO_3715 (O_3715,N_44937,N_45040);
xor UO_3716 (O_3716,N_44276,N_42029);
and UO_3717 (O_3717,N_47697,N_40344);
nand UO_3718 (O_3718,N_43729,N_45501);
or UO_3719 (O_3719,N_42513,N_42333);
xnor UO_3720 (O_3720,N_41259,N_41693);
or UO_3721 (O_3721,N_48784,N_45142);
xor UO_3722 (O_3722,N_44597,N_40095);
nor UO_3723 (O_3723,N_43483,N_48710);
nor UO_3724 (O_3724,N_45168,N_42346);
and UO_3725 (O_3725,N_46292,N_48178);
xnor UO_3726 (O_3726,N_44718,N_43789);
nand UO_3727 (O_3727,N_40887,N_41454);
xor UO_3728 (O_3728,N_43095,N_49884);
nand UO_3729 (O_3729,N_49614,N_45568);
and UO_3730 (O_3730,N_46115,N_47695);
and UO_3731 (O_3731,N_45436,N_49172);
nand UO_3732 (O_3732,N_40486,N_41838);
xor UO_3733 (O_3733,N_40985,N_45050);
nor UO_3734 (O_3734,N_45482,N_48669);
nand UO_3735 (O_3735,N_41030,N_48679);
nor UO_3736 (O_3736,N_49806,N_46042);
nand UO_3737 (O_3737,N_46864,N_40687);
nand UO_3738 (O_3738,N_43847,N_43641);
nand UO_3739 (O_3739,N_43386,N_49289);
nand UO_3740 (O_3740,N_45976,N_40975);
nor UO_3741 (O_3741,N_42813,N_48411);
nand UO_3742 (O_3742,N_42474,N_42827);
xnor UO_3743 (O_3743,N_45002,N_49788);
or UO_3744 (O_3744,N_47334,N_42739);
xor UO_3745 (O_3745,N_49834,N_40594);
xnor UO_3746 (O_3746,N_48360,N_45181);
and UO_3747 (O_3747,N_42026,N_48090);
nand UO_3748 (O_3748,N_43569,N_43437);
nor UO_3749 (O_3749,N_40285,N_41715);
or UO_3750 (O_3750,N_46999,N_48724);
xnor UO_3751 (O_3751,N_44310,N_43360);
nand UO_3752 (O_3752,N_47752,N_47351);
nand UO_3753 (O_3753,N_46259,N_49706);
and UO_3754 (O_3754,N_43598,N_43550);
xnor UO_3755 (O_3755,N_47512,N_45405);
or UO_3756 (O_3756,N_49619,N_49309);
nor UO_3757 (O_3757,N_48048,N_41116);
nor UO_3758 (O_3758,N_40233,N_44886);
nand UO_3759 (O_3759,N_40162,N_43619);
nor UO_3760 (O_3760,N_41671,N_46534);
nor UO_3761 (O_3761,N_41472,N_48334);
or UO_3762 (O_3762,N_48922,N_43045);
nand UO_3763 (O_3763,N_44618,N_40619);
or UO_3764 (O_3764,N_48434,N_44631);
or UO_3765 (O_3765,N_45578,N_46906);
xor UO_3766 (O_3766,N_47638,N_42140);
nor UO_3767 (O_3767,N_40049,N_49592);
or UO_3768 (O_3768,N_46047,N_48051);
nor UO_3769 (O_3769,N_40338,N_49944);
nand UO_3770 (O_3770,N_44895,N_44974);
nand UO_3771 (O_3771,N_47359,N_45995);
nand UO_3772 (O_3772,N_45433,N_43963);
and UO_3773 (O_3773,N_47057,N_40331);
nand UO_3774 (O_3774,N_41642,N_44450);
or UO_3775 (O_3775,N_49423,N_49576);
and UO_3776 (O_3776,N_42335,N_42117);
nand UO_3777 (O_3777,N_43858,N_48610);
nor UO_3778 (O_3778,N_43943,N_45851);
nor UO_3779 (O_3779,N_49441,N_47401);
nor UO_3780 (O_3780,N_49763,N_48172);
or UO_3781 (O_3781,N_41680,N_40500);
nand UO_3782 (O_3782,N_45688,N_42831);
nor UO_3783 (O_3783,N_49573,N_44202);
nor UO_3784 (O_3784,N_40800,N_49065);
nand UO_3785 (O_3785,N_44843,N_45759);
xnor UO_3786 (O_3786,N_45516,N_41905);
or UO_3787 (O_3787,N_43255,N_42947);
and UO_3788 (O_3788,N_40877,N_48019);
nor UO_3789 (O_3789,N_47059,N_43842);
nand UO_3790 (O_3790,N_49571,N_44035);
and UO_3791 (O_3791,N_45012,N_43281);
and UO_3792 (O_3792,N_44312,N_44134);
nand UO_3793 (O_3793,N_48717,N_41756);
xor UO_3794 (O_3794,N_47707,N_42939);
nand UO_3795 (O_3795,N_41169,N_47879);
xor UO_3796 (O_3796,N_47691,N_47413);
nor UO_3797 (O_3797,N_46889,N_44692);
or UO_3798 (O_3798,N_47927,N_47545);
and UO_3799 (O_3799,N_44353,N_43498);
and UO_3800 (O_3800,N_45157,N_45927);
and UO_3801 (O_3801,N_42717,N_46257);
xor UO_3802 (O_3802,N_49547,N_47101);
nand UO_3803 (O_3803,N_41931,N_43966);
xnor UO_3804 (O_3804,N_42708,N_42509);
nor UO_3805 (O_3805,N_47258,N_41720);
nor UO_3806 (O_3806,N_47394,N_43338);
or UO_3807 (O_3807,N_47801,N_45163);
xor UO_3808 (O_3808,N_41768,N_48349);
or UO_3809 (O_3809,N_44316,N_40815);
nand UO_3810 (O_3810,N_43640,N_42562);
nor UO_3811 (O_3811,N_41861,N_40934);
nor UO_3812 (O_3812,N_48668,N_41703);
xnor UO_3813 (O_3813,N_41601,N_42861);
nor UO_3814 (O_3814,N_46164,N_40424);
nor UO_3815 (O_3815,N_49832,N_49120);
xnor UO_3816 (O_3816,N_48902,N_41841);
xnor UO_3817 (O_3817,N_45153,N_43098);
and UO_3818 (O_3818,N_45484,N_47389);
nor UO_3819 (O_3819,N_49761,N_47210);
nand UO_3820 (O_3820,N_43563,N_43152);
and UO_3821 (O_3821,N_48688,N_42381);
nor UO_3822 (O_3822,N_45683,N_40138);
or UO_3823 (O_3823,N_49009,N_46381);
xor UO_3824 (O_3824,N_41448,N_44226);
nand UO_3825 (O_3825,N_49814,N_48174);
nand UO_3826 (O_3826,N_41814,N_46783);
nand UO_3827 (O_3827,N_46171,N_48739);
nor UO_3828 (O_3828,N_41342,N_42824);
nand UO_3829 (O_3829,N_46237,N_41156);
nand UO_3830 (O_3830,N_46378,N_46946);
xor UO_3831 (O_3831,N_49058,N_42582);
nand UO_3832 (O_3832,N_42940,N_42113);
or UO_3833 (O_3833,N_49090,N_42006);
and UO_3834 (O_3834,N_49458,N_45147);
and UO_3835 (O_3835,N_44173,N_42514);
nand UO_3836 (O_3836,N_46223,N_40135);
xor UO_3837 (O_3837,N_42053,N_41982);
and UO_3838 (O_3838,N_42748,N_47933);
xnor UO_3839 (O_3839,N_44349,N_48061);
nand UO_3840 (O_3840,N_47781,N_40302);
nor UO_3841 (O_3841,N_46015,N_41683);
and UO_3842 (O_3842,N_41754,N_42315);
xor UO_3843 (O_3843,N_42567,N_45452);
xnor UO_3844 (O_3844,N_47548,N_49393);
xor UO_3845 (O_3845,N_41113,N_43825);
nor UO_3846 (O_3846,N_45694,N_40867);
or UO_3847 (O_3847,N_44866,N_41166);
or UO_3848 (O_3848,N_41149,N_40890);
nand UO_3849 (O_3849,N_45342,N_45083);
xnor UO_3850 (O_3850,N_40227,N_48783);
or UO_3851 (O_3851,N_44000,N_48968);
or UO_3852 (O_3852,N_49765,N_48117);
and UO_3853 (O_3853,N_48131,N_47794);
nor UO_3854 (O_3854,N_48025,N_45275);
and UO_3855 (O_3855,N_46862,N_43479);
and UO_3856 (O_3856,N_40069,N_45280);
and UO_3857 (O_3857,N_48311,N_48530);
xor UO_3858 (O_3858,N_47073,N_47993);
nand UO_3859 (O_3859,N_42530,N_42215);
and UO_3860 (O_3860,N_45260,N_44999);
nor UO_3861 (O_3861,N_43553,N_46950);
and UO_3862 (O_3862,N_49247,N_41062);
and UO_3863 (O_3863,N_44902,N_42409);
or UO_3864 (O_3864,N_41480,N_41505);
or UO_3865 (O_3865,N_43582,N_44419);
nor UO_3866 (O_3866,N_43397,N_49040);
or UO_3867 (O_3867,N_46774,N_46401);
or UO_3868 (O_3868,N_44907,N_48265);
nor UO_3869 (O_3869,N_49103,N_49969);
nor UO_3870 (O_3870,N_42097,N_46345);
or UO_3871 (O_3871,N_41092,N_40924);
xor UO_3872 (O_3872,N_40383,N_41625);
and UO_3873 (O_3873,N_42578,N_41080);
or UO_3874 (O_3874,N_42457,N_43126);
nand UO_3875 (O_3875,N_42611,N_43673);
or UO_3876 (O_3876,N_47774,N_46151);
nor UO_3877 (O_3877,N_43365,N_44481);
or UO_3878 (O_3878,N_46726,N_41722);
xor UO_3879 (O_3879,N_41678,N_42572);
xnor UO_3880 (O_3880,N_44731,N_40469);
and UO_3881 (O_3881,N_43942,N_40818);
xnor UO_3882 (O_3882,N_42841,N_44342);
xnor UO_3883 (O_3883,N_46507,N_46372);
nand UO_3884 (O_3884,N_42360,N_43849);
xor UO_3885 (O_3885,N_43431,N_45284);
nor UO_3886 (O_3886,N_47465,N_42253);
or UO_3887 (O_3887,N_46016,N_41845);
and UO_3888 (O_3888,N_40826,N_42267);
nor UO_3889 (O_3889,N_45312,N_42575);
or UO_3890 (O_3890,N_46026,N_43103);
xnor UO_3891 (O_3891,N_44230,N_43381);
xnor UO_3892 (O_3892,N_41673,N_47531);
or UO_3893 (O_3893,N_49889,N_41349);
xor UO_3894 (O_3894,N_49056,N_44626);
xnor UO_3895 (O_3895,N_46586,N_45915);
xnor UO_3896 (O_3896,N_47128,N_47893);
nand UO_3897 (O_3897,N_42740,N_47305);
xnor UO_3898 (O_3898,N_42407,N_40005);
or UO_3899 (O_3899,N_45550,N_42292);
nor UO_3900 (O_3900,N_45611,N_47134);
xnor UO_3901 (O_3901,N_47534,N_42983);
or UO_3902 (O_3902,N_46448,N_44708);
nand UO_3903 (O_3903,N_46577,N_44635);
nand UO_3904 (O_3904,N_41716,N_49015);
or UO_3905 (O_3905,N_49085,N_42342);
nand UO_3906 (O_3906,N_46207,N_44001);
xnor UO_3907 (O_3907,N_40033,N_46713);
and UO_3908 (O_3908,N_49766,N_40692);
xor UO_3909 (O_3909,N_46423,N_49293);
and UO_3910 (O_3910,N_43300,N_48835);
or UO_3911 (O_3911,N_45540,N_49007);
xor UO_3912 (O_3912,N_46348,N_41275);
nand UO_3913 (O_3913,N_47812,N_46892);
or UO_3914 (O_3914,N_48925,N_47370);
xnor UO_3915 (O_3915,N_43889,N_45786);
nand UO_3916 (O_3916,N_48500,N_44536);
and UO_3917 (O_3917,N_44980,N_40395);
xnor UO_3918 (O_3918,N_43693,N_48261);
and UO_3919 (O_3919,N_46779,N_44723);
xor UO_3920 (O_3920,N_42867,N_44841);
or UO_3921 (O_3921,N_41461,N_49003);
or UO_3922 (O_3922,N_40305,N_47216);
nand UO_3923 (O_3923,N_48805,N_48726);
nand UO_3924 (O_3924,N_47844,N_48313);
and UO_3925 (O_3925,N_41946,N_49275);
xor UO_3926 (O_3926,N_45144,N_46181);
or UO_3927 (O_3927,N_48404,N_48940);
and UO_3928 (O_3928,N_49358,N_43843);
or UO_3929 (O_3929,N_47037,N_41512);
and UO_3930 (O_3930,N_46094,N_43319);
nand UO_3931 (O_3931,N_41894,N_44755);
nor UO_3932 (O_3932,N_47630,N_43274);
xor UO_3933 (O_3933,N_46329,N_48757);
nor UO_3934 (O_3934,N_44423,N_45606);
xnor UO_3935 (O_3935,N_41616,N_44438);
xor UO_3936 (O_3936,N_40962,N_46594);
nand UO_3937 (O_3937,N_46844,N_49262);
and UO_3938 (O_3938,N_45887,N_40124);
xor UO_3939 (O_3939,N_40822,N_42987);
and UO_3940 (O_3940,N_44826,N_45638);
nand UO_3941 (O_3941,N_40696,N_48300);
xor UO_3942 (O_3942,N_43631,N_42436);
xnor UO_3943 (O_3943,N_42527,N_41788);
nor UO_3944 (O_3944,N_44498,N_48161);
nor UO_3945 (O_3945,N_45101,N_44241);
and UO_3946 (O_3946,N_46855,N_47301);
or UO_3947 (O_3947,N_44819,N_47684);
or UO_3948 (O_3948,N_49146,N_44407);
nand UO_3949 (O_3949,N_40275,N_45642);
and UO_3950 (O_3950,N_40266,N_48187);
xnor UO_3951 (O_3951,N_42637,N_45671);
nor UO_3952 (O_3952,N_48453,N_46615);
nand UO_3953 (O_3953,N_43639,N_44193);
or UO_3954 (O_3954,N_41515,N_40226);
xor UO_3955 (O_3955,N_43938,N_40136);
xor UO_3956 (O_3956,N_45301,N_42393);
nor UO_3957 (O_3957,N_43960,N_44850);
nand UO_3958 (O_3958,N_48648,N_47552);
or UO_3959 (O_3959,N_44066,N_43277);
and UO_3960 (O_3960,N_46995,N_44789);
and UO_3961 (O_3961,N_45766,N_49530);
and UO_3962 (O_3962,N_46394,N_48155);
and UO_3963 (O_3963,N_47698,N_41041);
or UO_3964 (O_3964,N_43149,N_42325);
xnor UO_3965 (O_3965,N_42008,N_48565);
nor UO_3966 (O_3966,N_49062,N_40247);
or UO_3967 (O_3967,N_43433,N_49261);
and UO_3968 (O_3968,N_45080,N_41237);
or UO_3969 (O_3969,N_41696,N_45267);
xnor UO_3970 (O_3970,N_49585,N_40253);
nand UO_3971 (O_3971,N_49562,N_48363);
and UO_3972 (O_3972,N_44337,N_41016);
xor UO_3973 (O_3973,N_44489,N_48498);
nand UO_3974 (O_3974,N_44798,N_47658);
nor UO_3975 (O_3975,N_43947,N_43570);
xnor UO_3976 (O_3976,N_45912,N_40330);
xor UO_3977 (O_3977,N_43484,N_42449);
nand UO_3978 (O_3978,N_41327,N_44359);
nand UO_3979 (O_3979,N_42344,N_48127);
and UO_3980 (O_3980,N_47311,N_48170);
xnor UO_3981 (O_3981,N_44157,N_45222);
nor UO_3982 (O_3982,N_49705,N_44611);
nand UO_3983 (O_3983,N_47667,N_44188);
nand UO_3984 (O_3984,N_49353,N_44004);
or UO_3985 (O_3985,N_44158,N_43475);
or UO_3986 (O_3986,N_47424,N_41202);
and UO_3987 (O_3987,N_46251,N_40309);
nor UO_3988 (O_3988,N_48393,N_45754);
or UO_3989 (O_3989,N_43986,N_46002);
or UO_3990 (O_3990,N_45231,N_41155);
nand UO_3991 (O_3991,N_49648,N_46402);
or UO_3992 (O_3992,N_43974,N_47602);
xor UO_3993 (O_3993,N_46466,N_40252);
nor UO_3994 (O_3994,N_48173,N_47657);
nand UO_3995 (O_3995,N_48380,N_44368);
nand UO_3996 (O_3996,N_49335,N_42956);
or UO_3997 (O_3997,N_46973,N_44516);
xor UO_3998 (O_3998,N_48985,N_43575);
nor UO_3999 (O_3999,N_42014,N_47890);
or UO_4000 (O_4000,N_47051,N_48467);
xnor UO_4001 (O_4001,N_45467,N_45784);
nor UO_4002 (O_4002,N_47568,N_47222);
and UO_4003 (O_4003,N_49837,N_41044);
or UO_4004 (O_4004,N_42924,N_42584);
and UO_4005 (O_4005,N_41422,N_44780);
nor UO_4006 (O_4006,N_47504,N_48557);
xor UO_4007 (O_4007,N_45421,N_49963);
nor UO_4008 (O_4008,N_49029,N_40455);
nor UO_4009 (O_4009,N_49651,N_42952);
nand UO_4010 (O_4010,N_41956,N_42074);
xnor UO_4011 (O_4011,N_40288,N_46121);
xor UO_4012 (O_4012,N_40181,N_42364);
or UO_4013 (O_4013,N_47331,N_44273);
nor UO_4014 (O_4014,N_40329,N_45992);
and UO_4015 (O_4015,N_43500,N_49887);
or UO_4016 (O_4016,N_44365,N_42319);
nor UO_4017 (O_4017,N_41648,N_49215);
nand UO_4018 (O_4018,N_43902,N_49716);
xor UO_4019 (O_4019,N_45825,N_45030);
or UO_4020 (O_4020,N_46245,N_42656);
xor UO_4021 (O_4021,N_44304,N_43985);
nor UO_4022 (O_4022,N_45441,N_49764);
and UO_4023 (O_4023,N_47407,N_44816);
nor UO_4024 (O_4024,N_40016,N_40189);
xor UO_4025 (O_4025,N_41751,N_46503);
and UO_4026 (O_4026,N_44503,N_45259);
nand UO_4027 (O_4027,N_44771,N_41804);
nand UO_4028 (O_4028,N_43870,N_47159);
or UO_4029 (O_4029,N_41790,N_43297);
xor UO_4030 (O_4030,N_44565,N_47373);
xnor UO_4031 (O_4031,N_47951,N_49891);
xnor UO_4032 (O_4032,N_44726,N_42069);
and UO_4033 (O_4033,N_44306,N_43948);
nor UO_4034 (O_4034,N_47631,N_45980);
or UO_4035 (O_4035,N_45178,N_46508);
nand UO_4036 (O_4036,N_45886,N_46826);
nand UO_4037 (O_4037,N_44676,N_41304);
and UO_4038 (O_4038,N_41287,N_46476);
nor UO_4039 (O_4039,N_44085,N_42624);
xor UO_4040 (O_4040,N_41528,N_41358);
nor UO_4041 (O_4041,N_49171,N_47217);
nand UO_4042 (O_4042,N_43134,N_40869);
nor UO_4043 (O_4043,N_42898,N_40682);
nand UO_4044 (O_4044,N_43607,N_40956);
xor UO_4045 (O_4045,N_42903,N_44069);
nand UO_4046 (O_4046,N_40172,N_40456);
or UO_4047 (O_4047,N_42760,N_49304);
xor UO_4048 (O_4048,N_42807,N_48057);
nand UO_4049 (O_4049,N_40616,N_47264);
and UO_4050 (O_4050,N_44172,N_44739);
nand UO_4051 (O_4051,N_40460,N_46309);
xnor UO_4052 (O_4052,N_49069,N_41918);
and UO_4053 (O_4053,N_49264,N_44305);
xor UO_4054 (O_4054,N_48191,N_41875);
xnor UO_4055 (O_4055,N_46527,N_47600);
or UO_4056 (O_4056,N_43637,N_41086);
and UO_4057 (O_4057,N_43141,N_46708);
and UO_4058 (O_4058,N_48290,N_47769);
nand UO_4059 (O_4059,N_45928,N_45596);
nand UO_4060 (O_4060,N_49412,N_42128);
and UO_4061 (O_4061,N_48560,N_46550);
nand UO_4062 (O_4062,N_44641,N_48224);
xnor UO_4063 (O_4063,N_41109,N_49853);
or UO_4064 (O_4064,N_49326,N_47963);
and UO_4065 (O_4065,N_42667,N_49517);
xor UO_4066 (O_4066,N_44492,N_48010);
or UO_4067 (O_4067,N_40767,N_49157);
nand UO_4068 (O_4068,N_47880,N_42641);
xnor UO_4069 (O_4069,N_43015,N_48741);
nand UO_4070 (O_4070,N_49840,N_49527);
and UO_4071 (O_4071,N_42809,N_42354);
nand UO_4072 (O_4072,N_44754,N_40454);
nand UO_4073 (O_4073,N_49319,N_47452);
or UO_4074 (O_4074,N_48163,N_45038);
and UO_4075 (O_4075,N_43258,N_41537);
xnor UO_4076 (O_4076,N_45551,N_41557);
nand UO_4077 (O_4077,N_43382,N_47646);
or UO_4078 (O_4078,N_46879,N_49377);
and UO_4079 (O_4079,N_49101,N_45223);
xor UO_4080 (O_4080,N_42408,N_43705);
or UO_4081 (O_4081,N_43773,N_45156);
xnor UO_4082 (O_4082,N_43394,N_42534);
nor UO_4083 (O_4083,N_41697,N_41009);
and UO_4084 (O_4084,N_45703,N_46504);
and UO_4085 (O_4085,N_45833,N_43629);
or UO_4086 (O_4086,N_44922,N_47357);
and UO_4087 (O_4087,N_45389,N_40854);
nor UO_4088 (O_4088,N_48110,N_42976);
and UO_4089 (O_4089,N_48740,N_40482);
xor UO_4090 (O_4090,N_49691,N_44009);
nor UO_4091 (O_4091,N_40864,N_41540);
or UO_4092 (O_4092,N_40139,N_41940);
nand UO_4093 (O_4093,N_44526,N_43488);
nand UO_4094 (O_4094,N_43106,N_48146);
and UO_4095 (O_4095,N_41140,N_43795);
xor UO_4096 (O_4096,N_49396,N_42516);
xnor UO_4097 (O_4097,N_49244,N_47926);
nor UO_4098 (O_4098,N_46198,N_40999);
or UO_4099 (O_4099,N_44961,N_43335);
nor UO_4100 (O_4100,N_43634,N_42942);
xnor UO_4101 (O_4101,N_42210,N_44774);
nor UO_4102 (O_4102,N_47809,N_41533);
nor UO_4103 (O_4103,N_48266,N_46252);
nand UO_4104 (O_4104,N_43989,N_41127);
and UO_4105 (O_4105,N_46622,N_49553);
nand UO_4106 (O_4106,N_48678,N_46147);
nand UO_4107 (O_4107,N_42926,N_44615);
xor UO_4108 (O_4108,N_48225,N_42269);
nand UO_4109 (O_4109,N_45950,N_43259);
xor UO_4110 (O_4110,N_47681,N_40445);
nor UO_4111 (O_4111,N_44905,N_45228);
nor UO_4112 (O_4112,N_49132,N_44076);
nand UO_4113 (O_4113,N_46463,N_48681);
nor UO_4114 (O_4114,N_40463,N_41994);
nor UO_4115 (O_4115,N_49750,N_49639);
nor UO_4116 (O_4116,N_47014,N_43480);
xnor UO_4117 (O_4117,N_49791,N_49874);
and UO_4118 (O_4118,N_40670,N_43816);
nand UO_4119 (O_4119,N_41150,N_47870);
nand UO_4120 (O_4120,N_48613,N_46884);
or UO_4121 (O_4121,N_45476,N_45869);
and UO_4122 (O_4122,N_47475,N_49935);
and UO_4123 (O_4123,N_42164,N_43371);
nor UO_4124 (O_4124,N_43920,N_48721);
or UO_4125 (O_4125,N_42322,N_44149);
and UO_4126 (O_4126,N_49602,N_40296);
and UO_4127 (O_4127,N_44512,N_47309);
xor UO_4128 (O_4128,N_45729,N_43862);
xor UO_4129 (O_4129,N_42406,N_47150);
or UO_4130 (O_4130,N_46919,N_44343);
xor UO_4131 (O_4131,N_45942,N_41969);
xnor UO_4132 (O_4132,N_40833,N_49051);
and UO_4133 (O_4133,N_47620,N_41615);
or UO_4134 (O_4134,N_43218,N_47043);
or UO_4135 (O_4135,N_48956,N_41548);
or UO_4136 (O_4136,N_48033,N_47648);
and UO_4137 (O_4137,N_46313,N_43320);
nor UO_4138 (O_4138,N_44238,N_41186);
nand UO_4139 (O_4139,N_45076,N_44222);
nand UO_4140 (O_4140,N_44115,N_46808);
or UO_4141 (O_4141,N_49450,N_45732);
and UO_4142 (O_4142,N_46793,N_49729);
and UO_4143 (O_4143,N_44071,N_41176);
and UO_4144 (O_4144,N_40878,N_43770);
nor UO_4145 (O_4145,N_42089,N_49182);
nor UO_4146 (O_4146,N_46249,N_44908);
nand UO_4147 (O_4147,N_45346,N_43528);
nor UO_4148 (O_4148,N_45795,N_43220);
and UO_4149 (O_4149,N_45164,N_44147);
nor UO_4150 (O_4150,N_49539,N_43614);
xnor UO_4151 (O_4151,N_40790,N_45165);
xor UO_4152 (O_4152,N_44760,N_43176);
nor UO_4153 (O_4153,N_46670,N_46811);
nor UO_4154 (O_4154,N_40689,N_41273);
nand UO_4155 (O_4155,N_46533,N_49908);
and UO_4156 (O_4156,N_40708,N_43315);
and UO_4157 (O_4157,N_49266,N_47930);
or UO_4158 (O_4158,N_45592,N_46628);
or UO_4159 (O_4159,N_48965,N_40236);
and UO_4160 (O_4160,N_48058,N_47316);
xnor UO_4161 (O_4161,N_41249,N_48072);
or UO_4162 (O_4162,N_43063,N_43911);
and UO_4163 (O_4163,N_42525,N_44011);
xor UO_4164 (O_4164,N_48760,N_48082);
or UO_4165 (O_4165,N_47318,N_43053);
nor UO_4166 (O_4166,N_47682,N_43078);
nor UO_4167 (O_4167,N_45991,N_47590);
nor UO_4168 (O_4168,N_48488,N_46057);
or UO_4169 (O_4169,N_45173,N_40697);
xor UO_4170 (O_4170,N_42189,N_40580);
or UO_4171 (O_4171,N_44552,N_49551);
nand UO_4172 (O_4172,N_45232,N_41968);
xnor UO_4173 (O_4173,N_40323,N_40811);
and UO_4174 (O_4174,N_42522,N_41051);
or UO_4175 (O_4175,N_47567,N_49074);
nor UO_4176 (O_4176,N_49294,N_45409);
nand UO_4177 (O_4177,N_46709,N_44078);
xnor UO_4178 (O_4178,N_46475,N_46560);
and UO_4179 (O_4179,N_44683,N_49368);
and UO_4180 (O_4180,N_49725,N_47535);
and UO_4181 (O_4181,N_49845,N_48624);
nor UO_4182 (O_4182,N_49899,N_45576);
nor UO_4183 (O_4183,N_49495,N_40102);
and UO_4184 (O_4184,N_47383,N_42017);
xor UO_4185 (O_4185,N_41440,N_49567);
xnor UO_4186 (O_4186,N_42892,N_44227);
nand UO_4187 (O_4187,N_47763,N_42038);
xnor UO_4188 (O_4188,N_49930,N_47687);
xnor UO_4189 (O_4189,N_48320,N_44855);
or UO_4190 (O_4190,N_47818,N_43821);
xnor UO_4191 (O_4191,N_45382,N_43973);
or UO_4192 (O_4192,N_47747,N_42430);
nand UO_4193 (O_4193,N_43020,N_41309);
nor UO_4194 (O_4194,N_40662,N_45538);
nor UO_4195 (O_4195,N_40126,N_45404);
nand UO_4196 (O_4196,N_44973,N_47819);
nand UO_4197 (O_4197,N_49491,N_40387);
nand UO_4198 (O_4198,N_42007,N_48545);
nor UO_4199 (O_4199,N_46601,N_41757);
or UO_4200 (O_4200,N_44815,N_42482);
or UO_4201 (O_4201,N_48663,N_46832);
or UO_4202 (O_4202,N_44042,N_45932);
or UO_4203 (O_4203,N_48374,N_43801);
nand UO_4204 (O_4204,N_47471,N_40903);
and UO_4205 (O_4205,N_40475,N_40076);
and UO_4206 (O_4206,N_44370,N_42580);
nand UO_4207 (O_4207,N_48731,N_47958);
nand UO_4208 (O_4208,N_49762,N_40749);
xnor UO_4209 (O_4209,N_49801,N_45569);
xor UO_4210 (O_4210,N_41846,N_42726);
xor UO_4211 (O_4211,N_46290,N_45326);
and UO_4212 (O_4212,N_43030,N_40526);
nor UO_4213 (O_4213,N_48245,N_48126);
xor UO_4214 (O_4214,N_41911,N_46685);
or UO_4215 (O_4215,N_47439,N_49593);
xor UO_4216 (O_4216,N_41595,N_40894);
and UO_4217 (O_4217,N_46773,N_45493);
nor UO_4218 (O_4218,N_42945,N_40520);
xor UO_4219 (O_4219,N_40577,N_48494);
nand UO_4220 (O_4220,N_48183,N_47174);
nand UO_4221 (O_4221,N_49947,N_40665);
nor UO_4222 (O_4222,N_46455,N_43370);
or UO_4223 (O_4223,N_46828,N_49437);
and UO_4224 (O_4224,N_49298,N_47437);
xor UO_4225 (O_4225,N_45755,N_40188);
nor UO_4226 (O_4226,N_47834,N_46390);
xor UO_4227 (O_4227,N_43113,N_45416);
and UO_4228 (O_4228,N_40429,N_45047);
or UO_4229 (O_4229,N_40187,N_46936);
nand UO_4230 (O_4230,N_43542,N_43314);
xor UO_4231 (O_4231,N_48200,N_47399);
or UO_4232 (O_4232,N_46334,N_43344);
nand UO_4233 (O_4233,N_47533,N_40248);
nand UO_4234 (O_4234,N_48287,N_47485);
xor UO_4235 (O_4235,N_44496,N_46905);
nor UO_4236 (O_4236,N_45129,N_44743);
nand UO_4237 (O_4237,N_45190,N_41501);
xor UO_4238 (O_4238,N_47106,N_40173);
or UO_4239 (O_4239,N_46684,N_48700);
nor UO_4240 (O_4240,N_41384,N_46090);
or UO_4241 (O_4241,N_47474,N_41876);
xnor UO_4242 (O_4242,N_46176,N_42154);
or UO_4243 (O_4243,N_44415,N_43117);
nand UO_4244 (O_4244,N_40286,N_40153);
and UO_4245 (O_4245,N_43937,N_40481);
or UO_4246 (O_4246,N_45027,N_47225);
nor UO_4247 (O_4247,N_44080,N_46847);
nand UO_4248 (O_4248,N_40889,N_49582);
and UO_4249 (O_4249,N_42386,N_41394);
nand UO_4250 (O_4250,N_47688,N_49351);
nor UO_4251 (O_4251,N_43748,N_48876);
nand UO_4252 (O_4252,N_48044,N_41108);
xnor UO_4253 (O_4253,N_48599,N_43301);
and UO_4254 (O_4254,N_43180,N_48446);
nor UO_4255 (O_4255,N_49299,N_41387);
or UO_4256 (O_4256,N_42557,N_40939);
nor UO_4257 (O_4257,N_41554,N_40963);
or UO_4258 (O_4258,N_42620,N_40061);
xnor UO_4259 (O_4259,N_44187,N_40038);
nand UO_4260 (O_4260,N_42347,N_42710);
nor UO_4261 (O_4261,N_47292,N_45011);
nor UO_4262 (O_4262,N_49724,N_40267);
or UO_4263 (O_4263,N_47207,N_40426);
nand UO_4264 (O_4264,N_44801,N_45522);
and UO_4265 (O_4265,N_42576,N_41520);
and UO_4266 (O_4266,N_47045,N_49735);
or UO_4267 (O_4267,N_48075,N_49420);
or UO_4268 (O_4268,N_48848,N_47574);
and UO_4269 (O_4269,N_42110,N_49186);
xor UO_4270 (O_4270,N_41747,N_46935);
xnor UO_4271 (O_4271,N_45319,N_45941);
nand UO_4272 (O_4272,N_43490,N_42973);
nand UO_4273 (O_4273,N_42645,N_43599);
nand UO_4274 (O_4274,N_40715,N_43978);
or UO_4275 (O_4275,N_44510,N_41626);
and UO_4276 (O_4276,N_41409,N_49726);
or UO_4277 (O_4277,N_41164,N_41584);
xnor UO_4278 (O_4278,N_43420,N_48281);
nor UO_4279 (O_4279,N_49627,N_40819);
nand UO_4280 (O_4280,N_49929,N_40297);
or UO_4281 (O_4281,N_49613,N_41043);
xor UO_4282 (O_4282,N_42220,N_40568);
nand UO_4283 (O_4283,N_48537,N_46909);
nor UO_4284 (O_4284,N_49701,N_40047);
xor UO_4285 (O_4285,N_48451,N_42970);
and UO_4286 (O_4286,N_40298,N_44882);
or UO_4287 (O_4287,N_45206,N_41323);
or UO_4288 (O_4288,N_43341,N_42765);
nor UO_4289 (O_4289,N_48348,N_44234);
nand UO_4290 (O_4290,N_45937,N_46593);
nand UO_4291 (O_4291,N_47651,N_43893);
nand UO_4292 (O_4292,N_41707,N_40119);
xor UO_4293 (O_4293,N_49213,N_48185);
or UO_4294 (O_4294,N_43231,N_49064);
or UO_4295 (O_4295,N_48388,N_47627);
xnor UO_4296 (O_4296,N_48004,N_49642);
xor UO_4297 (O_4297,N_42417,N_47909);
and UO_4298 (O_4298,N_42772,N_42192);
nand UO_4299 (O_4299,N_47699,N_44392);
nand UO_4300 (O_4300,N_46979,N_46086);
and UO_4301 (O_4301,N_42536,N_45523);
nor UO_4302 (O_4302,N_41427,N_44245);
and UO_4303 (O_4303,N_40191,N_45398);
and UO_4304 (O_4304,N_46921,N_42174);
or UO_4305 (O_4305,N_40983,N_47922);
or UO_4306 (O_4306,N_46799,N_47107);
or UO_4307 (O_4307,N_41001,N_44079);
nand UO_4308 (O_4308,N_47189,N_46487);
nand UO_4309 (O_4309,N_40152,N_47734);
nand UO_4310 (O_4310,N_49752,N_46894);
nand UO_4311 (O_4311,N_42568,N_45361);
and UO_4312 (O_4312,N_40314,N_42738);
xnor UO_4313 (O_4313,N_45146,N_40246);
and UO_4314 (O_4314,N_43853,N_47901);
nor UO_4315 (O_4315,N_40642,N_45025);
nand UO_4316 (O_4316,N_48479,N_40240);
and UO_4317 (O_4317,N_45558,N_44707);
nand UO_4318 (O_4318,N_47009,N_42317);
and UO_4319 (O_4319,N_48598,N_42949);
xnor UO_4320 (O_4320,N_44574,N_45532);
or UO_4321 (O_4321,N_41798,N_40862);
or UO_4322 (O_4322,N_44702,N_45565);
nand UO_4323 (O_4323,N_45600,N_42234);
nand UO_4324 (O_4324,N_47164,N_43697);
and UO_4325 (O_4325,N_45334,N_46126);
or UO_4326 (O_4326,N_44583,N_44424);
nor UO_4327 (O_4327,N_46690,N_43024);
nand UO_4328 (O_4328,N_40947,N_46736);
or UO_4329 (O_4329,N_49438,N_43618);
xor UO_4330 (O_4330,N_41268,N_40466);
and UO_4331 (O_4331,N_47815,N_48456);
and UO_4332 (O_4332,N_44458,N_41403);
xor UO_4333 (O_4333,N_47775,N_42729);
nor UO_4334 (O_4334,N_42208,N_45895);
xor UO_4335 (O_4335,N_44610,N_47417);
nor UO_4336 (O_4336,N_45918,N_45195);
nand UO_4337 (O_4337,N_40134,N_46242);
and UO_4338 (O_4338,N_42828,N_48198);
nand UO_4339 (O_4339,N_40004,N_41657);
nor UO_4340 (O_4340,N_49095,N_47588);
and UO_4341 (O_4341,N_43833,N_41173);
or UO_4342 (O_4342,N_42338,N_45224);
nor UO_4343 (O_4343,N_41967,N_42188);
nor UO_4344 (O_4344,N_45119,N_40443);
xor UO_4345 (O_4345,N_42518,N_48116);
nand UO_4346 (O_4346,N_43606,N_45443);
or UO_4347 (O_4347,N_49688,N_49637);
xnor UO_4348 (O_4348,N_49121,N_43731);
xor UO_4349 (O_4349,N_49507,N_41878);
and UO_4350 (O_4350,N_45567,N_41295);
and UO_4351 (O_4351,N_46349,N_48574);
xor UO_4352 (O_4352,N_48745,N_49835);
nor UO_4353 (O_4353,N_42018,N_42484);
xnor UO_4354 (O_4354,N_42217,N_43781);
nand UO_4355 (O_4355,N_40294,N_43331);
and UO_4356 (O_4356,N_47136,N_49821);
nand UO_4357 (O_4357,N_44247,N_49108);
nand UO_4358 (O_4358,N_42786,N_42957);
nand UO_4359 (O_4359,N_42255,N_46824);
and UO_4360 (O_4360,N_44341,N_42483);
and UO_4361 (O_4361,N_45099,N_49463);
or UO_4362 (O_4362,N_49572,N_49505);
nor UO_4363 (O_4363,N_40610,N_45037);
nand UO_4364 (O_4364,N_41203,N_46228);
or UO_4365 (O_4365,N_41431,N_46032);
nor UO_4366 (O_4366,N_44605,N_40348);
xnor UO_4367 (O_4367,N_46872,N_46113);
nor UO_4368 (O_4368,N_49739,N_46434);
nand UO_4369 (O_4369,N_46118,N_44851);
nand UO_4370 (O_4370,N_41886,N_47521);
and UO_4371 (O_4371,N_42999,N_48013);
and UO_4372 (O_4372,N_42775,N_45368);
nor UO_4373 (O_4373,N_41800,N_40315);
or UO_4374 (O_4374,N_41130,N_47221);
nor UO_4375 (O_4375,N_42981,N_46128);
xnor UO_4376 (O_4376,N_44369,N_45700);
and UO_4377 (O_4377,N_42395,N_47232);
nor UO_4378 (O_4378,N_42820,N_49564);
or UO_4379 (O_4379,N_44250,N_43812);
nor UO_4380 (O_4380,N_44122,N_46003);
and UO_4381 (O_4381,N_45818,N_45020);
or UO_4382 (O_4382,N_41134,N_49638);
or UO_4383 (O_4383,N_46859,N_43845);
and UO_4384 (O_4384,N_41370,N_46530);
nor UO_4385 (O_4385,N_45358,N_41544);
xor UO_4386 (O_4386,N_43092,N_47259);
nand UO_4387 (O_4387,N_49698,N_42885);
nor UO_4388 (O_4388,N_40379,N_41541);
or UO_4389 (O_4389,N_43604,N_43501);
nand UO_4390 (O_4390,N_49329,N_45583);
xor UO_4391 (O_4391,N_43675,N_48675);
nor UO_4392 (O_4392,N_48343,N_40352);
xnor UO_4393 (O_4393,N_48394,N_42721);
nand UO_4394 (O_4394,N_46095,N_47849);
xor UO_4395 (O_4395,N_45556,N_44761);
nor UO_4396 (O_4396,N_49355,N_45662);
nand UO_4397 (O_4397,N_48994,N_47984);
nor UO_4398 (O_4398,N_46441,N_41269);
nand UO_4399 (O_4399,N_45507,N_47239);
nand UO_4400 (O_4400,N_44502,N_46866);
nand UO_4401 (O_4401,N_40184,N_47269);
or UO_4402 (O_4402,N_46135,N_48901);
nor UO_4403 (O_4403,N_48341,N_41829);
and UO_4404 (O_4404,N_41732,N_43442);
xor UO_4405 (O_4405,N_45503,N_40537);
nand UO_4406 (O_4406,N_47163,N_47152);
nand UO_4407 (O_4407,N_48099,N_46084);
nor UO_4408 (O_4408,N_41739,N_45650);
nor UO_4409 (O_4409,N_49082,N_45660);
nor UO_4410 (O_4410,N_47660,N_45357);
nand UO_4411 (O_4411,N_42532,N_47220);
or UO_4412 (O_4412,N_48483,N_45459);
xor UO_4413 (O_4413,N_44412,N_47033);
or UO_4414 (O_4414,N_47185,N_41631);
nand UO_4415 (O_4415,N_42313,N_40721);
and UO_4416 (O_4416,N_48386,N_44207);
xor UO_4417 (O_4417,N_45393,N_44804);
nand UO_4418 (O_4418,N_47962,N_43436);
and UO_4419 (O_4419,N_46585,N_46462);
and UO_4420 (O_4420,N_43694,N_43302);
nand UO_4421 (O_4421,N_47335,N_49550);
or UO_4422 (O_4422,N_47689,N_43084);
nor UO_4423 (O_4423,N_44811,N_44915);
and UO_4424 (O_4424,N_42529,N_43615);
xnor UO_4425 (O_4425,N_47607,N_49386);
and UO_4426 (O_4426,N_44976,N_41907);
or UO_4427 (O_4427,N_40795,N_41094);
or UO_4428 (O_4428,N_42411,N_46734);
nor UO_4429 (O_4429,N_49016,N_40223);
xnor UO_4430 (O_4430,N_42581,N_44039);
and UO_4431 (O_4431,N_44141,N_42823);
xnor UO_4432 (O_4432,N_44970,N_40845);
nand UO_4433 (O_4433,N_44783,N_45042);
and UO_4434 (O_4434,N_42764,N_49014);
nand UO_4435 (O_4435,N_45388,N_48990);
nand UO_4436 (O_4436,N_40560,N_42506);
nor UO_4437 (O_4437,N_42569,N_49414);
or UO_4438 (O_4438,N_48111,N_48632);
or UO_4439 (O_4439,N_47934,N_46792);
nand UO_4440 (O_4440,N_43796,N_46398);
and UO_4441 (O_4441,N_43743,N_42857);
nand UO_4442 (O_4442,N_48525,N_41666);
or UO_4443 (O_4443,N_44242,N_46360);
xnor UO_4444 (O_4444,N_46572,N_43984);
or UO_4445 (O_4445,N_43539,N_45225);
or UO_4446 (O_4446,N_45273,N_43378);
nor UO_4447 (O_4447,N_40533,N_47469);
nand UO_4448 (O_4448,N_46437,N_46679);
and UO_4449 (O_4449,N_47519,N_46624);
nor UO_4450 (O_4450,N_46385,N_46613);
xnor UO_4451 (O_4451,N_47199,N_43267);
and UO_4452 (O_4452,N_44991,N_48308);
nor UO_4453 (O_4453,N_46214,N_44894);
xnor UO_4454 (O_4454,N_49883,N_40703);
nand UO_4455 (O_4455,N_42416,N_49434);
nor UO_4456 (O_4456,N_43912,N_47942);
and UO_4457 (O_4457,N_44023,N_41769);
nor UO_4458 (O_4458,N_43493,N_46421);
or UO_4459 (O_4459,N_41717,N_46478);
nor UO_4460 (O_4460,N_46571,N_45100);
xor UO_4461 (O_4461,N_45068,N_47982);
xor UO_4462 (O_4462,N_45056,N_46124);
and UO_4463 (O_4463,N_41418,N_43109);
and UO_4464 (O_4464,N_44963,N_46157);
and UO_4465 (O_4465,N_43517,N_47081);
and UO_4466 (O_4466,N_43690,N_47772);
or UO_4467 (O_4467,N_40639,N_49684);
nand UO_4468 (O_4468,N_42571,N_49928);
nand UO_4469 (O_4469,N_48556,N_42936);
xnor UO_4470 (O_4470,N_40908,N_40510);
nor UO_4471 (O_4471,N_45678,N_49272);
or UO_4472 (O_4472,N_43594,N_42107);
nor UO_4473 (O_4473,N_42196,N_40072);
xor UO_4474 (O_4474,N_44740,N_41608);
or UO_4475 (O_4475,N_45494,N_40677);
and UO_4476 (O_4476,N_40059,N_46814);
xor UO_4477 (O_4477,N_43823,N_43580);
nand UO_4478 (O_4478,N_41209,N_40711);
and UO_4479 (O_4479,N_41449,N_45269);
or UO_4480 (O_4480,N_42019,N_40661);
and UO_4481 (O_4481,N_46648,N_49041);
nand UO_4482 (O_4482,N_44658,N_43967);
nor UO_4483 (O_4483,N_42891,N_48318);
and UO_4484 (O_4484,N_48319,N_42758);
nand UO_4485 (O_4485,N_42289,N_49174);
nand UO_4486 (O_4486,N_40228,N_40973);
or UO_4487 (O_4487,N_41036,N_44105);
nand UO_4488 (O_4488,N_49857,N_43196);
or UO_4489 (O_4489,N_49139,N_47506);
and UO_4490 (O_4490,N_46132,N_43983);
xnor UO_4491 (O_4491,N_40562,N_44714);
nand UO_4492 (O_4492,N_42080,N_40109);
xnor UO_4493 (O_4493,N_46185,N_43352);
nor UO_4494 (O_4494,N_40794,N_49488);
nor UO_4495 (O_4495,N_45192,N_45910);
nor UO_4496 (O_4496,N_49024,N_49337);
nor UO_4497 (O_4497,N_42094,N_40393);
or UO_4498 (O_4498,N_40645,N_43265);
nor UO_4499 (O_4499,N_41613,N_48695);
xor UO_4500 (O_4500,N_42912,N_49154);
nand UO_4501 (O_4501,N_47113,N_43727);
xnor UO_4502 (O_4502,N_40003,N_47209);
and UO_4503 (O_4503,N_43645,N_46159);
and UO_4504 (O_4504,N_48486,N_48907);
xnor UO_4505 (O_4505,N_42090,N_44251);
xnor UO_4506 (O_4506,N_49640,N_49931);
and UO_4507 (O_4507,N_43628,N_49493);
nor UO_4508 (O_4508,N_46278,N_44571);
and UO_4509 (O_4509,N_45657,N_42459);
and UO_4510 (O_4510,N_47878,N_46592);
or UO_4511 (O_4511,N_44647,N_48141);
xor UO_4512 (O_4512,N_40700,N_42168);
or UO_4513 (O_4513,N_45500,N_44218);
and UO_4514 (O_4514,N_48476,N_47252);
and UO_4515 (O_4515,N_47961,N_43797);
nor UO_4516 (O_4516,N_48752,N_40780);
xor UO_4517 (O_4517,N_40614,N_47008);
nor UO_4518 (O_4518,N_48417,N_42261);
nand UO_4519 (O_4519,N_49483,N_42998);
nor UO_4520 (O_4520,N_44357,N_43444);
nand UO_4521 (O_4521,N_47362,N_47409);
xor UO_4522 (O_4522,N_42767,N_47960);
nand UO_4523 (O_4523,N_44939,N_42157);
and UO_4524 (O_4524,N_43530,N_44216);
and UO_4525 (O_4525,N_48978,N_49302);
nand UO_4526 (O_4526,N_41192,N_46561);
nor UO_4527 (O_4527,N_47482,N_40523);
and UO_4528 (O_4528,N_46071,N_40485);
nor UO_4529 (O_4529,N_45511,N_40701);
and UO_4530 (O_4530,N_41566,N_48991);
nand UO_4531 (O_4531,N_40501,N_43913);
nor UO_4532 (O_4532,N_40809,N_47835);
and UO_4533 (O_4533,N_42412,N_46383);
and UO_4534 (O_4534,N_45123,N_41351);
nor UO_4535 (O_4535,N_48977,N_43882);
xor UO_4536 (O_4536,N_44097,N_42876);
nor UO_4537 (O_4537,N_40970,N_42724);
nand UO_4538 (O_4538,N_46236,N_42218);
nand UO_4539 (O_4539,N_44054,N_46540);
and UO_4540 (O_4540,N_44267,N_49961);
or UO_4541 (O_4541,N_49151,N_43788);
xor UO_4542 (O_4542,N_48209,N_47310);
or UO_4543 (O_4543,N_41020,N_42256);
and UO_4544 (O_4544,N_49995,N_48747);
nand UO_4545 (O_4545,N_48461,N_44329);
nand UO_4546 (O_4546,N_44713,N_48949);
nor UO_4547 (O_4547,N_44504,N_49268);
nand UO_4548 (O_4548,N_49901,N_46319);
and UO_4549 (O_4549,N_48744,N_48763);
and UO_4550 (O_4550,N_42022,N_48115);
nor UO_4551 (O_4551,N_42995,N_47948);
xnor UO_4552 (O_4552,N_48880,N_46008);
and UO_4553 (O_4553,N_49650,N_41934);
xor UO_4554 (O_4554,N_41007,N_48694);
xnor UO_4555 (O_4555,N_49116,N_46737);
or UO_4556 (O_4556,N_40130,N_42238);
nand UO_4557 (O_4557,N_48684,N_44933);
or UO_4558 (O_4558,N_49418,N_43306);
nor UO_4559 (O_4559,N_47076,N_49848);
nor UO_4560 (O_4560,N_48842,N_49617);
and UO_4561 (O_4561,N_49100,N_43076);
xnor UO_4562 (O_4562,N_45573,N_45866);
nor UO_4563 (O_4563,N_40255,N_40847);
xnor UO_4564 (O_4564,N_40385,N_46818);
nand UO_4565 (O_4565,N_49196,N_41880);
nand UO_4566 (O_4566,N_47372,N_45376);
nor UO_4567 (O_4567,N_49147,N_46749);
nor UO_4568 (O_4568,N_42247,N_43521);
or UO_4569 (O_4569,N_42402,N_41011);
nor UO_4570 (O_4570,N_42573,N_49680);
or UO_4571 (O_4571,N_45031,N_46021);
or UO_4572 (O_4572,N_42634,N_43410);
nand UO_4573 (O_4573,N_40591,N_48914);
and UO_4574 (O_4574,N_47290,N_41506);
xnor UO_4575 (O_4575,N_46842,N_40652);
and UO_4576 (O_4576,N_46020,N_44281);
xor UO_4577 (O_4577,N_43198,N_46595);
xor UO_4578 (O_4578,N_48759,N_47894);
and UO_4579 (O_4579,N_41434,N_41959);
xor UO_4580 (O_4580,N_49241,N_44983);
and UO_4581 (O_4581,N_48793,N_44601);
nand UO_4582 (O_4582,N_42318,N_40879);
or UO_4583 (O_4583,N_48214,N_49456);
nor UO_4584 (O_4584,N_41354,N_47329);
nor UO_4585 (O_4585,N_44014,N_45652);
nand UO_4586 (O_4586,N_40654,N_46197);
nand UO_4587 (O_4587,N_49955,N_47102);
and UO_4588 (O_4588,N_42076,N_44593);
and UO_4589 (O_4589,N_49894,N_40433);
nor UO_4590 (O_4590,N_43685,N_47974);
nor UO_4591 (O_4591,N_44589,N_42257);
nand UO_4592 (O_4592,N_40346,N_43395);
or UO_4593 (O_4593,N_42792,N_42727);
xor UO_4594 (O_4594,N_44511,N_42653);
nor UO_4595 (O_4595,N_43686,N_46716);
nand UO_4596 (O_4596,N_40000,N_40714);
nor UO_4597 (O_4597,N_43429,N_43636);
or UO_4598 (O_4598,N_45065,N_40075);
nand UO_4599 (O_4599,N_46911,N_42604);
and UO_4600 (O_4600,N_44284,N_47435);
or UO_4601 (O_4601,N_41033,N_40592);
nor UO_4602 (O_4602,N_46786,N_41276);
nand UO_4603 (O_4603,N_44192,N_48927);
xor UO_4604 (O_4604,N_40114,N_42778);
or UO_4605 (O_4605,N_47846,N_46220);
nor UO_4606 (O_4606,N_47459,N_47369);
nor UO_4607 (O_4607,N_45278,N_49306);
or UO_4608 (O_4608,N_46014,N_40536);
xor UO_4609 (O_4609,N_49161,N_45840);
or UO_4610 (O_4610,N_43540,N_41118);
or UO_4611 (O_4611,N_44213,N_40850);
xnor UO_4612 (O_4612,N_49870,N_42746);
nand UO_4613 (O_4613,N_44699,N_43617);
xnor UO_4614 (O_4614,N_48630,N_42864);
nor UO_4615 (O_4615,N_49421,N_40640);
nor UO_4616 (O_4616,N_43546,N_40828);
xnor UO_4617 (O_4617,N_43564,N_40872);
nor UO_4618 (O_4618,N_40997,N_47366);
nand UO_4619 (O_4619,N_48941,N_49481);
and UO_4620 (O_4620,N_45890,N_46314);
xnor UO_4621 (O_4621,N_44854,N_45411);
and UO_4622 (O_4622,N_43269,N_48714);
nor UO_4623 (O_4623,N_48084,N_48635);
xor UO_4624 (O_4624,N_40540,N_49879);
and UO_4625 (O_4625,N_45626,N_46666);
or UO_4626 (O_4626,N_48957,N_42914);
and UO_4627 (O_4627,N_43038,N_40214);
nor UO_4628 (O_4628,N_47621,N_45634);
xor UO_4629 (O_4629,N_46631,N_48002);
or UO_4630 (O_4630,N_47938,N_41735);
nand UO_4631 (O_4631,N_46358,N_42451);
nor UO_4632 (O_4632,N_45741,N_47028);
and UO_4633 (O_4633,N_46254,N_48984);
or UO_4634 (O_4634,N_40531,N_44585);
nor UO_4635 (O_4635,N_49805,N_42334);
nand UO_4636 (O_4636,N_47364,N_45764);
and UO_4637 (O_4637,N_47055,N_40885);
nand UO_4638 (O_4638,N_40612,N_45499);
nor UO_4639 (O_4639,N_40585,N_47524);
nand UO_4640 (O_4640,N_44824,N_43238);
xnor UO_4641 (O_4641,N_49148,N_49240);
nand UO_4642 (O_4642,N_45917,N_42787);
nor UO_4643 (O_4643,N_42209,N_40984);
nor UO_4644 (O_4644,N_45539,N_44240);
and UO_4645 (O_4645,N_44501,N_46280);
and UO_4646 (O_4646,N_43620,N_46672);
and UO_4647 (O_4647,N_40045,N_43775);
and UO_4648 (O_4648,N_48804,N_40105);
nand UO_4649 (O_4649,N_40972,N_44410);
xor UO_4650 (O_4650,N_46247,N_49050);
nor UO_4651 (O_4651,N_41167,N_48649);
and UO_4652 (O_4652,N_48189,N_42697);
nor UO_4653 (O_4653,N_46138,N_43373);
and UO_4654 (O_4654,N_40532,N_44507);
nor UO_4655 (O_4655,N_48095,N_44868);
xor UO_4656 (O_4656,N_48817,N_46759);
xnor UO_4657 (O_4657,N_43721,N_43337);
nand UO_4658 (O_4658,N_41046,N_44020);
nand UO_4659 (O_4659,N_45588,N_47314);
nor UO_4660 (O_4660,N_48032,N_48243);
or UO_4661 (O_4661,N_45881,N_45953);
or UO_4662 (O_4662,N_45646,N_43348);
xnor UO_4663 (O_4663,N_45579,N_40479);
or UO_4664 (O_4664,N_44972,N_47061);
and UO_4665 (O_4665,N_48512,N_46005);
nand UO_4666 (O_4666,N_44375,N_43425);
nor UO_4667 (O_4667,N_44703,N_45617);
xor UO_4668 (O_4668,N_45105,N_40683);
or UO_4669 (O_4669,N_44724,N_46546);
nor UO_4670 (O_4670,N_46557,N_45313);
or UO_4671 (O_4671,N_45194,N_43427);
and UO_4672 (O_4672,N_49284,N_43252);
or UO_4673 (O_4673,N_47759,N_43950);
nor UO_4674 (O_4674,N_46216,N_40897);
nand UO_4675 (O_4675,N_49917,N_47231);
nand UO_4676 (O_4676,N_49727,N_45006);
nor UO_4677 (O_4677,N_49250,N_42899);
nand UO_4678 (O_4678,N_46668,N_49002);
nand UO_4679 (O_4679,N_49332,N_41962);
nand UO_4680 (O_4680,N_45492,N_43254);
nand UO_4681 (O_4681,N_48361,N_46300);
or UO_4682 (O_4682,N_47096,N_43136);
nand UO_4683 (O_4683,N_43655,N_40846);
or UO_4684 (O_4684,N_45423,N_42284);
xnor UO_4685 (O_4685,N_48913,N_41250);
or UO_4686 (O_4686,N_44243,N_49771);
or UO_4687 (O_4687,N_40358,N_43512);
or UO_4688 (O_4688,N_47514,N_41958);
xnor UO_4689 (O_4689,N_44746,N_42415);
and UO_4690 (O_4690,N_48503,N_41760);
and UO_4691 (O_4691,N_44782,N_47625);
or UO_4692 (O_4692,N_47339,N_47348);
or UO_4693 (O_4693,N_46127,N_48620);
and UO_4694 (O_4694,N_43591,N_41590);
and UO_4695 (O_4695,N_47723,N_40375);
and UO_4696 (O_4696,N_45367,N_42883);
xnor UO_4697 (O_4697,N_41475,N_41068);
and UO_4698 (O_4698,N_48568,N_45332);
nor UO_4699 (O_4699,N_44533,N_40948);
nand UO_4700 (O_4700,N_48011,N_45064);
nor UO_4701 (O_4701,N_43414,N_42185);
nor UO_4702 (O_4702,N_49416,N_49407);
nand UO_4703 (O_4703,N_45316,N_49021);
nor UO_4704 (O_4704,N_44664,N_40257);
nor UO_4705 (O_4705,N_47341,N_42781);
xnor UO_4706 (O_4706,N_44201,N_47829);
and UO_4707 (O_4707,N_42138,N_42897);
and UO_4708 (O_4708,N_42389,N_46307);
or UO_4709 (O_4709,N_46388,N_42276);
and UO_4710 (O_4710,N_44435,N_44765);
or UO_4711 (O_4711,N_46190,N_48379);
nor UO_4712 (O_4712,N_44962,N_41365);
nor UO_4713 (O_4713,N_45351,N_49876);
nand UO_4714 (O_4714,N_40263,N_44948);
or UO_4715 (O_4715,N_45744,N_41872);
nand UO_4716 (O_4716,N_49496,N_46461);
nand UO_4717 (O_4717,N_49099,N_42574);
and UO_4718 (O_4718,N_44006,N_44590);
xnor UO_4719 (O_4719,N_40276,N_47778);
nor UO_4720 (O_4720,N_48415,N_45420);
and UO_4721 (O_4721,N_47381,N_43035);
nor UO_4722 (O_4722,N_47411,N_40431);
and UO_4723 (O_4723,N_43248,N_43970);
nor UO_4724 (O_4724,N_47742,N_40048);
nand UO_4725 (O_4725,N_42711,N_42755);
nand UO_4726 (O_4726,N_42681,N_44224);
and UO_4727 (O_4727,N_41665,N_47345);
and UO_4728 (O_4728,N_48015,N_40380);
nor UO_4729 (O_4729,N_47476,N_42160);
nand UO_4730 (O_4730,N_48018,N_49952);
nor UO_4731 (O_4731,N_41290,N_43468);
or UO_4732 (O_4732,N_42258,N_44090);
xor UO_4733 (O_4733,N_49338,N_48716);
and UO_4734 (O_4734,N_45904,N_48330);
or UO_4735 (O_4735,N_46701,N_41977);
nand UO_4736 (O_4736,N_44110,N_47241);
nand UO_4737 (O_4737,N_40096,N_48426);
nand UO_4738 (O_4738,N_41560,N_41589);
or UO_4739 (O_4739,N_46597,N_41624);
and UO_4740 (O_4740,N_43559,N_41972);
nor UO_4741 (O_4741,N_40178,N_46175);
nand UO_4742 (O_4742,N_49195,N_40921);
nor UO_4743 (O_4743,N_49663,N_45300);
and UO_4744 (O_4744,N_46304,N_41692);
xnor UO_4745 (O_4745,N_44309,N_43310);
and UO_4746 (O_4746,N_45241,N_41029);
and UO_4747 (O_4747,N_47591,N_46827);
xor UO_4748 (O_4748,N_42079,N_44921);
or UO_4749 (O_4749,N_46035,N_49080);
and UO_4750 (O_4750,N_41976,N_48321);
xnor UO_4751 (O_4751,N_48786,N_47099);
xor UO_4752 (O_4752,N_47985,N_46923);
nor UO_4753 (O_4753,N_45514,N_41569);
or UO_4754 (O_4754,N_40720,N_47865);
or UO_4755 (O_4755,N_48722,N_45018);
and UO_4756 (O_4756,N_43057,N_48781);
or UO_4757 (O_4757,N_41120,N_47847);
nor UO_4758 (O_4758,N_42776,N_46968);
nand UO_4759 (O_4759,N_45466,N_44351);
and UO_4760 (O_4760,N_46397,N_40932);
xnor UO_4761 (O_4761,N_44527,N_44101);
nor UO_4762 (O_4762,N_40954,N_47454);
or UO_4763 (O_4763,N_46447,N_47918);
or UO_4764 (O_4764,N_41417,N_48235);
nand UO_4765 (O_4765,N_41534,N_40390);
and UO_4766 (O_4766,N_46954,N_41893);
and UO_4767 (O_4767,N_42489,N_44404);
xnor UO_4768 (O_4768,N_48134,N_46410);
xor UO_4769 (O_4769,N_41098,N_45814);
nor UO_4770 (O_4770,N_47892,N_43186);
nand UO_4771 (O_4771,N_43202,N_43066);
or UO_4772 (O_4772,N_49317,N_49385);
and UO_4773 (O_4773,N_49465,N_44475);
and UO_4774 (O_4774,N_45537,N_41779);
nor UO_4775 (O_4775,N_47165,N_48552);
nor UO_4776 (O_4776,N_42934,N_42146);
and UO_4777 (O_4777,N_49350,N_45733);
nor UO_4778 (O_4778,N_40070,N_42084);
and UO_4779 (O_4779,N_41277,N_48046);
or UO_4780 (O_4780,N_45846,N_47219);
nor UO_4781 (O_4781,N_42098,N_42161);
nand UO_4782 (O_4782,N_44777,N_40574);
nand UO_4783 (O_4783,N_49896,N_47049);
and UO_4784 (O_4784,N_41271,N_46723);
xor UO_4785 (O_4785,N_43329,N_49559);
nand UO_4786 (O_4786,N_44645,N_46698);
xnor UO_4787 (O_4787,N_42744,N_42444);
nor UO_4788 (O_4788,N_42108,N_45907);
nand UO_4789 (O_4789,N_45643,N_44432);
and UO_4790 (O_4790,N_48887,N_41482);
and UO_4791 (O_4791,N_49018,N_40935);
or UO_4792 (O_4792,N_47406,N_45848);
xor UO_4793 (O_4793,N_44710,N_47509);
or UO_4794 (O_4794,N_42139,N_42135);
nor UO_4795 (O_4795,N_46240,N_48689);
xnor UO_4796 (O_4796,N_46922,N_40920);
xor UO_4797 (O_4797,N_41909,N_40474);
or UO_4798 (O_4798,N_41787,N_45564);
nor UO_4799 (O_4799,N_45209,N_41241);
and UO_4800 (O_4800,N_41835,N_41889);
nor UO_4801 (O_4801,N_40071,N_44673);
or UO_4802 (O_4802,N_41245,N_43073);
and UO_4803 (O_4803,N_45414,N_41373);
xnor UO_4804 (O_4804,N_42608,N_41194);
nand UO_4805 (O_4805,N_45255,N_44977);
or UO_4806 (O_4806,N_46431,N_41839);
or UO_4807 (O_4807,N_40576,N_42307);
xnor UO_4808 (O_4808,N_40440,N_41246);
nor UO_4809 (O_4809,N_45448,N_45036);
nand UO_4810 (O_4810,N_47525,N_43792);
and UO_4811 (O_4811,N_43562,N_48928);
nor UO_4812 (O_4812,N_48298,N_40373);
or UO_4813 (O_4813,N_42922,N_42985);
nor UO_4814 (O_4814,N_49233,N_43895);
nand UO_4815 (O_4815,N_49113,N_40078);
nor UO_4816 (O_4816,N_42666,N_47141);
and UO_4817 (O_4817,N_41987,N_43905);
or UO_4818 (O_4818,N_43813,N_48423);
or UO_4819 (O_4819,N_44875,N_49096);
nor UO_4820 (O_4820,N_45756,N_48728);
and UO_4821 (O_4821,N_49089,N_42688);
nand UO_4822 (O_4822,N_44176,N_49061);
nand UO_4823 (O_4823,N_49259,N_41573);
nand UO_4824 (O_4824,N_40942,N_45204);
and UO_4825 (O_4825,N_45853,N_40116);
xor UO_4826 (O_4826,N_43247,N_42733);
or UO_4827 (O_4827,N_45286,N_48812);
and UO_4828 (O_4828,N_47313,N_44956);
nand UO_4829 (O_4829,N_41006,N_41028);
or UO_4830 (O_4830,N_43932,N_40086);
and UO_4831 (O_4831,N_42993,N_47041);
or UO_4832 (O_4832,N_40313,N_49825);
nor UO_4833 (O_4833,N_47792,N_49953);
and UO_4834 (O_4834,N_43959,N_43022);
or UO_4835 (O_4835,N_47079,N_48944);
nand UO_4836 (O_4836,N_40215,N_41612);
xor UO_4837 (O_4837,N_45874,N_46989);
and UO_4838 (O_4838,N_47816,N_44598);
nand UO_4839 (O_4839,N_43295,N_41383);
nor UO_4840 (O_4840,N_44636,N_40035);
nor UO_4841 (O_4841,N_45320,N_44978);
nand UO_4842 (O_4842,N_46977,N_49536);
xor UO_4843 (O_4843,N_45323,N_49647);
nor UO_4844 (O_4844,N_48227,N_42101);
and UO_4845 (O_4845,N_47421,N_41111);
xor UO_4846 (O_4846,N_45885,N_46656);
nor UO_4847 (O_4847,N_48345,N_49073);
and UO_4848 (O_4848,N_45390,N_48303);
and UO_4849 (O_4849,N_44167,N_45951);
nor UO_4850 (O_4850,N_48577,N_43188);
nand UO_4851 (O_4851,N_40235,N_46742);
or UO_4852 (O_4852,N_49807,N_47899);
nor UO_4853 (O_4853,N_45929,N_46350);
or UO_4854 (O_4854,N_46675,N_41694);
nand UO_4855 (O_4855,N_45233,N_49542);
nand UO_4856 (O_4856,N_40785,N_49361);
xnor UO_4857 (O_4857,N_43326,N_49327);
or UO_4858 (O_4858,N_40230,N_43362);
nor UO_4859 (O_4859,N_48242,N_47275);
nand UO_4860 (O_4860,N_49320,N_40615);
and UO_4861 (O_4861,N_47202,N_43167);
nor UO_4862 (O_4862,N_42488,N_48454);
nand UO_4863 (O_4863,N_47888,N_47799);
or UO_4864 (O_4864,N_49398,N_46750);
nand UO_4865 (O_4865,N_47869,N_47131);
nor UO_4866 (O_4866,N_43284,N_49224);
nor UO_4867 (O_4867,N_45247,N_41159);
nand UO_4868 (O_4868,N_48890,N_48718);
xnor UO_4869 (O_4869,N_40413,N_42301);
nor UO_4870 (O_4870,N_45386,N_47593);
or UO_4871 (O_4871,N_44445,N_41726);
nor UO_4872 (O_4872,N_43928,N_40058);
and UO_4873 (O_4873,N_47609,N_49278);
nor UO_4874 (O_4874,N_44409,N_42539);
nor UO_4875 (O_4875,N_47067,N_42491);
nand UO_4876 (O_4876,N_48154,N_44515);
nand UO_4877 (O_4877,N_47462,N_47910);
nor UO_4878 (O_4878,N_43307,N_47171);
xor UO_4879 (O_4879,N_45593,N_43243);
and UO_4880 (O_4880,N_49878,N_40798);
and UO_4881 (O_4881,N_40304,N_44361);
nand UO_4882 (O_4882,N_41375,N_40125);
xnor UO_4883 (O_4883,N_41254,N_42519);
nand UO_4884 (O_4884,N_46785,N_41519);
nand UO_4885 (O_4885,N_45487,N_47104);
nor UO_4886 (O_4886,N_43869,N_45426);
nand UO_4887 (O_4887,N_47281,N_48399);
or UO_4888 (O_4888,N_48982,N_40558);
nor UO_4889 (O_4889,N_41791,N_45843);
and UO_4890 (O_4890,N_40583,N_46006);
and UO_4891 (O_4891,N_41215,N_43778);
or UO_4892 (O_4892,N_46153,N_42774);
or UO_4893 (O_4893,N_43170,N_42020);
nor UO_4894 (O_4894,N_40324,N_45722);
nand UO_4895 (O_4895,N_44558,N_40179);
or UO_4896 (O_4896,N_41070,N_43413);
nand UO_4897 (O_4897,N_46168,N_42275);
nor UO_4898 (O_4898,N_41727,N_40468);
or UO_4899 (O_4899,N_47988,N_48306);
or UO_4900 (O_4900,N_41859,N_45574);
xnor UO_4901 (O_4901,N_45891,N_48459);
and UO_4902 (O_4902,N_48036,N_44805);
nor UO_4903 (O_4903,N_42878,N_49452);
nor UO_4904 (O_4904,N_41289,N_45935);
xnor UO_4905 (O_4905,N_44350,N_43716);
or UO_4906 (O_4906,N_44588,N_47641);
or UO_4907 (O_4907,N_49119,N_49712);
nor UO_4908 (O_4908,N_46155,N_40199);
nor UO_4909 (O_4909,N_49122,N_41652);
nor UO_4910 (O_4910,N_42992,N_42297);
xor UO_4911 (O_4911,N_49144,N_46250);
nand UO_4912 (O_4912,N_48701,N_47393);
nand UO_4913 (O_4913,N_49030,N_42235);
nor UO_4914 (O_4914,N_43194,N_45966);
nand UO_4915 (O_4915,N_49057,N_42211);
and UO_4916 (O_4916,N_42788,N_43040);
or UO_4917 (O_4917,N_48039,N_43976);
and UO_4918 (O_4918,N_42734,N_47795);
or UO_4919 (O_4919,N_44812,N_41549);
nor UO_4920 (O_4920,N_47575,N_41366);
and UO_4921 (O_4921,N_49858,N_40675);
or UO_4922 (O_4922,N_40439,N_44648);
xnor UO_4923 (O_4923,N_43003,N_42001);
and UO_4924 (O_4924,N_48592,N_45902);
nor UO_4925 (O_4925,N_45175,N_48405);
nand UO_4926 (O_4926,N_42798,N_40320);
and UO_4927 (O_4927,N_41301,N_42919);
xnor UO_4928 (O_4928,N_40128,N_42643);
nand UO_4929 (O_4929,N_42671,N_44026);
nand UO_4930 (O_4930,N_42886,N_48653);
or UO_4931 (O_4931,N_41381,N_43807);
or UO_4932 (O_4932,N_41490,N_49609);
nor UO_4933 (O_4933,N_43868,N_42148);
xnor UO_4934 (O_4934,N_48136,N_42847);
nor UO_4935 (O_4935,N_44040,N_41989);
nor UO_4936 (O_4936,N_44892,N_43745);
or UO_4937 (O_4937,N_43523,N_48886);
or UO_4938 (O_4938,N_46746,N_48869);
xor UO_4939 (O_4939,N_49882,N_46403);
xor UO_4940 (O_4940,N_46170,N_43090);
nor UO_4941 (O_4941,N_48259,N_42314);
or UO_4942 (O_4942,N_40753,N_44476);
nand UO_4943 (O_4943,N_43212,N_44355);
or UO_4944 (O_4944,N_46438,N_45801);
or UO_4945 (O_4945,N_44153,N_44616);
xor UO_4946 (O_4946,N_40394,N_48970);
nand UO_4947 (O_4947,N_47913,N_43271);
or UO_4948 (O_4948,N_40381,N_47612);
or UO_4949 (O_4949,N_42829,N_46053);
nor UO_4950 (O_4950,N_45465,N_44559);
xor UO_4951 (O_4951,N_41873,N_48614);
xnor UO_4952 (O_4952,N_46655,N_49802);
nor UO_4953 (O_4953,N_40010,N_45713);
or UO_4954 (O_4954,N_47091,N_45093);
nand UO_4955 (O_4955,N_43440,N_49946);
or UO_4956 (O_4956,N_43899,N_42590);
nor UO_4957 (O_4957,N_40622,N_45428);
nor UO_4958 (O_4958,N_43389,N_41916);
or UO_4959 (O_4959,N_41103,N_48609);
nor UO_4960 (O_4960,N_47740,N_41438);
nor UO_4961 (O_4961,N_48768,N_44396);
nand UO_4962 (O_4962,N_44840,N_46564);
nor UO_4963 (O_4963,N_40995,N_48511);
or UO_4964 (O_4964,N_45089,N_44986);
and UO_4965 (O_4965,N_42062,N_40229);
nand UO_4966 (O_4966,N_45179,N_47986);
or UO_4967 (O_4967,N_47111,N_40950);
and UO_4968 (O_4968,N_46570,N_48277);
or UO_4969 (O_4969,N_43596,N_42720);
or UO_4970 (O_4970,N_46163,N_48326);
or UO_4971 (O_4971,N_49842,N_40209);
nand UO_4972 (O_4972,N_40873,N_40959);
xnor UO_4973 (O_4973,N_41221,N_45094);
xor UO_4974 (O_4974,N_47517,N_45235);
or UO_4975 (O_4975,N_42602,N_44257);
and UO_4976 (O_4976,N_42768,N_41662);
or UO_4977 (O_4977,N_49316,N_48507);
nor UO_4978 (O_4978,N_40834,N_47443);
xnor UO_4979 (O_4979,N_45971,N_40881);
or UO_4980 (O_4980,N_48093,N_44232);
nor UO_4981 (O_4981,N_47813,N_41218);
and UO_4982 (O_4982,N_45067,N_42909);
and UO_4983 (O_4983,N_47205,N_48933);
or UO_4984 (O_4984,N_49159,N_43798);
and UO_4985 (O_4985,N_41586,N_43927);
nor UO_4986 (O_4986,N_40515,N_41702);
nor UO_4987 (O_4987,N_42633,N_41606);
nand UO_4988 (O_4988,N_40410,N_49755);
and UO_4989 (O_4989,N_42401,N_45631);
and UO_4990 (O_4990,N_49661,N_44600);
nor UO_4991 (O_4991,N_48331,N_45488);
xor UO_4992 (O_4992,N_41378,N_45341);
nor UO_4993 (O_4993,N_40898,N_46917);
nand UO_4994 (O_4994,N_42153,N_42676);
nor UO_4995 (O_4995,N_45372,N_41809);
xor UO_4996 (O_4996,N_40776,N_40389);
nor UO_4997 (O_4997,N_47180,N_42077);
nor UO_4998 (O_4998,N_41819,N_41312);
or UO_4999 (O_4999,N_41833,N_47499);
endmodule