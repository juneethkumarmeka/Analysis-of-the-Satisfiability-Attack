module basic_1000_10000_1500_100_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_322,In_774);
or U1 (N_1,In_6,In_476);
nand U2 (N_2,In_118,In_240);
nor U3 (N_3,In_320,In_160);
xnor U4 (N_4,In_108,In_573);
nor U5 (N_5,In_687,In_655);
nand U6 (N_6,In_727,In_686);
and U7 (N_7,In_807,In_470);
xnor U8 (N_8,In_722,In_915);
xor U9 (N_9,In_795,In_839);
nor U10 (N_10,In_175,In_404);
nor U11 (N_11,In_95,In_783);
nor U12 (N_12,In_270,In_397);
and U13 (N_13,In_215,In_822);
nand U14 (N_14,In_842,In_164);
nor U15 (N_15,In_789,In_65);
or U16 (N_16,In_754,In_708);
nor U17 (N_17,In_134,In_582);
nand U18 (N_18,In_468,In_712);
xor U19 (N_19,In_970,In_55);
xor U20 (N_20,In_45,In_878);
nand U21 (N_21,In_58,In_291);
nor U22 (N_22,In_467,In_54);
or U23 (N_23,In_459,In_905);
nor U24 (N_24,In_618,In_988);
nand U25 (N_25,In_979,In_13);
and U26 (N_26,In_519,In_504);
nand U27 (N_27,In_244,In_833);
or U28 (N_28,In_870,In_953);
xnor U29 (N_29,In_121,In_876);
nor U30 (N_30,In_625,In_183);
xnor U31 (N_31,In_858,In_873);
nand U32 (N_32,In_697,In_318);
and U33 (N_33,In_414,In_493);
nand U34 (N_34,In_197,In_227);
or U35 (N_35,In_177,In_163);
and U36 (N_36,In_917,In_141);
nor U37 (N_37,In_604,In_838);
or U38 (N_38,In_828,In_739);
nand U39 (N_39,In_680,In_926);
nand U40 (N_40,In_555,In_460);
xnor U41 (N_41,In_332,In_17);
xnor U42 (N_42,In_14,In_957);
nand U43 (N_43,In_304,In_85);
and U44 (N_44,In_700,In_855);
and U45 (N_45,In_885,In_103);
nor U46 (N_46,In_997,In_2);
or U47 (N_47,In_880,In_360);
and U48 (N_48,In_330,In_362);
nor U49 (N_49,In_144,In_613);
nand U50 (N_50,In_978,In_530);
or U51 (N_51,In_740,In_678);
or U52 (N_52,In_66,In_268);
nor U53 (N_53,In_943,In_233);
nor U54 (N_54,In_338,In_348);
or U55 (N_55,In_76,In_196);
nor U56 (N_56,In_889,In_854);
nand U57 (N_57,In_384,In_882);
and U58 (N_58,In_863,In_714);
nor U59 (N_59,In_331,In_689);
nor U60 (N_60,In_374,In_225);
and U61 (N_61,In_888,In_831);
nor U62 (N_62,In_284,In_777);
or U63 (N_63,In_881,In_758);
nor U64 (N_64,In_531,In_26);
nor U65 (N_65,In_505,In_761);
nor U66 (N_66,In_825,In_168);
xor U67 (N_67,In_736,In_968);
nor U68 (N_68,In_329,In_550);
nand U69 (N_69,In_715,In_278);
nand U70 (N_70,In_817,In_796);
xnor U71 (N_71,In_602,In_998);
nor U72 (N_72,In_595,In_744);
nand U73 (N_73,In_829,In_934);
or U74 (N_74,In_326,In_986);
xnor U75 (N_75,In_238,In_96);
or U76 (N_76,In_371,In_907);
nor U77 (N_77,In_305,In_461);
and U78 (N_78,In_213,In_526);
nand U79 (N_79,In_773,In_436);
nor U80 (N_80,In_797,In_287);
nor U81 (N_81,In_21,In_308);
xnor U82 (N_82,In_241,In_67);
xor U83 (N_83,In_560,In_984);
and U84 (N_84,In_140,In_746);
nand U85 (N_85,In_69,In_852);
xor U86 (N_86,In_937,In_22);
and U87 (N_87,In_859,In_650);
and U88 (N_88,In_977,In_884);
nand U89 (N_89,In_200,In_11);
and U90 (N_90,In_895,In_10);
xor U91 (N_91,In_516,In_999);
nand U92 (N_92,In_276,In_192);
nor U93 (N_93,In_420,In_311);
and U94 (N_94,In_925,In_169);
xnor U95 (N_95,In_117,In_345);
nor U96 (N_96,In_283,In_851);
nor U97 (N_97,In_299,In_34);
or U98 (N_98,In_646,In_90);
xor U99 (N_99,In_656,In_622);
or U100 (N_100,In_63,In_313);
and U101 (N_101,In_8,In_229);
and U102 (N_102,In_166,N_33);
or U103 (N_103,In_205,In_563);
nor U104 (N_104,In_955,In_844);
nor U105 (N_105,N_79,In_540);
xnor U106 (N_106,In_632,In_690);
or U107 (N_107,In_378,In_503);
xor U108 (N_108,In_60,In_629);
nand U109 (N_109,In_472,In_853);
and U110 (N_110,In_517,In_931);
or U111 (N_111,In_285,In_152);
nor U112 (N_112,In_264,In_286);
nand U113 (N_113,N_78,In_927);
xor U114 (N_114,In_119,In_124);
or U115 (N_115,In_256,In_586);
nor U116 (N_116,In_228,In_257);
nand U117 (N_117,In_150,In_684);
nand U118 (N_118,In_790,In_428);
or U119 (N_119,In_91,In_969);
and U120 (N_120,In_403,In_94);
nand U121 (N_121,In_588,In_932);
nand U122 (N_122,N_26,In_778);
nand U123 (N_123,In_843,In_261);
nand U124 (N_124,In_958,In_510);
xnor U125 (N_125,In_438,In_897);
nor U126 (N_126,In_155,In_711);
and U127 (N_127,In_68,N_84);
xnor U128 (N_128,In_695,In_691);
nor U129 (N_129,N_55,In_989);
and U130 (N_130,In_146,In_20);
and U131 (N_131,In_661,In_966);
nand U132 (N_132,In_137,In_250);
nor U133 (N_133,In_395,In_993);
xnor U134 (N_134,N_87,In_487);
nand U135 (N_135,In_860,In_814);
nor U136 (N_136,In_741,N_41);
or U137 (N_137,In_914,In_439);
xor U138 (N_138,In_841,N_4);
or U139 (N_139,In_775,In_954);
xnor U140 (N_140,N_46,In_201);
and U141 (N_141,In_791,N_37);
or U142 (N_142,In_982,In_353);
nand U143 (N_143,In_537,In_832);
or U144 (N_144,In_56,In_755);
and U145 (N_145,In_748,N_97);
xnor U146 (N_146,In_801,In_370);
nand U147 (N_147,N_88,In_921);
xor U148 (N_148,In_587,In_845);
nor U149 (N_149,In_580,In_826);
nand U150 (N_150,In_142,In_612);
or U151 (N_151,In_725,In_543);
and U152 (N_152,N_22,In_802);
and U153 (N_153,In_593,N_60);
or U154 (N_154,In_62,In_617);
or U155 (N_155,In_309,In_433);
nor U156 (N_156,N_43,In_341);
nor U157 (N_157,In_713,In_992);
xnor U158 (N_158,In_938,In_449);
xnor U159 (N_159,In_407,In_116);
xor U160 (N_160,In_928,N_51);
xnor U161 (N_161,In_477,In_294);
nand U162 (N_162,In_385,In_749);
or U163 (N_163,In_834,In_527);
xnor U164 (N_164,In_717,In_640);
xor U165 (N_165,In_110,In_15);
nand U166 (N_166,In_962,In_770);
xnor U167 (N_167,In_728,In_699);
nand U168 (N_168,In_805,In_564);
and U169 (N_169,In_375,In_79);
nand U170 (N_170,N_7,In_806);
or U171 (N_171,In_597,In_138);
xor U172 (N_172,In_753,In_990);
nand U173 (N_173,N_99,In_923);
nand U174 (N_174,In_86,In_672);
and U175 (N_175,In_631,In_206);
xor U176 (N_176,N_66,In_98);
nor U177 (N_177,In_50,In_426);
or U178 (N_178,In_185,In_589);
nand U179 (N_179,In_887,In_871);
nand U180 (N_180,In_608,In_983);
or U181 (N_181,N_42,In_295);
and U182 (N_182,N_36,In_821);
xnor U183 (N_183,N_64,N_25);
and U184 (N_184,In_251,In_135);
and U185 (N_185,In_649,In_651);
nand U186 (N_186,In_275,In_377);
or U187 (N_187,In_751,In_660);
xor U188 (N_188,In_425,In_720);
and U189 (N_189,In_489,In_349);
or U190 (N_190,In_33,In_123);
or U191 (N_191,In_682,In_383);
and U192 (N_192,N_95,In_598);
and U193 (N_193,N_35,In_346);
nand U194 (N_194,In_867,In_130);
xnor U195 (N_195,In_752,In_974);
or U196 (N_196,In_894,In_764);
xnor U197 (N_197,In_165,N_59);
nand U198 (N_198,In_53,In_184);
nor U199 (N_199,N_1,In_359);
nand U200 (N_200,In_626,N_183);
nor U201 (N_201,In_223,In_226);
or U202 (N_202,In_47,N_62);
or U203 (N_203,In_388,In_418);
or U204 (N_204,N_14,In_702);
nand U205 (N_205,In_594,In_730);
or U206 (N_206,In_492,In_576);
and U207 (N_207,In_396,In_837);
and U208 (N_208,In_872,N_50);
or U209 (N_209,In_178,In_929);
or U210 (N_210,In_214,In_657);
or U211 (N_211,In_87,In_424);
and U212 (N_212,In_263,In_431);
xnor U213 (N_213,In_488,In_48);
or U214 (N_214,In_239,In_210);
and U215 (N_215,In_849,In_81);
or U216 (N_216,In_149,In_344);
nor U217 (N_217,In_366,In_782);
and U218 (N_218,In_333,In_18);
xor U219 (N_219,In_195,In_145);
and U220 (N_220,In_981,In_113);
or U221 (N_221,In_742,In_203);
or U222 (N_222,N_144,In_658);
nand U223 (N_223,In_231,In_965);
xnor U224 (N_224,In_731,N_111);
and U225 (N_225,In_158,In_495);
and U226 (N_226,N_34,In_198);
and U227 (N_227,In_951,In_514);
and U228 (N_228,In_552,N_149);
and U229 (N_229,N_175,In_167);
and U230 (N_230,In_599,N_75);
and U231 (N_231,In_281,In_181);
xnor U232 (N_232,N_184,In_562);
and U233 (N_233,In_78,In_128);
xor U234 (N_234,In_912,In_342);
nor U235 (N_235,In_232,In_217);
nand U236 (N_236,In_180,In_901);
and U237 (N_237,In_389,In_315);
nand U238 (N_238,In_452,In_445);
and U239 (N_239,In_558,N_118);
xor U240 (N_240,N_147,In_478);
or U241 (N_241,In_367,In_967);
and U242 (N_242,In_42,In_792);
or U243 (N_243,In_557,In_77);
and U244 (N_244,N_5,In_918);
or U245 (N_245,In_52,In_772);
nand U246 (N_246,In_539,In_653);
nor U247 (N_247,In_709,In_911);
nor U248 (N_248,In_960,In_413);
nor U249 (N_249,In_179,In_868);
or U250 (N_250,N_109,N_49);
xor U251 (N_251,In_502,In_642);
nor U252 (N_252,In_457,N_136);
xnor U253 (N_253,In_575,In_245);
xor U254 (N_254,In_447,In_781);
nor U255 (N_255,In_939,In_671);
and U256 (N_256,In_24,In_288);
nor U257 (N_257,N_13,In_886);
and U258 (N_258,N_23,N_176);
nand U259 (N_259,In_544,In_28);
and U260 (N_260,In_991,N_96);
nand U261 (N_261,In_952,N_137);
nor U262 (N_262,In_71,In_415);
and U263 (N_263,In_756,N_77);
and U264 (N_264,In_836,In_298);
nand U265 (N_265,In_664,In_601);
and U266 (N_266,In_767,In_600);
nor U267 (N_267,In_779,In_387);
nand U268 (N_268,In_857,In_328);
nor U269 (N_269,In_636,In_910);
xnor U270 (N_270,In_846,N_199);
nand U271 (N_271,In_316,N_141);
xor U272 (N_272,In_273,In_237);
or U273 (N_273,In_975,In_784);
nor U274 (N_274,In_199,In_898);
or U275 (N_275,N_94,In_75);
xnor U276 (N_276,N_105,N_101);
nand U277 (N_277,N_139,N_82);
nor U278 (N_278,In_464,In_920);
nor U279 (N_279,In_703,In_569);
or U280 (N_280,In_89,In_735);
xor U281 (N_281,In_485,In_64);
or U282 (N_282,In_698,In_515);
or U283 (N_283,N_172,In_693);
nor U284 (N_284,In_446,In_43);
or U285 (N_285,N_57,N_153);
nor U286 (N_286,In_31,In_339);
xnor U287 (N_287,In_314,In_49);
nand U288 (N_288,N_127,In_104);
or U289 (N_289,In_30,In_665);
xnor U290 (N_290,In_350,N_9);
xor U291 (N_291,In_463,In_83);
nor U292 (N_292,In_72,In_676);
and U293 (N_293,In_193,In_696);
nand U294 (N_294,In_547,N_72);
xor U295 (N_295,In_721,In_762);
xor U296 (N_296,In_584,In_368);
or U297 (N_297,In_260,In_961);
nand U298 (N_298,In_102,In_610);
or U299 (N_299,In_292,In_766);
or U300 (N_300,N_91,N_201);
nand U301 (N_301,In_706,In_498);
or U302 (N_302,In_624,In_716);
and U303 (N_303,In_379,N_15);
nor U304 (N_304,N_245,In_474);
xor U305 (N_305,In_209,In_819);
xor U306 (N_306,In_804,In_127);
nand U307 (N_307,In_143,In_139);
nor U308 (N_308,In_615,In_258);
xor U309 (N_309,In_606,In_820);
nor U310 (N_310,In_41,N_165);
nor U311 (N_311,In_16,In_361);
xnor U312 (N_312,N_298,N_234);
nand U313 (N_313,In_737,In_327);
nand U314 (N_314,In_173,In_572);
nor U315 (N_315,N_185,In_112);
and U316 (N_316,In_444,N_257);
nand U317 (N_317,In_211,In_216);
xor U318 (N_318,In_723,N_117);
xor U319 (N_319,In_466,N_295);
and U320 (N_320,In_620,N_269);
and U321 (N_321,In_635,In_114);
and U322 (N_322,In_99,In_808);
nor U323 (N_323,N_264,N_291);
or U324 (N_324,In_648,In_567);
xor U325 (N_325,In_818,In_490);
and U326 (N_326,In_9,In_701);
or U327 (N_327,In_964,In_132);
nand U328 (N_328,In_933,In_596);
or U329 (N_329,In_913,In_187);
or U330 (N_330,N_40,In_750);
xor U331 (N_331,N_28,In_638);
or U332 (N_332,In_824,N_250);
nand U333 (N_333,N_220,N_256);
and U334 (N_334,In_520,In_80);
nor U335 (N_335,N_261,In_306);
xnor U336 (N_336,In_394,In_101);
and U337 (N_337,In_335,In_337);
or U338 (N_338,In_948,In_985);
or U339 (N_339,In_451,In_351);
nor U340 (N_340,In_486,In_61);
nand U341 (N_341,N_100,N_266);
and U342 (N_342,In_724,In_518);
xor U343 (N_343,N_152,In_816);
nand U344 (N_344,In_521,N_159);
and U345 (N_345,In_535,In_681);
nor U346 (N_346,N_207,In_280);
or U347 (N_347,N_275,In_692);
nor U348 (N_348,In_266,In_236);
and U349 (N_349,In_565,In_522);
nor U350 (N_350,In_891,In_669);
and U351 (N_351,N_83,In_136);
nor U352 (N_352,In_553,In_729);
xor U353 (N_353,In_448,In_373);
xnor U354 (N_354,In_207,N_86);
nand U355 (N_355,In_949,In_399);
or U356 (N_356,N_272,In_409);
and U357 (N_357,In_482,In_592);
nor U358 (N_358,N_277,In_186);
nand U359 (N_359,N_52,N_65);
nand U360 (N_360,N_283,In_663);
nand U361 (N_361,N_222,In_369);
nand U362 (N_362,In_212,In_302);
nand U363 (N_363,In_365,In_507);
nor U364 (N_364,N_209,In_410);
nand U365 (N_365,N_54,In_19);
and U366 (N_366,N_69,N_268);
or U367 (N_367,In_92,N_204);
xnor U368 (N_368,In_434,In_44);
or U369 (N_369,In_246,In_471);
and U370 (N_370,N_293,In_903);
nor U371 (N_371,In_904,In_972);
and U372 (N_372,In_963,In_574);
nor U373 (N_373,N_126,In_614);
or U374 (N_374,N_262,N_196);
or U375 (N_375,N_19,N_189);
nand U376 (N_376,In_645,In_996);
and U377 (N_377,In_738,In_611);
nand U378 (N_378,In_390,In_190);
nor U379 (N_379,In_590,In_148);
nor U380 (N_380,In_255,N_58);
or U381 (N_381,In_946,N_120);
nand U382 (N_382,In_554,In_230);
nand U383 (N_383,In_391,In_443);
or U384 (N_384,N_239,In_812);
and U385 (N_385,In_39,In_513);
and U386 (N_386,In_456,In_234);
xor U387 (N_387,In_412,In_297);
nor U388 (N_388,N_21,In_267);
xnor U389 (N_389,N_211,N_107);
and U390 (N_390,N_228,In_710);
nand U391 (N_391,In_956,N_81);
nand U392 (N_392,In_29,In_799);
xnor U393 (N_393,N_255,In_381);
and U394 (N_394,N_267,N_71);
nand U395 (N_395,N_177,N_198);
nand U396 (N_396,N_212,N_223);
nand U397 (N_397,In_46,N_238);
and U398 (N_398,N_27,N_156);
nor U399 (N_399,N_202,N_39);
and U400 (N_400,N_383,N_205);
nor U401 (N_401,In_393,N_348);
nor U402 (N_402,In_890,N_6);
nand U403 (N_403,N_17,In_57);
and U404 (N_404,In_679,N_350);
or U405 (N_405,In_122,In_675);
xnor U406 (N_406,N_128,N_397);
or U407 (N_407,In_0,N_384);
nor U408 (N_408,N_8,N_394);
and U409 (N_409,In_902,N_258);
xnor U410 (N_410,N_192,N_296);
or U411 (N_411,In_242,In_97);
nand U412 (N_412,N_368,In_785);
xor U413 (N_413,In_204,N_382);
and U414 (N_414,In_462,N_381);
nor U415 (N_415,In_509,In_976);
or U416 (N_416,N_0,In_162);
and U417 (N_417,N_286,N_138);
xor U418 (N_418,In_759,N_186);
nor U419 (N_419,In_105,In_621);
and U420 (N_420,N_190,N_251);
nor U421 (N_421,N_326,In_93);
and U422 (N_422,N_370,In_936);
nor U423 (N_423,N_122,N_68);
xnor U424 (N_424,In_800,N_252);
xor U425 (N_425,N_325,In_659);
nor U426 (N_426,In_561,In_523);
xor U427 (N_427,In_652,N_310);
nor U428 (N_428,In_500,N_151);
and U429 (N_429,N_89,N_313);
nand U430 (N_430,N_339,N_30);
nand U431 (N_431,N_18,In_628);
nor U432 (N_432,In_533,N_284);
and U433 (N_433,In_469,In_793);
xor U434 (N_434,In_666,In_899);
nand U435 (N_435,In_623,N_387);
nand U436 (N_436,In_188,N_161);
or U437 (N_437,N_24,N_125);
nand U438 (N_438,N_215,In_823);
nand U439 (N_439,In_455,In_51);
nand U440 (N_440,N_154,In_347);
xnor U441 (N_441,N_174,N_113);
nor U442 (N_442,N_47,In_771);
xnor U443 (N_443,In_667,In_70);
xnor U444 (N_444,In_512,N_289);
nand U445 (N_445,In_830,In_82);
nand U446 (N_446,In_534,N_337);
xnor U447 (N_447,In_511,In_269);
xnor U448 (N_448,In_637,N_319);
and U449 (N_449,N_287,In_340);
xor U450 (N_450,N_398,N_320);
or U451 (N_451,N_306,N_301);
or U452 (N_452,N_106,N_32);
or U453 (N_453,In_354,In_271);
nor U454 (N_454,In_115,In_3);
xor U455 (N_455,In_566,In_685);
and U456 (N_456,N_243,N_352);
nor U457 (N_457,N_121,In_673);
or U458 (N_458,N_386,In_668);
xor U459 (N_459,In_191,In_363);
nor U460 (N_460,N_90,In_479);
xor U461 (N_461,In_532,In_111);
xnor U462 (N_462,N_242,In_290);
or U463 (N_463,In_607,N_203);
and U464 (N_464,N_200,In_609);
or U465 (N_465,In_25,In_528);
or U466 (N_466,In_277,N_335);
nand U467 (N_467,In_619,In_4);
or U468 (N_468,In_995,In_483);
nand U469 (N_469,N_341,N_232);
nand U470 (N_470,N_237,In_12);
and U471 (N_471,In_151,N_233);
nand U472 (N_472,N_210,In_296);
nand U473 (N_473,In_864,In_475);
nand U474 (N_474,In_760,N_70);
nor U475 (N_475,In_549,N_143);
nand U476 (N_476,N_173,In_506);
xnor U477 (N_477,In_571,In_411);
and U478 (N_478,N_132,In_325);
and U479 (N_479,N_351,N_235);
nor U480 (N_480,N_259,In_559);
or U481 (N_481,In_120,N_380);
or U482 (N_482,In_940,N_317);
xnor U483 (N_483,N_67,N_260);
and U484 (N_484,In_252,In_548);
nand U485 (N_485,In_253,N_116);
nand U486 (N_486,In_417,N_347);
nand U487 (N_487,N_373,In_38);
nand U488 (N_488,In_153,In_627);
or U489 (N_489,N_349,In_683);
nor U490 (N_490,N_169,N_327);
nand U491 (N_491,N_76,In_247);
or U492 (N_492,In_408,In_40);
nor U493 (N_493,In_88,In_950);
nor U494 (N_494,In_129,In_154);
and U495 (N_495,In_786,In_869);
nor U496 (N_496,In_194,N_390);
nand U497 (N_497,In_647,In_356);
nand U498 (N_498,N_240,In_133);
xnor U499 (N_499,N_364,N_247);
xnor U500 (N_500,In_484,N_363);
nand U501 (N_501,N_323,In_174);
xor U502 (N_502,N_112,N_400);
xor U503 (N_503,In_402,N_396);
or U504 (N_504,In_432,In_747);
xnor U505 (N_505,N_216,N_473);
xnor U506 (N_506,In_900,N_303);
nand U507 (N_507,In_357,N_288);
nor U508 (N_508,N_463,In_745);
xnor U509 (N_509,In_603,N_29);
nor U510 (N_510,In_37,In_674);
nor U511 (N_511,N_421,N_425);
nor U512 (N_512,N_464,N_497);
nor U513 (N_513,N_276,N_342);
nand U514 (N_514,N_433,In_922);
nand U515 (N_515,N_322,N_359);
nand U516 (N_516,N_218,N_290);
or U517 (N_517,N_443,In_427);
or U518 (N_518,In_570,In_172);
xor U519 (N_519,In_147,N_224);
nand U520 (N_520,N_470,In_546);
or U521 (N_521,N_230,N_119);
nor U522 (N_522,In_176,In_688);
and U523 (N_523,In_491,N_448);
nand U524 (N_524,N_451,In_879);
nand U525 (N_525,In_497,N_38);
or U526 (N_526,In_973,In_866);
and U527 (N_527,N_436,In_809);
nand U528 (N_528,N_478,In_862);
nand U529 (N_529,N_439,N_131);
and U530 (N_530,N_449,In_5);
xnor U531 (N_531,N_401,N_248);
nor U532 (N_532,N_333,N_155);
or U533 (N_533,N_182,N_494);
xnor U534 (N_534,In_896,N_31);
nand U535 (N_535,In_811,N_389);
nor U536 (N_536,In_780,N_442);
nand U537 (N_537,N_450,In_930);
nand U538 (N_538,In_170,N_358);
and U539 (N_539,In_450,N_366);
nor U540 (N_540,In_941,In_35);
xor U541 (N_541,N_444,In_581);
nor U542 (N_542,In_317,In_307);
nand U543 (N_543,N_56,N_10);
xnor U544 (N_544,In_171,N_74);
or U545 (N_545,N_180,In_303);
xor U546 (N_546,In_556,N_445);
and U547 (N_547,In_401,N_371);
nand U548 (N_548,In_481,N_282);
or U549 (N_549,In_794,In_243);
and U550 (N_550,In_892,In_787);
or U551 (N_551,N_110,In_616);
xnor U552 (N_552,In_437,N_465);
and U553 (N_553,N_221,N_455);
nand U554 (N_554,In_421,In_499);
nor U555 (N_555,In_776,N_20);
nor U556 (N_556,N_130,N_431);
or U557 (N_557,N_135,In_757);
nand U558 (N_558,N_369,N_332);
nor U559 (N_559,In_248,N_385);
nor U560 (N_560,N_360,In_249);
and U561 (N_561,N_480,In_835);
nor U562 (N_562,In_908,In_704);
or U563 (N_563,N_393,N_399);
nor U564 (N_564,N_2,In_768);
and U565 (N_565,In_161,In_100);
nand U566 (N_566,N_231,In_525);
nor U567 (N_567,N_12,N_429);
nand U568 (N_568,N_302,N_170);
and U569 (N_569,In_644,In_376);
or U570 (N_570,N_417,In_1);
nand U571 (N_571,N_278,In_909);
nor U572 (N_572,In_202,N_178);
nand U573 (N_573,N_422,N_468);
or U574 (N_574,In_458,N_430);
or U575 (N_575,N_437,In_480);
nor U576 (N_576,In_765,N_206);
xor U577 (N_577,N_488,N_194);
xor U578 (N_578,N_392,N_213);
nor U579 (N_579,In_850,N_53);
nor U580 (N_580,N_432,In_454);
and U581 (N_581,In_310,N_416);
and U582 (N_582,N_92,N_133);
or U583 (N_583,N_376,N_408);
xnor U584 (N_584,N_419,N_274);
nand U585 (N_585,In_189,In_254);
and U586 (N_586,N_489,N_324);
or U587 (N_587,N_476,N_158);
xnor U588 (N_588,N_440,N_285);
xnor U589 (N_589,N_481,N_361);
nand U590 (N_590,In_980,In_803);
or U591 (N_591,In_74,In_224);
and U592 (N_592,N_273,N_423);
or U593 (N_593,N_271,N_98);
xor U594 (N_594,N_11,In_406);
xor U595 (N_595,In_423,N_294);
nand U596 (N_596,In_352,In_182);
xnor U597 (N_597,N_453,In_639);
nor U598 (N_598,N_168,In_358);
nand U599 (N_599,In_501,N_309);
nand U600 (N_600,N_148,In_334);
xnor U601 (N_601,N_586,N_559);
nor U602 (N_602,N_409,N_410);
nand U603 (N_603,N_197,In_763);
and U604 (N_604,N_555,In_419);
nand U605 (N_605,N_441,N_395);
and U606 (N_606,N_564,N_541);
and U607 (N_607,N_483,In_159);
or U608 (N_608,In_947,In_707);
nor U609 (N_609,N_505,In_125);
nor U610 (N_610,N_501,N_466);
or U611 (N_611,N_93,In_405);
nor U612 (N_612,In_591,N_265);
xnor U613 (N_613,In_585,N_539);
nand U614 (N_614,N_535,In_827);
xor U615 (N_615,N_299,N_354);
xor U616 (N_616,N_556,In_959);
and U617 (N_617,In_293,In_274);
or U618 (N_618,N_458,N_527);
and U619 (N_619,N_241,N_581);
or U620 (N_620,N_146,In_994);
xor U621 (N_621,N_129,In_272);
nor U622 (N_622,N_150,In_578);
or U623 (N_623,N_580,N_588);
xnor U624 (N_624,N_362,N_508);
nor U625 (N_625,In_430,In_529);
nor U626 (N_626,In_453,In_355);
xnor U627 (N_627,N_160,In_630);
xor U628 (N_628,N_583,N_379);
nor U629 (N_629,N_479,N_281);
and U630 (N_630,N_340,N_405);
nor U631 (N_631,In_221,N_491);
nor U632 (N_632,N_114,In_126);
and U633 (N_633,N_518,N_344);
xnor U634 (N_634,N_574,N_193);
and U635 (N_635,In_73,N_187);
and U636 (N_636,In_84,N_402);
or U637 (N_637,In_874,N_515);
and U638 (N_638,In_7,N_315);
or U639 (N_639,In_893,N_590);
nor U640 (N_640,N_546,N_312);
xor U641 (N_641,N_456,N_343);
nand U642 (N_642,N_307,In_718);
nand U643 (N_643,N_3,N_500);
and U644 (N_644,N_597,In_798);
or U645 (N_645,In_694,In_633);
and U646 (N_646,In_924,In_473);
nor U647 (N_647,N_460,In_971);
nand U648 (N_648,N_577,N_571);
or U649 (N_649,In_551,N_63);
and U650 (N_650,In_440,N_578);
and U651 (N_651,In_380,N_486);
xor U652 (N_652,N_587,In_605);
xnor U653 (N_653,In_508,In_877);
and U654 (N_654,N_374,N_594);
nand U655 (N_655,N_164,N_208);
xor U656 (N_656,N_534,N_426);
nand U657 (N_657,In_321,N_569);
and U658 (N_658,N_502,In_465);
nand U659 (N_659,N_328,N_575);
nor U660 (N_660,N_311,In_156);
or U661 (N_661,N_179,N_411);
and U662 (N_662,N_512,N_438);
and U663 (N_663,N_498,N_124);
nand U664 (N_664,N_572,N_585);
nor U665 (N_665,N_514,In_856);
nand U666 (N_666,N_292,N_506);
and U667 (N_667,N_558,N_145);
nor U668 (N_668,In_262,In_131);
nor U669 (N_669,In_875,In_577);
xnor U670 (N_670,N_263,In_289);
or U671 (N_671,N_530,In_945);
and U672 (N_672,In_545,N_472);
nor U673 (N_673,In_634,N_434);
and U674 (N_674,N_528,In_300);
or U675 (N_675,N_44,In_705);
xor U676 (N_676,In_323,N_428);
nor U677 (N_677,In_847,N_533);
nand U678 (N_678,In_106,N_531);
xor U679 (N_679,In_541,In_641);
nor U680 (N_680,In_27,N_338);
nor U681 (N_681,N_48,In_848);
nand U682 (N_682,N_495,In_32);
and U683 (N_683,N_103,In_219);
nor U684 (N_684,N_477,N_280);
nand U685 (N_685,N_85,N_308);
nor U686 (N_686,N_345,In_109);
and U687 (N_687,N_454,In_935);
nor U688 (N_688,N_391,N_404);
nor U689 (N_689,N_521,N_522);
nand U690 (N_690,In_282,N_592);
xor U691 (N_691,In_235,N_142);
nor U692 (N_692,N_582,In_769);
or U693 (N_693,N_493,N_424);
or U694 (N_694,N_316,N_499);
or U695 (N_695,N_462,In_726);
and U696 (N_696,N_484,In_916);
or U697 (N_697,In_662,N_123);
and U698 (N_698,N_554,N_496);
nand U699 (N_699,N_517,In_208);
nor U700 (N_700,N_162,N_600);
nor U701 (N_701,In_568,N_418);
or U702 (N_702,N_102,N_675);
nor U703 (N_703,N_427,N_304);
or U704 (N_704,N_622,N_163);
or U705 (N_705,N_536,N_697);
nand U706 (N_706,In_944,In_59);
xnor U707 (N_707,N_599,N_690);
nand U708 (N_708,In_429,N_629);
nor U709 (N_709,N_61,N_679);
xnor U710 (N_710,N_457,N_104);
xnor U711 (N_711,N_646,N_188);
nand U712 (N_712,In_813,N_628);
and U713 (N_713,N_492,In_259);
or U714 (N_714,N_140,N_403);
nor U715 (N_715,N_562,N_167);
nor U716 (N_716,N_226,N_214);
nor U717 (N_717,N_545,N_699);
and U718 (N_718,N_652,In_496);
and U719 (N_719,N_643,N_615);
nor U720 (N_720,N_355,N_685);
nand U721 (N_721,In_442,N_407);
and U722 (N_722,N_557,N_694);
and U723 (N_723,N_565,N_482);
xnor U724 (N_724,N_336,In_441);
xor U725 (N_725,In_840,N_620);
xnor U726 (N_726,N_670,N_447);
nand U727 (N_727,N_452,N_603);
xnor U728 (N_728,N_191,N_642);
or U729 (N_729,In_733,N_516);
xor U730 (N_730,N_604,N_356);
and U731 (N_731,N_640,N_526);
and U732 (N_732,N_217,N_663);
and U733 (N_733,N_511,N_80);
or U734 (N_734,In_542,In_398);
xor U735 (N_735,N_524,N_669);
nor U736 (N_736,N_680,In_218);
nand U737 (N_737,N_321,N_529);
xnor U738 (N_738,In_319,In_324);
nor U739 (N_739,N_551,In_732);
and U740 (N_740,In_312,In_883);
nand U741 (N_741,N_510,N_297);
or U742 (N_742,N_543,N_672);
xor U743 (N_743,In_343,N_641);
nor U744 (N_744,N_696,N_157);
nand U745 (N_745,N_683,N_414);
or U746 (N_746,N_626,N_567);
nor U747 (N_747,In_301,N_375);
nor U748 (N_748,N_591,N_346);
xnor U749 (N_749,N_181,N_435);
xnor U750 (N_750,N_689,N_549);
nor U751 (N_751,N_606,N_377);
or U752 (N_752,N_613,In_810);
nor U753 (N_753,N_650,N_420);
xnor U754 (N_754,N_632,N_665);
nor U755 (N_755,N_579,N_548);
and U756 (N_756,N_623,N_682);
nor U757 (N_757,N_677,N_236);
or U758 (N_758,N_367,N_627);
and U759 (N_759,N_357,N_475);
or U760 (N_760,N_596,N_413);
or U761 (N_761,N_331,N_378);
xnor U762 (N_762,In_538,N_631);
or U763 (N_763,N_601,In_36);
nor U764 (N_764,N_353,N_372);
or U765 (N_765,N_563,In_400);
and U766 (N_766,N_412,In_435);
nor U767 (N_767,N_171,N_605);
xor U768 (N_768,N_693,N_471);
and U769 (N_769,N_621,N_330);
and U770 (N_770,N_612,N_630);
or U771 (N_771,N_589,N_648);
and U772 (N_772,N_542,N_584);
or U773 (N_773,N_538,N_246);
or U774 (N_774,N_647,N_513);
xnor U775 (N_775,N_523,N_568);
and U776 (N_776,N_550,N_610);
nand U777 (N_777,N_611,N_691);
xor U778 (N_778,In_364,In_386);
and U779 (N_779,N_537,In_734);
or U780 (N_780,N_686,N_253);
and U781 (N_781,N_474,N_618);
or U782 (N_782,N_608,N_676);
and U783 (N_783,In_815,N_684);
or U784 (N_784,In_524,In_654);
nor U785 (N_785,N_598,In_494);
or U786 (N_786,N_566,In_107);
nor U787 (N_787,N_459,In_677);
or U788 (N_788,N_688,N_249);
and U789 (N_789,N_305,In_416);
and U790 (N_790,N_16,N_687);
xor U791 (N_791,N_664,N_644);
or U792 (N_792,N_645,In_157);
xnor U793 (N_793,N_639,N_638);
or U794 (N_794,N_624,N_487);
xor U795 (N_795,N_560,N_655);
or U796 (N_796,N_520,N_552);
nand U797 (N_797,N_334,N_270);
nand U798 (N_798,In_865,N_678);
xnor U799 (N_799,N_661,N_254);
nand U800 (N_800,N_770,N_754);
xnor U801 (N_801,N_525,N_671);
nand U802 (N_802,N_752,N_743);
xnor U803 (N_803,N_712,N_314);
and U804 (N_804,N_607,N_504);
or U805 (N_805,N_625,N_616);
or U806 (N_806,N_791,N_774);
nand U807 (N_807,N_706,N_469);
nand U808 (N_808,N_219,N_724);
and U809 (N_809,N_720,In_670);
nand U810 (N_810,In_220,N_755);
nor U811 (N_811,N_742,N_570);
xnor U812 (N_812,N_758,N_734);
or U813 (N_813,N_244,N_637);
nor U814 (N_814,N_764,N_722);
nand U815 (N_815,N_718,N_593);
nor U816 (N_816,N_763,N_728);
or U817 (N_817,N_776,In_719);
xor U818 (N_818,N_777,N_732);
nand U819 (N_819,N_744,N_662);
or U820 (N_820,In_583,In_392);
nor U821 (N_821,N_798,N_657);
nor U822 (N_822,N_709,N_634);
xor U823 (N_823,In_265,N_619);
or U824 (N_824,In_422,N_753);
or U825 (N_825,N_617,N_707);
nand U826 (N_826,N_730,N_733);
or U827 (N_827,N_704,N_760);
xor U828 (N_828,In_987,N_653);
and U829 (N_829,N_726,N_797);
or U830 (N_830,N_771,N_773);
or U831 (N_831,N_746,N_767);
and U832 (N_832,N_544,N_446);
xor U833 (N_833,In_919,N_723);
and U834 (N_834,N_710,N_780);
nand U835 (N_835,N_794,N_415);
and U836 (N_836,N_769,N_750);
and U837 (N_837,N_654,N_788);
nor U838 (N_838,N_547,N_740);
nor U839 (N_839,N_674,N_756);
and U840 (N_840,N_792,N_365);
nor U841 (N_841,N_609,N_765);
xnor U842 (N_842,N_700,N_195);
nand U843 (N_843,N_717,N_781);
nor U844 (N_844,N_768,N_45);
and U845 (N_845,N_667,In_336);
and U846 (N_846,N_731,N_793);
nand U847 (N_847,N_737,N_503);
nor U848 (N_848,N_738,N_721);
nand U849 (N_849,N_108,N_711);
nor U850 (N_850,N_745,N_519);
nor U851 (N_851,N_736,N_681);
or U852 (N_852,N_633,N_719);
and U853 (N_853,N_799,N_698);
nand U854 (N_854,N_761,N_695);
nor U855 (N_855,N_741,N_762);
nor U856 (N_856,In_743,N_775);
xnor U857 (N_857,N_635,In_382);
and U858 (N_858,N_782,In_942);
xor U859 (N_859,In_643,N_595);
nand U860 (N_860,N_507,N_660);
nand U861 (N_861,In_579,N_751);
and U862 (N_862,N_166,N_713);
nor U863 (N_863,N_553,N_636);
or U864 (N_864,N_789,In_788);
xnor U865 (N_865,N_485,N_229);
nand U866 (N_866,N_279,N_614);
xnor U867 (N_867,N_329,N_739);
or U868 (N_868,N_651,N_796);
and U869 (N_869,N_749,N_715);
and U870 (N_870,N_714,N_766);
nor U871 (N_871,N_747,N_779);
and U872 (N_872,In_23,In_906);
nor U873 (N_873,N_659,In_372);
nand U874 (N_874,N_115,In_279);
or U875 (N_875,N_790,N_406);
nor U876 (N_876,N_727,N_703);
xor U877 (N_877,N_532,N_725);
xor U878 (N_878,N_778,N_602);
xor U879 (N_879,N_509,N_227);
nor U880 (N_880,N_784,N_748);
and U881 (N_881,N_673,N_772);
nor U882 (N_882,In_222,N_656);
and U883 (N_883,N_787,N_795);
nand U884 (N_884,N_735,N_388);
nand U885 (N_885,N_134,N_701);
and U886 (N_886,N_467,N_658);
nand U887 (N_887,N_786,N_540);
and U888 (N_888,N_561,N_716);
or U889 (N_889,N_73,In_536);
xor U890 (N_890,N_785,N_729);
nor U891 (N_891,N_708,N_702);
and U892 (N_892,N_692,N_757);
nand U893 (N_893,N_759,N_573);
xnor U894 (N_894,N_461,N_649);
or U895 (N_895,N_225,N_668);
xor U896 (N_896,In_861,N_783);
nand U897 (N_897,N_490,N_318);
nand U898 (N_898,N_576,N_300);
xor U899 (N_899,N_666,N_705);
nand U900 (N_900,N_855,N_822);
nor U901 (N_901,N_870,N_899);
nor U902 (N_902,N_872,N_812);
nand U903 (N_903,N_864,N_851);
nor U904 (N_904,N_847,N_805);
nand U905 (N_905,N_849,N_852);
or U906 (N_906,N_816,N_818);
nor U907 (N_907,N_843,N_842);
nand U908 (N_908,N_882,N_840);
nand U909 (N_909,N_820,N_827);
nand U910 (N_910,N_832,N_897);
or U911 (N_911,N_811,N_825);
and U912 (N_912,N_808,N_848);
nand U913 (N_913,N_859,N_844);
xnor U914 (N_914,N_831,N_880);
or U915 (N_915,N_815,N_821);
and U916 (N_916,N_846,N_858);
xnor U917 (N_917,N_857,N_850);
nand U918 (N_918,N_861,N_837);
or U919 (N_919,N_817,N_854);
nor U920 (N_920,N_838,N_841);
nor U921 (N_921,N_856,N_813);
xor U922 (N_922,N_892,N_835);
xnor U923 (N_923,N_868,N_875);
nand U924 (N_924,N_881,N_889);
or U925 (N_925,N_874,N_886);
nor U926 (N_926,N_804,N_833);
or U927 (N_927,N_823,N_884);
nand U928 (N_928,N_878,N_873);
nor U929 (N_929,N_862,N_800);
xnor U930 (N_930,N_891,N_887);
nor U931 (N_931,N_829,N_866);
xnor U932 (N_932,N_863,N_890);
or U933 (N_933,N_807,N_893);
or U934 (N_934,N_895,N_865);
or U935 (N_935,N_826,N_806);
xor U936 (N_936,N_876,N_885);
and U937 (N_937,N_869,N_853);
or U938 (N_938,N_803,N_896);
and U939 (N_939,N_819,N_860);
or U940 (N_940,N_888,N_834);
xor U941 (N_941,N_883,N_879);
nor U942 (N_942,N_802,N_801);
nand U943 (N_943,N_824,N_845);
or U944 (N_944,N_894,N_810);
or U945 (N_945,N_867,N_898);
xor U946 (N_946,N_814,N_877);
nand U947 (N_947,N_809,N_830);
nand U948 (N_948,N_836,N_839);
nand U949 (N_949,N_828,N_871);
xnor U950 (N_950,N_834,N_868);
or U951 (N_951,N_838,N_813);
and U952 (N_952,N_833,N_875);
or U953 (N_953,N_861,N_852);
or U954 (N_954,N_859,N_850);
xnor U955 (N_955,N_812,N_851);
or U956 (N_956,N_821,N_899);
or U957 (N_957,N_828,N_876);
and U958 (N_958,N_897,N_854);
nor U959 (N_959,N_834,N_845);
nand U960 (N_960,N_882,N_820);
or U961 (N_961,N_811,N_849);
nor U962 (N_962,N_812,N_809);
nand U963 (N_963,N_889,N_828);
xor U964 (N_964,N_859,N_892);
and U965 (N_965,N_806,N_848);
or U966 (N_966,N_859,N_843);
xnor U967 (N_967,N_802,N_868);
and U968 (N_968,N_826,N_823);
nand U969 (N_969,N_890,N_825);
or U970 (N_970,N_851,N_867);
xor U971 (N_971,N_830,N_857);
nand U972 (N_972,N_827,N_818);
and U973 (N_973,N_832,N_800);
nand U974 (N_974,N_849,N_805);
nand U975 (N_975,N_841,N_854);
and U976 (N_976,N_823,N_817);
or U977 (N_977,N_825,N_879);
and U978 (N_978,N_839,N_856);
or U979 (N_979,N_850,N_808);
xnor U980 (N_980,N_852,N_869);
nand U981 (N_981,N_820,N_898);
nor U982 (N_982,N_823,N_829);
nor U983 (N_983,N_869,N_884);
or U984 (N_984,N_895,N_879);
or U985 (N_985,N_851,N_827);
xor U986 (N_986,N_879,N_804);
or U987 (N_987,N_849,N_812);
and U988 (N_988,N_891,N_826);
nand U989 (N_989,N_815,N_843);
or U990 (N_990,N_816,N_801);
or U991 (N_991,N_896,N_893);
nand U992 (N_992,N_851,N_842);
nand U993 (N_993,N_885,N_804);
and U994 (N_994,N_868,N_806);
xor U995 (N_995,N_868,N_877);
or U996 (N_996,N_825,N_847);
xnor U997 (N_997,N_875,N_895);
or U998 (N_998,N_879,N_888);
xor U999 (N_999,N_824,N_803);
nand U1000 (N_1000,N_960,N_997);
xor U1001 (N_1001,N_966,N_957);
or U1002 (N_1002,N_953,N_906);
xnor U1003 (N_1003,N_900,N_927);
or U1004 (N_1004,N_998,N_921);
nor U1005 (N_1005,N_995,N_947);
or U1006 (N_1006,N_907,N_971);
nor U1007 (N_1007,N_990,N_976);
and U1008 (N_1008,N_996,N_929);
and U1009 (N_1009,N_949,N_977);
or U1010 (N_1010,N_931,N_994);
nand U1011 (N_1011,N_986,N_923);
or U1012 (N_1012,N_909,N_930);
and U1013 (N_1013,N_926,N_959);
nor U1014 (N_1014,N_914,N_924);
or U1015 (N_1015,N_991,N_941);
and U1016 (N_1016,N_967,N_911);
or U1017 (N_1017,N_963,N_904);
xnor U1018 (N_1018,N_938,N_937);
and U1019 (N_1019,N_970,N_917);
or U1020 (N_1020,N_942,N_928);
and U1021 (N_1021,N_969,N_939);
nor U1022 (N_1022,N_962,N_903);
xor U1023 (N_1023,N_908,N_979);
xnor U1024 (N_1024,N_918,N_919);
nor U1025 (N_1025,N_952,N_932);
or U1026 (N_1026,N_987,N_940);
xnor U1027 (N_1027,N_999,N_951);
nand U1028 (N_1028,N_950,N_975);
nand U1029 (N_1029,N_978,N_961);
nor U1030 (N_1030,N_905,N_913);
xnor U1031 (N_1031,N_992,N_901);
nor U1032 (N_1032,N_902,N_989);
xnor U1033 (N_1033,N_933,N_958);
and U1034 (N_1034,N_988,N_980);
xor U1035 (N_1035,N_915,N_935);
nand U1036 (N_1036,N_965,N_982);
and U1037 (N_1037,N_993,N_936);
and U1038 (N_1038,N_981,N_956);
or U1039 (N_1039,N_955,N_985);
and U1040 (N_1040,N_943,N_920);
xor U1041 (N_1041,N_910,N_946);
and U1042 (N_1042,N_954,N_973);
xor U1043 (N_1043,N_983,N_968);
nor U1044 (N_1044,N_922,N_964);
xnor U1045 (N_1045,N_925,N_984);
nand U1046 (N_1046,N_945,N_912);
and U1047 (N_1047,N_944,N_972);
xnor U1048 (N_1048,N_916,N_948);
nor U1049 (N_1049,N_934,N_974);
nor U1050 (N_1050,N_965,N_935);
nand U1051 (N_1051,N_937,N_982);
or U1052 (N_1052,N_946,N_909);
xor U1053 (N_1053,N_981,N_999);
nor U1054 (N_1054,N_906,N_931);
xor U1055 (N_1055,N_990,N_906);
nand U1056 (N_1056,N_926,N_984);
or U1057 (N_1057,N_927,N_920);
or U1058 (N_1058,N_942,N_920);
xor U1059 (N_1059,N_900,N_987);
nand U1060 (N_1060,N_975,N_907);
nand U1061 (N_1061,N_911,N_994);
nor U1062 (N_1062,N_970,N_959);
and U1063 (N_1063,N_900,N_981);
nor U1064 (N_1064,N_927,N_907);
and U1065 (N_1065,N_924,N_995);
xnor U1066 (N_1066,N_939,N_933);
nand U1067 (N_1067,N_959,N_952);
or U1068 (N_1068,N_963,N_926);
or U1069 (N_1069,N_915,N_968);
xnor U1070 (N_1070,N_925,N_908);
nor U1071 (N_1071,N_961,N_931);
nor U1072 (N_1072,N_966,N_988);
xor U1073 (N_1073,N_903,N_921);
nor U1074 (N_1074,N_955,N_904);
nor U1075 (N_1075,N_902,N_939);
nor U1076 (N_1076,N_922,N_965);
and U1077 (N_1077,N_960,N_993);
xnor U1078 (N_1078,N_907,N_968);
xnor U1079 (N_1079,N_962,N_915);
xnor U1080 (N_1080,N_911,N_938);
or U1081 (N_1081,N_902,N_977);
and U1082 (N_1082,N_942,N_972);
or U1083 (N_1083,N_992,N_934);
xnor U1084 (N_1084,N_963,N_929);
xnor U1085 (N_1085,N_945,N_957);
xnor U1086 (N_1086,N_982,N_908);
nor U1087 (N_1087,N_945,N_982);
nor U1088 (N_1088,N_938,N_907);
and U1089 (N_1089,N_921,N_923);
nand U1090 (N_1090,N_971,N_929);
nand U1091 (N_1091,N_988,N_958);
nor U1092 (N_1092,N_985,N_913);
nand U1093 (N_1093,N_958,N_965);
or U1094 (N_1094,N_919,N_936);
xnor U1095 (N_1095,N_914,N_969);
xor U1096 (N_1096,N_913,N_977);
or U1097 (N_1097,N_932,N_943);
nor U1098 (N_1098,N_945,N_971);
nand U1099 (N_1099,N_962,N_934);
and U1100 (N_1100,N_1094,N_1017);
nand U1101 (N_1101,N_1092,N_1077);
and U1102 (N_1102,N_1011,N_1057);
nand U1103 (N_1103,N_1071,N_1040);
nor U1104 (N_1104,N_1073,N_1021);
nor U1105 (N_1105,N_1086,N_1093);
or U1106 (N_1106,N_1062,N_1067);
xnor U1107 (N_1107,N_1048,N_1016);
or U1108 (N_1108,N_1045,N_1036);
xor U1109 (N_1109,N_1069,N_1004);
nand U1110 (N_1110,N_1090,N_1027);
and U1111 (N_1111,N_1078,N_1008);
and U1112 (N_1112,N_1015,N_1000);
nand U1113 (N_1113,N_1031,N_1097);
or U1114 (N_1114,N_1025,N_1059);
nor U1115 (N_1115,N_1074,N_1038);
xor U1116 (N_1116,N_1032,N_1005);
xor U1117 (N_1117,N_1009,N_1047);
nor U1118 (N_1118,N_1066,N_1099);
or U1119 (N_1119,N_1013,N_1055);
or U1120 (N_1120,N_1007,N_1024);
and U1121 (N_1121,N_1020,N_1001);
nand U1122 (N_1122,N_1050,N_1070);
or U1123 (N_1123,N_1030,N_1085);
nor U1124 (N_1124,N_1068,N_1053);
xor U1125 (N_1125,N_1054,N_1035);
nor U1126 (N_1126,N_1081,N_1010);
and U1127 (N_1127,N_1026,N_1064);
nor U1128 (N_1128,N_1044,N_1003);
and U1129 (N_1129,N_1051,N_1076);
and U1130 (N_1130,N_1046,N_1091);
nor U1131 (N_1131,N_1043,N_1063);
xnor U1132 (N_1132,N_1095,N_1056);
nor U1133 (N_1133,N_1072,N_1006);
or U1134 (N_1134,N_1034,N_1037);
xnor U1135 (N_1135,N_1002,N_1058);
or U1136 (N_1136,N_1088,N_1079);
nor U1137 (N_1137,N_1052,N_1018);
nor U1138 (N_1138,N_1041,N_1098);
and U1139 (N_1139,N_1019,N_1049);
nor U1140 (N_1140,N_1023,N_1082);
xor U1141 (N_1141,N_1061,N_1096);
nand U1142 (N_1142,N_1022,N_1014);
and U1143 (N_1143,N_1083,N_1089);
nor U1144 (N_1144,N_1060,N_1012);
nand U1145 (N_1145,N_1087,N_1039);
xnor U1146 (N_1146,N_1029,N_1028);
or U1147 (N_1147,N_1075,N_1080);
or U1148 (N_1148,N_1084,N_1033);
nor U1149 (N_1149,N_1042,N_1065);
nor U1150 (N_1150,N_1041,N_1016);
or U1151 (N_1151,N_1016,N_1080);
or U1152 (N_1152,N_1068,N_1084);
and U1153 (N_1153,N_1042,N_1073);
nand U1154 (N_1154,N_1007,N_1096);
xor U1155 (N_1155,N_1079,N_1038);
xnor U1156 (N_1156,N_1009,N_1067);
xor U1157 (N_1157,N_1009,N_1090);
or U1158 (N_1158,N_1025,N_1075);
and U1159 (N_1159,N_1092,N_1007);
nand U1160 (N_1160,N_1091,N_1021);
xnor U1161 (N_1161,N_1080,N_1038);
or U1162 (N_1162,N_1032,N_1092);
and U1163 (N_1163,N_1003,N_1002);
and U1164 (N_1164,N_1011,N_1067);
nand U1165 (N_1165,N_1012,N_1018);
and U1166 (N_1166,N_1007,N_1084);
xor U1167 (N_1167,N_1019,N_1073);
nand U1168 (N_1168,N_1099,N_1002);
xor U1169 (N_1169,N_1090,N_1047);
nor U1170 (N_1170,N_1053,N_1092);
and U1171 (N_1171,N_1082,N_1089);
nor U1172 (N_1172,N_1022,N_1050);
and U1173 (N_1173,N_1087,N_1045);
and U1174 (N_1174,N_1084,N_1046);
nor U1175 (N_1175,N_1065,N_1053);
or U1176 (N_1176,N_1065,N_1011);
nand U1177 (N_1177,N_1029,N_1071);
nor U1178 (N_1178,N_1084,N_1006);
nor U1179 (N_1179,N_1056,N_1028);
nor U1180 (N_1180,N_1096,N_1085);
nor U1181 (N_1181,N_1063,N_1036);
or U1182 (N_1182,N_1002,N_1059);
nand U1183 (N_1183,N_1021,N_1095);
nor U1184 (N_1184,N_1044,N_1048);
xnor U1185 (N_1185,N_1094,N_1084);
xnor U1186 (N_1186,N_1054,N_1077);
nand U1187 (N_1187,N_1009,N_1045);
and U1188 (N_1188,N_1082,N_1035);
and U1189 (N_1189,N_1076,N_1028);
nor U1190 (N_1190,N_1053,N_1022);
xnor U1191 (N_1191,N_1004,N_1035);
or U1192 (N_1192,N_1091,N_1025);
nor U1193 (N_1193,N_1025,N_1001);
nor U1194 (N_1194,N_1084,N_1052);
nor U1195 (N_1195,N_1098,N_1077);
and U1196 (N_1196,N_1062,N_1066);
nor U1197 (N_1197,N_1037,N_1032);
or U1198 (N_1198,N_1044,N_1063);
or U1199 (N_1199,N_1002,N_1088);
xor U1200 (N_1200,N_1110,N_1190);
nand U1201 (N_1201,N_1140,N_1189);
or U1202 (N_1202,N_1156,N_1160);
or U1203 (N_1203,N_1132,N_1158);
or U1204 (N_1204,N_1192,N_1131);
and U1205 (N_1205,N_1186,N_1122);
nor U1206 (N_1206,N_1143,N_1180);
or U1207 (N_1207,N_1134,N_1157);
nand U1208 (N_1208,N_1181,N_1178);
and U1209 (N_1209,N_1149,N_1197);
xor U1210 (N_1210,N_1126,N_1121);
nand U1211 (N_1211,N_1144,N_1108);
nand U1212 (N_1212,N_1135,N_1109);
xor U1213 (N_1213,N_1103,N_1127);
or U1214 (N_1214,N_1139,N_1111);
and U1215 (N_1215,N_1129,N_1137);
or U1216 (N_1216,N_1173,N_1183);
nor U1217 (N_1217,N_1145,N_1107);
and U1218 (N_1218,N_1123,N_1138);
or U1219 (N_1219,N_1136,N_1185);
nor U1220 (N_1220,N_1118,N_1104);
or U1221 (N_1221,N_1124,N_1174);
nand U1222 (N_1222,N_1198,N_1112);
xor U1223 (N_1223,N_1168,N_1142);
xnor U1224 (N_1224,N_1167,N_1120);
nor U1225 (N_1225,N_1102,N_1128);
or U1226 (N_1226,N_1147,N_1155);
nand U1227 (N_1227,N_1172,N_1117);
xnor U1228 (N_1228,N_1159,N_1170);
and U1229 (N_1229,N_1133,N_1164);
nor U1230 (N_1230,N_1199,N_1106);
nor U1231 (N_1231,N_1169,N_1105);
xor U1232 (N_1232,N_1196,N_1165);
and U1233 (N_1233,N_1154,N_1148);
and U1234 (N_1234,N_1179,N_1125);
or U1235 (N_1235,N_1113,N_1130);
or U1236 (N_1236,N_1187,N_1182);
and U1237 (N_1237,N_1176,N_1119);
xnor U1238 (N_1238,N_1177,N_1194);
and U1239 (N_1239,N_1146,N_1184);
nand U1240 (N_1240,N_1150,N_1171);
nor U1241 (N_1241,N_1191,N_1141);
nand U1242 (N_1242,N_1188,N_1195);
nand U1243 (N_1243,N_1162,N_1175);
or U1244 (N_1244,N_1114,N_1153);
xor U1245 (N_1245,N_1152,N_1166);
nor U1246 (N_1246,N_1116,N_1151);
or U1247 (N_1247,N_1193,N_1163);
or U1248 (N_1248,N_1101,N_1115);
and U1249 (N_1249,N_1100,N_1161);
and U1250 (N_1250,N_1130,N_1161);
xnor U1251 (N_1251,N_1110,N_1129);
and U1252 (N_1252,N_1168,N_1169);
nand U1253 (N_1253,N_1173,N_1159);
and U1254 (N_1254,N_1176,N_1188);
or U1255 (N_1255,N_1160,N_1188);
xor U1256 (N_1256,N_1139,N_1150);
and U1257 (N_1257,N_1100,N_1158);
and U1258 (N_1258,N_1187,N_1127);
nand U1259 (N_1259,N_1102,N_1116);
nor U1260 (N_1260,N_1175,N_1146);
or U1261 (N_1261,N_1134,N_1123);
xor U1262 (N_1262,N_1100,N_1109);
nor U1263 (N_1263,N_1174,N_1163);
nor U1264 (N_1264,N_1112,N_1134);
or U1265 (N_1265,N_1144,N_1185);
nand U1266 (N_1266,N_1105,N_1172);
or U1267 (N_1267,N_1131,N_1159);
xor U1268 (N_1268,N_1149,N_1180);
nor U1269 (N_1269,N_1152,N_1108);
nand U1270 (N_1270,N_1176,N_1123);
nor U1271 (N_1271,N_1117,N_1120);
xor U1272 (N_1272,N_1169,N_1100);
or U1273 (N_1273,N_1114,N_1181);
xor U1274 (N_1274,N_1178,N_1156);
nor U1275 (N_1275,N_1158,N_1194);
and U1276 (N_1276,N_1124,N_1197);
and U1277 (N_1277,N_1146,N_1167);
nand U1278 (N_1278,N_1104,N_1111);
or U1279 (N_1279,N_1183,N_1168);
and U1280 (N_1280,N_1115,N_1117);
or U1281 (N_1281,N_1148,N_1184);
xor U1282 (N_1282,N_1124,N_1188);
nor U1283 (N_1283,N_1151,N_1185);
nor U1284 (N_1284,N_1120,N_1130);
or U1285 (N_1285,N_1191,N_1185);
xor U1286 (N_1286,N_1118,N_1126);
xnor U1287 (N_1287,N_1119,N_1140);
nand U1288 (N_1288,N_1196,N_1158);
xnor U1289 (N_1289,N_1157,N_1181);
and U1290 (N_1290,N_1112,N_1108);
nand U1291 (N_1291,N_1120,N_1108);
xor U1292 (N_1292,N_1109,N_1170);
xnor U1293 (N_1293,N_1107,N_1187);
nor U1294 (N_1294,N_1192,N_1114);
nand U1295 (N_1295,N_1172,N_1114);
or U1296 (N_1296,N_1191,N_1157);
nand U1297 (N_1297,N_1194,N_1142);
and U1298 (N_1298,N_1161,N_1160);
nor U1299 (N_1299,N_1198,N_1108);
or U1300 (N_1300,N_1233,N_1270);
or U1301 (N_1301,N_1277,N_1248);
nor U1302 (N_1302,N_1272,N_1247);
nor U1303 (N_1303,N_1295,N_1261);
and U1304 (N_1304,N_1212,N_1210);
and U1305 (N_1305,N_1296,N_1227);
xnor U1306 (N_1306,N_1246,N_1282);
xor U1307 (N_1307,N_1240,N_1288);
nand U1308 (N_1308,N_1220,N_1285);
nor U1309 (N_1309,N_1278,N_1267);
or U1310 (N_1310,N_1203,N_1289);
and U1311 (N_1311,N_1218,N_1224);
or U1312 (N_1312,N_1244,N_1258);
nor U1313 (N_1313,N_1287,N_1207);
and U1314 (N_1314,N_1260,N_1259);
nor U1315 (N_1315,N_1226,N_1251);
or U1316 (N_1316,N_1235,N_1292);
nor U1317 (N_1317,N_1275,N_1214);
xor U1318 (N_1318,N_1294,N_1274);
nand U1319 (N_1319,N_1284,N_1256);
nor U1320 (N_1320,N_1269,N_1222);
nor U1321 (N_1321,N_1201,N_1252);
xor U1322 (N_1322,N_1211,N_1281);
and U1323 (N_1323,N_1209,N_1290);
nor U1324 (N_1324,N_1208,N_1228);
nor U1325 (N_1325,N_1242,N_1216);
nand U1326 (N_1326,N_1245,N_1230);
and U1327 (N_1327,N_1223,N_1239);
and U1328 (N_1328,N_1299,N_1243);
nand U1329 (N_1329,N_1279,N_1225);
nor U1330 (N_1330,N_1297,N_1262);
or U1331 (N_1331,N_1202,N_1205);
nand U1332 (N_1332,N_1241,N_1291);
and U1333 (N_1333,N_1221,N_1280);
nand U1334 (N_1334,N_1236,N_1231);
and U1335 (N_1335,N_1253,N_1217);
nor U1336 (N_1336,N_1298,N_1286);
nor U1337 (N_1337,N_1238,N_1257);
nor U1338 (N_1338,N_1213,N_1215);
or U1339 (N_1339,N_1255,N_1249);
xnor U1340 (N_1340,N_1234,N_1232);
or U1341 (N_1341,N_1237,N_1254);
and U1342 (N_1342,N_1264,N_1219);
or U1343 (N_1343,N_1229,N_1204);
and U1344 (N_1344,N_1250,N_1206);
nor U1345 (N_1345,N_1271,N_1200);
nand U1346 (N_1346,N_1293,N_1265);
nor U1347 (N_1347,N_1263,N_1283);
nor U1348 (N_1348,N_1276,N_1273);
nor U1349 (N_1349,N_1268,N_1266);
nor U1350 (N_1350,N_1292,N_1210);
or U1351 (N_1351,N_1287,N_1221);
or U1352 (N_1352,N_1274,N_1249);
and U1353 (N_1353,N_1238,N_1260);
and U1354 (N_1354,N_1294,N_1296);
xnor U1355 (N_1355,N_1220,N_1257);
nand U1356 (N_1356,N_1218,N_1211);
and U1357 (N_1357,N_1267,N_1203);
and U1358 (N_1358,N_1269,N_1292);
nor U1359 (N_1359,N_1238,N_1291);
xnor U1360 (N_1360,N_1201,N_1205);
nand U1361 (N_1361,N_1281,N_1262);
nor U1362 (N_1362,N_1265,N_1211);
xor U1363 (N_1363,N_1267,N_1213);
and U1364 (N_1364,N_1299,N_1290);
nor U1365 (N_1365,N_1287,N_1267);
xor U1366 (N_1366,N_1270,N_1200);
nor U1367 (N_1367,N_1276,N_1203);
or U1368 (N_1368,N_1232,N_1257);
xor U1369 (N_1369,N_1251,N_1201);
xor U1370 (N_1370,N_1258,N_1205);
nand U1371 (N_1371,N_1232,N_1240);
nand U1372 (N_1372,N_1246,N_1234);
nand U1373 (N_1373,N_1261,N_1232);
and U1374 (N_1374,N_1246,N_1254);
xor U1375 (N_1375,N_1269,N_1226);
xor U1376 (N_1376,N_1265,N_1203);
and U1377 (N_1377,N_1290,N_1294);
nand U1378 (N_1378,N_1241,N_1240);
nand U1379 (N_1379,N_1227,N_1271);
xnor U1380 (N_1380,N_1208,N_1232);
nor U1381 (N_1381,N_1284,N_1205);
xnor U1382 (N_1382,N_1298,N_1259);
nor U1383 (N_1383,N_1228,N_1261);
xor U1384 (N_1384,N_1270,N_1274);
xnor U1385 (N_1385,N_1224,N_1262);
xor U1386 (N_1386,N_1273,N_1261);
xor U1387 (N_1387,N_1278,N_1256);
or U1388 (N_1388,N_1277,N_1220);
xnor U1389 (N_1389,N_1201,N_1259);
xnor U1390 (N_1390,N_1233,N_1253);
and U1391 (N_1391,N_1229,N_1262);
nand U1392 (N_1392,N_1273,N_1246);
xor U1393 (N_1393,N_1225,N_1274);
nand U1394 (N_1394,N_1224,N_1248);
nor U1395 (N_1395,N_1254,N_1249);
xnor U1396 (N_1396,N_1275,N_1292);
xor U1397 (N_1397,N_1247,N_1202);
nand U1398 (N_1398,N_1251,N_1221);
xor U1399 (N_1399,N_1286,N_1267);
xnor U1400 (N_1400,N_1377,N_1381);
nor U1401 (N_1401,N_1395,N_1322);
and U1402 (N_1402,N_1343,N_1311);
xor U1403 (N_1403,N_1314,N_1359);
nor U1404 (N_1404,N_1386,N_1327);
or U1405 (N_1405,N_1358,N_1324);
nor U1406 (N_1406,N_1375,N_1387);
or U1407 (N_1407,N_1309,N_1344);
nor U1408 (N_1408,N_1396,N_1393);
or U1409 (N_1409,N_1326,N_1341);
and U1410 (N_1410,N_1329,N_1345);
or U1411 (N_1411,N_1335,N_1331);
and U1412 (N_1412,N_1370,N_1376);
nor U1413 (N_1413,N_1348,N_1338);
xor U1414 (N_1414,N_1332,N_1334);
or U1415 (N_1415,N_1354,N_1391);
nand U1416 (N_1416,N_1360,N_1306);
xnor U1417 (N_1417,N_1301,N_1371);
nand U1418 (N_1418,N_1365,N_1351);
xor U1419 (N_1419,N_1398,N_1328);
nor U1420 (N_1420,N_1361,N_1388);
or U1421 (N_1421,N_1353,N_1342);
xor U1422 (N_1422,N_1382,N_1355);
nand U1423 (N_1423,N_1369,N_1374);
or U1424 (N_1424,N_1333,N_1362);
nand U1425 (N_1425,N_1385,N_1321);
and U1426 (N_1426,N_1356,N_1317);
and U1427 (N_1427,N_1357,N_1378);
and U1428 (N_1428,N_1364,N_1316);
nor U1429 (N_1429,N_1330,N_1313);
and U1430 (N_1430,N_1363,N_1302);
nor U1431 (N_1431,N_1336,N_1392);
nor U1432 (N_1432,N_1315,N_1350);
or U1433 (N_1433,N_1352,N_1397);
nor U1434 (N_1434,N_1303,N_1337);
or U1435 (N_1435,N_1383,N_1305);
nor U1436 (N_1436,N_1380,N_1325);
or U1437 (N_1437,N_1340,N_1389);
and U1438 (N_1438,N_1384,N_1372);
xor U1439 (N_1439,N_1339,N_1304);
or U1440 (N_1440,N_1373,N_1394);
or U1441 (N_1441,N_1347,N_1366);
and U1442 (N_1442,N_1310,N_1368);
xnor U1443 (N_1443,N_1300,N_1318);
nand U1444 (N_1444,N_1308,N_1319);
xnor U1445 (N_1445,N_1307,N_1312);
nand U1446 (N_1446,N_1323,N_1399);
and U1447 (N_1447,N_1390,N_1349);
xnor U1448 (N_1448,N_1320,N_1367);
and U1449 (N_1449,N_1379,N_1346);
or U1450 (N_1450,N_1308,N_1314);
or U1451 (N_1451,N_1311,N_1328);
xnor U1452 (N_1452,N_1374,N_1349);
and U1453 (N_1453,N_1335,N_1347);
nor U1454 (N_1454,N_1373,N_1392);
and U1455 (N_1455,N_1320,N_1342);
nor U1456 (N_1456,N_1347,N_1336);
nor U1457 (N_1457,N_1389,N_1343);
nand U1458 (N_1458,N_1342,N_1375);
xnor U1459 (N_1459,N_1341,N_1351);
and U1460 (N_1460,N_1351,N_1352);
xnor U1461 (N_1461,N_1327,N_1303);
nor U1462 (N_1462,N_1321,N_1362);
and U1463 (N_1463,N_1316,N_1375);
nand U1464 (N_1464,N_1355,N_1331);
xnor U1465 (N_1465,N_1312,N_1343);
or U1466 (N_1466,N_1329,N_1367);
xnor U1467 (N_1467,N_1373,N_1302);
and U1468 (N_1468,N_1352,N_1323);
nor U1469 (N_1469,N_1345,N_1381);
xnor U1470 (N_1470,N_1331,N_1390);
or U1471 (N_1471,N_1322,N_1341);
nand U1472 (N_1472,N_1374,N_1312);
xor U1473 (N_1473,N_1378,N_1335);
nor U1474 (N_1474,N_1308,N_1380);
xor U1475 (N_1475,N_1362,N_1354);
nor U1476 (N_1476,N_1321,N_1302);
nand U1477 (N_1477,N_1340,N_1368);
nor U1478 (N_1478,N_1304,N_1340);
nand U1479 (N_1479,N_1375,N_1361);
xor U1480 (N_1480,N_1390,N_1303);
nand U1481 (N_1481,N_1334,N_1371);
nor U1482 (N_1482,N_1359,N_1334);
nor U1483 (N_1483,N_1353,N_1375);
xor U1484 (N_1484,N_1300,N_1306);
nor U1485 (N_1485,N_1346,N_1389);
and U1486 (N_1486,N_1348,N_1315);
nand U1487 (N_1487,N_1360,N_1351);
and U1488 (N_1488,N_1383,N_1379);
and U1489 (N_1489,N_1365,N_1350);
nand U1490 (N_1490,N_1319,N_1394);
and U1491 (N_1491,N_1304,N_1316);
nand U1492 (N_1492,N_1305,N_1379);
xor U1493 (N_1493,N_1304,N_1305);
nand U1494 (N_1494,N_1390,N_1375);
nand U1495 (N_1495,N_1377,N_1346);
or U1496 (N_1496,N_1365,N_1313);
and U1497 (N_1497,N_1383,N_1326);
and U1498 (N_1498,N_1357,N_1339);
xnor U1499 (N_1499,N_1326,N_1314);
xnor U1500 (N_1500,N_1487,N_1467);
nand U1501 (N_1501,N_1430,N_1400);
xor U1502 (N_1502,N_1417,N_1488);
nand U1503 (N_1503,N_1452,N_1440);
xnor U1504 (N_1504,N_1493,N_1425);
xnor U1505 (N_1505,N_1466,N_1406);
or U1506 (N_1506,N_1427,N_1485);
or U1507 (N_1507,N_1459,N_1473);
nor U1508 (N_1508,N_1471,N_1477);
and U1509 (N_1509,N_1486,N_1450);
nand U1510 (N_1510,N_1429,N_1476);
or U1511 (N_1511,N_1496,N_1423);
and U1512 (N_1512,N_1434,N_1437);
xnor U1513 (N_1513,N_1443,N_1461);
nor U1514 (N_1514,N_1428,N_1419);
xnor U1515 (N_1515,N_1449,N_1465);
nor U1516 (N_1516,N_1411,N_1405);
nor U1517 (N_1517,N_1447,N_1478);
xnor U1518 (N_1518,N_1495,N_1448);
or U1519 (N_1519,N_1414,N_1499);
nor U1520 (N_1520,N_1455,N_1446);
xnor U1521 (N_1521,N_1491,N_1444);
xor U1522 (N_1522,N_1462,N_1490);
or U1523 (N_1523,N_1432,N_1407);
xnor U1524 (N_1524,N_1460,N_1475);
or U1525 (N_1525,N_1409,N_1402);
and U1526 (N_1526,N_1484,N_1492);
and U1527 (N_1527,N_1472,N_1458);
or U1528 (N_1528,N_1479,N_1463);
and U1529 (N_1529,N_1420,N_1404);
nor U1530 (N_1530,N_1439,N_1415);
nand U1531 (N_1531,N_1468,N_1403);
nand U1532 (N_1532,N_1453,N_1451);
nand U1533 (N_1533,N_1498,N_1445);
and U1534 (N_1534,N_1436,N_1481);
xor U1535 (N_1535,N_1438,N_1422);
nor U1536 (N_1536,N_1483,N_1454);
or U1537 (N_1537,N_1497,N_1426);
nand U1538 (N_1538,N_1412,N_1469);
xor U1539 (N_1539,N_1474,N_1480);
xnor U1540 (N_1540,N_1424,N_1431);
or U1541 (N_1541,N_1442,N_1421);
nand U1542 (N_1542,N_1457,N_1416);
and U1543 (N_1543,N_1433,N_1401);
and U1544 (N_1544,N_1494,N_1418);
xor U1545 (N_1545,N_1482,N_1464);
and U1546 (N_1546,N_1435,N_1470);
or U1547 (N_1547,N_1456,N_1410);
nor U1548 (N_1548,N_1489,N_1408);
nor U1549 (N_1549,N_1413,N_1441);
nand U1550 (N_1550,N_1436,N_1485);
nor U1551 (N_1551,N_1479,N_1442);
nand U1552 (N_1552,N_1467,N_1450);
nor U1553 (N_1553,N_1480,N_1467);
nor U1554 (N_1554,N_1409,N_1449);
xor U1555 (N_1555,N_1410,N_1463);
nor U1556 (N_1556,N_1460,N_1458);
xor U1557 (N_1557,N_1417,N_1457);
and U1558 (N_1558,N_1423,N_1443);
nor U1559 (N_1559,N_1446,N_1406);
nand U1560 (N_1560,N_1413,N_1426);
nand U1561 (N_1561,N_1455,N_1474);
or U1562 (N_1562,N_1445,N_1471);
nor U1563 (N_1563,N_1418,N_1496);
or U1564 (N_1564,N_1479,N_1441);
nand U1565 (N_1565,N_1491,N_1431);
nor U1566 (N_1566,N_1478,N_1411);
or U1567 (N_1567,N_1432,N_1413);
or U1568 (N_1568,N_1485,N_1434);
nand U1569 (N_1569,N_1483,N_1414);
nand U1570 (N_1570,N_1430,N_1414);
nor U1571 (N_1571,N_1438,N_1498);
nor U1572 (N_1572,N_1448,N_1455);
or U1573 (N_1573,N_1492,N_1465);
or U1574 (N_1574,N_1407,N_1400);
nor U1575 (N_1575,N_1447,N_1453);
nor U1576 (N_1576,N_1451,N_1447);
or U1577 (N_1577,N_1481,N_1450);
nand U1578 (N_1578,N_1463,N_1483);
nor U1579 (N_1579,N_1473,N_1419);
nand U1580 (N_1580,N_1465,N_1451);
nor U1581 (N_1581,N_1429,N_1440);
and U1582 (N_1582,N_1428,N_1400);
and U1583 (N_1583,N_1475,N_1451);
or U1584 (N_1584,N_1483,N_1404);
nand U1585 (N_1585,N_1408,N_1473);
or U1586 (N_1586,N_1465,N_1444);
nor U1587 (N_1587,N_1433,N_1482);
or U1588 (N_1588,N_1432,N_1487);
or U1589 (N_1589,N_1419,N_1426);
nand U1590 (N_1590,N_1433,N_1414);
or U1591 (N_1591,N_1475,N_1426);
nand U1592 (N_1592,N_1424,N_1455);
and U1593 (N_1593,N_1466,N_1432);
xnor U1594 (N_1594,N_1494,N_1454);
and U1595 (N_1595,N_1467,N_1431);
and U1596 (N_1596,N_1483,N_1458);
or U1597 (N_1597,N_1455,N_1494);
or U1598 (N_1598,N_1415,N_1408);
nand U1599 (N_1599,N_1490,N_1433);
xnor U1600 (N_1600,N_1524,N_1585);
nand U1601 (N_1601,N_1553,N_1588);
xor U1602 (N_1602,N_1583,N_1574);
nand U1603 (N_1603,N_1577,N_1535);
or U1604 (N_1604,N_1506,N_1572);
nor U1605 (N_1605,N_1541,N_1537);
nand U1606 (N_1606,N_1550,N_1536);
or U1607 (N_1607,N_1549,N_1545);
xnor U1608 (N_1608,N_1519,N_1573);
nor U1609 (N_1609,N_1507,N_1597);
and U1610 (N_1610,N_1503,N_1589);
and U1611 (N_1611,N_1563,N_1599);
or U1612 (N_1612,N_1594,N_1569);
nor U1613 (N_1613,N_1516,N_1565);
or U1614 (N_1614,N_1532,N_1526);
xnor U1615 (N_1615,N_1544,N_1556);
xor U1616 (N_1616,N_1596,N_1540);
and U1617 (N_1617,N_1518,N_1543);
and U1618 (N_1618,N_1595,N_1575);
xnor U1619 (N_1619,N_1551,N_1531);
nand U1620 (N_1620,N_1557,N_1501);
or U1621 (N_1621,N_1513,N_1564);
and U1622 (N_1622,N_1542,N_1510);
nor U1623 (N_1623,N_1517,N_1511);
nand U1624 (N_1624,N_1582,N_1515);
xor U1625 (N_1625,N_1533,N_1568);
nor U1626 (N_1626,N_1548,N_1567);
nor U1627 (N_1627,N_1554,N_1528);
and U1628 (N_1628,N_1547,N_1521);
nor U1629 (N_1629,N_1500,N_1539);
nand U1630 (N_1630,N_1580,N_1566);
or U1631 (N_1631,N_1504,N_1581);
xnor U1632 (N_1632,N_1593,N_1530);
xor U1633 (N_1633,N_1576,N_1527);
xnor U1634 (N_1634,N_1578,N_1520);
or U1635 (N_1635,N_1514,N_1570);
xor U1636 (N_1636,N_1560,N_1558);
and U1637 (N_1637,N_1590,N_1591);
nand U1638 (N_1638,N_1534,N_1505);
nor U1639 (N_1639,N_1559,N_1592);
or U1640 (N_1640,N_1555,N_1562);
nor U1641 (N_1641,N_1508,N_1571);
or U1642 (N_1642,N_1587,N_1523);
nor U1643 (N_1643,N_1522,N_1561);
nor U1644 (N_1644,N_1525,N_1546);
xnor U1645 (N_1645,N_1552,N_1598);
nand U1646 (N_1646,N_1509,N_1584);
or U1647 (N_1647,N_1579,N_1502);
and U1648 (N_1648,N_1538,N_1512);
xnor U1649 (N_1649,N_1529,N_1586);
xnor U1650 (N_1650,N_1530,N_1522);
nand U1651 (N_1651,N_1566,N_1563);
or U1652 (N_1652,N_1515,N_1500);
nor U1653 (N_1653,N_1532,N_1590);
and U1654 (N_1654,N_1557,N_1555);
nor U1655 (N_1655,N_1536,N_1508);
and U1656 (N_1656,N_1549,N_1588);
xor U1657 (N_1657,N_1594,N_1531);
and U1658 (N_1658,N_1511,N_1530);
nand U1659 (N_1659,N_1506,N_1550);
and U1660 (N_1660,N_1573,N_1588);
or U1661 (N_1661,N_1577,N_1501);
nor U1662 (N_1662,N_1527,N_1583);
or U1663 (N_1663,N_1574,N_1523);
nand U1664 (N_1664,N_1573,N_1569);
xor U1665 (N_1665,N_1569,N_1512);
or U1666 (N_1666,N_1539,N_1519);
nor U1667 (N_1667,N_1569,N_1548);
nor U1668 (N_1668,N_1595,N_1510);
or U1669 (N_1669,N_1561,N_1567);
or U1670 (N_1670,N_1557,N_1548);
or U1671 (N_1671,N_1521,N_1527);
xnor U1672 (N_1672,N_1537,N_1568);
or U1673 (N_1673,N_1581,N_1584);
nand U1674 (N_1674,N_1539,N_1550);
nand U1675 (N_1675,N_1541,N_1552);
nand U1676 (N_1676,N_1536,N_1547);
nor U1677 (N_1677,N_1539,N_1562);
xnor U1678 (N_1678,N_1541,N_1578);
xor U1679 (N_1679,N_1527,N_1593);
nand U1680 (N_1680,N_1576,N_1583);
nor U1681 (N_1681,N_1511,N_1519);
nand U1682 (N_1682,N_1535,N_1512);
xnor U1683 (N_1683,N_1564,N_1546);
nand U1684 (N_1684,N_1590,N_1537);
and U1685 (N_1685,N_1531,N_1565);
xnor U1686 (N_1686,N_1507,N_1548);
xnor U1687 (N_1687,N_1535,N_1504);
nor U1688 (N_1688,N_1576,N_1596);
nand U1689 (N_1689,N_1520,N_1580);
xnor U1690 (N_1690,N_1548,N_1584);
or U1691 (N_1691,N_1503,N_1521);
xnor U1692 (N_1692,N_1575,N_1535);
nand U1693 (N_1693,N_1595,N_1584);
xor U1694 (N_1694,N_1544,N_1549);
or U1695 (N_1695,N_1506,N_1599);
or U1696 (N_1696,N_1516,N_1501);
or U1697 (N_1697,N_1523,N_1508);
xnor U1698 (N_1698,N_1585,N_1573);
xor U1699 (N_1699,N_1591,N_1536);
xnor U1700 (N_1700,N_1662,N_1652);
nor U1701 (N_1701,N_1602,N_1689);
nand U1702 (N_1702,N_1663,N_1621);
xor U1703 (N_1703,N_1645,N_1684);
nor U1704 (N_1704,N_1661,N_1695);
or U1705 (N_1705,N_1677,N_1649);
nand U1706 (N_1706,N_1686,N_1647);
or U1707 (N_1707,N_1631,N_1609);
xnor U1708 (N_1708,N_1690,N_1629);
nor U1709 (N_1709,N_1667,N_1638);
or U1710 (N_1710,N_1697,N_1613);
nand U1711 (N_1711,N_1611,N_1651);
nand U1712 (N_1712,N_1660,N_1632);
or U1713 (N_1713,N_1693,N_1620);
or U1714 (N_1714,N_1687,N_1622);
xnor U1715 (N_1715,N_1625,N_1671);
and U1716 (N_1716,N_1600,N_1666);
or U1717 (N_1717,N_1616,N_1615);
xor U1718 (N_1718,N_1627,N_1624);
nand U1719 (N_1719,N_1678,N_1655);
nand U1720 (N_1720,N_1640,N_1635);
and U1721 (N_1721,N_1641,N_1636);
and U1722 (N_1722,N_1656,N_1634);
nand U1723 (N_1723,N_1623,N_1619);
or U1724 (N_1724,N_1601,N_1683);
xnor U1725 (N_1725,N_1679,N_1654);
or U1726 (N_1726,N_1673,N_1642);
nand U1727 (N_1727,N_1676,N_1646);
or U1728 (N_1728,N_1669,N_1608);
nand U1729 (N_1729,N_1657,N_1696);
nor U1730 (N_1730,N_1603,N_1650);
and U1731 (N_1731,N_1688,N_1670);
and U1732 (N_1732,N_1659,N_1604);
or U1733 (N_1733,N_1692,N_1644);
or U1734 (N_1734,N_1643,N_1610);
or U1735 (N_1735,N_1614,N_1653);
and U1736 (N_1736,N_1628,N_1675);
or U1737 (N_1737,N_1607,N_1658);
nor U1738 (N_1738,N_1698,N_1699);
xor U1739 (N_1739,N_1606,N_1633);
and U1740 (N_1740,N_1630,N_1626);
xor U1741 (N_1741,N_1694,N_1681);
and U1742 (N_1742,N_1637,N_1664);
xor U1743 (N_1743,N_1682,N_1691);
xnor U1744 (N_1744,N_1612,N_1639);
xor U1745 (N_1745,N_1674,N_1617);
or U1746 (N_1746,N_1648,N_1668);
nor U1747 (N_1747,N_1680,N_1618);
nand U1748 (N_1748,N_1685,N_1672);
nor U1749 (N_1749,N_1605,N_1665);
or U1750 (N_1750,N_1680,N_1624);
nand U1751 (N_1751,N_1643,N_1605);
nor U1752 (N_1752,N_1618,N_1613);
and U1753 (N_1753,N_1667,N_1684);
nand U1754 (N_1754,N_1678,N_1683);
and U1755 (N_1755,N_1690,N_1674);
xnor U1756 (N_1756,N_1691,N_1609);
and U1757 (N_1757,N_1622,N_1658);
and U1758 (N_1758,N_1632,N_1620);
nand U1759 (N_1759,N_1609,N_1626);
nand U1760 (N_1760,N_1697,N_1661);
xor U1761 (N_1761,N_1699,N_1694);
xnor U1762 (N_1762,N_1683,N_1616);
and U1763 (N_1763,N_1684,N_1634);
nor U1764 (N_1764,N_1605,N_1613);
xor U1765 (N_1765,N_1649,N_1694);
or U1766 (N_1766,N_1639,N_1620);
nand U1767 (N_1767,N_1611,N_1660);
nand U1768 (N_1768,N_1614,N_1678);
or U1769 (N_1769,N_1690,N_1661);
xnor U1770 (N_1770,N_1659,N_1650);
xor U1771 (N_1771,N_1693,N_1638);
nand U1772 (N_1772,N_1627,N_1635);
xor U1773 (N_1773,N_1613,N_1617);
or U1774 (N_1774,N_1605,N_1641);
or U1775 (N_1775,N_1618,N_1693);
xor U1776 (N_1776,N_1671,N_1677);
or U1777 (N_1777,N_1631,N_1688);
nand U1778 (N_1778,N_1695,N_1666);
xnor U1779 (N_1779,N_1630,N_1658);
nand U1780 (N_1780,N_1669,N_1678);
nor U1781 (N_1781,N_1664,N_1608);
nor U1782 (N_1782,N_1641,N_1673);
nand U1783 (N_1783,N_1612,N_1690);
or U1784 (N_1784,N_1622,N_1610);
xnor U1785 (N_1785,N_1698,N_1689);
xnor U1786 (N_1786,N_1627,N_1665);
or U1787 (N_1787,N_1671,N_1634);
xor U1788 (N_1788,N_1618,N_1600);
xor U1789 (N_1789,N_1678,N_1673);
xor U1790 (N_1790,N_1689,N_1613);
nor U1791 (N_1791,N_1691,N_1639);
or U1792 (N_1792,N_1631,N_1673);
nand U1793 (N_1793,N_1646,N_1626);
or U1794 (N_1794,N_1638,N_1680);
nand U1795 (N_1795,N_1677,N_1667);
or U1796 (N_1796,N_1675,N_1605);
nor U1797 (N_1797,N_1685,N_1636);
nor U1798 (N_1798,N_1658,N_1678);
and U1799 (N_1799,N_1695,N_1635);
xor U1800 (N_1800,N_1737,N_1766);
nand U1801 (N_1801,N_1716,N_1752);
and U1802 (N_1802,N_1795,N_1732);
nand U1803 (N_1803,N_1725,N_1748);
xnor U1804 (N_1804,N_1793,N_1720);
or U1805 (N_1805,N_1742,N_1726);
nor U1806 (N_1806,N_1745,N_1723);
xor U1807 (N_1807,N_1746,N_1731);
nand U1808 (N_1808,N_1779,N_1713);
or U1809 (N_1809,N_1744,N_1717);
nor U1810 (N_1810,N_1734,N_1727);
or U1811 (N_1811,N_1751,N_1777);
xnor U1812 (N_1812,N_1741,N_1715);
nand U1813 (N_1813,N_1733,N_1761);
xor U1814 (N_1814,N_1778,N_1788);
xnor U1815 (N_1815,N_1722,N_1755);
xnor U1816 (N_1816,N_1771,N_1789);
xor U1817 (N_1817,N_1798,N_1711);
nor U1818 (N_1818,N_1762,N_1758);
or U1819 (N_1819,N_1792,N_1739);
nand U1820 (N_1820,N_1709,N_1756);
and U1821 (N_1821,N_1708,N_1760);
xnor U1822 (N_1822,N_1787,N_1712);
nor U1823 (N_1823,N_1710,N_1776);
nor U1824 (N_1824,N_1718,N_1774);
xor U1825 (N_1825,N_1714,N_1705);
xnor U1826 (N_1826,N_1747,N_1700);
or U1827 (N_1827,N_1753,N_1785);
and U1828 (N_1828,N_1706,N_1796);
and U1829 (N_1829,N_1768,N_1724);
nor U1830 (N_1830,N_1786,N_1719);
nand U1831 (N_1831,N_1772,N_1765);
nand U1832 (N_1832,N_1740,N_1729);
nor U1833 (N_1833,N_1728,N_1704);
nor U1834 (N_1834,N_1750,N_1783);
nor U1835 (N_1835,N_1780,N_1738);
nand U1836 (N_1836,N_1736,N_1707);
nand U1837 (N_1837,N_1701,N_1770);
and U1838 (N_1838,N_1757,N_1773);
or U1839 (N_1839,N_1784,N_1799);
nor U1840 (N_1840,N_1703,N_1759);
nand U1841 (N_1841,N_1797,N_1730);
and U1842 (N_1842,N_1702,N_1791);
nand U1843 (N_1843,N_1754,N_1735);
and U1844 (N_1844,N_1790,N_1763);
and U1845 (N_1845,N_1764,N_1794);
and U1846 (N_1846,N_1743,N_1749);
nand U1847 (N_1847,N_1721,N_1781);
xnor U1848 (N_1848,N_1775,N_1767);
nand U1849 (N_1849,N_1769,N_1782);
xor U1850 (N_1850,N_1700,N_1778);
and U1851 (N_1851,N_1791,N_1705);
or U1852 (N_1852,N_1779,N_1735);
nand U1853 (N_1853,N_1760,N_1705);
nand U1854 (N_1854,N_1737,N_1713);
xnor U1855 (N_1855,N_1757,N_1720);
xor U1856 (N_1856,N_1771,N_1784);
nor U1857 (N_1857,N_1759,N_1719);
and U1858 (N_1858,N_1726,N_1781);
or U1859 (N_1859,N_1783,N_1776);
or U1860 (N_1860,N_1753,N_1774);
xor U1861 (N_1861,N_1765,N_1759);
nand U1862 (N_1862,N_1702,N_1769);
nand U1863 (N_1863,N_1747,N_1722);
xnor U1864 (N_1864,N_1701,N_1763);
or U1865 (N_1865,N_1782,N_1713);
xor U1866 (N_1866,N_1748,N_1744);
and U1867 (N_1867,N_1788,N_1720);
and U1868 (N_1868,N_1744,N_1768);
nand U1869 (N_1869,N_1795,N_1769);
nor U1870 (N_1870,N_1712,N_1714);
nor U1871 (N_1871,N_1705,N_1718);
xnor U1872 (N_1872,N_1749,N_1728);
nor U1873 (N_1873,N_1723,N_1754);
nor U1874 (N_1874,N_1742,N_1769);
and U1875 (N_1875,N_1796,N_1768);
xor U1876 (N_1876,N_1726,N_1784);
and U1877 (N_1877,N_1737,N_1727);
or U1878 (N_1878,N_1753,N_1795);
nand U1879 (N_1879,N_1710,N_1701);
nand U1880 (N_1880,N_1726,N_1755);
and U1881 (N_1881,N_1798,N_1737);
nand U1882 (N_1882,N_1790,N_1717);
xnor U1883 (N_1883,N_1707,N_1753);
nor U1884 (N_1884,N_1712,N_1778);
nand U1885 (N_1885,N_1757,N_1791);
or U1886 (N_1886,N_1792,N_1756);
nor U1887 (N_1887,N_1738,N_1721);
and U1888 (N_1888,N_1782,N_1795);
and U1889 (N_1889,N_1700,N_1723);
or U1890 (N_1890,N_1787,N_1761);
nand U1891 (N_1891,N_1794,N_1717);
nand U1892 (N_1892,N_1777,N_1721);
or U1893 (N_1893,N_1750,N_1728);
and U1894 (N_1894,N_1773,N_1725);
nand U1895 (N_1895,N_1775,N_1764);
or U1896 (N_1896,N_1769,N_1746);
nor U1897 (N_1897,N_1770,N_1788);
nor U1898 (N_1898,N_1705,N_1752);
xor U1899 (N_1899,N_1729,N_1743);
and U1900 (N_1900,N_1851,N_1876);
nand U1901 (N_1901,N_1867,N_1833);
nand U1902 (N_1902,N_1828,N_1891);
or U1903 (N_1903,N_1842,N_1852);
nand U1904 (N_1904,N_1880,N_1834);
or U1905 (N_1905,N_1874,N_1870);
or U1906 (N_1906,N_1894,N_1873);
nand U1907 (N_1907,N_1872,N_1865);
nor U1908 (N_1908,N_1885,N_1810);
nor U1909 (N_1909,N_1840,N_1848);
nand U1910 (N_1910,N_1893,N_1802);
xor U1911 (N_1911,N_1814,N_1889);
xnor U1912 (N_1912,N_1849,N_1825);
or U1913 (N_1913,N_1822,N_1839);
or U1914 (N_1914,N_1801,N_1883);
nor U1915 (N_1915,N_1890,N_1815);
nand U1916 (N_1916,N_1807,N_1850);
nor U1917 (N_1917,N_1831,N_1812);
xnor U1918 (N_1918,N_1869,N_1843);
nor U1919 (N_1919,N_1844,N_1845);
xor U1920 (N_1920,N_1832,N_1868);
nor U1921 (N_1921,N_1847,N_1892);
xnor U1922 (N_1922,N_1817,N_1820);
and U1923 (N_1923,N_1838,N_1823);
or U1924 (N_1924,N_1836,N_1835);
or U1925 (N_1925,N_1856,N_1855);
or U1926 (N_1926,N_1857,N_1871);
nand U1927 (N_1927,N_1830,N_1808);
xnor U1928 (N_1928,N_1861,N_1862);
or U1929 (N_1929,N_1837,N_1829);
and U1930 (N_1930,N_1811,N_1897);
nor U1931 (N_1931,N_1821,N_1858);
nor U1932 (N_1932,N_1818,N_1886);
nor U1933 (N_1933,N_1884,N_1896);
nor U1934 (N_1934,N_1863,N_1898);
nor U1935 (N_1935,N_1859,N_1887);
nand U1936 (N_1936,N_1816,N_1866);
and U1937 (N_1937,N_1875,N_1809);
nor U1938 (N_1938,N_1882,N_1878);
or U1939 (N_1939,N_1895,N_1819);
nor U1940 (N_1940,N_1888,N_1877);
or U1941 (N_1941,N_1803,N_1879);
and U1942 (N_1942,N_1813,N_1826);
and U1943 (N_1943,N_1899,N_1800);
and U1944 (N_1944,N_1860,N_1846);
xor U1945 (N_1945,N_1881,N_1864);
and U1946 (N_1946,N_1806,N_1805);
or U1947 (N_1947,N_1854,N_1853);
nand U1948 (N_1948,N_1841,N_1804);
xnor U1949 (N_1949,N_1827,N_1824);
xnor U1950 (N_1950,N_1842,N_1889);
and U1951 (N_1951,N_1889,N_1836);
nand U1952 (N_1952,N_1898,N_1842);
or U1953 (N_1953,N_1889,N_1885);
or U1954 (N_1954,N_1802,N_1872);
xnor U1955 (N_1955,N_1816,N_1811);
nor U1956 (N_1956,N_1878,N_1822);
nor U1957 (N_1957,N_1814,N_1826);
or U1958 (N_1958,N_1823,N_1867);
and U1959 (N_1959,N_1862,N_1886);
and U1960 (N_1960,N_1850,N_1883);
and U1961 (N_1961,N_1857,N_1881);
or U1962 (N_1962,N_1893,N_1890);
and U1963 (N_1963,N_1897,N_1880);
xor U1964 (N_1964,N_1819,N_1808);
and U1965 (N_1965,N_1842,N_1872);
and U1966 (N_1966,N_1809,N_1805);
xnor U1967 (N_1967,N_1852,N_1832);
nor U1968 (N_1968,N_1846,N_1840);
nor U1969 (N_1969,N_1804,N_1818);
or U1970 (N_1970,N_1853,N_1827);
xor U1971 (N_1971,N_1806,N_1847);
nand U1972 (N_1972,N_1832,N_1877);
nand U1973 (N_1973,N_1884,N_1801);
or U1974 (N_1974,N_1839,N_1898);
or U1975 (N_1975,N_1897,N_1809);
xor U1976 (N_1976,N_1882,N_1858);
or U1977 (N_1977,N_1895,N_1808);
and U1978 (N_1978,N_1828,N_1823);
nand U1979 (N_1979,N_1855,N_1876);
nor U1980 (N_1980,N_1827,N_1829);
or U1981 (N_1981,N_1853,N_1828);
or U1982 (N_1982,N_1875,N_1814);
nand U1983 (N_1983,N_1858,N_1804);
and U1984 (N_1984,N_1866,N_1850);
xor U1985 (N_1985,N_1803,N_1849);
nor U1986 (N_1986,N_1802,N_1822);
and U1987 (N_1987,N_1871,N_1867);
nor U1988 (N_1988,N_1837,N_1854);
xnor U1989 (N_1989,N_1875,N_1882);
and U1990 (N_1990,N_1832,N_1869);
xnor U1991 (N_1991,N_1891,N_1802);
xor U1992 (N_1992,N_1820,N_1896);
and U1993 (N_1993,N_1894,N_1899);
or U1994 (N_1994,N_1819,N_1811);
xnor U1995 (N_1995,N_1855,N_1819);
nor U1996 (N_1996,N_1892,N_1886);
or U1997 (N_1997,N_1807,N_1875);
nor U1998 (N_1998,N_1888,N_1831);
or U1999 (N_1999,N_1811,N_1857);
and U2000 (N_2000,N_1972,N_1927);
or U2001 (N_2001,N_1999,N_1944);
nand U2002 (N_2002,N_1901,N_1984);
xor U2003 (N_2003,N_1953,N_1923);
nand U2004 (N_2004,N_1946,N_1977);
xnor U2005 (N_2005,N_1959,N_1920);
xor U2006 (N_2006,N_1940,N_1907);
nand U2007 (N_2007,N_1912,N_1910);
and U2008 (N_2008,N_1939,N_1934);
xor U2009 (N_2009,N_1950,N_1998);
xor U2010 (N_2010,N_1981,N_1976);
and U2011 (N_2011,N_1992,N_1971);
nand U2012 (N_2012,N_1989,N_1955);
xnor U2013 (N_2013,N_1904,N_1969);
or U2014 (N_2014,N_1974,N_1986);
nand U2015 (N_2015,N_1970,N_1937);
xnor U2016 (N_2016,N_1900,N_1963);
and U2017 (N_2017,N_1949,N_1947);
and U2018 (N_2018,N_1915,N_1983);
or U2019 (N_2019,N_1991,N_1964);
xnor U2020 (N_2020,N_1960,N_1911);
nand U2021 (N_2021,N_1996,N_1997);
nor U2022 (N_2022,N_1906,N_1935);
or U2023 (N_2023,N_1936,N_1929);
xnor U2024 (N_2024,N_1908,N_1903);
and U2025 (N_2025,N_1979,N_1925);
and U2026 (N_2026,N_1952,N_1932);
nand U2027 (N_2027,N_1928,N_1961);
nand U2028 (N_2028,N_1913,N_1978);
nor U2029 (N_2029,N_1993,N_1951);
xor U2030 (N_2030,N_1941,N_1994);
nor U2031 (N_2031,N_1987,N_1985);
xor U2032 (N_2032,N_1918,N_1966);
and U2033 (N_2033,N_1921,N_1965);
or U2034 (N_2034,N_1942,N_1967);
xor U2035 (N_2035,N_1917,N_1902);
and U2036 (N_2036,N_1943,N_1914);
nor U2037 (N_2037,N_1995,N_1922);
nor U2038 (N_2038,N_1973,N_1990);
nor U2039 (N_2039,N_1938,N_1909);
and U2040 (N_2040,N_1982,N_1926);
nor U2041 (N_2041,N_1916,N_1931);
nor U2042 (N_2042,N_1919,N_1924);
nor U2043 (N_2043,N_1948,N_1975);
nor U2044 (N_2044,N_1905,N_1945);
or U2045 (N_2045,N_1968,N_1957);
xnor U2046 (N_2046,N_1988,N_1933);
nor U2047 (N_2047,N_1980,N_1954);
nand U2048 (N_2048,N_1930,N_1962);
nor U2049 (N_2049,N_1956,N_1958);
or U2050 (N_2050,N_1986,N_1920);
nand U2051 (N_2051,N_1996,N_1922);
and U2052 (N_2052,N_1969,N_1997);
xnor U2053 (N_2053,N_1989,N_1923);
nor U2054 (N_2054,N_1924,N_1973);
nor U2055 (N_2055,N_1999,N_1988);
xnor U2056 (N_2056,N_1997,N_1909);
nor U2057 (N_2057,N_1942,N_1982);
and U2058 (N_2058,N_1935,N_1953);
or U2059 (N_2059,N_1999,N_1928);
nor U2060 (N_2060,N_1913,N_1908);
or U2061 (N_2061,N_1970,N_1944);
nand U2062 (N_2062,N_1988,N_1920);
xnor U2063 (N_2063,N_1954,N_1915);
xnor U2064 (N_2064,N_1930,N_1937);
or U2065 (N_2065,N_1969,N_1922);
and U2066 (N_2066,N_1976,N_1905);
nand U2067 (N_2067,N_1958,N_1955);
and U2068 (N_2068,N_1984,N_1990);
nor U2069 (N_2069,N_1995,N_1943);
or U2070 (N_2070,N_1917,N_1963);
xor U2071 (N_2071,N_1915,N_1957);
xnor U2072 (N_2072,N_1922,N_1982);
xnor U2073 (N_2073,N_1905,N_1954);
and U2074 (N_2074,N_1987,N_1976);
and U2075 (N_2075,N_1962,N_1972);
nand U2076 (N_2076,N_1965,N_1913);
nand U2077 (N_2077,N_1951,N_1962);
nor U2078 (N_2078,N_1930,N_1919);
nand U2079 (N_2079,N_1904,N_1914);
nand U2080 (N_2080,N_1996,N_1974);
and U2081 (N_2081,N_1935,N_1905);
xnor U2082 (N_2082,N_1981,N_1966);
nand U2083 (N_2083,N_1915,N_1988);
nand U2084 (N_2084,N_1995,N_1917);
or U2085 (N_2085,N_1923,N_1901);
xor U2086 (N_2086,N_1935,N_1925);
nor U2087 (N_2087,N_1995,N_1902);
and U2088 (N_2088,N_1966,N_1999);
nand U2089 (N_2089,N_1923,N_1977);
xor U2090 (N_2090,N_1939,N_1963);
and U2091 (N_2091,N_1990,N_1902);
and U2092 (N_2092,N_1938,N_1929);
and U2093 (N_2093,N_1954,N_1940);
xnor U2094 (N_2094,N_1959,N_1921);
xnor U2095 (N_2095,N_1934,N_1953);
and U2096 (N_2096,N_1969,N_1987);
nand U2097 (N_2097,N_1934,N_1984);
or U2098 (N_2098,N_1997,N_1919);
or U2099 (N_2099,N_1976,N_1925);
nor U2100 (N_2100,N_2005,N_2036);
or U2101 (N_2101,N_2014,N_2009);
nor U2102 (N_2102,N_2068,N_2074);
nor U2103 (N_2103,N_2093,N_2010);
nor U2104 (N_2104,N_2052,N_2043);
and U2105 (N_2105,N_2067,N_2091);
or U2106 (N_2106,N_2011,N_2024);
nor U2107 (N_2107,N_2085,N_2095);
nor U2108 (N_2108,N_2000,N_2094);
nor U2109 (N_2109,N_2057,N_2061);
and U2110 (N_2110,N_2071,N_2049);
nand U2111 (N_2111,N_2042,N_2055);
nand U2112 (N_2112,N_2064,N_2039);
and U2113 (N_2113,N_2044,N_2023);
nand U2114 (N_2114,N_2046,N_2001);
nor U2115 (N_2115,N_2027,N_2082);
nor U2116 (N_2116,N_2021,N_2086);
or U2117 (N_2117,N_2004,N_2054);
xnor U2118 (N_2118,N_2087,N_2077);
nor U2119 (N_2119,N_2020,N_2066);
nor U2120 (N_2120,N_2013,N_2070);
and U2121 (N_2121,N_2029,N_2099);
nor U2122 (N_2122,N_2003,N_2075);
or U2123 (N_2123,N_2048,N_2096);
or U2124 (N_2124,N_2006,N_2076);
or U2125 (N_2125,N_2050,N_2035);
and U2126 (N_2126,N_2079,N_2022);
nor U2127 (N_2127,N_2007,N_2034);
and U2128 (N_2128,N_2089,N_2090);
xnor U2129 (N_2129,N_2078,N_2062);
nand U2130 (N_2130,N_2080,N_2092);
nand U2131 (N_2131,N_2047,N_2059);
nor U2132 (N_2132,N_2069,N_2038);
xnor U2133 (N_2133,N_2041,N_2083);
nor U2134 (N_2134,N_2002,N_2051);
xnor U2135 (N_2135,N_2084,N_2097);
or U2136 (N_2136,N_2065,N_2030);
xnor U2137 (N_2137,N_2028,N_2081);
or U2138 (N_2138,N_2032,N_2025);
nand U2139 (N_2139,N_2063,N_2015);
xnor U2140 (N_2140,N_2045,N_2026);
nor U2141 (N_2141,N_2016,N_2040);
or U2142 (N_2142,N_2012,N_2033);
nor U2143 (N_2143,N_2088,N_2058);
or U2144 (N_2144,N_2018,N_2017);
and U2145 (N_2145,N_2056,N_2019);
and U2146 (N_2146,N_2098,N_2073);
xor U2147 (N_2147,N_2031,N_2008);
or U2148 (N_2148,N_2072,N_2053);
nand U2149 (N_2149,N_2037,N_2060);
xor U2150 (N_2150,N_2095,N_2071);
xor U2151 (N_2151,N_2001,N_2095);
nor U2152 (N_2152,N_2001,N_2035);
xnor U2153 (N_2153,N_2065,N_2050);
and U2154 (N_2154,N_2087,N_2071);
nor U2155 (N_2155,N_2018,N_2080);
nand U2156 (N_2156,N_2025,N_2096);
nand U2157 (N_2157,N_2024,N_2073);
or U2158 (N_2158,N_2034,N_2011);
xnor U2159 (N_2159,N_2021,N_2020);
nor U2160 (N_2160,N_2064,N_2012);
or U2161 (N_2161,N_2043,N_2020);
nand U2162 (N_2162,N_2024,N_2033);
xnor U2163 (N_2163,N_2086,N_2080);
and U2164 (N_2164,N_2078,N_2020);
xor U2165 (N_2165,N_2026,N_2076);
or U2166 (N_2166,N_2083,N_2029);
nand U2167 (N_2167,N_2006,N_2088);
or U2168 (N_2168,N_2059,N_2069);
and U2169 (N_2169,N_2074,N_2020);
nor U2170 (N_2170,N_2054,N_2096);
nor U2171 (N_2171,N_2050,N_2014);
nand U2172 (N_2172,N_2041,N_2029);
and U2173 (N_2173,N_2005,N_2015);
or U2174 (N_2174,N_2045,N_2016);
nor U2175 (N_2175,N_2021,N_2064);
nor U2176 (N_2176,N_2084,N_2018);
and U2177 (N_2177,N_2024,N_2066);
nor U2178 (N_2178,N_2001,N_2030);
nor U2179 (N_2179,N_2098,N_2090);
xnor U2180 (N_2180,N_2065,N_2002);
or U2181 (N_2181,N_2086,N_2037);
nand U2182 (N_2182,N_2081,N_2045);
or U2183 (N_2183,N_2075,N_2021);
nand U2184 (N_2184,N_2032,N_2066);
nor U2185 (N_2185,N_2071,N_2027);
nor U2186 (N_2186,N_2071,N_2004);
and U2187 (N_2187,N_2004,N_2096);
or U2188 (N_2188,N_2071,N_2009);
nor U2189 (N_2189,N_2044,N_2087);
and U2190 (N_2190,N_2020,N_2053);
xnor U2191 (N_2191,N_2058,N_2036);
and U2192 (N_2192,N_2045,N_2097);
and U2193 (N_2193,N_2072,N_2028);
nand U2194 (N_2194,N_2092,N_2025);
or U2195 (N_2195,N_2027,N_2010);
nand U2196 (N_2196,N_2036,N_2061);
xor U2197 (N_2197,N_2084,N_2023);
nor U2198 (N_2198,N_2064,N_2016);
or U2199 (N_2199,N_2084,N_2061);
xnor U2200 (N_2200,N_2182,N_2190);
nor U2201 (N_2201,N_2104,N_2108);
nor U2202 (N_2202,N_2166,N_2118);
or U2203 (N_2203,N_2106,N_2150);
nand U2204 (N_2204,N_2147,N_2122);
xnor U2205 (N_2205,N_2110,N_2185);
or U2206 (N_2206,N_2169,N_2162);
or U2207 (N_2207,N_2136,N_2157);
nor U2208 (N_2208,N_2111,N_2123);
and U2209 (N_2209,N_2139,N_2193);
nor U2210 (N_2210,N_2102,N_2181);
xnor U2211 (N_2211,N_2128,N_2120);
and U2212 (N_2212,N_2180,N_2187);
and U2213 (N_2213,N_2160,N_2119);
xor U2214 (N_2214,N_2153,N_2134);
nor U2215 (N_2215,N_2112,N_2141);
and U2216 (N_2216,N_2144,N_2196);
and U2217 (N_2217,N_2191,N_2197);
and U2218 (N_2218,N_2161,N_2199);
xnor U2219 (N_2219,N_2121,N_2163);
nand U2220 (N_2220,N_2177,N_2156);
xor U2221 (N_2221,N_2189,N_2132);
nand U2222 (N_2222,N_2101,N_2149);
and U2223 (N_2223,N_2135,N_2148);
xor U2224 (N_2224,N_2142,N_2194);
or U2225 (N_2225,N_2126,N_2103);
nand U2226 (N_2226,N_2145,N_2164);
nor U2227 (N_2227,N_2179,N_2170);
xor U2228 (N_2228,N_2155,N_2188);
nand U2229 (N_2229,N_2192,N_2146);
nor U2230 (N_2230,N_2127,N_2198);
or U2231 (N_2231,N_2174,N_2114);
nand U2232 (N_2232,N_2168,N_2117);
or U2233 (N_2233,N_2172,N_2159);
or U2234 (N_2234,N_2171,N_2115);
nor U2235 (N_2235,N_2131,N_2154);
xnor U2236 (N_2236,N_2184,N_2100);
and U2237 (N_2237,N_2137,N_2105);
or U2238 (N_2238,N_2167,N_2175);
or U2239 (N_2239,N_2158,N_2183);
nor U2240 (N_2240,N_2165,N_2113);
xnor U2241 (N_2241,N_2176,N_2138);
and U2242 (N_2242,N_2173,N_2143);
and U2243 (N_2243,N_2116,N_2133);
or U2244 (N_2244,N_2109,N_2124);
nand U2245 (N_2245,N_2130,N_2186);
nand U2246 (N_2246,N_2178,N_2140);
xnor U2247 (N_2247,N_2152,N_2125);
xor U2248 (N_2248,N_2151,N_2195);
xor U2249 (N_2249,N_2129,N_2107);
nor U2250 (N_2250,N_2120,N_2175);
and U2251 (N_2251,N_2100,N_2153);
xor U2252 (N_2252,N_2179,N_2122);
or U2253 (N_2253,N_2121,N_2151);
or U2254 (N_2254,N_2157,N_2138);
nand U2255 (N_2255,N_2138,N_2160);
xor U2256 (N_2256,N_2163,N_2158);
nand U2257 (N_2257,N_2192,N_2134);
nor U2258 (N_2258,N_2189,N_2196);
nand U2259 (N_2259,N_2152,N_2186);
nand U2260 (N_2260,N_2184,N_2153);
xnor U2261 (N_2261,N_2140,N_2142);
xor U2262 (N_2262,N_2170,N_2108);
nand U2263 (N_2263,N_2114,N_2178);
and U2264 (N_2264,N_2131,N_2122);
or U2265 (N_2265,N_2183,N_2117);
or U2266 (N_2266,N_2131,N_2137);
xor U2267 (N_2267,N_2177,N_2119);
xor U2268 (N_2268,N_2160,N_2146);
nor U2269 (N_2269,N_2105,N_2122);
and U2270 (N_2270,N_2163,N_2128);
nor U2271 (N_2271,N_2199,N_2149);
and U2272 (N_2272,N_2192,N_2174);
nand U2273 (N_2273,N_2169,N_2171);
and U2274 (N_2274,N_2192,N_2196);
and U2275 (N_2275,N_2120,N_2154);
nand U2276 (N_2276,N_2128,N_2114);
nor U2277 (N_2277,N_2111,N_2154);
nor U2278 (N_2278,N_2102,N_2198);
nand U2279 (N_2279,N_2169,N_2109);
or U2280 (N_2280,N_2127,N_2126);
xnor U2281 (N_2281,N_2190,N_2166);
nor U2282 (N_2282,N_2172,N_2175);
nand U2283 (N_2283,N_2143,N_2144);
xor U2284 (N_2284,N_2184,N_2165);
xor U2285 (N_2285,N_2110,N_2189);
nor U2286 (N_2286,N_2140,N_2154);
or U2287 (N_2287,N_2190,N_2148);
or U2288 (N_2288,N_2152,N_2173);
nand U2289 (N_2289,N_2170,N_2189);
or U2290 (N_2290,N_2199,N_2113);
or U2291 (N_2291,N_2144,N_2140);
nor U2292 (N_2292,N_2150,N_2183);
nor U2293 (N_2293,N_2113,N_2119);
nor U2294 (N_2294,N_2177,N_2187);
nor U2295 (N_2295,N_2178,N_2193);
and U2296 (N_2296,N_2149,N_2174);
nand U2297 (N_2297,N_2134,N_2142);
xnor U2298 (N_2298,N_2175,N_2118);
or U2299 (N_2299,N_2100,N_2142);
xnor U2300 (N_2300,N_2265,N_2200);
xor U2301 (N_2301,N_2239,N_2202);
nand U2302 (N_2302,N_2284,N_2291);
or U2303 (N_2303,N_2251,N_2249);
nand U2304 (N_2304,N_2296,N_2221);
or U2305 (N_2305,N_2277,N_2215);
nor U2306 (N_2306,N_2290,N_2297);
and U2307 (N_2307,N_2209,N_2260);
and U2308 (N_2308,N_2216,N_2224);
xor U2309 (N_2309,N_2207,N_2235);
xor U2310 (N_2310,N_2261,N_2263);
and U2311 (N_2311,N_2288,N_2243);
and U2312 (N_2312,N_2268,N_2272);
xor U2313 (N_2313,N_2279,N_2240);
nor U2314 (N_2314,N_2204,N_2231);
or U2315 (N_2315,N_2246,N_2250);
nor U2316 (N_2316,N_2254,N_2273);
or U2317 (N_2317,N_2230,N_2281);
nand U2318 (N_2318,N_2212,N_2282);
xnor U2319 (N_2319,N_2274,N_2294);
and U2320 (N_2320,N_2262,N_2201);
or U2321 (N_2321,N_2269,N_2226);
nor U2322 (N_2322,N_2219,N_2232);
and U2323 (N_2323,N_2255,N_2252);
or U2324 (N_2324,N_2227,N_2213);
xnor U2325 (N_2325,N_2275,N_2259);
nand U2326 (N_2326,N_2285,N_2238);
and U2327 (N_2327,N_2298,N_2217);
nor U2328 (N_2328,N_2244,N_2208);
or U2329 (N_2329,N_2283,N_2205);
xor U2330 (N_2330,N_2237,N_2228);
nor U2331 (N_2331,N_2218,N_2225);
or U2332 (N_2332,N_2248,N_2257);
xor U2333 (N_2333,N_2242,N_2258);
nand U2334 (N_2334,N_2287,N_2223);
nand U2335 (N_2335,N_2233,N_2276);
nand U2336 (N_2336,N_2271,N_2245);
or U2337 (N_2337,N_2203,N_2229);
or U2338 (N_2338,N_2210,N_2214);
and U2339 (N_2339,N_2256,N_2292);
and U2340 (N_2340,N_2280,N_2299);
nand U2341 (N_2341,N_2247,N_2266);
nor U2342 (N_2342,N_2220,N_2206);
and U2343 (N_2343,N_2222,N_2234);
or U2344 (N_2344,N_2270,N_2253);
xor U2345 (N_2345,N_2267,N_2295);
nor U2346 (N_2346,N_2211,N_2289);
nor U2347 (N_2347,N_2264,N_2278);
and U2348 (N_2348,N_2293,N_2286);
xnor U2349 (N_2349,N_2241,N_2236);
and U2350 (N_2350,N_2269,N_2268);
nor U2351 (N_2351,N_2262,N_2230);
nand U2352 (N_2352,N_2254,N_2235);
or U2353 (N_2353,N_2259,N_2244);
nor U2354 (N_2354,N_2206,N_2207);
xor U2355 (N_2355,N_2244,N_2242);
nand U2356 (N_2356,N_2232,N_2234);
or U2357 (N_2357,N_2228,N_2235);
nand U2358 (N_2358,N_2201,N_2213);
nand U2359 (N_2359,N_2203,N_2286);
nand U2360 (N_2360,N_2201,N_2273);
nor U2361 (N_2361,N_2249,N_2246);
xor U2362 (N_2362,N_2292,N_2215);
xnor U2363 (N_2363,N_2271,N_2252);
nand U2364 (N_2364,N_2233,N_2228);
and U2365 (N_2365,N_2287,N_2277);
or U2366 (N_2366,N_2269,N_2248);
nand U2367 (N_2367,N_2209,N_2298);
nand U2368 (N_2368,N_2284,N_2265);
or U2369 (N_2369,N_2240,N_2218);
xnor U2370 (N_2370,N_2203,N_2233);
or U2371 (N_2371,N_2243,N_2250);
nor U2372 (N_2372,N_2285,N_2220);
and U2373 (N_2373,N_2292,N_2233);
nor U2374 (N_2374,N_2262,N_2245);
nand U2375 (N_2375,N_2279,N_2238);
and U2376 (N_2376,N_2256,N_2223);
xor U2377 (N_2377,N_2201,N_2209);
or U2378 (N_2378,N_2239,N_2221);
nor U2379 (N_2379,N_2272,N_2291);
nor U2380 (N_2380,N_2296,N_2202);
or U2381 (N_2381,N_2233,N_2296);
xor U2382 (N_2382,N_2291,N_2220);
and U2383 (N_2383,N_2282,N_2292);
and U2384 (N_2384,N_2222,N_2210);
and U2385 (N_2385,N_2263,N_2236);
nor U2386 (N_2386,N_2250,N_2292);
and U2387 (N_2387,N_2289,N_2272);
nor U2388 (N_2388,N_2294,N_2260);
or U2389 (N_2389,N_2272,N_2294);
xor U2390 (N_2390,N_2212,N_2239);
nand U2391 (N_2391,N_2269,N_2281);
xor U2392 (N_2392,N_2224,N_2271);
nand U2393 (N_2393,N_2271,N_2259);
and U2394 (N_2394,N_2238,N_2269);
nor U2395 (N_2395,N_2207,N_2232);
nand U2396 (N_2396,N_2207,N_2241);
nor U2397 (N_2397,N_2289,N_2277);
nor U2398 (N_2398,N_2275,N_2274);
or U2399 (N_2399,N_2256,N_2251);
nand U2400 (N_2400,N_2327,N_2321);
nand U2401 (N_2401,N_2336,N_2353);
or U2402 (N_2402,N_2347,N_2385);
xnor U2403 (N_2403,N_2349,N_2384);
nand U2404 (N_2404,N_2367,N_2322);
nand U2405 (N_2405,N_2396,N_2343);
nand U2406 (N_2406,N_2360,N_2334);
or U2407 (N_2407,N_2309,N_2373);
nor U2408 (N_2408,N_2365,N_2366);
nor U2409 (N_2409,N_2328,N_2381);
nand U2410 (N_2410,N_2398,N_2318);
nor U2411 (N_2411,N_2325,N_2315);
and U2412 (N_2412,N_2362,N_2342);
nor U2413 (N_2413,N_2320,N_2339);
or U2414 (N_2414,N_2324,N_2391);
nand U2415 (N_2415,N_2394,N_2356);
nor U2416 (N_2416,N_2346,N_2313);
or U2417 (N_2417,N_2345,N_2372);
xnor U2418 (N_2418,N_2369,N_2351);
xnor U2419 (N_2419,N_2364,N_2329);
xnor U2420 (N_2420,N_2333,N_2359);
xor U2421 (N_2421,N_2377,N_2390);
and U2422 (N_2422,N_2340,N_2335);
nand U2423 (N_2423,N_2303,N_2352);
or U2424 (N_2424,N_2399,N_2387);
and U2425 (N_2425,N_2380,N_2341);
nand U2426 (N_2426,N_2310,N_2306);
or U2427 (N_2427,N_2331,N_2314);
nand U2428 (N_2428,N_2363,N_2393);
and U2429 (N_2429,N_2358,N_2307);
xor U2430 (N_2430,N_2301,N_2361);
nand U2431 (N_2431,N_2379,N_2348);
nand U2432 (N_2432,N_2350,N_2326);
nand U2433 (N_2433,N_2316,N_2337);
nor U2434 (N_2434,N_2338,N_2344);
nand U2435 (N_2435,N_2305,N_2370);
and U2436 (N_2436,N_2317,N_2323);
nor U2437 (N_2437,N_2392,N_2332);
and U2438 (N_2438,N_2374,N_2388);
and U2439 (N_2439,N_2354,N_2371);
or U2440 (N_2440,N_2395,N_2375);
and U2441 (N_2441,N_2368,N_2312);
and U2442 (N_2442,N_2355,N_2357);
and U2443 (N_2443,N_2302,N_2382);
or U2444 (N_2444,N_2397,N_2389);
xor U2445 (N_2445,N_2383,N_2304);
xnor U2446 (N_2446,N_2300,N_2319);
or U2447 (N_2447,N_2311,N_2330);
nor U2448 (N_2448,N_2386,N_2308);
xnor U2449 (N_2449,N_2376,N_2378);
or U2450 (N_2450,N_2303,N_2331);
or U2451 (N_2451,N_2353,N_2340);
nand U2452 (N_2452,N_2310,N_2309);
and U2453 (N_2453,N_2390,N_2359);
nand U2454 (N_2454,N_2338,N_2304);
and U2455 (N_2455,N_2330,N_2358);
and U2456 (N_2456,N_2369,N_2368);
and U2457 (N_2457,N_2343,N_2372);
and U2458 (N_2458,N_2362,N_2375);
and U2459 (N_2459,N_2305,N_2361);
or U2460 (N_2460,N_2359,N_2309);
nor U2461 (N_2461,N_2378,N_2315);
xnor U2462 (N_2462,N_2321,N_2389);
or U2463 (N_2463,N_2381,N_2324);
nor U2464 (N_2464,N_2309,N_2323);
or U2465 (N_2465,N_2351,N_2336);
and U2466 (N_2466,N_2337,N_2368);
nand U2467 (N_2467,N_2351,N_2361);
xnor U2468 (N_2468,N_2338,N_2306);
xnor U2469 (N_2469,N_2338,N_2383);
or U2470 (N_2470,N_2390,N_2381);
and U2471 (N_2471,N_2366,N_2341);
xnor U2472 (N_2472,N_2379,N_2326);
xor U2473 (N_2473,N_2379,N_2392);
or U2474 (N_2474,N_2333,N_2304);
and U2475 (N_2475,N_2356,N_2347);
nor U2476 (N_2476,N_2391,N_2381);
and U2477 (N_2477,N_2376,N_2362);
nor U2478 (N_2478,N_2315,N_2350);
nand U2479 (N_2479,N_2359,N_2378);
nor U2480 (N_2480,N_2321,N_2385);
or U2481 (N_2481,N_2349,N_2336);
nand U2482 (N_2482,N_2309,N_2329);
and U2483 (N_2483,N_2357,N_2387);
or U2484 (N_2484,N_2300,N_2368);
xnor U2485 (N_2485,N_2344,N_2378);
or U2486 (N_2486,N_2378,N_2381);
nand U2487 (N_2487,N_2378,N_2358);
xnor U2488 (N_2488,N_2349,N_2311);
nand U2489 (N_2489,N_2310,N_2373);
or U2490 (N_2490,N_2348,N_2382);
xnor U2491 (N_2491,N_2332,N_2361);
xnor U2492 (N_2492,N_2395,N_2374);
nand U2493 (N_2493,N_2349,N_2363);
xnor U2494 (N_2494,N_2366,N_2368);
xor U2495 (N_2495,N_2384,N_2388);
xnor U2496 (N_2496,N_2322,N_2388);
xnor U2497 (N_2497,N_2374,N_2330);
xnor U2498 (N_2498,N_2337,N_2393);
xnor U2499 (N_2499,N_2360,N_2354);
xor U2500 (N_2500,N_2413,N_2466);
nor U2501 (N_2501,N_2486,N_2433);
and U2502 (N_2502,N_2453,N_2409);
and U2503 (N_2503,N_2487,N_2457);
or U2504 (N_2504,N_2482,N_2475);
and U2505 (N_2505,N_2430,N_2480);
nor U2506 (N_2506,N_2418,N_2460);
xor U2507 (N_2507,N_2408,N_2499);
nand U2508 (N_2508,N_2417,N_2462);
xor U2509 (N_2509,N_2421,N_2426);
or U2510 (N_2510,N_2469,N_2410);
nand U2511 (N_2511,N_2479,N_2443);
xor U2512 (N_2512,N_2484,N_2424);
nor U2513 (N_2513,N_2445,N_2464);
xnor U2514 (N_2514,N_2447,N_2461);
or U2515 (N_2515,N_2490,N_2477);
xor U2516 (N_2516,N_2432,N_2496);
or U2517 (N_2517,N_2478,N_2428);
nand U2518 (N_2518,N_2444,N_2498);
and U2519 (N_2519,N_2470,N_2419);
xor U2520 (N_2520,N_2483,N_2436);
nand U2521 (N_2521,N_2423,N_2494);
nand U2522 (N_2522,N_2431,N_2454);
nand U2523 (N_2523,N_2429,N_2411);
xnor U2524 (N_2524,N_2488,N_2420);
nor U2525 (N_2525,N_2492,N_2491);
nor U2526 (N_2526,N_2400,N_2497);
or U2527 (N_2527,N_2434,N_2422);
nor U2528 (N_2528,N_2425,N_2463);
xor U2529 (N_2529,N_2468,N_2427);
and U2530 (N_2530,N_2416,N_2406);
xnor U2531 (N_2531,N_2414,N_2476);
nor U2532 (N_2532,N_2465,N_2437);
nand U2533 (N_2533,N_2415,N_2401);
nor U2534 (N_2534,N_2404,N_2438);
and U2535 (N_2535,N_2455,N_2450);
nand U2536 (N_2536,N_2456,N_2493);
or U2537 (N_2537,N_2446,N_2452);
or U2538 (N_2538,N_2440,N_2471);
nand U2539 (N_2539,N_2472,N_2474);
or U2540 (N_2540,N_2435,N_2449);
and U2541 (N_2541,N_2402,N_2448);
nand U2542 (N_2542,N_2451,N_2412);
nor U2543 (N_2543,N_2495,N_2489);
and U2544 (N_2544,N_2458,N_2441);
nor U2545 (N_2545,N_2407,N_2439);
nor U2546 (N_2546,N_2485,N_2481);
and U2547 (N_2547,N_2473,N_2405);
xnor U2548 (N_2548,N_2403,N_2459);
or U2549 (N_2549,N_2442,N_2467);
and U2550 (N_2550,N_2472,N_2489);
nor U2551 (N_2551,N_2473,N_2447);
nand U2552 (N_2552,N_2439,N_2456);
xnor U2553 (N_2553,N_2433,N_2470);
and U2554 (N_2554,N_2459,N_2494);
nor U2555 (N_2555,N_2467,N_2448);
xor U2556 (N_2556,N_2499,N_2421);
xor U2557 (N_2557,N_2439,N_2458);
xnor U2558 (N_2558,N_2469,N_2431);
nor U2559 (N_2559,N_2415,N_2424);
nor U2560 (N_2560,N_2416,N_2481);
or U2561 (N_2561,N_2467,N_2426);
or U2562 (N_2562,N_2402,N_2403);
or U2563 (N_2563,N_2430,N_2443);
nand U2564 (N_2564,N_2412,N_2431);
nor U2565 (N_2565,N_2476,N_2462);
and U2566 (N_2566,N_2495,N_2407);
xor U2567 (N_2567,N_2413,N_2427);
or U2568 (N_2568,N_2407,N_2401);
nor U2569 (N_2569,N_2443,N_2418);
xnor U2570 (N_2570,N_2403,N_2450);
xnor U2571 (N_2571,N_2404,N_2466);
nand U2572 (N_2572,N_2488,N_2477);
nand U2573 (N_2573,N_2422,N_2403);
or U2574 (N_2574,N_2400,N_2418);
or U2575 (N_2575,N_2473,N_2420);
xor U2576 (N_2576,N_2467,N_2480);
nor U2577 (N_2577,N_2472,N_2403);
nand U2578 (N_2578,N_2466,N_2467);
nor U2579 (N_2579,N_2407,N_2422);
or U2580 (N_2580,N_2473,N_2431);
xnor U2581 (N_2581,N_2465,N_2469);
and U2582 (N_2582,N_2430,N_2425);
xor U2583 (N_2583,N_2449,N_2455);
nand U2584 (N_2584,N_2439,N_2476);
xor U2585 (N_2585,N_2491,N_2445);
or U2586 (N_2586,N_2402,N_2484);
or U2587 (N_2587,N_2445,N_2456);
nor U2588 (N_2588,N_2402,N_2400);
or U2589 (N_2589,N_2492,N_2461);
and U2590 (N_2590,N_2446,N_2485);
nand U2591 (N_2591,N_2405,N_2490);
nand U2592 (N_2592,N_2461,N_2467);
xor U2593 (N_2593,N_2472,N_2477);
or U2594 (N_2594,N_2495,N_2494);
nand U2595 (N_2595,N_2410,N_2491);
xnor U2596 (N_2596,N_2421,N_2469);
nand U2597 (N_2597,N_2450,N_2496);
nor U2598 (N_2598,N_2416,N_2451);
nor U2599 (N_2599,N_2496,N_2480);
xnor U2600 (N_2600,N_2577,N_2592);
nor U2601 (N_2601,N_2583,N_2542);
xor U2602 (N_2602,N_2591,N_2585);
or U2603 (N_2603,N_2539,N_2533);
and U2604 (N_2604,N_2587,N_2553);
nand U2605 (N_2605,N_2546,N_2509);
or U2606 (N_2606,N_2516,N_2595);
xnor U2607 (N_2607,N_2570,N_2568);
xor U2608 (N_2608,N_2597,N_2565);
nand U2609 (N_2609,N_2525,N_2598);
or U2610 (N_2610,N_2596,N_2523);
nor U2611 (N_2611,N_2548,N_2529);
nand U2612 (N_2612,N_2573,N_2549);
nand U2613 (N_2613,N_2531,N_2547);
xnor U2614 (N_2614,N_2508,N_2518);
xor U2615 (N_2615,N_2505,N_2522);
and U2616 (N_2616,N_2504,N_2510);
or U2617 (N_2617,N_2528,N_2527);
xor U2618 (N_2618,N_2559,N_2562);
xnor U2619 (N_2619,N_2524,N_2590);
and U2620 (N_2620,N_2535,N_2519);
nand U2621 (N_2621,N_2575,N_2507);
xor U2622 (N_2622,N_2584,N_2555);
xnor U2623 (N_2623,N_2569,N_2566);
xnor U2624 (N_2624,N_2506,N_2579);
xor U2625 (N_2625,N_2551,N_2501);
nor U2626 (N_2626,N_2530,N_2594);
xnor U2627 (N_2627,N_2544,N_2572);
or U2628 (N_2628,N_2556,N_2580);
or U2629 (N_2629,N_2532,N_2526);
xnor U2630 (N_2630,N_2557,N_2538);
nand U2631 (N_2631,N_2558,N_2581);
nor U2632 (N_2632,N_2537,N_2599);
or U2633 (N_2633,N_2513,N_2520);
xnor U2634 (N_2634,N_2554,N_2571);
and U2635 (N_2635,N_2576,N_2545);
or U2636 (N_2636,N_2563,N_2582);
nand U2637 (N_2637,N_2514,N_2541);
or U2638 (N_2638,N_2586,N_2550);
or U2639 (N_2639,N_2543,N_2588);
nor U2640 (N_2640,N_2500,N_2561);
xor U2641 (N_2641,N_2540,N_2503);
nor U2642 (N_2642,N_2517,N_2536);
xor U2643 (N_2643,N_2589,N_2512);
nand U2644 (N_2644,N_2560,N_2574);
xor U2645 (N_2645,N_2552,N_2564);
nand U2646 (N_2646,N_2511,N_2578);
xor U2647 (N_2647,N_2502,N_2567);
xnor U2648 (N_2648,N_2593,N_2534);
xor U2649 (N_2649,N_2515,N_2521);
nand U2650 (N_2650,N_2550,N_2524);
and U2651 (N_2651,N_2596,N_2527);
xor U2652 (N_2652,N_2531,N_2530);
or U2653 (N_2653,N_2564,N_2596);
nor U2654 (N_2654,N_2554,N_2517);
or U2655 (N_2655,N_2589,N_2556);
and U2656 (N_2656,N_2598,N_2527);
nor U2657 (N_2657,N_2587,N_2543);
nor U2658 (N_2658,N_2568,N_2596);
or U2659 (N_2659,N_2545,N_2530);
and U2660 (N_2660,N_2563,N_2578);
nor U2661 (N_2661,N_2552,N_2545);
nand U2662 (N_2662,N_2565,N_2520);
nand U2663 (N_2663,N_2571,N_2535);
and U2664 (N_2664,N_2536,N_2542);
nand U2665 (N_2665,N_2559,N_2545);
and U2666 (N_2666,N_2574,N_2540);
nor U2667 (N_2667,N_2541,N_2562);
nand U2668 (N_2668,N_2599,N_2588);
nor U2669 (N_2669,N_2543,N_2528);
or U2670 (N_2670,N_2574,N_2568);
nand U2671 (N_2671,N_2538,N_2599);
nand U2672 (N_2672,N_2540,N_2530);
and U2673 (N_2673,N_2547,N_2580);
or U2674 (N_2674,N_2531,N_2585);
or U2675 (N_2675,N_2504,N_2524);
and U2676 (N_2676,N_2560,N_2526);
xor U2677 (N_2677,N_2503,N_2506);
and U2678 (N_2678,N_2544,N_2549);
nor U2679 (N_2679,N_2563,N_2549);
and U2680 (N_2680,N_2577,N_2557);
xor U2681 (N_2681,N_2506,N_2555);
xnor U2682 (N_2682,N_2572,N_2540);
xnor U2683 (N_2683,N_2586,N_2558);
and U2684 (N_2684,N_2569,N_2561);
or U2685 (N_2685,N_2520,N_2547);
xnor U2686 (N_2686,N_2509,N_2517);
or U2687 (N_2687,N_2501,N_2530);
nor U2688 (N_2688,N_2555,N_2573);
and U2689 (N_2689,N_2564,N_2597);
or U2690 (N_2690,N_2517,N_2599);
and U2691 (N_2691,N_2541,N_2535);
or U2692 (N_2692,N_2513,N_2592);
nand U2693 (N_2693,N_2532,N_2579);
and U2694 (N_2694,N_2542,N_2549);
nand U2695 (N_2695,N_2568,N_2508);
and U2696 (N_2696,N_2519,N_2595);
xnor U2697 (N_2697,N_2524,N_2575);
or U2698 (N_2698,N_2587,N_2513);
or U2699 (N_2699,N_2501,N_2568);
nand U2700 (N_2700,N_2646,N_2694);
and U2701 (N_2701,N_2618,N_2634);
nor U2702 (N_2702,N_2638,N_2656);
and U2703 (N_2703,N_2643,N_2636);
or U2704 (N_2704,N_2670,N_2673);
or U2705 (N_2705,N_2681,N_2691);
nor U2706 (N_2706,N_2655,N_2642);
and U2707 (N_2707,N_2606,N_2607);
or U2708 (N_2708,N_2689,N_2684);
nand U2709 (N_2709,N_2612,N_2664);
or U2710 (N_2710,N_2666,N_2662);
nand U2711 (N_2711,N_2668,N_2609);
and U2712 (N_2712,N_2680,N_2629);
and U2713 (N_2713,N_2660,N_2632);
or U2714 (N_2714,N_2617,N_2621);
xor U2715 (N_2715,N_2603,N_2635);
xor U2716 (N_2716,N_2672,N_2622);
nor U2717 (N_2717,N_2669,N_2644);
nor U2718 (N_2718,N_2663,N_2615);
xnor U2719 (N_2719,N_2611,N_2682);
xor U2720 (N_2720,N_2686,N_2678);
and U2721 (N_2721,N_2659,N_2688);
and U2722 (N_2722,N_2661,N_2639);
and U2723 (N_2723,N_2613,N_2625);
nand U2724 (N_2724,N_2647,N_2608);
nand U2725 (N_2725,N_2620,N_2696);
and U2726 (N_2726,N_2667,N_2619);
or U2727 (N_2727,N_2699,N_2674);
nor U2728 (N_2728,N_2693,N_2695);
nand U2729 (N_2729,N_2630,N_2627);
xnor U2730 (N_2730,N_2624,N_2623);
and U2731 (N_2731,N_2676,N_2601);
nand U2732 (N_2732,N_2645,N_2665);
nor U2733 (N_2733,N_2616,N_2654);
and U2734 (N_2734,N_2626,N_2604);
or U2735 (N_2735,N_2614,N_2657);
or U2736 (N_2736,N_2697,N_2675);
xor U2737 (N_2737,N_2602,N_2671);
xor U2738 (N_2738,N_2687,N_2658);
nor U2739 (N_2739,N_2677,N_2610);
nor U2740 (N_2740,N_2683,N_2633);
nand U2741 (N_2741,N_2631,N_2652);
nor U2742 (N_2742,N_2685,N_2640);
nand U2743 (N_2743,N_2679,N_2649);
nor U2744 (N_2744,N_2648,N_2651);
or U2745 (N_2745,N_2690,N_2628);
and U2746 (N_2746,N_2698,N_2641);
nand U2747 (N_2747,N_2605,N_2692);
nor U2748 (N_2748,N_2600,N_2637);
and U2749 (N_2749,N_2650,N_2653);
nand U2750 (N_2750,N_2693,N_2649);
nand U2751 (N_2751,N_2688,N_2681);
nor U2752 (N_2752,N_2632,N_2627);
nand U2753 (N_2753,N_2690,N_2603);
or U2754 (N_2754,N_2640,N_2677);
xnor U2755 (N_2755,N_2628,N_2699);
or U2756 (N_2756,N_2678,N_2654);
nand U2757 (N_2757,N_2659,N_2653);
nand U2758 (N_2758,N_2676,N_2645);
nand U2759 (N_2759,N_2622,N_2624);
nor U2760 (N_2760,N_2674,N_2610);
xnor U2761 (N_2761,N_2614,N_2621);
nand U2762 (N_2762,N_2682,N_2659);
nand U2763 (N_2763,N_2682,N_2601);
nor U2764 (N_2764,N_2678,N_2625);
nand U2765 (N_2765,N_2685,N_2605);
nand U2766 (N_2766,N_2694,N_2641);
or U2767 (N_2767,N_2610,N_2629);
and U2768 (N_2768,N_2696,N_2651);
or U2769 (N_2769,N_2604,N_2666);
or U2770 (N_2770,N_2632,N_2691);
nand U2771 (N_2771,N_2614,N_2660);
xor U2772 (N_2772,N_2636,N_2627);
and U2773 (N_2773,N_2692,N_2651);
nand U2774 (N_2774,N_2694,N_2693);
xor U2775 (N_2775,N_2681,N_2696);
nor U2776 (N_2776,N_2619,N_2693);
xnor U2777 (N_2777,N_2692,N_2608);
xnor U2778 (N_2778,N_2636,N_2698);
xnor U2779 (N_2779,N_2660,N_2616);
and U2780 (N_2780,N_2610,N_2625);
xor U2781 (N_2781,N_2645,N_2651);
or U2782 (N_2782,N_2631,N_2644);
and U2783 (N_2783,N_2681,N_2689);
and U2784 (N_2784,N_2607,N_2630);
nand U2785 (N_2785,N_2620,N_2644);
and U2786 (N_2786,N_2610,N_2611);
and U2787 (N_2787,N_2667,N_2674);
and U2788 (N_2788,N_2614,N_2688);
nor U2789 (N_2789,N_2680,N_2627);
or U2790 (N_2790,N_2636,N_2608);
nand U2791 (N_2791,N_2600,N_2638);
nand U2792 (N_2792,N_2642,N_2650);
or U2793 (N_2793,N_2662,N_2675);
xor U2794 (N_2794,N_2631,N_2680);
and U2795 (N_2795,N_2606,N_2662);
xnor U2796 (N_2796,N_2690,N_2658);
and U2797 (N_2797,N_2613,N_2621);
nand U2798 (N_2798,N_2609,N_2682);
nand U2799 (N_2799,N_2686,N_2614);
nand U2800 (N_2800,N_2715,N_2742);
xnor U2801 (N_2801,N_2754,N_2796);
and U2802 (N_2802,N_2767,N_2729);
or U2803 (N_2803,N_2787,N_2745);
nor U2804 (N_2804,N_2708,N_2722);
or U2805 (N_2805,N_2778,N_2785);
xor U2806 (N_2806,N_2721,N_2769);
nand U2807 (N_2807,N_2711,N_2720);
xor U2808 (N_2808,N_2730,N_2740);
and U2809 (N_2809,N_2726,N_2752);
and U2810 (N_2810,N_2779,N_2755);
or U2811 (N_2811,N_2723,N_2777);
or U2812 (N_2812,N_2797,N_2799);
or U2813 (N_2813,N_2763,N_2744);
and U2814 (N_2814,N_2756,N_2751);
and U2815 (N_2815,N_2737,N_2792);
nor U2816 (N_2816,N_2781,N_2725);
and U2817 (N_2817,N_2735,N_2790);
xnor U2818 (N_2818,N_2747,N_2704);
and U2819 (N_2819,N_2727,N_2789);
and U2820 (N_2820,N_2734,N_2702);
or U2821 (N_2821,N_2782,N_2770);
nand U2822 (N_2822,N_2793,N_2718);
nand U2823 (N_2823,N_2771,N_2757);
and U2824 (N_2824,N_2741,N_2716);
nand U2825 (N_2825,N_2713,N_2794);
or U2826 (N_2826,N_2709,N_2738);
and U2827 (N_2827,N_2766,N_2795);
nor U2828 (N_2828,N_2780,N_2791);
nand U2829 (N_2829,N_2701,N_2784);
nor U2830 (N_2830,N_2762,N_2774);
or U2831 (N_2831,N_2748,N_2759);
or U2832 (N_2832,N_2773,N_2710);
nand U2833 (N_2833,N_2706,N_2775);
or U2834 (N_2834,N_2750,N_2764);
nor U2835 (N_2835,N_2761,N_2736);
and U2836 (N_2836,N_2743,N_2703);
nor U2837 (N_2837,N_2724,N_2739);
xnor U2838 (N_2838,N_2765,N_2788);
nor U2839 (N_2839,N_2700,N_2749);
and U2840 (N_2840,N_2758,N_2753);
and U2841 (N_2841,N_2705,N_2786);
and U2842 (N_2842,N_2731,N_2776);
nor U2843 (N_2843,N_2798,N_2733);
xnor U2844 (N_2844,N_2712,N_2707);
nand U2845 (N_2845,N_2714,N_2746);
and U2846 (N_2846,N_2717,N_2783);
or U2847 (N_2847,N_2768,N_2772);
nand U2848 (N_2848,N_2719,N_2732);
or U2849 (N_2849,N_2760,N_2728);
or U2850 (N_2850,N_2739,N_2798);
nor U2851 (N_2851,N_2779,N_2711);
or U2852 (N_2852,N_2772,N_2730);
nand U2853 (N_2853,N_2737,N_2782);
and U2854 (N_2854,N_2741,N_2798);
or U2855 (N_2855,N_2765,N_2796);
xor U2856 (N_2856,N_2711,N_2728);
or U2857 (N_2857,N_2785,N_2750);
nor U2858 (N_2858,N_2746,N_2733);
nand U2859 (N_2859,N_2711,N_2767);
xnor U2860 (N_2860,N_2716,N_2799);
nor U2861 (N_2861,N_2706,N_2762);
or U2862 (N_2862,N_2762,N_2794);
or U2863 (N_2863,N_2786,N_2711);
or U2864 (N_2864,N_2713,N_2771);
xor U2865 (N_2865,N_2706,N_2788);
nor U2866 (N_2866,N_2754,N_2752);
nor U2867 (N_2867,N_2708,N_2768);
or U2868 (N_2868,N_2735,N_2722);
nor U2869 (N_2869,N_2760,N_2768);
or U2870 (N_2870,N_2726,N_2747);
nor U2871 (N_2871,N_2718,N_2777);
nand U2872 (N_2872,N_2737,N_2786);
nor U2873 (N_2873,N_2751,N_2739);
and U2874 (N_2874,N_2736,N_2758);
or U2875 (N_2875,N_2748,N_2724);
and U2876 (N_2876,N_2713,N_2710);
nand U2877 (N_2877,N_2775,N_2757);
nor U2878 (N_2878,N_2704,N_2724);
and U2879 (N_2879,N_2717,N_2782);
nand U2880 (N_2880,N_2706,N_2773);
and U2881 (N_2881,N_2737,N_2719);
or U2882 (N_2882,N_2764,N_2780);
nand U2883 (N_2883,N_2702,N_2773);
xnor U2884 (N_2884,N_2742,N_2721);
nor U2885 (N_2885,N_2763,N_2756);
or U2886 (N_2886,N_2725,N_2789);
or U2887 (N_2887,N_2730,N_2749);
nand U2888 (N_2888,N_2798,N_2771);
nand U2889 (N_2889,N_2759,N_2733);
nand U2890 (N_2890,N_2780,N_2746);
nor U2891 (N_2891,N_2729,N_2782);
or U2892 (N_2892,N_2762,N_2797);
nor U2893 (N_2893,N_2796,N_2747);
nor U2894 (N_2894,N_2718,N_2745);
and U2895 (N_2895,N_2779,N_2785);
nor U2896 (N_2896,N_2748,N_2703);
or U2897 (N_2897,N_2767,N_2753);
or U2898 (N_2898,N_2788,N_2770);
xor U2899 (N_2899,N_2799,N_2758);
nor U2900 (N_2900,N_2877,N_2882);
xnor U2901 (N_2901,N_2889,N_2870);
xnor U2902 (N_2902,N_2816,N_2842);
and U2903 (N_2903,N_2843,N_2828);
nor U2904 (N_2904,N_2850,N_2830);
nand U2905 (N_2905,N_2822,N_2886);
xor U2906 (N_2906,N_2846,N_2855);
or U2907 (N_2907,N_2865,N_2861);
nand U2908 (N_2908,N_2879,N_2835);
nand U2909 (N_2909,N_2864,N_2878);
or U2910 (N_2910,N_2807,N_2805);
nor U2911 (N_2911,N_2819,N_2876);
and U2912 (N_2912,N_2893,N_2853);
nor U2913 (N_2913,N_2852,N_2894);
nand U2914 (N_2914,N_2898,N_2887);
nand U2915 (N_2915,N_2862,N_2825);
and U2916 (N_2916,N_2845,N_2847);
and U2917 (N_2917,N_2856,N_2881);
nand U2918 (N_2918,N_2818,N_2806);
nand U2919 (N_2919,N_2868,N_2884);
or U2920 (N_2920,N_2871,N_2844);
nor U2921 (N_2921,N_2866,N_2896);
or U2922 (N_2922,N_2860,N_2812);
or U2923 (N_2923,N_2869,N_2817);
nor U2924 (N_2924,N_2829,N_2854);
xnor U2925 (N_2925,N_2815,N_2891);
nor U2926 (N_2926,N_2888,N_2841);
or U2927 (N_2927,N_2823,N_2831);
or U2928 (N_2928,N_2804,N_2851);
xnor U2929 (N_2929,N_2836,N_2813);
or U2930 (N_2930,N_2834,N_2827);
and U2931 (N_2931,N_2883,N_2837);
nor U2932 (N_2932,N_2859,N_2838);
xnor U2933 (N_2933,N_2857,N_2848);
or U2934 (N_2934,N_2899,N_2849);
nor U2935 (N_2935,N_2802,N_2803);
nor U2936 (N_2936,N_2880,N_2858);
or U2937 (N_2937,N_2810,N_2820);
and U2938 (N_2938,N_2839,N_2800);
and U2939 (N_2939,N_2885,N_2801);
nor U2940 (N_2940,N_2832,N_2863);
nor U2941 (N_2941,N_2809,N_2892);
or U2942 (N_2942,N_2874,N_2873);
or U2943 (N_2943,N_2811,N_2826);
and U2944 (N_2944,N_2840,N_2814);
nor U2945 (N_2945,N_2821,N_2872);
and U2946 (N_2946,N_2824,N_2890);
or U2947 (N_2947,N_2808,N_2895);
and U2948 (N_2948,N_2875,N_2867);
and U2949 (N_2949,N_2833,N_2897);
nor U2950 (N_2950,N_2898,N_2859);
nand U2951 (N_2951,N_2860,N_2846);
and U2952 (N_2952,N_2884,N_2806);
xnor U2953 (N_2953,N_2872,N_2856);
xor U2954 (N_2954,N_2856,N_2863);
nand U2955 (N_2955,N_2895,N_2834);
or U2956 (N_2956,N_2872,N_2855);
or U2957 (N_2957,N_2877,N_2876);
xnor U2958 (N_2958,N_2828,N_2825);
or U2959 (N_2959,N_2825,N_2851);
nor U2960 (N_2960,N_2829,N_2873);
and U2961 (N_2961,N_2830,N_2889);
and U2962 (N_2962,N_2829,N_2821);
nor U2963 (N_2963,N_2831,N_2844);
nor U2964 (N_2964,N_2896,N_2877);
nor U2965 (N_2965,N_2898,N_2899);
nor U2966 (N_2966,N_2850,N_2881);
nor U2967 (N_2967,N_2859,N_2844);
xnor U2968 (N_2968,N_2846,N_2826);
nand U2969 (N_2969,N_2888,N_2871);
nor U2970 (N_2970,N_2894,N_2887);
nor U2971 (N_2971,N_2823,N_2871);
nand U2972 (N_2972,N_2805,N_2886);
nor U2973 (N_2973,N_2850,N_2845);
nand U2974 (N_2974,N_2810,N_2800);
nand U2975 (N_2975,N_2841,N_2894);
or U2976 (N_2976,N_2877,N_2819);
xnor U2977 (N_2977,N_2821,N_2831);
and U2978 (N_2978,N_2881,N_2832);
xor U2979 (N_2979,N_2865,N_2801);
nand U2980 (N_2980,N_2890,N_2880);
nand U2981 (N_2981,N_2858,N_2877);
xor U2982 (N_2982,N_2898,N_2806);
and U2983 (N_2983,N_2842,N_2866);
nand U2984 (N_2984,N_2867,N_2880);
and U2985 (N_2985,N_2872,N_2816);
and U2986 (N_2986,N_2896,N_2820);
nand U2987 (N_2987,N_2858,N_2807);
or U2988 (N_2988,N_2840,N_2892);
nand U2989 (N_2989,N_2874,N_2857);
and U2990 (N_2990,N_2820,N_2850);
nand U2991 (N_2991,N_2878,N_2832);
or U2992 (N_2992,N_2861,N_2896);
xnor U2993 (N_2993,N_2812,N_2835);
or U2994 (N_2994,N_2884,N_2824);
and U2995 (N_2995,N_2811,N_2896);
nand U2996 (N_2996,N_2805,N_2870);
or U2997 (N_2997,N_2824,N_2867);
nand U2998 (N_2998,N_2883,N_2849);
and U2999 (N_2999,N_2848,N_2889);
nand U3000 (N_3000,N_2966,N_2901);
xor U3001 (N_3001,N_2915,N_2985);
nor U3002 (N_3002,N_2955,N_2958);
and U3003 (N_3003,N_2935,N_2991);
nand U3004 (N_3004,N_2971,N_2943);
nand U3005 (N_3005,N_2929,N_2983);
and U3006 (N_3006,N_2986,N_2946);
xor U3007 (N_3007,N_2988,N_2914);
and U3008 (N_3008,N_2924,N_2904);
nor U3009 (N_3009,N_2994,N_2930);
and U3010 (N_3010,N_2960,N_2941);
nand U3011 (N_3011,N_2997,N_2905);
and U3012 (N_3012,N_2931,N_2973);
xor U3013 (N_3013,N_2964,N_2993);
nor U3014 (N_3014,N_2977,N_2992);
or U3015 (N_3015,N_2974,N_2956);
nand U3016 (N_3016,N_2954,N_2945);
nand U3017 (N_3017,N_2987,N_2921);
nor U3018 (N_3018,N_2919,N_2989);
and U3019 (N_3019,N_2969,N_2912);
nor U3020 (N_3020,N_2976,N_2916);
xnor U3021 (N_3021,N_2962,N_2937);
nor U3022 (N_3022,N_2951,N_2996);
xor U3023 (N_3023,N_2952,N_2907);
nand U3024 (N_3024,N_2982,N_2963);
nor U3025 (N_3025,N_2910,N_2925);
or U3026 (N_3026,N_2970,N_2936);
nor U3027 (N_3027,N_2965,N_2984);
nor U3028 (N_3028,N_2926,N_2902);
nand U3029 (N_3029,N_2918,N_2940);
nor U3030 (N_3030,N_2903,N_2932);
nor U3031 (N_3031,N_2900,N_2959);
and U3032 (N_3032,N_2995,N_2979);
or U3033 (N_3033,N_2949,N_2933);
nor U3034 (N_3034,N_2980,N_2978);
nor U3035 (N_3035,N_2922,N_2981);
and U3036 (N_3036,N_2927,N_2938);
nand U3037 (N_3037,N_2906,N_2999);
nand U3038 (N_3038,N_2947,N_2948);
nand U3039 (N_3039,N_2967,N_2913);
or U3040 (N_3040,N_2961,N_2950);
or U3041 (N_3041,N_2968,N_2944);
nor U3042 (N_3042,N_2990,N_2957);
or U3043 (N_3043,N_2917,N_2908);
and U3044 (N_3044,N_2939,N_2909);
xor U3045 (N_3045,N_2998,N_2975);
and U3046 (N_3046,N_2923,N_2953);
and U3047 (N_3047,N_2934,N_2942);
and U3048 (N_3048,N_2972,N_2911);
nor U3049 (N_3049,N_2928,N_2920);
nand U3050 (N_3050,N_2910,N_2930);
nor U3051 (N_3051,N_2907,N_2981);
nor U3052 (N_3052,N_2915,N_2948);
or U3053 (N_3053,N_2906,N_2993);
nor U3054 (N_3054,N_2998,N_2916);
nor U3055 (N_3055,N_2962,N_2966);
and U3056 (N_3056,N_2989,N_2960);
nand U3057 (N_3057,N_2940,N_2964);
or U3058 (N_3058,N_2914,N_2900);
nor U3059 (N_3059,N_2930,N_2991);
xor U3060 (N_3060,N_2919,N_2960);
xor U3061 (N_3061,N_2958,N_2943);
and U3062 (N_3062,N_2956,N_2983);
and U3063 (N_3063,N_2999,N_2968);
or U3064 (N_3064,N_2997,N_2987);
or U3065 (N_3065,N_2912,N_2945);
or U3066 (N_3066,N_2964,N_2920);
nand U3067 (N_3067,N_2969,N_2990);
nor U3068 (N_3068,N_2974,N_2994);
nand U3069 (N_3069,N_2994,N_2916);
xnor U3070 (N_3070,N_2965,N_2950);
xor U3071 (N_3071,N_2983,N_2928);
and U3072 (N_3072,N_2985,N_2973);
xnor U3073 (N_3073,N_2961,N_2983);
and U3074 (N_3074,N_2996,N_2925);
xnor U3075 (N_3075,N_2988,N_2985);
nor U3076 (N_3076,N_2994,N_2981);
and U3077 (N_3077,N_2975,N_2935);
nor U3078 (N_3078,N_2964,N_2945);
and U3079 (N_3079,N_2964,N_2929);
and U3080 (N_3080,N_2945,N_2934);
xor U3081 (N_3081,N_2909,N_2902);
and U3082 (N_3082,N_2928,N_2903);
nand U3083 (N_3083,N_2976,N_2943);
or U3084 (N_3084,N_2939,N_2942);
nor U3085 (N_3085,N_2928,N_2932);
or U3086 (N_3086,N_2938,N_2919);
nand U3087 (N_3087,N_2989,N_2966);
and U3088 (N_3088,N_2942,N_2994);
or U3089 (N_3089,N_2962,N_2907);
and U3090 (N_3090,N_2955,N_2917);
xor U3091 (N_3091,N_2975,N_2989);
or U3092 (N_3092,N_2981,N_2923);
or U3093 (N_3093,N_2969,N_2929);
nand U3094 (N_3094,N_2975,N_2946);
xnor U3095 (N_3095,N_2971,N_2921);
nand U3096 (N_3096,N_2952,N_2900);
nand U3097 (N_3097,N_2934,N_2905);
nand U3098 (N_3098,N_2934,N_2929);
and U3099 (N_3099,N_2995,N_2919);
or U3100 (N_3100,N_3032,N_3052);
nand U3101 (N_3101,N_3029,N_3003);
nand U3102 (N_3102,N_3037,N_3038);
xnor U3103 (N_3103,N_3077,N_3014);
xor U3104 (N_3104,N_3082,N_3024);
xor U3105 (N_3105,N_3019,N_3027);
nor U3106 (N_3106,N_3018,N_3060);
nand U3107 (N_3107,N_3083,N_3086);
or U3108 (N_3108,N_3066,N_3084);
xnor U3109 (N_3109,N_3067,N_3042);
or U3110 (N_3110,N_3062,N_3061);
or U3111 (N_3111,N_3025,N_3089);
xor U3112 (N_3112,N_3046,N_3006);
xor U3113 (N_3113,N_3033,N_3043);
nor U3114 (N_3114,N_3073,N_3068);
and U3115 (N_3115,N_3090,N_3048);
nand U3116 (N_3116,N_3034,N_3064);
nor U3117 (N_3117,N_3041,N_3045);
xor U3118 (N_3118,N_3008,N_3055);
nand U3119 (N_3119,N_3030,N_3035);
or U3120 (N_3120,N_3007,N_3010);
nor U3121 (N_3121,N_3097,N_3092);
and U3122 (N_3122,N_3071,N_3085);
nor U3123 (N_3123,N_3004,N_3059);
nor U3124 (N_3124,N_3021,N_3031);
or U3125 (N_3125,N_3057,N_3050);
and U3126 (N_3126,N_3088,N_3076);
or U3127 (N_3127,N_3099,N_3087);
nor U3128 (N_3128,N_3074,N_3016);
nand U3129 (N_3129,N_3070,N_3023);
nor U3130 (N_3130,N_3056,N_3098);
or U3131 (N_3131,N_3000,N_3079);
xor U3132 (N_3132,N_3051,N_3081);
nor U3133 (N_3133,N_3040,N_3049);
and U3134 (N_3134,N_3095,N_3020);
nand U3135 (N_3135,N_3069,N_3065);
and U3136 (N_3136,N_3093,N_3053);
and U3137 (N_3137,N_3047,N_3080);
nor U3138 (N_3138,N_3044,N_3058);
and U3139 (N_3139,N_3096,N_3012);
nor U3140 (N_3140,N_3091,N_3054);
xor U3141 (N_3141,N_3001,N_3036);
nor U3142 (N_3142,N_3017,N_3094);
and U3143 (N_3143,N_3072,N_3026);
xor U3144 (N_3144,N_3009,N_3028);
xor U3145 (N_3145,N_3013,N_3005);
xor U3146 (N_3146,N_3075,N_3015);
or U3147 (N_3147,N_3039,N_3002);
or U3148 (N_3148,N_3011,N_3022);
nand U3149 (N_3149,N_3063,N_3078);
xor U3150 (N_3150,N_3081,N_3030);
and U3151 (N_3151,N_3068,N_3092);
or U3152 (N_3152,N_3084,N_3047);
or U3153 (N_3153,N_3095,N_3001);
nand U3154 (N_3154,N_3021,N_3004);
and U3155 (N_3155,N_3042,N_3091);
or U3156 (N_3156,N_3000,N_3039);
xor U3157 (N_3157,N_3034,N_3043);
xor U3158 (N_3158,N_3066,N_3047);
nor U3159 (N_3159,N_3060,N_3084);
and U3160 (N_3160,N_3061,N_3014);
or U3161 (N_3161,N_3087,N_3041);
and U3162 (N_3162,N_3002,N_3010);
or U3163 (N_3163,N_3016,N_3062);
nor U3164 (N_3164,N_3091,N_3045);
nor U3165 (N_3165,N_3016,N_3018);
and U3166 (N_3166,N_3038,N_3078);
and U3167 (N_3167,N_3074,N_3025);
or U3168 (N_3168,N_3034,N_3054);
xnor U3169 (N_3169,N_3043,N_3008);
xor U3170 (N_3170,N_3028,N_3012);
and U3171 (N_3171,N_3020,N_3021);
nand U3172 (N_3172,N_3056,N_3023);
or U3173 (N_3173,N_3029,N_3000);
nor U3174 (N_3174,N_3068,N_3001);
nand U3175 (N_3175,N_3074,N_3064);
or U3176 (N_3176,N_3025,N_3033);
and U3177 (N_3177,N_3054,N_3068);
xnor U3178 (N_3178,N_3069,N_3016);
nor U3179 (N_3179,N_3062,N_3056);
and U3180 (N_3180,N_3073,N_3005);
nor U3181 (N_3181,N_3091,N_3052);
xor U3182 (N_3182,N_3081,N_3002);
nand U3183 (N_3183,N_3092,N_3046);
xor U3184 (N_3184,N_3001,N_3094);
nand U3185 (N_3185,N_3048,N_3002);
nor U3186 (N_3186,N_3054,N_3021);
and U3187 (N_3187,N_3099,N_3034);
and U3188 (N_3188,N_3061,N_3019);
nand U3189 (N_3189,N_3075,N_3091);
xor U3190 (N_3190,N_3072,N_3004);
nor U3191 (N_3191,N_3014,N_3026);
or U3192 (N_3192,N_3026,N_3065);
xnor U3193 (N_3193,N_3057,N_3021);
nand U3194 (N_3194,N_3085,N_3060);
or U3195 (N_3195,N_3087,N_3002);
and U3196 (N_3196,N_3027,N_3078);
nand U3197 (N_3197,N_3099,N_3024);
nand U3198 (N_3198,N_3068,N_3007);
and U3199 (N_3199,N_3086,N_3074);
or U3200 (N_3200,N_3173,N_3135);
or U3201 (N_3201,N_3104,N_3124);
xnor U3202 (N_3202,N_3139,N_3133);
or U3203 (N_3203,N_3149,N_3161);
nand U3204 (N_3204,N_3136,N_3175);
nor U3205 (N_3205,N_3153,N_3103);
and U3206 (N_3206,N_3174,N_3163);
nor U3207 (N_3207,N_3188,N_3117);
nand U3208 (N_3208,N_3123,N_3154);
xor U3209 (N_3209,N_3162,N_3170);
or U3210 (N_3210,N_3131,N_3166);
xnor U3211 (N_3211,N_3197,N_3180);
nand U3212 (N_3212,N_3198,N_3119);
nand U3213 (N_3213,N_3129,N_3140);
nand U3214 (N_3214,N_3101,N_3191);
nor U3215 (N_3215,N_3179,N_3134);
and U3216 (N_3216,N_3195,N_3115);
or U3217 (N_3217,N_3107,N_3121);
or U3218 (N_3218,N_3185,N_3165);
nand U3219 (N_3219,N_3194,N_3110);
nor U3220 (N_3220,N_3168,N_3146);
and U3221 (N_3221,N_3184,N_3176);
nor U3222 (N_3222,N_3105,N_3177);
nor U3223 (N_3223,N_3196,N_3144);
or U3224 (N_3224,N_3187,N_3112);
nor U3225 (N_3225,N_3156,N_3141);
and U3226 (N_3226,N_3158,N_3169);
nor U3227 (N_3227,N_3199,N_3183);
nor U3228 (N_3228,N_3102,N_3147);
xor U3229 (N_3229,N_3152,N_3181);
or U3230 (N_3230,N_3108,N_3128);
and U3231 (N_3231,N_3172,N_3122);
and U3232 (N_3232,N_3125,N_3114);
and U3233 (N_3233,N_3137,N_3148);
nand U3234 (N_3234,N_3130,N_3171);
nor U3235 (N_3235,N_3145,N_3155);
nand U3236 (N_3236,N_3127,N_3150);
xor U3237 (N_3237,N_3100,N_3111);
and U3238 (N_3238,N_3157,N_3118);
and U3239 (N_3239,N_3106,N_3160);
or U3240 (N_3240,N_3109,N_3167);
or U3241 (N_3241,N_3126,N_3143);
nand U3242 (N_3242,N_3193,N_3113);
nand U3243 (N_3243,N_3189,N_3142);
nor U3244 (N_3244,N_3159,N_3178);
nor U3245 (N_3245,N_3138,N_3186);
xnor U3246 (N_3246,N_3190,N_3132);
xor U3247 (N_3247,N_3182,N_3120);
and U3248 (N_3248,N_3151,N_3116);
and U3249 (N_3249,N_3164,N_3192);
nand U3250 (N_3250,N_3191,N_3116);
or U3251 (N_3251,N_3106,N_3139);
nand U3252 (N_3252,N_3106,N_3166);
nor U3253 (N_3253,N_3148,N_3112);
xnor U3254 (N_3254,N_3170,N_3108);
or U3255 (N_3255,N_3193,N_3131);
and U3256 (N_3256,N_3160,N_3108);
nor U3257 (N_3257,N_3125,N_3187);
nand U3258 (N_3258,N_3144,N_3187);
nand U3259 (N_3259,N_3129,N_3144);
xnor U3260 (N_3260,N_3162,N_3193);
nand U3261 (N_3261,N_3163,N_3189);
nand U3262 (N_3262,N_3118,N_3165);
nand U3263 (N_3263,N_3110,N_3172);
nor U3264 (N_3264,N_3164,N_3188);
and U3265 (N_3265,N_3192,N_3156);
and U3266 (N_3266,N_3132,N_3127);
xor U3267 (N_3267,N_3105,N_3141);
or U3268 (N_3268,N_3190,N_3152);
or U3269 (N_3269,N_3105,N_3131);
and U3270 (N_3270,N_3181,N_3104);
and U3271 (N_3271,N_3143,N_3101);
xor U3272 (N_3272,N_3178,N_3193);
nand U3273 (N_3273,N_3183,N_3144);
nand U3274 (N_3274,N_3145,N_3162);
nor U3275 (N_3275,N_3116,N_3127);
xnor U3276 (N_3276,N_3114,N_3106);
xnor U3277 (N_3277,N_3182,N_3127);
or U3278 (N_3278,N_3162,N_3137);
nand U3279 (N_3279,N_3120,N_3103);
nor U3280 (N_3280,N_3122,N_3170);
xnor U3281 (N_3281,N_3177,N_3195);
xor U3282 (N_3282,N_3194,N_3149);
nand U3283 (N_3283,N_3182,N_3192);
nand U3284 (N_3284,N_3153,N_3135);
nand U3285 (N_3285,N_3181,N_3188);
nand U3286 (N_3286,N_3170,N_3105);
and U3287 (N_3287,N_3155,N_3159);
and U3288 (N_3288,N_3140,N_3138);
nor U3289 (N_3289,N_3140,N_3175);
nor U3290 (N_3290,N_3184,N_3177);
xor U3291 (N_3291,N_3188,N_3191);
nor U3292 (N_3292,N_3192,N_3128);
xor U3293 (N_3293,N_3154,N_3120);
or U3294 (N_3294,N_3188,N_3130);
nand U3295 (N_3295,N_3120,N_3138);
or U3296 (N_3296,N_3101,N_3152);
and U3297 (N_3297,N_3166,N_3119);
nor U3298 (N_3298,N_3147,N_3172);
or U3299 (N_3299,N_3191,N_3125);
nor U3300 (N_3300,N_3251,N_3289);
xnor U3301 (N_3301,N_3259,N_3287);
xnor U3302 (N_3302,N_3241,N_3204);
or U3303 (N_3303,N_3237,N_3214);
or U3304 (N_3304,N_3268,N_3239);
xor U3305 (N_3305,N_3226,N_3276);
or U3306 (N_3306,N_3200,N_3291);
or U3307 (N_3307,N_3299,N_3258);
nor U3308 (N_3308,N_3246,N_3283);
nand U3309 (N_3309,N_3278,N_3224);
and U3310 (N_3310,N_3247,N_3207);
and U3311 (N_3311,N_3218,N_3266);
nand U3312 (N_3312,N_3275,N_3231);
nand U3313 (N_3313,N_3205,N_3229);
nor U3314 (N_3314,N_3265,N_3220);
nor U3315 (N_3315,N_3236,N_3264);
xor U3316 (N_3316,N_3277,N_3271);
or U3317 (N_3317,N_3202,N_3263);
nor U3318 (N_3318,N_3221,N_3279);
nand U3319 (N_3319,N_3274,N_3296);
and U3320 (N_3320,N_3273,N_3282);
or U3321 (N_3321,N_3219,N_3222);
nand U3322 (N_3322,N_3206,N_3249);
nor U3323 (N_3323,N_3217,N_3216);
nand U3324 (N_3324,N_3234,N_3223);
xor U3325 (N_3325,N_3252,N_3248);
xnor U3326 (N_3326,N_3280,N_3250);
and U3327 (N_3327,N_3269,N_3244);
and U3328 (N_3328,N_3285,N_3215);
or U3329 (N_3329,N_3270,N_3213);
or U3330 (N_3330,N_3260,N_3209);
nand U3331 (N_3331,N_3211,N_3253);
xnor U3332 (N_3332,N_3230,N_3228);
nor U3333 (N_3333,N_3261,N_3243);
nor U3334 (N_3334,N_3297,N_3235);
nand U3335 (N_3335,N_3212,N_3293);
nor U3336 (N_3336,N_3290,N_3267);
nor U3337 (N_3337,N_3257,N_3281);
xor U3338 (N_3338,N_3262,N_3242);
xor U3339 (N_3339,N_3272,N_3295);
and U3340 (N_3340,N_3286,N_3238);
nor U3341 (N_3341,N_3294,N_3292);
nor U3342 (N_3342,N_3208,N_3288);
nor U3343 (N_3343,N_3255,N_3232);
xnor U3344 (N_3344,N_3245,N_3233);
and U3345 (N_3345,N_3203,N_3256);
xor U3346 (N_3346,N_3284,N_3298);
and U3347 (N_3347,N_3254,N_3225);
or U3348 (N_3348,N_3201,N_3227);
nor U3349 (N_3349,N_3240,N_3210);
and U3350 (N_3350,N_3211,N_3228);
or U3351 (N_3351,N_3267,N_3275);
or U3352 (N_3352,N_3287,N_3251);
and U3353 (N_3353,N_3294,N_3273);
and U3354 (N_3354,N_3213,N_3257);
xor U3355 (N_3355,N_3242,N_3217);
and U3356 (N_3356,N_3233,N_3282);
xnor U3357 (N_3357,N_3235,N_3261);
nand U3358 (N_3358,N_3211,N_3230);
xnor U3359 (N_3359,N_3244,N_3282);
nor U3360 (N_3360,N_3236,N_3258);
xor U3361 (N_3361,N_3265,N_3212);
nor U3362 (N_3362,N_3241,N_3297);
or U3363 (N_3363,N_3266,N_3206);
nor U3364 (N_3364,N_3261,N_3286);
nand U3365 (N_3365,N_3248,N_3233);
xnor U3366 (N_3366,N_3231,N_3237);
nand U3367 (N_3367,N_3221,N_3299);
nand U3368 (N_3368,N_3273,N_3200);
xnor U3369 (N_3369,N_3226,N_3245);
or U3370 (N_3370,N_3210,N_3262);
or U3371 (N_3371,N_3221,N_3298);
and U3372 (N_3372,N_3296,N_3277);
nor U3373 (N_3373,N_3289,N_3291);
and U3374 (N_3374,N_3211,N_3257);
nor U3375 (N_3375,N_3201,N_3287);
or U3376 (N_3376,N_3240,N_3278);
xnor U3377 (N_3377,N_3230,N_3284);
nor U3378 (N_3378,N_3234,N_3252);
nor U3379 (N_3379,N_3261,N_3238);
nor U3380 (N_3380,N_3205,N_3208);
or U3381 (N_3381,N_3284,N_3288);
xnor U3382 (N_3382,N_3285,N_3239);
or U3383 (N_3383,N_3218,N_3233);
nand U3384 (N_3384,N_3251,N_3248);
or U3385 (N_3385,N_3297,N_3252);
nand U3386 (N_3386,N_3230,N_3252);
nor U3387 (N_3387,N_3222,N_3206);
xnor U3388 (N_3388,N_3239,N_3243);
xor U3389 (N_3389,N_3273,N_3209);
xor U3390 (N_3390,N_3241,N_3266);
xnor U3391 (N_3391,N_3227,N_3276);
or U3392 (N_3392,N_3234,N_3278);
and U3393 (N_3393,N_3211,N_3284);
nor U3394 (N_3394,N_3265,N_3278);
nand U3395 (N_3395,N_3276,N_3206);
nand U3396 (N_3396,N_3258,N_3286);
or U3397 (N_3397,N_3233,N_3227);
nand U3398 (N_3398,N_3217,N_3200);
or U3399 (N_3399,N_3297,N_3261);
nand U3400 (N_3400,N_3306,N_3399);
and U3401 (N_3401,N_3325,N_3355);
xor U3402 (N_3402,N_3380,N_3385);
and U3403 (N_3403,N_3345,N_3395);
nor U3404 (N_3404,N_3330,N_3309);
nor U3405 (N_3405,N_3373,N_3313);
and U3406 (N_3406,N_3320,N_3369);
or U3407 (N_3407,N_3342,N_3336);
nor U3408 (N_3408,N_3370,N_3347);
nand U3409 (N_3409,N_3346,N_3358);
nand U3410 (N_3410,N_3311,N_3397);
or U3411 (N_3411,N_3322,N_3389);
or U3412 (N_3412,N_3337,N_3374);
nor U3413 (N_3413,N_3378,N_3367);
nor U3414 (N_3414,N_3383,N_3318);
nand U3415 (N_3415,N_3387,N_3398);
nor U3416 (N_3416,N_3390,N_3381);
or U3417 (N_3417,N_3308,N_3341);
xor U3418 (N_3418,N_3331,N_3328);
and U3419 (N_3419,N_3327,N_3365);
nand U3420 (N_3420,N_3307,N_3393);
or U3421 (N_3421,N_3363,N_3372);
nor U3422 (N_3422,N_3319,N_3377);
xor U3423 (N_3423,N_3379,N_3350);
nand U3424 (N_3424,N_3303,N_3302);
and U3425 (N_3425,N_3338,N_3304);
nand U3426 (N_3426,N_3315,N_3324);
or U3427 (N_3427,N_3368,N_3352);
nor U3428 (N_3428,N_3312,N_3386);
nand U3429 (N_3429,N_3332,N_3323);
and U3430 (N_3430,N_3366,N_3348);
and U3431 (N_3431,N_3344,N_3392);
nor U3432 (N_3432,N_3333,N_3305);
xnor U3433 (N_3433,N_3301,N_3317);
nor U3434 (N_3434,N_3354,N_3316);
nand U3435 (N_3435,N_3339,N_3310);
nor U3436 (N_3436,N_3340,N_3362);
xor U3437 (N_3437,N_3391,N_3357);
nand U3438 (N_3438,N_3382,N_3376);
or U3439 (N_3439,N_3353,N_3356);
and U3440 (N_3440,N_3351,N_3394);
and U3441 (N_3441,N_3321,N_3361);
and U3442 (N_3442,N_3375,N_3335);
and U3443 (N_3443,N_3371,N_3349);
or U3444 (N_3444,N_3343,N_3364);
nand U3445 (N_3445,N_3326,N_3360);
xnor U3446 (N_3446,N_3329,N_3334);
nand U3447 (N_3447,N_3359,N_3388);
nand U3448 (N_3448,N_3384,N_3396);
and U3449 (N_3449,N_3300,N_3314);
and U3450 (N_3450,N_3307,N_3357);
nor U3451 (N_3451,N_3399,N_3314);
xor U3452 (N_3452,N_3338,N_3320);
and U3453 (N_3453,N_3385,N_3350);
or U3454 (N_3454,N_3312,N_3367);
nand U3455 (N_3455,N_3306,N_3350);
or U3456 (N_3456,N_3302,N_3349);
and U3457 (N_3457,N_3309,N_3393);
and U3458 (N_3458,N_3355,N_3388);
and U3459 (N_3459,N_3324,N_3318);
nand U3460 (N_3460,N_3354,N_3389);
xor U3461 (N_3461,N_3367,N_3395);
and U3462 (N_3462,N_3313,N_3332);
and U3463 (N_3463,N_3339,N_3309);
and U3464 (N_3464,N_3374,N_3386);
xnor U3465 (N_3465,N_3391,N_3311);
nand U3466 (N_3466,N_3390,N_3373);
nand U3467 (N_3467,N_3300,N_3346);
and U3468 (N_3468,N_3385,N_3358);
nand U3469 (N_3469,N_3301,N_3367);
xor U3470 (N_3470,N_3366,N_3321);
xor U3471 (N_3471,N_3350,N_3381);
or U3472 (N_3472,N_3354,N_3362);
nor U3473 (N_3473,N_3343,N_3317);
nor U3474 (N_3474,N_3349,N_3398);
xor U3475 (N_3475,N_3352,N_3333);
and U3476 (N_3476,N_3327,N_3306);
nand U3477 (N_3477,N_3317,N_3313);
nand U3478 (N_3478,N_3357,N_3383);
nand U3479 (N_3479,N_3366,N_3342);
or U3480 (N_3480,N_3331,N_3387);
nor U3481 (N_3481,N_3348,N_3393);
and U3482 (N_3482,N_3319,N_3302);
and U3483 (N_3483,N_3339,N_3370);
and U3484 (N_3484,N_3322,N_3343);
nand U3485 (N_3485,N_3393,N_3391);
xor U3486 (N_3486,N_3302,N_3388);
nor U3487 (N_3487,N_3340,N_3361);
nand U3488 (N_3488,N_3361,N_3356);
xnor U3489 (N_3489,N_3326,N_3344);
xnor U3490 (N_3490,N_3331,N_3355);
xor U3491 (N_3491,N_3362,N_3376);
xor U3492 (N_3492,N_3389,N_3349);
or U3493 (N_3493,N_3360,N_3393);
xor U3494 (N_3494,N_3338,N_3315);
or U3495 (N_3495,N_3313,N_3327);
nor U3496 (N_3496,N_3337,N_3384);
xor U3497 (N_3497,N_3337,N_3350);
and U3498 (N_3498,N_3376,N_3313);
nand U3499 (N_3499,N_3335,N_3319);
nand U3500 (N_3500,N_3417,N_3438);
and U3501 (N_3501,N_3403,N_3428);
or U3502 (N_3502,N_3414,N_3466);
nand U3503 (N_3503,N_3456,N_3494);
nor U3504 (N_3504,N_3479,N_3446);
and U3505 (N_3505,N_3459,N_3483);
nand U3506 (N_3506,N_3407,N_3435);
and U3507 (N_3507,N_3468,N_3424);
nor U3508 (N_3508,N_3496,N_3411);
or U3509 (N_3509,N_3488,N_3493);
xor U3510 (N_3510,N_3465,N_3453);
nand U3511 (N_3511,N_3418,N_3480);
and U3512 (N_3512,N_3476,N_3422);
nor U3513 (N_3513,N_3463,N_3439);
nor U3514 (N_3514,N_3409,N_3481);
nor U3515 (N_3515,N_3487,N_3464);
xor U3516 (N_3516,N_3484,N_3499);
xnor U3517 (N_3517,N_3443,N_3477);
or U3518 (N_3518,N_3426,N_3400);
xor U3519 (N_3519,N_3490,N_3429);
xor U3520 (N_3520,N_3401,N_3420);
or U3521 (N_3521,N_3478,N_3469);
or U3522 (N_3522,N_3449,N_3437);
xnor U3523 (N_3523,N_3444,N_3408);
nor U3524 (N_3524,N_3434,N_3457);
or U3525 (N_3525,N_3460,N_3402);
and U3526 (N_3526,N_3495,N_3406);
nand U3527 (N_3527,N_3431,N_3492);
xnor U3528 (N_3528,N_3433,N_3410);
nor U3529 (N_3529,N_3421,N_3445);
nor U3530 (N_3530,N_3454,N_3455);
nand U3531 (N_3531,N_3472,N_3475);
nand U3532 (N_3532,N_3440,N_3427);
and U3533 (N_3533,N_3474,N_3497);
nor U3534 (N_3534,N_3432,N_3425);
xor U3535 (N_3535,N_3442,N_3451);
and U3536 (N_3536,N_3412,N_3467);
or U3537 (N_3537,N_3491,N_3489);
and U3538 (N_3538,N_3415,N_3405);
nor U3539 (N_3539,N_3419,N_3462);
or U3540 (N_3540,N_3447,N_3450);
nor U3541 (N_3541,N_3423,N_3482);
nor U3542 (N_3542,N_3498,N_3486);
nor U3543 (N_3543,N_3461,N_3473);
and U3544 (N_3544,N_3441,N_3452);
or U3545 (N_3545,N_3430,N_3416);
nand U3546 (N_3546,N_3470,N_3448);
and U3547 (N_3547,N_3485,N_3436);
xor U3548 (N_3548,N_3404,N_3458);
or U3549 (N_3549,N_3413,N_3471);
xnor U3550 (N_3550,N_3463,N_3425);
nor U3551 (N_3551,N_3418,N_3484);
or U3552 (N_3552,N_3495,N_3498);
and U3553 (N_3553,N_3461,N_3499);
and U3554 (N_3554,N_3412,N_3400);
nand U3555 (N_3555,N_3447,N_3416);
nor U3556 (N_3556,N_3494,N_3441);
xor U3557 (N_3557,N_3465,N_3488);
and U3558 (N_3558,N_3427,N_3442);
nor U3559 (N_3559,N_3494,N_3405);
nor U3560 (N_3560,N_3472,N_3479);
xor U3561 (N_3561,N_3460,N_3489);
nand U3562 (N_3562,N_3421,N_3451);
xnor U3563 (N_3563,N_3476,N_3497);
or U3564 (N_3564,N_3484,N_3472);
and U3565 (N_3565,N_3441,N_3474);
nor U3566 (N_3566,N_3430,N_3499);
nand U3567 (N_3567,N_3496,N_3456);
xor U3568 (N_3568,N_3410,N_3447);
or U3569 (N_3569,N_3472,N_3496);
xnor U3570 (N_3570,N_3495,N_3491);
or U3571 (N_3571,N_3499,N_3445);
nand U3572 (N_3572,N_3445,N_3454);
xnor U3573 (N_3573,N_3486,N_3482);
nand U3574 (N_3574,N_3459,N_3471);
xnor U3575 (N_3575,N_3435,N_3448);
and U3576 (N_3576,N_3473,N_3452);
xnor U3577 (N_3577,N_3483,N_3486);
nand U3578 (N_3578,N_3423,N_3481);
xnor U3579 (N_3579,N_3429,N_3413);
xor U3580 (N_3580,N_3441,N_3432);
xor U3581 (N_3581,N_3479,N_3495);
or U3582 (N_3582,N_3411,N_3484);
nor U3583 (N_3583,N_3481,N_3490);
and U3584 (N_3584,N_3430,N_3478);
nor U3585 (N_3585,N_3450,N_3451);
or U3586 (N_3586,N_3412,N_3480);
and U3587 (N_3587,N_3455,N_3496);
nand U3588 (N_3588,N_3476,N_3464);
xor U3589 (N_3589,N_3400,N_3414);
or U3590 (N_3590,N_3426,N_3415);
or U3591 (N_3591,N_3422,N_3407);
and U3592 (N_3592,N_3469,N_3402);
or U3593 (N_3593,N_3486,N_3466);
xnor U3594 (N_3594,N_3438,N_3436);
nor U3595 (N_3595,N_3414,N_3478);
nor U3596 (N_3596,N_3436,N_3454);
or U3597 (N_3597,N_3419,N_3485);
and U3598 (N_3598,N_3422,N_3430);
or U3599 (N_3599,N_3408,N_3463);
and U3600 (N_3600,N_3569,N_3572);
nor U3601 (N_3601,N_3511,N_3563);
and U3602 (N_3602,N_3500,N_3595);
nand U3603 (N_3603,N_3564,N_3545);
or U3604 (N_3604,N_3559,N_3532);
nor U3605 (N_3605,N_3503,N_3535);
and U3606 (N_3606,N_3538,N_3547);
or U3607 (N_3607,N_3591,N_3548);
nand U3608 (N_3608,N_3576,N_3558);
and U3609 (N_3609,N_3575,N_3554);
xnor U3610 (N_3610,N_3597,N_3593);
or U3611 (N_3611,N_3516,N_3555);
and U3612 (N_3612,N_3530,N_3537);
nand U3613 (N_3613,N_3514,N_3579);
or U3614 (N_3614,N_3562,N_3549);
xor U3615 (N_3615,N_3525,N_3501);
xor U3616 (N_3616,N_3574,N_3518);
and U3617 (N_3617,N_3542,N_3578);
and U3618 (N_3618,N_3567,N_3521);
nor U3619 (N_3619,N_3546,N_3517);
xor U3620 (N_3620,N_3539,N_3541);
nor U3621 (N_3621,N_3553,N_3582);
xnor U3622 (N_3622,N_3506,N_3589);
or U3623 (N_3623,N_3590,N_3533);
nor U3624 (N_3624,N_3510,N_3598);
nor U3625 (N_3625,N_3528,N_3580);
xnor U3626 (N_3626,N_3524,N_3534);
nor U3627 (N_3627,N_3504,N_3565);
nor U3628 (N_3628,N_3502,N_3543);
nand U3629 (N_3629,N_3592,N_3586);
nor U3630 (N_3630,N_3526,N_3568);
nand U3631 (N_3631,N_3512,N_3561);
or U3632 (N_3632,N_3581,N_3552);
or U3633 (N_3633,N_3573,N_3594);
nand U3634 (N_3634,N_3544,N_3570);
nand U3635 (N_3635,N_3588,N_3550);
or U3636 (N_3636,N_3523,N_3527);
and U3637 (N_3637,N_3505,N_3596);
xnor U3638 (N_3638,N_3515,N_3520);
and U3639 (N_3639,N_3566,N_3560);
and U3640 (N_3640,N_3599,N_3508);
and U3641 (N_3641,N_3540,N_3522);
xor U3642 (N_3642,N_3509,N_3513);
xor U3643 (N_3643,N_3583,N_3587);
and U3644 (N_3644,N_3585,N_3531);
nor U3645 (N_3645,N_3571,N_3577);
nor U3646 (N_3646,N_3584,N_3536);
and U3647 (N_3647,N_3551,N_3556);
xnor U3648 (N_3648,N_3529,N_3557);
or U3649 (N_3649,N_3507,N_3519);
nor U3650 (N_3650,N_3512,N_3510);
nand U3651 (N_3651,N_3586,N_3534);
nor U3652 (N_3652,N_3559,N_3586);
nand U3653 (N_3653,N_3558,N_3531);
and U3654 (N_3654,N_3538,N_3508);
nor U3655 (N_3655,N_3591,N_3516);
or U3656 (N_3656,N_3529,N_3560);
or U3657 (N_3657,N_3554,N_3595);
nand U3658 (N_3658,N_3501,N_3571);
and U3659 (N_3659,N_3569,N_3577);
and U3660 (N_3660,N_3568,N_3560);
xnor U3661 (N_3661,N_3531,N_3518);
nand U3662 (N_3662,N_3557,N_3522);
nor U3663 (N_3663,N_3594,N_3521);
nor U3664 (N_3664,N_3501,N_3534);
or U3665 (N_3665,N_3518,N_3532);
nor U3666 (N_3666,N_3568,N_3501);
or U3667 (N_3667,N_3580,N_3578);
xor U3668 (N_3668,N_3545,N_3582);
nand U3669 (N_3669,N_3536,N_3503);
nand U3670 (N_3670,N_3569,N_3588);
nand U3671 (N_3671,N_3554,N_3597);
or U3672 (N_3672,N_3536,N_3569);
xor U3673 (N_3673,N_3506,N_3563);
nor U3674 (N_3674,N_3542,N_3596);
nand U3675 (N_3675,N_3543,N_3532);
nand U3676 (N_3676,N_3585,N_3552);
or U3677 (N_3677,N_3587,N_3596);
nand U3678 (N_3678,N_3545,N_3549);
nor U3679 (N_3679,N_3500,N_3538);
nand U3680 (N_3680,N_3576,N_3582);
or U3681 (N_3681,N_3517,N_3563);
nor U3682 (N_3682,N_3553,N_3529);
nor U3683 (N_3683,N_3572,N_3531);
nor U3684 (N_3684,N_3501,N_3523);
nand U3685 (N_3685,N_3533,N_3578);
or U3686 (N_3686,N_3572,N_3597);
or U3687 (N_3687,N_3583,N_3542);
nand U3688 (N_3688,N_3531,N_3539);
and U3689 (N_3689,N_3555,N_3502);
or U3690 (N_3690,N_3507,N_3538);
and U3691 (N_3691,N_3520,N_3577);
nor U3692 (N_3692,N_3553,N_3594);
nor U3693 (N_3693,N_3543,N_3511);
nand U3694 (N_3694,N_3540,N_3520);
or U3695 (N_3695,N_3579,N_3510);
nor U3696 (N_3696,N_3561,N_3595);
and U3697 (N_3697,N_3509,N_3516);
nor U3698 (N_3698,N_3570,N_3512);
nor U3699 (N_3699,N_3576,N_3599);
and U3700 (N_3700,N_3608,N_3649);
and U3701 (N_3701,N_3601,N_3692);
and U3702 (N_3702,N_3616,N_3687);
nand U3703 (N_3703,N_3621,N_3619);
and U3704 (N_3704,N_3664,N_3684);
or U3705 (N_3705,N_3622,N_3633);
and U3706 (N_3706,N_3665,N_3634);
nand U3707 (N_3707,N_3615,N_3606);
nor U3708 (N_3708,N_3632,N_3609);
or U3709 (N_3709,N_3623,N_3671);
and U3710 (N_3710,N_3625,N_3689);
or U3711 (N_3711,N_3658,N_3691);
xor U3712 (N_3712,N_3676,N_3631);
or U3713 (N_3713,N_3600,N_3611);
xor U3714 (N_3714,N_3636,N_3697);
and U3715 (N_3715,N_3640,N_3659);
or U3716 (N_3716,N_3618,N_3675);
nand U3717 (N_3717,N_3668,N_3639);
nor U3718 (N_3718,N_3602,N_3674);
xor U3719 (N_3719,N_3661,N_3655);
and U3720 (N_3720,N_3654,N_3620);
xnor U3721 (N_3721,N_3642,N_3647);
or U3722 (N_3722,N_3698,N_3688);
nand U3723 (N_3723,N_3613,N_3624);
nor U3724 (N_3724,N_3696,N_3604);
and U3725 (N_3725,N_3635,N_3651);
nor U3726 (N_3726,N_3680,N_3641);
xor U3727 (N_3727,N_3627,N_3669);
nor U3728 (N_3728,N_3667,N_3672);
nor U3729 (N_3729,N_3628,N_3677);
and U3730 (N_3730,N_3646,N_3656);
and U3731 (N_3731,N_3699,N_3614);
and U3732 (N_3732,N_3679,N_3630);
and U3733 (N_3733,N_3653,N_3607);
or U3734 (N_3734,N_3644,N_3693);
nor U3735 (N_3735,N_3648,N_3605);
nor U3736 (N_3736,N_3652,N_3637);
and U3737 (N_3737,N_3678,N_3662);
nor U3738 (N_3738,N_3682,N_3643);
and U3739 (N_3739,N_3638,N_3690);
nand U3740 (N_3740,N_3694,N_3612);
nor U3741 (N_3741,N_3670,N_3681);
or U3742 (N_3742,N_3610,N_3603);
and U3743 (N_3743,N_3645,N_3666);
nor U3744 (N_3744,N_3617,N_3695);
xor U3745 (N_3745,N_3685,N_3657);
nand U3746 (N_3746,N_3673,N_3683);
xor U3747 (N_3747,N_3686,N_3663);
nor U3748 (N_3748,N_3629,N_3660);
nand U3749 (N_3749,N_3626,N_3650);
nor U3750 (N_3750,N_3633,N_3639);
nand U3751 (N_3751,N_3694,N_3640);
nor U3752 (N_3752,N_3655,N_3615);
and U3753 (N_3753,N_3649,N_3617);
xnor U3754 (N_3754,N_3677,N_3616);
nand U3755 (N_3755,N_3626,N_3698);
nor U3756 (N_3756,N_3693,N_3607);
and U3757 (N_3757,N_3658,N_3652);
nor U3758 (N_3758,N_3673,N_3696);
nand U3759 (N_3759,N_3694,N_3692);
nand U3760 (N_3760,N_3668,N_3603);
nand U3761 (N_3761,N_3619,N_3633);
nor U3762 (N_3762,N_3638,N_3696);
xnor U3763 (N_3763,N_3650,N_3697);
nor U3764 (N_3764,N_3664,N_3608);
nand U3765 (N_3765,N_3610,N_3656);
nor U3766 (N_3766,N_3604,N_3641);
nand U3767 (N_3767,N_3605,N_3672);
xnor U3768 (N_3768,N_3612,N_3622);
nor U3769 (N_3769,N_3652,N_3668);
xor U3770 (N_3770,N_3601,N_3600);
nand U3771 (N_3771,N_3625,N_3653);
nand U3772 (N_3772,N_3672,N_3658);
and U3773 (N_3773,N_3627,N_3648);
and U3774 (N_3774,N_3675,N_3622);
or U3775 (N_3775,N_3696,N_3608);
nand U3776 (N_3776,N_3610,N_3637);
xor U3777 (N_3777,N_3623,N_3678);
or U3778 (N_3778,N_3676,N_3616);
and U3779 (N_3779,N_3698,N_3604);
or U3780 (N_3780,N_3648,N_3634);
xor U3781 (N_3781,N_3695,N_3675);
nor U3782 (N_3782,N_3684,N_3652);
nor U3783 (N_3783,N_3662,N_3620);
or U3784 (N_3784,N_3656,N_3654);
or U3785 (N_3785,N_3667,N_3676);
xnor U3786 (N_3786,N_3632,N_3649);
or U3787 (N_3787,N_3616,N_3699);
or U3788 (N_3788,N_3615,N_3693);
xor U3789 (N_3789,N_3618,N_3615);
or U3790 (N_3790,N_3632,N_3679);
xnor U3791 (N_3791,N_3640,N_3689);
or U3792 (N_3792,N_3621,N_3626);
or U3793 (N_3793,N_3624,N_3679);
and U3794 (N_3794,N_3630,N_3695);
and U3795 (N_3795,N_3612,N_3675);
or U3796 (N_3796,N_3673,N_3691);
nand U3797 (N_3797,N_3637,N_3683);
nand U3798 (N_3798,N_3655,N_3609);
and U3799 (N_3799,N_3604,N_3699);
xor U3800 (N_3800,N_3727,N_3778);
and U3801 (N_3801,N_3780,N_3720);
or U3802 (N_3802,N_3704,N_3744);
and U3803 (N_3803,N_3758,N_3734);
xnor U3804 (N_3804,N_3796,N_3769);
xor U3805 (N_3805,N_3791,N_3748);
and U3806 (N_3806,N_3740,N_3718);
or U3807 (N_3807,N_3787,N_3733);
nor U3808 (N_3808,N_3750,N_3725);
or U3809 (N_3809,N_3707,N_3770);
xor U3810 (N_3810,N_3731,N_3736);
nor U3811 (N_3811,N_3701,N_3766);
xnor U3812 (N_3812,N_3747,N_3783);
nand U3813 (N_3813,N_3705,N_3776);
xor U3814 (N_3814,N_3793,N_3739);
or U3815 (N_3815,N_3768,N_3772);
nand U3816 (N_3816,N_3774,N_3723);
nand U3817 (N_3817,N_3716,N_3700);
nor U3818 (N_3818,N_3710,N_3792);
nand U3819 (N_3819,N_3741,N_3798);
xor U3820 (N_3820,N_3724,N_3761);
and U3821 (N_3821,N_3737,N_3703);
or U3822 (N_3822,N_3773,N_3795);
nand U3823 (N_3823,N_3789,N_3762);
nor U3824 (N_3824,N_3786,N_3729);
and U3825 (N_3825,N_3749,N_3711);
nand U3826 (N_3826,N_3712,N_3730);
or U3827 (N_3827,N_3757,N_3781);
nand U3828 (N_3828,N_3760,N_3753);
nor U3829 (N_3829,N_3756,N_3775);
xnor U3830 (N_3830,N_3788,N_3759);
nor U3831 (N_3831,N_3794,N_3771);
xor U3832 (N_3832,N_3738,N_3722);
nand U3833 (N_3833,N_3728,N_3702);
nand U3834 (N_3834,N_3742,N_3714);
xor U3835 (N_3835,N_3752,N_3755);
or U3836 (N_3836,N_3745,N_3790);
nor U3837 (N_3837,N_3721,N_3764);
or U3838 (N_3838,N_3785,N_3719);
nand U3839 (N_3839,N_3706,N_3765);
nor U3840 (N_3840,N_3799,N_3746);
nor U3841 (N_3841,N_3743,N_3726);
nor U3842 (N_3842,N_3797,N_3713);
nor U3843 (N_3843,N_3717,N_3754);
nor U3844 (N_3844,N_3782,N_3732);
xor U3845 (N_3845,N_3709,N_3777);
and U3846 (N_3846,N_3715,N_3735);
nand U3847 (N_3847,N_3708,N_3779);
xor U3848 (N_3848,N_3767,N_3784);
nor U3849 (N_3849,N_3751,N_3763);
or U3850 (N_3850,N_3749,N_3714);
xnor U3851 (N_3851,N_3752,N_3772);
nor U3852 (N_3852,N_3708,N_3723);
or U3853 (N_3853,N_3785,N_3794);
and U3854 (N_3854,N_3777,N_3712);
or U3855 (N_3855,N_3785,N_3774);
or U3856 (N_3856,N_3745,N_3731);
or U3857 (N_3857,N_3795,N_3799);
nor U3858 (N_3858,N_3725,N_3757);
and U3859 (N_3859,N_3744,N_3769);
or U3860 (N_3860,N_3751,N_3705);
xor U3861 (N_3861,N_3711,N_3772);
nand U3862 (N_3862,N_3748,N_3777);
nor U3863 (N_3863,N_3724,N_3716);
or U3864 (N_3864,N_3741,N_3773);
nand U3865 (N_3865,N_3734,N_3783);
xor U3866 (N_3866,N_3770,N_3733);
and U3867 (N_3867,N_3735,N_3754);
or U3868 (N_3868,N_3788,N_3706);
or U3869 (N_3869,N_3746,N_3797);
nor U3870 (N_3870,N_3798,N_3711);
nor U3871 (N_3871,N_3769,N_3780);
or U3872 (N_3872,N_3772,N_3738);
xnor U3873 (N_3873,N_3771,N_3776);
nor U3874 (N_3874,N_3705,N_3777);
and U3875 (N_3875,N_3779,N_3712);
xnor U3876 (N_3876,N_3723,N_3750);
and U3877 (N_3877,N_3790,N_3737);
nor U3878 (N_3878,N_3748,N_3737);
xor U3879 (N_3879,N_3795,N_3763);
or U3880 (N_3880,N_3737,N_3741);
nor U3881 (N_3881,N_3723,N_3710);
nand U3882 (N_3882,N_3780,N_3781);
or U3883 (N_3883,N_3746,N_3756);
and U3884 (N_3884,N_3734,N_3722);
nand U3885 (N_3885,N_3789,N_3761);
nor U3886 (N_3886,N_3791,N_3764);
and U3887 (N_3887,N_3747,N_3725);
or U3888 (N_3888,N_3769,N_3773);
xnor U3889 (N_3889,N_3764,N_3734);
or U3890 (N_3890,N_3786,N_3751);
and U3891 (N_3891,N_3794,N_3717);
and U3892 (N_3892,N_3710,N_3713);
nand U3893 (N_3893,N_3764,N_3746);
nor U3894 (N_3894,N_3721,N_3765);
and U3895 (N_3895,N_3705,N_3782);
and U3896 (N_3896,N_3797,N_3751);
nand U3897 (N_3897,N_3778,N_3770);
and U3898 (N_3898,N_3748,N_3710);
and U3899 (N_3899,N_3795,N_3740);
and U3900 (N_3900,N_3800,N_3812);
or U3901 (N_3901,N_3802,N_3827);
nand U3902 (N_3902,N_3840,N_3806);
and U3903 (N_3903,N_3869,N_3810);
nor U3904 (N_3904,N_3871,N_3804);
or U3905 (N_3905,N_3895,N_3899);
xor U3906 (N_3906,N_3876,N_3852);
xnor U3907 (N_3907,N_3874,N_3809);
nand U3908 (N_3908,N_3862,N_3811);
nor U3909 (N_3909,N_3822,N_3838);
xnor U3910 (N_3910,N_3868,N_3865);
xnor U3911 (N_3911,N_3855,N_3867);
nand U3912 (N_3912,N_3864,N_3891);
and U3913 (N_3913,N_3887,N_3828);
xnor U3914 (N_3914,N_3878,N_3858);
and U3915 (N_3915,N_3859,N_3815);
or U3916 (N_3916,N_3884,N_3879);
nor U3917 (N_3917,N_3814,N_3816);
nor U3918 (N_3918,N_3847,N_3854);
nor U3919 (N_3919,N_3842,N_3801);
xnor U3920 (N_3920,N_3863,N_3888);
xor U3921 (N_3921,N_3830,N_3819);
and U3922 (N_3922,N_3818,N_3832);
xor U3923 (N_3923,N_3889,N_3896);
nand U3924 (N_3924,N_3848,N_3875);
nor U3925 (N_3925,N_3831,N_3870);
nand U3926 (N_3926,N_3860,N_3856);
xor U3927 (N_3927,N_3866,N_3883);
nand U3928 (N_3928,N_3861,N_3820);
or U3929 (N_3929,N_3833,N_3873);
xnor U3930 (N_3930,N_3823,N_3890);
and U3931 (N_3931,N_3826,N_3829);
nor U3932 (N_3932,N_3813,N_3844);
nand U3933 (N_3933,N_3845,N_3803);
nand U3934 (N_3934,N_3851,N_3825);
xor U3935 (N_3935,N_3805,N_3893);
or U3936 (N_3936,N_3880,N_3872);
nand U3937 (N_3937,N_3817,N_3824);
xor U3938 (N_3938,N_3839,N_3897);
and U3939 (N_3939,N_3841,N_3877);
xnor U3940 (N_3940,N_3821,N_3886);
and U3941 (N_3941,N_3892,N_3834);
and U3942 (N_3942,N_3885,N_3850);
nor U3943 (N_3943,N_3881,N_3846);
nand U3944 (N_3944,N_3882,N_3853);
and U3945 (N_3945,N_3837,N_3849);
nand U3946 (N_3946,N_3857,N_3836);
or U3947 (N_3947,N_3843,N_3808);
nor U3948 (N_3948,N_3807,N_3898);
nor U3949 (N_3949,N_3894,N_3835);
or U3950 (N_3950,N_3881,N_3820);
and U3951 (N_3951,N_3824,N_3809);
nand U3952 (N_3952,N_3817,N_3890);
xnor U3953 (N_3953,N_3888,N_3875);
and U3954 (N_3954,N_3866,N_3897);
and U3955 (N_3955,N_3867,N_3825);
nand U3956 (N_3956,N_3819,N_3894);
xnor U3957 (N_3957,N_3808,N_3823);
and U3958 (N_3958,N_3812,N_3821);
xnor U3959 (N_3959,N_3835,N_3871);
nand U3960 (N_3960,N_3817,N_3809);
nand U3961 (N_3961,N_3833,N_3804);
nand U3962 (N_3962,N_3838,N_3850);
xnor U3963 (N_3963,N_3839,N_3828);
nand U3964 (N_3964,N_3859,N_3812);
or U3965 (N_3965,N_3887,N_3867);
nand U3966 (N_3966,N_3895,N_3866);
or U3967 (N_3967,N_3825,N_3817);
nor U3968 (N_3968,N_3887,N_3859);
and U3969 (N_3969,N_3803,N_3872);
xor U3970 (N_3970,N_3872,N_3866);
and U3971 (N_3971,N_3885,N_3866);
nand U3972 (N_3972,N_3843,N_3837);
xor U3973 (N_3973,N_3851,N_3890);
nand U3974 (N_3974,N_3825,N_3811);
nand U3975 (N_3975,N_3896,N_3867);
nor U3976 (N_3976,N_3872,N_3870);
nand U3977 (N_3977,N_3811,N_3831);
xnor U3978 (N_3978,N_3863,N_3885);
nand U3979 (N_3979,N_3842,N_3814);
and U3980 (N_3980,N_3857,N_3806);
nand U3981 (N_3981,N_3890,N_3809);
xor U3982 (N_3982,N_3800,N_3852);
nor U3983 (N_3983,N_3826,N_3887);
or U3984 (N_3984,N_3862,N_3850);
nand U3985 (N_3985,N_3865,N_3857);
nand U3986 (N_3986,N_3838,N_3896);
nor U3987 (N_3987,N_3820,N_3811);
xor U3988 (N_3988,N_3878,N_3845);
and U3989 (N_3989,N_3862,N_3837);
and U3990 (N_3990,N_3888,N_3821);
and U3991 (N_3991,N_3844,N_3896);
and U3992 (N_3992,N_3883,N_3884);
nor U3993 (N_3993,N_3889,N_3865);
or U3994 (N_3994,N_3811,N_3875);
xor U3995 (N_3995,N_3867,N_3826);
and U3996 (N_3996,N_3840,N_3827);
xnor U3997 (N_3997,N_3816,N_3870);
xnor U3998 (N_3998,N_3857,N_3845);
or U3999 (N_3999,N_3850,N_3821);
or U4000 (N_4000,N_3906,N_3991);
or U4001 (N_4001,N_3984,N_3912);
xnor U4002 (N_4002,N_3986,N_3908);
xnor U4003 (N_4003,N_3970,N_3947);
or U4004 (N_4004,N_3921,N_3989);
and U4005 (N_4005,N_3954,N_3976);
nand U4006 (N_4006,N_3928,N_3969);
and U4007 (N_4007,N_3958,N_3946);
or U4008 (N_4008,N_3927,N_3940);
nand U4009 (N_4009,N_3961,N_3933);
and U4010 (N_4010,N_3965,N_3994);
nor U4011 (N_4011,N_3949,N_3997);
nor U4012 (N_4012,N_3992,N_3981);
or U4013 (N_4013,N_3964,N_3996);
nand U4014 (N_4014,N_3934,N_3952);
and U4015 (N_4015,N_3944,N_3995);
nor U4016 (N_4016,N_3902,N_3972);
and U4017 (N_4017,N_3963,N_3936);
nor U4018 (N_4018,N_3978,N_3983);
and U4019 (N_4019,N_3929,N_3990);
and U4020 (N_4020,N_3915,N_3962);
nor U4021 (N_4021,N_3911,N_3913);
nand U4022 (N_4022,N_3926,N_3980);
xor U4023 (N_4023,N_3907,N_3901);
and U4024 (N_4024,N_3960,N_3903);
xnor U4025 (N_4025,N_3959,N_3945);
nor U4026 (N_4026,N_3937,N_3932);
or U4027 (N_4027,N_3920,N_3993);
and U4028 (N_4028,N_3971,N_3974);
and U4029 (N_4029,N_3924,N_3966);
or U4030 (N_4030,N_3975,N_3919);
nand U4031 (N_4031,N_3987,N_3998);
xnor U4032 (N_4032,N_3951,N_3982);
xnor U4033 (N_4033,N_3985,N_3948);
or U4034 (N_4034,N_3988,N_3904);
xor U4035 (N_4035,N_3938,N_3909);
or U4036 (N_4036,N_3923,N_3941);
or U4037 (N_4037,N_3916,N_3905);
nor U4038 (N_4038,N_3968,N_3943);
xor U4039 (N_4039,N_3957,N_3953);
nand U4040 (N_4040,N_3935,N_3900);
nor U4041 (N_4041,N_3918,N_3955);
and U4042 (N_4042,N_3917,N_3973);
nand U4043 (N_4043,N_3942,N_3931);
nand U4044 (N_4044,N_3956,N_3979);
or U4045 (N_4045,N_3925,N_3939);
nor U4046 (N_4046,N_3910,N_3999);
xor U4047 (N_4047,N_3950,N_3914);
or U4048 (N_4048,N_3977,N_3930);
nand U4049 (N_4049,N_3922,N_3967);
and U4050 (N_4050,N_3961,N_3992);
and U4051 (N_4051,N_3976,N_3905);
or U4052 (N_4052,N_3943,N_3932);
or U4053 (N_4053,N_3925,N_3943);
xnor U4054 (N_4054,N_3911,N_3996);
or U4055 (N_4055,N_3967,N_3933);
nand U4056 (N_4056,N_3948,N_3910);
nor U4057 (N_4057,N_3978,N_3931);
and U4058 (N_4058,N_3911,N_3901);
and U4059 (N_4059,N_3954,N_3909);
or U4060 (N_4060,N_3963,N_3935);
and U4061 (N_4061,N_3991,N_3956);
nand U4062 (N_4062,N_3948,N_3958);
or U4063 (N_4063,N_3936,N_3923);
or U4064 (N_4064,N_3956,N_3910);
and U4065 (N_4065,N_3935,N_3981);
xor U4066 (N_4066,N_3941,N_3961);
xnor U4067 (N_4067,N_3977,N_3955);
nor U4068 (N_4068,N_3909,N_3929);
xnor U4069 (N_4069,N_3964,N_3927);
nand U4070 (N_4070,N_3923,N_3950);
nand U4071 (N_4071,N_3932,N_3954);
nor U4072 (N_4072,N_3911,N_3937);
and U4073 (N_4073,N_3936,N_3997);
and U4074 (N_4074,N_3901,N_3950);
and U4075 (N_4075,N_3987,N_3984);
nand U4076 (N_4076,N_3945,N_3955);
and U4077 (N_4077,N_3949,N_3909);
or U4078 (N_4078,N_3902,N_3955);
nand U4079 (N_4079,N_3917,N_3948);
nand U4080 (N_4080,N_3910,N_3922);
nor U4081 (N_4081,N_3963,N_3965);
xor U4082 (N_4082,N_3937,N_3933);
nor U4083 (N_4083,N_3937,N_3962);
xor U4084 (N_4084,N_3923,N_3900);
xor U4085 (N_4085,N_3936,N_3916);
xnor U4086 (N_4086,N_3907,N_3934);
nor U4087 (N_4087,N_3925,N_3996);
and U4088 (N_4088,N_3956,N_3948);
xnor U4089 (N_4089,N_3962,N_3925);
nand U4090 (N_4090,N_3971,N_3920);
xnor U4091 (N_4091,N_3950,N_3933);
nand U4092 (N_4092,N_3943,N_3991);
and U4093 (N_4093,N_3908,N_3956);
and U4094 (N_4094,N_3921,N_3903);
or U4095 (N_4095,N_3912,N_3928);
nor U4096 (N_4096,N_3928,N_3940);
nor U4097 (N_4097,N_3981,N_3948);
and U4098 (N_4098,N_3973,N_3957);
or U4099 (N_4099,N_3921,N_3996);
or U4100 (N_4100,N_4089,N_4042);
or U4101 (N_4101,N_4055,N_4007);
nor U4102 (N_4102,N_4014,N_4020);
and U4103 (N_4103,N_4053,N_4091);
nor U4104 (N_4104,N_4029,N_4021);
nand U4105 (N_4105,N_4035,N_4012);
or U4106 (N_4106,N_4018,N_4058);
xor U4107 (N_4107,N_4071,N_4025);
or U4108 (N_4108,N_4050,N_4087);
or U4109 (N_4109,N_4019,N_4028);
xnor U4110 (N_4110,N_4097,N_4000);
nor U4111 (N_4111,N_4092,N_4076);
xor U4112 (N_4112,N_4057,N_4033);
and U4113 (N_4113,N_4099,N_4088);
or U4114 (N_4114,N_4095,N_4067);
nor U4115 (N_4115,N_4036,N_4090);
or U4116 (N_4116,N_4054,N_4061);
nand U4117 (N_4117,N_4068,N_4082);
nor U4118 (N_4118,N_4073,N_4046);
nor U4119 (N_4119,N_4017,N_4009);
and U4120 (N_4120,N_4049,N_4085);
and U4121 (N_4121,N_4056,N_4063);
and U4122 (N_4122,N_4043,N_4031);
xor U4123 (N_4123,N_4022,N_4081);
nand U4124 (N_4124,N_4030,N_4048);
xor U4125 (N_4125,N_4002,N_4010);
nand U4126 (N_4126,N_4004,N_4069);
nand U4127 (N_4127,N_4038,N_4086);
nand U4128 (N_4128,N_4006,N_4079);
or U4129 (N_4129,N_4005,N_4051);
nor U4130 (N_4130,N_4066,N_4074);
and U4131 (N_4131,N_4045,N_4084);
xor U4132 (N_4132,N_4072,N_4052);
nand U4133 (N_4133,N_4041,N_4040);
and U4134 (N_4134,N_4093,N_4078);
nor U4135 (N_4135,N_4013,N_4096);
or U4136 (N_4136,N_4011,N_4016);
xor U4137 (N_4137,N_4037,N_4015);
xor U4138 (N_4138,N_4039,N_4023);
nand U4139 (N_4139,N_4064,N_4032);
nand U4140 (N_4140,N_4077,N_4094);
and U4141 (N_4141,N_4062,N_4059);
xnor U4142 (N_4142,N_4001,N_4060);
and U4143 (N_4143,N_4080,N_4027);
or U4144 (N_4144,N_4034,N_4026);
or U4145 (N_4145,N_4008,N_4098);
and U4146 (N_4146,N_4075,N_4003);
and U4147 (N_4147,N_4070,N_4065);
nand U4148 (N_4148,N_4047,N_4044);
nor U4149 (N_4149,N_4083,N_4024);
nand U4150 (N_4150,N_4008,N_4060);
and U4151 (N_4151,N_4031,N_4098);
nor U4152 (N_4152,N_4027,N_4090);
or U4153 (N_4153,N_4028,N_4054);
and U4154 (N_4154,N_4021,N_4070);
or U4155 (N_4155,N_4023,N_4009);
nand U4156 (N_4156,N_4049,N_4069);
xor U4157 (N_4157,N_4036,N_4023);
and U4158 (N_4158,N_4071,N_4091);
nor U4159 (N_4159,N_4012,N_4092);
nand U4160 (N_4160,N_4082,N_4065);
xor U4161 (N_4161,N_4041,N_4037);
nand U4162 (N_4162,N_4076,N_4089);
nand U4163 (N_4163,N_4028,N_4058);
xor U4164 (N_4164,N_4047,N_4039);
xnor U4165 (N_4165,N_4087,N_4038);
nand U4166 (N_4166,N_4076,N_4042);
or U4167 (N_4167,N_4061,N_4007);
nor U4168 (N_4168,N_4069,N_4089);
nand U4169 (N_4169,N_4096,N_4060);
nor U4170 (N_4170,N_4021,N_4094);
nor U4171 (N_4171,N_4035,N_4033);
and U4172 (N_4172,N_4032,N_4043);
nand U4173 (N_4173,N_4033,N_4056);
and U4174 (N_4174,N_4079,N_4097);
nor U4175 (N_4175,N_4029,N_4005);
nand U4176 (N_4176,N_4038,N_4097);
and U4177 (N_4177,N_4080,N_4009);
xnor U4178 (N_4178,N_4009,N_4054);
nor U4179 (N_4179,N_4015,N_4066);
nand U4180 (N_4180,N_4013,N_4030);
nand U4181 (N_4181,N_4034,N_4027);
nor U4182 (N_4182,N_4054,N_4005);
xnor U4183 (N_4183,N_4012,N_4077);
and U4184 (N_4184,N_4063,N_4024);
or U4185 (N_4185,N_4018,N_4009);
and U4186 (N_4186,N_4011,N_4059);
nor U4187 (N_4187,N_4072,N_4095);
nor U4188 (N_4188,N_4044,N_4061);
nand U4189 (N_4189,N_4013,N_4051);
nand U4190 (N_4190,N_4079,N_4048);
or U4191 (N_4191,N_4034,N_4006);
and U4192 (N_4192,N_4063,N_4009);
nand U4193 (N_4193,N_4081,N_4093);
nor U4194 (N_4194,N_4005,N_4079);
or U4195 (N_4195,N_4012,N_4009);
and U4196 (N_4196,N_4002,N_4042);
nand U4197 (N_4197,N_4024,N_4050);
nor U4198 (N_4198,N_4049,N_4024);
and U4199 (N_4199,N_4093,N_4056);
nand U4200 (N_4200,N_4145,N_4158);
or U4201 (N_4201,N_4194,N_4159);
and U4202 (N_4202,N_4146,N_4168);
and U4203 (N_4203,N_4143,N_4155);
and U4204 (N_4204,N_4142,N_4189);
xnor U4205 (N_4205,N_4196,N_4154);
and U4206 (N_4206,N_4153,N_4170);
xor U4207 (N_4207,N_4130,N_4149);
xor U4208 (N_4208,N_4115,N_4123);
and U4209 (N_4209,N_4114,N_4167);
nand U4210 (N_4210,N_4144,N_4160);
xor U4211 (N_4211,N_4103,N_4122);
or U4212 (N_4212,N_4151,N_4131);
and U4213 (N_4213,N_4129,N_4173);
or U4214 (N_4214,N_4148,N_4110);
nor U4215 (N_4215,N_4125,N_4135);
nor U4216 (N_4216,N_4185,N_4166);
and U4217 (N_4217,N_4126,N_4139);
and U4218 (N_4218,N_4165,N_4152);
xor U4219 (N_4219,N_4141,N_4133);
nand U4220 (N_4220,N_4118,N_4175);
and U4221 (N_4221,N_4140,N_4198);
xor U4222 (N_4222,N_4162,N_4182);
nand U4223 (N_4223,N_4187,N_4107);
xnor U4224 (N_4224,N_4104,N_4179);
nand U4225 (N_4225,N_4119,N_4184);
and U4226 (N_4226,N_4183,N_4164);
nor U4227 (N_4227,N_4188,N_4134);
or U4228 (N_4228,N_4120,N_4181);
nor U4229 (N_4229,N_4156,N_4136);
nand U4230 (N_4230,N_4127,N_4171);
xnor U4231 (N_4231,N_4116,N_4147);
nand U4232 (N_4232,N_4112,N_4186);
nor U4233 (N_4233,N_4111,N_4161);
and U4234 (N_4234,N_4193,N_4105);
or U4235 (N_4235,N_4197,N_4113);
nor U4236 (N_4236,N_4121,N_4157);
xnor U4237 (N_4237,N_4128,N_4192);
and U4238 (N_4238,N_4132,N_4169);
nor U4239 (N_4239,N_4172,N_4180);
nor U4240 (N_4240,N_4150,N_4124);
or U4241 (N_4241,N_4137,N_4191);
nor U4242 (N_4242,N_4100,N_4199);
and U4243 (N_4243,N_4101,N_4178);
or U4244 (N_4244,N_4117,N_4176);
or U4245 (N_4245,N_4190,N_4138);
nor U4246 (N_4246,N_4108,N_4177);
and U4247 (N_4247,N_4174,N_4106);
nor U4248 (N_4248,N_4102,N_4195);
and U4249 (N_4249,N_4163,N_4109);
or U4250 (N_4250,N_4162,N_4166);
and U4251 (N_4251,N_4121,N_4113);
or U4252 (N_4252,N_4147,N_4118);
or U4253 (N_4253,N_4117,N_4127);
or U4254 (N_4254,N_4151,N_4178);
xnor U4255 (N_4255,N_4170,N_4194);
nand U4256 (N_4256,N_4181,N_4143);
nor U4257 (N_4257,N_4161,N_4171);
nor U4258 (N_4258,N_4115,N_4135);
and U4259 (N_4259,N_4178,N_4185);
nor U4260 (N_4260,N_4136,N_4133);
nand U4261 (N_4261,N_4136,N_4143);
nor U4262 (N_4262,N_4157,N_4183);
xor U4263 (N_4263,N_4172,N_4129);
or U4264 (N_4264,N_4179,N_4164);
nand U4265 (N_4265,N_4195,N_4193);
nor U4266 (N_4266,N_4163,N_4158);
nand U4267 (N_4267,N_4139,N_4172);
nor U4268 (N_4268,N_4118,N_4190);
xor U4269 (N_4269,N_4161,N_4178);
nand U4270 (N_4270,N_4110,N_4125);
or U4271 (N_4271,N_4147,N_4194);
nor U4272 (N_4272,N_4173,N_4175);
or U4273 (N_4273,N_4180,N_4106);
xnor U4274 (N_4274,N_4151,N_4171);
nand U4275 (N_4275,N_4181,N_4161);
or U4276 (N_4276,N_4150,N_4181);
or U4277 (N_4277,N_4155,N_4183);
or U4278 (N_4278,N_4120,N_4132);
nor U4279 (N_4279,N_4147,N_4120);
and U4280 (N_4280,N_4159,N_4141);
nand U4281 (N_4281,N_4111,N_4107);
nor U4282 (N_4282,N_4189,N_4111);
xnor U4283 (N_4283,N_4173,N_4152);
nand U4284 (N_4284,N_4117,N_4129);
nand U4285 (N_4285,N_4197,N_4178);
nand U4286 (N_4286,N_4168,N_4186);
and U4287 (N_4287,N_4147,N_4188);
nor U4288 (N_4288,N_4180,N_4133);
nor U4289 (N_4289,N_4167,N_4107);
or U4290 (N_4290,N_4183,N_4127);
nor U4291 (N_4291,N_4163,N_4179);
or U4292 (N_4292,N_4151,N_4176);
xor U4293 (N_4293,N_4121,N_4108);
and U4294 (N_4294,N_4167,N_4148);
nand U4295 (N_4295,N_4139,N_4135);
xor U4296 (N_4296,N_4172,N_4186);
nor U4297 (N_4297,N_4101,N_4166);
xnor U4298 (N_4298,N_4170,N_4197);
or U4299 (N_4299,N_4156,N_4160);
nor U4300 (N_4300,N_4234,N_4258);
or U4301 (N_4301,N_4205,N_4208);
nand U4302 (N_4302,N_4231,N_4276);
nand U4303 (N_4303,N_4275,N_4272);
or U4304 (N_4304,N_4222,N_4219);
nor U4305 (N_4305,N_4221,N_4257);
nand U4306 (N_4306,N_4228,N_4287);
nor U4307 (N_4307,N_4255,N_4215);
xor U4308 (N_4308,N_4271,N_4212);
xnor U4309 (N_4309,N_4295,N_4264);
or U4310 (N_4310,N_4296,N_4236);
nor U4311 (N_4311,N_4243,N_4278);
nor U4312 (N_4312,N_4297,N_4210);
or U4313 (N_4313,N_4263,N_4245);
nor U4314 (N_4314,N_4277,N_4229);
nand U4315 (N_4315,N_4273,N_4202);
nor U4316 (N_4316,N_4200,N_4290);
xor U4317 (N_4317,N_4281,N_4265);
nor U4318 (N_4318,N_4279,N_4254);
and U4319 (N_4319,N_4294,N_4248);
xnor U4320 (N_4320,N_4220,N_4267);
or U4321 (N_4321,N_4209,N_4230);
nor U4322 (N_4322,N_4237,N_4283);
nor U4323 (N_4323,N_4206,N_4225);
and U4324 (N_4324,N_4211,N_4201);
or U4325 (N_4325,N_4288,N_4232);
nand U4326 (N_4326,N_4242,N_4266);
nand U4327 (N_4327,N_4285,N_4216);
nand U4328 (N_4328,N_4252,N_4233);
nor U4329 (N_4329,N_4213,N_4269);
and U4330 (N_4330,N_4284,N_4280);
or U4331 (N_4331,N_4289,N_4253);
nand U4332 (N_4332,N_4214,N_4238);
nor U4333 (N_4333,N_4207,N_4217);
or U4334 (N_4334,N_4223,N_4259);
and U4335 (N_4335,N_4251,N_4299);
nand U4336 (N_4336,N_4291,N_4282);
nand U4337 (N_4337,N_4203,N_4226);
nand U4338 (N_4338,N_4241,N_4224);
or U4339 (N_4339,N_4247,N_4204);
and U4340 (N_4340,N_4240,N_4286);
nand U4341 (N_4341,N_4292,N_4227);
nand U4342 (N_4342,N_4260,N_4235);
nor U4343 (N_4343,N_4250,N_4274);
and U4344 (N_4344,N_4268,N_4218);
xnor U4345 (N_4345,N_4261,N_4262);
nand U4346 (N_4346,N_4293,N_4298);
or U4347 (N_4347,N_4239,N_4246);
and U4348 (N_4348,N_4249,N_4244);
and U4349 (N_4349,N_4270,N_4256);
or U4350 (N_4350,N_4211,N_4229);
nand U4351 (N_4351,N_4258,N_4213);
and U4352 (N_4352,N_4250,N_4217);
and U4353 (N_4353,N_4240,N_4210);
nand U4354 (N_4354,N_4238,N_4222);
and U4355 (N_4355,N_4271,N_4209);
nand U4356 (N_4356,N_4295,N_4254);
nand U4357 (N_4357,N_4283,N_4215);
and U4358 (N_4358,N_4262,N_4289);
and U4359 (N_4359,N_4290,N_4259);
xnor U4360 (N_4360,N_4229,N_4200);
or U4361 (N_4361,N_4211,N_4287);
xnor U4362 (N_4362,N_4200,N_4253);
nand U4363 (N_4363,N_4248,N_4204);
or U4364 (N_4364,N_4226,N_4253);
nand U4365 (N_4365,N_4244,N_4236);
or U4366 (N_4366,N_4275,N_4230);
and U4367 (N_4367,N_4236,N_4285);
xor U4368 (N_4368,N_4226,N_4263);
or U4369 (N_4369,N_4266,N_4260);
or U4370 (N_4370,N_4211,N_4235);
nand U4371 (N_4371,N_4253,N_4268);
and U4372 (N_4372,N_4286,N_4202);
nand U4373 (N_4373,N_4286,N_4291);
or U4374 (N_4374,N_4220,N_4216);
and U4375 (N_4375,N_4228,N_4210);
and U4376 (N_4376,N_4286,N_4293);
or U4377 (N_4377,N_4272,N_4247);
nand U4378 (N_4378,N_4244,N_4222);
and U4379 (N_4379,N_4264,N_4244);
and U4380 (N_4380,N_4237,N_4248);
and U4381 (N_4381,N_4235,N_4213);
or U4382 (N_4382,N_4205,N_4206);
nand U4383 (N_4383,N_4209,N_4270);
or U4384 (N_4384,N_4259,N_4264);
or U4385 (N_4385,N_4225,N_4286);
or U4386 (N_4386,N_4275,N_4214);
nor U4387 (N_4387,N_4221,N_4265);
nand U4388 (N_4388,N_4244,N_4240);
xnor U4389 (N_4389,N_4251,N_4252);
or U4390 (N_4390,N_4285,N_4281);
nand U4391 (N_4391,N_4268,N_4271);
or U4392 (N_4392,N_4277,N_4267);
xor U4393 (N_4393,N_4256,N_4253);
xnor U4394 (N_4394,N_4244,N_4225);
and U4395 (N_4395,N_4247,N_4200);
nor U4396 (N_4396,N_4222,N_4255);
or U4397 (N_4397,N_4255,N_4245);
and U4398 (N_4398,N_4280,N_4204);
nand U4399 (N_4399,N_4211,N_4228);
xnor U4400 (N_4400,N_4332,N_4369);
or U4401 (N_4401,N_4321,N_4316);
xnor U4402 (N_4402,N_4356,N_4361);
nor U4403 (N_4403,N_4396,N_4343);
and U4404 (N_4404,N_4354,N_4308);
or U4405 (N_4405,N_4390,N_4309);
and U4406 (N_4406,N_4323,N_4364);
nand U4407 (N_4407,N_4315,N_4345);
xnor U4408 (N_4408,N_4312,N_4398);
xnor U4409 (N_4409,N_4357,N_4300);
nor U4410 (N_4410,N_4381,N_4338);
xnor U4411 (N_4411,N_4392,N_4346);
nand U4412 (N_4412,N_4348,N_4342);
or U4413 (N_4413,N_4333,N_4305);
xnor U4414 (N_4414,N_4336,N_4386);
or U4415 (N_4415,N_4344,N_4370);
xor U4416 (N_4416,N_4314,N_4399);
xor U4417 (N_4417,N_4382,N_4310);
or U4418 (N_4418,N_4331,N_4341);
nor U4419 (N_4419,N_4365,N_4384);
nand U4420 (N_4420,N_4380,N_4363);
and U4421 (N_4421,N_4330,N_4347);
nor U4422 (N_4422,N_4368,N_4349);
nand U4423 (N_4423,N_4371,N_4327);
or U4424 (N_4424,N_4350,N_4329);
nand U4425 (N_4425,N_4302,N_4358);
and U4426 (N_4426,N_4360,N_4374);
or U4427 (N_4427,N_4367,N_4393);
nand U4428 (N_4428,N_4324,N_4387);
nand U4429 (N_4429,N_4352,N_4394);
nor U4430 (N_4430,N_4307,N_4376);
nand U4431 (N_4431,N_4355,N_4397);
xor U4432 (N_4432,N_4334,N_4366);
xnor U4433 (N_4433,N_4351,N_4301);
or U4434 (N_4434,N_4317,N_4306);
and U4435 (N_4435,N_4389,N_4303);
and U4436 (N_4436,N_4337,N_4362);
xor U4437 (N_4437,N_4304,N_4377);
and U4438 (N_4438,N_4328,N_4325);
xnor U4439 (N_4439,N_4385,N_4359);
nand U4440 (N_4440,N_4391,N_4372);
or U4441 (N_4441,N_4339,N_4318);
or U4442 (N_4442,N_4373,N_4378);
xor U4443 (N_4443,N_4311,N_4319);
and U4444 (N_4444,N_4320,N_4383);
nor U4445 (N_4445,N_4313,N_4322);
nand U4446 (N_4446,N_4395,N_4335);
nor U4447 (N_4447,N_4326,N_4340);
nand U4448 (N_4448,N_4353,N_4379);
xnor U4449 (N_4449,N_4388,N_4375);
nand U4450 (N_4450,N_4391,N_4358);
and U4451 (N_4451,N_4361,N_4350);
or U4452 (N_4452,N_4331,N_4387);
and U4453 (N_4453,N_4396,N_4311);
xor U4454 (N_4454,N_4379,N_4347);
and U4455 (N_4455,N_4347,N_4332);
nand U4456 (N_4456,N_4341,N_4384);
or U4457 (N_4457,N_4371,N_4343);
or U4458 (N_4458,N_4390,N_4365);
nor U4459 (N_4459,N_4338,N_4371);
nor U4460 (N_4460,N_4312,N_4355);
xor U4461 (N_4461,N_4341,N_4314);
xor U4462 (N_4462,N_4317,N_4304);
xnor U4463 (N_4463,N_4339,N_4345);
or U4464 (N_4464,N_4344,N_4313);
and U4465 (N_4465,N_4301,N_4329);
or U4466 (N_4466,N_4399,N_4305);
nor U4467 (N_4467,N_4366,N_4308);
or U4468 (N_4468,N_4389,N_4350);
or U4469 (N_4469,N_4335,N_4329);
xor U4470 (N_4470,N_4361,N_4306);
nor U4471 (N_4471,N_4319,N_4348);
and U4472 (N_4472,N_4308,N_4320);
nor U4473 (N_4473,N_4316,N_4389);
or U4474 (N_4474,N_4397,N_4396);
nor U4475 (N_4475,N_4304,N_4399);
xor U4476 (N_4476,N_4375,N_4380);
nand U4477 (N_4477,N_4369,N_4338);
xor U4478 (N_4478,N_4387,N_4385);
nor U4479 (N_4479,N_4338,N_4393);
nand U4480 (N_4480,N_4358,N_4340);
or U4481 (N_4481,N_4354,N_4383);
or U4482 (N_4482,N_4319,N_4364);
nor U4483 (N_4483,N_4317,N_4341);
nand U4484 (N_4484,N_4365,N_4369);
nor U4485 (N_4485,N_4363,N_4311);
xnor U4486 (N_4486,N_4390,N_4338);
or U4487 (N_4487,N_4359,N_4331);
or U4488 (N_4488,N_4312,N_4359);
xnor U4489 (N_4489,N_4303,N_4336);
and U4490 (N_4490,N_4365,N_4353);
or U4491 (N_4491,N_4327,N_4360);
and U4492 (N_4492,N_4375,N_4383);
or U4493 (N_4493,N_4303,N_4381);
xor U4494 (N_4494,N_4312,N_4336);
nand U4495 (N_4495,N_4389,N_4358);
or U4496 (N_4496,N_4341,N_4385);
xnor U4497 (N_4497,N_4314,N_4323);
nand U4498 (N_4498,N_4352,N_4301);
nand U4499 (N_4499,N_4311,N_4398);
nand U4500 (N_4500,N_4457,N_4491);
nor U4501 (N_4501,N_4419,N_4415);
and U4502 (N_4502,N_4452,N_4404);
nand U4503 (N_4503,N_4406,N_4474);
and U4504 (N_4504,N_4401,N_4447);
and U4505 (N_4505,N_4418,N_4466);
nor U4506 (N_4506,N_4482,N_4496);
and U4507 (N_4507,N_4484,N_4473);
xor U4508 (N_4508,N_4463,N_4437);
nor U4509 (N_4509,N_4460,N_4451);
nand U4510 (N_4510,N_4449,N_4443);
xnor U4511 (N_4511,N_4445,N_4487);
nand U4512 (N_4512,N_4462,N_4407);
nand U4513 (N_4513,N_4420,N_4476);
xnor U4514 (N_4514,N_4475,N_4428);
xor U4515 (N_4515,N_4446,N_4412);
nor U4516 (N_4516,N_4433,N_4467);
and U4517 (N_4517,N_4417,N_4441);
nand U4518 (N_4518,N_4480,N_4471);
nand U4519 (N_4519,N_4490,N_4450);
nor U4520 (N_4520,N_4425,N_4436);
xnor U4521 (N_4521,N_4493,N_4416);
and U4522 (N_4522,N_4400,N_4421);
and U4523 (N_4523,N_4444,N_4461);
or U4524 (N_4524,N_4477,N_4488);
xor U4525 (N_4525,N_4494,N_4483);
or U4526 (N_4526,N_4434,N_4495);
xnor U4527 (N_4527,N_4486,N_4429);
and U4528 (N_4528,N_4465,N_4498);
nor U4529 (N_4529,N_4424,N_4478);
xnor U4530 (N_4530,N_4472,N_4497);
nand U4531 (N_4531,N_4402,N_4459);
xnor U4532 (N_4532,N_4479,N_4439);
nand U4533 (N_4533,N_4403,N_4448);
nand U4534 (N_4534,N_4454,N_4431);
xor U4535 (N_4535,N_4435,N_4458);
xor U4536 (N_4536,N_4468,N_4469);
or U4537 (N_4537,N_4422,N_4411);
nand U4538 (N_4538,N_4499,N_4423);
nand U4539 (N_4539,N_4408,N_4464);
xnor U4540 (N_4540,N_4427,N_4432);
and U4541 (N_4541,N_4442,N_4405);
nor U4542 (N_4542,N_4489,N_4453);
or U4543 (N_4543,N_4438,N_4409);
or U4544 (N_4544,N_4492,N_4455);
nor U4545 (N_4545,N_4430,N_4470);
or U4546 (N_4546,N_4410,N_4456);
xnor U4547 (N_4547,N_4426,N_4440);
and U4548 (N_4548,N_4481,N_4485);
nor U4549 (N_4549,N_4413,N_4414);
nor U4550 (N_4550,N_4441,N_4487);
and U4551 (N_4551,N_4445,N_4420);
and U4552 (N_4552,N_4498,N_4411);
or U4553 (N_4553,N_4441,N_4489);
nor U4554 (N_4554,N_4408,N_4469);
and U4555 (N_4555,N_4437,N_4466);
or U4556 (N_4556,N_4424,N_4456);
or U4557 (N_4557,N_4402,N_4447);
xor U4558 (N_4558,N_4403,N_4485);
xnor U4559 (N_4559,N_4445,N_4476);
or U4560 (N_4560,N_4461,N_4450);
nor U4561 (N_4561,N_4458,N_4464);
nor U4562 (N_4562,N_4436,N_4404);
nand U4563 (N_4563,N_4441,N_4442);
and U4564 (N_4564,N_4434,N_4490);
or U4565 (N_4565,N_4499,N_4403);
nor U4566 (N_4566,N_4452,N_4458);
nand U4567 (N_4567,N_4470,N_4464);
and U4568 (N_4568,N_4430,N_4446);
and U4569 (N_4569,N_4493,N_4468);
nand U4570 (N_4570,N_4426,N_4477);
nand U4571 (N_4571,N_4424,N_4492);
nand U4572 (N_4572,N_4483,N_4484);
xor U4573 (N_4573,N_4463,N_4475);
nor U4574 (N_4574,N_4449,N_4491);
xor U4575 (N_4575,N_4412,N_4465);
or U4576 (N_4576,N_4469,N_4402);
or U4577 (N_4577,N_4470,N_4479);
xor U4578 (N_4578,N_4456,N_4494);
nor U4579 (N_4579,N_4479,N_4468);
xnor U4580 (N_4580,N_4483,N_4453);
nand U4581 (N_4581,N_4401,N_4434);
nand U4582 (N_4582,N_4439,N_4467);
and U4583 (N_4583,N_4473,N_4427);
xnor U4584 (N_4584,N_4467,N_4488);
xnor U4585 (N_4585,N_4482,N_4413);
nor U4586 (N_4586,N_4441,N_4439);
xnor U4587 (N_4587,N_4428,N_4496);
xnor U4588 (N_4588,N_4451,N_4473);
nand U4589 (N_4589,N_4466,N_4442);
and U4590 (N_4590,N_4486,N_4478);
nor U4591 (N_4591,N_4470,N_4445);
nor U4592 (N_4592,N_4416,N_4444);
nor U4593 (N_4593,N_4409,N_4499);
nor U4594 (N_4594,N_4417,N_4450);
or U4595 (N_4595,N_4406,N_4440);
nand U4596 (N_4596,N_4437,N_4407);
nor U4597 (N_4597,N_4492,N_4495);
xnor U4598 (N_4598,N_4441,N_4436);
and U4599 (N_4599,N_4449,N_4468);
and U4600 (N_4600,N_4585,N_4539);
and U4601 (N_4601,N_4518,N_4531);
xor U4602 (N_4602,N_4586,N_4578);
and U4603 (N_4603,N_4530,N_4589);
and U4604 (N_4604,N_4579,N_4517);
nor U4605 (N_4605,N_4587,N_4506);
nand U4606 (N_4606,N_4521,N_4553);
nor U4607 (N_4607,N_4545,N_4573);
nand U4608 (N_4608,N_4528,N_4583);
and U4609 (N_4609,N_4564,N_4563);
or U4610 (N_4610,N_4592,N_4549);
or U4611 (N_4611,N_4535,N_4559);
nand U4612 (N_4612,N_4581,N_4567);
nand U4613 (N_4613,N_4577,N_4522);
nor U4614 (N_4614,N_4593,N_4524);
xnor U4615 (N_4615,N_4571,N_4576);
xor U4616 (N_4616,N_4594,N_4512);
and U4617 (N_4617,N_4566,N_4514);
xnor U4618 (N_4618,N_4582,N_4548);
or U4619 (N_4619,N_4596,N_4523);
nand U4620 (N_4620,N_4542,N_4546);
and U4621 (N_4621,N_4544,N_4558);
or U4622 (N_4622,N_4557,N_4525);
xnor U4623 (N_4623,N_4516,N_4541);
nor U4624 (N_4624,N_4503,N_4588);
nand U4625 (N_4625,N_4507,N_4561);
or U4626 (N_4626,N_4580,N_4591);
nor U4627 (N_4627,N_4501,N_4500);
or U4628 (N_4628,N_4519,N_4562);
nand U4629 (N_4629,N_4534,N_4554);
and U4630 (N_4630,N_4552,N_4575);
nor U4631 (N_4631,N_4508,N_4536);
nor U4632 (N_4632,N_4513,N_4556);
nand U4633 (N_4633,N_4590,N_4574);
xnor U4634 (N_4634,N_4568,N_4511);
xor U4635 (N_4635,N_4505,N_4565);
or U4636 (N_4636,N_4543,N_4527);
nor U4637 (N_4637,N_4551,N_4509);
or U4638 (N_4638,N_4504,N_4547);
or U4639 (N_4639,N_4555,N_4540);
nor U4640 (N_4640,N_4572,N_4510);
xnor U4641 (N_4641,N_4560,N_4599);
or U4642 (N_4642,N_4502,N_4569);
or U4643 (N_4643,N_4515,N_4570);
and U4644 (N_4644,N_4538,N_4529);
and U4645 (N_4645,N_4520,N_4532);
xor U4646 (N_4646,N_4526,N_4537);
nor U4647 (N_4647,N_4584,N_4595);
xor U4648 (N_4648,N_4533,N_4550);
nand U4649 (N_4649,N_4598,N_4597);
nor U4650 (N_4650,N_4549,N_4595);
nor U4651 (N_4651,N_4529,N_4516);
and U4652 (N_4652,N_4576,N_4545);
or U4653 (N_4653,N_4545,N_4539);
nor U4654 (N_4654,N_4534,N_4558);
and U4655 (N_4655,N_4530,N_4511);
and U4656 (N_4656,N_4551,N_4588);
nand U4657 (N_4657,N_4568,N_4597);
and U4658 (N_4658,N_4524,N_4580);
and U4659 (N_4659,N_4568,N_4578);
or U4660 (N_4660,N_4576,N_4503);
or U4661 (N_4661,N_4524,N_4537);
nor U4662 (N_4662,N_4576,N_4510);
nand U4663 (N_4663,N_4549,N_4582);
xor U4664 (N_4664,N_4525,N_4581);
nor U4665 (N_4665,N_4551,N_4589);
nor U4666 (N_4666,N_4585,N_4570);
nand U4667 (N_4667,N_4506,N_4586);
nand U4668 (N_4668,N_4503,N_4547);
xnor U4669 (N_4669,N_4519,N_4567);
nor U4670 (N_4670,N_4579,N_4571);
nand U4671 (N_4671,N_4586,N_4503);
and U4672 (N_4672,N_4546,N_4509);
or U4673 (N_4673,N_4541,N_4576);
or U4674 (N_4674,N_4520,N_4565);
nand U4675 (N_4675,N_4536,N_4588);
nor U4676 (N_4676,N_4580,N_4585);
nand U4677 (N_4677,N_4573,N_4500);
nor U4678 (N_4678,N_4585,N_4553);
nor U4679 (N_4679,N_4567,N_4593);
or U4680 (N_4680,N_4573,N_4556);
and U4681 (N_4681,N_4554,N_4582);
nor U4682 (N_4682,N_4597,N_4595);
and U4683 (N_4683,N_4515,N_4597);
and U4684 (N_4684,N_4581,N_4504);
and U4685 (N_4685,N_4512,N_4545);
and U4686 (N_4686,N_4538,N_4569);
and U4687 (N_4687,N_4590,N_4510);
or U4688 (N_4688,N_4598,N_4539);
nand U4689 (N_4689,N_4563,N_4533);
xnor U4690 (N_4690,N_4597,N_4559);
nand U4691 (N_4691,N_4512,N_4537);
xor U4692 (N_4692,N_4586,N_4558);
nand U4693 (N_4693,N_4516,N_4535);
or U4694 (N_4694,N_4508,N_4548);
and U4695 (N_4695,N_4546,N_4552);
nand U4696 (N_4696,N_4585,N_4536);
nand U4697 (N_4697,N_4500,N_4597);
nor U4698 (N_4698,N_4582,N_4505);
xor U4699 (N_4699,N_4574,N_4507);
or U4700 (N_4700,N_4673,N_4644);
or U4701 (N_4701,N_4637,N_4664);
nand U4702 (N_4702,N_4655,N_4636);
and U4703 (N_4703,N_4683,N_4617);
and U4704 (N_4704,N_4616,N_4698);
and U4705 (N_4705,N_4696,N_4661);
xnor U4706 (N_4706,N_4690,N_4632);
and U4707 (N_4707,N_4658,N_4640);
nor U4708 (N_4708,N_4675,N_4600);
xor U4709 (N_4709,N_4680,N_4672);
and U4710 (N_4710,N_4693,N_4666);
xnor U4711 (N_4711,N_4626,N_4692);
and U4712 (N_4712,N_4678,N_4685);
or U4713 (N_4713,N_4684,N_4614);
xor U4714 (N_4714,N_4646,N_4631);
nand U4715 (N_4715,N_4689,N_4629);
xor U4716 (N_4716,N_4653,N_4652);
xor U4717 (N_4717,N_4662,N_4687);
nand U4718 (N_4718,N_4603,N_4628);
or U4719 (N_4719,N_4639,N_4665);
nand U4720 (N_4720,N_4668,N_4610);
nor U4721 (N_4721,N_4604,N_4677);
xor U4722 (N_4722,N_4618,N_4633);
and U4723 (N_4723,N_4630,N_4697);
nand U4724 (N_4724,N_4695,N_4623);
nor U4725 (N_4725,N_4624,N_4635);
or U4726 (N_4726,N_4670,N_4627);
or U4727 (N_4727,N_4679,N_4657);
or U4728 (N_4728,N_4602,N_4642);
or U4729 (N_4729,N_4619,N_4608);
nor U4730 (N_4730,N_4620,N_4621);
nor U4731 (N_4731,N_4625,N_4613);
and U4732 (N_4732,N_4615,N_4648);
xor U4733 (N_4733,N_4609,N_4611);
and U4734 (N_4734,N_4686,N_4601);
nor U4735 (N_4735,N_4669,N_4651);
xor U4736 (N_4736,N_4622,N_4643);
xnor U4737 (N_4737,N_4649,N_4663);
nor U4738 (N_4738,N_4659,N_4650);
nand U4739 (N_4739,N_4671,N_4660);
nand U4740 (N_4740,N_4605,N_4656);
nor U4741 (N_4741,N_4667,N_4645);
and U4742 (N_4742,N_4638,N_4691);
nand U4743 (N_4743,N_4688,N_4699);
nand U4744 (N_4744,N_4654,N_4647);
xnor U4745 (N_4745,N_4681,N_4641);
xor U4746 (N_4746,N_4694,N_4612);
nand U4747 (N_4747,N_4607,N_4674);
and U4748 (N_4748,N_4682,N_4634);
nand U4749 (N_4749,N_4606,N_4676);
or U4750 (N_4750,N_4608,N_4604);
nor U4751 (N_4751,N_4613,N_4667);
or U4752 (N_4752,N_4662,N_4653);
and U4753 (N_4753,N_4633,N_4661);
and U4754 (N_4754,N_4686,N_4619);
and U4755 (N_4755,N_4631,N_4637);
xor U4756 (N_4756,N_4682,N_4636);
or U4757 (N_4757,N_4686,N_4663);
or U4758 (N_4758,N_4693,N_4648);
nor U4759 (N_4759,N_4635,N_4631);
nand U4760 (N_4760,N_4618,N_4667);
and U4761 (N_4761,N_4655,N_4686);
or U4762 (N_4762,N_4627,N_4635);
nor U4763 (N_4763,N_4601,N_4642);
nand U4764 (N_4764,N_4603,N_4675);
and U4765 (N_4765,N_4611,N_4663);
nand U4766 (N_4766,N_4691,N_4674);
or U4767 (N_4767,N_4670,N_4642);
nand U4768 (N_4768,N_4651,N_4622);
xor U4769 (N_4769,N_4677,N_4606);
and U4770 (N_4770,N_4683,N_4671);
xnor U4771 (N_4771,N_4661,N_4638);
xnor U4772 (N_4772,N_4657,N_4677);
nor U4773 (N_4773,N_4656,N_4639);
nand U4774 (N_4774,N_4693,N_4645);
nand U4775 (N_4775,N_4625,N_4691);
and U4776 (N_4776,N_4644,N_4691);
nand U4777 (N_4777,N_4694,N_4605);
and U4778 (N_4778,N_4623,N_4643);
nor U4779 (N_4779,N_4618,N_4665);
nand U4780 (N_4780,N_4624,N_4668);
or U4781 (N_4781,N_4698,N_4686);
xnor U4782 (N_4782,N_4653,N_4648);
and U4783 (N_4783,N_4648,N_4602);
nand U4784 (N_4784,N_4671,N_4669);
and U4785 (N_4785,N_4611,N_4699);
or U4786 (N_4786,N_4606,N_4656);
or U4787 (N_4787,N_4689,N_4698);
xor U4788 (N_4788,N_4656,N_4686);
xnor U4789 (N_4789,N_4633,N_4676);
nor U4790 (N_4790,N_4614,N_4628);
nand U4791 (N_4791,N_4609,N_4664);
or U4792 (N_4792,N_4603,N_4665);
nor U4793 (N_4793,N_4616,N_4603);
nand U4794 (N_4794,N_4612,N_4637);
and U4795 (N_4795,N_4620,N_4618);
xnor U4796 (N_4796,N_4655,N_4664);
nand U4797 (N_4797,N_4689,N_4660);
nand U4798 (N_4798,N_4646,N_4698);
nor U4799 (N_4799,N_4658,N_4660);
or U4800 (N_4800,N_4753,N_4726);
nand U4801 (N_4801,N_4762,N_4787);
nand U4802 (N_4802,N_4752,N_4722);
xor U4803 (N_4803,N_4713,N_4741);
nor U4804 (N_4804,N_4767,N_4792);
or U4805 (N_4805,N_4789,N_4750);
nand U4806 (N_4806,N_4764,N_4772);
nand U4807 (N_4807,N_4725,N_4755);
or U4808 (N_4808,N_4735,N_4745);
xnor U4809 (N_4809,N_4791,N_4718);
xor U4810 (N_4810,N_4758,N_4721);
nor U4811 (N_4811,N_4784,N_4723);
nand U4812 (N_4812,N_4714,N_4786);
or U4813 (N_4813,N_4731,N_4727);
nand U4814 (N_4814,N_4742,N_4773);
nor U4815 (N_4815,N_4782,N_4740);
xnor U4816 (N_4816,N_4790,N_4747);
xnor U4817 (N_4817,N_4738,N_4770);
nand U4818 (N_4818,N_4730,N_4719);
nor U4819 (N_4819,N_4724,N_4701);
or U4820 (N_4820,N_4748,N_4708);
and U4821 (N_4821,N_4785,N_4761);
and U4822 (N_4822,N_4771,N_4715);
nand U4823 (N_4823,N_4768,N_4759);
and U4824 (N_4824,N_4795,N_4799);
nor U4825 (N_4825,N_4706,N_4728);
nor U4826 (N_4826,N_4756,N_4775);
nor U4827 (N_4827,N_4705,N_4797);
and U4828 (N_4828,N_4788,N_4746);
nor U4829 (N_4829,N_4707,N_4776);
or U4830 (N_4830,N_4751,N_4736);
and U4831 (N_4831,N_4757,N_4783);
nor U4832 (N_4832,N_4737,N_4765);
xor U4833 (N_4833,N_4743,N_4754);
xnor U4834 (N_4834,N_4702,N_4717);
or U4835 (N_4835,N_4739,N_4734);
and U4836 (N_4836,N_4793,N_4774);
xnor U4837 (N_4837,N_4744,N_4777);
xor U4838 (N_4838,N_4704,N_4766);
and U4839 (N_4839,N_4749,N_4763);
xor U4840 (N_4840,N_4778,N_4798);
xnor U4841 (N_4841,N_4779,N_4712);
nor U4842 (N_4842,N_4711,N_4703);
nor U4843 (N_4843,N_4794,N_4760);
nand U4844 (N_4844,N_4732,N_4700);
and U4845 (N_4845,N_4780,N_4781);
or U4846 (N_4846,N_4720,N_4716);
nor U4847 (N_4847,N_4769,N_4710);
nand U4848 (N_4848,N_4709,N_4733);
nor U4849 (N_4849,N_4729,N_4796);
or U4850 (N_4850,N_4775,N_4786);
or U4851 (N_4851,N_4720,N_4742);
nor U4852 (N_4852,N_4796,N_4784);
or U4853 (N_4853,N_4783,N_4746);
and U4854 (N_4854,N_4778,N_4773);
nand U4855 (N_4855,N_4719,N_4706);
xor U4856 (N_4856,N_4753,N_4766);
or U4857 (N_4857,N_4747,N_4736);
or U4858 (N_4858,N_4730,N_4785);
nor U4859 (N_4859,N_4713,N_4757);
nor U4860 (N_4860,N_4755,N_4720);
and U4861 (N_4861,N_4725,N_4759);
or U4862 (N_4862,N_4752,N_4718);
and U4863 (N_4863,N_4764,N_4722);
and U4864 (N_4864,N_4738,N_4732);
and U4865 (N_4865,N_4706,N_4701);
or U4866 (N_4866,N_4703,N_4727);
nor U4867 (N_4867,N_4779,N_4760);
or U4868 (N_4868,N_4712,N_4781);
nand U4869 (N_4869,N_4727,N_4734);
or U4870 (N_4870,N_4760,N_4791);
xnor U4871 (N_4871,N_4752,N_4704);
or U4872 (N_4872,N_4791,N_4712);
or U4873 (N_4873,N_4797,N_4741);
nor U4874 (N_4874,N_4736,N_4778);
or U4875 (N_4875,N_4722,N_4744);
or U4876 (N_4876,N_4771,N_4724);
nor U4877 (N_4877,N_4741,N_4779);
nor U4878 (N_4878,N_4738,N_4702);
nand U4879 (N_4879,N_4763,N_4788);
and U4880 (N_4880,N_4778,N_4760);
nand U4881 (N_4881,N_4701,N_4708);
or U4882 (N_4882,N_4739,N_4708);
nor U4883 (N_4883,N_4799,N_4701);
xnor U4884 (N_4884,N_4797,N_4737);
nor U4885 (N_4885,N_4718,N_4710);
xnor U4886 (N_4886,N_4707,N_4751);
xnor U4887 (N_4887,N_4751,N_4740);
nor U4888 (N_4888,N_4730,N_4722);
nor U4889 (N_4889,N_4723,N_4772);
nor U4890 (N_4890,N_4764,N_4736);
xnor U4891 (N_4891,N_4756,N_4706);
xor U4892 (N_4892,N_4733,N_4720);
nand U4893 (N_4893,N_4706,N_4704);
nand U4894 (N_4894,N_4715,N_4770);
or U4895 (N_4895,N_4721,N_4792);
nand U4896 (N_4896,N_4761,N_4731);
and U4897 (N_4897,N_4752,N_4779);
and U4898 (N_4898,N_4739,N_4779);
nand U4899 (N_4899,N_4712,N_4740);
nor U4900 (N_4900,N_4842,N_4898);
or U4901 (N_4901,N_4822,N_4875);
xor U4902 (N_4902,N_4834,N_4829);
nor U4903 (N_4903,N_4819,N_4899);
xnor U4904 (N_4904,N_4877,N_4856);
or U4905 (N_4905,N_4806,N_4845);
nor U4906 (N_4906,N_4886,N_4867);
xor U4907 (N_4907,N_4801,N_4866);
and U4908 (N_4908,N_4804,N_4884);
or U4909 (N_4909,N_4817,N_4827);
nand U4910 (N_4910,N_4812,N_4835);
or U4911 (N_4911,N_4839,N_4805);
and U4912 (N_4912,N_4854,N_4873);
or U4913 (N_4913,N_4855,N_4870);
nor U4914 (N_4914,N_4864,N_4825);
and U4915 (N_4915,N_4815,N_4888);
nor U4916 (N_4916,N_4860,N_4879);
xor U4917 (N_4917,N_4897,N_4844);
or U4918 (N_4918,N_4818,N_4865);
nand U4919 (N_4919,N_4826,N_4803);
nor U4920 (N_4920,N_4871,N_4807);
nor U4921 (N_4921,N_4885,N_4861);
and U4922 (N_4922,N_4894,N_4892);
or U4923 (N_4923,N_4830,N_4832);
and U4924 (N_4924,N_4893,N_4810);
nor U4925 (N_4925,N_4838,N_4802);
xnor U4926 (N_4926,N_4828,N_4800);
nand U4927 (N_4927,N_4851,N_4863);
or U4928 (N_4928,N_4895,N_4824);
and U4929 (N_4929,N_4883,N_4869);
nor U4930 (N_4930,N_4882,N_4813);
xnor U4931 (N_4931,N_4823,N_4889);
nor U4932 (N_4932,N_4859,N_4831);
xnor U4933 (N_4933,N_4808,N_4833);
xnor U4934 (N_4934,N_4816,N_4847);
nand U4935 (N_4935,N_4857,N_4858);
nand U4936 (N_4936,N_4896,N_4821);
nor U4937 (N_4937,N_4891,N_4846);
and U4938 (N_4938,N_4850,N_4880);
and U4939 (N_4939,N_4862,N_4848);
xnor U4940 (N_4940,N_4814,N_4820);
and U4941 (N_4941,N_4890,N_4872);
xnor U4942 (N_4942,N_4811,N_4840);
nand U4943 (N_4943,N_4852,N_4878);
and U4944 (N_4944,N_4837,N_4881);
or U4945 (N_4945,N_4887,N_4836);
xor U4946 (N_4946,N_4849,N_4874);
xor U4947 (N_4947,N_4809,N_4853);
and U4948 (N_4948,N_4876,N_4868);
or U4949 (N_4949,N_4843,N_4841);
or U4950 (N_4950,N_4836,N_4825);
nand U4951 (N_4951,N_4841,N_4879);
and U4952 (N_4952,N_4870,N_4877);
or U4953 (N_4953,N_4871,N_4824);
xnor U4954 (N_4954,N_4848,N_4831);
or U4955 (N_4955,N_4803,N_4871);
or U4956 (N_4956,N_4850,N_4873);
nor U4957 (N_4957,N_4865,N_4888);
nand U4958 (N_4958,N_4840,N_4851);
nand U4959 (N_4959,N_4880,N_4814);
and U4960 (N_4960,N_4887,N_4868);
or U4961 (N_4961,N_4818,N_4868);
or U4962 (N_4962,N_4880,N_4867);
and U4963 (N_4963,N_4812,N_4831);
and U4964 (N_4964,N_4822,N_4879);
or U4965 (N_4965,N_4843,N_4828);
and U4966 (N_4966,N_4899,N_4867);
nand U4967 (N_4967,N_4820,N_4862);
or U4968 (N_4968,N_4876,N_4857);
xnor U4969 (N_4969,N_4888,N_4818);
nand U4970 (N_4970,N_4832,N_4851);
xnor U4971 (N_4971,N_4813,N_4822);
and U4972 (N_4972,N_4858,N_4803);
nor U4973 (N_4973,N_4843,N_4875);
or U4974 (N_4974,N_4832,N_4874);
xor U4975 (N_4975,N_4898,N_4890);
or U4976 (N_4976,N_4849,N_4898);
nand U4977 (N_4977,N_4802,N_4827);
or U4978 (N_4978,N_4846,N_4818);
xnor U4979 (N_4979,N_4805,N_4823);
nand U4980 (N_4980,N_4825,N_4820);
or U4981 (N_4981,N_4898,N_4891);
and U4982 (N_4982,N_4866,N_4820);
or U4983 (N_4983,N_4884,N_4894);
nand U4984 (N_4984,N_4841,N_4803);
or U4985 (N_4985,N_4859,N_4892);
and U4986 (N_4986,N_4895,N_4866);
xor U4987 (N_4987,N_4825,N_4845);
nor U4988 (N_4988,N_4859,N_4829);
nor U4989 (N_4989,N_4864,N_4892);
xor U4990 (N_4990,N_4867,N_4846);
nand U4991 (N_4991,N_4836,N_4822);
nor U4992 (N_4992,N_4802,N_4806);
nor U4993 (N_4993,N_4808,N_4896);
nor U4994 (N_4994,N_4874,N_4868);
nand U4995 (N_4995,N_4858,N_4853);
or U4996 (N_4996,N_4816,N_4882);
nor U4997 (N_4997,N_4838,N_4885);
and U4998 (N_4998,N_4810,N_4885);
xnor U4999 (N_4999,N_4872,N_4816);
nand U5000 (N_5000,N_4994,N_4982);
or U5001 (N_5001,N_4956,N_4924);
nor U5002 (N_5002,N_4983,N_4915);
nor U5003 (N_5003,N_4954,N_4977);
nor U5004 (N_5004,N_4930,N_4973);
or U5005 (N_5005,N_4993,N_4996);
nand U5006 (N_5006,N_4905,N_4918);
or U5007 (N_5007,N_4914,N_4942);
and U5008 (N_5008,N_4992,N_4951);
nor U5009 (N_5009,N_4969,N_4921);
xor U5010 (N_5010,N_4980,N_4974);
nand U5011 (N_5011,N_4900,N_4986);
nor U5012 (N_5012,N_4988,N_4941);
nor U5013 (N_5013,N_4984,N_4943);
xor U5014 (N_5014,N_4923,N_4965);
nor U5015 (N_5015,N_4932,N_4995);
nand U5016 (N_5016,N_4935,N_4937);
or U5017 (N_5017,N_4911,N_4902);
and U5018 (N_5018,N_4945,N_4931);
or U5019 (N_5019,N_4952,N_4946);
xor U5020 (N_5020,N_4957,N_4916);
nor U5021 (N_5021,N_4936,N_4949);
nand U5022 (N_5022,N_4978,N_4987);
nand U5023 (N_5023,N_4958,N_4925);
nand U5024 (N_5024,N_4922,N_4960);
xor U5025 (N_5025,N_4997,N_4990);
xor U5026 (N_5026,N_4967,N_4939);
or U5027 (N_5027,N_4962,N_4908);
and U5028 (N_5028,N_4947,N_4975);
and U5029 (N_5029,N_4991,N_4964);
nor U5030 (N_5030,N_4940,N_4929);
xor U5031 (N_5031,N_4981,N_4913);
nor U5032 (N_5032,N_4955,N_4917);
xor U5033 (N_5033,N_4959,N_4919);
or U5034 (N_5034,N_4933,N_4934);
or U5035 (N_5035,N_4903,N_4901);
and U5036 (N_5036,N_4944,N_4904);
xnor U5037 (N_5037,N_4961,N_4907);
nand U5038 (N_5038,N_4910,N_4948);
or U5039 (N_5039,N_4999,N_4953);
or U5040 (N_5040,N_4971,N_4985);
or U5041 (N_5041,N_4979,N_4920);
and U5042 (N_5042,N_4906,N_4938);
xnor U5043 (N_5043,N_4998,N_4928);
xor U5044 (N_5044,N_4966,N_4912);
nand U5045 (N_5045,N_4970,N_4989);
nor U5046 (N_5046,N_4927,N_4976);
and U5047 (N_5047,N_4963,N_4968);
nand U5048 (N_5048,N_4926,N_4909);
and U5049 (N_5049,N_4950,N_4972);
xnor U5050 (N_5050,N_4984,N_4972);
xor U5051 (N_5051,N_4995,N_4904);
and U5052 (N_5052,N_4961,N_4955);
xnor U5053 (N_5053,N_4984,N_4974);
xnor U5054 (N_5054,N_4955,N_4948);
or U5055 (N_5055,N_4974,N_4931);
or U5056 (N_5056,N_4946,N_4943);
nand U5057 (N_5057,N_4917,N_4999);
nand U5058 (N_5058,N_4938,N_4927);
nand U5059 (N_5059,N_4938,N_4954);
nor U5060 (N_5060,N_4960,N_4968);
nor U5061 (N_5061,N_4920,N_4922);
xor U5062 (N_5062,N_4902,N_4984);
nand U5063 (N_5063,N_4994,N_4977);
nand U5064 (N_5064,N_4948,N_4915);
nand U5065 (N_5065,N_4997,N_4949);
nand U5066 (N_5066,N_4916,N_4917);
and U5067 (N_5067,N_4924,N_4952);
and U5068 (N_5068,N_4928,N_4930);
nand U5069 (N_5069,N_4953,N_4904);
or U5070 (N_5070,N_4941,N_4911);
nand U5071 (N_5071,N_4997,N_4945);
nand U5072 (N_5072,N_4970,N_4931);
or U5073 (N_5073,N_4957,N_4909);
xor U5074 (N_5074,N_4924,N_4958);
or U5075 (N_5075,N_4998,N_4916);
or U5076 (N_5076,N_4957,N_4992);
and U5077 (N_5077,N_4903,N_4974);
and U5078 (N_5078,N_4959,N_4926);
or U5079 (N_5079,N_4948,N_4981);
or U5080 (N_5080,N_4998,N_4932);
xnor U5081 (N_5081,N_4902,N_4960);
and U5082 (N_5082,N_4981,N_4953);
and U5083 (N_5083,N_4988,N_4976);
nand U5084 (N_5084,N_4951,N_4925);
nor U5085 (N_5085,N_4916,N_4903);
nand U5086 (N_5086,N_4916,N_4949);
nand U5087 (N_5087,N_4949,N_4953);
nand U5088 (N_5088,N_4982,N_4956);
and U5089 (N_5089,N_4905,N_4953);
nand U5090 (N_5090,N_4915,N_4936);
and U5091 (N_5091,N_4957,N_4925);
nand U5092 (N_5092,N_4941,N_4903);
and U5093 (N_5093,N_4963,N_4993);
and U5094 (N_5094,N_4985,N_4907);
nor U5095 (N_5095,N_4926,N_4994);
or U5096 (N_5096,N_4967,N_4996);
xor U5097 (N_5097,N_4980,N_4956);
or U5098 (N_5098,N_4940,N_4942);
nor U5099 (N_5099,N_4939,N_4973);
xnor U5100 (N_5100,N_5042,N_5075);
or U5101 (N_5101,N_5007,N_5016);
xor U5102 (N_5102,N_5090,N_5023);
xnor U5103 (N_5103,N_5089,N_5085);
nor U5104 (N_5104,N_5098,N_5040);
or U5105 (N_5105,N_5044,N_5011);
or U5106 (N_5106,N_5019,N_5045);
and U5107 (N_5107,N_5022,N_5035);
and U5108 (N_5108,N_5029,N_5036);
nor U5109 (N_5109,N_5084,N_5061);
nand U5110 (N_5110,N_5058,N_5021);
and U5111 (N_5111,N_5073,N_5010);
nand U5112 (N_5112,N_5081,N_5018);
xor U5113 (N_5113,N_5039,N_5052);
nand U5114 (N_5114,N_5067,N_5094);
and U5115 (N_5115,N_5064,N_5009);
and U5116 (N_5116,N_5063,N_5051);
xor U5117 (N_5117,N_5031,N_5096);
nor U5118 (N_5118,N_5093,N_5032);
and U5119 (N_5119,N_5095,N_5088);
nor U5120 (N_5120,N_5086,N_5001);
nor U5121 (N_5121,N_5078,N_5028);
nand U5122 (N_5122,N_5015,N_5097);
or U5123 (N_5123,N_5047,N_5072);
and U5124 (N_5124,N_5087,N_5082);
and U5125 (N_5125,N_5079,N_5033);
and U5126 (N_5126,N_5092,N_5099);
or U5127 (N_5127,N_5025,N_5002);
nor U5128 (N_5128,N_5062,N_5026);
nand U5129 (N_5129,N_5020,N_5043);
and U5130 (N_5130,N_5012,N_5059);
xnor U5131 (N_5131,N_5048,N_5037);
nor U5132 (N_5132,N_5068,N_5046);
or U5133 (N_5133,N_5041,N_5038);
or U5134 (N_5134,N_5076,N_5006);
xnor U5135 (N_5135,N_5008,N_5024);
and U5136 (N_5136,N_5066,N_5083);
xnor U5137 (N_5137,N_5074,N_5049);
nand U5138 (N_5138,N_5014,N_5034);
and U5139 (N_5139,N_5091,N_5060);
or U5140 (N_5140,N_5056,N_5005);
nor U5141 (N_5141,N_5003,N_5077);
nor U5142 (N_5142,N_5070,N_5004);
or U5143 (N_5143,N_5071,N_5069);
nand U5144 (N_5144,N_5053,N_5055);
nor U5145 (N_5145,N_5050,N_5017);
and U5146 (N_5146,N_5057,N_5030);
xnor U5147 (N_5147,N_5080,N_5013);
nand U5148 (N_5148,N_5065,N_5054);
xor U5149 (N_5149,N_5000,N_5027);
xor U5150 (N_5150,N_5021,N_5013);
or U5151 (N_5151,N_5067,N_5076);
or U5152 (N_5152,N_5087,N_5062);
and U5153 (N_5153,N_5012,N_5002);
and U5154 (N_5154,N_5018,N_5095);
or U5155 (N_5155,N_5055,N_5040);
and U5156 (N_5156,N_5096,N_5078);
and U5157 (N_5157,N_5047,N_5035);
or U5158 (N_5158,N_5049,N_5004);
nor U5159 (N_5159,N_5051,N_5049);
nand U5160 (N_5160,N_5018,N_5045);
xnor U5161 (N_5161,N_5064,N_5012);
or U5162 (N_5162,N_5002,N_5042);
nand U5163 (N_5163,N_5002,N_5043);
and U5164 (N_5164,N_5004,N_5054);
xor U5165 (N_5165,N_5047,N_5060);
nand U5166 (N_5166,N_5042,N_5047);
and U5167 (N_5167,N_5017,N_5073);
or U5168 (N_5168,N_5004,N_5095);
nand U5169 (N_5169,N_5066,N_5011);
and U5170 (N_5170,N_5039,N_5071);
nor U5171 (N_5171,N_5011,N_5050);
xor U5172 (N_5172,N_5060,N_5016);
nor U5173 (N_5173,N_5079,N_5088);
and U5174 (N_5174,N_5067,N_5026);
nand U5175 (N_5175,N_5008,N_5026);
nor U5176 (N_5176,N_5056,N_5023);
and U5177 (N_5177,N_5045,N_5066);
xor U5178 (N_5178,N_5050,N_5002);
or U5179 (N_5179,N_5019,N_5032);
and U5180 (N_5180,N_5092,N_5025);
and U5181 (N_5181,N_5081,N_5085);
nor U5182 (N_5182,N_5073,N_5055);
nand U5183 (N_5183,N_5096,N_5075);
xnor U5184 (N_5184,N_5034,N_5079);
nand U5185 (N_5185,N_5080,N_5033);
nand U5186 (N_5186,N_5090,N_5085);
and U5187 (N_5187,N_5044,N_5037);
xnor U5188 (N_5188,N_5093,N_5067);
nor U5189 (N_5189,N_5063,N_5014);
nor U5190 (N_5190,N_5020,N_5036);
nand U5191 (N_5191,N_5054,N_5029);
nand U5192 (N_5192,N_5016,N_5071);
xor U5193 (N_5193,N_5052,N_5021);
nand U5194 (N_5194,N_5000,N_5064);
and U5195 (N_5195,N_5071,N_5091);
xnor U5196 (N_5196,N_5063,N_5054);
nor U5197 (N_5197,N_5019,N_5038);
or U5198 (N_5198,N_5040,N_5081);
xnor U5199 (N_5199,N_5082,N_5077);
or U5200 (N_5200,N_5108,N_5120);
and U5201 (N_5201,N_5174,N_5106);
xor U5202 (N_5202,N_5117,N_5175);
nand U5203 (N_5203,N_5109,N_5156);
nor U5204 (N_5204,N_5180,N_5190);
nor U5205 (N_5205,N_5199,N_5164);
and U5206 (N_5206,N_5144,N_5196);
or U5207 (N_5207,N_5100,N_5188);
and U5208 (N_5208,N_5126,N_5197);
nor U5209 (N_5209,N_5158,N_5107);
or U5210 (N_5210,N_5162,N_5134);
nor U5211 (N_5211,N_5194,N_5157);
nand U5212 (N_5212,N_5123,N_5142);
or U5213 (N_5213,N_5119,N_5130);
and U5214 (N_5214,N_5104,N_5133);
nor U5215 (N_5215,N_5148,N_5193);
xor U5216 (N_5216,N_5121,N_5176);
or U5217 (N_5217,N_5150,N_5173);
xnor U5218 (N_5218,N_5113,N_5165);
or U5219 (N_5219,N_5186,N_5184);
and U5220 (N_5220,N_5139,N_5127);
nand U5221 (N_5221,N_5140,N_5131);
nor U5222 (N_5222,N_5163,N_5195);
xor U5223 (N_5223,N_5198,N_5161);
xor U5224 (N_5224,N_5122,N_5118);
and U5225 (N_5225,N_5181,N_5103);
or U5226 (N_5226,N_5101,N_5114);
and U5227 (N_5227,N_5179,N_5149);
or U5228 (N_5228,N_5124,N_5137);
nor U5229 (N_5229,N_5129,N_5125);
xnor U5230 (N_5230,N_5151,N_5182);
or U5231 (N_5231,N_5155,N_5105);
xnor U5232 (N_5232,N_5135,N_5168);
xnor U5233 (N_5233,N_5160,N_5171);
or U5234 (N_5234,N_5183,N_5159);
xnor U5235 (N_5235,N_5146,N_5153);
or U5236 (N_5236,N_5141,N_5110);
and U5237 (N_5237,N_5128,N_5143);
or U5238 (N_5238,N_5187,N_5132);
or U5239 (N_5239,N_5167,N_5154);
or U5240 (N_5240,N_5170,N_5115);
nor U5241 (N_5241,N_5169,N_5177);
or U5242 (N_5242,N_5147,N_5166);
nand U5243 (N_5243,N_5145,N_5185);
xnor U5244 (N_5244,N_5116,N_5102);
or U5245 (N_5245,N_5192,N_5112);
or U5246 (N_5246,N_5136,N_5191);
nor U5247 (N_5247,N_5138,N_5178);
or U5248 (N_5248,N_5111,N_5172);
nand U5249 (N_5249,N_5189,N_5152);
and U5250 (N_5250,N_5101,N_5168);
xnor U5251 (N_5251,N_5138,N_5165);
nand U5252 (N_5252,N_5103,N_5126);
and U5253 (N_5253,N_5174,N_5154);
xor U5254 (N_5254,N_5151,N_5122);
xnor U5255 (N_5255,N_5123,N_5199);
and U5256 (N_5256,N_5135,N_5111);
xor U5257 (N_5257,N_5166,N_5157);
and U5258 (N_5258,N_5131,N_5196);
nor U5259 (N_5259,N_5144,N_5120);
nand U5260 (N_5260,N_5121,N_5103);
xor U5261 (N_5261,N_5193,N_5144);
nor U5262 (N_5262,N_5191,N_5198);
xor U5263 (N_5263,N_5111,N_5129);
nand U5264 (N_5264,N_5134,N_5174);
and U5265 (N_5265,N_5155,N_5111);
xor U5266 (N_5266,N_5160,N_5153);
nand U5267 (N_5267,N_5107,N_5184);
or U5268 (N_5268,N_5159,N_5157);
nand U5269 (N_5269,N_5116,N_5167);
nor U5270 (N_5270,N_5182,N_5183);
or U5271 (N_5271,N_5145,N_5144);
nor U5272 (N_5272,N_5179,N_5110);
or U5273 (N_5273,N_5116,N_5194);
nand U5274 (N_5274,N_5123,N_5185);
nand U5275 (N_5275,N_5197,N_5181);
and U5276 (N_5276,N_5130,N_5199);
xor U5277 (N_5277,N_5110,N_5148);
or U5278 (N_5278,N_5198,N_5114);
nand U5279 (N_5279,N_5101,N_5108);
or U5280 (N_5280,N_5121,N_5110);
xnor U5281 (N_5281,N_5121,N_5171);
or U5282 (N_5282,N_5170,N_5154);
and U5283 (N_5283,N_5180,N_5126);
nand U5284 (N_5284,N_5131,N_5149);
or U5285 (N_5285,N_5180,N_5170);
nor U5286 (N_5286,N_5128,N_5101);
xnor U5287 (N_5287,N_5153,N_5107);
and U5288 (N_5288,N_5141,N_5191);
xnor U5289 (N_5289,N_5166,N_5129);
nand U5290 (N_5290,N_5117,N_5179);
nor U5291 (N_5291,N_5169,N_5100);
nand U5292 (N_5292,N_5114,N_5144);
nor U5293 (N_5293,N_5103,N_5101);
and U5294 (N_5294,N_5108,N_5165);
nand U5295 (N_5295,N_5199,N_5137);
nor U5296 (N_5296,N_5119,N_5114);
nor U5297 (N_5297,N_5152,N_5108);
and U5298 (N_5298,N_5183,N_5178);
xnor U5299 (N_5299,N_5102,N_5101);
or U5300 (N_5300,N_5220,N_5210);
nor U5301 (N_5301,N_5225,N_5260);
xor U5302 (N_5302,N_5270,N_5258);
nand U5303 (N_5303,N_5293,N_5217);
and U5304 (N_5304,N_5268,N_5246);
or U5305 (N_5305,N_5266,N_5205);
nand U5306 (N_5306,N_5292,N_5255);
nand U5307 (N_5307,N_5243,N_5227);
and U5308 (N_5308,N_5263,N_5213);
nand U5309 (N_5309,N_5275,N_5272);
or U5310 (N_5310,N_5233,N_5276);
or U5311 (N_5311,N_5207,N_5239);
nor U5312 (N_5312,N_5242,N_5256);
nor U5313 (N_5313,N_5281,N_5222);
or U5314 (N_5314,N_5261,N_5248);
or U5315 (N_5315,N_5271,N_5278);
nor U5316 (N_5316,N_5259,N_5228);
or U5317 (N_5317,N_5290,N_5234);
nand U5318 (N_5318,N_5282,N_5201);
or U5319 (N_5319,N_5286,N_5264);
xor U5320 (N_5320,N_5288,N_5229);
xnor U5321 (N_5321,N_5257,N_5279);
nor U5322 (N_5322,N_5235,N_5251);
nor U5323 (N_5323,N_5262,N_5216);
nand U5324 (N_5324,N_5203,N_5218);
and U5325 (N_5325,N_5249,N_5223);
nand U5326 (N_5326,N_5244,N_5224);
nor U5327 (N_5327,N_5232,N_5284);
nor U5328 (N_5328,N_5231,N_5206);
and U5329 (N_5329,N_5245,N_5287);
nand U5330 (N_5330,N_5267,N_5208);
xor U5331 (N_5331,N_5285,N_5202);
and U5332 (N_5332,N_5219,N_5280);
xor U5333 (N_5333,N_5241,N_5226);
nand U5334 (N_5334,N_5291,N_5294);
xor U5335 (N_5335,N_5265,N_5215);
nor U5336 (N_5336,N_5273,N_5277);
nand U5337 (N_5337,N_5240,N_5297);
nor U5338 (N_5338,N_5253,N_5254);
or U5339 (N_5339,N_5238,N_5211);
xnor U5340 (N_5340,N_5299,N_5214);
nor U5341 (N_5341,N_5237,N_5298);
and U5342 (N_5342,N_5212,N_5274);
nor U5343 (N_5343,N_5230,N_5289);
and U5344 (N_5344,N_5283,N_5252);
nand U5345 (N_5345,N_5269,N_5209);
and U5346 (N_5346,N_5250,N_5296);
nor U5347 (N_5347,N_5221,N_5236);
and U5348 (N_5348,N_5200,N_5247);
nor U5349 (N_5349,N_5204,N_5295);
nand U5350 (N_5350,N_5229,N_5265);
nor U5351 (N_5351,N_5278,N_5269);
xor U5352 (N_5352,N_5211,N_5254);
and U5353 (N_5353,N_5200,N_5218);
and U5354 (N_5354,N_5271,N_5290);
and U5355 (N_5355,N_5294,N_5296);
xnor U5356 (N_5356,N_5219,N_5208);
nand U5357 (N_5357,N_5286,N_5202);
or U5358 (N_5358,N_5287,N_5229);
nand U5359 (N_5359,N_5236,N_5232);
nor U5360 (N_5360,N_5209,N_5257);
nor U5361 (N_5361,N_5201,N_5213);
nand U5362 (N_5362,N_5278,N_5280);
and U5363 (N_5363,N_5275,N_5203);
or U5364 (N_5364,N_5209,N_5297);
or U5365 (N_5365,N_5219,N_5251);
xor U5366 (N_5366,N_5223,N_5286);
and U5367 (N_5367,N_5205,N_5235);
or U5368 (N_5368,N_5225,N_5210);
and U5369 (N_5369,N_5280,N_5216);
xor U5370 (N_5370,N_5226,N_5278);
or U5371 (N_5371,N_5230,N_5219);
or U5372 (N_5372,N_5257,N_5298);
or U5373 (N_5373,N_5204,N_5261);
xor U5374 (N_5374,N_5216,N_5256);
and U5375 (N_5375,N_5275,N_5292);
and U5376 (N_5376,N_5233,N_5256);
nand U5377 (N_5377,N_5214,N_5264);
and U5378 (N_5378,N_5218,N_5291);
nor U5379 (N_5379,N_5270,N_5293);
or U5380 (N_5380,N_5267,N_5283);
or U5381 (N_5381,N_5290,N_5257);
xnor U5382 (N_5382,N_5265,N_5288);
and U5383 (N_5383,N_5299,N_5288);
nand U5384 (N_5384,N_5220,N_5272);
xnor U5385 (N_5385,N_5261,N_5260);
or U5386 (N_5386,N_5244,N_5226);
nor U5387 (N_5387,N_5284,N_5299);
nand U5388 (N_5388,N_5250,N_5259);
nor U5389 (N_5389,N_5255,N_5248);
nor U5390 (N_5390,N_5208,N_5284);
nor U5391 (N_5391,N_5202,N_5250);
nand U5392 (N_5392,N_5240,N_5280);
nand U5393 (N_5393,N_5243,N_5274);
xor U5394 (N_5394,N_5212,N_5266);
xor U5395 (N_5395,N_5280,N_5215);
xor U5396 (N_5396,N_5284,N_5278);
xnor U5397 (N_5397,N_5293,N_5259);
nor U5398 (N_5398,N_5269,N_5212);
and U5399 (N_5399,N_5244,N_5205);
xor U5400 (N_5400,N_5388,N_5380);
nor U5401 (N_5401,N_5373,N_5360);
and U5402 (N_5402,N_5311,N_5361);
nand U5403 (N_5403,N_5399,N_5301);
or U5404 (N_5404,N_5332,N_5384);
nand U5405 (N_5405,N_5346,N_5371);
nand U5406 (N_5406,N_5328,N_5302);
and U5407 (N_5407,N_5353,N_5336);
or U5408 (N_5408,N_5350,N_5303);
and U5409 (N_5409,N_5342,N_5349);
nand U5410 (N_5410,N_5321,N_5369);
or U5411 (N_5411,N_5397,N_5306);
nand U5412 (N_5412,N_5318,N_5387);
nor U5413 (N_5413,N_5385,N_5312);
nand U5414 (N_5414,N_5366,N_5313);
xnor U5415 (N_5415,N_5368,N_5338);
or U5416 (N_5416,N_5364,N_5381);
or U5417 (N_5417,N_5314,N_5330);
and U5418 (N_5418,N_5355,N_5395);
nand U5419 (N_5419,N_5370,N_5320);
nand U5420 (N_5420,N_5343,N_5383);
xnor U5421 (N_5421,N_5341,N_5316);
nor U5422 (N_5422,N_5374,N_5365);
nand U5423 (N_5423,N_5304,N_5325);
nor U5424 (N_5424,N_5323,N_5348);
and U5425 (N_5425,N_5386,N_5390);
and U5426 (N_5426,N_5334,N_5398);
nand U5427 (N_5427,N_5372,N_5335);
nand U5428 (N_5428,N_5319,N_5363);
or U5429 (N_5429,N_5367,N_5376);
or U5430 (N_5430,N_5375,N_5307);
nor U5431 (N_5431,N_5392,N_5357);
or U5432 (N_5432,N_5359,N_5305);
and U5433 (N_5433,N_5333,N_5329);
nand U5434 (N_5434,N_5378,N_5331);
nand U5435 (N_5435,N_5310,N_5352);
nor U5436 (N_5436,N_5351,N_5396);
nor U5437 (N_5437,N_5327,N_5326);
xor U5438 (N_5438,N_5344,N_5356);
nand U5439 (N_5439,N_5324,N_5354);
and U5440 (N_5440,N_5322,N_5308);
or U5441 (N_5441,N_5379,N_5347);
xor U5442 (N_5442,N_5309,N_5317);
or U5443 (N_5443,N_5337,N_5340);
xor U5444 (N_5444,N_5300,N_5345);
or U5445 (N_5445,N_5393,N_5377);
nor U5446 (N_5446,N_5339,N_5389);
xor U5447 (N_5447,N_5358,N_5315);
xor U5448 (N_5448,N_5382,N_5394);
nand U5449 (N_5449,N_5391,N_5362);
nand U5450 (N_5450,N_5367,N_5322);
nor U5451 (N_5451,N_5389,N_5312);
xnor U5452 (N_5452,N_5359,N_5339);
nand U5453 (N_5453,N_5349,N_5329);
or U5454 (N_5454,N_5304,N_5361);
xnor U5455 (N_5455,N_5332,N_5369);
nand U5456 (N_5456,N_5308,N_5329);
nand U5457 (N_5457,N_5382,N_5340);
xnor U5458 (N_5458,N_5366,N_5325);
xnor U5459 (N_5459,N_5327,N_5339);
and U5460 (N_5460,N_5327,N_5375);
xnor U5461 (N_5461,N_5316,N_5354);
or U5462 (N_5462,N_5377,N_5383);
xnor U5463 (N_5463,N_5321,N_5333);
or U5464 (N_5464,N_5395,N_5386);
nor U5465 (N_5465,N_5308,N_5390);
nor U5466 (N_5466,N_5374,N_5371);
nand U5467 (N_5467,N_5330,N_5308);
and U5468 (N_5468,N_5357,N_5395);
nor U5469 (N_5469,N_5355,N_5381);
or U5470 (N_5470,N_5325,N_5383);
nor U5471 (N_5471,N_5327,N_5341);
or U5472 (N_5472,N_5320,N_5356);
xnor U5473 (N_5473,N_5306,N_5367);
and U5474 (N_5474,N_5306,N_5369);
and U5475 (N_5475,N_5327,N_5385);
xnor U5476 (N_5476,N_5358,N_5354);
or U5477 (N_5477,N_5388,N_5305);
nand U5478 (N_5478,N_5351,N_5304);
nor U5479 (N_5479,N_5336,N_5343);
or U5480 (N_5480,N_5312,N_5353);
and U5481 (N_5481,N_5360,N_5320);
nor U5482 (N_5482,N_5355,N_5385);
nor U5483 (N_5483,N_5391,N_5358);
nand U5484 (N_5484,N_5348,N_5320);
nor U5485 (N_5485,N_5399,N_5315);
xnor U5486 (N_5486,N_5369,N_5361);
nand U5487 (N_5487,N_5377,N_5394);
or U5488 (N_5488,N_5315,N_5309);
xnor U5489 (N_5489,N_5398,N_5365);
xnor U5490 (N_5490,N_5392,N_5340);
nor U5491 (N_5491,N_5353,N_5397);
and U5492 (N_5492,N_5341,N_5372);
or U5493 (N_5493,N_5308,N_5348);
or U5494 (N_5494,N_5329,N_5371);
xnor U5495 (N_5495,N_5330,N_5361);
nor U5496 (N_5496,N_5379,N_5338);
nor U5497 (N_5497,N_5309,N_5313);
nor U5498 (N_5498,N_5330,N_5335);
and U5499 (N_5499,N_5354,N_5379);
xor U5500 (N_5500,N_5459,N_5493);
and U5501 (N_5501,N_5427,N_5436);
or U5502 (N_5502,N_5421,N_5444);
or U5503 (N_5503,N_5453,N_5475);
xor U5504 (N_5504,N_5490,N_5413);
and U5505 (N_5505,N_5462,N_5423);
nor U5506 (N_5506,N_5476,N_5430);
and U5507 (N_5507,N_5495,N_5412);
nor U5508 (N_5508,N_5466,N_5420);
xnor U5509 (N_5509,N_5410,N_5446);
nor U5510 (N_5510,N_5415,N_5422);
nor U5511 (N_5511,N_5404,N_5431);
xor U5512 (N_5512,N_5408,N_5473);
nor U5513 (N_5513,N_5451,N_5479);
and U5514 (N_5514,N_5460,N_5488);
xor U5515 (N_5515,N_5440,N_5449);
xor U5516 (N_5516,N_5491,N_5492);
and U5517 (N_5517,N_5458,N_5435);
nand U5518 (N_5518,N_5499,N_5401);
xnor U5519 (N_5519,N_5437,N_5487);
and U5520 (N_5520,N_5472,N_5405);
nor U5521 (N_5521,N_5496,N_5433);
or U5522 (N_5522,N_5418,N_5474);
and U5523 (N_5523,N_5483,N_5402);
nor U5524 (N_5524,N_5447,N_5455);
nor U5525 (N_5525,N_5419,N_5463);
nor U5526 (N_5526,N_5461,N_5406);
xor U5527 (N_5527,N_5478,N_5457);
or U5528 (N_5528,N_5480,N_5482);
and U5529 (N_5529,N_5400,N_5417);
xnor U5530 (N_5530,N_5425,N_5416);
or U5531 (N_5531,N_5469,N_5494);
xnor U5532 (N_5532,N_5443,N_5407);
or U5533 (N_5533,N_5414,N_5434);
nand U5534 (N_5534,N_5429,N_5454);
xor U5535 (N_5535,N_5403,N_5409);
nor U5536 (N_5536,N_5438,N_5486);
xor U5537 (N_5537,N_5497,N_5426);
and U5538 (N_5538,N_5470,N_5464);
xnor U5539 (N_5539,N_5428,N_5471);
and U5540 (N_5540,N_5441,N_5477);
or U5541 (N_5541,N_5456,N_5481);
or U5542 (N_5542,N_5485,N_5442);
nor U5543 (N_5543,N_5498,N_5439);
xor U5544 (N_5544,N_5411,N_5445);
nand U5545 (N_5545,N_5448,N_5489);
xnor U5546 (N_5546,N_5484,N_5432);
nand U5547 (N_5547,N_5450,N_5424);
nor U5548 (N_5548,N_5452,N_5468);
or U5549 (N_5549,N_5465,N_5467);
and U5550 (N_5550,N_5477,N_5494);
xor U5551 (N_5551,N_5462,N_5403);
xnor U5552 (N_5552,N_5401,N_5445);
nor U5553 (N_5553,N_5461,N_5403);
xor U5554 (N_5554,N_5477,N_5476);
xnor U5555 (N_5555,N_5498,N_5431);
and U5556 (N_5556,N_5454,N_5441);
or U5557 (N_5557,N_5427,N_5402);
and U5558 (N_5558,N_5456,N_5421);
and U5559 (N_5559,N_5497,N_5400);
and U5560 (N_5560,N_5402,N_5410);
xnor U5561 (N_5561,N_5476,N_5495);
nand U5562 (N_5562,N_5487,N_5475);
xnor U5563 (N_5563,N_5400,N_5495);
and U5564 (N_5564,N_5427,N_5481);
xor U5565 (N_5565,N_5423,N_5434);
xnor U5566 (N_5566,N_5491,N_5451);
nand U5567 (N_5567,N_5422,N_5410);
xnor U5568 (N_5568,N_5418,N_5406);
nand U5569 (N_5569,N_5473,N_5430);
xor U5570 (N_5570,N_5459,N_5482);
nor U5571 (N_5571,N_5479,N_5489);
nor U5572 (N_5572,N_5455,N_5478);
nand U5573 (N_5573,N_5472,N_5473);
nand U5574 (N_5574,N_5417,N_5495);
or U5575 (N_5575,N_5479,N_5403);
xnor U5576 (N_5576,N_5495,N_5420);
and U5577 (N_5577,N_5493,N_5407);
and U5578 (N_5578,N_5401,N_5427);
and U5579 (N_5579,N_5454,N_5497);
and U5580 (N_5580,N_5400,N_5412);
xor U5581 (N_5581,N_5484,N_5401);
and U5582 (N_5582,N_5411,N_5401);
xor U5583 (N_5583,N_5408,N_5417);
nand U5584 (N_5584,N_5402,N_5456);
xnor U5585 (N_5585,N_5461,N_5436);
nand U5586 (N_5586,N_5430,N_5414);
and U5587 (N_5587,N_5417,N_5469);
and U5588 (N_5588,N_5426,N_5491);
nor U5589 (N_5589,N_5441,N_5436);
nand U5590 (N_5590,N_5416,N_5480);
xnor U5591 (N_5591,N_5406,N_5499);
nand U5592 (N_5592,N_5416,N_5469);
xnor U5593 (N_5593,N_5492,N_5499);
and U5594 (N_5594,N_5499,N_5467);
and U5595 (N_5595,N_5407,N_5473);
nand U5596 (N_5596,N_5494,N_5493);
and U5597 (N_5597,N_5415,N_5416);
nand U5598 (N_5598,N_5435,N_5410);
nand U5599 (N_5599,N_5450,N_5418);
nor U5600 (N_5600,N_5538,N_5525);
and U5601 (N_5601,N_5575,N_5522);
and U5602 (N_5602,N_5570,N_5577);
nand U5603 (N_5603,N_5580,N_5579);
and U5604 (N_5604,N_5598,N_5550);
xnor U5605 (N_5605,N_5533,N_5590);
nand U5606 (N_5606,N_5591,N_5541);
nor U5607 (N_5607,N_5514,N_5558);
nand U5608 (N_5608,N_5542,N_5516);
nand U5609 (N_5609,N_5500,N_5544);
nand U5610 (N_5610,N_5594,N_5546);
nor U5611 (N_5611,N_5583,N_5555);
xnor U5612 (N_5612,N_5597,N_5585);
or U5613 (N_5613,N_5534,N_5552);
xnor U5614 (N_5614,N_5578,N_5586);
or U5615 (N_5615,N_5537,N_5561);
nor U5616 (N_5616,N_5510,N_5504);
nor U5617 (N_5617,N_5564,N_5571);
xor U5618 (N_5618,N_5569,N_5536);
xor U5619 (N_5619,N_5519,N_5560);
nand U5620 (N_5620,N_5506,N_5524);
and U5621 (N_5621,N_5513,N_5566);
nand U5622 (N_5622,N_5572,N_5521);
and U5623 (N_5623,N_5501,N_5547);
xor U5624 (N_5624,N_5589,N_5503);
nand U5625 (N_5625,N_5502,N_5512);
and U5626 (N_5626,N_5554,N_5557);
nand U5627 (N_5627,N_5532,N_5520);
or U5628 (N_5628,N_5539,N_5528);
and U5629 (N_5629,N_5595,N_5596);
nor U5630 (N_5630,N_5530,N_5556);
and U5631 (N_5631,N_5548,N_5584);
nand U5632 (N_5632,N_5518,N_5573);
or U5633 (N_5633,N_5587,N_5545);
and U5634 (N_5634,N_5553,N_5515);
nor U5635 (N_5635,N_5531,N_5517);
nor U5636 (N_5636,N_5527,N_5523);
nand U5637 (N_5637,N_5582,N_5551);
and U5638 (N_5638,N_5592,N_5563);
xnor U5639 (N_5639,N_5535,N_5511);
xnor U5640 (N_5640,N_5599,N_5559);
nand U5641 (N_5641,N_5567,N_5526);
or U5642 (N_5642,N_5529,N_5549);
and U5643 (N_5643,N_5568,N_5505);
nand U5644 (N_5644,N_5543,N_5508);
and U5645 (N_5645,N_5565,N_5540);
nand U5646 (N_5646,N_5574,N_5509);
xor U5647 (N_5647,N_5581,N_5562);
and U5648 (N_5648,N_5507,N_5576);
xnor U5649 (N_5649,N_5593,N_5588);
or U5650 (N_5650,N_5597,N_5506);
xnor U5651 (N_5651,N_5557,N_5539);
and U5652 (N_5652,N_5589,N_5552);
xor U5653 (N_5653,N_5555,N_5523);
nor U5654 (N_5654,N_5538,N_5507);
nor U5655 (N_5655,N_5531,N_5565);
nand U5656 (N_5656,N_5589,N_5579);
xor U5657 (N_5657,N_5546,N_5581);
and U5658 (N_5658,N_5597,N_5583);
nor U5659 (N_5659,N_5569,N_5509);
nand U5660 (N_5660,N_5575,N_5512);
xor U5661 (N_5661,N_5591,N_5514);
xnor U5662 (N_5662,N_5574,N_5531);
or U5663 (N_5663,N_5516,N_5559);
or U5664 (N_5664,N_5548,N_5536);
or U5665 (N_5665,N_5539,N_5532);
nand U5666 (N_5666,N_5556,N_5578);
xor U5667 (N_5667,N_5518,N_5574);
and U5668 (N_5668,N_5527,N_5588);
nand U5669 (N_5669,N_5572,N_5502);
nor U5670 (N_5670,N_5576,N_5592);
and U5671 (N_5671,N_5537,N_5566);
or U5672 (N_5672,N_5599,N_5596);
or U5673 (N_5673,N_5538,N_5595);
or U5674 (N_5674,N_5521,N_5533);
and U5675 (N_5675,N_5501,N_5535);
nand U5676 (N_5676,N_5588,N_5540);
or U5677 (N_5677,N_5575,N_5585);
nor U5678 (N_5678,N_5541,N_5512);
or U5679 (N_5679,N_5569,N_5581);
nor U5680 (N_5680,N_5501,N_5595);
nand U5681 (N_5681,N_5545,N_5522);
xor U5682 (N_5682,N_5594,N_5576);
and U5683 (N_5683,N_5584,N_5557);
nand U5684 (N_5684,N_5514,N_5590);
nor U5685 (N_5685,N_5512,N_5576);
nand U5686 (N_5686,N_5557,N_5573);
xor U5687 (N_5687,N_5555,N_5501);
nand U5688 (N_5688,N_5520,N_5595);
or U5689 (N_5689,N_5524,N_5582);
nor U5690 (N_5690,N_5538,N_5571);
or U5691 (N_5691,N_5590,N_5548);
nand U5692 (N_5692,N_5595,N_5552);
and U5693 (N_5693,N_5516,N_5549);
nand U5694 (N_5694,N_5503,N_5526);
and U5695 (N_5695,N_5550,N_5519);
and U5696 (N_5696,N_5586,N_5502);
nand U5697 (N_5697,N_5541,N_5548);
nand U5698 (N_5698,N_5549,N_5515);
nand U5699 (N_5699,N_5536,N_5511);
or U5700 (N_5700,N_5670,N_5658);
or U5701 (N_5701,N_5694,N_5675);
nor U5702 (N_5702,N_5685,N_5653);
xnor U5703 (N_5703,N_5639,N_5635);
nor U5704 (N_5704,N_5609,N_5693);
and U5705 (N_5705,N_5610,N_5611);
nor U5706 (N_5706,N_5679,N_5606);
xnor U5707 (N_5707,N_5651,N_5664);
nor U5708 (N_5708,N_5631,N_5607);
or U5709 (N_5709,N_5601,N_5605);
and U5710 (N_5710,N_5627,N_5663);
and U5711 (N_5711,N_5613,N_5689);
nand U5712 (N_5712,N_5608,N_5640);
nor U5713 (N_5713,N_5665,N_5686);
or U5714 (N_5714,N_5682,N_5646);
nor U5715 (N_5715,N_5697,N_5695);
nand U5716 (N_5716,N_5677,N_5662);
xor U5717 (N_5717,N_5621,N_5661);
and U5718 (N_5718,N_5644,N_5643);
nor U5719 (N_5719,N_5623,N_5692);
nand U5720 (N_5720,N_5614,N_5668);
nand U5721 (N_5721,N_5654,N_5622);
nor U5722 (N_5722,N_5647,N_5612);
and U5723 (N_5723,N_5688,N_5600);
nand U5724 (N_5724,N_5669,N_5656);
nor U5725 (N_5725,N_5674,N_5659);
xor U5726 (N_5726,N_5642,N_5696);
xnor U5727 (N_5727,N_5626,N_5676);
nand U5728 (N_5728,N_5618,N_5660);
nand U5729 (N_5729,N_5615,N_5624);
nand U5730 (N_5730,N_5684,N_5671);
nand U5731 (N_5731,N_5617,N_5690);
nand U5732 (N_5732,N_5634,N_5632);
nand U5733 (N_5733,N_5681,N_5699);
xnor U5734 (N_5734,N_5625,N_5667);
or U5735 (N_5735,N_5648,N_5604);
xor U5736 (N_5736,N_5691,N_5619);
or U5737 (N_5737,N_5616,N_5630);
nand U5738 (N_5738,N_5698,N_5678);
nor U5739 (N_5739,N_5680,N_5641);
or U5740 (N_5740,N_5649,N_5620);
and U5741 (N_5741,N_5603,N_5655);
or U5742 (N_5742,N_5636,N_5637);
nor U5743 (N_5743,N_5629,N_5687);
nor U5744 (N_5744,N_5683,N_5673);
nand U5745 (N_5745,N_5633,N_5638);
and U5746 (N_5746,N_5650,N_5652);
xnor U5747 (N_5747,N_5657,N_5645);
xnor U5748 (N_5748,N_5628,N_5602);
xor U5749 (N_5749,N_5666,N_5672);
xnor U5750 (N_5750,N_5658,N_5617);
nor U5751 (N_5751,N_5659,N_5646);
xnor U5752 (N_5752,N_5691,N_5679);
nor U5753 (N_5753,N_5691,N_5614);
nor U5754 (N_5754,N_5680,N_5670);
nor U5755 (N_5755,N_5633,N_5698);
nor U5756 (N_5756,N_5603,N_5648);
nor U5757 (N_5757,N_5677,N_5679);
or U5758 (N_5758,N_5651,N_5618);
xnor U5759 (N_5759,N_5616,N_5637);
nand U5760 (N_5760,N_5602,N_5675);
nand U5761 (N_5761,N_5676,N_5695);
xnor U5762 (N_5762,N_5639,N_5664);
nor U5763 (N_5763,N_5667,N_5645);
or U5764 (N_5764,N_5618,N_5607);
nor U5765 (N_5765,N_5673,N_5697);
or U5766 (N_5766,N_5609,N_5608);
and U5767 (N_5767,N_5639,N_5649);
xor U5768 (N_5768,N_5655,N_5604);
and U5769 (N_5769,N_5683,N_5604);
and U5770 (N_5770,N_5662,N_5634);
or U5771 (N_5771,N_5618,N_5650);
nor U5772 (N_5772,N_5679,N_5663);
or U5773 (N_5773,N_5675,N_5684);
and U5774 (N_5774,N_5670,N_5697);
xnor U5775 (N_5775,N_5624,N_5677);
and U5776 (N_5776,N_5695,N_5689);
nand U5777 (N_5777,N_5618,N_5628);
or U5778 (N_5778,N_5658,N_5601);
nand U5779 (N_5779,N_5615,N_5617);
nor U5780 (N_5780,N_5613,N_5624);
and U5781 (N_5781,N_5644,N_5693);
nor U5782 (N_5782,N_5613,N_5664);
nand U5783 (N_5783,N_5629,N_5683);
xor U5784 (N_5784,N_5605,N_5697);
nor U5785 (N_5785,N_5617,N_5691);
or U5786 (N_5786,N_5648,N_5657);
or U5787 (N_5787,N_5660,N_5642);
and U5788 (N_5788,N_5669,N_5646);
nand U5789 (N_5789,N_5670,N_5619);
xnor U5790 (N_5790,N_5616,N_5695);
nand U5791 (N_5791,N_5610,N_5613);
nor U5792 (N_5792,N_5693,N_5653);
xor U5793 (N_5793,N_5671,N_5641);
or U5794 (N_5794,N_5658,N_5695);
nor U5795 (N_5795,N_5676,N_5649);
nand U5796 (N_5796,N_5669,N_5635);
nand U5797 (N_5797,N_5655,N_5602);
or U5798 (N_5798,N_5695,N_5625);
and U5799 (N_5799,N_5689,N_5694);
xor U5800 (N_5800,N_5708,N_5728);
xor U5801 (N_5801,N_5754,N_5777);
or U5802 (N_5802,N_5714,N_5742);
xnor U5803 (N_5803,N_5776,N_5747);
nand U5804 (N_5804,N_5784,N_5718);
nand U5805 (N_5805,N_5797,N_5722);
nand U5806 (N_5806,N_5798,N_5727);
or U5807 (N_5807,N_5774,N_5756);
xnor U5808 (N_5808,N_5703,N_5790);
nand U5809 (N_5809,N_5759,N_5702);
nand U5810 (N_5810,N_5796,N_5701);
and U5811 (N_5811,N_5766,N_5710);
xnor U5812 (N_5812,N_5734,N_5721);
and U5813 (N_5813,N_5749,N_5735);
and U5814 (N_5814,N_5786,N_5723);
nand U5815 (N_5815,N_5724,N_5771);
and U5816 (N_5816,N_5799,N_5720);
xor U5817 (N_5817,N_5711,N_5795);
nand U5818 (N_5818,N_5741,N_5707);
and U5819 (N_5819,N_5764,N_5767);
nand U5820 (N_5820,N_5794,N_5744);
nand U5821 (N_5821,N_5713,N_5789);
xnor U5822 (N_5822,N_5730,N_5748);
and U5823 (N_5823,N_5740,N_5715);
or U5824 (N_5824,N_5733,N_5763);
or U5825 (N_5825,N_5751,N_5750);
nor U5826 (N_5826,N_5785,N_5792);
nor U5827 (N_5827,N_5773,N_5743);
nor U5828 (N_5828,N_5769,N_5726);
nor U5829 (N_5829,N_5717,N_5768);
xor U5830 (N_5830,N_5752,N_5782);
or U5831 (N_5831,N_5762,N_5775);
nand U5832 (N_5832,N_5746,N_5739);
xnor U5833 (N_5833,N_5712,N_5706);
nor U5834 (N_5834,N_5791,N_5729);
xnor U5835 (N_5835,N_5705,N_5793);
or U5836 (N_5836,N_5781,N_5787);
nor U5837 (N_5837,N_5745,N_5716);
nor U5838 (N_5838,N_5731,N_5778);
xor U5839 (N_5839,N_5737,N_5755);
or U5840 (N_5840,N_5779,N_5736);
or U5841 (N_5841,N_5783,N_5761);
and U5842 (N_5842,N_5738,N_5700);
xor U5843 (N_5843,N_5788,N_5757);
xnor U5844 (N_5844,N_5772,N_5709);
xor U5845 (N_5845,N_5725,N_5704);
xnor U5846 (N_5846,N_5770,N_5765);
nor U5847 (N_5847,N_5719,N_5780);
and U5848 (N_5848,N_5753,N_5758);
nand U5849 (N_5849,N_5732,N_5760);
and U5850 (N_5850,N_5776,N_5726);
nand U5851 (N_5851,N_5713,N_5704);
nor U5852 (N_5852,N_5727,N_5712);
xnor U5853 (N_5853,N_5784,N_5751);
xor U5854 (N_5854,N_5776,N_5715);
nor U5855 (N_5855,N_5757,N_5701);
and U5856 (N_5856,N_5719,N_5702);
nand U5857 (N_5857,N_5720,N_5727);
or U5858 (N_5858,N_5786,N_5783);
nand U5859 (N_5859,N_5784,N_5782);
or U5860 (N_5860,N_5779,N_5757);
and U5861 (N_5861,N_5725,N_5791);
or U5862 (N_5862,N_5733,N_5741);
nor U5863 (N_5863,N_5752,N_5798);
or U5864 (N_5864,N_5764,N_5756);
nor U5865 (N_5865,N_5777,N_5749);
xor U5866 (N_5866,N_5796,N_5774);
nand U5867 (N_5867,N_5724,N_5703);
nand U5868 (N_5868,N_5719,N_5736);
nor U5869 (N_5869,N_5785,N_5712);
xnor U5870 (N_5870,N_5741,N_5754);
xor U5871 (N_5871,N_5760,N_5750);
xnor U5872 (N_5872,N_5733,N_5794);
or U5873 (N_5873,N_5700,N_5795);
and U5874 (N_5874,N_5745,N_5790);
xnor U5875 (N_5875,N_5774,N_5763);
nor U5876 (N_5876,N_5760,N_5757);
and U5877 (N_5877,N_5759,N_5782);
and U5878 (N_5878,N_5768,N_5704);
or U5879 (N_5879,N_5701,N_5793);
or U5880 (N_5880,N_5757,N_5700);
nor U5881 (N_5881,N_5792,N_5702);
and U5882 (N_5882,N_5792,N_5774);
nand U5883 (N_5883,N_5701,N_5781);
or U5884 (N_5884,N_5713,N_5717);
nor U5885 (N_5885,N_5714,N_5753);
and U5886 (N_5886,N_5788,N_5786);
and U5887 (N_5887,N_5744,N_5793);
and U5888 (N_5888,N_5780,N_5755);
nor U5889 (N_5889,N_5702,N_5710);
or U5890 (N_5890,N_5758,N_5741);
nor U5891 (N_5891,N_5738,N_5778);
nor U5892 (N_5892,N_5760,N_5799);
and U5893 (N_5893,N_5758,N_5701);
and U5894 (N_5894,N_5714,N_5730);
nor U5895 (N_5895,N_5781,N_5727);
nor U5896 (N_5896,N_5719,N_5784);
xor U5897 (N_5897,N_5784,N_5736);
or U5898 (N_5898,N_5789,N_5747);
nand U5899 (N_5899,N_5735,N_5788);
nand U5900 (N_5900,N_5827,N_5896);
or U5901 (N_5901,N_5812,N_5899);
or U5902 (N_5902,N_5857,N_5852);
or U5903 (N_5903,N_5887,N_5847);
nand U5904 (N_5904,N_5860,N_5830);
or U5905 (N_5905,N_5844,N_5819);
nor U5906 (N_5906,N_5892,N_5856);
nand U5907 (N_5907,N_5880,N_5806);
nand U5908 (N_5908,N_5837,N_5802);
and U5909 (N_5909,N_5842,N_5850);
nand U5910 (N_5910,N_5883,N_5890);
nand U5911 (N_5911,N_5831,N_5813);
nor U5912 (N_5912,N_5836,N_5851);
nor U5913 (N_5913,N_5833,N_5893);
and U5914 (N_5914,N_5849,N_5826);
xnor U5915 (N_5915,N_5810,N_5804);
nor U5916 (N_5916,N_5858,N_5828);
nor U5917 (N_5917,N_5863,N_5895);
nand U5918 (N_5918,N_5861,N_5821);
xnor U5919 (N_5919,N_5815,N_5838);
xor U5920 (N_5920,N_5877,N_5801);
nor U5921 (N_5921,N_5878,N_5888);
nand U5922 (N_5922,N_5848,N_5834);
or U5923 (N_5923,N_5839,N_5800);
and U5924 (N_5924,N_5872,N_5884);
nand U5925 (N_5925,N_5886,N_5823);
and U5926 (N_5926,N_5843,N_5853);
or U5927 (N_5927,N_5862,N_5845);
or U5928 (N_5928,N_5889,N_5879);
nor U5929 (N_5929,N_5809,N_5820);
xnor U5930 (N_5930,N_5816,N_5868);
nand U5931 (N_5931,N_5885,N_5841);
or U5932 (N_5932,N_5866,N_5835);
and U5933 (N_5933,N_5891,N_5807);
nand U5934 (N_5934,N_5829,N_5867);
xnor U5935 (N_5935,N_5811,N_5869);
and U5936 (N_5936,N_5855,N_5873);
or U5937 (N_5937,N_5874,N_5894);
nand U5938 (N_5938,N_5870,N_5897);
nor U5939 (N_5939,N_5898,N_5825);
or U5940 (N_5940,N_5824,N_5859);
or U5941 (N_5941,N_5846,N_5881);
or U5942 (N_5942,N_5808,N_5875);
or U5943 (N_5943,N_5818,N_5840);
and U5944 (N_5944,N_5805,N_5817);
xnor U5945 (N_5945,N_5832,N_5876);
nand U5946 (N_5946,N_5864,N_5822);
or U5947 (N_5947,N_5865,N_5814);
and U5948 (N_5948,N_5882,N_5871);
nor U5949 (N_5949,N_5854,N_5803);
nand U5950 (N_5950,N_5895,N_5889);
nor U5951 (N_5951,N_5822,N_5873);
xor U5952 (N_5952,N_5830,N_5804);
xor U5953 (N_5953,N_5839,N_5822);
nand U5954 (N_5954,N_5828,N_5881);
xnor U5955 (N_5955,N_5829,N_5888);
and U5956 (N_5956,N_5861,N_5856);
nand U5957 (N_5957,N_5804,N_5802);
nor U5958 (N_5958,N_5878,N_5841);
and U5959 (N_5959,N_5865,N_5894);
xor U5960 (N_5960,N_5827,N_5821);
or U5961 (N_5961,N_5852,N_5856);
xnor U5962 (N_5962,N_5867,N_5819);
xnor U5963 (N_5963,N_5861,N_5858);
and U5964 (N_5964,N_5880,N_5832);
xnor U5965 (N_5965,N_5887,N_5890);
xnor U5966 (N_5966,N_5835,N_5865);
xnor U5967 (N_5967,N_5890,N_5840);
xor U5968 (N_5968,N_5843,N_5855);
xor U5969 (N_5969,N_5838,N_5899);
xor U5970 (N_5970,N_5803,N_5820);
xnor U5971 (N_5971,N_5849,N_5887);
nor U5972 (N_5972,N_5859,N_5838);
xor U5973 (N_5973,N_5851,N_5868);
nand U5974 (N_5974,N_5844,N_5885);
xnor U5975 (N_5975,N_5839,N_5814);
nand U5976 (N_5976,N_5850,N_5836);
xnor U5977 (N_5977,N_5831,N_5832);
nor U5978 (N_5978,N_5868,N_5884);
and U5979 (N_5979,N_5830,N_5884);
and U5980 (N_5980,N_5846,N_5865);
and U5981 (N_5981,N_5823,N_5812);
or U5982 (N_5982,N_5829,N_5809);
nand U5983 (N_5983,N_5857,N_5816);
nor U5984 (N_5984,N_5831,N_5848);
or U5985 (N_5985,N_5831,N_5893);
xor U5986 (N_5986,N_5806,N_5858);
or U5987 (N_5987,N_5816,N_5856);
nor U5988 (N_5988,N_5801,N_5827);
xor U5989 (N_5989,N_5875,N_5800);
nor U5990 (N_5990,N_5871,N_5844);
and U5991 (N_5991,N_5832,N_5853);
nor U5992 (N_5992,N_5823,N_5849);
nor U5993 (N_5993,N_5838,N_5823);
xor U5994 (N_5994,N_5855,N_5881);
nor U5995 (N_5995,N_5899,N_5841);
or U5996 (N_5996,N_5815,N_5836);
or U5997 (N_5997,N_5857,N_5825);
xnor U5998 (N_5998,N_5828,N_5804);
and U5999 (N_5999,N_5886,N_5844);
xnor U6000 (N_6000,N_5959,N_5916);
nand U6001 (N_6001,N_5963,N_5902);
and U6002 (N_6002,N_5908,N_5962);
xor U6003 (N_6003,N_5945,N_5986);
nand U6004 (N_6004,N_5942,N_5967);
and U6005 (N_6005,N_5964,N_5985);
nand U6006 (N_6006,N_5936,N_5991);
nor U6007 (N_6007,N_5988,N_5981);
xnor U6008 (N_6008,N_5927,N_5955);
nand U6009 (N_6009,N_5903,N_5953);
nand U6010 (N_6010,N_5989,N_5934);
nor U6011 (N_6011,N_5925,N_5919);
or U6012 (N_6012,N_5971,N_5939);
nor U6013 (N_6013,N_5998,N_5920);
or U6014 (N_6014,N_5935,N_5928);
nor U6015 (N_6015,N_5976,N_5948);
nand U6016 (N_6016,N_5924,N_5979);
or U6017 (N_6017,N_5907,N_5904);
nand U6018 (N_6018,N_5956,N_5906);
nor U6019 (N_6019,N_5926,N_5983);
and U6020 (N_6020,N_5980,N_5987);
xnor U6021 (N_6021,N_5997,N_5958);
nand U6022 (N_6022,N_5933,N_5930);
xnor U6023 (N_6023,N_5912,N_5937);
nand U6024 (N_6024,N_5960,N_5909);
or U6025 (N_6025,N_5946,N_5961);
nand U6026 (N_6026,N_5978,N_5992);
nand U6027 (N_6027,N_5974,N_5913);
and U6028 (N_6028,N_5995,N_5921);
nor U6029 (N_6029,N_5957,N_5918);
nand U6030 (N_6030,N_5922,N_5990);
xnor U6031 (N_6031,N_5905,N_5943);
nand U6032 (N_6032,N_5966,N_5917);
nand U6033 (N_6033,N_5910,N_5914);
nand U6034 (N_6034,N_5947,N_5901);
or U6035 (N_6035,N_5940,N_5975);
xnor U6036 (N_6036,N_5977,N_5996);
nor U6037 (N_6037,N_5929,N_5915);
nand U6038 (N_6038,N_5951,N_5941);
xnor U6039 (N_6039,N_5932,N_5931);
and U6040 (N_6040,N_5984,N_5994);
or U6041 (N_6041,N_5973,N_5938);
or U6042 (N_6042,N_5923,N_5949);
xnor U6043 (N_6043,N_5950,N_5952);
nor U6044 (N_6044,N_5954,N_5900);
and U6045 (N_6045,N_5968,N_5969);
or U6046 (N_6046,N_5965,N_5993);
nand U6047 (N_6047,N_5972,N_5944);
and U6048 (N_6048,N_5999,N_5970);
xor U6049 (N_6049,N_5982,N_5911);
xor U6050 (N_6050,N_5942,N_5957);
xor U6051 (N_6051,N_5960,N_5965);
xor U6052 (N_6052,N_5983,N_5922);
and U6053 (N_6053,N_5911,N_5913);
nor U6054 (N_6054,N_5990,N_5975);
or U6055 (N_6055,N_5917,N_5901);
nand U6056 (N_6056,N_5988,N_5906);
and U6057 (N_6057,N_5919,N_5952);
xor U6058 (N_6058,N_5922,N_5915);
or U6059 (N_6059,N_5992,N_5958);
xnor U6060 (N_6060,N_5946,N_5919);
and U6061 (N_6061,N_5913,N_5945);
and U6062 (N_6062,N_5955,N_5962);
nor U6063 (N_6063,N_5931,N_5974);
and U6064 (N_6064,N_5935,N_5994);
nor U6065 (N_6065,N_5940,N_5980);
and U6066 (N_6066,N_5916,N_5987);
nand U6067 (N_6067,N_5974,N_5907);
nand U6068 (N_6068,N_5998,N_5959);
nand U6069 (N_6069,N_5908,N_5905);
xnor U6070 (N_6070,N_5993,N_5964);
and U6071 (N_6071,N_5950,N_5963);
nor U6072 (N_6072,N_5968,N_5990);
or U6073 (N_6073,N_5933,N_5965);
and U6074 (N_6074,N_5930,N_5974);
nor U6075 (N_6075,N_5921,N_5936);
nor U6076 (N_6076,N_5958,N_5982);
or U6077 (N_6077,N_5962,N_5913);
nand U6078 (N_6078,N_5989,N_5901);
or U6079 (N_6079,N_5988,N_5947);
nand U6080 (N_6080,N_5950,N_5911);
nand U6081 (N_6081,N_5906,N_5975);
or U6082 (N_6082,N_5967,N_5911);
nand U6083 (N_6083,N_5913,N_5966);
nand U6084 (N_6084,N_5923,N_5972);
or U6085 (N_6085,N_5909,N_5925);
xnor U6086 (N_6086,N_5957,N_5979);
or U6087 (N_6087,N_5954,N_5971);
nor U6088 (N_6088,N_5997,N_5950);
or U6089 (N_6089,N_5937,N_5995);
xor U6090 (N_6090,N_5903,N_5949);
nand U6091 (N_6091,N_5902,N_5927);
xnor U6092 (N_6092,N_5900,N_5940);
or U6093 (N_6093,N_5908,N_5974);
or U6094 (N_6094,N_5958,N_5978);
and U6095 (N_6095,N_5987,N_5962);
nand U6096 (N_6096,N_5944,N_5906);
nor U6097 (N_6097,N_5963,N_5913);
or U6098 (N_6098,N_5985,N_5925);
xor U6099 (N_6099,N_5995,N_5980);
nand U6100 (N_6100,N_6088,N_6029);
nand U6101 (N_6101,N_6081,N_6043);
xnor U6102 (N_6102,N_6011,N_6074);
xor U6103 (N_6103,N_6060,N_6001);
nor U6104 (N_6104,N_6061,N_6097);
or U6105 (N_6105,N_6030,N_6004);
nand U6106 (N_6106,N_6027,N_6048);
or U6107 (N_6107,N_6069,N_6058);
nand U6108 (N_6108,N_6094,N_6067);
or U6109 (N_6109,N_6023,N_6035);
nor U6110 (N_6110,N_6072,N_6024);
nand U6111 (N_6111,N_6092,N_6098);
xor U6112 (N_6112,N_6066,N_6078);
nand U6113 (N_6113,N_6087,N_6070);
and U6114 (N_6114,N_6041,N_6083);
or U6115 (N_6115,N_6017,N_6054);
or U6116 (N_6116,N_6019,N_6089);
and U6117 (N_6117,N_6002,N_6042);
and U6118 (N_6118,N_6051,N_6018);
or U6119 (N_6119,N_6044,N_6085);
nor U6120 (N_6120,N_6059,N_6084);
nor U6121 (N_6121,N_6033,N_6090);
or U6122 (N_6122,N_6080,N_6010);
nand U6123 (N_6123,N_6093,N_6031);
or U6124 (N_6124,N_6038,N_6049);
xnor U6125 (N_6125,N_6037,N_6056);
nand U6126 (N_6126,N_6071,N_6028);
xor U6127 (N_6127,N_6040,N_6065);
xnor U6128 (N_6128,N_6021,N_6022);
or U6129 (N_6129,N_6005,N_6036);
nor U6130 (N_6130,N_6077,N_6099);
and U6131 (N_6131,N_6075,N_6008);
nor U6132 (N_6132,N_6034,N_6046);
nor U6133 (N_6133,N_6076,N_6032);
and U6134 (N_6134,N_6007,N_6073);
and U6135 (N_6135,N_6013,N_6068);
nor U6136 (N_6136,N_6009,N_6095);
nand U6137 (N_6137,N_6047,N_6082);
or U6138 (N_6138,N_6015,N_6016);
and U6139 (N_6139,N_6063,N_6006);
or U6140 (N_6140,N_6000,N_6014);
xor U6141 (N_6141,N_6012,N_6055);
and U6142 (N_6142,N_6053,N_6039);
or U6143 (N_6143,N_6050,N_6045);
and U6144 (N_6144,N_6057,N_6026);
and U6145 (N_6145,N_6086,N_6003);
xor U6146 (N_6146,N_6096,N_6025);
xnor U6147 (N_6147,N_6079,N_6020);
and U6148 (N_6148,N_6064,N_6052);
or U6149 (N_6149,N_6091,N_6062);
xor U6150 (N_6150,N_6074,N_6061);
nor U6151 (N_6151,N_6085,N_6056);
nand U6152 (N_6152,N_6004,N_6038);
xor U6153 (N_6153,N_6022,N_6090);
nor U6154 (N_6154,N_6051,N_6064);
nand U6155 (N_6155,N_6032,N_6036);
xor U6156 (N_6156,N_6045,N_6085);
nand U6157 (N_6157,N_6010,N_6090);
nor U6158 (N_6158,N_6042,N_6035);
nand U6159 (N_6159,N_6069,N_6057);
nand U6160 (N_6160,N_6048,N_6058);
or U6161 (N_6161,N_6049,N_6082);
or U6162 (N_6162,N_6088,N_6050);
nor U6163 (N_6163,N_6076,N_6045);
and U6164 (N_6164,N_6099,N_6024);
xnor U6165 (N_6165,N_6055,N_6065);
nor U6166 (N_6166,N_6081,N_6013);
xor U6167 (N_6167,N_6005,N_6097);
or U6168 (N_6168,N_6066,N_6026);
nor U6169 (N_6169,N_6099,N_6043);
or U6170 (N_6170,N_6047,N_6086);
nor U6171 (N_6171,N_6064,N_6099);
or U6172 (N_6172,N_6076,N_6065);
or U6173 (N_6173,N_6083,N_6077);
xor U6174 (N_6174,N_6089,N_6096);
nor U6175 (N_6175,N_6063,N_6058);
nor U6176 (N_6176,N_6065,N_6035);
or U6177 (N_6177,N_6080,N_6072);
nor U6178 (N_6178,N_6034,N_6037);
xnor U6179 (N_6179,N_6098,N_6094);
xor U6180 (N_6180,N_6018,N_6014);
nor U6181 (N_6181,N_6022,N_6078);
nand U6182 (N_6182,N_6065,N_6044);
and U6183 (N_6183,N_6073,N_6029);
or U6184 (N_6184,N_6097,N_6001);
nand U6185 (N_6185,N_6056,N_6009);
or U6186 (N_6186,N_6018,N_6000);
and U6187 (N_6187,N_6066,N_6045);
xor U6188 (N_6188,N_6016,N_6097);
nand U6189 (N_6189,N_6071,N_6063);
and U6190 (N_6190,N_6073,N_6033);
nor U6191 (N_6191,N_6065,N_6067);
xor U6192 (N_6192,N_6072,N_6088);
nor U6193 (N_6193,N_6097,N_6057);
nand U6194 (N_6194,N_6078,N_6044);
or U6195 (N_6195,N_6001,N_6064);
nor U6196 (N_6196,N_6072,N_6056);
nand U6197 (N_6197,N_6042,N_6096);
xor U6198 (N_6198,N_6024,N_6017);
and U6199 (N_6199,N_6037,N_6099);
or U6200 (N_6200,N_6135,N_6131);
nand U6201 (N_6201,N_6118,N_6198);
xnor U6202 (N_6202,N_6144,N_6101);
or U6203 (N_6203,N_6184,N_6127);
nand U6204 (N_6204,N_6141,N_6130);
xnor U6205 (N_6205,N_6134,N_6104);
nand U6206 (N_6206,N_6197,N_6129);
nor U6207 (N_6207,N_6140,N_6167);
or U6208 (N_6208,N_6150,N_6139);
nand U6209 (N_6209,N_6152,N_6149);
nand U6210 (N_6210,N_6146,N_6168);
nand U6211 (N_6211,N_6166,N_6164);
and U6212 (N_6212,N_6154,N_6102);
nand U6213 (N_6213,N_6157,N_6151);
xor U6214 (N_6214,N_6175,N_6195);
nor U6215 (N_6215,N_6136,N_6100);
xor U6216 (N_6216,N_6147,N_6156);
nand U6217 (N_6217,N_6174,N_6191);
xnor U6218 (N_6218,N_6119,N_6143);
xnor U6219 (N_6219,N_6177,N_6117);
and U6220 (N_6220,N_6179,N_6145);
or U6221 (N_6221,N_6112,N_6138);
nor U6222 (N_6222,N_6155,N_6142);
and U6223 (N_6223,N_6109,N_6107);
or U6224 (N_6224,N_6196,N_6132);
nor U6225 (N_6225,N_6176,N_6180);
nand U6226 (N_6226,N_6108,N_6199);
xor U6227 (N_6227,N_6161,N_6181);
or U6228 (N_6228,N_6182,N_6173);
and U6229 (N_6229,N_6162,N_6186);
and U6230 (N_6230,N_6137,N_6171);
or U6231 (N_6231,N_6163,N_6110);
nor U6232 (N_6232,N_6190,N_6106);
or U6233 (N_6233,N_6183,N_6124);
nand U6234 (N_6234,N_6165,N_6148);
nand U6235 (N_6235,N_6188,N_6133);
nor U6236 (N_6236,N_6178,N_6103);
and U6237 (N_6237,N_6192,N_6113);
nand U6238 (N_6238,N_6114,N_6159);
nor U6239 (N_6239,N_6121,N_6111);
xnor U6240 (N_6240,N_6105,N_6189);
nor U6241 (N_6241,N_6123,N_6185);
xnor U6242 (N_6242,N_6125,N_6172);
and U6243 (N_6243,N_6115,N_6170);
and U6244 (N_6244,N_6128,N_6153);
xnor U6245 (N_6245,N_6169,N_6160);
nor U6246 (N_6246,N_6120,N_6122);
nor U6247 (N_6247,N_6126,N_6193);
nand U6248 (N_6248,N_6187,N_6158);
or U6249 (N_6249,N_6116,N_6194);
nor U6250 (N_6250,N_6173,N_6105);
nor U6251 (N_6251,N_6131,N_6199);
and U6252 (N_6252,N_6166,N_6129);
xnor U6253 (N_6253,N_6143,N_6156);
and U6254 (N_6254,N_6132,N_6191);
nand U6255 (N_6255,N_6158,N_6117);
xor U6256 (N_6256,N_6189,N_6181);
xor U6257 (N_6257,N_6107,N_6118);
xor U6258 (N_6258,N_6135,N_6116);
xor U6259 (N_6259,N_6161,N_6178);
or U6260 (N_6260,N_6127,N_6178);
nor U6261 (N_6261,N_6156,N_6144);
nor U6262 (N_6262,N_6158,N_6129);
xor U6263 (N_6263,N_6177,N_6158);
nand U6264 (N_6264,N_6157,N_6189);
nor U6265 (N_6265,N_6193,N_6148);
and U6266 (N_6266,N_6160,N_6119);
xnor U6267 (N_6267,N_6199,N_6175);
nor U6268 (N_6268,N_6122,N_6176);
xor U6269 (N_6269,N_6171,N_6184);
and U6270 (N_6270,N_6182,N_6150);
nor U6271 (N_6271,N_6173,N_6152);
and U6272 (N_6272,N_6113,N_6128);
and U6273 (N_6273,N_6196,N_6194);
xnor U6274 (N_6274,N_6166,N_6193);
xor U6275 (N_6275,N_6191,N_6157);
or U6276 (N_6276,N_6185,N_6170);
or U6277 (N_6277,N_6170,N_6129);
nand U6278 (N_6278,N_6101,N_6116);
and U6279 (N_6279,N_6143,N_6198);
or U6280 (N_6280,N_6143,N_6110);
xnor U6281 (N_6281,N_6176,N_6194);
nor U6282 (N_6282,N_6182,N_6113);
nand U6283 (N_6283,N_6126,N_6131);
xor U6284 (N_6284,N_6133,N_6163);
and U6285 (N_6285,N_6124,N_6165);
and U6286 (N_6286,N_6187,N_6110);
or U6287 (N_6287,N_6137,N_6111);
nor U6288 (N_6288,N_6191,N_6135);
and U6289 (N_6289,N_6191,N_6159);
nor U6290 (N_6290,N_6136,N_6161);
xor U6291 (N_6291,N_6171,N_6189);
nand U6292 (N_6292,N_6115,N_6168);
nor U6293 (N_6293,N_6187,N_6155);
xor U6294 (N_6294,N_6147,N_6199);
xnor U6295 (N_6295,N_6170,N_6195);
nor U6296 (N_6296,N_6147,N_6121);
nor U6297 (N_6297,N_6126,N_6130);
nor U6298 (N_6298,N_6157,N_6124);
nor U6299 (N_6299,N_6133,N_6154);
or U6300 (N_6300,N_6220,N_6232);
and U6301 (N_6301,N_6218,N_6203);
or U6302 (N_6302,N_6274,N_6252);
nand U6303 (N_6303,N_6290,N_6223);
nor U6304 (N_6304,N_6224,N_6201);
xor U6305 (N_6305,N_6281,N_6238);
nor U6306 (N_6306,N_6257,N_6267);
or U6307 (N_6307,N_6222,N_6256);
or U6308 (N_6308,N_6284,N_6233);
xnor U6309 (N_6309,N_6260,N_6227);
or U6310 (N_6310,N_6234,N_6235);
and U6311 (N_6311,N_6264,N_6245);
xor U6312 (N_6312,N_6214,N_6276);
and U6313 (N_6313,N_6221,N_6254);
nand U6314 (N_6314,N_6250,N_6248);
or U6315 (N_6315,N_6273,N_6282);
and U6316 (N_6316,N_6261,N_6263);
nor U6317 (N_6317,N_6292,N_6275);
nor U6318 (N_6318,N_6278,N_6280);
nor U6319 (N_6319,N_6246,N_6225);
and U6320 (N_6320,N_6287,N_6247);
nor U6321 (N_6321,N_6219,N_6206);
or U6322 (N_6322,N_6208,N_6226);
xnor U6323 (N_6323,N_6285,N_6207);
nor U6324 (N_6324,N_6293,N_6251);
and U6325 (N_6325,N_6253,N_6268);
or U6326 (N_6326,N_6271,N_6265);
nor U6327 (N_6327,N_6262,N_6229);
or U6328 (N_6328,N_6241,N_6295);
nor U6329 (N_6329,N_6205,N_6279);
xnor U6330 (N_6330,N_6243,N_6277);
nand U6331 (N_6331,N_6228,N_6289);
and U6332 (N_6332,N_6259,N_6288);
nand U6333 (N_6333,N_6231,N_6249);
xor U6334 (N_6334,N_6272,N_6240);
or U6335 (N_6335,N_6215,N_6202);
or U6336 (N_6336,N_6258,N_6239);
nor U6337 (N_6337,N_6242,N_6294);
nor U6338 (N_6338,N_6283,N_6212);
and U6339 (N_6339,N_6200,N_6204);
and U6340 (N_6340,N_6230,N_6210);
and U6341 (N_6341,N_6291,N_6299);
nor U6342 (N_6342,N_6216,N_6266);
xnor U6343 (N_6343,N_6213,N_6211);
and U6344 (N_6344,N_6244,N_6298);
and U6345 (N_6345,N_6237,N_6255);
xnor U6346 (N_6346,N_6270,N_6209);
nor U6347 (N_6347,N_6217,N_6236);
nor U6348 (N_6348,N_6286,N_6297);
and U6349 (N_6349,N_6296,N_6269);
xnor U6350 (N_6350,N_6215,N_6271);
nand U6351 (N_6351,N_6239,N_6222);
or U6352 (N_6352,N_6261,N_6271);
xor U6353 (N_6353,N_6296,N_6253);
nand U6354 (N_6354,N_6253,N_6227);
or U6355 (N_6355,N_6238,N_6205);
xnor U6356 (N_6356,N_6247,N_6297);
nor U6357 (N_6357,N_6278,N_6298);
or U6358 (N_6358,N_6248,N_6292);
nand U6359 (N_6359,N_6262,N_6227);
or U6360 (N_6360,N_6295,N_6228);
xor U6361 (N_6361,N_6214,N_6217);
xor U6362 (N_6362,N_6208,N_6248);
and U6363 (N_6363,N_6271,N_6259);
nor U6364 (N_6364,N_6203,N_6235);
xor U6365 (N_6365,N_6272,N_6245);
or U6366 (N_6366,N_6221,N_6290);
nand U6367 (N_6367,N_6230,N_6265);
nand U6368 (N_6368,N_6262,N_6207);
nand U6369 (N_6369,N_6288,N_6268);
xor U6370 (N_6370,N_6263,N_6218);
xnor U6371 (N_6371,N_6272,N_6287);
nor U6372 (N_6372,N_6239,N_6253);
xor U6373 (N_6373,N_6289,N_6215);
and U6374 (N_6374,N_6255,N_6265);
and U6375 (N_6375,N_6260,N_6244);
and U6376 (N_6376,N_6284,N_6219);
or U6377 (N_6377,N_6228,N_6258);
xor U6378 (N_6378,N_6261,N_6248);
or U6379 (N_6379,N_6229,N_6202);
nor U6380 (N_6380,N_6289,N_6273);
nor U6381 (N_6381,N_6277,N_6260);
nor U6382 (N_6382,N_6266,N_6233);
nor U6383 (N_6383,N_6295,N_6223);
or U6384 (N_6384,N_6272,N_6200);
and U6385 (N_6385,N_6240,N_6263);
or U6386 (N_6386,N_6203,N_6267);
nor U6387 (N_6387,N_6285,N_6294);
nand U6388 (N_6388,N_6289,N_6252);
or U6389 (N_6389,N_6207,N_6290);
nand U6390 (N_6390,N_6261,N_6250);
nor U6391 (N_6391,N_6286,N_6258);
and U6392 (N_6392,N_6252,N_6264);
xor U6393 (N_6393,N_6201,N_6283);
or U6394 (N_6394,N_6257,N_6245);
xnor U6395 (N_6395,N_6264,N_6230);
and U6396 (N_6396,N_6268,N_6298);
nor U6397 (N_6397,N_6296,N_6220);
or U6398 (N_6398,N_6255,N_6217);
and U6399 (N_6399,N_6206,N_6276);
xnor U6400 (N_6400,N_6324,N_6352);
nor U6401 (N_6401,N_6316,N_6390);
and U6402 (N_6402,N_6383,N_6351);
xnor U6403 (N_6403,N_6360,N_6317);
and U6404 (N_6404,N_6381,N_6378);
xnor U6405 (N_6405,N_6327,N_6362);
and U6406 (N_6406,N_6312,N_6386);
and U6407 (N_6407,N_6338,N_6380);
and U6408 (N_6408,N_6335,N_6398);
and U6409 (N_6409,N_6303,N_6376);
and U6410 (N_6410,N_6379,N_6363);
xnor U6411 (N_6411,N_6354,N_6394);
and U6412 (N_6412,N_6393,N_6375);
nand U6413 (N_6413,N_6388,N_6321);
nor U6414 (N_6414,N_6330,N_6391);
or U6415 (N_6415,N_6346,N_6314);
nand U6416 (N_6416,N_6369,N_6302);
nand U6417 (N_6417,N_6355,N_6311);
nand U6418 (N_6418,N_6364,N_6345);
xnor U6419 (N_6419,N_6342,N_6357);
nor U6420 (N_6420,N_6305,N_6353);
nand U6421 (N_6421,N_6350,N_6361);
nand U6422 (N_6422,N_6358,N_6304);
nand U6423 (N_6423,N_6368,N_6373);
nand U6424 (N_6424,N_6337,N_6318);
or U6425 (N_6425,N_6366,N_6356);
nand U6426 (N_6426,N_6377,N_6310);
nor U6427 (N_6427,N_6372,N_6320);
and U6428 (N_6428,N_6323,N_6392);
nor U6429 (N_6429,N_6306,N_6348);
xor U6430 (N_6430,N_6336,N_6382);
xor U6431 (N_6431,N_6349,N_6344);
xor U6432 (N_6432,N_6384,N_6308);
and U6433 (N_6433,N_6332,N_6339);
nand U6434 (N_6434,N_6397,N_6300);
or U6435 (N_6435,N_6322,N_6359);
nor U6436 (N_6436,N_6367,N_6333);
xor U6437 (N_6437,N_6307,N_6374);
xor U6438 (N_6438,N_6387,N_6309);
nand U6439 (N_6439,N_6395,N_6331);
and U6440 (N_6440,N_6370,N_6319);
nor U6441 (N_6441,N_6399,N_6340);
or U6442 (N_6442,N_6389,N_6396);
and U6443 (N_6443,N_6328,N_6347);
and U6444 (N_6444,N_6315,N_6313);
and U6445 (N_6445,N_6385,N_6341);
or U6446 (N_6446,N_6365,N_6325);
and U6447 (N_6447,N_6326,N_6334);
and U6448 (N_6448,N_6371,N_6301);
nor U6449 (N_6449,N_6343,N_6329);
nand U6450 (N_6450,N_6350,N_6329);
nor U6451 (N_6451,N_6363,N_6344);
or U6452 (N_6452,N_6364,N_6308);
or U6453 (N_6453,N_6352,N_6307);
nor U6454 (N_6454,N_6367,N_6372);
or U6455 (N_6455,N_6375,N_6321);
nand U6456 (N_6456,N_6303,N_6391);
nor U6457 (N_6457,N_6351,N_6359);
xnor U6458 (N_6458,N_6338,N_6361);
and U6459 (N_6459,N_6336,N_6325);
nor U6460 (N_6460,N_6311,N_6343);
nor U6461 (N_6461,N_6368,N_6381);
nand U6462 (N_6462,N_6391,N_6398);
and U6463 (N_6463,N_6350,N_6322);
and U6464 (N_6464,N_6377,N_6337);
nand U6465 (N_6465,N_6302,N_6392);
nor U6466 (N_6466,N_6305,N_6351);
or U6467 (N_6467,N_6356,N_6395);
or U6468 (N_6468,N_6390,N_6383);
xor U6469 (N_6469,N_6370,N_6318);
and U6470 (N_6470,N_6343,N_6351);
or U6471 (N_6471,N_6388,N_6326);
and U6472 (N_6472,N_6390,N_6347);
or U6473 (N_6473,N_6315,N_6350);
nand U6474 (N_6474,N_6303,N_6379);
and U6475 (N_6475,N_6368,N_6362);
nor U6476 (N_6476,N_6362,N_6345);
or U6477 (N_6477,N_6343,N_6371);
nor U6478 (N_6478,N_6320,N_6392);
nor U6479 (N_6479,N_6388,N_6322);
and U6480 (N_6480,N_6391,N_6358);
nor U6481 (N_6481,N_6378,N_6380);
xnor U6482 (N_6482,N_6351,N_6397);
or U6483 (N_6483,N_6300,N_6323);
and U6484 (N_6484,N_6349,N_6328);
nand U6485 (N_6485,N_6378,N_6379);
or U6486 (N_6486,N_6348,N_6385);
nand U6487 (N_6487,N_6366,N_6305);
or U6488 (N_6488,N_6313,N_6378);
nand U6489 (N_6489,N_6393,N_6326);
and U6490 (N_6490,N_6349,N_6335);
nand U6491 (N_6491,N_6340,N_6359);
nor U6492 (N_6492,N_6310,N_6303);
xnor U6493 (N_6493,N_6367,N_6363);
or U6494 (N_6494,N_6355,N_6384);
and U6495 (N_6495,N_6351,N_6362);
or U6496 (N_6496,N_6385,N_6349);
xnor U6497 (N_6497,N_6312,N_6389);
and U6498 (N_6498,N_6333,N_6341);
or U6499 (N_6499,N_6343,N_6336);
xor U6500 (N_6500,N_6488,N_6427);
nor U6501 (N_6501,N_6449,N_6483);
and U6502 (N_6502,N_6439,N_6413);
nor U6503 (N_6503,N_6489,N_6431);
and U6504 (N_6504,N_6480,N_6410);
and U6505 (N_6505,N_6428,N_6475);
nand U6506 (N_6506,N_6482,N_6448);
or U6507 (N_6507,N_6442,N_6409);
nor U6508 (N_6508,N_6469,N_6497);
nand U6509 (N_6509,N_6496,N_6425);
xnor U6510 (N_6510,N_6408,N_6451);
nor U6511 (N_6511,N_6464,N_6402);
xor U6512 (N_6512,N_6471,N_6433);
xnor U6513 (N_6513,N_6485,N_6404);
or U6514 (N_6514,N_6456,N_6461);
or U6515 (N_6515,N_6453,N_6498);
and U6516 (N_6516,N_6452,N_6484);
nand U6517 (N_6517,N_6499,N_6486);
xor U6518 (N_6518,N_6458,N_6420);
or U6519 (N_6519,N_6440,N_6481);
nor U6520 (N_6520,N_6478,N_6403);
and U6521 (N_6521,N_6407,N_6443);
or U6522 (N_6522,N_6424,N_6444);
nand U6523 (N_6523,N_6419,N_6470);
or U6524 (N_6524,N_6491,N_6487);
and U6525 (N_6525,N_6473,N_6492);
or U6526 (N_6526,N_6437,N_6455);
xor U6527 (N_6527,N_6457,N_6454);
and U6528 (N_6528,N_6468,N_6426);
xor U6529 (N_6529,N_6417,N_6436);
nand U6530 (N_6530,N_6472,N_6412);
nand U6531 (N_6531,N_6435,N_6421);
and U6532 (N_6532,N_6465,N_6445);
nand U6533 (N_6533,N_6474,N_6414);
nand U6534 (N_6534,N_6418,N_6406);
or U6535 (N_6535,N_6438,N_6466);
xor U6536 (N_6536,N_6459,N_6447);
nand U6537 (N_6537,N_6416,N_6415);
and U6538 (N_6538,N_6450,N_6463);
nor U6539 (N_6539,N_6446,N_6400);
xor U6540 (N_6540,N_6495,N_6467);
or U6541 (N_6541,N_6479,N_6423);
nor U6542 (N_6542,N_6422,N_6434);
nor U6543 (N_6543,N_6432,N_6429);
or U6544 (N_6544,N_6401,N_6405);
or U6545 (N_6545,N_6411,N_6477);
and U6546 (N_6546,N_6493,N_6460);
xor U6547 (N_6547,N_6476,N_6441);
and U6548 (N_6548,N_6430,N_6490);
xnor U6549 (N_6549,N_6494,N_6462);
or U6550 (N_6550,N_6434,N_6476);
xor U6551 (N_6551,N_6446,N_6450);
and U6552 (N_6552,N_6481,N_6470);
and U6553 (N_6553,N_6440,N_6419);
and U6554 (N_6554,N_6404,N_6425);
or U6555 (N_6555,N_6499,N_6420);
xor U6556 (N_6556,N_6484,N_6438);
nand U6557 (N_6557,N_6402,N_6495);
xor U6558 (N_6558,N_6470,N_6451);
nand U6559 (N_6559,N_6478,N_6483);
nand U6560 (N_6560,N_6469,N_6472);
xnor U6561 (N_6561,N_6444,N_6491);
nor U6562 (N_6562,N_6444,N_6488);
nor U6563 (N_6563,N_6474,N_6455);
and U6564 (N_6564,N_6425,N_6417);
xor U6565 (N_6565,N_6449,N_6495);
nor U6566 (N_6566,N_6402,N_6451);
or U6567 (N_6567,N_6424,N_6492);
nand U6568 (N_6568,N_6403,N_6458);
and U6569 (N_6569,N_6468,N_6475);
nand U6570 (N_6570,N_6483,N_6437);
xnor U6571 (N_6571,N_6430,N_6459);
or U6572 (N_6572,N_6421,N_6487);
nand U6573 (N_6573,N_6444,N_6472);
xnor U6574 (N_6574,N_6423,N_6403);
and U6575 (N_6575,N_6490,N_6441);
nand U6576 (N_6576,N_6481,N_6486);
and U6577 (N_6577,N_6446,N_6456);
and U6578 (N_6578,N_6409,N_6411);
and U6579 (N_6579,N_6402,N_6483);
nand U6580 (N_6580,N_6405,N_6410);
nor U6581 (N_6581,N_6491,N_6407);
nand U6582 (N_6582,N_6480,N_6470);
and U6583 (N_6583,N_6439,N_6473);
xor U6584 (N_6584,N_6425,N_6498);
and U6585 (N_6585,N_6441,N_6496);
nand U6586 (N_6586,N_6476,N_6431);
or U6587 (N_6587,N_6441,N_6462);
and U6588 (N_6588,N_6455,N_6457);
or U6589 (N_6589,N_6423,N_6457);
and U6590 (N_6590,N_6435,N_6473);
nor U6591 (N_6591,N_6446,N_6402);
nand U6592 (N_6592,N_6410,N_6400);
nor U6593 (N_6593,N_6447,N_6448);
or U6594 (N_6594,N_6433,N_6454);
nand U6595 (N_6595,N_6435,N_6459);
nor U6596 (N_6596,N_6402,N_6425);
xor U6597 (N_6597,N_6457,N_6412);
nand U6598 (N_6598,N_6494,N_6425);
nor U6599 (N_6599,N_6428,N_6471);
xnor U6600 (N_6600,N_6507,N_6552);
or U6601 (N_6601,N_6574,N_6516);
and U6602 (N_6602,N_6522,N_6526);
nor U6603 (N_6603,N_6504,N_6580);
nand U6604 (N_6604,N_6539,N_6554);
xor U6605 (N_6605,N_6509,N_6532);
or U6606 (N_6606,N_6584,N_6521);
xor U6607 (N_6607,N_6589,N_6594);
nand U6608 (N_6608,N_6536,N_6579);
and U6609 (N_6609,N_6520,N_6556);
nor U6610 (N_6610,N_6555,N_6548);
or U6611 (N_6611,N_6567,N_6577);
nor U6612 (N_6612,N_6588,N_6550);
xnor U6613 (N_6613,N_6544,N_6585);
xor U6614 (N_6614,N_6518,N_6595);
or U6615 (N_6615,N_6529,N_6575);
or U6616 (N_6616,N_6559,N_6511);
nand U6617 (N_6617,N_6578,N_6524);
xor U6618 (N_6618,N_6563,N_6596);
xnor U6619 (N_6619,N_6591,N_6525);
xnor U6620 (N_6620,N_6569,N_6535);
or U6621 (N_6621,N_6592,N_6506);
or U6622 (N_6622,N_6531,N_6515);
nor U6623 (N_6623,N_6564,N_6553);
xnor U6624 (N_6624,N_6543,N_6505);
nor U6625 (N_6625,N_6549,N_6570);
or U6626 (N_6626,N_6571,N_6513);
or U6627 (N_6627,N_6514,N_6587);
nor U6628 (N_6628,N_6537,N_6546);
xor U6629 (N_6629,N_6542,N_6573);
nor U6630 (N_6630,N_6583,N_6508);
nor U6631 (N_6631,N_6545,N_6510);
and U6632 (N_6632,N_6547,N_6551);
or U6633 (N_6633,N_6565,N_6566);
nand U6634 (N_6634,N_6572,N_6530);
xnor U6635 (N_6635,N_6560,N_6541);
or U6636 (N_6636,N_6599,N_6586);
xor U6637 (N_6637,N_6598,N_6568);
and U6638 (N_6638,N_6527,N_6503);
and U6639 (N_6639,N_6590,N_6519);
nand U6640 (N_6640,N_6597,N_6561);
xnor U6641 (N_6641,N_6517,N_6533);
nor U6642 (N_6642,N_6581,N_6501);
or U6643 (N_6643,N_6540,N_6500);
xnor U6644 (N_6644,N_6528,N_6557);
nand U6645 (N_6645,N_6502,N_6538);
nand U6646 (N_6646,N_6582,N_6576);
and U6647 (N_6647,N_6558,N_6534);
nand U6648 (N_6648,N_6512,N_6593);
nand U6649 (N_6649,N_6523,N_6562);
or U6650 (N_6650,N_6524,N_6545);
or U6651 (N_6651,N_6559,N_6542);
and U6652 (N_6652,N_6541,N_6551);
nor U6653 (N_6653,N_6584,N_6586);
or U6654 (N_6654,N_6566,N_6563);
and U6655 (N_6655,N_6555,N_6553);
nor U6656 (N_6656,N_6533,N_6551);
xor U6657 (N_6657,N_6551,N_6584);
and U6658 (N_6658,N_6504,N_6567);
or U6659 (N_6659,N_6554,N_6569);
and U6660 (N_6660,N_6545,N_6550);
or U6661 (N_6661,N_6544,N_6574);
and U6662 (N_6662,N_6579,N_6507);
xor U6663 (N_6663,N_6593,N_6598);
nand U6664 (N_6664,N_6568,N_6586);
nor U6665 (N_6665,N_6585,N_6567);
xor U6666 (N_6666,N_6551,N_6512);
or U6667 (N_6667,N_6545,N_6551);
nor U6668 (N_6668,N_6534,N_6596);
and U6669 (N_6669,N_6565,N_6504);
nand U6670 (N_6670,N_6500,N_6515);
and U6671 (N_6671,N_6509,N_6527);
nand U6672 (N_6672,N_6529,N_6516);
xor U6673 (N_6673,N_6532,N_6522);
xor U6674 (N_6674,N_6570,N_6551);
nor U6675 (N_6675,N_6564,N_6590);
nor U6676 (N_6676,N_6546,N_6560);
xor U6677 (N_6677,N_6533,N_6546);
or U6678 (N_6678,N_6527,N_6541);
nand U6679 (N_6679,N_6543,N_6562);
and U6680 (N_6680,N_6526,N_6505);
and U6681 (N_6681,N_6510,N_6570);
nand U6682 (N_6682,N_6535,N_6590);
and U6683 (N_6683,N_6513,N_6556);
nor U6684 (N_6684,N_6557,N_6559);
and U6685 (N_6685,N_6537,N_6555);
nand U6686 (N_6686,N_6513,N_6576);
and U6687 (N_6687,N_6513,N_6548);
nand U6688 (N_6688,N_6569,N_6523);
xnor U6689 (N_6689,N_6556,N_6533);
nand U6690 (N_6690,N_6565,N_6540);
xnor U6691 (N_6691,N_6546,N_6597);
nand U6692 (N_6692,N_6534,N_6566);
nor U6693 (N_6693,N_6559,N_6551);
nor U6694 (N_6694,N_6548,N_6536);
nor U6695 (N_6695,N_6556,N_6559);
or U6696 (N_6696,N_6515,N_6511);
and U6697 (N_6697,N_6574,N_6528);
nor U6698 (N_6698,N_6570,N_6548);
and U6699 (N_6699,N_6526,N_6520);
or U6700 (N_6700,N_6649,N_6659);
and U6701 (N_6701,N_6679,N_6678);
nand U6702 (N_6702,N_6640,N_6631);
xor U6703 (N_6703,N_6615,N_6664);
nand U6704 (N_6704,N_6637,N_6619);
and U6705 (N_6705,N_6639,N_6625);
and U6706 (N_6706,N_6653,N_6606);
nor U6707 (N_6707,N_6668,N_6692);
or U6708 (N_6708,N_6618,N_6630);
or U6709 (N_6709,N_6609,N_6646);
nand U6710 (N_6710,N_6641,N_6654);
or U6711 (N_6711,N_6636,N_6663);
nor U6712 (N_6712,N_6658,N_6614);
nor U6713 (N_6713,N_6695,N_6674);
or U6714 (N_6714,N_6699,N_6608);
nor U6715 (N_6715,N_6655,N_6642);
xnor U6716 (N_6716,N_6666,N_6656);
xnor U6717 (N_6717,N_6647,N_6671);
nand U6718 (N_6718,N_6660,N_6613);
nor U6719 (N_6719,N_6673,N_6675);
or U6720 (N_6720,N_6650,N_6643);
nor U6721 (N_6721,N_6682,N_6605);
or U6722 (N_6722,N_6690,N_6627);
and U6723 (N_6723,N_6634,N_6698);
xor U6724 (N_6724,N_6681,N_6648);
nor U6725 (N_6725,N_6693,N_6623);
nor U6726 (N_6726,N_6622,N_6661);
or U6727 (N_6727,N_6662,N_6620);
xor U6728 (N_6728,N_6617,N_6638);
nor U6729 (N_6729,N_6633,N_6632);
xor U6730 (N_6730,N_6657,N_6628);
or U6731 (N_6731,N_6645,N_6624);
and U6732 (N_6732,N_6689,N_6626);
xor U6733 (N_6733,N_6685,N_6684);
nor U6734 (N_6734,N_6691,N_6697);
nand U6735 (N_6735,N_6686,N_6612);
or U6736 (N_6736,N_6651,N_6644);
or U6737 (N_6737,N_6683,N_6669);
and U6738 (N_6738,N_6621,N_6600);
or U6739 (N_6739,N_6604,N_6602);
xor U6740 (N_6740,N_6629,N_6687);
or U6741 (N_6741,N_6667,N_6616);
nand U6742 (N_6742,N_6601,N_6635);
xor U6743 (N_6743,N_6611,N_6694);
nand U6744 (N_6744,N_6610,N_6665);
nor U6745 (N_6745,N_6670,N_6672);
or U6746 (N_6746,N_6677,N_6603);
nand U6747 (N_6747,N_6652,N_6676);
nand U6748 (N_6748,N_6680,N_6688);
xor U6749 (N_6749,N_6607,N_6696);
xor U6750 (N_6750,N_6678,N_6660);
nor U6751 (N_6751,N_6608,N_6607);
xor U6752 (N_6752,N_6654,N_6678);
and U6753 (N_6753,N_6692,N_6644);
xor U6754 (N_6754,N_6620,N_6648);
xnor U6755 (N_6755,N_6642,N_6650);
or U6756 (N_6756,N_6606,N_6648);
xor U6757 (N_6757,N_6661,N_6692);
nand U6758 (N_6758,N_6608,N_6657);
xnor U6759 (N_6759,N_6678,N_6630);
nor U6760 (N_6760,N_6610,N_6675);
nor U6761 (N_6761,N_6659,N_6695);
nand U6762 (N_6762,N_6647,N_6649);
nand U6763 (N_6763,N_6618,N_6696);
xor U6764 (N_6764,N_6606,N_6654);
nand U6765 (N_6765,N_6666,N_6628);
nand U6766 (N_6766,N_6661,N_6653);
xnor U6767 (N_6767,N_6655,N_6622);
xnor U6768 (N_6768,N_6607,N_6660);
nor U6769 (N_6769,N_6657,N_6661);
or U6770 (N_6770,N_6695,N_6618);
or U6771 (N_6771,N_6656,N_6695);
or U6772 (N_6772,N_6617,N_6609);
nor U6773 (N_6773,N_6670,N_6651);
and U6774 (N_6774,N_6632,N_6685);
or U6775 (N_6775,N_6667,N_6698);
and U6776 (N_6776,N_6691,N_6604);
or U6777 (N_6777,N_6612,N_6692);
xnor U6778 (N_6778,N_6690,N_6631);
and U6779 (N_6779,N_6600,N_6612);
and U6780 (N_6780,N_6662,N_6656);
or U6781 (N_6781,N_6687,N_6650);
xor U6782 (N_6782,N_6668,N_6603);
xnor U6783 (N_6783,N_6604,N_6660);
nor U6784 (N_6784,N_6673,N_6642);
nand U6785 (N_6785,N_6666,N_6616);
or U6786 (N_6786,N_6608,N_6698);
nor U6787 (N_6787,N_6646,N_6604);
and U6788 (N_6788,N_6629,N_6674);
xnor U6789 (N_6789,N_6698,N_6694);
or U6790 (N_6790,N_6631,N_6605);
nand U6791 (N_6791,N_6679,N_6620);
nor U6792 (N_6792,N_6687,N_6609);
and U6793 (N_6793,N_6632,N_6638);
xor U6794 (N_6794,N_6685,N_6672);
nand U6795 (N_6795,N_6638,N_6670);
and U6796 (N_6796,N_6653,N_6691);
nand U6797 (N_6797,N_6604,N_6611);
xnor U6798 (N_6798,N_6649,N_6601);
nor U6799 (N_6799,N_6612,N_6640);
or U6800 (N_6800,N_6758,N_6725);
nand U6801 (N_6801,N_6770,N_6736);
nand U6802 (N_6802,N_6795,N_6718);
nor U6803 (N_6803,N_6757,N_6777);
nand U6804 (N_6804,N_6721,N_6752);
nand U6805 (N_6805,N_6793,N_6734);
nand U6806 (N_6806,N_6747,N_6765);
nor U6807 (N_6807,N_6705,N_6733);
xnor U6808 (N_6808,N_6751,N_6701);
nand U6809 (N_6809,N_6763,N_6719);
nand U6810 (N_6810,N_6781,N_6788);
nor U6811 (N_6811,N_6766,N_6710);
nand U6812 (N_6812,N_6776,N_6741);
or U6813 (N_6813,N_6742,N_6700);
or U6814 (N_6814,N_6755,N_6798);
nor U6815 (N_6815,N_6782,N_6759);
xor U6816 (N_6816,N_6756,N_6762);
xor U6817 (N_6817,N_6787,N_6711);
and U6818 (N_6818,N_6717,N_6707);
nor U6819 (N_6819,N_6729,N_6774);
and U6820 (N_6820,N_6789,N_6792);
nor U6821 (N_6821,N_6761,N_6713);
xnor U6822 (N_6822,N_6764,N_6775);
and U6823 (N_6823,N_6784,N_6780);
nand U6824 (N_6824,N_6732,N_6738);
nor U6825 (N_6825,N_6767,N_6743);
and U6826 (N_6826,N_6712,N_6708);
or U6827 (N_6827,N_6728,N_6786);
xnor U6828 (N_6828,N_6706,N_6797);
nand U6829 (N_6829,N_6702,N_6704);
nor U6830 (N_6830,N_6771,N_6796);
and U6831 (N_6831,N_6748,N_6754);
xnor U6832 (N_6832,N_6731,N_6722);
nand U6833 (N_6833,N_6714,N_6720);
nor U6834 (N_6834,N_6783,N_6772);
or U6835 (N_6835,N_6749,N_6744);
and U6836 (N_6836,N_6737,N_6799);
xnor U6837 (N_6837,N_6769,N_6723);
or U6838 (N_6838,N_6791,N_6735);
or U6839 (N_6839,N_6790,N_6726);
nor U6840 (N_6840,N_6727,N_6753);
xnor U6841 (N_6841,N_6715,N_6778);
and U6842 (N_6842,N_6709,N_6750);
nor U6843 (N_6843,N_6768,N_6779);
or U6844 (N_6844,N_6746,N_6716);
or U6845 (N_6845,N_6745,N_6739);
xnor U6846 (N_6846,N_6760,N_6740);
nand U6847 (N_6847,N_6703,N_6773);
xnor U6848 (N_6848,N_6785,N_6794);
xor U6849 (N_6849,N_6730,N_6724);
nand U6850 (N_6850,N_6737,N_6758);
nand U6851 (N_6851,N_6758,N_6779);
nand U6852 (N_6852,N_6764,N_6799);
nand U6853 (N_6853,N_6766,N_6700);
or U6854 (N_6854,N_6773,N_6732);
and U6855 (N_6855,N_6796,N_6731);
xnor U6856 (N_6856,N_6710,N_6740);
nor U6857 (N_6857,N_6712,N_6703);
nor U6858 (N_6858,N_6751,N_6700);
nor U6859 (N_6859,N_6778,N_6799);
nor U6860 (N_6860,N_6792,N_6771);
nand U6861 (N_6861,N_6762,N_6722);
xnor U6862 (N_6862,N_6784,N_6779);
xnor U6863 (N_6863,N_6728,N_6741);
nor U6864 (N_6864,N_6778,N_6703);
nand U6865 (N_6865,N_6770,N_6704);
xnor U6866 (N_6866,N_6718,N_6724);
and U6867 (N_6867,N_6771,N_6798);
nor U6868 (N_6868,N_6781,N_6769);
and U6869 (N_6869,N_6760,N_6729);
or U6870 (N_6870,N_6768,N_6726);
and U6871 (N_6871,N_6771,N_6732);
nor U6872 (N_6872,N_6782,N_6733);
nand U6873 (N_6873,N_6741,N_6700);
xnor U6874 (N_6874,N_6742,N_6793);
and U6875 (N_6875,N_6760,N_6724);
nand U6876 (N_6876,N_6716,N_6781);
nor U6877 (N_6877,N_6779,N_6763);
or U6878 (N_6878,N_6766,N_6748);
nand U6879 (N_6879,N_6762,N_6778);
and U6880 (N_6880,N_6787,N_6753);
nor U6881 (N_6881,N_6770,N_6746);
and U6882 (N_6882,N_6719,N_6735);
and U6883 (N_6883,N_6787,N_6707);
nand U6884 (N_6884,N_6790,N_6704);
xnor U6885 (N_6885,N_6732,N_6788);
xnor U6886 (N_6886,N_6757,N_6722);
xnor U6887 (N_6887,N_6795,N_6702);
xnor U6888 (N_6888,N_6708,N_6794);
xnor U6889 (N_6889,N_6728,N_6748);
or U6890 (N_6890,N_6737,N_6796);
xor U6891 (N_6891,N_6757,N_6710);
nor U6892 (N_6892,N_6765,N_6793);
or U6893 (N_6893,N_6763,N_6726);
xor U6894 (N_6894,N_6776,N_6703);
nand U6895 (N_6895,N_6773,N_6738);
or U6896 (N_6896,N_6734,N_6762);
xnor U6897 (N_6897,N_6741,N_6726);
nand U6898 (N_6898,N_6744,N_6757);
xor U6899 (N_6899,N_6797,N_6735);
nand U6900 (N_6900,N_6801,N_6871);
nor U6901 (N_6901,N_6849,N_6853);
nor U6902 (N_6902,N_6803,N_6800);
nor U6903 (N_6903,N_6838,N_6822);
and U6904 (N_6904,N_6844,N_6887);
nor U6905 (N_6905,N_6892,N_6863);
or U6906 (N_6906,N_6835,N_6855);
xnor U6907 (N_6907,N_6873,N_6852);
nand U6908 (N_6908,N_6826,N_6809);
xor U6909 (N_6909,N_6832,N_6859);
or U6910 (N_6910,N_6879,N_6827);
and U6911 (N_6911,N_6829,N_6866);
and U6912 (N_6912,N_6804,N_6897);
and U6913 (N_6913,N_6865,N_6895);
nand U6914 (N_6914,N_6840,N_6875);
or U6915 (N_6915,N_6815,N_6812);
and U6916 (N_6916,N_6872,N_6867);
or U6917 (N_6917,N_6882,N_6884);
or U6918 (N_6918,N_6810,N_6837);
and U6919 (N_6919,N_6823,N_6828);
and U6920 (N_6920,N_6845,N_6802);
nor U6921 (N_6921,N_6807,N_6896);
xnor U6922 (N_6922,N_6850,N_6841);
and U6923 (N_6923,N_6808,N_6898);
and U6924 (N_6924,N_6858,N_6877);
xnor U6925 (N_6925,N_6883,N_6819);
xor U6926 (N_6926,N_6864,N_6861);
nand U6927 (N_6927,N_6833,N_6857);
and U6928 (N_6928,N_6820,N_6894);
nand U6929 (N_6929,N_6856,N_6824);
or U6930 (N_6930,N_6848,N_6881);
nor U6931 (N_6931,N_6805,N_6830);
and U6932 (N_6932,N_6889,N_6825);
nor U6933 (N_6933,N_6869,N_6868);
and U6934 (N_6934,N_6811,N_6821);
nand U6935 (N_6935,N_6870,N_6817);
xnor U6936 (N_6936,N_6885,N_6831);
xnor U6937 (N_6937,N_6891,N_6876);
or U6938 (N_6938,N_6836,N_6893);
nand U6939 (N_6939,N_6851,N_6806);
nand U6940 (N_6940,N_6854,N_6846);
or U6941 (N_6941,N_6862,N_6880);
or U6942 (N_6942,N_6834,N_6839);
nor U6943 (N_6943,N_6878,N_6888);
xnor U6944 (N_6944,N_6813,N_6886);
nor U6945 (N_6945,N_6899,N_6814);
nor U6946 (N_6946,N_6842,N_6818);
nor U6947 (N_6947,N_6890,N_6860);
and U6948 (N_6948,N_6843,N_6847);
and U6949 (N_6949,N_6816,N_6874);
xor U6950 (N_6950,N_6873,N_6859);
and U6951 (N_6951,N_6858,N_6859);
nor U6952 (N_6952,N_6819,N_6827);
xor U6953 (N_6953,N_6893,N_6820);
and U6954 (N_6954,N_6812,N_6867);
nand U6955 (N_6955,N_6849,N_6855);
nand U6956 (N_6956,N_6846,N_6899);
or U6957 (N_6957,N_6879,N_6855);
nand U6958 (N_6958,N_6885,N_6833);
xnor U6959 (N_6959,N_6831,N_6892);
and U6960 (N_6960,N_6828,N_6899);
xnor U6961 (N_6961,N_6872,N_6864);
xnor U6962 (N_6962,N_6855,N_6802);
nand U6963 (N_6963,N_6889,N_6806);
nand U6964 (N_6964,N_6855,N_6831);
xnor U6965 (N_6965,N_6882,N_6853);
xnor U6966 (N_6966,N_6881,N_6806);
or U6967 (N_6967,N_6841,N_6800);
and U6968 (N_6968,N_6826,N_6856);
nor U6969 (N_6969,N_6825,N_6820);
nand U6970 (N_6970,N_6866,N_6894);
or U6971 (N_6971,N_6883,N_6895);
xor U6972 (N_6972,N_6865,N_6816);
nor U6973 (N_6973,N_6812,N_6831);
nor U6974 (N_6974,N_6880,N_6842);
xor U6975 (N_6975,N_6819,N_6896);
nand U6976 (N_6976,N_6830,N_6850);
xor U6977 (N_6977,N_6878,N_6893);
nand U6978 (N_6978,N_6848,N_6892);
xnor U6979 (N_6979,N_6863,N_6880);
nor U6980 (N_6980,N_6804,N_6853);
xnor U6981 (N_6981,N_6872,N_6823);
nand U6982 (N_6982,N_6890,N_6807);
nand U6983 (N_6983,N_6886,N_6811);
xnor U6984 (N_6984,N_6875,N_6868);
xor U6985 (N_6985,N_6827,N_6892);
or U6986 (N_6986,N_6841,N_6832);
and U6987 (N_6987,N_6870,N_6809);
xnor U6988 (N_6988,N_6825,N_6875);
xnor U6989 (N_6989,N_6810,N_6829);
and U6990 (N_6990,N_6882,N_6848);
nand U6991 (N_6991,N_6806,N_6855);
xnor U6992 (N_6992,N_6801,N_6887);
and U6993 (N_6993,N_6806,N_6812);
or U6994 (N_6994,N_6821,N_6802);
nor U6995 (N_6995,N_6855,N_6854);
nor U6996 (N_6996,N_6830,N_6854);
nand U6997 (N_6997,N_6866,N_6869);
and U6998 (N_6998,N_6860,N_6872);
xor U6999 (N_6999,N_6823,N_6841);
xnor U7000 (N_7000,N_6909,N_6936);
or U7001 (N_7001,N_6961,N_6989);
and U7002 (N_7002,N_6971,N_6946);
nand U7003 (N_7003,N_6978,N_6900);
or U7004 (N_7004,N_6905,N_6917);
nand U7005 (N_7005,N_6982,N_6951);
nand U7006 (N_7006,N_6907,N_6981);
xnor U7007 (N_7007,N_6970,N_6906);
xor U7008 (N_7008,N_6930,N_6975);
xor U7009 (N_7009,N_6990,N_6974);
nor U7010 (N_7010,N_6944,N_6995);
xnor U7011 (N_7011,N_6920,N_6940);
and U7012 (N_7012,N_6926,N_6957);
or U7013 (N_7013,N_6999,N_6992);
or U7014 (N_7014,N_6949,N_6924);
xnor U7015 (N_7015,N_6985,N_6954);
nor U7016 (N_7016,N_6903,N_6908);
nor U7017 (N_7017,N_6913,N_6925);
or U7018 (N_7018,N_6972,N_6953);
nand U7019 (N_7019,N_6929,N_6963);
or U7020 (N_7020,N_6967,N_6956);
or U7021 (N_7021,N_6923,N_6916);
or U7022 (N_7022,N_6996,N_6934);
nand U7023 (N_7023,N_6904,N_6968);
xnor U7024 (N_7024,N_6922,N_6901);
or U7025 (N_7025,N_6939,N_6935);
xor U7026 (N_7026,N_6948,N_6994);
nor U7027 (N_7027,N_6931,N_6959);
xor U7028 (N_7028,N_6943,N_6911);
xnor U7029 (N_7029,N_6933,N_6984);
and U7030 (N_7030,N_6973,N_6962);
nand U7031 (N_7031,N_6942,N_6993);
nor U7032 (N_7032,N_6919,N_6902);
and U7033 (N_7033,N_6945,N_6979);
nor U7034 (N_7034,N_6938,N_6988);
or U7035 (N_7035,N_6997,N_6937);
nand U7036 (N_7036,N_6912,N_6915);
nor U7037 (N_7037,N_6958,N_6977);
and U7038 (N_7038,N_6960,N_6976);
or U7039 (N_7039,N_6987,N_6986);
and U7040 (N_7040,N_6952,N_6965);
xnor U7041 (N_7041,N_6980,N_6927);
and U7042 (N_7042,N_6998,N_6991);
or U7043 (N_7043,N_6918,N_6955);
nand U7044 (N_7044,N_6914,N_6947);
nand U7045 (N_7045,N_6950,N_6966);
xnor U7046 (N_7046,N_6941,N_6921);
nand U7047 (N_7047,N_6969,N_6983);
or U7048 (N_7048,N_6964,N_6928);
and U7049 (N_7049,N_6932,N_6910);
and U7050 (N_7050,N_6917,N_6956);
nor U7051 (N_7051,N_6935,N_6913);
and U7052 (N_7052,N_6987,N_6965);
nor U7053 (N_7053,N_6951,N_6965);
or U7054 (N_7054,N_6992,N_6977);
or U7055 (N_7055,N_6959,N_6995);
nand U7056 (N_7056,N_6909,N_6929);
or U7057 (N_7057,N_6964,N_6900);
nor U7058 (N_7058,N_6934,N_6949);
xor U7059 (N_7059,N_6963,N_6935);
or U7060 (N_7060,N_6918,N_6937);
and U7061 (N_7061,N_6908,N_6934);
nor U7062 (N_7062,N_6968,N_6927);
or U7063 (N_7063,N_6971,N_6921);
and U7064 (N_7064,N_6912,N_6908);
nor U7065 (N_7065,N_6945,N_6955);
and U7066 (N_7066,N_6917,N_6923);
nand U7067 (N_7067,N_6955,N_6995);
and U7068 (N_7068,N_6917,N_6927);
or U7069 (N_7069,N_6997,N_6901);
xor U7070 (N_7070,N_6979,N_6941);
nor U7071 (N_7071,N_6913,N_6927);
and U7072 (N_7072,N_6914,N_6956);
nor U7073 (N_7073,N_6948,N_6951);
xnor U7074 (N_7074,N_6950,N_6919);
xnor U7075 (N_7075,N_6996,N_6969);
and U7076 (N_7076,N_6975,N_6999);
or U7077 (N_7077,N_6992,N_6958);
nand U7078 (N_7078,N_6981,N_6968);
nand U7079 (N_7079,N_6933,N_6987);
nand U7080 (N_7080,N_6974,N_6951);
xnor U7081 (N_7081,N_6947,N_6901);
nor U7082 (N_7082,N_6961,N_6993);
nand U7083 (N_7083,N_6985,N_6948);
nor U7084 (N_7084,N_6914,N_6944);
nand U7085 (N_7085,N_6900,N_6912);
xnor U7086 (N_7086,N_6993,N_6925);
and U7087 (N_7087,N_6949,N_6972);
xnor U7088 (N_7088,N_6953,N_6928);
and U7089 (N_7089,N_6902,N_6998);
nand U7090 (N_7090,N_6994,N_6989);
nand U7091 (N_7091,N_6940,N_6921);
nor U7092 (N_7092,N_6978,N_6985);
nand U7093 (N_7093,N_6950,N_6995);
nor U7094 (N_7094,N_6961,N_6933);
and U7095 (N_7095,N_6925,N_6962);
or U7096 (N_7096,N_6965,N_6949);
nand U7097 (N_7097,N_6902,N_6952);
nand U7098 (N_7098,N_6972,N_6964);
nor U7099 (N_7099,N_6991,N_6914);
xor U7100 (N_7100,N_7058,N_7043);
and U7101 (N_7101,N_7066,N_7007);
nor U7102 (N_7102,N_7042,N_7060);
xnor U7103 (N_7103,N_7009,N_7073);
nor U7104 (N_7104,N_7098,N_7019);
and U7105 (N_7105,N_7056,N_7036);
nor U7106 (N_7106,N_7051,N_7024);
xor U7107 (N_7107,N_7085,N_7059);
nor U7108 (N_7108,N_7029,N_7040);
nor U7109 (N_7109,N_7050,N_7054);
or U7110 (N_7110,N_7084,N_7083);
or U7111 (N_7111,N_7017,N_7065);
nand U7112 (N_7112,N_7074,N_7090);
xnor U7113 (N_7113,N_7021,N_7047);
and U7114 (N_7114,N_7082,N_7016);
xnor U7115 (N_7115,N_7034,N_7039);
or U7116 (N_7116,N_7055,N_7089);
nand U7117 (N_7117,N_7070,N_7092);
and U7118 (N_7118,N_7001,N_7008);
nand U7119 (N_7119,N_7067,N_7096);
nand U7120 (N_7120,N_7038,N_7062);
nor U7121 (N_7121,N_7013,N_7094);
xnor U7122 (N_7122,N_7061,N_7068);
nand U7123 (N_7123,N_7014,N_7004);
and U7124 (N_7124,N_7025,N_7032);
nand U7125 (N_7125,N_7088,N_7046);
xor U7126 (N_7126,N_7018,N_7078);
xor U7127 (N_7127,N_7028,N_7097);
or U7128 (N_7128,N_7010,N_7037);
nand U7129 (N_7129,N_7022,N_7093);
nor U7130 (N_7130,N_7079,N_7076);
nor U7131 (N_7131,N_7006,N_7031);
or U7132 (N_7132,N_7023,N_7086);
and U7133 (N_7133,N_7049,N_7035);
xnor U7134 (N_7134,N_7020,N_7099);
xnor U7135 (N_7135,N_7077,N_7000);
nand U7136 (N_7136,N_7081,N_7091);
and U7137 (N_7137,N_7053,N_7003);
and U7138 (N_7138,N_7011,N_7052);
or U7139 (N_7139,N_7071,N_7063);
nor U7140 (N_7140,N_7026,N_7087);
or U7141 (N_7141,N_7069,N_7095);
nor U7142 (N_7142,N_7064,N_7072);
nand U7143 (N_7143,N_7041,N_7033);
and U7144 (N_7144,N_7080,N_7002);
or U7145 (N_7145,N_7057,N_7044);
and U7146 (N_7146,N_7005,N_7027);
nand U7147 (N_7147,N_7030,N_7012);
or U7148 (N_7148,N_7048,N_7075);
nand U7149 (N_7149,N_7015,N_7045);
nor U7150 (N_7150,N_7088,N_7056);
xnor U7151 (N_7151,N_7023,N_7048);
and U7152 (N_7152,N_7076,N_7088);
and U7153 (N_7153,N_7075,N_7083);
and U7154 (N_7154,N_7016,N_7064);
nor U7155 (N_7155,N_7076,N_7058);
nor U7156 (N_7156,N_7096,N_7034);
xnor U7157 (N_7157,N_7074,N_7003);
nor U7158 (N_7158,N_7062,N_7049);
and U7159 (N_7159,N_7056,N_7060);
nand U7160 (N_7160,N_7002,N_7075);
nand U7161 (N_7161,N_7022,N_7060);
or U7162 (N_7162,N_7082,N_7014);
nand U7163 (N_7163,N_7036,N_7082);
xor U7164 (N_7164,N_7033,N_7095);
and U7165 (N_7165,N_7024,N_7049);
and U7166 (N_7166,N_7053,N_7044);
xor U7167 (N_7167,N_7063,N_7037);
xnor U7168 (N_7168,N_7001,N_7000);
xnor U7169 (N_7169,N_7007,N_7093);
and U7170 (N_7170,N_7039,N_7077);
or U7171 (N_7171,N_7074,N_7072);
and U7172 (N_7172,N_7099,N_7027);
or U7173 (N_7173,N_7086,N_7034);
and U7174 (N_7174,N_7038,N_7081);
xor U7175 (N_7175,N_7074,N_7033);
nand U7176 (N_7176,N_7047,N_7067);
nor U7177 (N_7177,N_7016,N_7045);
nor U7178 (N_7178,N_7025,N_7089);
and U7179 (N_7179,N_7004,N_7081);
xor U7180 (N_7180,N_7088,N_7098);
xnor U7181 (N_7181,N_7067,N_7055);
and U7182 (N_7182,N_7025,N_7085);
nand U7183 (N_7183,N_7003,N_7008);
nand U7184 (N_7184,N_7061,N_7090);
xor U7185 (N_7185,N_7003,N_7052);
xnor U7186 (N_7186,N_7097,N_7024);
nand U7187 (N_7187,N_7090,N_7038);
or U7188 (N_7188,N_7086,N_7061);
xnor U7189 (N_7189,N_7094,N_7057);
or U7190 (N_7190,N_7094,N_7098);
nand U7191 (N_7191,N_7091,N_7082);
or U7192 (N_7192,N_7051,N_7097);
or U7193 (N_7193,N_7096,N_7040);
and U7194 (N_7194,N_7018,N_7023);
xor U7195 (N_7195,N_7082,N_7048);
xnor U7196 (N_7196,N_7049,N_7012);
and U7197 (N_7197,N_7080,N_7000);
or U7198 (N_7198,N_7079,N_7088);
nor U7199 (N_7199,N_7011,N_7077);
or U7200 (N_7200,N_7175,N_7111);
and U7201 (N_7201,N_7116,N_7119);
or U7202 (N_7202,N_7178,N_7196);
and U7203 (N_7203,N_7161,N_7127);
xor U7204 (N_7204,N_7185,N_7193);
xor U7205 (N_7205,N_7112,N_7136);
and U7206 (N_7206,N_7142,N_7129);
and U7207 (N_7207,N_7105,N_7192);
nand U7208 (N_7208,N_7152,N_7138);
and U7209 (N_7209,N_7160,N_7102);
nor U7210 (N_7210,N_7176,N_7191);
nand U7211 (N_7211,N_7155,N_7184);
or U7212 (N_7212,N_7110,N_7169);
nand U7213 (N_7213,N_7144,N_7179);
or U7214 (N_7214,N_7130,N_7123);
nand U7215 (N_7215,N_7114,N_7125);
or U7216 (N_7216,N_7139,N_7137);
nor U7217 (N_7217,N_7199,N_7104);
or U7218 (N_7218,N_7168,N_7162);
or U7219 (N_7219,N_7121,N_7132);
nand U7220 (N_7220,N_7189,N_7170);
and U7221 (N_7221,N_7126,N_7107);
and U7222 (N_7222,N_7157,N_7171);
nor U7223 (N_7223,N_7134,N_7145);
and U7224 (N_7224,N_7194,N_7147);
nand U7225 (N_7225,N_7124,N_7109);
and U7226 (N_7226,N_7198,N_7150);
nand U7227 (N_7227,N_7122,N_7131);
xnor U7228 (N_7228,N_7154,N_7167);
nor U7229 (N_7229,N_7135,N_7165);
and U7230 (N_7230,N_7172,N_7183);
and U7231 (N_7231,N_7186,N_7180);
xor U7232 (N_7232,N_7141,N_7118);
nor U7233 (N_7233,N_7158,N_7166);
nor U7234 (N_7234,N_7140,N_7181);
nand U7235 (N_7235,N_7115,N_7197);
nand U7236 (N_7236,N_7128,N_7108);
or U7237 (N_7237,N_7100,N_7177);
xor U7238 (N_7238,N_7190,N_7120);
xor U7239 (N_7239,N_7182,N_7148);
and U7240 (N_7240,N_7103,N_7164);
nor U7241 (N_7241,N_7163,N_7101);
nor U7242 (N_7242,N_7133,N_7156);
xor U7243 (N_7243,N_7188,N_7146);
xnor U7244 (N_7244,N_7174,N_7117);
xnor U7245 (N_7245,N_7151,N_7143);
or U7246 (N_7246,N_7153,N_7195);
or U7247 (N_7247,N_7173,N_7159);
or U7248 (N_7248,N_7113,N_7149);
nand U7249 (N_7249,N_7187,N_7106);
nand U7250 (N_7250,N_7110,N_7175);
or U7251 (N_7251,N_7153,N_7178);
and U7252 (N_7252,N_7169,N_7197);
nand U7253 (N_7253,N_7128,N_7147);
nor U7254 (N_7254,N_7166,N_7104);
nand U7255 (N_7255,N_7134,N_7152);
or U7256 (N_7256,N_7146,N_7187);
or U7257 (N_7257,N_7140,N_7143);
nor U7258 (N_7258,N_7102,N_7166);
xnor U7259 (N_7259,N_7146,N_7177);
nor U7260 (N_7260,N_7163,N_7139);
nor U7261 (N_7261,N_7153,N_7121);
xor U7262 (N_7262,N_7130,N_7159);
or U7263 (N_7263,N_7166,N_7112);
xor U7264 (N_7264,N_7186,N_7187);
nand U7265 (N_7265,N_7169,N_7142);
nor U7266 (N_7266,N_7175,N_7145);
nor U7267 (N_7267,N_7176,N_7199);
and U7268 (N_7268,N_7134,N_7198);
or U7269 (N_7269,N_7108,N_7106);
nor U7270 (N_7270,N_7199,N_7185);
or U7271 (N_7271,N_7104,N_7115);
or U7272 (N_7272,N_7114,N_7188);
nor U7273 (N_7273,N_7153,N_7130);
and U7274 (N_7274,N_7162,N_7113);
nand U7275 (N_7275,N_7108,N_7123);
nor U7276 (N_7276,N_7158,N_7177);
xnor U7277 (N_7277,N_7111,N_7163);
nand U7278 (N_7278,N_7134,N_7151);
nand U7279 (N_7279,N_7107,N_7185);
and U7280 (N_7280,N_7196,N_7156);
xnor U7281 (N_7281,N_7138,N_7114);
xnor U7282 (N_7282,N_7121,N_7128);
or U7283 (N_7283,N_7195,N_7179);
and U7284 (N_7284,N_7158,N_7180);
nor U7285 (N_7285,N_7179,N_7112);
xnor U7286 (N_7286,N_7151,N_7146);
nand U7287 (N_7287,N_7132,N_7152);
nor U7288 (N_7288,N_7144,N_7134);
or U7289 (N_7289,N_7110,N_7170);
and U7290 (N_7290,N_7176,N_7182);
or U7291 (N_7291,N_7139,N_7118);
or U7292 (N_7292,N_7160,N_7191);
nand U7293 (N_7293,N_7175,N_7102);
and U7294 (N_7294,N_7120,N_7108);
nor U7295 (N_7295,N_7151,N_7187);
xor U7296 (N_7296,N_7192,N_7164);
and U7297 (N_7297,N_7167,N_7159);
or U7298 (N_7298,N_7198,N_7100);
and U7299 (N_7299,N_7119,N_7102);
nand U7300 (N_7300,N_7200,N_7275);
nand U7301 (N_7301,N_7251,N_7206);
nand U7302 (N_7302,N_7269,N_7262);
or U7303 (N_7303,N_7268,N_7236);
nor U7304 (N_7304,N_7221,N_7224);
nor U7305 (N_7305,N_7225,N_7226);
nand U7306 (N_7306,N_7273,N_7228);
or U7307 (N_7307,N_7218,N_7209);
or U7308 (N_7308,N_7292,N_7213);
nor U7309 (N_7309,N_7238,N_7253);
xor U7310 (N_7310,N_7286,N_7239);
nor U7311 (N_7311,N_7289,N_7274);
xor U7312 (N_7312,N_7246,N_7223);
xor U7313 (N_7313,N_7235,N_7281);
or U7314 (N_7314,N_7288,N_7214);
nand U7315 (N_7315,N_7242,N_7215);
and U7316 (N_7316,N_7266,N_7270);
nor U7317 (N_7317,N_7222,N_7276);
xor U7318 (N_7318,N_7207,N_7241);
or U7319 (N_7319,N_7243,N_7201);
xor U7320 (N_7320,N_7227,N_7202);
nand U7321 (N_7321,N_7231,N_7219);
nand U7322 (N_7322,N_7260,N_7217);
xor U7323 (N_7323,N_7257,N_7296);
xor U7324 (N_7324,N_7264,N_7234);
and U7325 (N_7325,N_7252,N_7232);
xnor U7326 (N_7326,N_7290,N_7229);
nand U7327 (N_7327,N_7263,N_7267);
and U7328 (N_7328,N_7282,N_7250);
and U7329 (N_7329,N_7259,N_7255);
nand U7330 (N_7330,N_7240,N_7298);
and U7331 (N_7331,N_7287,N_7204);
xor U7332 (N_7332,N_7203,N_7244);
and U7333 (N_7333,N_7271,N_7210);
and U7334 (N_7334,N_7258,N_7277);
and U7335 (N_7335,N_7299,N_7297);
nor U7336 (N_7336,N_7249,N_7293);
xnor U7337 (N_7337,N_7285,N_7237);
nand U7338 (N_7338,N_7256,N_7265);
xor U7339 (N_7339,N_7254,N_7248);
and U7340 (N_7340,N_7212,N_7230);
and U7341 (N_7341,N_7233,N_7280);
or U7342 (N_7342,N_7294,N_7278);
or U7343 (N_7343,N_7220,N_7283);
and U7344 (N_7344,N_7279,N_7205);
nor U7345 (N_7345,N_7216,N_7208);
and U7346 (N_7346,N_7247,N_7211);
nand U7347 (N_7347,N_7245,N_7295);
nand U7348 (N_7348,N_7291,N_7272);
or U7349 (N_7349,N_7261,N_7284);
and U7350 (N_7350,N_7275,N_7298);
or U7351 (N_7351,N_7274,N_7232);
nor U7352 (N_7352,N_7257,N_7266);
and U7353 (N_7353,N_7273,N_7271);
nand U7354 (N_7354,N_7296,N_7222);
and U7355 (N_7355,N_7245,N_7217);
nor U7356 (N_7356,N_7256,N_7233);
nand U7357 (N_7357,N_7205,N_7225);
and U7358 (N_7358,N_7287,N_7291);
nor U7359 (N_7359,N_7252,N_7228);
xnor U7360 (N_7360,N_7202,N_7223);
xnor U7361 (N_7361,N_7230,N_7282);
nor U7362 (N_7362,N_7220,N_7260);
or U7363 (N_7363,N_7256,N_7214);
and U7364 (N_7364,N_7256,N_7242);
or U7365 (N_7365,N_7269,N_7290);
or U7366 (N_7366,N_7271,N_7213);
and U7367 (N_7367,N_7211,N_7280);
nand U7368 (N_7368,N_7278,N_7232);
or U7369 (N_7369,N_7201,N_7280);
xnor U7370 (N_7370,N_7224,N_7294);
nor U7371 (N_7371,N_7268,N_7273);
xor U7372 (N_7372,N_7253,N_7283);
xnor U7373 (N_7373,N_7295,N_7208);
and U7374 (N_7374,N_7260,N_7225);
and U7375 (N_7375,N_7210,N_7221);
xnor U7376 (N_7376,N_7288,N_7220);
nand U7377 (N_7377,N_7243,N_7296);
or U7378 (N_7378,N_7271,N_7250);
nor U7379 (N_7379,N_7241,N_7262);
nor U7380 (N_7380,N_7277,N_7231);
nor U7381 (N_7381,N_7256,N_7273);
or U7382 (N_7382,N_7223,N_7242);
xnor U7383 (N_7383,N_7247,N_7280);
nand U7384 (N_7384,N_7263,N_7254);
and U7385 (N_7385,N_7294,N_7211);
or U7386 (N_7386,N_7222,N_7250);
and U7387 (N_7387,N_7285,N_7215);
nor U7388 (N_7388,N_7204,N_7262);
nand U7389 (N_7389,N_7285,N_7271);
xnor U7390 (N_7390,N_7299,N_7248);
and U7391 (N_7391,N_7296,N_7206);
nor U7392 (N_7392,N_7222,N_7221);
or U7393 (N_7393,N_7213,N_7227);
xnor U7394 (N_7394,N_7292,N_7295);
nor U7395 (N_7395,N_7221,N_7213);
and U7396 (N_7396,N_7269,N_7288);
and U7397 (N_7397,N_7203,N_7276);
nor U7398 (N_7398,N_7290,N_7286);
nand U7399 (N_7399,N_7294,N_7247);
nand U7400 (N_7400,N_7319,N_7317);
and U7401 (N_7401,N_7325,N_7322);
and U7402 (N_7402,N_7375,N_7369);
and U7403 (N_7403,N_7306,N_7347);
nand U7404 (N_7404,N_7393,N_7376);
and U7405 (N_7405,N_7320,N_7340);
nand U7406 (N_7406,N_7372,N_7323);
nor U7407 (N_7407,N_7315,N_7331);
nand U7408 (N_7408,N_7396,N_7371);
xnor U7409 (N_7409,N_7381,N_7316);
or U7410 (N_7410,N_7353,N_7350);
or U7411 (N_7411,N_7355,N_7344);
xnor U7412 (N_7412,N_7332,N_7337);
nand U7413 (N_7413,N_7309,N_7326);
nor U7414 (N_7414,N_7310,N_7394);
or U7415 (N_7415,N_7362,N_7374);
xnor U7416 (N_7416,N_7330,N_7370);
or U7417 (N_7417,N_7358,N_7399);
xor U7418 (N_7418,N_7377,N_7302);
and U7419 (N_7419,N_7389,N_7367);
nand U7420 (N_7420,N_7334,N_7307);
xor U7421 (N_7421,N_7318,N_7301);
nor U7422 (N_7422,N_7333,N_7342);
nand U7423 (N_7423,N_7305,N_7314);
nand U7424 (N_7424,N_7339,N_7395);
nor U7425 (N_7425,N_7388,N_7397);
or U7426 (N_7426,N_7359,N_7364);
or U7427 (N_7427,N_7329,N_7357);
xor U7428 (N_7428,N_7365,N_7343);
or U7429 (N_7429,N_7383,N_7386);
nor U7430 (N_7430,N_7308,N_7335);
and U7431 (N_7431,N_7327,N_7382);
or U7432 (N_7432,N_7352,N_7368);
and U7433 (N_7433,N_7321,N_7354);
or U7434 (N_7434,N_7336,N_7385);
and U7435 (N_7435,N_7360,N_7348);
and U7436 (N_7436,N_7378,N_7384);
or U7437 (N_7437,N_7390,N_7380);
xor U7438 (N_7438,N_7303,N_7338);
and U7439 (N_7439,N_7324,N_7373);
or U7440 (N_7440,N_7363,N_7351);
xor U7441 (N_7441,N_7328,N_7341);
nor U7442 (N_7442,N_7387,N_7311);
nand U7443 (N_7443,N_7379,N_7345);
nor U7444 (N_7444,N_7304,N_7398);
xor U7445 (N_7445,N_7349,N_7300);
xor U7446 (N_7446,N_7361,N_7313);
xor U7447 (N_7447,N_7356,N_7346);
or U7448 (N_7448,N_7392,N_7366);
nand U7449 (N_7449,N_7391,N_7312);
nor U7450 (N_7450,N_7377,N_7394);
nand U7451 (N_7451,N_7354,N_7335);
nand U7452 (N_7452,N_7387,N_7352);
nor U7453 (N_7453,N_7337,N_7348);
nor U7454 (N_7454,N_7397,N_7375);
and U7455 (N_7455,N_7374,N_7364);
nand U7456 (N_7456,N_7362,N_7333);
and U7457 (N_7457,N_7386,N_7398);
nand U7458 (N_7458,N_7386,N_7357);
and U7459 (N_7459,N_7346,N_7382);
or U7460 (N_7460,N_7390,N_7360);
nand U7461 (N_7461,N_7336,N_7369);
xor U7462 (N_7462,N_7363,N_7326);
and U7463 (N_7463,N_7319,N_7354);
nand U7464 (N_7464,N_7324,N_7333);
nor U7465 (N_7465,N_7362,N_7375);
nand U7466 (N_7466,N_7381,N_7340);
nor U7467 (N_7467,N_7390,N_7373);
or U7468 (N_7468,N_7310,N_7375);
and U7469 (N_7469,N_7397,N_7354);
nor U7470 (N_7470,N_7334,N_7318);
nor U7471 (N_7471,N_7333,N_7338);
or U7472 (N_7472,N_7360,N_7355);
xnor U7473 (N_7473,N_7398,N_7347);
nor U7474 (N_7474,N_7336,N_7305);
and U7475 (N_7475,N_7359,N_7382);
nand U7476 (N_7476,N_7334,N_7381);
xnor U7477 (N_7477,N_7391,N_7356);
xor U7478 (N_7478,N_7314,N_7329);
xor U7479 (N_7479,N_7330,N_7302);
nor U7480 (N_7480,N_7341,N_7392);
or U7481 (N_7481,N_7393,N_7319);
nor U7482 (N_7482,N_7324,N_7326);
or U7483 (N_7483,N_7392,N_7301);
and U7484 (N_7484,N_7377,N_7386);
nor U7485 (N_7485,N_7383,N_7362);
or U7486 (N_7486,N_7363,N_7368);
or U7487 (N_7487,N_7329,N_7379);
nand U7488 (N_7488,N_7382,N_7336);
xnor U7489 (N_7489,N_7351,N_7352);
nand U7490 (N_7490,N_7342,N_7318);
or U7491 (N_7491,N_7374,N_7350);
and U7492 (N_7492,N_7303,N_7382);
nor U7493 (N_7493,N_7360,N_7381);
nand U7494 (N_7494,N_7330,N_7340);
nand U7495 (N_7495,N_7382,N_7330);
and U7496 (N_7496,N_7321,N_7318);
xor U7497 (N_7497,N_7304,N_7390);
nor U7498 (N_7498,N_7357,N_7362);
nand U7499 (N_7499,N_7349,N_7345);
xnor U7500 (N_7500,N_7484,N_7437);
nand U7501 (N_7501,N_7433,N_7499);
or U7502 (N_7502,N_7400,N_7407);
xnor U7503 (N_7503,N_7451,N_7424);
nor U7504 (N_7504,N_7419,N_7434);
nor U7505 (N_7505,N_7438,N_7413);
and U7506 (N_7506,N_7473,N_7480);
and U7507 (N_7507,N_7429,N_7493);
nand U7508 (N_7508,N_7445,N_7488);
nand U7509 (N_7509,N_7471,N_7491);
or U7510 (N_7510,N_7494,N_7450);
xor U7511 (N_7511,N_7467,N_7464);
nor U7512 (N_7512,N_7418,N_7486);
nand U7513 (N_7513,N_7420,N_7447);
nand U7514 (N_7514,N_7468,N_7401);
xnor U7515 (N_7515,N_7474,N_7446);
or U7516 (N_7516,N_7430,N_7477);
nand U7517 (N_7517,N_7470,N_7402);
or U7518 (N_7518,N_7492,N_7426);
nor U7519 (N_7519,N_7404,N_7485);
or U7520 (N_7520,N_7479,N_7403);
nor U7521 (N_7521,N_7476,N_7462);
xor U7522 (N_7522,N_7482,N_7469);
and U7523 (N_7523,N_7481,N_7455);
or U7524 (N_7524,N_7472,N_7435);
nor U7525 (N_7525,N_7457,N_7478);
xor U7526 (N_7526,N_7463,N_7495);
or U7527 (N_7527,N_7456,N_7496);
nand U7528 (N_7528,N_7436,N_7415);
xnor U7529 (N_7529,N_7449,N_7459);
and U7530 (N_7530,N_7440,N_7483);
and U7531 (N_7531,N_7417,N_7416);
nor U7532 (N_7532,N_7422,N_7461);
or U7533 (N_7533,N_7412,N_7411);
nand U7534 (N_7534,N_7453,N_7497);
nor U7535 (N_7535,N_7409,N_7425);
and U7536 (N_7536,N_7405,N_7489);
nand U7537 (N_7537,N_7490,N_7427);
nand U7538 (N_7538,N_7465,N_7458);
nor U7539 (N_7539,N_7439,N_7421);
xor U7540 (N_7540,N_7414,N_7444);
nand U7541 (N_7541,N_7406,N_7475);
nand U7542 (N_7542,N_7441,N_7466);
or U7543 (N_7543,N_7448,N_7410);
nand U7544 (N_7544,N_7442,N_7423);
nand U7545 (N_7545,N_7487,N_7432);
nor U7546 (N_7546,N_7454,N_7431);
nand U7547 (N_7547,N_7498,N_7443);
nor U7548 (N_7548,N_7408,N_7460);
xor U7549 (N_7549,N_7428,N_7452);
nor U7550 (N_7550,N_7449,N_7424);
xnor U7551 (N_7551,N_7441,N_7481);
and U7552 (N_7552,N_7441,N_7429);
or U7553 (N_7553,N_7457,N_7490);
nor U7554 (N_7554,N_7478,N_7490);
or U7555 (N_7555,N_7426,N_7458);
or U7556 (N_7556,N_7437,N_7486);
or U7557 (N_7557,N_7422,N_7471);
xnor U7558 (N_7558,N_7495,N_7450);
nor U7559 (N_7559,N_7458,N_7414);
nand U7560 (N_7560,N_7431,N_7466);
xnor U7561 (N_7561,N_7413,N_7421);
nand U7562 (N_7562,N_7404,N_7433);
nor U7563 (N_7563,N_7428,N_7442);
or U7564 (N_7564,N_7471,N_7443);
and U7565 (N_7565,N_7427,N_7464);
nand U7566 (N_7566,N_7419,N_7429);
xor U7567 (N_7567,N_7468,N_7421);
nor U7568 (N_7568,N_7438,N_7475);
xor U7569 (N_7569,N_7455,N_7411);
xor U7570 (N_7570,N_7452,N_7409);
nor U7571 (N_7571,N_7427,N_7496);
xnor U7572 (N_7572,N_7431,N_7427);
xnor U7573 (N_7573,N_7426,N_7479);
xor U7574 (N_7574,N_7420,N_7459);
or U7575 (N_7575,N_7451,N_7438);
xnor U7576 (N_7576,N_7425,N_7424);
or U7577 (N_7577,N_7440,N_7474);
nand U7578 (N_7578,N_7459,N_7400);
nor U7579 (N_7579,N_7472,N_7465);
xor U7580 (N_7580,N_7478,N_7499);
nand U7581 (N_7581,N_7493,N_7432);
nor U7582 (N_7582,N_7464,N_7412);
or U7583 (N_7583,N_7414,N_7451);
nor U7584 (N_7584,N_7483,N_7412);
xnor U7585 (N_7585,N_7417,N_7460);
and U7586 (N_7586,N_7460,N_7443);
nand U7587 (N_7587,N_7428,N_7444);
nand U7588 (N_7588,N_7424,N_7489);
xnor U7589 (N_7589,N_7440,N_7482);
or U7590 (N_7590,N_7440,N_7467);
or U7591 (N_7591,N_7408,N_7458);
nand U7592 (N_7592,N_7443,N_7421);
nand U7593 (N_7593,N_7449,N_7451);
xnor U7594 (N_7594,N_7412,N_7429);
xor U7595 (N_7595,N_7409,N_7432);
or U7596 (N_7596,N_7498,N_7478);
or U7597 (N_7597,N_7460,N_7475);
xnor U7598 (N_7598,N_7493,N_7480);
or U7599 (N_7599,N_7457,N_7400);
or U7600 (N_7600,N_7566,N_7516);
xnor U7601 (N_7601,N_7553,N_7544);
nor U7602 (N_7602,N_7571,N_7537);
and U7603 (N_7603,N_7554,N_7533);
nand U7604 (N_7604,N_7555,N_7560);
or U7605 (N_7605,N_7584,N_7526);
or U7606 (N_7606,N_7540,N_7502);
and U7607 (N_7607,N_7585,N_7565);
or U7608 (N_7608,N_7579,N_7569);
xnor U7609 (N_7609,N_7511,N_7534);
nand U7610 (N_7610,N_7589,N_7590);
xor U7611 (N_7611,N_7514,N_7536);
or U7612 (N_7612,N_7577,N_7532);
xnor U7613 (N_7613,N_7591,N_7558);
or U7614 (N_7614,N_7559,N_7500);
and U7615 (N_7615,N_7586,N_7598);
and U7616 (N_7616,N_7570,N_7547);
nor U7617 (N_7617,N_7568,N_7531);
nand U7618 (N_7618,N_7517,N_7510);
nand U7619 (N_7619,N_7563,N_7539);
or U7620 (N_7620,N_7567,N_7541);
xnor U7621 (N_7621,N_7529,N_7546);
nand U7622 (N_7622,N_7506,N_7576);
or U7623 (N_7623,N_7599,N_7521);
nor U7624 (N_7624,N_7513,N_7582);
xnor U7625 (N_7625,N_7587,N_7538);
or U7626 (N_7626,N_7549,N_7575);
nor U7627 (N_7627,N_7520,N_7505);
xor U7628 (N_7628,N_7581,N_7518);
nor U7629 (N_7629,N_7530,N_7524);
xnor U7630 (N_7630,N_7528,N_7527);
xnor U7631 (N_7631,N_7550,N_7504);
xnor U7632 (N_7632,N_7597,N_7583);
and U7633 (N_7633,N_7552,N_7535);
nor U7634 (N_7634,N_7522,N_7557);
xnor U7635 (N_7635,N_7562,N_7595);
nor U7636 (N_7636,N_7525,N_7551);
xor U7637 (N_7637,N_7503,N_7542);
nand U7638 (N_7638,N_7507,N_7561);
nand U7639 (N_7639,N_7578,N_7593);
nand U7640 (N_7640,N_7512,N_7580);
nand U7641 (N_7641,N_7523,N_7574);
or U7642 (N_7642,N_7572,N_7509);
or U7643 (N_7643,N_7556,N_7543);
nor U7644 (N_7644,N_7588,N_7573);
or U7645 (N_7645,N_7519,N_7501);
nor U7646 (N_7646,N_7545,N_7596);
xor U7647 (N_7647,N_7592,N_7515);
nand U7648 (N_7648,N_7564,N_7548);
nor U7649 (N_7649,N_7594,N_7508);
nand U7650 (N_7650,N_7515,N_7522);
nor U7651 (N_7651,N_7526,N_7504);
and U7652 (N_7652,N_7552,N_7527);
and U7653 (N_7653,N_7529,N_7531);
or U7654 (N_7654,N_7577,N_7515);
nand U7655 (N_7655,N_7523,N_7593);
nand U7656 (N_7656,N_7562,N_7594);
xor U7657 (N_7657,N_7554,N_7564);
and U7658 (N_7658,N_7590,N_7584);
xor U7659 (N_7659,N_7551,N_7589);
nor U7660 (N_7660,N_7545,N_7550);
xnor U7661 (N_7661,N_7543,N_7582);
nor U7662 (N_7662,N_7515,N_7505);
nand U7663 (N_7663,N_7530,N_7558);
nor U7664 (N_7664,N_7524,N_7533);
xnor U7665 (N_7665,N_7507,N_7567);
nand U7666 (N_7666,N_7542,N_7505);
or U7667 (N_7667,N_7586,N_7552);
or U7668 (N_7668,N_7537,N_7511);
or U7669 (N_7669,N_7521,N_7500);
or U7670 (N_7670,N_7504,N_7534);
nand U7671 (N_7671,N_7596,N_7583);
nand U7672 (N_7672,N_7526,N_7589);
nand U7673 (N_7673,N_7561,N_7569);
xnor U7674 (N_7674,N_7567,N_7583);
nand U7675 (N_7675,N_7576,N_7505);
and U7676 (N_7676,N_7578,N_7527);
xor U7677 (N_7677,N_7598,N_7515);
and U7678 (N_7678,N_7564,N_7593);
and U7679 (N_7679,N_7584,N_7542);
nand U7680 (N_7680,N_7532,N_7553);
and U7681 (N_7681,N_7544,N_7537);
and U7682 (N_7682,N_7507,N_7563);
or U7683 (N_7683,N_7526,N_7547);
or U7684 (N_7684,N_7529,N_7535);
and U7685 (N_7685,N_7591,N_7543);
nor U7686 (N_7686,N_7583,N_7561);
or U7687 (N_7687,N_7597,N_7585);
xnor U7688 (N_7688,N_7562,N_7549);
xnor U7689 (N_7689,N_7532,N_7583);
nor U7690 (N_7690,N_7566,N_7500);
and U7691 (N_7691,N_7579,N_7595);
and U7692 (N_7692,N_7552,N_7537);
or U7693 (N_7693,N_7584,N_7565);
nand U7694 (N_7694,N_7521,N_7505);
nor U7695 (N_7695,N_7538,N_7545);
or U7696 (N_7696,N_7570,N_7521);
xnor U7697 (N_7697,N_7521,N_7522);
nor U7698 (N_7698,N_7564,N_7546);
xnor U7699 (N_7699,N_7524,N_7594);
nor U7700 (N_7700,N_7642,N_7639);
nand U7701 (N_7701,N_7647,N_7622);
and U7702 (N_7702,N_7634,N_7689);
xnor U7703 (N_7703,N_7625,N_7605);
or U7704 (N_7704,N_7648,N_7602);
nand U7705 (N_7705,N_7619,N_7617);
nor U7706 (N_7706,N_7646,N_7669);
nor U7707 (N_7707,N_7684,N_7601);
and U7708 (N_7708,N_7632,N_7627);
nor U7709 (N_7709,N_7638,N_7628);
nand U7710 (N_7710,N_7685,N_7673);
xor U7711 (N_7711,N_7616,N_7676);
or U7712 (N_7712,N_7658,N_7623);
xnor U7713 (N_7713,N_7645,N_7699);
or U7714 (N_7714,N_7644,N_7614);
xnor U7715 (N_7715,N_7697,N_7670);
xnor U7716 (N_7716,N_7678,N_7694);
nor U7717 (N_7717,N_7615,N_7629);
xnor U7718 (N_7718,N_7661,N_7611);
xor U7719 (N_7719,N_7663,N_7640);
and U7720 (N_7720,N_7613,N_7696);
and U7721 (N_7721,N_7677,N_7651);
xnor U7722 (N_7722,N_7695,N_7687);
or U7723 (N_7723,N_7655,N_7679);
nor U7724 (N_7724,N_7667,N_7603);
nor U7725 (N_7725,N_7660,N_7652);
and U7726 (N_7726,N_7693,N_7688);
xor U7727 (N_7727,N_7609,N_7630);
or U7728 (N_7728,N_7683,N_7620);
nor U7729 (N_7729,N_7633,N_7656);
nand U7730 (N_7730,N_7672,N_7682);
nor U7731 (N_7731,N_7659,N_7621);
xnor U7732 (N_7732,N_7653,N_7604);
nor U7733 (N_7733,N_7635,N_7649);
nor U7734 (N_7734,N_7666,N_7691);
xor U7735 (N_7735,N_7610,N_7641);
nor U7736 (N_7736,N_7607,N_7626);
nand U7737 (N_7737,N_7698,N_7624);
xnor U7738 (N_7738,N_7657,N_7664);
and U7739 (N_7739,N_7650,N_7637);
nor U7740 (N_7740,N_7631,N_7671);
or U7741 (N_7741,N_7681,N_7668);
nand U7742 (N_7742,N_7686,N_7680);
nand U7743 (N_7743,N_7618,N_7690);
nor U7744 (N_7744,N_7606,N_7692);
and U7745 (N_7745,N_7612,N_7675);
or U7746 (N_7746,N_7654,N_7608);
nor U7747 (N_7747,N_7662,N_7665);
and U7748 (N_7748,N_7674,N_7600);
or U7749 (N_7749,N_7643,N_7636);
or U7750 (N_7750,N_7692,N_7630);
nor U7751 (N_7751,N_7646,N_7695);
or U7752 (N_7752,N_7627,N_7631);
xnor U7753 (N_7753,N_7669,N_7643);
nand U7754 (N_7754,N_7669,N_7632);
and U7755 (N_7755,N_7611,N_7673);
and U7756 (N_7756,N_7603,N_7676);
nand U7757 (N_7757,N_7655,N_7611);
nand U7758 (N_7758,N_7699,N_7644);
nor U7759 (N_7759,N_7673,N_7663);
or U7760 (N_7760,N_7610,N_7699);
nor U7761 (N_7761,N_7694,N_7651);
xnor U7762 (N_7762,N_7649,N_7654);
xnor U7763 (N_7763,N_7666,N_7697);
or U7764 (N_7764,N_7632,N_7675);
xor U7765 (N_7765,N_7667,N_7629);
nand U7766 (N_7766,N_7697,N_7682);
and U7767 (N_7767,N_7608,N_7684);
nand U7768 (N_7768,N_7678,N_7646);
nand U7769 (N_7769,N_7638,N_7694);
xor U7770 (N_7770,N_7674,N_7659);
xnor U7771 (N_7771,N_7650,N_7609);
or U7772 (N_7772,N_7632,N_7639);
nand U7773 (N_7773,N_7617,N_7602);
or U7774 (N_7774,N_7676,N_7692);
nand U7775 (N_7775,N_7671,N_7678);
nand U7776 (N_7776,N_7625,N_7684);
or U7777 (N_7777,N_7610,N_7652);
nor U7778 (N_7778,N_7613,N_7633);
or U7779 (N_7779,N_7628,N_7683);
or U7780 (N_7780,N_7692,N_7684);
or U7781 (N_7781,N_7631,N_7602);
xor U7782 (N_7782,N_7687,N_7615);
or U7783 (N_7783,N_7699,N_7623);
or U7784 (N_7784,N_7676,N_7695);
or U7785 (N_7785,N_7624,N_7645);
or U7786 (N_7786,N_7687,N_7662);
or U7787 (N_7787,N_7682,N_7694);
and U7788 (N_7788,N_7620,N_7628);
and U7789 (N_7789,N_7606,N_7687);
nor U7790 (N_7790,N_7618,N_7681);
nor U7791 (N_7791,N_7683,N_7694);
xnor U7792 (N_7792,N_7693,N_7672);
or U7793 (N_7793,N_7668,N_7631);
and U7794 (N_7794,N_7682,N_7681);
and U7795 (N_7795,N_7648,N_7618);
xor U7796 (N_7796,N_7619,N_7669);
xor U7797 (N_7797,N_7650,N_7657);
xnor U7798 (N_7798,N_7651,N_7690);
and U7799 (N_7799,N_7697,N_7622);
or U7800 (N_7800,N_7722,N_7735);
nor U7801 (N_7801,N_7756,N_7742);
and U7802 (N_7802,N_7749,N_7733);
or U7803 (N_7803,N_7720,N_7762);
xnor U7804 (N_7804,N_7753,N_7763);
or U7805 (N_7805,N_7715,N_7711);
xnor U7806 (N_7806,N_7752,N_7743);
xnor U7807 (N_7807,N_7773,N_7751);
nand U7808 (N_7808,N_7701,N_7709);
or U7809 (N_7809,N_7794,N_7737);
or U7810 (N_7810,N_7727,N_7769);
nor U7811 (N_7811,N_7778,N_7780);
or U7812 (N_7812,N_7775,N_7700);
or U7813 (N_7813,N_7790,N_7706);
nor U7814 (N_7814,N_7746,N_7719);
or U7815 (N_7815,N_7772,N_7789);
and U7816 (N_7816,N_7717,N_7765);
nand U7817 (N_7817,N_7758,N_7787);
and U7818 (N_7818,N_7738,N_7740);
nor U7819 (N_7819,N_7708,N_7707);
xnor U7820 (N_7820,N_7736,N_7766);
nor U7821 (N_7821,N_7705,N_7741);
or U7822 (N_7822,N_7729,N_7712);
and U7823 (N_7823,N_7797,N_7760);
nand U7824 (N_7824,N_7776,N_7748);
nand U7825 (N_7825,N_7713,N_7774);
and U7826 (N_7826,N_7771,N_7783);
nand U7827 (N_7827,N_7770,N_7728);
or U7828 (N_7828,N_7744,N_7721);
and U7829 (N_7829,N_7714,N_7796);
nand U7830 (N_7830,N_7734,N_7750);
nand U7831 (N_7831,N_7759,N_7730);
and U7832 (N_7832,N_7795,N_7731);
nor U7833 (N_7833,N_7739,N_7723);
or U7834 (N_7834,N_7799,N_7798);
xor U7835 (N_7835,N_7767,N_7732);
and U7836 (N_7836,N_7724,N_7784);
xor U7837 (N_7837,N_7702,N_7768);
or U7838 (N_7838,N_7777,N_7716);
xnor U7839 (N_7839,N_7710,N_7703);
nor U7840 (N_7840,N_7747,N_7726);
nor U7841 (N_7841,N_7788,N_7725);
nor U7842 (N_7842,N_7791,N_7718);
and U7843 (N_7843,N_7745,N_7781);
or U7844 (N_7844,N_7764,N_7754);
xnor U7845 (N_7845,N_7792,N_7785);
xor U7846 (N_7846,N_7779,N_7782);
or U7847 (N_7847,N_7704,N_7793);
and U7848 (N_7848,N_7757,N_7786);
xnor U7849 (N_7849,N_7755,N_7761);
nand U7850 (N_7850,N_7759,N_7756);
or U7851 (N_7851,N_7761,N_7767);
nand U7852 (N_7852,N_7793,N_7767);
xor U7853 (N_7853,N_7764,N_7714);
and U7854 (N_7854,N_7752,N_7756);
or U7855 (N_7855,N_7750,N_7783);
or U7856 (N_7856,N_7745,N_7744);
nand U7857 (N_7857,N_7775,N_7701);
nor U7858 (N_7858,N_7712,N_7719);
nor U7859 (N_7859,N_7733,N_7751);
and U7860 (N_7860,N_7751,N_7763);
or U7861 (N_7861,N_7713,N_7704);
or U7862 (N_7862,N_7773,N_7703);
nor U7863 (N_7863,N_7730,N_7764);
or U7864 (N_7864,N_7718,N_7780);
or U7865 (N_7865,N_7792,N_7736);
nand U7866 (N_7866,N_7778,N_7709);
nor U7867 (N_7867,N_7790,N_7791);
or U7868 (N_7868,N_7709,N_7728);
nand U7869 (N_7869,N_7793,N_7757);
nor U7870 (N_7870,N_7723,N_7708);
xor U7871 (N_7871,N_7784,N_7773);
or U7872 (N_7872,N_7728,N_7711);
or U7873 (N_7873,N_7786,N_7798);
nor U7874 (N_7874,N_7710,N_7713);
or U7875 (N_7875,N_7755,N_7780);
nor U7876 (N_7876,N_7770,N_7784);
and U7877 (N_7877,N_7742,N_7715);
nand U7878 (N_7878,N_7755,N_7704);
nor U7879 (N_7879,N_7705,N_7724);
nand U7880 (N_7880,N_7763,N_7799);
xor U7881 (N_7881,N_7747,N_7775);
and U7882 (N_7882,N_7722,N_7723);
nand U7883 (N_7883,N_7794,N_7742);
and U7884 (N_7884,N_7767,N_7704);
nand U7885 (N_7885,N_7744,N_7776);
and U7886 (N_7886,N_7725,N_7711);
xnor U7887 (N_7887,N_7710,N_7717);
nand U7888 (N_7888,N_7739,N_7726);
nor U7889 (N_7889,N_7727,N_7720);
or U7890 (N_7890,N_7740,N_7792);
xor U7891 (N_7891,N_7732,N_7792);
xor U7892 (N_7892,N_7736,N_7764);
nor U7893 (N_7893,N_7779,N_7799);
nand U7894 (N_7894,N_7724,N_7753);
and U7895 (N_7895,N_7780,N_7725);
nor U7896 (N_7896,N_7768,N_7738);
or U7897 (N_7897,N_7758,N_7710);
and U7898 (N_7898,N_7750,N_7728);
and U7899 (N_7899,N_7739,N_7760);
nand U7900 (N_7900,N_7841,N_7887);
nand U7901 (N_7901,N_7800,N_7861);
nand U7902 (N_7902,N_7806,N_7865);
nand U7903 (N_7903,N_7829,N_7888);
xor U7904 (N_7904,N_7803,N_7896);
xnor U7905 (N_7905,N_7847,N_7895);
nand U7906 (N_7906,N_7838,N_7801);
and U7907 (N_7907,N_7851,N_7818);
xnor U7908 (N_7908,N_7884,N_7832);
nor U7909 (N_7909,N_7817,N_7805);
nor U7910 (N_7910,N_7849,N_7893);
and U7911 (N_7911,N_7837,N_7862);
nor U7912 (N_7912,N_7842,N_7811);
or U7913 (N_7913,N_7879,N_7894);
or U7914 (N_7914,N_7844,N_7857);
or U7915 (N_7915,N_7813,N_7814);
xnor U7916 (N_7916,N_7881,N_7886);
or U7917 (N_7917,N_7853,N_7872);
and U7918 (N_7918,N_7870,N_7822);
or U7919 (N_7919,N_7854,N_7874);
nand U7920 (N_7920,N_7812,N_7808);
xnor U7921 (N_7921,N_7880,N_7807);
or U7922 (N_7922,N_7864,N_7848);
nor U7923 (N_7923,N_7831,N_7897);
xnor U7924 (N_7924,N_7834,N_7873);
nor U7925 (N_7925,N_7875,N_7898);
xnor U7926 (N_7926,N_7821,N_7858);
or U7927 (N_7927,N_7869,N_7855);
and U7928 (N_7928,N_7892,N_7802);
or U7929 (N_7929,N_7816,N_7846);
xnor U7930 (N_7930,N_7840,N_7889);
or U7931 (N_7931,N_7859,N_7882);
and U7932 (N_7932,N_7827,N_7826);
and U7933 (N_7933,N_7876,N_7867);
or U7934 (N_7934,N_7883,N_7890);
nand U7935 (N_7935,N_7824,N_7899);
xor U7936 (N_7936,N_7843,N_7877);
nor U7937 (N_7937,N_7863,N_7856);
and U7938 (N_7938,N_7804,N_7885);
xnor U7939 (N_7939,N_7878,N_7825);
xor U7940 (N_7940,N_7835,N_7823);
or U7941 (N_7941,N_7839,N_7868);
or U7942 (N_7942,N_7819,N_7860);
nand U7943 (N_7943,N_7845,N_7866);
nand U7944 (N_7944,N_7850,N_7891);
nand U7945 (N_7945,N_7820,N_7809);
nor U7946 (N_7946,N_7836,N_7871);
or U7947 (N_7947,N_7828,N_7815);
xnor U7948 (N_7948,N_7833,N_7830);
and U7949 (N_7949,N_7852,N_7810);
and U7950 (N_7950,N_7876,N_7805);
nand U7951 (N_7951,N_7836,N_7832);
nor U7952 (N_7952,N_7828,N_7875);
nor U7953 (N_7953,N_7834,N_7824);
or U7954 (N_7954,N_7834,N_7804);
xnor U7955 (N_7955,N_7815,N_7802);
or U7956 (N_7956,N_7862,N_7839);
or U7957 (N_7957,N_7849,N_7844);
and U7958 (N_7958,N_7814,N_7809);
nor U7959 (N_7959,N_7866,N_7856);
nor U7960 (N_7960,N_7833,N_7866);
xnor U7961 (N_7961,N_7897,N_7880);
nor U7962 (N_7962,N_7844,N_7863);
and U7963 (N_7963,N_7847,N_7882);
nor U7964 (N_7964,N_7820,N_7803);
and U7965 (N_7965,N_7861,N_7815);
or U7966 (N_7966,N_7892,N_7824);
or U7967 (N_7967,N_7894,N_7842);
and U7968 (N_7968,N_7844,N_7833);
nand U7969 (N_7969,N_7829,N_7851);
xor U7970 (N_7970,N_7892,N_7817);
or U7971 (N_7971,N_7831,N_7833);
nand U7972 (N_7972,N_7865,N_7809);
and U7973 (N_7973,N_7819,N_7865);
and U7974 (N_7974,N_7856,N_7889);
and U7975 (N_7975,N_7899,N_7837);
xnor U7976 (N_7976,N_7868,N_7828);
and U7977 (N_7977,N_7842,N_7862);
or U7978 (N_7978,N_7879,N_7811);
nand U7979 (N_7979,N_7874,N_7898);
nor U7980 (N_7980,N_7817,N_7807);
nand U7981 (N_7981,N_7813,N_7899);
nor U7982 (N_7982,N_7815,N_7895);
nand U7983 (N_7983,N_7808,N_7816);
nand U7984 (N_7984,N_7816,N_7885);
nor U7985 (N_7985,N_7892,N_7875);
xor U7986 (N_7986,N_7848,N_7852);
and U7987 (N_7987,N_7863,N_7818);
xnor U7988 (N_7988,N_7868,N_7833);
xor U7989 (N_7989,N_7831,N_7809);
xnor U7990 (N_7990,N_7860,N_7891);
and U7991 (N_7991,N_7892,N_7822);
nor U7992 (N_7992,N_7865,N_7859);
or U7993 (N_7993,N_7809,N_7825);
nor U7994 (N_7994,N_7830,N_7829);
or U7995 (N_7995,N_7844,N_7838);
nand U7996 (N_7996,N_7868,N_7846);
nor U7997 (N_7997,N_7820,N_7899);
and U7998 (N_7998,N_7809,N_7810);
or U7999 (N_7999,N_7885,N_7801);
nand U8000 (N_8000,N_7993,N_7916);
and U8001 (N_8001,N_7981,N_7920);
nand U8002 (N_8002,N_7901,N_7986);
nand U8003 (N_8003,N_7951,N_7938);
or U8004 (N_8004,N_7962,N_7989);
nand U8005 (N_8005,N_7964,N_7982);
nand U8006 (N_8006,N_7996,N_7932);
nor U8007 (N_8007,N_7945,N_7966);
or U8008 (N_8008,N_7943,N_7912);
nor U8009 (N_8009,N_7934,N_7969);
nor U8010 (N_8010,N_7922,N_7998);
or U8011 (N_8011,N_7959,N_7995);
and U8012 (N_8012,N_7936,N_7958);
nand U8013 (N_8013,N_7963,N_7970);
or U8014 (N_8014,N_7968,N_7950);
nand U8015 (N_8015,N_7911,N_7980);
and U8016 (N_8016,N_7944,N_7952);
and U8017 (N_8017,N_7992,N_7908);
and U8018 (N_8018,N_7999,N_7927);
xnor U8019 (N_8019,N_7987,N_7914);
nand U8020 (N_8020,N_7918,N_7967);
or U8021 (N_8021,N_7955,N_7948);
nor U8022 (N_8022,N_7972,N_7930);
or U8023 (N_8023,N_7942,N_7974);
nor U8024 (N_8024,N_7965,N_7984);
and U8025 (N_8025,N_7913,N_7900);
nand U8026 (N_8026,N_7940,N_7909);
and U8027 (N_8027,N_7907,N_7991);
nand U8028 (N_8028,N_7937,N_7905);
xor U8029 (N_8029,N_7935,N_7975);
xor U8030 (N_8030,N_7947,N_7921);
nor U8031 (N_8031,N_7961,N_7983);
nand U8032 (N_8032,N_7933,N_7903);
and U8033 (N_8033,N_7956,N_7990);
and U8034 (N_8034,N_7925,N_7928);
xor U8035 (N_8035,N_7929,N_7949);
and U8036 (N_8036,N_7977,N_7988);
nor U8037 (N_8037,N_7904,N_7931);
nand U8038 (N_8038,N_7915,N_7939);
and U8039 (N_8039,N_7902,N_7941);
or U8040 (N_8040,N_7997,N_7994);
nand U8041 (N_8041,N_7923,N_7946);
and U8042 (N_8042,N_7960,N_7917);
or U8043 (N_8043,N_7910,N_7985);
nor U8044 (N_8044,N_7971,N_7924);
or U8045 (N_8045,N_7973,N_7979);
nor U8046 (N_8046,N_7926,N_7954);
nor U8047 (N_8047,N_7919,N_7953);
and U8048 (N_8048,N_7976,N_7906);
nor U8049 (N_8049,N_7978,N_7957);
nand U8050 (N_8050,N_7902,N_7915);
xnor U8051 (N_8051,N_7922,N_7997);
nand U8052 (N_8052,N_7927,N_7947);
and U8053 (N_8053,N_7965,N_7994);
xnor U8054 (N_8054,N_7912,N_7950);
nand U8055 (N_8055,N_7961,N_7909);
nor U8056 (N_8056,N_7910,N_7911);
or U8057 (N_8057,N_7995,N_7940);
nor U8058 (N_8058,N_7912,N_7907);
nand U8059 (N_8059,N_7905,N_7944);
and U8060 (N_8060,N_7937,N_7966);
or U8061 (N_8061,N_7989,N_7990);
and U8062 (N_8062,N_7929,N_7922);
nor U8063 (N_8063,N_7918,N_7937);
or U8064 (N_8064,N_7988,N_7997);
nand U8065 (N_8065,N_7962,N_7957);
xor U8066 (N_8066,N_7979,N_7948);
or U8067 (N_8067,N_7960,N_7965);
and U8068 (N_8068,N_7942,N_7936);
nor U8069 (N_8069,N_7931,N_7944);
or U8070 (N_8070,N_7965,N_7950);
nor U8071 (N_8071,N_7981,N_7968);
nand U8072 (N_8072,N_7919,N_7994);
nor U8073 (N_8073,N_7930,N_7981);
and U8074 (N_8074,N_7909,N_7960);
or U8075 (N_8075,N_7973,N_7946);
nor U8076 (N_8076,N_7962,N_7978);
nand U8077 (N_8077,N_7944,N_7984);
xor U8078 (N_8078,N_7941,N_7900);
xnor U8079 (N_8079,N_7970,N_7945);
nor U8080 (N_8080,N_7939,N_7934);
or U8081 (N_8081,N_7929,N_7950);
and U8082 (N_8082,N_7925,N_7918);
nand U8083 (N_8083,N_7992,N_7978);
nor U8084 (N_8084,N_7922,N_7938);
and U8085 (N_8085,N_7947,N_7941);
or U8086 (N_8086,N_7941,N_7925);
xnor U8087 (N_8087,N_7972,N_7971);
nand U8088 (N_8088,N_7935,N_7937);
nand U8089 (N_8089,N_7964,N_7965);
xnor U8090 (N_8090,N_7905,N_7947);
nor U8091 (N_8091,N_7987,N_7966);
or U8092 (N_8092,N_7926,N_7962);
xor U8093 (N_8093,N_7964,N_7942);
nor U8094 (N_8094,N_7980,N_7989);
nand U8095 (N_8095,N_7983,N_7943);
and U8096 (N_8096,N_7905,N_7976);
xnor U8097 (N_8097,N_7983,N_7993);
or U8098 (N_8098,N_7998,N_7925);
and U8099 (N_8099,N_7980,N_7936);
or U8100 (N_8100,N_8051,N_8072);
and U8101 (N_8101,N_8083,N_8023);
nor U8102 (N_8102,N_8054,N_8022);
nor U8103 (N_8103,N_8005,N_8025);
nor U8104 (N_8104,N_8027,N_8093);
or U8105 (N_8105,N_8036,N_8089);
nand U8106 (N_8106,N_8053,N_8032);
nor U8107 (N_8107,N_8012,N_8029);
xnor U8108 (N_8108,N_8099,N_8047);
and U8109 (N_8109,N_8007,N_8028);
or U8110 (N_8110,N_8079,N_8008);
nor U8111 (N_8111,N_8086,N_8010);
or U8112 (N_8112,N_8073,N_8002);
xnor U8113 (N_8113,N_8039,N_8038);
nand U8114 (N_8114,N_8065,N_8069);
xor U8115 (N_8115,N_8078,N_8020);
nand U8116 (N_8116,N_8049,N_8055);
and U8117 (N_8117,N_8033,N_8000);
xor U8118 (N_8118,N_8026,N_8096);
nor U8119 (N_8119,N_8016,N_8052);
xnor U8120 (N_8120,N_8043,N_8013);
nand U8121 (N_8121,N_8035,N_8057);
nor U8122 (N_8122,N_8024,N_8067);
nor U8123 (N_8123,N_8044,N_8015);
or U8124 (N_8124,N_8058,N_8003);
and U8125 (N_8125,N_8092,N_8021);
xor U8126 (N_8126,N_8048,N_8070);
and U8127 (N_8127,N_8071,N_8041);
xnor U8128 (N_8128,N_8031,N_8097);
nand U8129 (N_8129,N_8091,N_8088);
xnor U8130 (N_8130,N_8074,N_8077);
xor U8131 (N_8131,N_8040,N_8068);
or U8132 (N_8132,N_8094,N_8090);
or U8133 (N_8133,N_8063,N_8050);
xor U8134 (N_8134,N_8001,N_8014);
nand U8135 (N_8135,N_8059,N_8085);
nor U8136 (N_8136,N_8017,N_8060);
and U8137 (N_8137,N_8006,N_8098);
nor U8138 (N_8138,N_8084,N_8062);
nand U8139 (N_8139,N_8087,N_8075);
nor U8140 (N_8140,N_8064,N_8019);
nor U8141 (N_8141,N_8045,N_8009);
or U8142 (N_8142,N_8042,N_8095);
nor U8143 (N_8143,N_8056,N_8004);
and U8144 (N_8144,N_8030,N_8037);
nand U8145 (N_8145,N_8082,N_8081);
or U8146 (N_8146,N_8046,N_8011);
nor U8147 (N_8147,N_8034,N_8076);
or U8148 (N_8148,N_8061,N_8018);
nand U8149 (N_8149,N_8066,N_8080);
nor U8150 (N_8150,N_8038,N_8079);
or U8151 (N_8151,N_8077,N_8046);
nor U8152 (N_8152,N_8034,N_8082);
xor U8153 (N_8153,N_8029,N_8034);
or U8154 (N_8154,N_8061,N_8029);
nand U8155 (N_8155,N_8049,N_8072);
xor U8156 (N_8156,N_8049,N_8013);
xor U8157 (N_8157,N_8078,N_8029);
and U8158 (N_8158,N_8008,N_8000);
or U8159 (N_8159,N_8060,N_8016);
nand U8160 (N_8160,N_8052,N_8086);
nand U8161 (N_8161,N_8038,N_8008);
nand U8162 (N_8162,N_8070,N_8093);
and U8163 (N_8163,N_8080,N_8044);
nor U8164 (N_8164,N_8039,N_8062);
or U8165 (N_8165,N_8020,N_8030);
and U8166 (N_8166,N_8028,N_8034);
and U8167 (N_8167,N_8029,N_8069);
or U8168 (N_8168,N_8061,N_8034);
and U8169 (N_8169,N_8088,N_8010);
nor U8170 (N_8170,N_8042,N_8098);
and U8171 (N_8171,N_8076,N_8097);
nand U8172 (N_8172,N_8008,N_8087);
or U8173 (N_8173,N_8040,N_8074);
or U8174 (N_8174,N_8065,N_8075);
nor U8175 (N_8175,N_8016,N_8047);
nand U8176 (N_8176,N_8042,N_8063);
or U8177 (N_8177,N_8043,N_8066);
or U8178 (N_8178,N_8094,N_8045);
nand U8179 (N_8179,N_8040,N_8043);
xor U8180 (N_8180,N_8031,N_8064);
or U8181 (N_8181,N_8072,N_8053);
nor U8182 (N_8182,N_8031,N_8033);
nor U8183 (N_8183,N_8082,N_8061);
or U8184 (N_8184,N_8070,N_8064);
nor U8185 (N_8185,N_8051,N_8000);
xor U8186 (N_8186,N_8099,N_8088);
or U8187 (N_8187,N_8057,N_8092);
xor U8188 (N_8188,N_8067,N_8023);
or U8189 (N_8189,N_8008,N_8004);
and U8190 (N_8190,N_8037,N_8023);
and U8191 (N_8191,N_8068,N_8022);
nand U8192 (N_8192,N_8005,N_8091);
and U8193 (N_8193,N_8012,N_8054);
xor U8194 (N_8194,N_8047,N_8044);
and U8195 (N_8195,N_8027,N_8060);
and U8196 (N_8196,N_8062,N_8036);
and U8197 (N_8197,N_8037,N_8060);
or U8198 (N_8198,N_8094,N_8042);
nand U8199 (N_8199,N_8020,N_8037);
nor U8200 (N_8200,N_8177,N_8193);
xor U8201 (N_8201,N_8135,N_8132);
and U8202 (N_8202,N_8195,N_8164);
xnor U8203 (N_8203,N_8185,N_8182);
or U8204 (N_8204,N_8137,N_8129);
xnor U8205 (N_8205,N_8161,N_8108);
nor U8206 (N_8206,N_8163,N_8138);
nor U8207 (N_8207,N_8159,N_8141);
or U8208 (N_8208,N_8117,N_8173);
and U8209 (N_8209,N_8118,N_8111);
or U8210 (N_8210,N_8166,N_8110);
nand U8211 (N_8211,N_8142,N_8187);
or U8212 (N_8212,N_8122,N_8186);
nand U8213 (N_8213,N_8178,N_8162);
xnor U8214 (N_8214,N_8145,N_8107);
nor U8215 (N_8215,N_8174,N_8181);
xnor U8216 (N_8216,N_8123,N_8171);
xnor U8217 (N_8217,N_8146,N_8115);
xnor U8218 (N_8218,N_8152,N_8130);
and U8219 (N_8219,N_8140,N_8197);
or U8220 (N_8220,N_8106,N_8184);
and U8221 (N_8221,N_8167,N_8172);
xor U8222 (N_8222,N_8103,N_8160);
and U8223 (N_8223,N_8155,N_8183);
and U8224 (N_8224,N_8144,N_8104);
nor U8225 (N_8225,N_8196,N_8194);
and U8226 (N_8226,N_8170,N_8168);
nand U8227 (N_8227,N_8114,N_8179);
nand U8228 (N_8228,N_8190,N_8156);
nor U8229 (N_8229,N_8143,N_8149);
or U8230 (N_8230,N_8191,N_8153);
and U8231 (N_8231,N_8151,N_8113);
and U8232 (N_8232,N_8165,N_8112);
or U8233 (N_8233,N_8124,N_8148);
xor U8234 (N_8234,N_8150,N_8175);
and U8235 (N_8235,N_8192,N_8127);
and U8236 (N_8236,N_8136,N_8102);
or U8237 (N_8237,N_8116,N_8157);
or U8238 (N_8238,N_8169,N_8180);
nand U8239 (N_8239,N_8134,N_8126);
or U8240 (N_8240,N_8189,N_8101);
nand U8241 (N_8241,N_8133,N_8128);
or U8242 (N_8242,N_8109,N_8176);
xnor U8243 (N_8243,N_8100,N_8199);
xnor U8244 (N_8244,N_8120,N_8147);
xnor U8245 (N_8245,N_8198,N_8188);
xor U8246 (N_8246,N_8131,N_8154);
nand U8247 (N_8247,N_8121,N_8119);
or U8248 (N_8248,N_8158,N_8105);
nor U8249 (N_8249,N_8125,N_8139);
or U8250 (N_8250,N_8194,N_8110);
and U8251 (N_8251,N_8141,N_8102);
and U8252 (N_8252,N_8156,N_8149);
nand U8253 (N_8253,N_8105,N_8126);
or U8254 (N_8254,N_8175,N_8162);
nand U8255 (N_8255,N_8199,N_8155);
or U8256 (N_8256,N_8166,N_8160);
nor U8257 (N_8257,N_8194,N_8132);
xor U8258 (N_8258,N_8153,N_8166);
and U8259 (N_8259,N_8104,N_8193);
nor U8260 (N_8260,N_8177,N_8109);
xor U8261 (N_8261,N_8157,N_8126);
xnor U8262 (N_8262,N_8146,N_8190);
nand U8263 (N_8263,N_8168,N_8192);
nor U8264 (N_8264,N_8108,N_8186);
nor U8265 (N_8265,N_8125,N_8105);
nor U8266 (N_8266,N_8101,N_8181);
or U8267 (N_8267,N_8162,N_8172);
xor U8268 (N_8268,N_8183,N_8160);
or U8269 (N_8269,N_8164,N_8110);
and U8270 (N_8270,N_8155,N_8167);
nand U8271 (N_8271,N_8131,N_8105);
xnor U8272 (N_8272,N_8189,N_8193);
and U8273 (N_8273,N_8171,N_8195);
and U8274 (N_8274,N_8129,N_8139);
and U8275 (N_8275,N_8105,N_8197);
xnor U8276 (N_8276,N_8168,N_8179);
nand U8277 (N_8277,N_8112,N_8158);
xor U8278 (N_8278,N_8174,N_8179);
or U8279 (N_8279,N_8196,N_8135);
xor U8280 (N_8280,N_8148,N_8197);
xor U8281 (N_8281,N_8110,N_8176);
nor U8282 (N_8282,N_8182,N_8177);
nor U8283 (N_8283,N_8136,N_8121);
xnor U8284 (N_8284,N_8131,N_8176);
and U8285 (N_8285,N_8105,N_8170);
xnor U8286 (N_8286,N_8184,N_8103);
or U8287 (N_8287,N_8195,N_8147);
nor U8288 (N_8288,N_8146,N_8108);
nor U8289 (N_8289,N_8150,N_8159);
xnor U8290 (N_8290,N_8106,N_8177);
nand U8291 (N_8291,N_8126,N_8128);
xor U8292 (N_8292,N_8123,N_8134);
and U8293 (N_8293,N_8190,N_8118);
xor U8294 (N_8294,N_8129,N_8173);
xor U8295 (N_8295,N_8133,N_8137);
xor U8296 (N_8296,N_8174,N_8190);
nor U8297 (N_8297,N_8193,N_8119);
or U8298 (N_8298,N_8143,N_8123);
nand U8299 (N_8299,N_8134,N_8128);
xor U8300 (N_8300,N_8283,N_8295);
and U8301 (N_8301,N_8281,N_8246);
nand U8302 (N_8302,N_8292,N_8220);
or U8303 (N_8303,N_8286,N_8228);
nor U8304 (N_8304,N_8208,N_8231);
nor U8305 (N_8305,N_8278,N_8296);
or U8306 (N_8306,N_8259,N_8212);
xor U8307 (N_8307,N_8289,N_8282);
or U8308 (N_8308,N_8233,N_8235);
and U8309 (N_8309,N_8265,N_8218);
or U8310 (N_8310,N_8294,N_8248);
and U8311 (N_8311,N_8270,N_8239);
nand U8312 (N_8312,N_8277,N_8240);
and U8313 (N_8313,N_8272,N_8209);
and U8314 (N_8314,N_8249,N_8293);
nor U8315 (N_8315,N_8200,N_8285);
and U8316 (N_8316,N_8276,N_8269);
nand U8317 (N_8317,N_8266,N_8238);
or U8318 (N_8318,N_8262,N_8274);
nand U8319 (N_8319,N_8210,N_8229);
or U8320 (N_8320,N_8280,N_8298);
and U8321 (N_8321,N_8232,N_8207);
or U8322 (N_8322,N_8253,N_8299);
and U8323 (N_8323,N_8214,N_8217);
nor U8324 (N_8324,N_8288,N_8211);
and U8325 (N_8325,N_8250,N_8247);
and U8326 (N_8326,N_8219,N_8241);
or U8327 (N_8327,N_8273,N_8201);
nor U8328 (N_8328,N_8215,N_8225);
or U8329 (N_8329,N_8263,N_8290);
and U8330 (N_8330,N_8279,N_8255);
and U8331 (N_8331,N_8254,N_8258);
and U8332 (N_8332,N_8224,N_8216);
and U8333 (N_8333,N_8223,N_8245);
nor U8334 (N_8334,N_8243,N_8261);
nor U8335 (N_8335,N_8244,N_8297);
xnor U8336 (N_8336,N_8237,N_8202);
nor U8337 (N_8337,N_8204,N_8287);
nor U8338 (N_8338,N_8236,N_8234);
nor U8339 (N_8339,N_8203,N_8284);
and U8340 (N_8340,N_8242,N_8251);
or U8341 (N_8341,N_8206,N_8257);
or U8342 (N_8342,N_8264,N_8222);
nand U8343 (N_8343,N_8267,N_8275);
xnor U8344 (N_8344,N_8227,N_8230);
xor U8345 (N_8345,N_8205,N_8213);
or U8346 (N_8346,N_8268,N_8256);
nor U8347 (N_8347,N_8226,N_8221);
nand U8348 (N_8348,N_8291,N_8252);
or U8349 (N_8349,N_8271,N_8260);
or U8350 (N_8350,N_8273,N_8286);
nor U8351 (N_8351,N_8298,N_8241);
nor U8352 (N_8352,N_8200,N_8274);
xnor U8353 (N_8353,N_8270,N_8244);
or U8354 (N_8354,N_8200,N_8278);
nand U8355 (N_8355,N_8221,N_8288);
xor U8356 (N_8356,N_8226,N_8283);
nand U8357 (N_8357,N_8270,N_8263);
nand U8358 (N_8358,N_8284,N_8224);
or U8359 (N_8359,N_8210,N_8294);
nor U8360 (N_8360,N_8230,N_8283);
xor U8361 (N_8361,N_8280,N_8255);
xor U8362 (N_8362,N_8263,N_8207);
nand U8363 (N_8363,N_8261,N_8213);
nand U8364 (N_8364,N_8292,N_8294);
nand U8365 (N_8365,N_8294,N_8284);
or U8366 (N_8366,N_8251,N_8253);
and U8367 (N_8367,N_8284,N_8251);
and U8368 (N_8368,N_8253,N_8242);
nor U8369 (N_8369,N_8279,N_8260);
nor U8370 (N_8370,N_8270,N_8252);
nand U8371 (N_8371,N_8273,N_8229);
nand U8372 (N_8372,N_8239,N_8233);
nor U8373 (N_8373,N_8274,N_8212);
nor U8374 (N_8374,N_8286,N_8284);
nand U8375 (N_8375,N_8288,N_8298);
or U8376 (N_8376,N_8299,N_8284);
xor U8377 (N_8377,N_8280,N_8229);
nor U8378 (N_8378,N_8285,N_8258);
or U8379 (N_8379,N_8267,N_8206);
nor U8380 (N_8380,N_8211,N_8245);
and U8381 (N_8381,N_8238,N_8210);
nor U8382 (N_8382,N_8203,N_8261);
nand U8383 (N_8383,N_8259,N_8239);
or U8384 (N_8384,N_8291,N_8213);
xor U8385 (N_8385,N_8249,N_8261);
and U8386 (N_8386,N_8272,N_8215);
and U8387 (N_8387,N_8236,N_8205);
and U8388 (N_8388,N_8253,N_8289);
xor U8389 (N_8389,N_8214,N_8247);
xnor U8390 (N_8390,N_8297,N_8229);
or U8391 (N_8391,N_8273,N_8270);
nand U8392 (N_8392,N_8246,N_8293);
and U8393 (N_8393,N_8201,N_8271);
nand U8394 (N_8394,N_8200,N_8279);
nor U8395 (N_8395,N_8285,N_8273);
or U8396 (N_8396,N_8256,N_8275);
and U8397 (N_8397,N_8298,N_8269);
xnor U8398 (N_8398,N_8238,N_8226);
nand U8399 (N_8399,N_8225,N_8272);
and U8400 (N_8400,N_8303,N_8373);
nor U8401 (N_8401,N_8360,N_8322);
nor U8402 (N_8402,N_8362,N_8316);
and U8403 (N_8403,N_8306,N_8361);
xor U8404 (N_8404,N_8374,N_8355);
or U8405 (N_8405,N_8378,N_8309);
and U8406 (N_8406,N_8324,N_8387);
xnor U8407 (N_8407,N_8381,N_8386);
nor U8408 (N_8408,N_8375,N_8302);
xnor U8409 (N_8409,N_8395,N_8333);
xnor U8410 (N_8410,N_8337,N_8339);
xnor U8411 (N_8411,N_8383,N_8328);
or U8412 (N_8412,N_8393,N_8349);
nand U8413 (N_8413,N_8326,N_8342);
or U8414 (N_8414,N_8390,N_8335);
xnor U8415 (N_8415,N_8394,N_8338);
nand U8416 (N_8416,N_8385,N_8318);
and U8417 (N_8417,N_8356,N_8369);
and U8418 (N_8418,N_8392,N_8352);
or U8419 (N_8419,N_8305,N_8377);
xnor U8420 (N_8420,N_8331,N_8317);
nand U8421 (N_8421,N_8325,N_8398);
xnor U8422 (N_8422,N_8365,N_8300);
xnor U8423 (N_8423,N_8384,N_8334);
and U8424 (N_8424,N_8379,N_8347);
and U8425 (N_8425,N_8366,N_8319);
nor U8426 (N_8426,N_8327,N_8348);
xor U8427 (N_8427,N_8312,N_8332);
or U8428 (N_8428,N_8344,N_8350);
nand U8429 (N_8429,N_8367,N_8396);
or U8430 (N_8430,N_8376,N_8389);
xnor U8431 (N_8431,N_8359,N_8351);
xnor U8432 (N_8432,N_8358,N_8340);
xor U8433 (N_8433,N_8336,N_8371);
xnor U8434 (N_8434,N_8308,N_8314);
xnor U8435 (N_8435,N_8397,N_8364);
xor U8436 (N_8436,N_8323,N_8320);
xnor U8437 (N_8437,N_8354,N_8341);
nand U8438 (N_8438,N_8343,N_8330);
nor U8439 (N_8439,N_8315,N_8313);
or U8440 (N_8440,N_8372,N_8346);
nand U8441 (N_8441,N_8307,N_8388);
or U8442 (N_8442,N_8380,N_8382);
or U8443 (N_8443,N_8311,N_8321);
nand U8444 (N_8444,N_8391,N_8370);
or U8445 (N_8445,N_8310,N_8363);
xor U8446 (N_8446,N_8329,N_8345);
nor U8447 (N_8447,N_8357,N_8353);
nand U8448 (N_8448,N_8301,N_8399);
or U8449 (N_8449,N_8304,N_8368);
xor U8450 (N_8450,N_8358,N_8367);
and U8451 (N_8451,N_8358,N_8374);
xor U8452 (N_8452,N_8348,N_8339);
and U8453 (N_8453,N_8378,N_8312);
or U8454 (N_8454,N_8348,N_8335);
nand U8455 (N_8455,N_8386,N_8336);
xor U8456 (N_8456,N_8335,N_8325);
nand U8457 (N_8457,N_8372,N_8365);
nor U8458 (N_8458,N_8360,N_8389);
nor U8459 (N_8459,N_8330,N_8397);
nand U8460 (N_8460,N_8340,N_8343);
and U8461 (N_8461,N_8349,N_8303);
nand U8462 (N_8462,N_8322,N_8328);
nand U8463 (N_8463,N_8376,N_8346);
or U8464 (N_8464,N_8319,N_8349);
or U8465 (N_8465,N_8315,N_8364);
or U8466 (N_8466,N_8358,N_8357);
or U8467 (N_8467,N_8308,N_8366);
nor U8468 (N_8468,N_8360,N_8350);
xnor U8469 (N_8469,N_8398,N_8347);
nand U8470 (N_8470,N_8329,N_8375);
nand U8471 (N_8471,N_8364,N_8336);
or U8472 (N_8472,N_8337,N_8356);
and U8473 (N_8473,N_8323,N_8324);
and U8474 (N_8474,N_8314,N_8367);
nand U8475 (N_8475,N_8308,N_8357);
nand U8476 (N_8476,N_8343,N_8325);
xor U8477 (N_8477,N_8393,N_8361);
xor U8478 (N_8478,N_8397,N_8319);
or U8479 (N_8479,N_8383,N_8339);
nor U8480 (N_8480,N_8307,N_8346);
xor U8481 (N_8481,N_8348,N_8389);
or U8482 (N_8482,N_8307,N_8326);
or U8483 (N_8483,N_8347,N_8354);
and U8484 (N_8484,N_8305,N_8363);
xnor U8485 (N_8485,N_8322,N_8354);
or U8486 (N_8486,N_8301,N_8372);
xnor U8487 (N_8487,N_8394,N_8347);
and U8488 (N_8488,N_8334,N_8306);
nor U8489 (N_8489,N_8384,N_8329);
xor U8490 (N_8490,N_8372,N_8395);
nand U8491 (N_8491,N_8310,N_8376);
or U8492 (N_8492,N_8334,N_8366);
or U8493 (N_8493,N_8319,N_8356);
or U8494 (N_8494,N_8392,N_8322);
and U8495 (N_8495,N_8372,N_8347);
and U8496 (N_8496,N_8353,N_8379);
xnor U8497 (N_8497,N_8389,N_8366);
nor U8498 (N_8498,N_8303,N_8374);
nor U8499 (N_8499,N_8317,N_8384);
xor U8500 (N_8500,N_8496,N_8409);
or U8501 (N_8501,N_8460,N_8429);
and U8502 (N_8502,N_8411,N_8441);
nor U8503 (N_8503,N_8483,N_8470);
nand U8504 (N_8504,N_8493,N_8431);
or U8505 (N_8505,N_8400,N_8443);
and U8506 (N_8506,N_8476,N_8471);
nand U8507 (N_8507,N_8419,N_8424);
or U8508 (N_8508,N_8485,N_8402);
xor U8509 (N_8509,N_8427,N_8405);
nand U8510 (N_8510,N_8490,N_8484);
or U8511 (N_8511,N_8401,N_8440);
or U8512 (N_8512,N_8478,N_8477);
nor U8513 (N_8513,N_8486,N_8499);
or U8514 (N_8514,N_8454,N_8455);
nor U8515 (N_8515,N_8472,N_8436);
nor U8516 (N_8516,N_8421,N_8406);
xnor U8517 (N_8517,N_8426,N_8488);
and U8518 (N_8518,N_8491,N_8479);
xor U8519 (N_8519,N_8456,N_8494);
or U8520 (N_8520,N_8432,N_8458);
xnor U8521 (N_8521,N_8464,N_8415);
nor U8522 (N_8522,N_8416,N_8462);
and U8523 (N_8523,N_8497,N_8467);
xor U8524 (N_8524,N_8414,N_8423);
xor U8525 (N_8525,N_8482,N_8412);
xor U8526 (N_8526,N_8438,N_8404);
and U8527 (N_8527,N_8447,N_8466);
or U8528 (N_8528,N_8469,N_8428);
and U8529 (N_8529,N_8468,N_8480);
xnor U8530 (N_8530,N_8474,N_8433);
and U8531 (N_8531,N_8452,N_8457);
xnor U8532 (N_8532,N_8449,N_8413);
and U8533 (N_8533,N_8465,N_8450);
xnor U8534 (N_8534,N_8439,N_8495);
xor U8535 (N_8535,N_8444,N_8492);
nand U8536 (N_8536,N_8437,N_8487);
or U8537 (N_8537,N_8430,N_8403);
nand U8538 (N_8538,N_8489,N_8498);
nand U8539 (N_8539,N_8451,N_8417);
xor U8540 (N_8540,N_8434,N_8418);
and U8541 (N_8541,N_8410,N_8420);
nand U8542 (N_8542,N_8407,N_8408);
or U8543 (N_8543,N_8425,N_8435);
xor U8544 (N_8544,N_8473,N_8481);
nand U8545 (N_8545,N_8448,N_8463);
and U8546 (N_8546,N_8445,N_8461);
and U8547 (N_8547,N_8459,N_8446);
or U8548 (N_8548,N_8475,N_8442);
nand U8549 (N_8549,N_8422,N_8453);
and U8550 (N_8550,N_8424,N_8483);
nor U8551 (N_8551,N_8481,N_8420);
and U8552 (N_8552,N_8435,N_8432);
or U8553 (N_8553,N_8445,N_8417);
nand U8554 (N_8554,N_8414,N_8471);
nand U8555 (N_8555,N_8426,N_8480);
nand U8556 (N_8556,N_8405,N_8439);
nand U8557 (N_8557,N_8416,N_8408);
nor U8558 (N_8558,N_8414,N_8413);
nand U8559 (N_8559,N_8436,N_8469);
nor U8560 (N_8560,N_8463,N_8412);
and U8561 (N_8561,N_8471,N_8446);
or U8562 (N_8562,N_8495,N_8469);
nand U8563 (N_8563,N_8498,N_8471);
or U8564 (N_8564,N_8487,N_8457);
nor U8565 (N_8565,N_8424,N_8451);
or U8566 (N_8566,N_8497,N_8470);
xnor U8567 (N_8567,N_8440,N_8467);
nand U8568 (N_8568,N_8409,N_8487);
nand U8569 (N_8569,N_8422,N_8403);
or U8570 (N_8570,N_8484,N_8447);
nand U8571 (N_8571,N_8447,N_8440);
xnor U8572 (N_8572,N_8425,N_8408);
nor U8573 (N_8573,N_8456,N_8458);
or U8574 (N_8574,N_8490,N_8447);
or U8575 (N_8575,N_8493,N_8433);
or U8576 (N_8576,N_8484,N_8472);
and U8577 (N_8577,N_8449,N_8453);
nor U8578 (N_8578,N_8431,N_8482);
nand U8579 (N_8579,N_8477,N_8472);
and U8580 (N_8580,N_8421,N_8496);
and U8581 (N_8581,N_8448,N_8467);
or U8582 (N_8582,N_8455,N_8492);
nor U8583 (N_8583,N_8494,N_8442);
nor U8584 (N_8584,N_8462,N_8487);
and U8585 (N_8585,N_8486,N_8477);
or U8586 (N_8586,N_8461,N_8407);
or U8587 (N_8587,N_8484,N_8469);
nor U8588 (N_8588,N_8484,N_8429);
nor U8589 (N_8589,N_8452,N_8425);
or U8590 (N_8590,N_8459,N_8441);
nor U8591 (N_8591,N_8497,N_8496);
xor U8592 (N_8592,N_8445,N_8413);
nor U8593 (N_8593,N_8431,N_8468);
and U8594 (N_8594,N_8489,N_8450);
nor U8595 (N_8595,N_8494,N_8484);
nand U8596 (N_8596,N_8450,N_8415);
and U8597 (N_8597,N_8462,N_8449);
and U8598 (N_8598,N_8415,N_8428);
nor U8599 (N_8599,N_8401,N_8459);
nand U8600 (N_8600,N_8533,N_8505);
xor U8601 (N_8601,N_8511,N_8548);
or U8602 (N_8602,N_8549,N_8576);
nor U8603 (N_8603,N_8513,N_8518);
or U8604 (N_8604,N_8598,N_8545);
and U8605 (N_8605,N_8512,N_8582);
or U8606 (N_8606,N_8547,N_8516);
or U8607 (N_8607,N_8532,N_8517);
xor U8608 (N_8608,N_8595,N_8597);
or U8609 (N_8609,N_8501,N_8592);
xor U8610 (N_8610,N_8589,N_8515);
xnor U8611 (N_8611,N_8590,N_8557);
xor U8612 (N_8612,N_8573,N_8571);
or U8613 (N_8613,N_8519,N_8540);
xor U8614 (N_8614,N_8556,N_8504);
and U8615 (N_8615,N_8526,N_8553);
nor U8616 (N_8616,N_8552,N_8534);
xnor U8617 (N_8617,N_8536,N_8500);
or U8618 (N_8618,N_8562,N_8537);
nand U8619 (N_8619,N_8544,N_8528);
or U8620 (N_8620,N_8563,N_8522);
and U8621 (N_8621,N_8567,N_8572);
nand U8622 (N_8622,N_8543,N_8503);
nor U8623 (N_8623,N_8530,N_8535);
xnor U8624 (N_8624,N_8507,N_8575);
and U8625 (N_8625,N_8509,N_8580);
nand U8626 (N_8626,N_8531,N_8588);
nand U8627 (N_8627,N_8554,N_8546);
xnor U8628 (N_8628,N_8524,N_8559);
nor U8629 (N_8629,N_8579,N_8506);
and U8630 (N_8630,N_8570,N_8584);
xor U8631 (N_8631,N_8551,N_8569);
xor U8632 (N_8632,N_8539,N_8583);
or U8633 (N_8633,N_8541,N_8542);
nor U8634 (N_8634,N_8577,N_8578);
and U8635 (N_8635,N_8561,N_8585);
or U8636 (N_8636,N_8596,N_8574);
and U8637 (N_8637,N_8527,N_8565);
or U8638 (N_8638,N_8550,N_8523);
nand U8639 (N_8639,N_8529,N_8525);
or U8640 (N_8640,N_8514,N_8538);
or U8641 (N_8641,N_8510,N_8593);
or U8642 (N_8642,N_8568,N_8599);
nor U8643 (N_8643,N_8581,N_8555);
and U8644 (N_8644,N_8560,N_8566);
nand U8645 (N_8645,N_8564,N_8520);
nor U8646 (N_8646,N_8502,N_8594);
and U8647 (N_8647,N_8508,N_8587);
and U8648 (N_8648,N_8521,N_8591);
nor U8649 (N_8649,N_8586,N_8558);
and U8650 (N_8650,N_8524,N_8567);
and U8651 (N_8651,N_8580,N_8599);
nand U8652 (N_8652,N_8530,N_8538);
nor U8653 (N_8653,N_8568,N_8576);
nor U8654 (N_8654,N_8505,N_8555);
or U8655 (N_8655,N_8555,N_8516);
nand U8656 (N_8656,N_8558,N_8519);
and U8657 (N_8657,N_8579,N_8570);
nand U8658 (N_8658,N_8587,N_8512);
nand U8659 (N_8659,N_8545,N_8554);
nand U8660 (N_8660,N_8558,N_8514);
or U8661 (N_8661,N_8589,N_8537);
and U8662 (N_8662,N_8591,N_8569);
nand U8663 (N_8663,N_8578,N_8579);
xor U8664 (N_8664,N_8551,N_8532);
nor U8665 (N_8665,N_8565,N_8559);
nand U8666 (N_8666,N_8584,N_8505);
or U8667 (N_8667,N_8506,N_8521);
xor U8668 (N_8668,N_8537,N_8587);
xor U8669 (N_8669,N_8569,N_8587);
or U8670 (N_8670,N_8531,N_8560);
xor U8671 (N_8671,N_8569,N_8546);
or U8672 (N_8672,N_8538,N_8552);
and U8673 (N_8673,N_8509,N_8533);
nor U8674 (N_8674,N_8583,N_8572);
nor U8675 (N_8675,N_8519,N_8593);
nor U8676 (N_8676,N_8537,N_8543);
nand U8677 (N_8677,N_8516,N_8571);
nand U8678 (N_8678,N_8599,N_8564);
nand U8679 (N_8679,N_8527,N_8519);
nand U8680 (N_8680,N_8508,N_8547);
nand U8681 (N_8681,N_8522,N_8517);
nand U8682 (N_8682,N_8591,N_8578);
or U8683 (N_8683,N_8567,N_8520);
xnor U8684 (N_8684,N_8579,N_8539);
nor U8685 (N_8685,N_8598,N_8558);
nor U8686 (N_8686,N_8582,N_8598);
and U8687 (N_8687,N_8561,N_8582);
nor U8688 (N_8688,N_8540,N_8584);
xor U8689 (N_8689,N_8545,N_8503);
or U8690 (N_8690,N_8538,N_8500);
xnor U8691 (N_8691,N_8519,N_8504);
nand U8692 (N_8692,N_8571,N_8500);
nand U8693 (N_8693,N_8587,N_8526);
nand U8694 (N_8694,N_8596,N_8508);
nand U8695 (N_8695,N_8502,N_8504);
nand U8696 (N_8696,N_8585,N_8518);
nor U8697 (N_8697,N_8565,N_8524);
nor U8698 (N_8698,N_8538,N_8506);
or U8699 (N_8699,N_8548,N_8598);
nor U8700 (N_8700,N_8632,N_8673);
nand U8701 (N_8701,N_8628,N_8631);
nor U8702 (N_8702,N_8688,N_8624);
nor U8703 (N_8703,N_8671,N_8640);
xor U8704 (N_8704,N_8670,N_8650);
nor U8705 (N_8705,N_8699,N_8695);
nor U8706 (N_8706,N_8644,N_8656);
nor U8707 (N_8707,N_8630,N_8681);
nand U8708 (N_8708,N_8641,N_8619);
xnor U8709 (N_8709,N_8643,N_8639);
nand U8710 (N_8710,N_8667,N_8633);
and U8711 (N_8711,N_8604,N_8677);
and U8712 (N_8712,N_8658,N_8614);
or U8713 (N_8713,N_8648,N_8689);
or U8714 (N_8714,N_8605,N_8646);
and U8715 (N_8715,N_8616,N_8663);
nor U8716 (N_8716,N_8622,N_8607);
nor U8717 (N_8717,N_8625,N_8680);
xor U8718 (N_8718,N_8665,N_8654);
nand U8719 (N_8719,N_8642,N_8606);
and U8720 (N_8720,N_8666,N_8678);
nor U8721 (N_8721,N_8621,N_8601);
nand U8722 (N_8722,N_8683,N_8685);
nor U8723 (N_8723,N_8676,N_8674);
and U8724 (N_8724,N_8668,N_8600);
nor U8725 (N_8725,N_8693,N_8691);
nor U8726 (N_8726,N_8602,N_8651);
or U8727 (N_8727,N_8603,N_8612);
nor U8728 (N_8728,N_8608,N_8655);
nor U8729 (N_8729,N_8687,N_8661);
xnor U8730 (N_8730,N_8627,N_8609);
nor U8731 (N_8731,N_8620,N_8694);
nand U8732 (N_8732,N_8690,N_8617);
or U8733 (N_8733,N_8649,N_8615);
or U8734 (N_8734,N_8634,N_8669);
nand U8735 (N_8735,N_8653,N_8629);
xor U8736 (N_8736,N_8659,N_8647);
and U8737 (N_8737,N_8675,N_8684);
and U8738 (N_8738,N_8618,N_8636);
xor U8739 (N_8739,N_8610,N_8682);
or U8740 (N_8740,N_8686,N_8638);
and U8741 (N_8741,N_8662,N_8613);
nand U8742 (N_8742,N_8626,N_8623);
nor U8743 (N_8743,N_8698,N_8697);
or U8744 (N_8744,N_8664,N_8660);
or U8745 (N_8745,N_8692,N_8657);
nand U8746 (N_8746,N_8696,N_8611);
nor U8747 (N_8747,N_8652,N_8637);
or U8748 (N_8748,N_8635,N_8672);
nor U8749 (N_8749,N_8679,N_8645);
xor U8750 (N_8750,N_8606,N_8664);
or U8751 (N_8751,N_8672,N_8677);
and U8752 (N_8752,N_8666,N_8620);
xnor U8753 (N_8753,N_8635,N_8628);
xor U8754 (N_8754,N_8645,N_8621);
xnor U8755 (N_8755,N_8605,N_8694);
nor U8756 (N_8756,N_8676,N_8603);
or U8757 (N_8757,N_8628,N_8693);
and U8758 (N_8758,N_8658,N_8681);
or U8759 (N_8759,N_8678,N_8697);
or U8760 (N_8760,N_8692,N_8630);
or U8761 (N_8761,N_8639,N_8692);
and U8762 (N_8762,N_8638,N_8609);
and U8763 (N_8763,N_8647,N_8654);
and U8764 (N_8764,N_8629,N_8606);
or U8765 (N_8765,N_8693,N_8639);
and U8766 (N_8766,N_8684,N_8665);
or U8767 (N_8767,N_8605,N_8612);
and U8768 (N_8768,N_8662,N_8628);
nand U8769 (N_8769,N_8677,N_8683);
xor U8770 (N_8770,N_8629,N_8640);
and U8771 (N_8771,N_8669,N_8692);
xnor U8772 (N_8772,N_8615,N_8635);
or U8773 (N_8773,N_8647,N_8605);
and U8774 (N_8774,N_8641,N_8636);
nand U8775 (N_8775,N_8635,N_8668);
nor U8776 (N_8776,N_8674,N_8683);
nor U8777 (N_8777,N_8670,N_8686);
nor U8778 (N_8778,N_8626,N_8643);
nand U8779 (N_8779,N_8617,N_8652);
and U8780 (N_8780,N_8675,N_8655);
and U8781 (N_8781,N_8611,N_8684);
and U8782 (N_8782,N_8653,N_8602);
and U8783 (N_8783,N_8675,N_8672);
nand U8784 (N_8784,N_8614,N_8633);
xnor U8785 (N_8785,N_8681,N_8614);
nor U8786 (N_8786,N_8613,N_8623);
nor U8787 (N_8787,N_8631,N_8668);
xor U8788 (N_8788,N_8637,N_8616);
nand U8789 (N_8789,N_8641,N_8652);
or U8790 (N_8790,N_8651,N_8610);
or U8791 (N_8791,N_8631,N_8643);
or U8792 (N_8792,N_8635,N_8636);
nor U8793 (N_8793,N_8620,N_8647);
nand U8794 (N_8794,N_8667,N_8660);
nor U8795 (N_8795,N_8624,N_8682);
and U8796 (N_8796,N_8669,N_8653);
xnor U8797 (N_8797,N_8673,N_8621);
nor U8798 (N_8798,N_8676,N_8648);
xor U8799 (N_8799,N_8604,N_8694);
xor U8800 (N_8800,N_8799,N_8715);
and U8801 (N_8801,N_8792,N_8753);
nor U8802 (N_8802,N_8709,N_8784);
nand U8803 (N_8803,N_8751,N_8782);
or U8804 (N_8804,N_8789,N_8771);
and U8805 (N_8805,N_8783,N_8764);
nand U8806 (N_8806,N_8756,N_8700);
and U8807 (N_8807,N_8729,N_8749);
xnor U8808 (N_8808,N_8724,N_8763);
or U8809 (N_8809,N_8769,N_8745);
xor U8810 (N_8810,N_8739,N_8710);
nand U8811 (N_8811,N_8713,N_8777);
nand U8812 (N_8812,N_8741,N_8781);
xor U8813 (N_8813,N_8701,N_8740);
and U8814 (N_8814,N_8744,N_8704);
nand U8815 (N_8815,N_8797,N_8737);
nor U8816 (N_8816,N_8727,N_8786);
nand U8817 (N_8817,N_8733,N_8721);
xor U8818 (N_8818,N_8761,N_8774);
nand U8819 (N_8819,N_8747,N_8767);
nor U8820 (N_8820,N_8711,N_8706);
nor U8821 (N_8821,N_8742,N_8796);
xnor U8822 (N_8822,N_8716,N_8798);
nor U8823 (N_8823,N_8773,N_8728);
xor U8824 (N_8824,N_8719,N_8702);
xor U8825 (N_8825,N_8752,N_8772);
nor U8826 (N_8826,N_8757,N_8703);
or U8827 (N_8827,N_8776,N_8730);
xor U8828 (N_8828,N_8768,N_8746);
xnor U8829 (N_8829,N_8743,N_8760);
nor U8830 (N_8830,N_8714,N_8795);
and U8831 (N_8831,N_8791,N_8705);
and U8832 (N_8832,N_8793,N_8720);
xor U8833 (N_8833,N_8750,N_8759);
xnor U8834 (N_8834,N_8788,N_8725);
or U8835 (N_8835,N_8766,N_8770);
xnor U8836 (N_8836,N_8785,N_8707);
or U8837 (N_8837,N_8787,N_8731);
nand U8838 (N_8838,N_8734,N_8762);
nand U8839 (N_8839,N_8708,N_8726);
nand U8840 (N_8840,N_8765,N_8790);
and U8841 (N_8841,N_8794,N_8775);
nand U8842 (N_8842,N_8778,N_8735);
nor U8843 (N_8843,N_8754,N_8736);
nor U8844 (N_8844,N_8758,N_8722);
or U8845 (N_8845,N_8780,N_8718);
nand U8846 (N_8846,N_8748,N_8738);
and U8847 (N_8847,N_8712,N_8779);
or U8848 (N_8848,N_8755,N_8732);
nor U8849 (N_8849,N_8723,N_8717);
nor U8850 (N_8850,N_8724,N_8729);
or U8851 (N_8851,N_8700,N_8721);
and U8852 (N_8852,N_8743,N_8728);
xor U8853 (N_8853,N_8709,N_8717);
or U8854 (N_8854,N_8738,N_8792);
xnor U8855 (N_8855,N_8772,N_8756);
and U8856 (N_8856,N_8773,N_8712);
and U8857 (N_8857,N_8796,N_8722);
or U8858 (N_8858,N_8706,N_8761);
nor U8859 (N_8859,N_8775,N_8771);
and U8860 (N_8860,N_8736,N_8702);
and U8861 (N_8861,N_8747,N_8711);
or U8862 (N_8862,N_8720,N_8727);
and U8863 (N_8863,N_8784,N_8736);
or U8864 (N_8864,N_8772,N_8765);
or U8865 (N_8865,N_8744,N_8711);
and U8866 (N_8866,N_8700,N_8715);
nor U8867 (N_8867,N_8734,N_8772);
nand U8868 (N_8868,N_8724,N_8734);
or U8869 (N_8869,N_8710,N_8784);
or U8870 (N_8870,N_8749,N_8755);
nand U8871 (N_8871,N_8791,N_8798);
nand U8872 (N_8872,N_8762,N_8721);
and U8873 (N_8873,N_8737,N_8745);
and U8874 (N_8874,N_8739,N_8741);
nand U8875 (N_8875,N_8769,N_8760);
or U8876 (N_8876,N_8765,N_8774);
xor U8877 (N_8877,N_8777,N_8750);
and U8878 (N_8878,N_8758,N_8785);
nand U8879 (N_8879,N_8700,N_8795);
and U8880 (N_8880,N_8793,N_8777);
and U8881 (N_8881,N_8703,N_8720);
xnor U8882 (N_8882,N_8724,N_8776);
nand U8883 (N_8883,N_8746,N_8789);
xnor U8884 (N_8884,N_8788,N_8701);
nor U8885 (N_8885,N_8763,N_8741);
or U8886 (N_8886,N_8718,N_8782);
and U8887 (N_8887,N_8707,N_8723);
xor U8888 (N_8888,N_8799,N_8716);
xor U8889 (N_8889,N_8780,N_8799);
nor U8890 (N_8890,N_8717,N_8791);
xor U8891 (N_8891,N_8745,N_8778);
xor U8892 (N_8892,N_8774,N_8781);
or U8893 (N_8893,N_8704,N_8730);
nor U8894 (N_8894,N_8739,N_8738);
xor U8895 (N_8895,N_8780,N_8740);
and U8896 (N_8896,N_8772,N_8744);
xor U8897 (N_8897,N_8724,N_8700);
nor U8898 (N_8898,N_8702,N_8706);
xnor U8899 (N_8899,N_8750,N_8771);
nor U8900 (N_8900,N_8870,N_8806);
and U8901 (N_8901,N_8852,N_8875);
nor U8902 (N_8902,N_8845,N_8889);
and U8903 (N_8903,N_8853,N_8854);
xor U8904 (N_8904,N_8856,N_8872);
nor U8905 (N_8905,N_8801,N_8891);
or U8906 (N_8906,N_8808,N_8871);
xor U8907 (N_8907,N_8867,N_8887);
or U8908 (N_8908,N_8894,N_8868);
and U8909 (N_8909,N_8848,N_8820);
or U8910 (N_8910,N_8814,N_8837);
nor U8911 (N_8911,N_8890,N_8843);
nand U8912 (N_8912,N_8807,N_8859);
and U8913 (N_8913,N_8863,N_8884);
and U8914 (N_8914,N_8850,N_8883);
xnor U8915 (N_8915,N_8827,N_8831);
or U8916 (N_8916,N_8838,N_8885);
nand U8917 (N_8917,N_8834,N_8832);
and U8918 (N_8918,N_8895,N_8858);
or U8919 (N_8919,N_8886,N_8824);
and U8920 (N_8920,N_8802,N_8835);
and U8921 (N_8921,N_8879,N_8860);
nand U8922 (N_8922,N_8805,N_8816);
nor U8923 (N_8923,N_8817,N_8865);
and U8924 (N_8924,N_8829,N_8804);
and U8925 (N_8925,N_8899,N_8819);
and U8926 (N_8926,N_8851,N_8847);
and U8927 (N_8927,N_8822,N_8811);
nor U8928 (N_8928,N_8812,N_8840);
nand U8929 (N_8929,N_8803,N_8892);
or U8930 (N_8930,N_8876,N_8846);
nor U8931 (N_8931,N_8842,N_8833);
nand U8932 (N_8932,N_8825,N_8836);
xnor U8933 (N_8933,N_8830,N_8897);
nand U8934 (N_8934,N_8873,N_8877);
nand U8935 (N_8935,N_8841,N_8888);
nor U8936 (N_8936,N_8881,N_8818);
nor U8937 (N_8937,N_8878,N_8862);
or U8938 (N_8938,N_8882,N_8809);
xnor U8939 (N_8939,N_8857,N_8898);
and U8940 (N_8940,N_8813,N_8823);
xor U8941 (N_8941,N_8810,N_8896);
nand U8942 (N_8942,N_8826,N_8893);
xnor U8943 (N_8943,N_8861,N_8800);
nand U8944 (N_8944,N_8864,N_8849);
and U8945 (N_8945,N_8855,N_8821);
or U8946 (N_8946,N_8874,N_8815);
nor U8947 (N_8947,N_8844,N_8869);
or U8948 (N_8948,N_8839,N_8880);
nand U8949 (N_8949,N_8866,N_8828);
nand U8950 (N_8950,N_8871,N_8873);
xor U8951 (N_8951,N_8828,N_8833);
nand U8952 (N_8952,N_8883,N_8814);
and U8953 (N_8953,N_8860,N_8806);
xnor U8954 (N_8954,N_8849,N_8884);
or U8955 (N_8955,N_8808,N_8847);
nor U8956 (N_8956,N_8851,N_8805);
nor U8957 (N_8957,N_8854,N_8873);
or U8958 (N_8958,N_8824,N_8818);
and U8959 (N_8959,N_8843,N_8879);
or U8960 (N_8960,N_8844,N_8866);
nor U8961 (N_8961,N_8836,N_8818);
nand U8962 (N_8962,N_8840,N_8822);
and U8963 (N_8963,N_8826,N_8836);
xnor U8964 (N_8964,N_8869,N_8810);
nor U8965 (N_8965,N_8823,N_8801);
xnor U8966 (N_8966,N_8870,N_8882);
nand U8967 (N_8967,N_8805,N_8812);
nand U8968 (N_8968,N_8888,N_8831);
nand U8969 (N_8969,N_8840,N_8834);
and U8970 (N_8970,N_8879,N_8868);
nand U8971 (N_8971,N_8890,N_8871);
xnor U8972 (N_8972,N_8855,N_8864);
or U8973 (N_8973,N_8853,N_8846);
xnor U8974 (N_8974,N_8888,N_8879);
and U8975 (N_8975,N_8895,N_8808);
or U8976 (N_8976,N_8883,N_8864);
xor U8977 (N_8977,N_8889,N_8839);
nand U8978 (N_8978,N_8857,N_8843);
and U8979 (N_8979,N_8881,N_8865);
nand U8980 (N_8980,N_8817,N_8829);
nand U8981 (N_8981,N_8823,N_8888);
or U8982 (N_8982,N_8811,N_8834);
or U8983 (N_8983,N_8868,N_8841);
or U8984 (N_8984,N_8802,N_8820);
or U8985 (N_8985,N_8850,N_8859);
and U8986 (N_8986,N_8820,N_8878);
nor U8987 (N_8987,N_8804,N_8854);
or U8988 (N_8988,N_8818,N_8873);
nor U8989 (N_8989,N_8820,N_8847);
or U8990 (N_8990,N_8865,N_8800);
nor U8991 (N_8991,N_8850,N_8838);
nor U8992 (N_8992,N_8819,N_8873);
or U8993 (N_8993,N_8824,N_8889);
nand U8994 (N_8994,N_8880,N_8881);
or U8995 (N_8995,N_8828,N_8868);
nor U8996 (N_8996,N_8807,N_8849);
xor U8997 (N_8997,N_8806,N_8830);
nor U8998 (N_8998,N_8886,N_8859);
and U8999 (N_8999,N_8869,N_8890);
nor U9000 (N_9000,N_8989,N_8966);
or U9001 (N_9001,N_8922,N_8950);
xor U9002 (N_9002,N_8956,N_8945);
or U9003 (N_9003,N_8931,N_8997);
xnor U9004 (N_9004,N_8957,N_8918);
xnor U9005 (N_9005,N_8976,N_8963);
xor U9006 (N_9006,N_8936,N_8967);
and U9007 (N_9007,N_8939,N_8933);
xnor U9008 (N_9008,N_8993,N_8942);
or U9009 (N_9009,N_8973,N_8944);
xor U9010 (N_9010,N_8979,N_8961);
nand U9011 (N_9011,N_8907,N_8971);
xor U9012 (N_9012,N_8964,N_8975);
or U9013 (N_9013,N_8938,N_8968);
and U9014 (N_9014,N_8915,N_8994);
xnor U9015 (N_9015,N_8991,N_8955);
and U9016 (N_9016,N_8949,N_8958);
nand U9017 (N_9017,N_8940,N_8978);
xnor U9018 (N_9018,N_8986,N_8930);
nor U9019 (N_9019,N_8988,N_8959);
nand U9020 (N_9020,N_8926,N_8977);
nand U9021 (N_9021,N_8990,N_8913);
nor U9022 (N_9022,N_8946,N_8952);
or U9023 (N_9023,N_8974,N_8916);
nand U9024 (N_9024,N_8925,N_8904);
xor U9025 (N_9025,N_8983,N_8919);
xor U9026 (N_9026,N_8987,N_8948);
nor U9027 (N_9027,N_8970,N_8982);
xor U9028 (N_9028,N_8984,N_8992);
or U9029 (N_9029,N_8996,N_8902);
or U9030 (N_9030,N_8981,N_8929);
or U9031 (N_9031,N_8917,N_8924);
nor U9032 (N_9032,N_8901,N_8927);
and U9033 (N_9033,N_8911,N_8969);
nor U9034 (N_9034,N_8998,N_8912);
and U9035 (N_9035,N_8921,N_8985);
and U9036 (N_9036,N_8923,N_8999);
xnor U9037 (N_9037,N_8920,N_8965);
xnor U9038 (N_9038,N_8951,N_8937);
and U9039 (N_9039,N_8980,N_8995);
and U9040 (N_9040,N_8908,N_8905);
or U9041 (N_9041,N_8906,N_8954);
nor U9042 (N_9042,N_8900,N_8953);
nand U9043 (N_9043,N_8903,N_8962);
or U9044 (N_9044,N_8943,N_8972);
or U9045 (N_9045,N_8960,N_8935);
or U9046 (N_9046,N_8941,N_8914);
nor U9047 (N_9047,N_8910,N_8928);
nor U9048 (N_9048,N_8909,N_8932);
nand U9049 (N_9049,N_8934,N_8947);
and U9050 (N_9050,N_8977,N_8920);
xor U9051 (N_9051,N_8937,N_8997);
xor U9052 (N_9052,N_8961,N_8963);
nand U9053 (N_9053,N_8961,N_8962);
xnor U9054 (N_9054,N_8979,N_8957);
or U9055 (N_9055,N_8932,N_8991);
or U9056 (N_9056,N_8954,N_8936);
xnor U9057 (N_9057,N_8965,N_8961);
nand U9058 (N_9058,N_8927,N_8961);
and U9059 (N_9059,N_8979,N_8934);
nand U9060 (N_9060,N_8999,N_8983);
nand U9061 (N_9061,N_8954,N_8998);
and U9062 (N_9062,N_8998,N_8961);
nand U9063 (N_9063,N_8925,N_8947);
or U9064 (N_9064,N_8936,N_8964);
nor U9065 (N_9065,N_8997,N_8996);
and U9066 (N_9066,N_8986,N_8946);
xor U9067 (N_9067,N_8940,N_8909);
and U9068 (N_9068,N_8967,N_8919);
xor U9069 (N_9069,N_8953,N_8972);
and U9070 (N_9070,N_8949,N_8959);
or U9071 (N_9071,N_8971,N_8945);
nand U9072 (N_9072,N_8973,N_8935);
nor U9073 (N_9073,N_8983,N_8902);
or U9074 (N_9074,N_8987,N_8961);
nor U9075 (N_9075,N_8934,N_8930);
nor U9076 (N_9076,N_8949,N_8985);
nand U9077 (N_9077,N_8993,N_8952);
nor U9078 (N_9078,N_8993,N_8928);
nand U9079 (N_9079,N_8960,N_8908);
nand U9080 (N_9080,N_8912,N_8916);
or U9081 (N_9081,N_8968,N_8937);
and U9082 (N_9082,N_8914,N_8917);
or U9083 (N_9083,N_8944,N_8946);
nand U9084 (N_9084,N_8921,N_8918);
xor U9085 (N_9085,N_8934,N_8980);
or U9086 (N_9086,N_8972,N_8930);
xnor U9087 (N_9087,N_8984,N_8932);
nand U9088 (N_9088,N_8961,N_8917);
nor U9089 (N_9089,N_8910,N_8940);
xor U9090 (N_9090,N_8991,N_8961);
xnor U9091 (N_9091,N_8953,N_8938);
or U9092 (N_9092,N_8911,N_8928);
and U9093 (N_9093,N_8990,N_8989);
or U9094 (N_9094,N_8986,N_8970);
or U9095 (N_9095,N_8981,N_8912);
and U9096 (N_9096,N_8935,N_8902);
or U9097 (N_9097,N_8972,N_8990);
and U9098 (N_9098,N_8932,N_8907);
and U9099 (N_9099,N_8990,N_8947);
nor U9100 (N_9100,N_9012,N_9067);
and U9101 (N_9101,N_9047,N_9097);
nor U9102 (N_9102,N_9018,N_9044);
nand U9103 (N_9103,N_9016,N_9028);
or U9104 (N_9104,N_9034,N_9073);
and U9105 (N_9105,N_9087,N_9008);
or U9106 (N_9106,N_9070,N_9026);
or U9107 (N_9107,N_9053,N_9086);
nor U9108 (N_9108,N_9099,N_9048);
or U9109 (N_9109,N_9045,N_9088);
xor U9110 (N_9110,N_9036,N_9057);
nor U9111 (N_9111,N_9060,N_9000);
nor U9112 (N_9112,N_9024,N_9051);
nand U9113 (N_9113,N_9011,N_9093);
and U9114 (N_9114,N_9063,N_9031);
nor U9115 (N_9115,N_9043,N_9019);
and U9116 (N_9116,N_9066,N_9085);
and U9117 (N_9117,N_9096,N_9072);
or U9118 (N_9118,N_9091,N_9065);
and U9119 (N_9119,N_9039,N_9081);
or U9120 (N_9120,N_9095,N_9014);
nor U9121 (N_9121,N_9015,N_9089);
and U9122 (N_9122,N_9004,N_9007);
nor U9123 (N_9123,N_9090,N_9033);
and U9124 (N_9124,N_9055,N_9049);
and U9125 (N_9125,N_9013,N_9076);
or U9126 (N_9126,N_9083,N_9074);
nand U9127 (N_9127,N_9038,N_9035);
nor U9128 (N_9128,N_9094,N_9003);
nor U9129 (N_9129,N_9037,N_9069);
or U9130 (N_9130,N_9005,N_9021);
or U9131 (N_9131,N_9042,N_9027);
or U9132 (N_9132,N_9078,N_9062);
xnor U9133 (N_9133,N_9006,N_9002);
or U9134 (N_9134,N_9064,N_9056);
nand U9135 (N_9135,N_9054,N_9098);
and U9136 (N_9136,N_9020,N_9009);
nand U9137 (N_9137,N_9029,N_9052);
and U9138 (N_9138,N_9032,N_9041);
xnor U9139 (N_9139,N_9025,N_9001);
nand U9140 (N_9140,N_9058,N_9023);
and U9141 (N_9141,N_9017,N_9040);
nor U9142 (N_9142,N_9084,N_9075);
xnor U9143 (N_9143,N_9079,N_9030);
and U9144 (N_9144,N_9010,N_9071);
nand U9145 (N_9145,N_9046,N_9050);
or U9146 (N_9146,N_9059,N_9082);
or U9147 (N_9147,N_9068,N_9080);
xor U9148 (N_9148,N_9061,N_9077);
nor U9149 (N_9149,N_9022,N_9092);
nand U9150 (N_9150,N_9093,N_9065);
and U9151 (N_9151,N_9057,N_9061);
nand U9152 (N_9152,N_9083,N_9026);
nor U9153 (N_9153,N_9093,N_9068);
nor U9154 (N_9154,N_9072,N_9070);
xnor U9155 (N_9155,N_9024,N_9001);
xnor U9156 (N_9156,N_9001,N_9046);
nand U9157 (N_9157,N_9031,N_9010);
and U9158 (N_9158,N_9044,N_9050);
xnor U9159 (N_9159,N_9093,N_9072);
and U9160 (N_9160,N_9067,N_9073);
nor U9161 (N_9161,N_9066,N_9077);
nor U9162 (N_9162,N_9044,N_9008);
xnor U9163 (N_9163,N_9032,N_9063);
and U9164 (N_9164,N_9067,N_9062);
xor U9165 (N_9165,N_9022,N_9038);
xor U9166 (N_9166,N_9042,N_9091);
nand U9167 (N_9167,N_9059,N_9012);
xnor U9168 (N_9168,N_9062,N_9014);
xor U9169 (N_9169,N_9047,N_9089);
nor U9170 (N_9170,N_9006,N_9065);
and U9171 (N_9171,N_9036,N_9053);
and U9172 (N_9172,N_9055,N_9056);
xor U9173 (N_9173,N_9070,N_9039);
xnor U9174 (N_9174,N_9077,N_9060);
nor U9175 (N_9175,N_9051,N_9080);
and U9176 (N_9176,N_9050,N_9087);
or U9177 (N_9177,N_9088,N_9071);
and U9178 (N_9178,N_9032,N_9072);
or U9179 (N_9179,N_9061,N_9032);
and U9180 (N_9180,N_9038,N_9058);
and U9181 (N_9181,N_9024,N_9094);
nor U9182 (N_9182,N_9024,N_9030);
or U9183 (N_9183,N_9044,N_9015);
xor U9184 (N_9184,N_9085,N_9048);
and U9185 (N_9185,N_9069,N_9003);
xnor U9186 (N_9186,N_9079,N_9039);
nor U9187 (N_9187,N_9068,N_9085);
nor U9188 (N_9188,N_9009,N_9095);
xnor U9189 (N_9189,N_9013,N_9064);
or U9190 (N_9190,N_9042,N_9040);
xor U9191 (N_9191,N_9091,N_9076);
and U9192 (N_9192,N_9078,N_9001);
xor U9193 (N_9193,N_9012,N_9006);
nor U9194 (N_9194,N_9031,N_9047);
nand U9195 (N_9195,N_9022,N_9059);
nor U9196 (N_9196,N_9053,N_9061);
and U9197 (N_9197,N_9080,N_9090);
or U9198 (N_9198,N_9059,N_9014);
and U9199 (N_9199,N_9078,N_9029);
nor U9200 (N_9200,N_9140,N_9165);
xor U9201 (N_9201,N_9185,N_9127);
xnor U9202 (N_9202,N_9179,N_9199);
nor U9203 (N_9203,N_9131,N_9117);
nor U9204 (N_9204,N_9174,N_9129);
or U9205 (N_9205,N_9189,N_9190);
nor U9206 (N_9206,N_9126,N_9102);
nor U9207 (N_9207,N_9183,N_9146);
and U9208 (N_9208,N_9105,N_9196);
nor U9209 (N_9209,N_9103,N_9144);
nand U9210 (N_9210,N_9121,N_9119);
nand U9211 (N_9211,N_9137,N_9192);
nor U9212 (N_9212,N_9182,N_9187);
xor U9213 (N_9213,N_9170,N_9154);
or U9214 (N_9214,N_9194,N_9191);
nor U9215 (N_9215,N_9157,N_9136);
nor U9216 (N_9216,N_9100,N_9109);
and U9217 (N_9217,N_9116,N_9167);
nor U9218 (N_9218,N_9101,N_9135);
or U9219 (N_9219,N_9139,N_9113);
and U9220 (N_9220,N_9149,N_9143);
or U9221 (N_9221,N_9173,N_9188);
or U9222 (N_9222,N_9176,N_9110);
or U9223 (N_9223,N_9123,N_9147);
nand U9224 (N_9224,N_9156,N_9164);
or U9225 (N_9225,N_9114,N_9178);
and U9226 (N_9226,N_9195,N_9130);
nor U9227 (N_9227,N_9168,N_9160);
or U9228 (N_9228,N_9172,N_9152);
nand U9229 (N_9229,N_9197,N_9166);
or U9230 (N_9230,N_9158,N_9153);
nand U9231 (N_9231,N_9128,N_9120);
xnor U9232 (N_9232,N_9124,N_9159);
and U9233 (N_9233,N_9177,N_9112);
nand U9234 (N_9234,N_9171,N_9132);
nor U9235 (N_9235,N_9162,N_9111);
xnor U9236 (N_9236,N_9138,N_9161);
nor U9237 (N_9237,N_9118,N_9175);
nor U9238 (N_9238,N_9106,N_9169);
or U9239 (N_9239,N_9108,N_9122);
nand U9240 (N_9240,N_9125,N_9193);
xor U9241 (N_9241,N_9133,N_9134);
or U9242 (N_9242,N_9155,N_9145);
xor U9243 (N_9243,N_9141,N_9148);
and U9244 (N_9244,N_9198,N_9181);
or U9245 (N_9245,N_9184,N_9180);
nor U9246 (N_9246,N_9142,N_9107);
or U9247 (N_9247,N_9186,N_9150);
or U9248 (N_9248,N_9104,N_9163);
xor U9249 (N_9249,N_9115,N_9151);
xor U9250 (N_9250,N_9163,N_9191);
nor U9251 (N_9251,N_9183,N_9197);
and U9252 (N_9252,N_9199,N_9178);
nand U9253 (N_9253,N_9162,N_9143);
and U9254 (N_9254,N_9109,N_9146);
nor U9255 (N_9255,N_9185,N_9155);
xor U9256 (N_9256,N_9106,N_9124);
nor U9257 (N_9257,N_9163,N_9169);
or U9258 (N_9258,N_9106,N_9167);
and U9259 (N_9259,N_9125,N_9106);
xor U9260 (N_9260,N_9144,N_9140);
nand U9261 (N_9261,N_9135,N_9107);
or U9262 (N_9262,N_9119,N_9132);
or U9263 (N_9263,N_9126,N_9112);
xnor U9264 (N_9264,N_9111,N_9181);
and U9265 (N_9265,N_9174,N_9197);
nand U9266 (N_9266,N_9116,N_9143);
and U9267 (N_9267,N_9108,N_9135);
nor U9268 (N_9268,N_9185,N_9110);
and U9269 (N_9269,N_9172,N_9162);
nand U9270 (N_9270,N_9176,N_9179);
xnor U9271 (N_9271,N_9136,N_9197);
nor U9272 (N_9272,N_9161,N_9112);
nor U9273 (N_9273,N_9172,N_9174);
or U9274 (N_9274,N_9106,N_9113);
xor U9275 (N_9275,N_9186,N_9164);
or U9276 (N_9276,N_9143,N_9144);
nand U9277 (N_9277,N_9161,N_9126);
nor U9278 (N_9278,N_9106,N_9142);
or U9279 (N_9279,N_9146,N_9129);
nor U9280 (N_9280,N_9178,N_9140);
and U9281 (N_9281,N_9167,N_9151);
nand U9282 (N_9282,N_9150,N_9111);
nor U9283 (N_9283,N_9118,N_9148);
or U9284 (N_9284,N_9157,N_9167);
xnor U9285 (N_9285,N_9135,N_9123);
or U9286 (N_9286,N_9191,N_9120);
or U9287 (N_9287,N_9188,N_9125);
and U9288 (N_9288,N_9162,N_9191);
nand U9289 (N_9289,N_9183,N_9124);
nand U9290 (N_9290,N_9158,N_9197);
and U9291 (N_9291,N_9154,N_9137);
and U9292 (N_9292,N_9165,N_9107);
nand U9293 (N_9293,N_9145,N_9115);
or U9294 (N_9294,N_9158,N_9179);
or U9295 (N_9295,N_9124,N_9135);
or U9296 (N_9296,N_9191,N_9164);
or U9297 (N_9297,N_9175,N_9115);
or U9298 (N_9298,N_9113,N_9199);
nand U9299 (N_9299,N_9153,N_9194);
and U9300 (N_9300,N_9236,N_9211);
or U9301 (N_9301,N_9270,N_9271);
nor U9302 (N_9302,N_9246,N_9275);
nand U9303 (N_9303,N_9255,N_9227);
xor U9304 (N_9304,N_9296,N_9219);
nand U9305 (N_9305,N_9282,N_9245);
or U9306 (N_9306,N_9288,N_9203);
nand U9307 (N_9307,N_9252,N_9265);
or U9308 (N_9308,N_9278,N_9292);
or U9309 (N_9309,N_9268,N_9264);
and U9310 (N_9310,N_9279,N_9286);
xnor U9311 (N_9311,N_9298,N_9244);
nand U9312 (N_9312,N_9206,N_9243);
nand U9313 (N_9313,N_9263,N_9225);
xor U9314 (N_9314,N_9208,N_9238);
and U9315 (N_9315,N_9267,N_9201);
xor U9316 (N_9316,N_9259,N_9251);
xor U9317 (N_9317,N_9248,N_9289);
xor U9318 (N_9318,N_9202,N_9261);
nand U9319 (N_9319,N_9232,N_9253);
nor U9320 (N_9320,N_9204,N_9281);
nand U9321 (N_9321,N_9249,N_9229);
or U9322 (N_9322,N_9299,N_9221);
and U9323 (N_9323,N_9277,N_9220);
xnor U9324 (N_9324,N_9266,N_9224);
nand U9325 (N_9325,N_9250,N_9200);
nor U9326 (N_9326,N_9274,N_9212);
and U9327 (N_9327,N_9280,N_9273);
and U9328 (N_9328,N_9205,N_9242);
or U9329 (N_9329,N_9256,N_9294);
or U9330 (N_9330,N_9269,N_9240);
xnor U9331 (N_9331,N_9231,N_9257);
nor U9332 (N_9332,N_9287,N_9222);
nor U9333 (N_9333,N_9218,N_9254);
nor U9334 (N_9334,N_9235,N_9213);
nor U9335 (N_9335,N_9233,N_9247);
and U9336 (N_9336,N_9285,N_9230);
and U9337 (N_9337,N_9262,N_9283);
and U9338 (N_9338,N_9214,N_9239);
nand U9339 (N_9339,N_9241,N_9217);
nor U9340 (N_9340,N_9215,N_9258);
or U9341 (N_9341,N_9207,N_9228);
nor U9342 (N_9342,N_9237,N_9216);
nor U9343 (N_9343,N_9272,N_9284);
and U9344 (N_9344,N_9293,N_9260);
or U9345 (N_9345,N_9234,N_9297);
xnor U9346 (N_9346,N_9210,N_9295);
or U9347 (N_9347,N_9209,N_9223);
or U9348 (N_9348,N_9276,N_9226);
nor U9349 (N_9349,N_9290,N_9291);
xor U9350 (N_9350,N_9211,N_9283);
nor U9351 (N_9351,N_9205,N_9269);
xor U9352 (N_9352,N_9289,N_9213);
or U9353 (N_9353,N_9260,N_9274);
or U9354 (N_9354,N_9254,N_9219);
nor U9355 (N_9355,N_9289,N_9279);
and U9356 (N_9356,N_9247,N_9290);
nor U9357 (N_9357,N_9297,N_9242);
and U9358 (N_9358,N_9260,N_9214);
or U9359 (N_9359,N_9287,N_9289);
xnor U9360 (N_9360,N_9286,N_9229);
xor U9361 (N_9361,N_9229,N_9214);
xor U9362 (N_9362,N_9209,N_9238);
nand U9363 (N_9363,N_9226,N_9208);
xnor U9364 (N_9364,N_9214,N_9247);
nor U9365 (N_9365,N_9218,N_9286);
nor U9366 (N_9366,N_9270,N_9246);
xor U9367 (N_9367,N_9295,N_9264);
and U9368 (N_9368,N_9268,N_9217);
and U9369 (N_9369,N_9238,N_9239);
xnor U9370 (N_9370,N_9207,N_9235);
nand U9371 (N_9371,N_9259,N_9286);
nor U9372 (N_9372,N_9257,N_9295);
nand U9373 (N_9373,N_9236,N_9287);
and U9374 (N_9374,N_9233,N_9252);
nor U9375 (N_9375,N_9281,N_9226);
xor U9376 (N_9376,N_9283,N_9232);
xor U9377 (N_9377,N_9217,N_9290);
nand U9378 (N_9378,N_9208,N_9265);
or U9379 (N_9379,N_9239,N_9281);
nand U9380 (N_9380,N_9244,N_9214);
xnor U9381 (N_9381,N_9265,N_9238);
nor U9382 (N_9382,N_9220,N_9228);
or U9383 (N_9383,N_9268,N_9246);
xor U9384 (N_9384,N_9285,N_9296);
nand U9385 (N_9385,N_9285,N_9273);
or U9386 (N_9386,N_9217,N_9296);
or U9387 (N_9387,N_9217,N_9286);
nand U9388 (N_9388,N_9215,N_9218);
or U9389 (N_9389,N_9212,N_9279);
or U9390 (N_9390,N_9242,N_9234);
xnor U9391 (N_9391,N_9222,N_9246);
and U9392 (N_9392,N_9242,N_9240);
or U9393 (N_9393,N_9233,N_9244);
or U9394 (N_9394,N_9233,N_9249);
or U9395 (N_9395,N_9266,N_9297);
and U9396 (N_9396,N_9259,N_9210);
xnor U9397 (N_9397,N_9270,N_9223);
and U9398 (N_9398,N_9296,N_9231);
and U9399 (N_9399,N_9207,N_9296);
nor U9400 (N_9400,N_9358,N_9395);
nand U9401 (N_9401,N_9321,N_9386);
and U9402 (N_9402,N_9337,N_9368);
xnor U9403 (N_9403,N_9336,N_9326);
nand U9404 (N_9404,N_9302,N_9312);
nor U9405 (N_9405,N_9399,N_9367);
xor U9406 (N_9406,N_9398,N_9363);
xor U9407 (N_9407,N_9392,N_9330);
nor U9408 (N_9408,N_9301,N_9327);
nor U9409 (N_9409,N_9356,N_9306);
nor U9410 (N_9410,N_9317,N_9360);
nand U9411 (N_9411,N_9366,N_9318);
and U9412 (N_9412,N_9383,N_9307);
nand U9413 (N_9413,N_9365,N_9350);
xnor U9414 (N_9414,N_9319,N_9380);
nor U9415 (N_9415,N_9308,N_9305);
or U9416 (N_9416,N_9344,N_9377);
nor U9417 (N_9417,N_9372,N_9374);
and U9418 (N_9418,N_9373,N_9390);
and U9419 (N_9419,N_9359,N_9388);
and U9420 (N_9420,N_9339,N_9353);
and U9421 (N_9421,N_9340,N_9331);
nor U9422 (N_9422,N_9316,N_9385);
and U9423 (N_9423,N_9393,N_9333);
xor U9424 (N_9424,N_9314,N_9361);
xor U9425 (N_9425,N_9349,N_9397);
and U9426 (N_9426,N_9351,N_9364);
and U9427 (N_9427,N_9389,N_9313);
nand U9428 (N_9428,N_9310,N_9352);
xor U9429 (N_9429,N_9341,N_9370);
xor U9430 (N_9430,N_9348,N_9396);
nand U9431 (N_9431,N_9300,N_9309);
or U9432 (N_9432,N_9322,N_9328);
nand U9433 (N_9433,N_9335,N_9345);
and U9434 (N_9434,N_9346,N_9357);
or U9435 (N_9435,N_9375,N_9343);
nand U9436 (N_9436,N_9342,N_9371);
nor U9437 (N_9437,N_9379,N_9384);
nand U9438 (N_9438,N_9382,N_9315);
xor U9439 (N_9439,N_9362,N_9394);
nand U9440 (N_9440,N_9354,N_9376);
or U9441 (N_9441,N_9369,N_9332);
or U9442 (N_9442,N_9304,N_9355);
nor U9443 (N_9443,N_9347,N_9324);
nand U9444 (N_9444,N_9311,N_9387);
and U9445 (N_9445,N_9338,N_9334);
or U9446 (N_9446,N_9381,N_9303);
and U9447 (N_9447,N_9329,N_9378);
nand U9448 (N_9448,N_9323,N_9320);
xor U9449 (N_9449,N_9391,N_9325);
xor U9450 (N_9450,N_9335,N_9355);
nand U9451 (N_9451,N_9368,N_9386);
or U9452 (N_9452,N_9356,N_9326);
and U9453 (N_9453,N_9324,N_9395);
nor U9454 (N_9454,N_9351,N_9325);
or U9455 (N_9455,N_9384,N_9368);
nand U9456 (N_9456,N_9387,N_9348);
xnor U9457 (N_9457,N_9344,N_9310);
or U9458 (N_9458,N_9387,N_9393);
nand U9459 (N_9459,N_9334,N_9305);
and U9460 (N_9460,N_9389,N_9328);
xor U9461 (N_9461,N_9360,N_9372);
and U9462 (N_9462,N_9340,N_9316);
and U9463 (N_9463,N_9326,N_9386);
nor U9464 (N_9464,N_9349,N_9394);
nor U9465 (N_9465,N_9309,N_9306);
xnor U9466 (N_9466,N_9333,N_9370);
and U9467 (N_9467,N_9372,N_9392);
nand U9468 (N_9468,N_9346,N_9302);
nand U9469 (N_9469,N_9310,N_9380);
nand U9470 (N_9470,N_9384,N_9364);
nand U9471 (N_9471,N_9360,N_9361);
or U9472 (N_9472,N_9309,N_9346);
nand U9473 (N_9473,N_9359,N_9364);
nand U9474 (N_9474,N_9368,N_9398);
or U9475 (N_9475,N_9388,N_9384);
and U9476 (N_9476,N_9340,N_9312);
and U9477 (N_9477,N_9342,N_9318);
or U9478 (N_9478,N_9367,N_9303);
nand U9479 (N_9479,N_9352,N_9365);
nor U9480 (N_9480,N_9388,N_9335);
xor U9481 (N_9481,N_9338,N_9322);
nor U9482 (N_9482,N_9399,N_9352);
xnor U9483 (N_9483,N_9328,N_9376);
nand U9484 (N_9484,N_9313,N_9371);
nor U9485 (N_9485,N_9309,N_9388);
or U9486 (N_9486,N_9352,N_9311);
nand U9487 (N_9487,N_9349,N_9332);
nor U9488 (N_9488,N_9351,N_9344);
and U9489 (N_9489,N_9368,N_9321);
nor U9490 (N_9490,N_9386,N_9357);
or U9491 (N_9491,N_9343,N_9383);
and U9492 (N_9492,N_9397,N_9312);
nor U9493 (N_9493,N_9368,N_9392);
nor U9494 (N_9494,N_9358,N_9374);
xor U9495 (N_9495,N_9340,N_9321);
or U9496 (N_9496,N_9386,N_9397);
xor U9497 (N_9497,N_9371,N_9366);
nor U9498 (N_9498,N_9362,N_9357);
and U9499 (N_9499,N_9368,N_9311);
and U9500 (N_9500,N_9426,N_9446);
or U9501 (N_9501,N_9490,N_9419);
nand U9502 (N_9502,N_9448,N_9413);
nor U9503 (N_9503,N_9484,N_9441);
and U9504 (N_9504,N_9486,N_9435);
nor U9505 (N_9505,N_9407,N_9422);
or U9506 (N_9506,N_9497,N_9440);
or U9507 (N_9507,N_9453,N_9491);
and U9508 (N_9508,N_9437,N_9408);
and U9509 (N_9509,N_9481,N_9474);
and U9510 (N_9510,N_9496,N_9452);
nand U9511 (N_9511,N_9409,N_9480);
xnor U9512 (N_9512,N_9431,N_9468);
nor U9513 (N_9513,N_9457,N_9429);
nand U9514 (N_9514,N_9401,N_9466);
or U9515 (N_9515,N_9430,N_9428);
nor U9516 (N_9516,N_9462,N_9421);
or U9517 (N_9517,N_9488,N_9471);
or U9518 (N_9518,N_9454,N_9434);
nand U9519 (N_9519,N_9447,N_9479);
nor U9520 (N_9520,N_9499,N_9494);
or U9521 (N_9521,N_9414,N_9476);
and U9522 (N_9522,N_9423,N_9492);
xor U9523 (N_9523,N_9439,N_9498);
or U9524 (N_9524,N_9469,N_9472);
and U9525 (N_9525,N_9443,N_9473);
nand U9526 (N_9526,N_9402,N_9482);
or U9527 (N_9527,N_9417,N_9455);
nand U9528 (N_9528,N_9442,N_9424);
or U9529 (N_9529,N_9493,N_9467);
xnor U9530 (N_9530,N_9451,N_9412);
xor U9531 (N_9531,N_9475,N_9425);
or U9532 (N_9532,N_9495,N_9400);
nand U9533 (N_9533,N_9411,N_9410);
xor U9534 (N_9534,N_9483,N_9478);
nor U9535 (N_9535,N_9458,N_9485);
nor U9536 (N_9536,N_9450,N_9436);
nor U9537 (N_9537,N_9449,N_9445);
xnor U9538 (N_9538,N_9432,N_9433);
nand U9539 (N_9539,N_9456,N_9420);
or U9540 (N_9540,N_9444,N_9438);
nor U9541 (N_9541,N_9405,N_9463);
or U9542 (N_9542,N_9470,N_9416);
and U9543 (N_9543,N_9465,N_9461);
xnor U9544 (N_9544,N_9415,N_9464);
and U9545 (N_9545,N_9403,N_9459);
nor U9546 (N_9546,N_9404,N_9487);
or U9547 (N_9547,N_9427,N_9489);
and U9548 (N_9548,N_9406,N_9477);
nor U9549 (N_9549,N_9460,N_9418);
nor U9550 (N_9550,N_9410,N_9440);
xnor U9551 (N_9551,N_9412,N_9455);
xor U9552 (N_9552,N_9434,N_9421);
or U9553 (N_9553,N_9435,N_9420);
xnor U9554 (N_9554,N_9427,N_9418);
nand U9555 (N_9555,N_9405,N_9454);
xnor U9556 (N_9556,N_9442,N_9444);
nand U9557 (N_9557,N_9450,N_9469);
nand U9558 (N_9558,N_9483,N_9485);
xnor U9559 (N_9559,N_9437,N_9407);
and U9560 (N_9560,N_9443,N_9467);
nor U9561 (N_9561,N_9457,N_9497);
and U9562 (N_9562,N_9460,N_9426);
nand U9563 (N_9563,N_9464,N_9457);
xor U9564 (N_9564,N_9465,N_9452);
or U9565 (N_9565,N_9409,N_9436);
xor U9566 (N_9566,N_9422,N_9427);
nand U9567 (N_9567,N_9485,N_9461);
nand U9568 (N_9568,N_9428,N_9435);
and U9569 (N_9569,N_9482,N_9498);
or U9570 (N_9570,N_9444,N_9452);
or U9571 (N_9571,N_9432,N_9462);
xnor U9572 (N_9572,N_9404,N_9457);
or U9573 (N_9573,N_9467,N_9430);
and U9574 (N_9574,N_9435,N_9409);
and U9575 (N_9575,N_9477,N_9464);
nor U9576 (N_9576,N_9416,N_9445);
and U9577 (N_9577,N_9476,N_9462);
nor U9578 (N_9578,N_9431,N_9406);
or U9579 (N_9579,N_9404,N_9455);
and U9580 (N_9580,N_9427,N_9444);
xnor U9581 (N_9581,N_9471,N_9447);
or U9582 (N_9582,N_9490,N_9485);
nor U9583 (N_9583,N_9460,N_9414);
nand U9584 (N_9584,N_9400,N_9468);
nor U9585 (N_9585,N_9491,N_9402);
or U9586 (N_9586,N_9459,N_9420);
or U9587 (N_9587,N_9490,N_9492);
nand U9588 (N_9588,N_9467,N_9401);
and U9589 (N_9589,N_9464,N_9459);
nor U9590 (N_9590,N_9449,N_9418);
or U9591 (N_9591,N_9421,N_9482);
nand U9592 (N_9592,N_9443,N_9422);
and U9593 (N_9593,N_9446,N_9465);
nand U9594 (N_9594,N_9468,N_9490);
nor U9595 (N_9595,N_9436,N_9413);
and U9596 (N_9596,N_9436,N_9404);
nand U9597 (N_9597,N_9410,N_9469);
nor U9598 (N_9598,N_9431,N_9497);
or U9599 (N_9599,N_9411,N_9449);
and U9600 (N_9600,N_9544,N_9551);
xor U9601 (N_9601,N_9597,N_9598);
or U9602 (N_9602,N_9515,N_9521);
xnor U9603 (N_9603,N_9582,N_9554);
and U9604 (N_9604,N_9596,N_9584);
or U9605 (N_9605,N_9532,N_9502);
nand U9606 (N_9606,N_9507,N_9510);
nor U9607 (N_9607,N_9514,N_9567);
xor U9608 (N_9608,N_9526,N_9503);
and U9609 (N_9609,N_9574,N_9566);
xor U9610 (N_9610,N_9555,N_9550);
nand U9611 (N_9611,N_9535,N_9558);
nor U9612 (N_9612,N_9505,N_9516);
and U9613 (N_9613,N_9571,N_9540);
or U9614 (N_9614,N_9501,N_9511);
or U9615 (N_9615,N_9534,N_9541);
and U9616 (N_9616,N_9563,N_9577);
nand U9617 (N_9617,N_9561,N_9583);
xor U9618 (N_9618,N_9560,N_9565);
xnor U9619 (N_9619,N_9517,N_9576);
nand U9620 (N_9620,N_9508,N_9549);
or U9621 (N_9621,N_9529,N_9509);
nor U9622 (N_9622,N_9586,N_9581);
and U9623 (N_9623,N_9556,N_9530);
xnor U9624 (N_9624,N_9547,N_9537);
nand U9625 (N_9625,N_9538,N_9506);
and U9626 (N_9626,N_9585,N_9542);
xnor U9627 (N_9627,N_9504,N_9545);
nor U9628 (N_9628,N_9559,N_9579);
or U9629 (N_9629,N_9575,N_9564);
nand U9630 (N_9630,N_9500,N_9536);
nor U9631 (N_9631,N_9589,N_9593);
nand U9632 (N_9632,N_9569,N_9523);
or U9633 (N_9633,N_9522,N_9548);
nand U9634 (N_9634,N_9513,N_9525);
or U9635 (N_9635,N_9520,N_9546);
or U9636 (N_9636,N_9553,N_9518);
or U9637 (N_9637,N_9562,N_9573);
nand U9638 (N_9638,N_9592,N_9572);
or U9639 (N_9639,N_9568,N_9531);
or U9640 (N_9640,N_9590,N_9588);
or U9641 (N_9641,N_9528,N_9543);
and U9642 (N_9642,N_9552,N_9587);
xnor U9643 (N_9643,N_9578,N_9539);
and U9644 (N_9644,N_9557,N_9524);
nand U9645 (N_9645,N_9591,N_9570);
nand U9646 (N_9646,N_9512,N_9599);
xor U9647 (N_9647,N_9533,N_9519);
or U9648 (N_9648,N_9527,N_9580);
xnor U9649 (N_9649,N_9595,N_9594);
and U9650 (N_9650,N_9597,N_9595);
or U9651 (N_9651,N_9523,N_9545);
and U9652 (N_9652,N_9594,N_9596);
and U9653 (N_9653,N_9567,N_9518);
and U9654 (N_9654,N_9569,N_9561);
or U9655 (N_9655,N_9547,N_9541);
or U9656 (N_9656,N_9552,N_9515);
nor U9657 (N_9657,N_9545,N_9557);
nand U9658 (N_9658,N_9524,N_9522);
and U9659 (N_9659,N_9544,N_9558);
xor U9660 (N_9660,N_9536,N_9558);
or U9661 (N_9661,N_9525,N_9501);
and U9662 (N_9662,N_9524,N_9531);
or U9663 (N_9663,N_9543,N_9530);
nor U9664 (N_9664,N_9556,N_9571);
or U9665 (N_9665,N_9559,N_9541);
or U9666 (N_9666,N_9590,N_9557);
or U9667 (N_9667,N_9578,N_9531);
or U9668 (N_9668,N_9500,N_9539);
nor U9669 (N_9669,N_9596,N_9550);
nor U9670 (N_9670,N_9582,N_9541);
xnor U9671 (N_9671,N_9506,N_9555);
nor U9672 (N_9672,N_9591,N_9550);
nor U9673 (N_9673,N_9556,N_9539);
nor U9674 (N_9674,N_9583,N_9542);
nand U9675 (N_9675,N_9548,N_9530);
nor U9676 (N_9676,N_9501,N_9571);
and U9677 (N_9677,N_9512,N_9560);
or U9678 (N_9678,N_9596,N_9535);
nand U9679 (N_9679,N_9506,N_9545);
and U9680 (N_9680,N_9520,N_9594);
or U9681 (N_9681,N_9502,N_9563);
nand U9682 (N_9682,N_9547,N_9550);
and U9683 (N_9683,N_9549,N_9588);
and U9684 (N_9684,N_9521,N_9503);
or U9685 (N_9685,N_9583,N_9563);
nor U9686 (N_9686,N_9588,N_9572);
nand U9687 (N_9687,N_9568,N_9517);
or U9688 (N_9688,N_9596,N_9583);
nand U9689 (N_9689,N_9502,N_9587);
nand U9690 (N_9690,N_9513,N_9546);
and U9691 (N_9691,N_9585,N_9520);
nand U9692 (N_9692,N_9557,N_9538);
nand U9693 (N_9693,N_9583,N_9550);
nor U9694 (N_9694,N_9590,N_9558);
or U9695 (N_9695,N_9597,N_9599);
nor U9696 (N_9696,N_9530,N_9593);
nor U9697 (N_9697,N_9507,N_9597);
nand U9698 (N_9698,N_9569,N_9596);
nand U9699 (N_9699,N_9549,N_9536);
or U9700 (N_9700,N_9689,N_9663);
nand U9701 (N_9701,N_9651,N_9629);
nor U9702 (N_9702,N_9615,N_9636);
and U9703 (N_9703,N_9611,N_9683);
nor U9704 (N_9704,N_9682,N_9687);
or U9705 (N_9705,N_9698,N_9603);
nand U9706 (N_9706,N_9628,N_9622);
or U9707 (N_9707,N_9623,N_9601);
and U9708 (N_9708,N_9618,N_9690);
xor U9709 (N_9709,N_9645,N_9613);
or U9710 (N_9710,N_9681,N_9608);
and U9711 (N_9711,N_9648,N_9652);
or U9712 (N_9712,N_9624,N_9695);
nand U9713 (N_9713,N_9678,N_9659);
nand U9714 (N_9714,N_9602,N_9642);
and U9715 (N_9715,N_9685,N_9697);
or U9716 (N_9716,N_9649,N_9639);
nand U9717 (N_9717,N_9604,N_9664);
or U9718 (N_9718,N_9609,N_9699);
nand U9719 (N_9719,N_9661,N_9653);
nor U9720 (N_9720,N_9675,N_9633);
xnor U9721 (N_9721,N_9671,N_9632);
xnor U9722 (N_9722,N_9650,N_9638);
or U9723 (N_9723,N_9617,N_9676);
xnor U9724 (N_9724,N_9605,N_9672);
nand U9725 (N_9725,N_9677,N_9626);
and U9726 (N_9726,N_9647,N_9686);
xnor U9727 (N_9727,N_9688,N_9665);
nor U9728 (N_9728,N_9641,N_9684);
or U9729 (N_9729,N_9693,N_9666);
or U9730 (N_9730,N_9621,N_9692);
or U9731 (N_9731,N_9627,N_9620);
xnor U9732 (N_9732,N_9614,N_9600);
or U9733 (N_9733,N_9631,N_9646);
xor U9734 (N_9734,N_9696,N_9654);
or U9735 (N_9735,N_9606,N_9643);
xor U9736 (N_9736,N_9607,N_9612);
or U9737 (N_9737,N_9610,N_9673);
nand U9738 (N_9738,N_9644,N_9660);
xnor U9739 (N_9739,N_9619,N_9625);
and U9740 (N_9740,N_9634,N_9616);
or U9741 (N_9741,N_9655,N_9662);
xnor U9742 (N_9742,N_9657,N_9670);
or U9743 (N_9743,N_9679,N_9630);
nor U9744 (N_9744,N_9680,N_9656);
xor U9745 (N_9745,N_9667,N_9635);
xor U9746 (N_9746,N_9669,N_9691);
nand U9747 (N_9747,N_9668,N_9694);
nor U9748 (N_9748,N_9658,N_9674);
xor U9749 (N_9749,N_9637,N_9640);
xnor U9750 (N_9750,N_9690,N_9631);
nor U9751 (N_9751,N_9698,N_9694);
or U9752 (N_9752,N_9681,N_9651);
or U9753 (N_9753,N_9657,N_9611);
nor U9754 (N_9754,N_9674,N_9690);
xor U9755 (N_9755,N_9622,N_9666);
nand U9756 (N_9756,N_9686,N_9617);
nand U9757 (N_9757,N_9614,N_9682);
nor U9758 (N_9758,N_9669,N_9639);
or U9759 (N_9759,N_9625,N_9667);
xnor U9760 (N_9760,N_9679,N_9686);
nor U9761 (N_9761,N_9671,N_9637);
nor U9762 (N_9762,N_9675,N_9696);
xnor U9763 (N_9763,N_9611,N_9686);
nor U9764 (N_9764,N_9639,N_9638);
or U9765 (N_9765,N_9615,N_9670);
xor U9766 (N_9766,N_9682,N_9610);
and U9767 (N_9767,N_9616,N_9694);
xor U9768 (N_9768,N_9659,N_9693);
nand U9769 (N_9769,N_9661,N_9643);
nor U9770 (N_9770,N_9675,N_9637);
xnor U9771 (N_9771,N_9687,N_9606);
nand U9772 (N_9772,N_9644,N_9606);
nor U9773 (N_9773,N_9601,N_9682);
nand U9774 (N_9774,N_9647,N_9666);
nor U9775 (N_9775,N_9668,N_9657);
nand U9776 (N_9776,N_9699,N_9630);
or U9777 (N_9777,N_9685,N_9655);
nor U9778 (N_9778,N_9661,N_9642);
nand U9779 (N_9779,N_9635,N_9658);
nor U9780 (N_9780,N_9602,N_9629);
nand U9781 (N_9781,N_9665,N_9627);
or U9782 (N_9782,N_9687,N_9680);
nand U9783 (N_9783,N_9695,N_9620);
or U9784 (N_9784,N_9616,N_9630);
nand U9785 (N_9785,N_9693,N_9694);
xnor U9786 (N_9786,N_9600,N_9678);
xnor U9787 (N_9787,N_9692,N_9607);
or U9788 (N_9788,N_9603,N_9677);
nor U9789 (N_9789,N_9663,N_9615);
xor U9790 (N_9790,N_9636,N_9633);
nand U9791 (N_9791,N_9672,N_9680);
xnor U9792 (N_9792,N_9666,N_9673);
xnor U9793 (N_9793,N_9630,N_9632);
nor U9794 (N_9794,N_9614,N_9675);
xor U9795 (N_9795,N_9690,N_9641);
nand U9796 (N_9796,N_9677,N_9649);
xor U9797 (N_9797,N_9616,N_9695);
nand U9798 (N_9798,N_9637,N_9691);
nor U9799 (N_9799,N_9611,N_9609);
nor U9800 (N_9800,N_9766,N_9733);
nor U9801 (N_9801,N_9707,N_9782);
xor U9802 (N_9802,N_9780,N_9792);
nand U9803 (N_9803,N_9778,N_9789);
nand U9804 (N_9804,N_9755,N_9713);
nand U9805 (N_9805,N_9781,N_9734);
nand U9806 (N_9806,N_9729,N_9718);
nand U9807 (N_9807,N_9701,N_9720);
or U9808 (N_9808,N_9764,N_9706);
and U9809 (N_9809,N_9716,N_9738);
nor U9810 (N_9810,N_9711,N_9749);
or U9811 (N_9811,N_9793,N_9726);
nor U9812 (N_9812,N_9772,N_9747);
xor U9813 (N_9813,N_9771,N_9743);
and U9814 (N_9814,N_9784,N_9730);
or U9815 (N_9815,N_9760,N_9753);
nor U9816 (N_9816,N_9737,N_9731);
xnor U9817 (N_9817,N_9769,N_9761);
xnor U9818 (N_9818,N_9714,N_9758);
or U9819 (N_9819,N_9775,N_9739);
xor U9820 (N_9820,N_9790,N_9709);
or U9821 (N_9821,N_9774,N_9708);
or U9822 (N_9822,N_9705,N_9791);
xor U9823 (N_9823,N_9723,N_9777);
xor U9824 (N_9824,N_9759,N_9797);
xor U9825 (N_9825,N_9712,N_9768);
nand U9826 (N_9826,N_9745,N_9779);
or U9827 (N_9827,N_9719,N_9736);
xnor U9828 (N_9828,N_9783,N_9702);
nor U9829 (N_9829,N_9752,N_9762);
xnor U9830 (N_9830,N_9754,N_9748);
xnor U9831 (N_9831,N_9796,N_9735);
nand U9832 (N_9832,N_9785,N_9741);
nand U9833 (N_9833,N_9717,N_9710);
nor U9834 (N_9834,N_9776,N_9724);
and U9835 (N_9835,N_9799,N_9765);
and U9836 (N_9836,N_9722,N_9732);
nand U9837 (N_9837,N_9725,N_9757);
xor U9838 (N_9838,N_9795,N_9787);
and U9839 (N_9839,N_9721,N_9740);
nor U9840 (N_9840,N_9744,N_9746);
or U9841 (N_9841,N_9742,N_9794);
nand U9842 (N_9842,N_9727,N_9700);
and U9843 (N_9843,N_9750,N_9715);
nand U9844 (N_9844,N_9788,N_9786);
nand U9845 (N_9845,N_9751,N_9763);
nand U9846 (N_9846,N_9770,N_9728);
nand U9847 (N_9847,N_9767,N_9703);
or U9848 (N_9848,N_9704,N_9773);
nor U9849 (N_9849,N_9756,N_9798);
or U9850 (N_9850,N_9742,N_9775);
and U9851 (N_9851,N_9723,N_9730);
xor U9852 (N_9852,N_9706,N_9709);
and U9853 (N_9853,N_9754,N_9711);
and U9854 (N_9854,N_9765,N_9736);
nand U9855 (N_9855,N_9703,N_9718);
and U9856 (N_9856,N_9756,N_9788);
or U9857 (N_9857,N_9734,N_9709);
nor U9858 (N_9858,N_9716,N_9744);
xnor U9859 (N_9859,N_9738,N_9743);
xor U9860 (N_9860,N_9731,N_9715);
or U9861 (N_9861,N_9731,N_9716);
and U9862 (N_9862,N_9725,N_9778);
xor U9863 (N_9863,N_9719,N_9794);
xnor U9864 (N_9864,N_9706,N_9746);
xnor U9865 (N_9865,N_9792,N_9775);
and U9866 (N_9866,N_9745,N_9728);
or U9867 (N_9867,N_9774,N_9775);
or U9868 (N_9868,N_9704,N_9703);
nand U9869 (N_9869,N_9725,N_9775);
nand U9870 (N_9870,N_9707,N_9745);
or U9871 (N_9871,N_9724,N_9701);
xnor U9872 (N_9872,N_9795,N_9725);
and U9873 (N_9873,N_9773,N_9710);
nand U9874 (N_9874,N_9723,N_9713);
xnor U9875 (N_9875,N_9787,N_9703);
nor U9876 (N_9876,N_9788,N_9770);
and U9877 (N_9877,N_9791,N_9709);
nand U9878 (N_9878,N_9713,N_9745);
nand U9879 (N_9879,N_9719,N_9781);
or U9880 (N_9880,N_9793,N_9766);
nand U9881 (N_9881,N_9781,N_9750);
xnor U9882 (N_9882,N_9714,N_9712);
nand U9883 (N_9883,N_9749,N_9738);
nand U9884 (N_9884,N_9728,N_9739);
and U9885 (N_9885,N_9711,N_9797);
nand U9886 (N_9886,N_9730,N_9710);
nand U9887 (N_9887,N_9788,N_9706);
xnor U9888 (N_9888,N_9739,N_9752);
nand U9889 (N_9889,N_9770,N_9723);
nand U9890 (N_9890,N_9719,N_9757);
nand U9891 (N_9891,N_9747,N_9752);
or U9892 (N_9892,N_9733,N_9778);
nand U9893 (N_9893,N_9771,N_9706);
and U9894 (N_9894,N_9743,N_9781);
and U9895 (N_9895,N_9781,N_9772);
or U9896 (N_9896,N_9719,N_9747);
and U9897 (N_9897,N_9752,N_9757);
xnor U9898 (N_9898,N_9752,N_9701);
or U9899 (N_9899,N_9742,N_9784);
xor U9900 (N_9900,N_9838,N_9844);
and U9901 (N_9901,N_9807,N_9812);
xnor U9902 (N_9902,N_9818,N_9836);
xor U9903 (N_9903,N_9864,N_9881);
nor U9904 (N_9904,N_9852,N_9847);
nor U9905 (N_9905,N_9822,N_9872);
xor U9906 (N_9906,N_9845,N_9829);
nor U9907 (N_9907,N_9825,N_9816);
or U9908 (N_9908,N_9899,N_9811);
nand U9909 (N_9909,N_9806,N_9809);
and U9910 (N_9910,N_9866,N_9857);
nor U9911 (N_9911,N_9892,N_9887);
and U9912 (N_9912,N_9804,N_9833);
xnor U9913 (N_9913,N_9898,N_9851);
nor U9914 (N_9914,N_9875,N_9839);
nor U9915 (N_9915,N_9870,N_9873);
nand U9916 (N_9916,N_9874,N_9858);
or U9917 (N_9917,N_9882,N_9835);
xnor U9918 (N_9918,N_9869,N_9859);
or U9919 (N_9919,N_9850,N_9867);
nand U9920 (N_9920,N_9800,N_9805);
or U9921 (N_9921,N_9840,N_9827);
nor U9922 (N_9922,N_9877,N_9841);
or U9923 (N_9923,N_9830,N_9897);
or U9924 (N_9924,N_9876,N_9890);
xnor U9925 (N_9925,N_9863,N_9878);
nor U9926 (N_9926,N_9837,N_9884);
or U9927 (N_9927,N_9823,N_9808);
nor U9928 (N_9928,N_9801,N_9848);
and U9929 (N_9929,N_9853,N_9893);
nor U9930 (N_9930,N_9846,N_9813);
nor U9931 (N_9931,N_9826,N_9842);
nor U9932 (N_9932,N_9860,N_9802);
or U9933 (N_9933,N_9849,N_9828);
nand U9934 (N_9934,N_9819,N_9894);
xnor U9935 (N_9935,N_9824,N_9817);
nand U9936 (N_9936,N_9843,N_9831);
and U9937 (N_9937,N_9856,N_9865);
nor U9938 (N_9938,N_9810,N_9891);
nand U9939 (N_9939,N_9820,N_9886);
or U9940 (N_9940,N_9871,N_9861);
nor U9941 (N_9941,N_9896,N_9868);
and U9942 (N_9942,N_9885,N_9832);
nor U9943 (N_9943,N_9888,N_9855);
xnor U9944 (N_9944,N_9803,N_9895);
nand U9945 (N_9945,N_9814,N_9879);
nor U9946 (N_9946,N_9821,N_9815);
and U9947 (N_9947,N_9880,N_9889);
and U9948 (N_9948,N_9883,N_9862);
xor U9949 (N_9949,N_9854,N_9834);
and U9950 (N_9950,N_9808,N_9878);
and U9951 (N_9951,N_9803,N_9824);
or U9952 (N_9952,N_9889,N_9833);
nor U9953 (N_9953,N_9898,N_9825);
nor U9954 (N_9954,N_9858,N_9890);
xor U9955 (N_9955,N_9877,N_9866);
nand U9956 (N_9956,N_9818,N_9853);
xnor U9957 (N_9957,N_9858,N_9875);
nor U9958 (N_9958,N_9803,N_9887);
nor U9959 (N_9959,N_9883,N_9885);
and U9960 (N_9960,N_9860,N_9888);
and U9961 (N_9961,N_9882,N_9817);
or U9962 (N_9962,N_9843,N_9813);
and U9963 (N_9963,N_9824,N_9882);
nand U9964 (N_9964,N_9817,N_9883);
xnor U9965 (N_9965,N_9872,N_9846);
nor U9966 (N_9966,N_9823,N_9871);
and U9967 (N_9967,N_9815,N_9890);
xor U9968 (N_9968,N_9810,N_9851);
nand U9969 (N_9969,N_9845,N_9885);
xnor U9970 (N_9970,N_9883,N_9847);
and U9971 (N_9971,N_9857,N_9813);
nor U9972 (N_9972,N_9831,N_9806);
nor U9973 (N_9973,N_9850,N_9891);
and U9974 (N_9974,N_9884,N_9861);
or U9975 (N_9975,N_9804,N_9823);
or U9976 (N_9976,N_9851,N_9874);
nand U9977 (N_9977,N_9849,N_9835);
or U9978 (N_9978,N_9873,N_9807);
or U9979 (N_9979,N_9884,N_9848);
nor U9980 (N_9980,N_9896,N_9899);
nand U9981 (N_9981,N_9880,N_9811);
nand U9982 (N_9982,N_9831,N_9854);
and U9983 (N_9983,N_9862,N_9831);
xnor U9984 (N_9984,N_9869,N_9893);
nand U9985 (N_9985,N_9849,N_9881);
and U9986 (N_9986,N_9886,N_9822);
or U9987 (N_9987,N_9895,N_9847);
nor U9988 (N_9988,N_9891,N_9899);
xor U9989 (N_9989,N_9828,N_9864);
xor U9990 (N_9990,N_9854,N_9876);
nand U9991 (N_9991,N_9884,N_9818);
nor U9992 (N_9992,N_9889,N_9816);
nor U9993 (N_9993,N_9870,N_9813);
nor U9994 (N_9994,N_9852,N_9863);
or U9995 (N_9995,N_9836,N_9824);
or U9996 (N_9996,N_9800,N_9834);
or U9997 (N_9997,N_9824,N_9860);
or U9998 (N_9998,N_9814,N_9832);
nor U9999 (N_9999,N_9894,N_9849);
nor UO_0 (O_0,N_9905,N_9972);
or UO_1 (O_1,N_9992,N_9941);
and UO_2 (O_2,N_9961,N_9919);
nand UO_3 (O_3,N_9901,N_9999);
nor UO_4 (O_4,N_9978,N_9913);
xor UO_5 (O_5,N_9957,N_9944);
and UO_6 (O_6,N_9929,N_9998);
or UO_7 (O_7,N_9994,N_9937);
and UO_8 (O_8,N_9907,N_9977);
or UO_9 (O_9,N_9952,N_9946);
or UO_10 (O_10,N_9993,N_9967);
xnor UO_11 (O_11,N_9960,N_9908);
nand UO_12 (O_12,N_9911,N_9902);
and UO_13 (O_13,N_9951,N_9940);
xnor UO_14 (O_14,N_9943,N_9949);
and UO_15 (O_15,N_9931,N_9922);
and UO_16 (O_16,N_9932,N_9981);
or UO_17 (O_17,N_9950,N_9991);
nand UO_18 (O_18,N_9997,N_9973);
or UO_19 (O_19,N_9953,N_9924);
nor UO_20 (O_20,N_9984,N_9986);
xnor UO_21 (O_21,N_9926,N_9916);
nand UO_22 (O_22,N_9923,N_9963);
and UO_23 (O_23,N_9910,N_9959);
nor UO_24 (O_24,N_9955,N_9915);
nand UO_25 (O_25,N_9996,N_9925);
nor UO_26 (O_26,N_9975,N_9964);
or UO_27 (O_27,N_9939,N_9930);
nor UO_28 (O_28,N_9969,N_9983);
xnor UO_29 (O_29,N_9979,N_9980);
nor UO_30 (O_30,N_9935,N_9938);
or UO_31 (O_31,N_9965,N_9914);
nand UO_32 (O_32,N_9958,N_9968);
nor UO_33 (O_33,N_9985,N_9921);
and UO_34 (O_34,N_9989,N_9966);
and UO_35 (O_35,N_9962,N_9927);
nand UO_36 (O_36,N_9945,N_9900);
nand UO_37 (O_37,N_9912,N_9909);
or UO_38 (O_38,N_9948,N_9904);
and UO_39 (O_39,N_9920,N_9974);
xnor UO_40 (O_40,N_9990,N_9956);
nor UO_41 (O_41,N_9995,N_9934);
xnor UO_42 (O_42,N_9954,N_9988);
nor UO_43 (O_43,N_9982,N_9917);
nand UO_44 (O_44,N_9976,N_9942);
or UO_45 (O_45,N_9906,N_9918);
xor UO_46 (O_46,N_9933,N_9903);
and UO_47 (O_47,N_9971,N_9987);
or UO_48 (O_48,N_9936,N_9947);
xor UO_49 (O_49,N_9928,N_9970);
nor UO_50 (O_50,N_9965,N_9980);
or UO_51 (O_51,N_9975,N_9954);
and UO_52 (O_52,N_9951,N_9921);
nand UO_53 (O_53,N_9975,N_9921);
nand UO_54 (O_54,N_9988,N_9975);
and UO_55 (O_55,N_9940,N_9971);
or UO_56 (O_56,N_9964,N_9943);
and UO_57 (O_57,N_9931,N_9928);
and UO_58 (O_58,N_9933,N_9938);
nor UO_59 (O_59,N_9983,N_9900);
and UO_60 (O_60,N_9990,N_9964);
or UO_61 (O_61,N_9999,N_9916);
nand UO_62 (O_62,N_9947,N_9990);
nor UO_63 (O_63,N_9958,N_9900);
nor UO_64 (O_64,N_9915,N_9987);
nor UO_65 (O_65,N_9966,N_9994);
xnor UO_66 (O_66,N_9979,N_9928);
and UO_67 (O_67,N_9992,N_9924);
xnor UO_68 (O_68,N_9911,N_9972);
nor UO_69 (O_69,N_9937,N_9947);
nand UO_70 (O_70,N_9957,N_9902);
or UO_71 (O_71,N_9916,N_9925);
and UO_72 (O_72,N_9951,N_9965);
or UO_73 (O_73,N_9949,N_9909);
nor UO_74 (O_74,N_9942,N_9909);
nor UO_75 (O_75,N_9946,N_9916);
nand UO_76 (O_76,N_9938,N_9950);
and UO_77 (O_77,N_9925,N_9909);
xnor UO_78 (O_78,N_9956,N_9928);
nand UO_79 (O_79,N_9985,N_9940);
and UO_80 (O_80,N_9963,N_9995);
or UO_81 (O_81,N_9938,N_9966);
and UO_82 (O_82,N_9983,N_9953);
xor UO_83 (O_83,N_9990,N_9908);
xnor UO_84 (O_84,N_9947,N_9974);
nand UO_85 (O_85,N_9949,N_9983);
xnor UO_86 (O_86,N_9997,N_9946);
nand UO_87 (O_87,N_9902,N_9963);
nand UO_88 (O_88,N_9998,N_9995);
nand UO_89 (O_89,N_9910,N_9994);
nor UO_90 (O_90,N_9966,N_9996);
nor UO_91 (O_91,N_9912,N_9928);
and UO_92 (O_92,N_9940,N_9911);
and UO_93 (O_93,N_9966,N_9984);
or UO_94 (O_94,N_9947,N_9972);
nor UO_95 (O_95,N_9923,N_9913);
and UO_96 (O_96,N_9924,N_9919);
nand UO_97 (O_97,N_9995,N_9990);
nor UO_98 (O_98,N_9963,N_9996);
nor UO_99 (O_99,N_9918,N_9967);
xor UO_100 (O_100,N_9944,N_9964);
or UO_101 (O_101,N_9937,N_9987);
nand UO_102 (O_102,N_9923,N_9951);
xor UO_103 (O_103,N_9988,N_9913);
and UO_104 (O_104,N_9963,N_9929);
or UO_105 (O_105,N_9907,N_9957);
and UO_106 (O_106,N_9980,N_9929);
or UO_107 (O_107,N_9946,N_9945);
and UO_108 (O_108,N_9931,N_9919);
and UO_109 (O_109,N_9936,N_9950);
nor UO_110 (O_110,N_9959,N_9980);
nand UO_111 (O_111,N_9988,N_9945);
nor UO_112 (O_112,N_9908,N_9959);
nand UO_113 (O_113,N_9998,N_9949);
or UO_114 (O_114,N_9914,N_9912);
nor UO_115 (O_115,N_9934,N_9979);
xnor UO_116 (O_116,N_9952,N_9975);
xor UO_117 (O_117,N_9917,N_9996);
nand UO_118 (O_118,N_9909,N_9984);
and UO_119 (O_119,N_9979,N_9989);
nor UO_120 (O_120,N_9926,N_9999);
nand UO_121 (O_121,N_9948,N_9980);
and UO_122 (O_122,N_9995,N_9930);
or UO_123 (O_123,N_9968,N_9937);
xor UO_124 (O_124,N_9938,N_9908);
nor UO_125 (O_125,N_9926,N_9980);
nor UO_126 (O_126,N_9956,N_9907);
nand UO_127 (O_127,N_9968,N_9960);
and UO_128 (O_128,N_9946,N_9964);
nand UO_129 (O_129,N_9991,N_9934);
nor UO_130 (O_130,N_9947,N_9907);
xor UO_131 (O_131,N_9914,N_9952);
and UO_132 (O_132,N_9974,N_9906);
or UO_133 (O_133,N_9966,N_9981);
and UO_134 (O_134,N_9903,N_9959);
nand UO_135 (O_135,N_9935,N_9902);
and UO_136 (O_136,N_9961,N_9909);
nand UO_137 (O_137,N_9908,N_9911);
nor UO_138 (O_138,N_9916,N_9953);
nor UO_139 (O_139,N_9982,N_9933);
nand UO_140 (O_140,N_9992,N_9949);
xor UO_141 (O_141,N_9996,N_9989);
nor UO_142 (O_142,N_9901,N_9935);
and UO_143 (O_143,N_9916,N_9903);
xor UO_144 (O_144,N_9915,N_9971);
nor UO_145 (O_145,N_9993,N_9948);
nand UO_146 (O_146,N_9958,N_9961);
and UO_147 (O_147,N_9901,N_9914);
and UO_148 (O_148,N_9904,N_9956);
xnor UO_149 (O_149,N_9978,N_9909);
nand UO_150 (O_150,N_9936,N_9991);
nor UO_151 (O_151,N_9930,N_9971);
and UO_152 (O_152,N_9969,N_9933);
nor UO_153 (O_153,N_9937,N_9989);
nor UO_154 (O_154,N_9988,N_9948);
nor UO_155 (O_155,N_9945,N_9906);
nand UO_156 (O_156,N_9906,N_9900);
and UO_157 (O_157,N_9980,N_9925);
xor UO_158 (O_158,N_9906,N_9926);
or UO_159 (O_159,N_9989,N_9939);
or UO_160 (O_160,N_9992,N_9943);
xnor UO_161 (O_161,N_9979,N_9969);
or UO_162 (O_162,N_9921,N_9995);
nor UO_163 (O_163,N_9928,N_9980);
xor UO_164 (O_164,N_9983,N_9936);
nor UO_165 (O_165,N_9992,N_9974);
nor UO_166 (O_166,N_9921,N_9970);
nor UO_167 (O_167,N_9952,N_9937);
and UO_168 (O_168,N_9958,N_9934);
nand UO_169 (O_169,N_9974,N_9971);
and UO_170 (O_170,N_9920,N_9991);
or UO_171 (O_171,N_9947,N_9956);
xor UO_172 (O_172,N_9996,N_9927);
xnor UO_173 (O_173,N_9930,N_9976);
or UO_174 (O_174,N_9965,N_9915);
nor UO_175 (O_175,N_9950,N_9947);
nor UO_176 (O_176,N_9987,N_9926);
and UO_177 (O_177,N_9961,N_9987);
and UO_178 (O_178,N_9956,N_9931);
nor UO_179 (O_179,N_9941,N_9996);
and UO_180 (O_180,N_9931,N_9913);
nand UO_181 (O_181,N_9901,N_9930);
nand UO_182 (O_182,N_9980,N_9919);
nor UO_183 (O_183,N_9965,N_9982);
or UO_184 (O_184,N_9900,N_9959);
nor UO_185 (O_185,N_9943,N_9932);
nand UO_186 (O_186,N_9955,N_9971);
and UO_187 (O_187,N_9968,N_9946);
or UO_188 (O_188,N_9983,N_9979);
xnor UO_189 (O_189,N_9983,N_9929);
or UO_190 (O_190,N_9948,N_9900);
or UO_191 (O_191,N_9974,N_9969);
nand UO_192 (O_192,N_9919,N_9979);
nor UO_193 (O_193,N_9943,N_9958);
nand UO_194 (O_194,N_9917,N_9962);
nor UO_195 (O_195,N_9915,N_9984);
or UO_196 (O_196,N_9976,N_9964);
nand UO_197 (O_197,N_9958,N_9903);
nand UO_198 (O_198,N_9953,N_9905);
xor UO_199 (O_199,N_9922,N_9932);
nor UO_200 (O_200,N_9907,N_9948);
xor UO_201 (O_201,N_9915,N_9928);
and UO_202 (O_202,N_9963,N_9960);
or UO_203 (O_203,N_9947,N_9942);
nand UO_204 (O_204,N_9934,N_9904);
nand UO_205 (O_205,N_9945,N_9964);
xor UO_206 (O_206,N_9993,N_9920);
nand UO_207 (O_207,N_9970,N_9922);
nor UO_208 (O_208,N_9945,N_9905);
and UO_209 (O_209,N_9901,N_9922);
or UO_210 (O_210,N_9917,N_9943);
or UO_211 (O_211,N_9911,N_9971);
xor UO_212 (O_212,N_9941,N_9962);
and UO_213 (O_213,N_9915,N_9916);
and UO_214 (O_214,N_9974,N_9988);
nand UO_215 (O_215,N_9947,N_9922);
or UO_216 (O_216,N_9962,N_9988);
or UO_217 (O_217,N_9945,N_9904);
xor UO_218 (O_218,N_9953,N_9941);
and UO_219 (O_219,N_9950,N_9902);
or UO_220 (O_220,N_9908,N_9912);
and UO_221 (O_221,N_9963,N_9987);
xnor UO_222 (O_222,N_9968,N_9987);
or UO_223 (O_223,N_9980,N_9997);
nor UO_224 (O_224,N_9948,N_9938);
nand UO_225 (O_225,N_9972,N_9914);
xnor UO_226 (O_226,N_9974,N_9952);
and UO_227 (O_227,N_9959,N_9911);
nor UO_228 (O_228,N_9908,N_9968);
or UO_229 (O_229,N_9966,N_9970);
nand UO_230 (O_230,N_9931,N_9989);
nand UO_231 (O_231,N_9992,N_9906);
and UO_232 (O_232,N_9908,N_9977);
nand UO_233 (O_233,N_9908,N_9997);
or UO_234 (O_234,N_9959,N_9930);
nor UO_235 (O_235,N_9950,N_9971);
and UO_236 (O_236,N_9957,N_9964);
nor UO_237 (O_237,N_9921,N_9914);
xor UO_238 (O_238,N_9921,N_9987);
nor UO_239 (O_239,N_9938,N_9936);
xnor UO_240 (O_240,N_9936,N_9990);
nand UO_241 (O_241,N_9938,N_9904);
nor UO_242 (O_242,N_9995,N_9964);
or UO_243 (O_243,N_9976,N_9952);
or UO_244 (O_244,N_9971,N_9936);
or UO_245 (O_245,N_9963,N_9969);
xnor UO_246 (O_246,N_9958,N_9920);
and UO_247 (O_247,N_9923,N_9986);
and UO_248 (O_248,N_9989,N_9960);
and UO_249 (O_249,N_9903,N_9975);
nor UO_250 (O_250,N_9991,N_9958);
and UO_251 (O_251,N_9915,N_9927);
nand UO_252 (O_252,N_9965,N_9938);
and UO_253 (O_253,N_9979,N_9924);
nand UO_254 (O_254,N_9944,N_9956);
nor UO_255 (O_255,N_9939,N_9976);
nand UO_256 (O_256,N_9962,N_9959);
nand UO_257 (O_257,N_9925,N_9952);
nor UO_258 (O_258,N_9977,N_9972);
or UO_259 (O_259,N_9934,N_9980);
xnor UO_260 (O_260,N_9922,N_9958);
nor UO_261 (O_261,N_9925,N_9904);
or UO_262 (O_262,N_9911,N_9977);
xor UO_263 (O_263,N_9957,N_9972);
xnor UO_264 (O_264,N_9910,N_9945);
nor UO_265 (O_265,N_9967,N_9938);
nor UO_266 (O_266,N_9927,N_9955);
xnor UO_267 (O_267,N_9999,N_9909);
nor UO_268 (O_268,N_9909,N_9990);
xnor UO_269 (O_269,N_9909,N_9953);
xor UO_270 (O_270,N_9967,N_9969);
or UO_271 (O_271,N_9924,N_9949);
nor UO_272 (O_272,N_9985,N_9999);
nand UO_273 (O_273,N_9940,N_9917);
or UO_274 (O_274,N_9924,N_9925);
and UO_275 (O_275,N_9913,N_9998);
xor UO_276 (O_276,N_9928,N_9945);
and UO_277 (O_277,N_9924,N_9975);
or UO_278 (O_278,N_9961,N_9989);
xor UO_279 (O_279,N_9908,N_9939);
and UO_280 (O_280,N_9951,N_9984);
or UO_281 (O_281,N_9914,N_9900);
and UO_282 (O_282,N_9990,N_9920);
xnor UO_283 (O_283,N_9909,N_9951);
or UO_284 (O_284,N_9943,N_9980);
nor UO_285 (O_285,N_9984,N_9970);
nand UO_286 (O_286,N_9903,N_9979);
nor UO_287 (O_287,N_9922,N_9912);
nor UO_288 (O_288,N_9959,N_9949);
nand UO_289 (O_289,N_9909,N_9960);
and UO_290 (O_290,N_9981,N_9952);
or UO_291 (O_291,N_9972,N_9993);
nand UO_292 (O_292,N_9923,N_9919);
nand UO_293 (O_293,N_9941,N_9995);
and UO_294 (O_294,N_9910,N_9915);
and UO_295 (O_295,N_9972,N_9959);
or UO_296 (O_296,N_9975,N_9927);
xor UO_297 (O_297,N_9959,N_9923);
xor UO_298 (O_298,N_9995,N_9960);
xnor UO_299 (O_299,N_9911,N_9904);
xnor UO_300 (O_300,N_9952,N_9945);
or UO_301 (O_301,N_9974,N_9909);
and UO_302 (O_302,N_9996,N_9919);
nor UO_303 (O_303,N_9967,N_9957);
xor UO_304 (O_304,N_9916,N_9921);
and UO_305 (O_305,N_9922,N_9915);
xor UO_306 (O_306,N_9934,N_9914);
xor UO_307 (O_307,N_9950,N_9953);
or UO_308 (O_308,N_9956,N_9996);
nand UO_309 (O_309,N_9941,N_9936);
nor UO_310 (O_310,N_9915,N_9979);
xnor UO_311 (O_311,N_9955,N_9901);
nand UO_312 (O_312,N_9934,N_9933);
nand UO_313 (O_313,N_9913,N_9902);
and UO_314 (O_314,N_9982,N_9931);
nand UO_315 (O_315,N_9957,N_9982);
and UO_316 (O_316,N_9908,N_9963);
or UO_317 (O_317,N_9907,N_9917);
xor UO_318 (O_318,N_9912,N_9905);
xnor UO_319 (O_319,N_9997,N_9917);
xor UO_320 (O_320,N_9911,N_9942);
xnor UO_321 (O_321,N_9951,N_9982);
or UO_322 (O_322,N_9952,N_9907);
xnor UO_323 (O_323,N_9904,N_9933);
nor UO_324 (O_324,N_9982,N_9922);
nor UO_325 (O_325,N_9958,N_9907);
or UO_326 (O_326,N_9992,N_9960);
or UO_327 (O_327,N_9908,N_9953);
nor UO_328 (O_328,N_9952,N_9930);
nor UO_329 (O_329,N_9997,N_9919);
nor UO_330 (O_330,N_9916,N_9992);
xnor UO_331 (O_331,N_9926,N_9990);
and UO_332 (O_332,N_9921,N_9933);
and UO_333 (O_333,N_9995,N_9931);
nor UO_334 (O_334,N_9954,N_9941);
and UO_335 (O_335,N_9917,N_9988);
nor UO_336 (O_336,N_9980,N_9903);
nor UO_337 (O_337,N_9978,N_9933);
xnor UO_338 (O_338,N_9984,N_9954);
nand UO_339 (O_339,N_9936,N_9902);
and UO_340 (O_340,N_9988,N_9936);
xor UO_341 (O_341,N_9913,N_9951);
or UO_342 (O_342,N_9986,N_9916);
nor UO_343 (O_343,N_9909,N_9924);
and UO_344 (O_344,N_9997,N_9979);
and UO_345 (O_345,N_9990,N_9954);
and UO_346 (O_346,N_9957,N_9900);
and UO_347 (O_347,N_9902,N_9920);
and UO_348 (O_348,N_9966,N_9988);
nand UO_349 (O_349,N_9968,N_9972);
and UO_350 (O_350,N_9975,N_9941);
nand UO_351 (O_351,N_9909,N_9986);
nor UO_352 (O_352,N_9978,N_9929);
xnor UO_353 (O_353,N_9981,N_9910);
or UO_354 (O_354,N_9951,N_9928);
nand UO_355 (O_355,N_9963,N_9989);
or UO_356 (O_356,N_9969,N_9957);
and UO_357 (O_357,N_9975,N_9904);
and UO_358 (O_358,N_9986,N_9921);
and UO_359 (O_359,N_9956,N_9971);
nor UO_360 (O_360,N_9947,N_9951);
nand UO_361 (O_361,N_9961,N_9944);
xor UO_362 (O_362,N_9914,N_9976);
or UO_363 (O_363,N_9956,N_9942);
xor UO_364 (O_364,N_9925,N_9912);
and UO_365 (O_365,N_9983,N_9928);
or UO_366 (O_366,N_9985,N_9971);
and UO_367 (O_367,N_9967,N_9964);
nand UO_368 (O_368,N_9928,N_9905);
nand UO_369 (O_369,N_9994,N_9963);
and UO_370 (O_370,N_9953,N_9990);
nand UO_371 (O_371,N_9923,N_9912);
xnor UO_372 (O_372,N_9980,N_9990);
and UO_373 (O_373,N_9986,N_9922);
nor UO_374 (O_374,N_9909,N_9991);
nand UO_375 (O_375,N_9960,N_9971);
or UO_376 (O_376,N_9966,N_9949);
and UO_377 (O_377,N_9977,N_9943);
or UO_378 (O_378,N_9983,N_9990);
nand UO_379 (O_379,N_9931,N_9920);
and UO_380 (O_380,N_9968,N_9916);
xnor UO_381 (O_381,N_9958,N_9963);
or UO_382 (O_382,N_9914,N_9948);
nand UO_383 (O_383,N_9916,N_9997);
or UO_384 (O_384,N_9921,N_9946);
nand UO_385 (O_385,N_9900,N_9984);
or UO_386 (O_386,N_9934,N_9984);
xnor UO_387 (O_387,N_9921,N_9948);
and UO_388 (O_388,N_9965,N_9930);
or UO_389 (O_389,N_9903,N_9950);
nand UO_390 (O_390,N_9977,N_9906);
and UO_391 (O_391,N_9974,N_9989);
nor UO_392 (O_392,N_9935,N_9928);
nand UO_393 (O_393,N_9966,N_9977);
or UO_394 (O_394,N_9939,N_9997);
and UO_395 (O_395,N_9928,N_9952);
or UO_396 (O_396,N_9913,N_9989);
or UO_397 (O_397,N_9917,N_9995);
or UO_398 (O_398,N_9998,N_9918);
or UO_399 (O_399,N_9995,N_9961);
nand UO_400 (O_400,N_9991,N_9954);
nand UO_401 (O_401,N_9945,N_9917);
or UO_402 (O_402,N_9962,N_9923);
nor UO_403 (O_403,N_9958,N_9953);
or UO_404 (O_404,N_9953,N_9960);
xor UO_405 (O_405,N_9928,N_9991);
nor UO_406 (O_406,N_9989,N_9955);
nand UO_407 (O_407,N_9910,N_9966);
nand UO_408 (O_408,N_9930,N_9932);
xnor UO_409 (O_409,N_9984,N_9962);
xnor UO_410 (O_410,N_9991,N_9977);
or UO_411 (O_411,N_9960,N_9927);
nand UO_412 (O_412,N_9904,N_9950);
or UO_413 (O_413,N_9976,N_9919);
and UO_414 (O_414,N_9955,N_9912);
nand UO_415 (O_415,N_9901,N_9945);
nor UO_416 (O_416,N_9999,N_9968);
nand UO_417 (O_417,N_9967,N_9970);
and UO_418 (O_418,N_9996,N_9955);
nand UO_419 (O_419,N_9930,N_9960);
nor UO_420 (O_420,N_9949,N_9914);
or UO_421 (O_421,N_9986,N_9962);
and UO_422 (O_422,N_9932,N_9948);
and UO_423 (O_423,N_9935,N_9939);
and UO_424 (O_424,N_9995,N_9977);
and UO_425 (O_425,N_9973,N_9924);
nand UO_426 (O_426,N_9971,N_9964);
nor UO_427 (O_427,N_9928,N_9907);
nor UO_428 (O_428,N_9970,N_9947);
nand UO_429 (O_429,N_9976,N_9913);
and UO_430 (O_430,N_9927,N_9994);
nand UO_431 (O_431,N_9944,N_9963);
nand UO_432 (O_432,N_9972,N_9951);
or UO_433 (O_433,N_9996,N_9949);
or UO_434 (O_434,N_9941,N_9932);
xnor UO_435 (O_435,N_9977,N_9936);
and UO_436 (O_436,N_9995,N_9944);
and UO_437 (O_437,N_9971,N_9961);
nand UO_438 (O_438,N_9994,N_9942);
and UO_439 (O_439,N_9978,N_9932);
nor UO_440 (O_440,N_9996,N_9924);
nor UO_441 (O_441,N_9951,N_9910);
nand UO_442 (O_442,N_9964,N_9925);
nor UO_443 (O_443,N_9984,N_9941);
xnor UO_444 (O_444,N_9904,N_9942);
or UO_445 (O_445,N_9960,N_9999);
nand UO_446 (O_446,N_9955,N_9924);
xor UO_447 (O_447,N_9986,N_9950);
or UO_448 (O_448,N_9971,N_9967);
xnor UO_449 (O_449,N_9916,N_9962);
nor UO_450 (O_450,N_9926,N_9963);
or UO_451 (O_451,N_9968,N_9953);
and UO_452 (O_452,N_9961,N_9998);
xnor UO_453 (O_453,N_9906,N_9944);
xnor UO_454 (O_454,N_9917,N_9909);
nand UO_455 (O_455,N_9945,N_9971);
xor UO_456 (O_456,N_9932,N_9931);
nor UO_457 (O_457,N_9994,N_9948);
or UO_458 (O_458,N_9974,N_9943);
xnor UO_459 (O_459,N_9940,N_9991);
nor UO_460 (O_460,N_9997,N_9925);
nor UO_461 (O_461,N_9938,N_9984);
or UO_462 (O_462,N_9936,N_9915);
nand UO_463 (O_463,N_9986,N_9987);
xor UO_464 (O_464,N_9900,N_9966);
nor UO_465 (O_465,N_9949,N_9933);
nand UO_466 (O_466,N_9919,N_9913);
xor UO_467 (O_467,N_9935,N_9921);
or UO_468 (O_468,N_9960,N_9951);
and UO_469 (O_469,N_9995,N_9908);
xnor UO_470 (O_470,N_9964,N_9908);
nor UO_471 (O_471,N_9936,N_9953);
nor UO_472 (O_472,N_9994,N_9939);
xor UO_473 (O_473,N_9988,N_9914);
and UO_474 (O_474,N_9967,N_9921);
nand UO_475 (O_475,N_9996,N_9935);
and UO_476 (O_476,N_9980,N_9961);
nor UO_477 (O_477,N_9926,N_9940);
or UO_478 (O_478,N_9902,N_9908);
xor UO_479 (O_479,N_9976,N_9967);
and UO_480 (O_480,N_9951,N_9920);
or UO_481 (O_481,N_9944,N_9962);
xor UO_482 (O_482,N_9971,N_9980);
nor UO_483 (O_483,N_9930,N_9902);
nor UO_484 (O_484,N_9964,N_9914);
or UO_485 (O_485,N_9982,N_9921);
or UO_486 (O_486,N_9941,N_9955);
and UO_487 (O_487,N_9997,N_9943);
xnor UO_488 (O_488,N_9982,N_9963);
nor UO_489 (O_489,N_9947,N_9949);
or UO_490 (O_490,N_9913,N_9927);
xor UO_491 (O_491,N_9901,N_9903);
or UO_492 (O_492,N_9933,N_9984);
xor UO_493 (O_493,N_9936,N_9944);
or UO_494 (O_494,N_9961,N_9933);
and UO_495 (O_495,N_9901,N_9978);
or UO_496 (O_496,N_9910,N_9950);
nand UO_497 (O_497,N_9926,N_9938);
nor UO_498 (O_498,N_9981,N_9904);
or UO_499 (O_499,N_9981,N_9901);
xnor UO_500 (O_500,N_9948,N_9970);
or UO_501 (O_501,N_9929,N_9976);
nand UO_502 (O_502,N_9949,N_9930);
nand UO_503 (O_503,N_9939,N_9983);
nand UO_504 (O_504,N_9968,N_9982);
and UO_505 (O_505,N_9963,N_9912);
and UO_506 (O_506,N_9972,N_9956);
nand UO_507 (O_507,N_9983,N_9958);
or UO_508 (O_508,N_9953,N_9964);
nor UO_509 (O_509,N_9913,N_9983);
and UO_510 (O_510,N_9918,N_9949);
or UO_511 (O_511,N_9920,N_9972);
or UO_512 (O_512,N_9927,N_9901);
and UO_513 (O_513,N_9949,N_9929);
or UO_514 (O_514,N_9917,N_9928);
and UO_515 (O_515,N_9936,N_9910);
and UO_516 (O_516,N_9961,N_9941);
and UO_517 (O_517,N_9961,N_9924);
nor UO_518 (O_518,N_9914,N_9905);
or UO_519 (O_519,N_9929,N_9920);
xnor UO_520 (O_520,N_9940,N_9960);
xnor UO_521 (O_521,N_9967,N_9960);
nand UO_522 (O_522,N_9919,N_9991);
nand UO_523 (O_523,N_9912,N_9988);
or UO_524 (O_524,N_9935,N_9931);
nor UO_525 (O_525,N_9979,N_9927);
nor UO_526 (O_526,N_9923,N_9960);
xor UO_527 (O_527,N_9967,N_9950);
nand UO_528 (O_528,N_9955,N_9968);
xnor UO_529 (O_529,N_9916,N_9932);
xnor UO_530 (O_530,N_9912,N_9990);
and UO_531 (O_531,N_9980,N_9927);
nand UO_532 (O_532,N_9974,N_9983);
nand UO_533 (O_533,N_9937,N_9940);
nor UO_534 (O_534,N_9936,N_9957);
xnor UO_535 (O_535,N_9962,N_9958);
nand UO_536 (O_536,N_9933,N_9919);
or UO_537 (O_537,N_9958,N_9904);
nor UO_538 (O_538,N_9908,N_9986);
nand UO_539 (O_539,N_9928,N_9976);
and UO_540 (O_540,N_9979,N_9972);
nand UO_541 (O_541,N_9983,N_9947);
xor UO_542 (O_542,N_9905,N_9951);
nand UO_543 (O_543,N_9985,N_9981);
nand UO_544 (O_544,N_9901,N_9932);
and UO_545 (O_545,N_9950,N_9993);
xor UO_546 (O_546,N_9985,N_9950);
and UO_547 (O_547,N_9902,N_9997);
nor UO_548 (O_548,N_9989,N_9970);
nor UO_549 (O_549,N_9926,N_9958);
and UO_550 (O_550,N_9922,N_9972);
nor UO_551 (O_551,N_9907,N_9975);
nand UO_552 (O_552,N_9918,N_9985);
and UO_553 (O_553,N_9980,N_9976);
nor UO_554 (O_554,N_9945,N_9944);
or UO_555 (O_555,N_9906,N_9904);
xor UO_556 (O_556,N_9913,N_9905);
nor UO_557 (O_557,N_9987,N_9902);
nor UO_558 (O_558,N_9915,N_9989);
xor UO_559 (O_559,N_9906,N_9953);
xor UO_560 (O_560,N_9924,N_9991);
and UO_561 (O_561,N_9949,N_9912);
nor UO_562 (O_562,N_9907,N_9960);
and UO_563 (O_563,N_9912,N_9944);
or UO_564 (O_564,N_9969,N_9962);
and UO_565 (O_565,N_9926,N_9966);
xor UO_566 (O_566,N_9963,N_9953);
or UO_567 (O_567,N_9907,N_9905);
xor UO_568 (O_568,N_9980,N_9988);
xor UO_569 (O_569,N_9931,N_9949);
xnor UO_570 (O_570,N_9904,N_9917);
nand UO_571 (O_571,N_9928,N_9995);
nand UO_572 (O_572,N_9921,N_9913);
and UO_573 (O_573,N_9968,N_9996);
and UO_574 (O_574,N_9952,N_9938);
nand UO_575 (O_575,N_9933,N_9925);
and UO_576 (O_576,N_9993,N_9971);
or UO_577 (O_577,N_9992,N_9902);
and UO_578 (O_578,N_9943,N_9983);
nor UO_579 (O_579,N_9932,N_9909);
nand UO_580 (O_580,N_9973,N_9959);
nand UO_581 (O_581,N_9978,N_9939);
xor UO_582 (O_582,N_9911,N_9955);
xor UO_583 (O_583,N_9949,N_9980);
or UO_584 (O_584,N_9910,N_9961);
and UO_585 (O_585,N_9981,N_9975);
or UO_586 (O_586,N_9928,N_9924);
nand UO_587 (O_587,N_9947,N_9903);
nand UO_588 (O_588,N_9990,N_9931);
and UO_589 (O_589,N_9965,N_9956);
or UO_590 (O_590,N_9958,N_9937);
xor UO_591 (O_591,N_9964,N_9997);
or UO_592 (O_592,N_9915,N_9990);
nand UO_593 (O_593,N_9954,N_9970);
nand UO_594 (O_594,N_9920,N_9976);
or UO_595 (O_595,N_9952,N_9910);
xnor UO_596 (O_596,N_9986,N_9911);
or UO_597 (O_597,N_9956,N_9901);
and UO_598 (O_598,N_9906,N_9907);
xnor UO_599 (O_599,N_9928,N_9959);
nand UO_600 (O_600,N_9980,N_9954);
nor UO_601 (O_601,N_9909,N_9983);
or UO_602 (O_602,N_9991,N_9993);
nand UO_603 (O_603,N_9996,N_9930);
nor UO_604 (O_604,N_9972,N_9954);
xor UO_605 (O_605,N_9996,N_9940);
and UO_606 (O_606,N_9905,N_9938);
or UO_607 (O_607,N_9940,N_9962);
and UO_608 (O_608,N_9977,N_9996);
nor UO_609 (O_609,N_9920,N_9941);
xnor UO_610 (O_610,N_9923,N_9920);
and UO_611 (O_611,N_9911,N_9913);
xor UO_612 (O_612,N_9960,N_9966);
or UO_613 (O_613,N_9987,N_9930);
or UO_614 (O_614,N_9900,N_9976);
nor UO_615 (O_615,N_9927,N_9900);
nor UO_616 (O_616,N_9976,N_9925);
xnor UO_617 (O_617,N_9995,N_9927);
nor UO_618 (O_618,N_9924,N_9910);
xor UO_619 (O_619,N_9919,N_9902);
xor UO_620 (O_620,N_9903,N_9921);
nand UO_621 (O_621,N_9957,N_9973);
xor UO_622 (O_622,N_9903,N_9977);
or UO_623 (O_623,N_9937,N_9909);
xor UO_624 (O_624,N_9918,N_9912);
or UO_625 (O_625,N_9951,N_9998);
xor UO_626 (O_626,N_9911,N_9999);
xor UO_627 (O_627,N_9934,N_9963);
and UO_628 (O_628,N_9962,N_9973);
nor UO_629 (O_629,N_9932,N_9950);
and UO_630 (O_630,N_9934,N_9928);
and UO_631 (O_631,N_9985,N_9907);
nand UO_632 (O_632,N_9913,N_9906);
nor UO_633 (O_633,N_9907,N_9989);
nor UO_634 (O_634,N_9941,N_9933);
or UO_635 (O_635,N_9924,N_9965);
xor UO_636 (O_636,N_9990,N_9942);
or UO_637 (O_637,N_9991,N_9943);
nand UO_638 (O_638,N_9990,N_9994);
nor UO_639 (O_639,N_9969,N_9901);
nand UO_640 (O_640,N_9968,N_9941);
xor UO_641 (O_641,N_9984,N_9920);
or UO_642 (O_642,N_9946,N_9962);
nand UO_643 (O_643,N_9982,N_9918);
nand UO_644 (O_644,N_9955,N_9947);
and UO_645 (O_645,N_9960,N_9915);
nor UO_646 (O_646,N_9919,N_9975);
or UO_647 (O_647,N_9949,N_9923);
or UO_648 (O_648,N_9930,N_9967);
xor UO_649 (O_649,N_9910,N_9967);
and UO_650 (O_650,N_9995,N_9994);
nor UO_651 (O_651,N_9907,N_9976);
nor UO_652 (O_652,N_9980,N_9987);
xnor UO_653 (O_653,N_9992,N_9998);
and UO_654 (O_654,N_9936,N_9945);
and UO_655 (O_655,N_9922,N_9974);
and UO_656 (O_656,N_9929,N_9926);
nor UO_657 (O_657,N_9995,N_9965);
nand UO_658 (O_658,N_9968,N_9934);
and UO_659 (O_659,N_9913,N_9903);
nand UO_660 (O_660,N_9940,N_9980);
xnor UO_661 (O_661,N_9957,N_9927);
nand UO_662 (O_662,N_9953,N_9994);
nor UO_663 (O_663,N_9902,N_9976);
xnor UO_664 (O_664,N_9975,N_9939);
xor UO_665 (O_665,N_9918,N_9900);
or UO_666 (O_666,N_9976,N_9991);
and UO_667 (O_667,N_9958,N_9995);
xnor UO_668 (O_668,N_9985,N_9942);
xnor UO_669 (O_669,N_9993,N_9941);
and UO_670 (O_670,N_9991,N_9980);
xor UO_671 (O_671,N_9985,N_9995);
xor UO_672 (O_672,N_9937,N_9929);
nor UO_673 (O_673,N_9902,N_9979);
or UO_674 (O_674,N_9997,N_9938);
nand UO_675 (O_675,N_9973,N_9917);
nor UO_676 (O_676,N_9901,N_9915);
xor UO_677 (O_677,N_9957,N_9920);
and UO_678 (O_678,N_9979,N_9998);
or UO_679 (O_679,N_9949,N_9927);
and UO_680 (O_680,N_9908,N_9903);
and UO_681 (O_681,N_9912,N_9948);
xor UO_682 (O_682,N_9917,N_9946);
and UO_683 (O_683,N_9990,N_9929);
nor UO_684 (O_684,N_9923,N_9999);
nand UO_685 (O_685,N_9928,N_9901);
or UO_686 (O_686,N_9925,N_9918);
nand UO_687 (O_687,N_9983,N_9952);
or UO_688 (O_688,N_9905,N_9960);
and UO_689 (O_689,N_9929,N_9936);
xor UO_690 (O_690,N_9908,N_9970);
or UO_691 (O_691,N_9963,N_9932);
nor UO_692 (O_692,N_9923,N_9901);
or UO_693 (O_693,N_9971,N_9963);
nor UO_694 (O_694,N_9932,N_9957);
nor UO_695 (O_695,N_9946,N_9920);
or UO_696 (O_696,N_9934,N_9931);
nor UO_697 (O_697,N_9927,N_9917);
xnor UO_698 (O_698,N_9971,N_9996);
or UO_699 (O_699,N_9904,N_9901);
and UO_700 (O_700,N_9915,N_9993);
or UO_701 (O_701,N_9969,N_9926);
nor UO_702 (O_702,N_9978,N_9912);
and UO_703 (O_703,N_9980,N_9901);
or UO_704 (O_704,N_9911,N_9981);
or UO_705 (O_705,N_9956,N_9934);
nand UO_706 (O_706,N_9927,N_9934);
xnor UO_707 (O_707,N_9994,N_9922);
or UO_708 (O_708,N_9939,N_9907);
xor UO_709 (O_709,N_9915,N_9959);
or UO_710 (O_710,N_9990,N_9998);
nand UO_711 (O_711,N_9904,N_9954);
and UO_712 (O_712,N_9929,N_9905);
nor UO_713 (O_713,N_9915,N_9947);
xnor UO_714 (O_714,N_9997,N_9935);
and UO_715 (O_715,N_9975,N_9985);
or UO_716 (O_716,N_9935,N_9926);
nor UO_717 (O_717,N_9920,N_9927);
nor UO_718 (O_718,N_9986,N_9994);
or UO_719 (O_719,N_9921,N_9938);
or UO_720 (O_720,N_9963,N_9946);
and UO_721 (O_721,N_9940,N_9997);
or UO_722 (O_722,N_9941,N_9988);
nand UO_723 (O_723,N_9957,N_9903);
nor UO_724 (O_724,N_9929,N_9939);
xor UO_725 (O_725,N_9901,N_9987);
nor UO_726 (O_726,N_9917,N_9974);
nor UO_727 (O_727,N_9938,N_9998);
and UO_728 (O_728,N_9935,N_9937);
nor UO_729 (O_729,N_9943,N_9972);
xnor UO_730 (O_730,N_9929,N_9911);
xnor UO_731 (O_731,N_9925,N_9914);
xnor UO_732 (O_732,N_9975,N_9945);
or UO_733 (O_733,N_9910,N_9993);
and UO_734 (O_734,N_9937,N_9907);
or UO_735 (O_735,N_9967,N_9968);
or UO_736 (O_736,N_9936,N_9979);
or UO_737 (O_737,N_9930,N_9981);
nand UO_738 (O_738,N_9962,N_9928);
and UO_739 (O_739,N_9963,N_9972);
xnor UO_740 (O_740,N_9935,N_9914);
nor UO_741 (O_741,N_9959,N_9902);
and UO_742 (O_742,N_9900,N_9949);
nor UO_743 (O_743,N_9953,N_9914);
xor UO_744 (O_744,N_9955,N_9910);
xor UO_745 (O_745,N_9930,N_9924);
xor UO_746 (O_746,N_9910,N_9953);
or UO_747 (O_747,N_9993,N_9924);
nor UO_748 (O_748,N_9906,N_9997);
xnor UO_749 (O_749,N_9944,N_9913);
or UO_750 (O_750,N_9964,N_9930);
and UO_751 (O_751,N_9943,N_9971);
nor UO_752 (O_752,N_9952,N_9915);
nand UO_753 (O_753,N_9974,N_9980);
nand UO_754 (O_754,N_9940,N_9930);
and UO_755 (O_755,N_9987,N_9966);
or UO_756 (O_756,N_9976,N_9906);
nor UO_757 (O_757,N_9921,N_9943);
nand UO_758 (O_758,N_9944,N_9978);
xor UO_759 (O_759,N_9998,N_9964);
or UO_760 (O_760,N_9906,N_9983);
xor UO_761 (O_761,N_9918,N_9981);
nand UO_762 (O_762,N_9906,N_9937);
nor UO_763 (O_763,N_9948,N_9995);
or UO_764 (O_764,N_9960,N_9932);
nor UO_765 (O_765,N_9974,N_9951);
xor UO_766 (O_766,N_9987,N_9990);
nand UO_767 (O_767,N_9973,N_9968);
and UO_768 (O_768,N_9997,N_9920);
and UO_769 (O_769,N_9932,N_9994);
and UO_770 (O_770,N_9911,N_9970);
nand UO_771 (O_771,N_9984,N_9947);
and UO_772 (O_772,N_9950,N_9915);
and UO_773 (O_773,N_9912,N_9983);
nand UO_774 (O_774,N_9936,N_9978);
or UO_775 (O_775,N_9977,N_9935);
and UO_776 (O_776,N_9931,N_9969);
xnor UO_777 (O_777,N_9922,N_9989);
nor UO_778 (O_778,N_9908,N_9917);
xnor UO_779 (O_779,N_9968,N_9978);
nand UO_780 (O_780,N_9959,N_9935);
xor UO_781 (O_781,N_9942,N_9923);
xor UO_782 (O_782,N_9947,N_9933);
nor UO_783 (O_783,N_9971,N_9937);
and UO_784 (O_784,N_9969,N_9978);
and UO_785 (O_785,N_9923,N_9925);
xor UO_786 (O_786,N_9960,N_9913);
nand UO_787 (O_787,N_9936,N_9992);
or UO_788 (O_788,N_9919,N_9981);
xnor UO_789 (O_789,N_9965,N_9955);
nand UO_790 (O_790,N_9918,N_9996);
nor UO_791 (O_791,N_9943,N_9965);
and UO_792 (O_792,N_9943,N_9973);
or UO_793 (O_793,N_9978,N_9983);
nor UO_794 (O_794,N_9966,N_9907);
or UO_795 (O_795,N_9930,N_9975);
and UO_796 (O_796,N_9987,N_9920);
or UO_797 (O_797,N_9918,N_9974);
xnor UO_798 (O_798,N_9942,N_9965);
and UO_799 (O_799,N_9933,N_9915);
nand UO_800 (O_800,N_9990,N_9975);
or UO_801 (O_801,N_9981,N_9942);
nand UO_802 (O_802,N_9959,N_9993);
xor UO_803 (O_803,N_9905,N_9999);
nor UO_804 (O_804,N_9996,N_9922);
or UO_805 (O_805,N_9905,N_9970);
nor UO_806 (O_806,N_9982,N_9960);
xor UO_807 (O_807,N_9981,N_9948);
or UO_808 (O_808,N_9938,N_9913);
nor UO_809 (O_809,N_9920,N_9939);
xnor UO_810 (O_810,N_9926,N_9948);
nand UO_811 (O_811,N_9922,N_9977);
nor UO_812 (O_812,N_9918,N_9908);
xor UO_813 (O_813,N_9957,N_9965);
xor UO_814 (O_814,N_9935,N_9961);
and UO_815 (O_815,N_9922,N_9963);
xnor UO_816 (O_816,N_9907,N_9959);
xnor UO_817 (O_817,N_9927,N_9972);
and UO_818 (O_818,N_9947,N_9982);
nor UO_819 (O_819,N_9979,N_9948);
nor UO_820 (O_820,N_9950,N_9926);
xnor UO_821 (O_821,N_9973,N_9953);
and UO_822 (O_822,N_9983,N_9908);
or UO_823 (O_823,N_9929,N_9904);
or UO_824 (O_824,N_9943,N_9999);
and UO_825 (O_825,N_9913,N_9991);
xnor UO_826 (O_826,N_9967,N_9981);
xor UO_827 (O_827,N_9993,N_9999);
xnor UO_828 (O_828,N_9906,N_9970);
or UO_829 (O_829,N_9993,N_9908);
nand UO_830 (O_830,N_9966,N_9998);
and UO_831 (O_831,N_9901,N_9949);
nor UO_832 (O_832,N_9906,N_9950);
xnor UO_833 (O_833,N_9924,N_9981);
or UO_834 (O_834,N_9925,N_9900);
or UO_835 (O_835,N_9935,N_9908);
xnor UO_836 (O_836,N_9933,N_9975);
and UO_837 (O_837,N_9932,N_9992);
nand UO_838 (O_838,N_9998,N_9928);
or UO_839 (O_839,N_9985,N_9937);
and UO_840 (O_840,N_9934,N_9920);
nor UO_841 (O_841,N_9915,N_9940);
and UO_842 (O_842,N_9962,N_9921);
nand UO_843 (O_843,N_9994,N_9969);
nor UO_844 (O_844,N_9990,N_9925);
nor UO_845 (O_845,N_9909,N_9959);
or UO_846 (O_846,N_9952,N_9951);
nor UO_847 (O_847,N_9953,N_9988);
nor UO_848 (O_848,N_9952,N_9953);
nand UO_849 (O_849,N_9942,N_9959);
nor UO_850 (O_850,N_9930,N_9915);
nor UO_851 (O_851,N_9993,N_9998);
nor UO_852 (O_852,N_9989,N_9901);
nor UO_853 (O_853,N_9920,N_9935);
and UO_854 (O_854,N_9952,N_9989);
or UO_855 (O_855,N_9953,N_9900);
nand UO_856 (O_856,N_9916,N_9938);
xor UO_857 (O_857,N_9974,N_9968);
xor UO_858 (O_858,N_9902,N_9942);
or UO_859 (O_859,N_9950,N_9956);
nand UO_860 (O_860,N_9971,N_9917);
xor UO_861 (O_861,N_9906,N_9902);
and UO_862 (O_862,N_9907,N_9980);
nand UO_863 (O_863,N_9928,N_9972);
nand UO_864 (O_864,N_9965,N_9907);
nor UO_865 (O_865,N_9910,N_9909);
xor UO_866 (O_866,N_9916,N_9939);
nor UO_867 (O_867,N_9986,N_9983);
xnor UO_868 (O_868,N_9933,N_9976);
or UO_869 (O_869,N_9944,N_9993);
nor UO_870 (O_870,N_9960,N_9978);
or UO_871 (O_871,N_9939,N_9967);
nand UO_872 (O_872,N_9989,N_9928);
nand UO_873 (O_873,N_9986,N_9947);
xor UO_874 (O_874,N_9944,N_9918);
nor UO_875 (O_875,N_9974,N_9913);
nand UO_876 (O_876,N_9907,N_9974);
nand UO_877 (O_877,N_9971,N_9907);
nand UO_878 (O_878,N_9987,N_9908);
or UO_879 (O_879,N_9970,N_9990);
or UO_880 (O_880,N_9908,N_9927);
xnor UO_881 (O_881,N_9903,N_9911);
nand UO_882 (O_882,N_9903,N_9922);
xnor UO_883 (O_883,N_9999,N_9913);
nor UO_884 (O_884,N_9991,N_9965);
xnor UO_885 (O_885,N_9917,N_9951);
nand UO_886 (O_886,N_9926,N_9928);
nand UO_887 (O_887,N_9970,N_9903);
or UO_888 (O_888,N_9907,N_9993);
xor UO_889 (O_889,N_9933,N_9924);
xnor UO_890 (O_890,N_9957,N_9989);
or UO_891 (O_891,N_9939,N_9919);
nor UO_892 (O_892,N_9988,N_9930);
nand UO_893 (O_893,N_9985,N_9930);
and UO_894 (O_894,N_9953,N_9974);
nor UO_895 (O_895,N_9910,N_9912);
xor UO_896 (O_896,N_9924,N_9939);
xor UO_897 (O_897,N_9903,N_9928);
and UO_898 (O_898,N_9955,N_9946);
nor UO_899 (O_899,N_9989,N_9916);
nand UO_900 (O_900,N_9901,N_9933);
nor UO_901 (O_901,N_9919,N_9903);
and UO_902 (O_902,N_9935,N_9954);
and UO_903 (O_903,N_9953,N_9946);
nand UO_904 (O_904,N_9920,N_9948);
or UO_905 (O_905,N_9965,N_9973);
xnor UO_906 (O_906,N_9941,N_9928);
nand UO_907 (O_907,N_9986,N_9978);
nor UO_908 (O_908,N_9952,N_9991);
or UO_909 (O_909,N_9973,N_9914);
or UO_910 (O_910,N_9951,N_9995);
or UO_911 (O_911,N_9937,N_9991);
or UO_912 (O_912,N_9976,N_9904);
nor UO_913 (O_913,N_9913,N_9980);
nor UO_914 (O_914,N_9984,N_9910);
or UO_915 (O_915,N_9935,N_9906);
nand UO_916 (O_916,N_9976,N_9940);
nor UO_917 (O_917,N_9934,N_9964);
nor UO_918 (O_918,N_9993,N_9973);
xor UO_919 (O_919,N_9944,N_9980);
nand UO_920 (O_920,N_9953,N_9980);
nor UO_921 (O_921,N_9996,N_9998);
nand UO_922 (O_922,N_9998,N_9904);
or UO_923 (O_923,N_9956,N_9977);
nor UO_924 (O_924,N_9940,N_9949);
xor UO_925 (O_925,N_9917,N_9919);
xnor UO_926 (O_926,N_9921,N_9908);
xor UO_927 (O_927,N_9929,N_9907);
or UO_928 (O_928,N_9941,N_9939);
nor UO_929 (O_929,N_9919,N_9970);
and UO_930 (O_930,N_9951,N_9935);
xor UO_931 (O_931,N_9910,N_9937);
or UO_932 (O_932,N_9953,N_9978);
xnor UO_933 (O_933,N_9960,N_9920);
nor UO_934 (O_934,N_9996,N_9987);
nand UO_935 (O_935,N_9958,N_9956);
nor UO_936 (O_936,N_9940,N_9977);
nor UO_937 (O_937,N_9901,N_9938);
and UO_938 (O_938,N_9926,N_9977);
or UO_939 (O_939,N_9976,N_9994);
nor UO_940 (O_940,N_9957,N_9942);
and UO_941 (O_941,N_9930,N_9905);
nand UO_942 (O_942,N_9980,N_9935);
and UO_943 (O_943,N_9998,N_9943);
nor UO_944 (O_944,N_9937,N_9903);
xor UO_945 (O_945,N_9959,N_9999);
and UO_946 (O_946,N_9931,N_9980);
nor UO_947 (O_947,N_9929,N_9901);
or UO_948 (O_948,N_9927,N_9907);
nand UO_949 (O_949,N_9924,N_9918);
xnor UO_950 (O_950,N_9953,N_9921);
nor UO_951 (O_951,N_9906,N_9954);
or UO_952 (O_952,N_9964,N_9921);
or UO_953 (O_953,N_9914,N_9930);
nand UO_954 (O_954,N_9982,N_9926);
nor UO_955 (O_955,N_9998,N_9903);
and UO_956 (O_956,N_9914,N_9999);
nand UO_957 (O_957,N_9914,N_9975);
nand UO_958 (O_958,N_9987,N_9997);
xor UO_959 (O_959,N_9928,N_9965);
or UO_960 (O_960,N_9922,N_9924);
or UO_961 (O_961,N_9964,N_9996);
xnor UO_962 (O_962,N_9929,N_9918);
nor UO_963 (O_963,N_9998,N_9909);
nor UO_964 (O_964,N_9947,N_9925);
xnor UO_965 (O_965,N_9904,N_9916);
nand UO_966 (O_966,N_9942,N_9945);
and UO_967 (O_967,N_9900,N_9917);
and UO_968 (O_968,N_9966,N_9952);
xor UO_969 (O_969,N_9916,N_9909);
nor UO_970 (O_970,N_9953,N_9955);
nor UO_971 (O_971,N_9919,N_9920);
xnor UO_972 (O_972,N_9928,N_9913);
nand UO_973 (O_973,N_9961,N_9973);
nor UO_974 (O_974,N_9970,N_9907);
xor UO_975 (O_975,N_9955,N_9932);
or UO_976 (O_976,N_9922,N_9908);
nor UO_977 (O_977,N_9947,N_9978);
or UO_978 (O_978,N_9925,N_9913);
xnor UO_979 (O_979,N_9994,N_9918);
nor UO_980 (O_980,N_9957,N_9995);
and UO_981 (O_981,N_9975,N_9901);
xnor UO_982 (O_982,N_9963,N_9924);
or UO_983 (O_983,N_9977,N_9975);
and UO_984 (O_984,N_9920,N_9954);
or UO_985 (O_985,N_9947,N_9920);
nor UO_986 (O_986,N_9945,N_9913);
or UO_987 (O_987,N_9910,N_9956);
and UO_988 (O_988,N_9935,N_9930);
nand UO_989 (O_989,N_9902,N_9978);
xnor UO_990 (O_990,N_9935,N_9944);
nand UO_991 (O_991,N_9933,N_9927);
nand UO_992 (O_992,N_9954,N_9903);
and UO_993 (O_993,N_9946,N_9915);
or UO_994 (O_994,N_9972,N_9949);
nand UO_995 (O_995,N_9998,N_9930);
xnor UO_996 (O_996,N_9946,N_9987);
or UO_997 (O_997,N_9996,N_9904);
nand UO_998 (O_998,N_9976,N_9931);
nand UO_999 (O_999,N_9977,N_9964);
and UO_1000 (O_1000,N_9909,N_9987);
nand UO_1001 (O_1001,N_9967,N_9994);
or UO_1002 (O_1002,N_9984,N_9978);
nand UO_1003 (O_1003,N_9953,N_9982);
nand UO_1004 (O_1004,N_9998,N_9906);
nor UO_1005 (O_1005,N_9990,N_9973);
and UO_1006 (O_1006,N_9976,N_9948);
nand UO_1007 (O_1007,N_9954,N_9974);
xnor UO_1008 (O_1008,N_9971,N_9942);
nor UO_1009 (O_1009,N_9979,N_9954);
nor UO_1010 (O_1010,N_9917,N_9979);
nand UO_1011 (O_1011,N_9967,N_9959);
or UO_1012 (O_1012,N_9960,N_9901);
nand UO_1013 (O_1013,N_9947,N_9948);
or UO_1014 (O_1014,N_9978,N_9981);
xor UO_1015 (O_1015,N_9974,N_9941);
and UO_1016 (O_1016,N_9940,N_9910);
nand UO_1017 (O_1017,N_9908,N_9933);
and UO_1018 (O_1018,N_9920,N_9915);
xnor UO_1019 (O_1019,N_9930,N_9904);
nand UO_1020 (O_1020,N_9912,N_9984);
xor UO_1021 (O_1021,N_9963,N_9980);
and UO_1022 (O_1022,N_9965,N_9927);
nor UO_1023 (O_1023,N_9905,N_9948);
and UO_1024 (O_1024,N_9908,N_9950);
xnor UO_1025 (O_1025,N_9980,N_9950);
nand UO_1026 (O_1026,N_9971,N_9951);
and UO_1027 (O_1027,N_9974,N_9945);
and UO_1028 (O_1028,N_9924,N_9946);
or UO_1029 (O_1029,N_9944,N_9967);
xnor UO_1030 (O_1030,N_9943,N_9906);
or UO_1031 (O_1031,N_9918,N_9916);
and UO_1032 (O_1032,N_9922,N_9969);
nor UO_1033 (O_1033,N_9999,N_9953);
nand UO_1034 (O_1034,N_9999,N_9958);
and UO_1035 (O_1035,N_9993,N_9933);
and UO_1036 (O_1036,N_9966,N_9912);
xnor UO_1037 (O_1037,N_9966,N_9980);
nand UO_1038 (O_1038,N_9940,N_9957);
or UO_1039 (O_1039,N_9998,N_9972);
and UO_1040 (O_1040,N_9960,N_9985);
and UO_1041 (O_1041,N_9923,N_9990);
xnor UO_1042 (O_1042,N_9984,N_9971);
nand UO_1043 (O_1043,N_9967,N_9991);
nand UO_1044 (O_1044,N_9984,N_9911);
xor UO_1045 (O_1045,N_9999,N_9966);
and UO_1046 (O_1046,N_9997,N_9905);
xnor UO_1047 (O_1047,N_9976,N_9968);
or UO_1048 (O_1048,N_9998,N_9934);
or UO_1049 (O_1049,N_9960,N_9981);
nand UO_1050 (O_1050,N_9981,N_9934);
or UO_1051 (O_1051,N_9980,N_9986);
nand UO_1052 (O_1052,N_9927,N_9981);
xor UO_1053 (O_1053,N_9938,N_9986);
xnor UO_1054 (O_1054,N_9937,N_9981);
nor UO_1055 (O_1055,N_9951,N_9953);
xor UO_1056 (O_1056,N_9997,N_9901);
nor UO_1057 (O_1057,N_9992,N_9948);
and UO_1058 (O_1058,N_9944,N_9986);
nor UO_1059 (O_1059,N_9993,N_9914);
nand UO_1060 (O_1060,N_9910,N_9905);
xor UO_1061 (O_1061,N_9933,N_9985);
nor UO_1062 (O_1062,N_9944,N_9940);
nand UO_1063 (O_1063,N_9984,N_9998);
or UO_1064 (O_1064,N_9968,N_9995);
or UO_1065 (O_1065,N_9986,N_9975);
or UO_1066 (O_1066,N_9930,N_9956);
or UO_1067 (O_1067,N_9929,N_9922);
and UO_1068 (O_1068,N_9932,N_9924);
xor UO_1069 (O_1069,N_9976,N_9912);
or UO_1070 (O_1070,N_9972,N_9971);
nand UO_1071 (O_1071,N_9986,N_9981);
nand UO_1072 (O_1072,N_9972,N_9939);
xor UO_1073 (O_1073,N_9961,N_9947);
or UO_1074 (O_1074,N_9954,N_9992);
nand UO_1075 (O_1075,N_9987,N_9931);
xnor UO_1076 (O_1076,N_9930,N_9974);
nor UO_1077 (O_1077,N_9926,N_9918);
nor UO_1078 (O_1078,N_9918,N_9976);
or UO_1079 (O_1079,N_9938,N_9996);
and UO_1080 (O_1080,N_9922,N_9946);
xnor UO_1081 (O_1081,N_9973,N_9949);
or UO_1082 (O_1082,N_9976,N_9924);
xnor UO_1083 (O_1083,N_9938,N_9910);
xnor UO_1084 (O_1084,N_9902,N_9993);
nand UO_1085 (O_1085,N_9981,N_9962);
nor UO_1086 (O_1086,N_9931,N_9925);
xnor UO_1087 (O_1087,N_9992,N_9993);
nor UO_1088 (O_1088,N_9905,N_9902);
or UO_1089 (O_1089,N_9965,N_9979);
or UO_1090 (O_1090,N_9967,N_9903);
nor UO_1091 (O_1091,N_9941,N_9938);
or UO_1092 (O_1092,N_9941,N_9981);
xnor UO_1093 (O_1093,N_9932,N_9920);
and UO_1094 (O_1094,N_9979,N_9993);
nand UO_1095 (O_1095,N_9939,N_9982);
or UO_1096 (O_1096,N_9935,N_9969);
xnor UO_1097 (O_1097,N_9951,N_9915);
nand UO_1098 (O_1098,N_9999,N_9967);
nand UO_1099 (O_1099,N_9986,N_9973);
or UO_1100 (O_1100,N_9959,N_9938);
and UO_1101 (O_1101,N_9913,N_9958);
xor UO_1102 (O_1102,N_9938,N_9925);
xnor UO_1103 (O_1103,N_9992,N_9989);
nor UO_1104 (O_1104,N_9918,N_9977);
xnor UO_1105 (O_1105,N_9907,N_9903);
xnor UO_1106 (O_1106,N_9922,N_9955);
nor UO_1107 (O_1107,N_9902,N_9982);
or UO_1108 (O_1108,N_9932,N_9982);
or UO_1109 (O_1109,N_9902,N_9956);
nor UO_1110 (O_1110,N_9900,N_9989);
nand UO_1111 (O_1111,N_9942,N_9953);
or UO_1112 (O_1112,N_9929,N_9987);
nor UO_1113 (O_1113,N_9973,N_9942);
xor UO_1114 (O_1114,N_9941,N_9960);
nand UO_1115 (O_1115,N_9961,N_9975);
or UO_1116 (O_1116,N_9958,N_9928);
or UO_1117 (O_1117,N_9946,N_9908);
and UO_1118 (O_1118,N_9955,N_9931);
nor UO_1119 (O_1119,N_9948,N_9906);
xor UO_1120 (O_1120,N_9985,N_9906);
nand UO_1121 (O_1121,N_9967,N_9902);
or UO_1122 (O_1122,N_9964,N_9947);
and UO_1123 (O_1123,N_9909,N_9956);
nand UO_1124 (O_1124,N_9941,N_9973);
and UO_1125 (O_1125,N_9949,N_9961);
nand UO_1126 (O_1126,N_9933,N_9935);
nor UO_1127 (O_1127,N_9968,N_9912);
and UO_1128 (O_1128,N_9941,N_9947);
or UO_1129 (O_1129,N_9952,N_9977);
or UO_1130 (O_1130,N_9952,N_9935);
nand UO_1131 (O_1131,N_9924,N_9904);
and UO_1132 (O_1132,N_9970,N_9926);
nor UO_1133 (O_1133,N_9976,N_9946);
nor UO_1134 (O_1134,N_9987,N_9924);
xnor UO_1135 (O_1135,N_9979,N_9964);
nor UO_1136 (O_1136,N_9968,N_9954);
and UO_1137 (O_1137,N_9940,N_9935);
xor UO_1138 (O_1138,N_9935,N_9955);
nor UO_1139 (O_1139,N_9935,N_9913);
or UO_1140 (O_1140,N_9937,N_9916);
nor UO_1141 (O_1141,N_9981,N_9991);
xor UO_1142 (O_1142,N_9979,N_9905);
nand UO_1143 (O_1143,N_9916,N_9963);
nand UO_1144 (O_1144,N_9944,N_9938);
nand UO_1145 (O_1145,N_9916,N_9934);
or UO_1146 (O_1146,N_9990,N_9963);
and UO_1147 (O_1147,N_9965,N_9963);
or UO_1148 (O_1148,N_9925,N_9960);
xnor UO_1149 (O_1149,N_9988,N_9925);
and UO_1150 (O_1150,N_9954,N_9914);
and UO_1151 (O_1151,N_9996,N_9902);
nor UO_1152 (O_1152,N_9929,N_9960);
nor UO_1153 (O_1153,N_9909,N_9922);
nand UO_1154 (O_1154,N_9940,N_9989);
nand UO_1155 (O_1155,N_9936,N_9901);
or UO_1156 (O_1156,N_9910,N_9919);
and UO_1157 (O_1157,N_9989,N_9990);
nand UO_1158 (O_1158,N_9933,N_9960);
nor UO_1159 (O_1159,N_9977,N_9960);
nor UO_1160 (O_1160,N_9958,N_9992);
or UO_1161 (O_1161,N_9917,N_9958);
or UO_1162 (O_1162,N_9945,N_9920);
nand UO_1163 (O_1163,N_9997,N_9965);
and UO_1164 (O_1164,N_9900,N_9926);
xor UO_1165 (O_1165,N_9926,N_9967);
xnor UO_1166 (O_1166,N_9957,N_9980);
nor UO_1167 (O_1167,N_9962,N_9965);
nor UO_1168 (O_1168,N_9942,N_9969);
and UO_1169 (O_1169,N_9961,N_9970);
nor UO_1170 (O_1170,N_9958,N_9909);
nand UO_1171 (O_1171,N_9949,N_9962);
and UO_1172 (O_1172,N_9980,N_9952);
xor UO_1173 (O_1173,N_9982,N_9979);
and UO_1174 (O_1174,N_9970,N_9902);
nand UO_1175 (O_1175,N_9931,N_9959);
or UO_1176 (O_1176,N_9916,N_9961);
or UO_1177 (O_1177,N_9921,N_9972);
and UO_1178 (O_1178,N_9951,N_9967);
or UO_1179 (O_1179,N_9923,N_9987);
nor UO_1180 (O_1180,N_9984,N_9940);
nand UO_1181 (O_1181,N_9938,N_9980);
and UO_1182 (O_1182,N_9962,N_9948);
and UO_1183 (O_1183,N_9937,N_9995);
nand UO_1184 (O_1184,N_9997,N_9918);
nor UO_1185 (O_1185,N_9936,N_9951);
nor UO_1186 (O_1186,N_9939,N_9923);
or UO_1187 (O_1187,N_9916,N_9969);
nor UO_1188 (O_1188,N_9929,N_9968);
xnor UO_1189 (O_1189,N_9999,N_9962);
and UO_1190 (O_1190,N_9943,N_9956);
nor UO_1191 (O_1191,N_9927,N_9926);
and UO_1192 (O_1192,N_9965,N_9904);
nand UO_1193 (O_1193,N_9990,N_9997);
nand UO_1194 (O_1194,N_9987,N_9950);
and UO_1195 (O_1195,N_9932,N_9910);
xnor UO_1196 (O_1196,N_9953,N_9975);
and UO_1197 (O_1197,N_9952,N_9943);
and UO_1198 (O_1198,N_9987,N_9978);
or UO_1199 (O_1199,N_9961,N_9934);
or UO_1200 (O_1200,N_9924,N_9916);
nor UO_1201 (O_1201,N_9964,N_9912);
or UO_1202 (O_1202,N_9964,N_9922);
and UO_1203 (O_1203,N_9970,N_9934);
xnor UO_1204 (O_1204,N_9966,N_9958);
or UO_1205 (O_1205,N_9964,N_9962);
xor UO_1206 (O_1206,N_9906,N_9960);
and UO_1207 (O_1207,N_9954,N_9994);
or UO_1208 (O_1208,N_9945,N_9963);
or UO_1209 (O_1209,N_9920,N_9937);
nand UO_1210 (O_1210,N_9971,N_9983);
xnor UO_1211 (O_1211,N_9963,N_9976);
xor UO_1212 (O_1212,N_9909,N_9982);
or UO_1213 (O_1213,N_9960,N_9922);
or UO_1214 (O_1214,N_9928,N_9910);
nand UO_1215 (O_1215,N_9932,N_9990);
nand UO_1216 (O_1216,N_9972,N_9964);
or UO_1217 (O_1217,N_9951,N_9961);
xnor UO_1218 (O_1218,N_9915,N_9908);
or UO_1219 (O_1219,N_9990,N_9928);
nand UO_1220 (O_1220,N_9905,N_9961);
and UO_1221 (O_1221,N_9904,N_9946);
nor UO_1222 (O_1222,N_9986,N_9957);
or UO_1223 (O_1223,N_9969,N_9976);
xnor UO_1224 (O_1224,N_9947,N_9935);
nor UO_1225 (O_1225,N_9996,N_9970);
and UO_1226 (O_1226,N_9938,N_9953);
or UO_1227 (O_1227,N_9995,N_9942);
nand UO_1228 (O_1228,N_9974,N_9962);
nor UO_1229 (O_1229,N_9994,N_9980);
xor UO_1230 (O_1230,N_9907,N_9931);
or UO_1231 (O_1231,N_9939,N_9934);
nor UO_1232 (O_1232,N_9976,N_9974);
nand UO_1233 (O_1233,N_9926,N_9995);
nor UO_1234 (O_1234,N_9994,N_9975);
or UO_1235 (O_1235,N_9910,N_9954);
nor UO_1236 (O_1236,N_9913,N_9933);
nand UO_1237 (O_1237,N_9976,N_9954);
nor UO_1238 (O_1238,N_9957,N_9981);
and UO_1239 (O_1239,N_9905,N_9927);
xor UO_1240 (O_1240,N_9949,N_9954);
xnor UO_1241 (O_1241,N_9996,N_9914);
xor UO_1242 (O_1242,N_9995,N_9971);
or UO_1243 (O_1243,N_9960,N_9939);
and UO_1244 (O_1244,N_9934,N_9947);
nor UO_1245 (O_1245,N_9973,N_9932);
nor UO_1246 (O_1246,N_9945,N_9933);
nand UO_1247 (O_1247,N_9988,N_9944);
and UO_1248 (O_1248,N_9959,N_9916);
nand UO_1249 (O_1249,N_9995,N_9955);
and UO_1250 (O_1250,N_9926,N_9924);
nand UO_1251 (O_1251,N_9972,N_9910);
or UO_1252 (O_1252,N_9960,N_9994);
or UO_1253 (O_1253,N_9933,N_9922);
or UO_1254 (O_1254,N_9913,N_9994);
or UO_1255 (O_1255,N_9996,N_9911);
nand UO_1256 (O_1256,N_9981,N_9947);
and UO_1257 (O_1257,N_9922,N_9900);
xnor UO_1258 (O_1258,N_9947,N_9979);
or UO_1259 (O_1259,N_9914,N_9906);
or UO_1260 (O_1260,N_9912,N_9975);
or UO_1261 (O_1261,N_9915,N_9929);
or UO_1262 (O_1262,N_9992,N_9928);
xnor UO_1263 (O_1263,N_9949,N_9955);
nor UO_1264 (O_1264,N_9973,N_9947);
and UO_1265 (O_1265,N_9917,N_9903);
nand UO_1266 (O_1266,N_9989,N_9991);
nand UO_1267 (O_1267,N_9973,N_9982);
xor UO_1268 (O_1268,N_9969,N_9934);
xnor UO_1269 (O_1269,N_9964,N_9969);
and UO_1270 (O_1270,N_9911,N_9993);
and UO_1271 (O_1271,N_9940,N_9931);
nor UO_1272 (O_1272,N_9939,N_9963);
xnor UO_1273 (O_1273,N_9929,N_9959);
and UO_1274 (O_1274,N_9958,N_9994);
and UO_1275 (O_1275,N_9951,N_9911);
or UO_1276 (O_1276,N_9940,N_9998);
nand UO_1277 (O_1277,N_9977,N_9900);
xor UO_1278 (O_1278,N_9935,N_9904);
xnor UO_1279 (O_1279,N_9940,N_9963);
or UO_1280 (O_1280,N_9962,N_9905);
or UO_1281 (O_1281,N_9962,N_9956);
and UO_1282 (O_1282,N_9965,N_9901);
nor UO_1283 (O_1283,N_9943,N_9916);
nor UO_1284 (O_1284,N_9910,N_9934);
xnor UO_1285 (O_1285,N_9919,N_9950);
nor UO_1286 (O_1286,N_9985,N_9994);
nand UO_1287 (O_1287,N_9939,N_9987);
nand UO_1288 (O_1288,N_9959,N_9996);
or UO_1289 (O_1289,N_9996,N_9929);
nor UO_1290 (O_1290,N_9976,N_9984);
xnor UO_1291 (O_1291,N_9934,N_9993);
nand UO_1292 (O_1292,N_9946,N_9919);
nor UO_1293 (O_1293,N_9979,N_9955);
xnor UO_1294 (O_1294,N_9972,N_9983);
xnor UO_1295 (O_1295,N_9911,N_9982);
or UO_1296 (O_1296,N_9926,N_9912);
and UO_1297 (O_1297,N_9901,N_9947);
nand UO_1298 (O_1298,N_9982,N_9990);
nor UO_1299 (O_1299,N_9964,N_9902);
and UO_1300 (O_1300,N_9945,N_9918);
and UO_1301 (O_1301,N_9908,N_9940);
or UO_1302 (O_1302,N_9900,N_9960);
xnor UO_1303 (O_1303,N_9970,N_9933);
or UO_1304 (O_1304,N_9958,N_9939);
xnor UO_1305 (O_1305,N_9964,N_9910);
nand UO_1306 (O_1306,N_9993,N_9984);
and UO_1307 (O_1307,N_9917,N_9911);
nor UO_1308 (O_1308,N_9955,N_9960);
and UO_1309 (O_1309,N_9939,N_9952);
or UO_1310 (O_1310,N_9983,N_9951);
or UO_1311 (O_1311,N_9957,N_9928);
xor UO_1312 (O_1312,N_9915,N_9948);
nor UO_1313 (O_1313,N_9937,N_9932);
nor UO_1314 (O_1314,N_9948,N_9930);
xnor UO_1315 (O_1315,N_9941,N_9909);
nand UO_1316 (O_1316,N_9920,N_9955);
or UO_1317 (O_1317,N_9999,N_9981);
or UO_1318 (O_1318,N_9923,N_9931);
nor UO_1319 (O_1319,N_9993,N_9945);
and UO_1320 (O_1320,N_9953,N_9932);
xnor UO_1321 (O_1321,N_9975,N_9918);
and UO_1322 (O_1322,N_9926,N_9993);
nand UO_1323 (O_1323,N_9976,N_9941);
or UO_1324 (O_1324,N_9950,N_9964);
and UO_1325 (O_1325,N_9971,N_9959);
or UO_1326 (O_1326,N_9900,N_9943);
or UO_1327 (O_1327,N_9998,N_9987);
nor UO_1328 (O_1328,N_9997,N_9983);
nand UO_1329 (O_1329,N_9952,N_9948);
or UO_1330 (O_1330,N_9978,N_9931);
nor UO_1331 (O_1331,N_9935,N_9975);
nor UO_1332 (O_1332,N_9962,N_9932);
and UO_1333 (O_1333,N_9992,N_9912);
or UO_1334 (O_1334,N_9957,N_9906);
nand UO_1335 (O_1335,N_9927,N_9931);
and UO_1336 (O_1336,N_9918,N_9938);
and UO_1337 (O_1337,N_9992,N_9923);
xor UO_1338 (O_1338,N_9911,N_9937);
xnor UO_1339 (O_1339,N_9982,N_9945);
or UO_1340 (O_1340,N_9939,N_9974);
or UO_1341 (O_1341,N_9932,N_9970);
nor UO_1342 (O_1342,N_9998,N_9959);
or UO_1343 (O_1343,N_9943,N_9968);
nand UO_1344 (O_1344,N_9924,N_9901);
xor UO_1345 (O_1345,N_9932,N_9938);
nor UO_1346 (O_1346,N_9931,N_9914);
and UO_1347 (O_1347,N_9974,N_9977);
nand UO_1348 (O_1348,N_9988,N_9999);
and UO_1349 (O_1349,N_9907,N_9981);
xnor UO_1350 (O_1350,N_9913,N_9950);
and UO_1351 (O_1351,N_9918,N_9995);
or UO_1352 (O_1352,N_9924,N_9989);
or UO_1353 (O_1353,N_9931,N_9963);
xnor UO_1354 (O_1354,N_9982,N_9994);
and UO_1355 (O_1355,N_9993,N_9923);
nor UO_1356 (O_1356,N_9938,N_9930);
nor UO_1357 (O_1357,N_9910,N_9907);
nand UO_1358 (O_1358,N_9903,N_9982);
nand UO_1359 (O_1359,N_9961,N_9918);
xnor UO_1360 (O_1360,N_9970,N_9987);
nor UO_1361 (O_1361,N_9918,N_9922);
xnor UO_1362 (O_1362,N_9982,N_9930);
xnor UO_1363 (O_1363,N_9921,N_9939);
nand UO_1364 (O_1364,N_9982,N_9907);
and UO_1365 (O_1365,N_9941,N_9911);
xnor UO_1366 (O_1366,N_9911,N_9974);
and UO_1367 (O_1367,N_9984,N_9901);
xnor UO_1368 (O_1368,N_9954,N_9985);
nor UO_1369 (O_1369,N_9961,N_9915);
xor UO_1370 (O_1370,N_9989,N_9902);
nor UO_1371 (O_1371,N_9991,N_9947);
xnor UO_1372 (O_1372,N_9989,N_9999);
nor UO_1373 (O_1373,N_9963,N_9981);
nor UO_1374 (O_1374,N_9905,N_9920);
and UO_1375 (O_1375,N_9998,N_9932);
nand UO_1376 (O_1376,N_9985,N_9947);
or UO_1377 (O_1377,N_9922,N_9971);
nor UO_1378 (O_1378,N_9961,N_9932);
nand UO_1379 (O_1379,N_9963,N_9997);
xor UO_1380 (O_1380,N_9986,N_9900);
nor UO_1381 (O_1381,N_9956,N_9932);
nand UO_1382 (O_1382,N_9917,N_9920);
and UO_1383 (O_1383,N_9928,N_9950);
or UO_1384 (O_1384,N_9965,N_9916);
nand UO_1385 (O_1385,N_9935,N_9918);
or UO_1386 (O_1386,N_9952,N_9900);
nand UO_1387 (O_1387,N_9972,N_9958);
and UO_1388 (O_1388,N_9996,N_9907);
nor UO_1389 (O_1389,N_9967,N_9913);
nand UO_1390 (O_1390,N_9907,N_9936);
nor UO_1391 (O_1391,N_9922,N_9976);
or UO_1392 (O_1392,N_9968,N_9915);
nor UO_1393 (O_1393,N_9938,N_9989);
nor UO_1394 (O_1394,N_9923,N_9918);
or UO_1395 (O_1395,N_9926,N_9989);
nor UO_1396 (O_1396,N_9900,N_9904);
xor UO_1397 (O_1397,N_9914,N_9982);
nand UO_1398 (O_1398,N_9926,N_9978);
xor UO_1399 (O_1399,N_9996,N_9909);
nor UO_1400 (O_1400,N_9912,N_9995);
and UO_1401 (O_1401,N_9930,N_9955);
nor UO_1402 (O_1402,N_9998,N_9921);
or UO_1403 (O_1403,N_9996,N_9923);
xor UO_1404 (O_1404,N_9978,N_9930);
xnor UO_1405 (O_1405,N_9991,N_9983);
nand UO_1406 (O_1406,N_9948,N_9973);
nand UO_1407 (O_1407,N_9918,N_9919);
nand UO_1408 (O_1408,N_9965,N_9919);
nor UO_1409 (O_1409,N_9960,N_9936);
xnor UO_1410 (O_1410,N_9967,N_9989);
xor UO_1411 (O_1411,N_9950,N_9918);
and UO_1412 (O_1412,N_9927,N_9985);
nor UO_1413 (O_1413,N_9953,N_9943);
or UO_1414 (O_1414,N_9942,N_9931);
and UO_1415 (O_1415,N_9965,N_9922);
and UO_1416 (O_1416,N_9975,N_9944);
or UO_1417 (O_1417,N_9975,N_9928);
nor UO_1418 (O_1418,N_9967,N_9990);
xnor UO_1419 (O_1419,N_9985,N_9990);
xor UO_1420 (O_1420,N_9969,N_9911);
and UO_1421 (O_1421,N_9946,N_9992);
xor UO_1422 (O_1422,N_9984,N_9906);
xor UO_1423 (O_1423,N_9916,N_9954);
or UO_1424 (O_1424,N_9937,N_9931);
xnor UO_1425 (O_1425,N_9953,N_9947);
and UO_1426 (O_1426,N_9942,N_9907);
and UO_1427 (O_1427,N_9942,N_9999);
nand UO_1428 (O_1428,N_9901,N_9900);
nand UO_1429 (O_1429,N_9980,N_9922);
xnor UO_1430 (O_1430,N_9971,N_9969);
xnor UO_1431 (O_1431,N_9987,N_9914);
nor UO_1432 (O_1432,N_9957,N_9949);
nand UO_1433 (O_1433,N_9942,N_9914);
or UO_1434 (O_1434,N_9949,N_9997);
and UO_1435 (O_1435,N_9962,N_9994);
nor UO_1436 (O_1436,N_9960,N_9931);
or UO_1437 (O_1437,N_9992,N_9938);
or UO_1438 (O_1438,N_9934,N_9978);
or UO_1439 (O_1439,N_9907,N_9934);
and UO_1440 (O_1440,N_9941,N_9980);
or UO_1441 (O_1441,N_9990,N_9958);
xnor UO_1442 (O_1442,N_9984,N_9952);
and UO_1443 (O_1443,N_9972,N_9973);
xnor UO_1444 (O_1444,N_9902,N_9917);
xnor UO_1445 (O_1445,N_9964,N_9986);
xnor UO_1446 (O_1446,N_9931,N_9958);
and UO_1447 (O_1447,N_9922,N_9928);
nand UO_1448 (O_1448,N_9975,N_9915);
or UO_1449 (O_1449,N_9912,N_9939);
nor UO_1450 (O_1450,N_9946,N_9977);
or UO_1451 (O_1451,N_9955,N_9916);
and UO_1452 (O_1452,N_9968,N_9923);
nand UO_1453 (O_1453,N_9911,N_9975);
nand UO_1454 (O_1454,N_9911,N_9983);
nor UO_1455 (O_1455,N_9953,N_9915);
nand UO_1456 (O_1456,N_9905,N_9946);
xor UO_1457 (O_1457,N_9931,N_9951);
and UO_1458 (O_1458,N_9977,N_9998);
xnor UO_1459 (O_1459,N_9906,N_9973);
or UO_1460 (O_1460,N_9956,N_9967);
xor UO_1461 (O_1461,N_9984,N_9958);
nor UO_1462 (O_1462,N_9947,N_9944);
nor UO_1463 (O_1463,N_9946,N_9959);
and UO_1464 (O_1464,N_9910,N_9943);
nand UO_1465 (O_1465,N_9914,N_9916);
and UO_1466 (O_1466,N_9927,N_9916);
nor UO_1467 (O_1467,N_9935,N_9960);
nand UO_1468 (O_1468,N_9920,N_9912);
or UO_1469 (O_1469,N_9949,N_9917);
or UO_1470 (O_1470,N_9912,N_9950);
xor UO_1471 (O_1471,N_9956,N_9964);
xor UO_1472 (O_1472,N_9918,N_9937);
or UO_1473 (O_1473,N_9959,N_9921);
nor UO_1474 (O_1474,N_9943,N_9937);
and UO_1475 (O_1475,N_9995,N_9959);
and UO_1476 (O_1476,N_9905,N_9980);
and UO_1477 (O_1477,N_9911,N_9948);
nand UO_1478 (O_1478,N_9936,N_9919);
and UO_1479 (O_1479,N_9982,N_9985);
and UO_1480 (O_1480,N_9988,N_9905);
xor UO_1481 (O_1481,N_9982,N_9920);
nor UO_1482 (O_1482,N_9994,N_9934);
and UO_1483 (O_1483,N_9978,N_9966);
or UO_1484 (O_1484,N_9986,N_9979);
nor UO_1485 (O_1485,N_9931,N_9985);
nand UO_1486 (O_1486,N_9917,N_9964);
and UO_1487 (O_1487,N_9955,N_9939);
xnor UO_1488 (O_1488,N_9930,N_9989);
or UO_1489 (O_1489,N_9910,N_9982);
nor UO_1490 (O_1490,N_9905,N_9966);
nor UO_1491 (O_1491,N_9968,N_9930);
xor UO_1492 (O_1492,N_9965,N_9954);
nor UO_1493 (O_1493,N_9915,N_9976);
nand UO_1494 (O_1494,N_9919,N_9915);
or UO_1495 (O_1495,N_9914,N_9956);
nand UO_1496 (O_1496,N_9959,N_9906);
nor UO_1497 (O_1497,N_9999,N_9939);
nand UO_1498 (O_1498,N_9976,N_9970);
nor UO_1499 (O_1499,N_9901,N_9962);
endmodule